* File: sky130_fd_sc_hdll__xnor2_2.pxi.spice
* Created: Wed Sep  2 08:53:44 2020
* 
x_PM_SKY130_FD_SC_HDLL__XNOR2_2%B N_B_c_95_n N_B_M1007_g N_B_c_102_n N_B_M1005_g
+ N_B_c_103_n N_B_M1016_g N_B_c_96_n N_B_M1017_g N_B_c_97_n N_B_M1004_g
+ N_B_c_104_n N_B_M1015_g N_B_c_105_n N_B_M1019_g N_B_c_98_n N_B_M1014_g
+ N_B_c_128_p N_B_c_106_n N_B_c_107_n N_B_c_124_p N_B_c_99_n N_B_c_108_n
+ N_B_c_109_n B N_B_c_100_n N_B_c_101_n B PM_SKY130_FD_SC_HDLL__XNOR2_2%B
x_PM_SKY130_FD_SC_HDLL__XNOR2_2%A N_A_c_211_n N_A_M1002_g N_A_c_218_n
+ N_A_M1009_g N_A_c_212_n N_A_M1003_g N_A_c_219_n N_A_M1012_g N_A_c_213_n
+ N_A_M1011_g N_A_c_220_n N_A_M1000_g N_A_c_221_n N_A_M1006_g N_A_c_214_n
+ N_A_M1018_g N_A_c_215_n N_A_c_216_n A N_A_c_217_n N_A_c_245_n
+ PM_SKY130_FD_SC_HDLL__XNOR2_2%A
x_PM_SKY130_FD_SC_HDLL__XNOR2_2%A_27_297# N_A_27_297#_M1007_s
+ N_A_27_297#_M1005_s N_A_27_297#_M1016_s N_A_27_297#_M1012_d
+ N_A_27_297#_c_304_n N_A_27_297#_M1001_g N_A_27_297#_c_313_n
+ N_A_27_297#_M1008_g N_A_27_297#_c_314_n N_A_27_297#_M1010_g
+ N_A_27_297#_c_305_n N_A_27_297#_M1013_g N_A_27_297#_c_306_n
+ N_A_27_297#_c_307_n N_A_27_297#_c_308_n N_A_27_297#_c_332_n
+ N_A_27_297#_c_338_n N_A_27_297#_c_316_n N_A_27_297#_c_357_n
+ N_A_27_297#_c_317_n N_A_27_297#_c_318_n N_A_27_297#_c_309_n
+ N_A_27_297#_c_310_n N_A_27_297#_c_311_n N_A_27_297#_c_320_n
+ N_A_27_297#_c_350_n N_A_27_297#_c_351_n N_A_27_297#_c_312_n
+ PM_SKY130_FD_SC_HDLL__XNOR2_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__XNOR2_2%VPWR N_VPWR_M1005_d N_VPWR_M1009_s
+ N_VPWR_M1000_s N_VPWR_M1008_d N_VPWR_M1010_d N_VPWR_c_445_n N_VPWR_c_446_n
+ N_VPWR_c_447_n N_VPWR_c_448_n N_VPWR_c_449_n N_VPWR_c_450_n N_VPWR_c_451_n
+ N_VPWR_c_452_n N_VPWR_c_453_n N_VPWR_c_454_n N_VPWR_c_455_n VPWR
+ N_VPWR_c_456_n N_VPWR_c_457_n N_VPWR_c_458_n N_VPWR_c_444_n
+ PM_SKY130_FD_SC_HDLL__XNOR2_2%VPWR
x_PM_SKY130_FD_SC_HDLL__XNOR2_2%A_514_297# N_A_514_297#_M1000_d
+ N_A_514_297#_M1006_d N_A_514_297#_M1019_s N_A_514_297#_c_550_n
+ N_A_514_297#_c_580_n N_A_514_297#_c_556_n N_A_514_297#_c_558_n
+ N_A_514_297#_c_569_n N_A_514_297#_c_552_n N_A_514_297#_c_554_n
+ PM_SKY130_FD_SC_HDLL__XNOR2_2%A_514_297#
x_PM_SKY130_FD_SC_HDLL__XNOR2_2%Y N_Y_M1001_d N_Y_M1013_d N_Y_M1015_d
+ N_Y_M1008_s N_Y_c_608_n N_Y_c_605_n N_Y_c_637_n N_Y_c_606_n N_Y_c_607_n
+ N_Y_c_623_n Y PM_SKY130_FD_SC_HDLL__XNOR2_2%Y
x_PM_SKY130_FD_SC_HDLL__XNOR2_2%A_27_47# N_A_27_47#_M1007_d N_A_27_47#_M1017_d
+ N_A_27_47#_M1003_d N_A_27_47#_c_660_n N_A_27_47#_c_669_n N_A_27_47#_c_661_n
+ N_A_27_47#_c_662_n N_A_27_47#_c_663_n PM_SKY130_FD_SC_HDLL__XNOR2_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__XNOR2_2%VGND N_VGND_M1002_s N_VGND_M1011_d
+ N_VGND_M1018_d N_VGND_M1014_d N_VGND_c_704_n N_VGND_c_705_n N_VGND_c_706_n
+ N_VGND_c_707_n N_VGND_c_708_n N_VGND_c_709_n N_VGND_c_710_n N_VGND_c_711_n
+ N_VGND_c_712_n N_VGND_c_713_n VGND N_VGND_c_714_n N_VGND_c_715_n
+ N_VGND_c_716_n N_VGND_c_717_n PM_SKY130_FD_SC_HDLL__XNOR2_2%VGND
x_PM_SKY130_FD_SC_HDLL__XNOR2_2%A_600_47# N_A_600_47#_M1011_s
+ N_A_600_47#_M1004_s N_A_600_47#_M1001_s N_A_600_47#_c_808_n
+ N_A_600_47#_c_794_n N_A_600_47#_c_795_n N_A_600_47#_c_803_n
+ N_A_600_47#_c_796_n N_A_600_47#_c_797_n N_A_600_47#_c_798_n
+ PM_SKY130_FD_SC_HDLL__XNOR2_2%A_600_47#
cc_1 VNB N_B_c_95_n 0.0200643f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_2 VNB N_B_c_96_n 0.0171406f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=0.995
cc_3 VNB N_B_c_97_n 0.0172187f $X=-0.19 $Y=-0.24 $X2=3.865 $Y2=0.995
cc_4 VNB N_B_c_98_n 0.0226999f $X=-0.19 $Y=-0.24 $X2=4.42 $Y2=0.995
cc_5 VNB N_B_c_99_n 0.00545644f $X=-0.19 $Y=-0.24 $X2=4.105 $Y2=1.16
cc_6 VNB N_B_c_100_n 0.0403029f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=1.202
cc_7 VNB N_B_c_101_n 0.0453222f $X=-0.19 $Y=-0.24 $X2=4.395 $Y2=1.202
cc_8 VNB N_A_c_211_n 0.0164927f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_9 VNB N_A_c_212_n 0.0219568f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=1.41
cc_10 VNB N_A_c_213_n 0.0222857f $X=-0.19 $Y=-0.24 $X2=3.865 $Y2=0.995
cc_11 VNB N_A_c_214_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=4.42 $Y2=0.995
cc_12 VNB N_A_c_215_n 0.0521692f $X=-0.19 $Y=-0.24 $X2=0.84 $Y2=1.18
cc_13 VNB N_A_c_216_n 0.0311503f $X=-0.19 $Y=-0.24 $X2=0.7 $Y2=1.16
cc_14 VNB N_A_c_217_n 0.031367f $X=-0.19 $Y=-0.24 $X2=3.265 $Y2=1.285
cc_15 VNB N_A_27_297#_c_304_n 0.022408f $X=-0.19 $Y=-0.24 $X2=3.865 $Y2=0.995
cc_16 VNB N_A_27_297#_c_305_n 0.0208584f $X=-0.19 $Y=-0.24 $X2=4.42 $Y2=0.995
cc_17 VNB N_A_27_297#_c_306_n 0.0205172f $X=-0.19 $Y=-0.24 $X2=0.7 $Y2=1.18
cc_18 VNB N_A_27_297#_c_307_n 0.0112022f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_297#_c_308_n 0.00613798f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=1.445
cc_20 VNB N_A_27_297#_c_309_n 0.0014749f $X=-0.19 $Y=-0.24 $X2=3.865 $Y2=1.202
cc_21 VNB N_A_27_297#_c_310_n 0.00469016f $X=-0.19 $Y=-0.24 $X2=3.89 $Y2=1.202
cc_22 VNB N_A_27_297#_c_311_n 0.00192645f $X=-0.19 $Y=-0.24 $X2=4.395 $Y2=1.202
cc_23 VNB N_A_27_297#_c_312_n 0.0460527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_444_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_Y_c_605_n 0.00241737f $X=-0.19 $Y=-0.24 $X2=3.865 $Y2=0.56
cc_26 VNB N_Y_c_606_n 0.00870355f $X=-0.19 $Y=-0.24 $X2=4.395 $Y2=1.985
cc_27 VNB N_Y_c_607_n 0.0365788f $X=-0.19 $Y=-0.24 $X2=4.42 $Y2=0.995
cc_28 VNB N_A_27_47#_c_660_n 0.00961138f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=0.995
cc_29 VNB N_A_27_47#_c_661_n 0.00359399f $X=-0.19 $Y=-0.24 $X2=3.865 $Y2=0.56
cc_30 VNB N_A_27_47#_c_662_n 0.00668696f $X=-0.19 $Y=-0.24 $X2=3.89 $Y2=1.41
cc_31 VNB N_A_27_47#_c_663_n 0.00473791f $X=-0.19 $Y=-0.24 $X2=4.395 $Y2=1.985
cc_32 VNB N_VGND_c_704_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=3.865 $Y2=0.56
cc_33 VNB N_VGND_c_705_n 0.0061705f $X=-0.19 $Y=-0.24 $X2=4.395 $Y2=1.41
cc_34 VNB N_VGND_c_706_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=4.42 $Y2=0.56
cc_35 VNB N_VGND_c_707_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0.7 $Y2=1.16
cc_36 VNB N_VGND_c_708_n 0.022981f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=1.285
cc_37 VNB N_VGND_c_709_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=1.445
cc_38 VNB N_VGND_c_710_n 0.0199314f $X=-0.19 $Y=-0.24 $X2=3.265 $Y2=1.445
cc_39 VNB N_VGND_c_711_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=3.35 $Y2=1.18
cc_40 VNB N_VGND_c_712_n 0.0200753f $X=-0.19 $Y=-0.24 $X2=4.105 $Y2=1.16
cc_41 VNB N_VGND_c_713_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=4.105 $Y2=1.16
cc_42 VNB N_VGND_c_714_n 0.0397774f $X=-0.19 $Y=-0.24 $X2=3.18 $Y2=1.53
cc_43 VNB N_VGND_c_715_n 0.0444932f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_716_n 0.329131f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_717_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_600_47#_c_794_n 0.00265754f $X=-0.19 $Y=-0.24 $X2=3.865 $Y2=0.56
cc_47 VNB N_A_600_47#_c_795_n 0.00345369f $X=-0.19 $Y=-0.24 $X2=3.865 $Y2=0.56
cc_48 VNB N_A_600_47#_c_796_n 0.00296989f $X=-0.19 $Y=-0.24 $X2=4.42 $Y2=0.995
cc_49 VNB N_A_600_47#_c_797_n 0.00254255f $X=-0.19 $Y=-0.24 $X2=4.42 $Y2=0.56
cc_50 VNB N_A_600_47#_c_798_n 0.016375f $X=-0.19 $Y=-0.24 $X2=0.84 $Y2=1.18
cc_51 VPB N_B_c_102_n 0.019152f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.41
cc_52 VPB N_B_c_103_n 0.0158458f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.41
cc_53 VPB N_B_c_104_n 0.0163836f $X=-0.19 $Y=1.305 $X2=3.89 $Y2=1.41
cc_54 VPB N_B_c_105_n 0.0197756f $X=-0.19 $Y=1.305 $X2=4.395 $Y2=1.41
cc_55 VPB N_B_c_106_n 0.00110906f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.445
cc_56 VPB N_B_c_107_n 0.00111619f $X=-0.19 $Y=1.305 $X2=3.265 $Y2=1.445
cc_57 VPB N_B_c_108_n 3.75749e-19 $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.53
cc_58 VPB N_B_c_109_n 0.0174163f $X=-0.19 $Y=1.305 $X2=3.18 $Y2=1.53
cc_59 VPB N_B_c_100_n 0.0211369f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.202
cc_60 VPB N_B_c_101_n 0.0218116f $X=-0.19 $Y=1.305 $X2=4.395 $Y2=1.202
cc_61 VPB N_A_c_218_n 0.0159819f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.41
cc_62 VPB N_A_c_219_n 0.0201091f $X=-0.19 $Y=1.305 $X2=1.005 $Y2=0.995
cc_63 VPB N_A_c_220_n 0.0200815f $X=-0.19 $Y=1.305 $X2=3.89 $Y2=1.41
cc_64 VPB N_A_c_221_n 0.0160958f $X=-0.19 $Y=1.305 $X2=4.395 $Y2=1.41
cc_65 VPB N_A_c_215_n 0.0215169f $X=-0.19 $Y=1.305 $X2=0.84 $Y2=1.18
cc_66 VPB N_A_c_216_n 0.0218747f $X=-0.19 $Y=1.305 $X2=0.7 $Y2=1.16
cc_67 VPB N_A_c_217_n 0.0216533f $X=-0.19 $Y=1.305 $X2=3.265 $Y2=1.285
cc_68 VPB N_A_27_297#_c_313_n 0.019044f $X=-0.19 $Y=1.305 $X2=3.89 $Y2=1.41
cc_69 VPB N_A_27_297#_c_314_n 0.0191634f $X=-0.19 $Y=1.305 $X2=4.395 $Y2=1.41
cc_70 VPB N_A_27_297#_c_306_n 0.0206721f $X=-0.19 $Y=1.305 $X2=0.7 $Y2=1.18
cc_71 VPB N_A_27_297#_c_316_n 0.0079379f $X=-0.19 $Y=1.305 $X2=1.06 $Y2=1.445
cc_72 VPB N_A_27_297#_c_317_n 0.0150054f $X=-0.19 $Y=1.305 $X2=0.7 $Y2=1.202
cc_73 VPB N_A_27_297#_c_318_n 0.00179402f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.202
cc_74 VPB N_A_27_297#_c_309_n 0.00375635f $X=-0.19 $Y=1.305 $X2=3.865 $Y2=1.202
cc_75 VPB N_A_27_297#_c_320_n 0.0274163f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.53
cc_76 VPB N_A_27_297#_c_312_n 0.0207963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_445_n 0.00516582f $X=-0.19 $Y=1.305 $X2=4.395 $Y2=1.985
cc_78 VPB N_VPWR_c_446_n 0.0180033f $X=-0.19 $Y=1.305 $X2=4.42 $Y2=0.995
cc_79 VPB N_VPWR_c_447_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0.7 $Y2=1.18
cc_80 VPB N_VPWR_c_448_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.285
cc_81 VPB N_VPWR_c_449_n 0.00518f $X=-0.19 $Y=1.305 $X2=3.35 $Y2=1.18
cc_82 VPB N_VPWR_c_450_n 0.012578f $X=-0.19 $Y=1.305 $X2=4.105 $Y2=1.16
cc_83 VPB N_VPWR_c_451_n 0.0355081f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_452_n 0.0342691f $X=-0.19 $Y=1.305 $X2=1.06 $Y2=1.445
cc_85 VPB N_VPWR_c_453_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_454_n 0.0417393f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.202
cc_87 VPB N_VPWR_c_455_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0.7 $Y2=1.202
cc_88 VPB N_VPWR_c_456_n 0.0199228f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_457_n 0.0229322f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_458_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_444_n 0.0514084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_Y_c_608_n 0.0081428f $X=-0.19 $Y=1.305 $X2=3.865 $Y2=0.995
cc_93 VPB N_Y_c_607_n 0.00617194f $X=-0.19 $Y=1.305 $X2=4.42 $Y2=0.995
cc_94 VPB Y 0.0139784f $X=-0.19 $Y=1.305 $X2=3.265 $Y2=1.285
cc_95 N_B_c_96_n N_A_c_211_n 0.0174641f $X=1.005 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_96 N_B_c_103_n N_A_c_218_n 0.0227815f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_97 N_B_c_109_n N_A_c_218_n 0.0118596f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_98 N_B_c_109_n N_A_c_219_n 0.0139024f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_99 N_B_c_107_n N_A_c_220_n 7.38573e-19 $X=3.265 $Y=1.445 $X2=0 $Y2=0
cc_100 N_B_c_109_n N_A_c_220_n 0.0167584f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_101 N_B_c_104_n N_A_c_221_n 0.0339574f $X=3.89 $Y=1.41 $X2=0 $Y2=0
cc_102 N_B_c_107_n N_A_c_221_n 8.28383e-19 $X=3.265 $Y=1.445 $X2=0 $Y2=0
cc_103 N_B_c_109_n N_A_c_221_n 0.00458999f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_104 N_B_c_97_n N_A_c_214_n 0.0240039f $X=3.865 $Y=0.995 $X2=0 $Y2=0
cc_105 N_B_c_109_n N_A_c_215_n 0.0202172f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_106 N_B_c_107_n N_A_c_216_n 0.00991248f $X=3.265 $Y=1.445 $X2=0 $Y2=0
cc_107 N_B_c_124_p N_A_c_216_n 0.00936469f $X=3.35 $Y=1.18 $X2=0 $Y2=0
cc_108 N_B_c_99_n N_A_c_216_n 0.0121981f $X=4.105 $Y=1.16 $X2=0 $Y2=0
cc_109 N_B_c_109_n N_A_c_216_n 0.00446101f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_110 N_B_c_101_n N_A_c_216_n 0.0240039f $X=4.395 $Y=1.202 $X2=0 $Y2=0
cc_111 N_B_c_128_p N_A_c_217_n 8.65006e-19 $X=0.84 $Y=1.18 $X2=0 $Y2=0
cc_112 N_B_c_106_n N_A_c_217_n 7.38579e-19 $X=0.925 $Y=1.445 $X2=0 $Y2=0
cc_113 N_B_c_109_n N_A_c_217_n 0.00822315f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_114 N_B_c_100_n N_A_c_217_n 0.0174641f $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_115 N_B_c_128_p N_A_c_245_n 0.00934672f $X=0.84 $Y=1.18 $X2=0 $Y2=0
cc_116 N_B_c_124_p N_A_c_245_n 0.0114522f $X=3.35 $Y=1.18 $X2=0 $Y2=0
cc_117 N_B_c_109_n N_A_c_245_n 0.111043f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_118 N_B_c_100_n N_A_c_245_n 8.98834e-19 $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_119 N_B_c_109_n N_A_27_297#_M1016_s 0.00187091f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_120 N_B_c_109_n N_A_27_297#_M1012_d 0.00326277f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_121 N_B_c_95_n N_A_27_297#_c_306_n 0.0171172f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_122 N_B_c_102_n N_A_27_297#_c_306_n 0.0115243f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_123 N_B_c_128_p N_A_27_297#_c_306_n 0.0166521f $X=0.84 $Y=1.18 $X2=0 $Y2=0
cc_124 N_B_c_106_n N_A_27_297#_c_306_n 0.00542123f $X=0.925 $Y=1.445 $X2=0 $Y2=0
cc_125 N_B_c_108_n N_A_27_297#_c_306_n 0.00367293f $X=1.01 $Y=1.53 $X2=0 $Y2=0
cc_126 N_B_c_95_n N_A_27_297#_c_308_n 0.01524f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_127 N_B_c_128_p N_A_27_297#_c_308_n 0.0305592f $X=0.84 $Y=1.18 $X2=0 $Y2=0
cc_128 N_B_c_100_n N_A_27_297#_c_308_n 0.00470019f $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_129 N_B_c_102_n N_A_27_297#_c_332_n 0.0155661f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_130 N_B_c_103_n N_A_27_297#_c_332_n 0.012299f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_131 N_B_c_128_p N_A_27_297#_c_332_n 0.00967248f $X=0.84 $Y=1.18 $X2=0 $Y2=0
cc_132 N_B_c_108_n N_A_27_297#_c_332_n 0.00896222f $X=1.01 $Y=1.53 $X2=0 $Y2=0
cc_133 N_B_c_109_n N_A_27_297#_c_332_n 0.00401671f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_134 N_B_c_100_n N_A_27_297#_c_332_n 0.00416568f $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_135 N_B_c_109_n N_A_27_297#_c_338_n 0.0372789f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_136 N_B_c_99_n N_A_27_297#_c_316_n 0.00704997f $X=4.105 $Y=1.16 $X2=0 $Y2=0
cc_137 N_B_c_109_n N_A_27_297#_c_316_n 0.0642896f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_138 N_B_c_104_n N_A_27_297#_c_317_n 0.0138603f $X=3.89 $Y=1.41 $X2=0 $Y2=0
cc_139 N_B_c_105_n N_A_27_297#_c_317_n 0.0162885f $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_140 N_B_c_99_n N_A_27_297#_c_317_n 0.0374638f $X=4.105 $Y=1.16 $X2=0 $Y2=0
cc_141 N_B_c_101_n N_A_27_297#_c_317_n 0.00876763f $X=4.395 $Y=1.202 $X2=0 $Y2=0
cc_142 N_B_c_99_n N_A_27_297#_c_318_n 0.0142097f $X=4.105 $Y=1.16 $X2=0 $Y2=0
cc_143 N_B_c_109_n N_A_27_297#_c_318_n 0.0101184f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_144 N_B_c_105_n N_A_27_297#_c_309_n 0.00103459f $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_145 N_B_c_101_n N_A_27_297#_c_309_n 0.00428171f $X=4.395 $Y=1.202 $X2=0 $Y2=0
cc_146 N_B_c_101_n N_A_27_297#_c_310_n 0.0055665f $X=4.395 $Y=1.202 $X2=0 $Y2=0
cc_147 N_B_c_109_n N_A_27_297#_c_350_n 0.0143191f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_148 N_B_c_109_n N_A_27_297#_c_351_n 0.0173294f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_149 N_B_c_109_n N_VPWR_M1009_s 0.00187547f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_150 N_B_c_109_n N_VPWR_M1000_s 0.00186066f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_151 N_B_c_102_n N_VPWR_c_445_n 0.00300743f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_152 N_B_c_103_n N_VPWR_c_445_n 0.00300743f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_153 N_B_c_103_n N_VPWR_c_446_n 0.0053025f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_154 N_B_c_105_n N_VPWR_c_449_n 0.00213395f $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_155 N_B_c_104_n N_VPWR_c_454_n 0.00430894f $X=3.89 $Y=1.41 $X2=0 $Y2=0
cc_156 N_B_c_105_n N_VPWR_c_454_n 0.00429453f $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_157 N_B_c_102_n N_VPWR_c_457_n 0.0053025f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_158 N_B_c_102_n N_VPWR_c_444_n 0.00783005f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_159 N_B_c_103_n N_VPWR_c_444_n 0.00693014f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_160 N_B_c_104_n N_VPWR_c_444_n 0.00573936f $X=3.89 $Y=1.41 $X2=0 $Y2=0
cc_161 N_B_c_105_n N_VPWR_c_444_n 0.00743743f $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_162 N_B_c_109_n N_A_514_297#_M1000_d 0.00321556f $X=3.18 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_163 N_B_c_104_n N_A_514_297#_c_550_n 0.00877428f $X=3.89 $Y=1.41 $X2=0 $Y2=0
cc_164 N_B_c_105_n N_A_514_297#_c_550_n 0.0101571f $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_165 N_B_c_104_n N_A_514_297#_c_552_n 0.00423898f $X=3.89 $Y=1.41 $X2=0 $Y2=0
cc_166 N_B_c_105_n N_A_514_297#_c_552_n 8.12765e-19 $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_167 N_B_c_104_n N_A_514_297#_c_554_n 0.0057248f $X=3.89 $Y=1.41 $X2=0 $Y2=0
cc_168 N_B_c_105_n N_A_514_297#_c_554_n 7.7891e-19 $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_169 N_B_c_105_n N_Y_c_608_n 0.0128257f $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_170 N_B_c_95_n N_A_27_47#_c_660_n 0.00964761f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_171 N_B_c_96_n N_A_27_47#_c_660_n 0.0129372f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B_c_128_p N_A_27_47#_c_660_n 0.00242422f $X=0.84 $Y=1.18 $X2=0 $Y2=0
cc_173 N_B_c_96_n N_A_27_47#_c_661_n 4.25198e-19 $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_174 N_B_c_109_n N_A_27_47#_c_661_n 0.00848395f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_175 N_B_c_97_n N_VGND_c_706_n 0.00268723f $X=3.865 $Y=0.995 $X2=0 $Y2=0
cc_176 N_B_c_98_n N_VGND_c_707_n 0.00438629f $X=4.42 $Y=0.995 $X2=0 $Y2=0
cc_177 N_B_c_97_n N_VGND_c_712_n 0.00423334f $X=3.865 $Y=0.995 $X2=0 $Y2=0
cc_178 N_B_c_98_n N_VGND_c_712_n 0.00437852f $X=4.42 $Y=0.995 $X2=0 $Y2=0
cc_179 N_B_c_95_n N_VGND_c_714_n 0.00357877f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_180 N_B_c_96_n N_VGND_c_714_n 0.00357877f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_181 N_B_c_95_n N_VGND_c_716_n 0.00644512f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_182 N_B_c_96_n N_VGND_c_716_n 0.005504f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_183 N_B_c_97_n N_VGND_c_716_n 0.00611128f $X=3.865 $Y=0.995 $X2=0 $Y2=0
cc_184 N_B_c_98_n N_VGND_c_716_n 0.00752949f $X=4.42 $Y=0.995 $X2=0 $Y2=0
cc_185 N_B_c_97_n N_A_600_47#_c_794_n 0.00865686f $X=3.865 $Y=0.995 $X2=0 $Y2=0
cc_186 N_B_c_99_n N_A_600_47#_c_794_n 0.0407882f $X=4.105 $Y=1.16 $X2=0 $Y2=0
cc_187 N_B_c_124_p N_A_600_47#_c_795_n 0.0148552f $X=3.35 $Y=1.18 $X2=0 $Y2=0
cc_188 N_B_c_109_n N_A_600_47#_c_795_n 0.00744432f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_189 N_B_c_97_n N_A_600_47#_c_803_n 0.013155f $X=3.865 $Y=0.995 $X2=0 $Y2=0
cc_190 N_B_c_97_n N_A_600_47#_c_796_n 0.00377905f $X=3.865 $Y=0.995 $X2=0 $Y2=0
cc_191 N_B_c_99_n N_A_600_47#_c_796_n 0.0320564f $X=4.105 $Y=1.16 $X2=0 $Y2=0
cc_192 N_B_c_101_n N_A_600_47#_c_796_n 0.00575847f $X=4.395 $Y=1.202 $X2=0 $Y2=0
cc_193 N_B_c_98_n N_A_600_47#_c_798_n 0.0147453f $X=4.42 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_c_218_n N_A_27_297#_c_338_n 0.0123176f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A_c_219_n N_A_27_297#_c_338_n 0.0123176f $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A_c_220_n N_A_27_297#_c_316_n 0.014186f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A_c_221_n N_A_27_297#_c_316_n 0.0136013f $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_c_216_n N_A_27_297#_c_316_n 5.77563e-19 $X=3.42 $Y=1.202 $X2=0 $Y2=0
cc_199 N_A_c_221_n N_A_27_297#_c_357_n 0.00361661f $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_200 N_A_c_221_n N_A_27_297#_c_318_n 0.00178809f $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A_c_220_n N_A_27_297#_c_351_n 0.00447768f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A_c_218_n N_VPWR_c_446_n 0.0053025f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A_c_218_n N_VPWR_c_447_n 0.00300743f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A_c_219_n N_VPWR_c_447_n 0.00300743f $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A_c_220_n N_VPWR_c_448_n 0.00324888f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A_c_221_n N_VPWR_c_448_n 0.00324888f $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A_c_219_n N_VPWR_c_452_n 0.0053025f $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A_c_220_n N_VPWR_c_452_n 0.00702461f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A_c_221_n N_VPWR_c_454_n 0.00702461f $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A_c_218_n N_VPWR_c_444_n 0.00693014f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A_c_219_n N_VPWR_c_444_n 0.00818727f $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A_c_220_n N_VPWR_c_444_n 0.00689121f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_213 N_A_c_221_n N_VPWR_c_444_n 0.0056586f $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A_c_220_n N_A_514_297#_c_556_n 0.00243733f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A_c_221_n N_A_514_297#_c_556_n 0.00300011f $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A_c_220_n N_A_514_297#_c_558_n 0.00176867f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_217 N_A_c_221_n N_A_514_297#_c_552_n 4.31774e-19 $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A_c_211_n N_A_27_47#_c_669_n 0.00282739f $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A_c_211_n N_A_27_47#_c_661_n 0.00513431f $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_c_212_n N_A_27_47#_c_661_n 4.74935e-19 $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A_c_245_n N_A_27_47#_c_661_n 0.00185207f $X=1.52 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A_c_211_n N_A_27_47#_c_662_n 0.00901254f $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A_c_212_n N_A_27_47#_c_662_n 0.010262f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A_c_215_n N_A_27_47#_c_662_n 0.00664936f $X=2.85 $Y=1.16 $X2=0 $Y2=0
cc_225 N_A_c_217_n N_A_27_47#_c_662_n 0.00345343f $X=2.02 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A_c_245_n N_A_27_47#_c_662_n 0.070814f $X=1.52 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A_c_211_n N_A_27_47#_c_663_n 5.24597e-19 $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A_c_212_n N_A_27_47#_c_663_n 0.00651696f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A_c_211_n N_VGND_c_704_n 0.00378935f $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A_c_212_n N_VGND_c_704_n 0.00276126f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A_c_212_n N_VGND_c_705_n 0.00274593f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_c_213_n N_VGND_c_705_n 0.00482457f $X=2.925 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_c_215_n N_VGND_c_705_n 0.00330968f $X=2.85 $Y=1.16 $X2=0 $Y2=0
cc_234 N_A_c_245_n N_VGND_c_705_n 0.0137693f $X=1.52 $Y=1.16 $X2=0 $Y2=0
cc_235 N_A_c_214_n N_VGND_c_706_n 0.00268723f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A_c_212_n N_VGND_c_708_n 0.00423334f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A_c_213_n N_VGND_c_710_n 0.00541359f $X=2.925 $Y=0.995 $X2=0 $Y2=0
cc_238 N_A_c_214_n N_VGND_c_710_n 0.00437852f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A_c_211_n N_VGND_c_714_n 0.00421816f $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A_c_211_n N_VGND_c_716_n 0.00600232f $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A_c_212_n N_VGND_c_716_n 0.00716934f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_c_213_n N_VGND_c_716_n 0.0110699f $X=2.925 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A_c_214_n N_VGND_c_716_n 0.00615622f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_c_213_n N_A_600_47#_c_808_n 0.00539651f $X=2.925 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A_c_214_n N_A_600_47#_c_794_n 0.0106151f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_c_213_n N_A_600_47#_c_795_n 0.00306677f $X=2.925 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A_c_216_n N_A_600_47#_c_795_n 0.00540411f $X=3.42 $Y=1.202 $X2=0 $Y2=0
cc_248 N_A_c_214_n N_A_600_47#_c_803_n 5.31699e-19 $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A_27_297#_c_332_n N_VPWR_M1005_d 0.0044785f $X=1.09 $Y=1.875 $X2=-0.19
+ $Y2=-0.24
cc_250 N_A_27_297#_c_338_n N_VPWR_M1009_s 0.00348321f $X=2.03 $Y=1.875 $X2=0
+ $Y2=0
cc_251 N_A_27_297#_c_316_n N_VPWR_M1000_s 0.00337791f $X=3.61 $Y=1.87 $X2=0
+ $Y2=0
cc_252 N_A_27_297#_c_317_n N_VPWR_M1008_d 0.0047706f $X=5.035 $Y=1.54 $X2=0
+ $Y2=0
cc_253 N_A_27_297#_c_332_n N_VPWR_c_445_n 0.0139299f $X=1.09 $Y=1.875 $X2=0
+ $Y2=0
cc_254 N_A_27_297#_c_332_n N_VPWR_c_446_n 0.00254499f $X=1.09 $Y=1.875 $X2=0
+ $Y2=0
cc_255 N_A_27_297#_c_338_n N_VPWR_c_446_n 0.00254499f $X=2.03 $Y=1.875 $X2=0
+ $Y2=0
cc_256 N_A_27_297#_c_350_n N_VPWR_c_446_n 0.0149311f $X=1.215 $Y=1.96 $X2=0
+ $Y2=0
cc_257 N_A_27_297#_c_338_n N_VPWR_c_447_n 0.0139299f $X=2.03 $Y=1.875 $X2=0
+ $Y2=0
cc_258 N_A_27_297#_c_316_n N_VPWR_c_448_n 0.0124746f $X=3.61 $Y=1.87 $X2=0 $Y2=0
cc_259 N_A_27_297#_c_313_n N_VPWR_c_449_n 0.00479105f $X=5.385 $Y=1.41 $X2=0
+ $Y2=0
cc_260 N_A_27_297#_c_314_n N_VPWR_c_451_n 0.00491766f $X=5.855 $Y=1.41 $X2=0
+ $Y2=0
cc_261 N_A_27_297#_c_338_n N_VPWR_c_452_n 0.00254499f $X=2.03 $Y=1.875 $X2=0
+ $Y2=0
cc_262 N_A_27_297#_c_351_n N_VPWR_c_452_n 0.0161853f $X=2.155 $Y=1.96 $X2=0
+ $Y2=0
cc_263 N_A_27_297#_c_313_n N_VPWR_c_456_n 0.0053025f $X=5.385 $Y=1.41 $X2=0
+ $Y2=0
cc_264 N_A_27_297#_c_314_n N_VPWR_c_456_n 0.00702461f $X=5.855 $Y=1.41 $X2=0
+ $Y2=0
cc_265 N_A_27_297#_c_332_n N_VPWR_c_457_n 0.00254499f $X=1.09 $Y=1.875 $X2=0
+ $Y2=0
cc_266 N_A_27_297#_c_320_n N_VPWR_c_457_n 0.0208235f $X=0.275 $Y=1.96 $X2=0
+ $Y2=0
cc_267 N_A_27_297#_M1005_s N_VPWR_c_444_n 0.00239308f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_268 N_A_27_297#_M1016_s N_VPWR_c_444_n 0.00250248f $X=1.07 $Y=1.485 $X2=0
+ $Y2=0
cc_269 N_A_27_297#_M1012_d N_VPWR_c_444_n 0.00253742f $X=2.01 $Y=1.485 $X2=0
+ $Y2=0
cc_270 N_A_27_297#_c_313_n N_VPWR_c_444_n 0.00823423f $X=5.385 $Y=1.41 $X2=0
+ $Y2=0
cc_271 N_A_27_297#_c_314_n N_VPWR_c_444_n 0.013472f $X=5.855 $Y=1.41 $X2=0 $Y2=0
cc_272 N_A_27_297#_c_332_n N_VPWR_c_444_n 0.0103134f $X=1.09 $Y=1.875 $X2=0
+ $Y2=0
cc_273 N_A_27_297#_c_338_n N_VPWR_c_444_n 0.0103134f $X=2.03 $Y=1.875 $X2=0
+ $Y2=0
cc_274 N_A_27_297#_c_316_n N_VPWR_c_444_n 0.0117978f $X=3.61 $Y=1.87 $X2=0 $Y2=0
cc_275 N_A_27_297#_c_320_n N_VPWR_c_444_n 0.0120542f $X=0.275 $Y=1.96 $X2=0
+ $Y2=0
cc_276 N_A_27_297#_c_350_n N_VPWR_c_444_n 0.00955092f $X=1.215 $Y=1.96 $X2=0
+ $Y2=0
cc_277 N_A_27_297#_c_351_n N_VPWR_c_444_n 0.00955092f $X=2.155 $Y=1.96 $X2=0
+ $Y2=0
cc_278 N_A_27_297#_c_316_n N_A_514_297#_M1000_d 0.00563848f $X=3.61 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_279 N_A_27_297#_c_316_n N_A_514_297#_M1006_d 0.00289412f $X=3.61 $Y=1.87
+ $X2=0 $Y2=0
cc_280 N_A_27_297#_c_357_n N_A_514_297#_M1006_d 0.00176276f $X=3.695 $Y=1.785
+ $X2=0 $Y2=0
cc_281 N_A_27_297#_c_318_n N_A_514_297#_M1006_d 0.00150347f $X=3.78 $Y=1.54
+ $X2=0 $Y2=0
cc_282 N_A_27_297#_c_317_n N_A_514_297#_M1019_s 0.00295153f $X=5.035 $Y=1.54
+ $X2=0 $Y2=0
cc_283 N_A_27_297#_c_317_n N_A_514_297#_c_550_n 0.00296639f $X=5.035 $Y=1.54
+ $X2=0 $Y2=0
cc_284 N_A_27_297#_c_316_n N_A_514_297#_c_556_n 0.0172782f $X=3.61 $Y=1.87 $X2=0
+ $Y2=0
cc_285 N_A_27_297#_c_316_n N_A_514_297#_c_558_n 0.00913267f $X=3.61 $Y=1.87
+ $X2=0 $Y2=0
cc_286 N_A_27_297#_c_351_n N_A_514_297#_c_558_n 0.00270019f $X=2.155 $Y=1.96
+ $X2=0 $Y2=0
cc_287 N_A_27_297#_c_316_n N_A_514_297#_c_569_n 0.0144404f $X=3.61 $Y=1.87 $X2=0
+ $Y2=0
cc_288 N_A_27_297#_c_351_n N_A_514_297#_c_569_n 0.0152341f $X=2.155 $Y=1.96
+ $X2=0 $Y2=0
cc_289 N_A_27_297#_c_316_n N_A_514_297#_c_552_n 0.0045174f $X=3.61 $Y=1.87 $X2=0
+ $Y2=0
cc_290 N_A_27_297#_c_317_n N_A_514_297#_c_552_n 0.00264455f $X=5.035 $Y=1.54
+ $X2=0 $Y2=0
cc_291 N_A_27_297#_c_316_n N_A_514_297#_c_554_n 0.0130614f $X=3.61 $Y=1.87 $X2=0
+ $Y2=0
cc_292 N_A_27_297#_c_317_n N_A_514_297#_c_554_n 9.8802e-19 $X=5.035 $Y=1.54
+ $X2=0 $Y2=0
cc_293 N_A_27_297#_c_317_n N_Y_M1015_d 0.00265147f $X=5.035 $Y=1.54 $X2=0 $Y2=0
cc_294 N_A_27_297#_c_313_n N_Y_c_608_n 0.0162359f $X=5.385 $Y=1.41 $X2=0 $Y2=0
cc_295 N_A_27_297#_c_317_n N_Y_c_608_n 0.0622533f $X=5.035 $Y=1.54 $X2=0 $Y2=0
cc_296 N_A_27_297#_c_311_n N_Y_c_608_n 0.00684602f $X=5.58 $Y=1.16 $X2=0 $Y2=0
cc_297 N_A_27_297#_c_304_n N_Y_c_605_n 0.00888424f $X=5.36 $Y=0.995 $X2=0 $Y2=0
cc_298 N_A_27_297#_c_305_n N_Y_c_605_n 0.012708f $X=5.88 $Y=0.995 $X2=0 $Y2=0
cc_299 N_A_27_297#_c_304_n N_Y_c_607_n 9.90894e-19 $X=5.36 $Y=0.995 $X2=0 $Y2=0
cc_300 N_A_27_297#_c_314_n N_Y_c_607_n 2.10127e-19 $X=5.855 $Y=1.41 $X2=0 $Y2=0
cc_301 N_A_27_297#_c_305_n N_Y_c_607_n 0.00955064f $X=5.88 $Y=0.995 $X2=0 $Y2=0
cc_302 N_A_27_297#_c_311_n N_Y_c_607_n 0.0117164f $X=5.58 $Y=1.16 $X2=0 $Y2=0
cc_303 N_A_27_297#_c_312_n N_Y_c_607_n 0.0211036f $X=5.855 $Y=1.202 $X2=0 $Y2=0
cc_304 N_A_27_297#_c_317_n N_Y_c_623_n 0.0132087f $X=5.035 $Y=1.54 $X2=0 $Y2=0
cc_305 N_A_27_297#_c_313_n Y 7.92403e-19 $X=5.385 $Y=1.41 $X2=0 $Y2=0
cc_306 N_A_27_297#_c_314_n Y 0.0249314f $X=5.855 $Y=1.41 $X2=0 $Y2=0
cc_307 N_A_27_297#_c_317_n Y 0.00610927f $X=5.035 $Y=1.54 $X2=0 $Y2=0
cc_308 N_A_27_297#_c_309_n Y 0.00223824f $X=5.12 $Y=1.455 $X2=0 $Y2=0
cc_309 N_A_27_297#_c_311_n Y 0.0181862f $X=5.58 $Y=1.16 $X2=0 $Y2=0
cc_310 N_A_27_297#_c_312_n Y 0.00759803f $X=5.855 $Y=1.202 $X2=0 $Y2=0
cc_311 N_A_27_297#_c_307_n N_A_27_47#_M1007_d 0.00318623f $X=0.315 $Y=0.77
+ $X2=-0.19 $Y2=-0.24
cc_312 N_A_27_297#_c_308_n N_A_27_47#_M1007_d 3.84519e-19 $X=0.745 $Y=0.73
+ $X2=-0.19 $Y2=-0.24
cc_313 N_A_27_297#_M1007_s N_A_27_47#_c_660_n 0.00507817f $X=0.56 $Y=0.235 $X2=0
+ $Y2=0
cc_314 N_A_27_297#_c_307_n N_A_27_47#_c_660_n 0.0165567f $X=0.315 $Y=0.77 $X2=0
+ $Y2=0
cc_315 N_A_27_297#_c_308_n N_A_27_47#_c_660_n 0.0313423f $X=0.745 $Y=0.73 $X2=0
+ $Y2=0
cc_316 N_A_27_297#_c_308_n N_A_27_47#_c_661_n 6.23806e-19 $X=0.745 $Y=0.73 $X2=0
+ $Y2=0
cc_317 N_A_27_297#_c_304_n N_VGND_c_707_n 0.00252945f $X=5.36 $Y=0.995 $X2=0
+ $Y2=0
cc_318 N_A_27_297#_c_307_n N_VGND_c_714_n 3.97819e-19 $X=0.315 $Y=0.77 $X2=0
+ $Y2=0
cc_319 N_A_27_297#_c_304_n N_VGND_c_715_n 0.00368123f $X=5.36 $Y=0.995 $X2=0
+ $Y2=0
cc_320 N_A_27_297#_c_305_n N_VGND_c_715_n 0.00368116f $X=5.88 $Y=0.995 $X2=0
+ $Y2=0
cc_321 N_A_27_297#_M1007_s N_VGND_c_716_n 0.00297142f $X=0.56 $Y=0.235 $X2=0
+ $Y2=0
cc_322 N_A_27_297#_c_304_n N_VGND_c_716_n 0.00682404f $X=5.36 $Y=0.995 $X2=0
+ $Y2=0
cc_323 N_A_27_297#_c_305_n N_VGND_c_716_n 0.00649112f $X=5.88 $Y=0.995 $X2=0
+ $Y2=0
cc_324 N_A_27_297#_c_307_n N_VGND_c_716_n 0.00112342f $X=0.315 $Y=0.77 $X2=0
+ $Y2=0
cc_325 N_A_27_297#_c_317_n N_A_600_47#_c_796_n 6.68497e-19 $X=5.035 $Y=1.54
+ $X2=0 $Y2=0
cc_326 N_A_27_297#_c_304_n N_A_600_47#_c_797_n 0.00502358f $X=5.36 $Y=0.995
+ $X2=0 $Y2=0
cc_327 N_A_27_297#_c_305_n N_A_600_47#_c_797_n 0.00147798f $X=5.88 $Y=0.995
+ $X2=0 $Y2=0
cc_328 N_A_27_297#_c_312_n N_A_600_47#_c_797_n 0.0047334f $X=5.855 $Y=1.202
+ $X2=0 $Y2=0
cc_329 N_A_27_297#_c_304_n N_A_600_47#_c_798_n 0.00990301f $X=5.36 $Y=0.995
+ $X2=0 $Y2=0
cc_330 N_A_27_297#_c_317_n N_A_600_47#_c_798_n 0.0225866f $X=5.035 $Y=1.54 $X2=0
+ $Y2=0
cc_331 N_A_27_297#_c_310_n N_A_600_47#_c_798_n 0.0141654f $X=5.205 $Y=1.16 $X2=0
+ $Y2=0
cc_332 N_A_27_297#_c_311_n N_A_600_47#_c_798_n 0.0392005f $X=5.58 $Y=1.16 $X2=0
+ $Y2=0
cc_333 N_VPWR_c_444_n N_A_514_297#_M1000_d 0.00151936f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_334 N_VPWR_c_444_n N_A_514_297#_M1006_d 0.00128721f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_335 N_VPWR_c_444_n N_A_514_297#_M1019_s 0.00215913f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_336 N_VPWR_c_454_n N_A_514_297#_c_550_n 0.0368378f $X=5.025 $Y=2.72 $X2=0
+ $Y2=0
cc_337 N_VPWR_c_444_n N_A_514_297#_c_550_n 0.0212317f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_338 N_VPWR_c_449_n N_A_514_297#_c_580_n 0.0180653f $X=5.15 $Y=2.3 $X2=0 $Y2=0
cc_339 N_VPWR_c_454_n N_A_514_297#_c_580_n 0.0154343f $X=5.025 $Y=2.72 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_444_n N_A_514_297#_c_580_n 0.00938089f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_341 N_VPWR_M1000_s N_A_514_297#_c_556_n 4.93802e-19 $X=3.04 $Y=1.485 $X2=0
+ $Y2=0
cc_342 N_VPWR_c_448_n N_A_514_297#_c_556_n 0.0139466f $X=3.185 $Y=2.3 $X2=0
+ $Y2=0
cc_343 N_VPWR_c_452_n N_A_514_297#_c_556_n 7.89352e-19 $X=3.06 $Y=2.72 $X2=0
+ $Y2=0
cc_344 N_VPWR_c_454_n N_A_514_297#_c_556_n 0.00112424f $X=5.025 $Y=2.72 $X2=0
+ $Y2=0
cc_345 N_VPWR_c_444_n N_A_514_297#_c_556_n 0.060737f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_346 N_VPWR_c_448_n N_A_514_297#_c_558_n 0.0012986f $X=3.185 $Y=2.3 $X2=0
+ $Y2=0
cc_347 N_VPWR_c_452_n N_A_514_297#_c_558_n 4.39771e-19 $X=3.06 $Y=2.72 $X2=0
+ $Y2=0
cc_348 N_VPWR_c_444_n N_A_514_297#_c_558_n 0.028281f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_349 N_VPWR_c_448_n N_A_514_297#_c_569_n 0.00457308f $X=3.185 $Y=2.3 $X2=0
+ $Y2=0
cc_350 N_VPWR_c_452_n N_A_514_297#_c_569_n 0.0154637f $X=3.06 $Y=2.72 $X2=0
+ $Y2=0
cc_351 N_VPWR_c_444_n N_A_514_297#_c_569_n 0.00264208f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_352 N_VPWR_c_448_n N_A_514_297#_c_552_n 3.06455e-19 $X=3.185 $Y=2.3 $X2=0
+ $Y2=0
cc_353 N_VPWR_c_444_n N_A_514_297#_c_552_n 0.0281012f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_354 N_VPWR_c_448_n N_A_514_297#_c_554_n 0.00389626f $X=3.185 $Y=2.3 $X2=0
+ $Y2=0
cc_355 N_VPWR_c_454_n N_A_514_297#_c_554_n 0.0185527f $X=5.025 $Y=2.72 $X2=0
+ $Y2=0
cc_356 N_VPWR_c_444_n N_A_514_297#_c_554_n 0.0029493f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_357 N_VPWR_c_444_n N_Y_M1015_d 0.002602f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_358 N_VPWR_c_444_n N_Y_M1008_s 0.00389781f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_359 N_VPWR_M1008_d N_Y_c_608_n 0.00558454f $X=5.025 $Y=1.485 $X2=0 $Y2=0
cc_360 N_VPWR_c_449_n N_Y_c_608_n 0.016717f $X=5.15 $Y=2.3 $X2=0 $Y2=0
cc_361 N_VPWR_c_454_n N_Y_c_608_n 0.0039015f $X=5.025 $Y=2.72 $X2=0 $Y2=0
cc_362 N_VPWR_c_456_n N_Y_c_608_n 0.00253649f $X=5.965 $Y=2.72 $X2=0 $Y2=0
cc_363 N_VPWR_c_444_n N_Y_c_608_n 0.0135959f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_364 N_VPWR_c_456_n N_Y_c_637_n 0.00444396f $X=5.965 $Y=2.72 $X2=0 $Y2=0
cc_365 N_VPWR_c_444_n N_Y_c_637_n 0.00763999f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_366 N_VPWR_M1010_d Y 0.00328122f $X=5.945 $Y=1.485 $X2=0 $Y2=0
cc_367 N_VPWR_c_451_n Y 0.0281423f $X=6.09 $Y=1.96 $X2=0 $Y2=0
cc_368 N_A_514_297#_c_550_n N_Y_M1015_d 0.0046332f $X=4.505 $Y=2.38 $X2=0.485
+ $Y2=0.56
cc_369 N_A_514_297#_M1019_s N_Y_c_608_n 0.0053134f $X=4.485 $Y=1.485 $X2=3.865
+ $Y2=0.995
cc_370 N_A_514_297#_c_550_n N_Y_c_608_n 0.00625304f $X=4.505 $Y=2.38 $X2=3.865
+ $Y2=0.995
cc_371 N_A_514_297#_c_580_n N_Y_c_608_n 0.0157703f $X=4.63 $Y=2.3 $X2=3.865
+ $Y2=0.995
cc_372 N_A_514_297#_c_550_n N_Y_c_623_n 0.012411f $X=4.505 $Y=2.38 $X2=4.42
+ $Y2=0.56
cc_373 N_A_514_297#_c_552_n N_Y_c_623_n 0.00139207f $X=3.77 $Y=2.21 $X2=4.42
+ $Y2=0.56
cc_374 N_Y_c_605_n N_VGND_c_707_n 0.0100248f $X=5.95 $Y=0.39 $X2=0 $Y2=0
cc_375 N_Y_c_605_n N_VGND_c_715_n 0.0423892f $X=5.95 $Y=0.39 $X2=0 $Y2=0
cc_376 N_Y_c_606_n N_VGND_c_715_n 0.0193947f $X=6.145 $Y=0.475 $X2=0 $Y2=0
cc_377 N_Y_M1001_d N_VGND_c_716_n 0.0021262f $X=5.025 $Y=0.235 $X2=0 $Y2=0
cc_378 N_Y_M1013_d N_VGND_c_716_n 0.00212516f $X=5.955 $Y=0.235 $X2=0 $Y2=0
cc_379 N_Y_c_605_n N_VGND_c_716_n 0.0333931f $X=5.95 $Y=0.39 $X2=0 $Y2=0
cc_380 N_Y_c_606_n N_VGND_c_716_n 0.0145499f $X=6.145 $Y=0.475 $X2=0 $Y2=0
cc_381 N_Y_c_605_n N_A_600_47#_M1001_s 0.00524752f $X=5.95 $Y=0.39 $X2=0 $Y2=0
cc_382 N_Y_c_605_n N_A_600_47#_c_797_n 0.0201898f $X=5.95 $Y=0.39 $X2=0 $Y2=0
cc_383 N_Y_c_607_n N_A_600_47#_c_797_n 0.00969616f $X=6.145 $Y=1.415 $X2=0 $Y2=0
cc_384 Y N_A_600_47#_c_797_n 3.67648e-19 $X=6.11 $Y=1.445 $X2=0 $Y2=0
cc_385 N_Y_M1001_d N_A_600_47#_c_798_n 0.00319929f $X=5.025 $Y=0.235 $X2=0 $Y2=0
cc_386 N_Y_c_605_n N_A_600_47#_c_798_n 0.0177508f $X=5.95 $Y=0.39 $X2=0 $Y2=0
cc_387 N_A_27_47#_c_662_n N_VGND_M1002_s 0.00251047f $X=1.94 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_388 N_A_27_47#_c_669_n N_VGND_c_704_n 0.0141571f $X=1.255 $Y=0.475 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_c_661_n N_VGND_c_704_n 0.00471242f $X=1.255 $Y=0.725 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_c_662_n N_VGND_c_704_n 0.0127273f $X=1.94 $Y=0.815 $X2=0 $Y2=0
cc_391 N_A_27_47#_c_662_n N_VGND_c_705_n 0.00976974f $X=1.94 $Y=0.815 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_663_n N_VGND_c_705_n 0.0241299f $X=2.155 $Y=0.39 $X2=0 $Y2=0
cc_393 N_A_27_47#_c_662_n N_VGND_c_708_n 0.00198695f $X=1.94 $Y=0.815 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_c_663_n N_VGND_c_708_n 0.0244523f $X=2.155 $Y=0.39 $X2=0 $Y2=0
cc_395 N_A_27_47#_c_660_n N_VGND_c_714_n 0.0590541f $X=1.13 $Y=0.365 $X2=0 $Y2=0
cc_396 N_A_27_47#_c_669_n N_VGND_c_714_n 0.0152108f $X=1.255 $Y=0.475 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_c_662_n N_VGND_c_714_n 0.00266636f $X=1.94 $Y=0.815 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_M1007_d N_VGND_c_716_n 0.00221642f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_M1017_d N_VGND_c_716_n 0.00215206f $X=1.08 $Y=0.235 $X2=0
+ $Y2=0
cc_400 N_A_27_47#_M1003_d N_VGND_c_716_n 0.00266705f $X=1.97 $Y=0.235 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_c_660_n N_VGND_c_716_n 0.036878f $X=1.13 $Y=0.365 $X2=0 $Y2=0
cc_402 N_A_27_47#_c_669_n N_VGND_c_716_n 0.00940698f $X=1.255 $Y=0.475 $X2=0
+ $Y2=0
cc_403 N_A_27_47#_c_662_n N_VGND_c_716_n 0.00972452f $X=1.94 $Y=0.815 $X2=0
+ $Y2=0
cc_404 N_A_27_47#_c_663_n N_VGND_c_716_n 0.0143352f $X=2.155 $Y=0.39 $X2=0 $Y2=0
cc_405 N_VGND_c_716_n N_A_600_47#_M1011_s 0.00304143f $X=6.21 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_406 N_VGND_c_716_n N_A_600_47#_M1004_s 0.0033305f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_407 N_VGND_c_716_n N_A_600_47#_M1001_s 0.00301822f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_408 N_VGND_c_710_n N_A_600_47#_c_808_n 0.0231806f $X=3.57 $Y=0 $X2=0 $Y2=0
cc_409 N_VGND_c_716_n N_A_600_47#_c_808_n 0.0143352f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_410 N_VGND_M1018_d N_A_600_47#_c_794_n 0.00162089f $X=3.52 $Y=0.235 $X2=0
+ $Y2=0
cc_411 N_VGND_c_706_n N_A_600_47#_c_794_n 0.0122559f $X=3.655 $Y=0.39 $X2=0
+ $Y2=0
cc_412 N_VGND_c_710_n N_A_600_47#_c_794_n 0.00254521f $X=3.57 $Y=0 $X2=0 $Y2=0
cc_413 N_VGND_c_712_n N_A_600_47#_c_794_n 0.00198695f $X=4.545 $Y=0 $X2=0 $Y2=0
cc_414 N_VGND_c_716_n N_A_600_47#_c_794_n 0.0094839f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_415 N_VGND_c_705_n N_A_600_47#_c_795_n 0.00830019f $X=2.715 $Y=0.39 $X2=0
+ $Y2=0
cc_416 N_VGND_c_712_n N_A_600_47#_c_803_n 0.0256662f $X=4.545 $Y=0 $X2=0 $Y2=0
cc_417 N_VGND_c_716_n N_A_600_47#_c_803_n 0.0157539f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_418 N_VGND_M1014_d N_A_600_47#_c_798_n 0.00315681f $X=4.495 $Y=0.235 $X2=0
+ $Y2=0
cc_419 N_VGND_c_707_n N_A_600_47#_c_798_n 0.0127273f $X=4.63 $Y=0.39 $X2=0 $Y2=0
cc_420 N_VGND_c_712_n N_A_600_47#_c_798_n 0.00254521f $X=4.545 $Y=0 $X2=0 $Y2=0
cc_421 N_VGND_c_715_n N_A_600_47#_c_798_n 0.00409419f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_422 N_VGND_c_716_n N_A_600_47#_c_798_n 0.0137746f $X=6.21 $Y=0 $X2=0 $Y2=0
