* NGSPICE file created from sky130_fd_sc_hdll__and2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__and2b_2 A_N B VGND VNB VPB VPWR X
M1000 VPWR a_230_413# X VPB phighvt w=1e+06u l=180000u
+  ad=9.248e+11p pd=7.78e+06u as=4.5e+11p ps=2.9e+06u
M1001 VPWR A_N a_27_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1002 VGND B a_327_47# VNB nshort w=420000u l=150000u
+  ad=5.4195e+11p pd=5.38e+06u as=1.344e+11p ps=1.48e+06u
M1003 VPWR B a_230_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1004 VGND a_230_413# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.12e+11p ps=2.26e+06u
M1005 a_327_47# a_27_413# a_230_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1006 a_27_413# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1007 X a_230_413# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_230_413# a_27_413# VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_230_413# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

