* File: sky130_fd_sc_hdll__clkbuf_4.pex.spice
* Created: Wed Sep  2 08:25:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_4%A 1 3 6 8 9
c33 1 0 1.51211e-19 $X=0.5 $Y=1.41
r34 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r35 9 14 0.864332 $w=3.98e-07 $l=3e-08 $layer=LI1_cond $X=0.625 $Y=1.19
+ $X2=0.625 $Y2=1.16
r36 8 14 8.93143 $w=3.98e-07 $l=3.1e-07 $layer=LI1_cond $X=0.625 $Y=0.85
+ $X2=0.625 $Y2=1.16
r37 4 13 38.5462 $w=3.19e-07 $l=1.67481e-07 $layer=POLY_cond $X=0.525 $Y=0.995
+ $X2=0.52 $Y2=1.16
r38 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.525 $Y=0.995
+ $X2=0.525 $Y2=0.445
r39 1 13 46.8511 $w=3.19e-07 $l=2.59808e-07 $layer=POLY_cond $X=0.5 $Y=1.41
+ $X2=0.52 $Y2=1.16
r40 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_4%A_27_47# 1 2 9 11 13 16 18 20 21 25 27 29
+ 30 32 34 37 40 41 42 43 45 48 50 53 54 59 60 65 67
c106 54 0 1.51211e-19 $X=1.215 $Y=1.16
c107 53 0 2.11231e-19 $X=1.105 $Y=1.495
c108 27 0 2.35182e-20 $X=1.99 $Y=1.41
r109 62 65 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.17 $Y=0.42 $X2=0.26
+ $Y2=0.42
r110 59 60 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.07
+ $Y=1.16 $X2=2.07 $Y2=1.16
r111 56 59 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.34 $Y=1.16
+ $X2=2.07 $Y2=1.16
r112 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.34
+ $Y=1.16 $X2=1.34 $Y2=1.16
r113 54 56 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.215 $Y=1.16
+ $X2=1.34 $Y2=1.16
r114 52 54 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.105 $Y=1.245
+ $X2=1.215 $Y2=1.16
r115 52 53 13.0959 $w=2.18e-07 $l=2.5e-07 $layer=LI1_cond $X=1.105 $Y=1.245
+ $X2=1.105 $Y2=1.495
r116 51 67 2.60907 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.395 $Y=1.58
+ $X2=0.24 $Y2=1.58
r117 50 53 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.995 $Y=1.58
+ $X2=1.105 $Y2=1.495
r118 50 51 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=0.995 $Y=1.58
+ $X2=0.395 $Y2=1.58
r119 46 67 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=1.58
r120 46 48 0.92939 $w=3.08e-07 $l=2.5e-08 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=1.69
r121 45 67 3.84343 $w=2.4e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.17 $Y=1.495
+ $X2=0.24 $Y2=1.58
r122 44 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.17 $Y2=0.42
r123 44 45 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.17 $Y2=1.495
r124 41 57 15.2694 $w=2.75e-07 $l=7e-08 $layer=POLY_cond $X=1.41 $Y=1.157
+ $X2=1.34 $Y2=1.157
r125 41 42 6.52665 $w=2.75e-07 $l=1.25698e-07 $layer=POLY_cond $X=1.41 $Y=1.157
+ $X2=1.51 $Y2=1.215
r126 39 57 45.8082 $w=2.75e-07 $l=2.1e-07 $layer=POLY_cond $X=1.13 $Y=1.157
+ $X2=1.34 $Y2=1.157
r127 39 40 1.63566 $w=2.75e-07 $l=1.25698e-07 $layer=POLY_cond $X=1.13 $Y=1.157
+ $X2=1.03 $Y2=1.215
r128 35 43 30.4925 $w=1.65e-07 $l=2.07123e-07 $layer=POLY_cond $X=2.495 $Y=1.02
+ $X2=2.47 $Y2=1.215
r129 35 37 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.495 $Y=1.02
+ $X2=2.495 $Y2=0.445
r130 32 43 30.4925 $w=1.65e-07 $l=1.95e-07 $layer=POLY_cond $X=2.47 $Y=1.41
+ $X2=2.47 $Y2=1.215
r131 32 34 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.47 $Y=1.41
+ $X2=2.47 $Y2=1.985
r132 31 60 6.52665 $w=2.75e-07 $l=1.25698e-07 $layer=POLY_cond $X=2.09 $Y=1.157
+ $X2=1.99 $Y2=1.215
r133 30 43 1.63566 $w=2.75e-07 $l=1.25698e-07 $layer=POLY_cond $X=2.37 $Y=1.157
+ $X2=2.47 $Y2=1.215
r134 30 31 61.0776 $w=2.75e-07 $l=2.8e-07 $layer=POLY_cond $X=2.37 $Y=1.157
+ $X2=2.09 $Y2=1.157
r135 27 60 18.6979 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=1.99 $Y=1.41
+ $X2=1.99 $Y2=1.215
r136 27 29 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.99 $Y=1.41
+ $X2=1.99 $Y2=1.985
r137 23 60 18.6979 $w=1.5e-07 $l=2.04756e-07 $layer=POLY_cond $X=1.97 $Y=1.02
+ $X2=1.99 $Y2=1.215
r138 23 25 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.97 $Y=1.02
+ $X2=1.97 $Y2=0.445
r139 22 42 6.52665 $w=2.75e-07 $l=1.25698e-07 $layer=POLY_cond $X=1.61 $Y=1.157
+ $X2=1.51 $Y2=1.215
r140 21 60 6.52665 $w=2.75e-07 $l=1.25698e-07 $layer=POLY_cond $X=1.89 $Y=1.157
+ $X2=1.99 $Y2=1.215
r141 21 22 61.0776 $w=2.75e-07 $l=2.8e-07 $layer=POLY_cond $X=1.89 $Y=1.157
+ $X2=1.61 $Y2=1.157
r142 18 42 18.6979 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=1.51 $Y=1.41
+ $X2=1.51 $Y2=1.215
r143 18 20 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.51 $Y=1.41
+ $X2=1.51 $Y2=1.985
r144 14 42 18.6979 $w=1.5e-07 $l=2.04756e-07 $layer=POLY_cond $X=1.49 $Y=1.02
+ $X2=1.51 $Y2=1.215
r145 14 16 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.49 $Y=1.02
+ $X2=1.49 $Y2=0.445
r146 11 40 30.4925 $w=1.65e-07 $l=1.95e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.03 $Y2=1.215
r147 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.03 $Y2=1.985
r148 7 40 30.4925 $w=1.65e-07 $l=2.07123e-07 $layer=POLY_cond $X=1.005 $Y=1.02
+ $X2=1.03 $Y2=1.215
r149 7 9 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.005 $Y=1.02
+ $X2=1.005 $Y2=0.445
r150 2 48 300 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.69
r151 1 65 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_4%VPWR 1 2 3 14 18 22 25 26 28 29 30 40 41
+ 44
r45 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r46 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r47 38 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r48 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r49 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r50 35 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r51 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r52 32 44 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=0.77 $Y2=2.72
r53 32 34 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=1.61 $Y2=2.72
r54 30 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r55 28 37 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.53 $Y2=2.72
r56 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.71 $Y2=2.72
r57 27 40 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.875 $Y=2.72
+ $X2=2.99 $Y2=2.72
r58 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=2.72
+ $X2=2.71 $Y2=2.72
r59 25 34 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.625 $Y=2.72
+ $X2=1.61 $Y2=2.72
r60 25 26 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.625 $Y=2.72
+ $X2=1.752 $Y2=2.72
r61 24 37 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.88 $Y=2.72
+ $X2=2.53 $Y2=2.72
r62 24 26 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.88 $Y=2.72
+ $X2=1.752 $Y2=2.72
r63 20 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=2.635
+ $X2=2.71 $Y2=2.72
r64 20 22 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=2.71 $Y=2.635
+ $X2=2.71 $Y2=1.93
r65 16 26 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.752 $Y=2.635
+ $X2=1.752 $Y2=2.72
r66 16 18 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=1.752 $Y=2.635
+ $X2=1.752 $Y2=2.34
r67 12 44 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=2.635
+ $X2=0.77 $Y2=2.72
r68 12 14 23.6065 $w=3.08e-07 $l=6.35e-07 $layer=LI1_cond $X=0.77 $Y=2.635
+ $X2=0.77 $Y2=2
r69 3 22 300 $w=1.7e-07 $l=5.14563e-07 $layer=licon1_PDIFF $count=2 $X=2.56
+ $Y=1.485 $X2=2.71 $Y2=1.93
r70 2 18 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.6
+ $Y=1.485 $X2=1.75 $Y2=2.34
r71 1 14 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=1.485 $X2=0.74 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_4%X 1 2 3 4 15 19 21 22 23 24 27 34 35 36
+ 37 43
c70 36 0 2.35182e-20 $X=2.79 $Y=0.85
c71 3 0 1.10391e-19 $X=1.12 $Y=1.485
r72 37 43 5.38235 $w=4.98e-07 $l=2.25e-07 $layer=LI1_cond $X=2.66 $Y=1.19
+ $X2=2.66 $Y2=1.415
r73 36 42 2.53623 $w=3.8e-07 $l=1.90825e-07 $layer=LI1_cond $X=2.507 $Y=0.82
+ $X2=2.66 $Y2=0.905
r74 36 37 6.45882 $w=4.98e-07 $l=2.7e-07 $layer=LI1_cond $X=2.66 $Y=0.92
+ $X2=2.66 $Y2=1.19
r75 36 42 0.358824 $w=4.98e-07 $l=1.5e-08 $layer=LI1_cond $X=2.66 $Y=0.92
+ $X2=2.66 $Y2=0.905
r76 35 43 19.1257 $w=2.33e-07 $l=3.9e-07 $layer=LI1_cond $X=2.27 $Y=1.532
+ $X2=2.66 $Y2=1.532
r77 35 48 1.96161 $w=2.33e-07 $l=4e-08 $layer=LI1_cond $X=2.27 $Y=1.532 $X2=2.23
+ $Y2=1.532
r78 30 34 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.235 $Y=1.835
+ $X2=2.235 $Y2=1.92
r79 29 48 0.0901955 $w=2.6e-07 $l=1.20474e-07 $layer=LI1_cond $X=2.235 $Y=1.65
+ $X2=2.23 $Y2=1.532
r80 29 30 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=2.235 $Y=1.65
+ $X2=2.235 $Y2=1.835
r81 25 36 2.53623 $w=3.8e-07 $l=3.11615e-07 $layer=LI1_cond $X=2.235 $Y=0.735
+ $X2=2.507 $Y2=0.82
r82 25 27 9.97306 $w=2.58e-07 $l=2.25e-07 $layer=LI1_cond $X=2.235 $Y=0.735
+ $X2=2.235 $Y2=0.51
r83 23 34 2.90867 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.105 $Y=1.92
+ $X2=2.235 $Y2=1.92
r84 23 24 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.105 $Y=1.92
+ $X2=1.405 $Y2=1.92
r85 21 36 4.34722 $w=1.7e-07 $l=4.02e-07 $layer=LI1_cond $X=2.105 $Y=0.82
+ $X2=2.507 $Y2=0.82
r86 21 22 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.105 $Y=0.82
+ $X2=1.405 $Y2=0.82
r87 17 24 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.275 $Y=2.005
+ $X2=1.405 $Y2=1.92
r88 17 19 7.09196 $w=2.58e-07 $l=1.6e-07 $layer=LI1_cond $X=1.275 $Y=2.005
+ $X2=1.275 $Y2=2.165
r89 13 22 7.97992 $w=1.7e-07 $l=2.16365e-07 $layer=LI1_cond $X=1.227 $Y=0.735
+ $X2=1.405 $Y2=0.82
r90 13 15 7.30422 $w=3.53e-07 $l=2.25e-07 $layer=LI1_cond $X=1.227 $Y=0.735
+ $X2=1.227 $Y2=0.51
r91 4 48 600 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=1 $X=2.08
+ $Y=1.485 $X2=2.23 $Y2=1.62
r92 4 34 300 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=2 $X=2.08
+ $Y=1.485 $X2=2.23 $Y2=1.96
r93 3 19 600 $w=1.7e-07 $l=7.51266e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.485 $X2=1.27 $Y2=2.165
r94 2 27 182 $w=1.7e-07 $l=3.57596e-07 $layer=licon1_NDIFF $count=1 $X=2.045
+ $Y=0.235 $X2=2.235 $Y2=0.51
r95 1 15 182 $w=1.7e-07 $l=3.59514e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.235 $X2=1.275 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_4%VGND 1 2 3 12 16 20 23 24 26 27 28 30 43
+ 44 47
r47 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r48 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r49 41 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r50 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r51 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r52 38 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r53 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r54 35 47 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.742
+ $Y2=0
r55 35 37 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=1.61
+ $Y2=0
r56 30 47 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.742
+ $Y2=0
r57 30 32 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.23
+ $Y2=0
r58 28 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r59 28 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r60 26 40 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.585 $Y=0 $X2=2.53
+ $Y2=0
r61 26 27 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.585 $Y=0 $X2=2.725
+ $Y2=0
r62 25 43 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.99
+ $Y2=0
r63 25 27 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.725
+ $Y2=0
r64 23 37 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.625 $Y=0 $X2=1.61
+ $Y2=0
r65 23 24 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.625 $Y=0 $X2=1.752
+ $Y2=0
r66 22 40 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=2.53
+ $Y2=0
r67 22 24 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=1.752
+ $Y2=0
r68 18 27 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=0.085
+ $X2=2.725 $Y2=0
r69 18 20 12.965 $w=2.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.725 $Y=0.085
+ $X2=2.725 $Y2=0.4
r70 14 24 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.752 $Y=0.085
+ $X2=1.752 $Y2=0
r71 14 16 14.2361 $w=2.53e-07 $l=3.15e-07 $layer=LI1_cond $X=1.752 $Y=0.085
+ $X2=1.752 $Y2=0.4
r72 10 47 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.742 $Y=0.085
+ $X2=0.742 $Y2=0
r73 10 12 13.2007 $w=2.73e-07 $l=3.15e-07 $layer=LI1_cond $X=0.742 $Y=0.085
+ $X2=0.742 $Y2=0.4
r74 3 20 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=2.57
+ $Y=0.235 $X2=2.715 $Y2=0.4
r75 2 16 182 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_NDIFF $count=1 $X=1.565
+ $Y=0.235 $X2=1.755 $Y2=0.4
r76 1 12 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.235 $X2=0.74 $Y2=0.4
.ends

