* File: sky130_fd_sc_hdll__nand2_1.pxi.spice
* Created: Wed Sep  2 08:36:36 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND2_1%B N_B_c_31_n N_B_M1000_g N_B_c_28_n N_B_M1002_g
+ B N_B_c_30_n PM_SKY130_FD_SC_HDLL__NAND2_1%B
x_PM_SKY130_FD_SC_HDLL__NAND2_1%A N_A_c_52_n N_A_M1001_g N_A_c_53_n N_A_M1003_g
+ A PM_SKY130_FD_SC_HDLL__NAND2_1%A
x_PM_SKY130_FD_SC_HDLL__NAND2_1%VPWR N_VPWR_M1000_s N_VPWR_M1003_d N_VPWR_c_75_n
+ N_VPWR_c_76_n N_VPWR_c_77_n N_VPWR_c_78_n VPWR N_VPWR_c_79_n N_VPWR_c_74_n
+ N_VPWR_c_81_n PM_SKY130_FD_SC_HDLL__NAND2_1%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND2_1%Y N_Y_M1001_d N_Y_M1000_d Y Y Y Y Y N_Y_c_99_n
+ PM_SKY130_FD_SC_HDLL__NAND2_1%Y
x_PM_SKY130_FD_SC_HDLL__NAND2_1%VGND N_VGND_M1002_s N_VGND_c_126_n
+ N_VGND_c_127_n VGND N_VGND_c_128_n N_VGND_c_129_n VGND
+ PM_SKY130_FD_SC_HDLL__NAND2_1%VGND
cc_1 VNB N_B_c_28_n 0.0221895f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_2 VNB B 0.00939618f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_3 VNB N_B_c_30_n 0.0436531f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_4 VNB N_A_c_52_n 0.0221092f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_5 VNB N_A_c_53_n 0.0409484f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_6 VNB A 0.0087026f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_7 VNB N_VPWR_c_74_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB Y 0.00793185f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_9 VNB N_Y_c_99_n 0.0276021f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_VGND_c_126_n 0.0108751f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_11 VNB N_VGND_c_127_n 0.0330625f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.56
cc_12 VNB N_VGND_c_128_n 0.0409804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VGND_c_129_n 0.137581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VPB N_B_c_31_n 0.0212147f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_15 VPB B 8.02347e-19 $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_16 VPB N_B_c_30_n 0.0191277f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_17 VPB N_A_c_53_n 0.039824f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_18 VPB A 7.2205e-19 $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_19 VPB N_VPWR_c_75_n 0.0102689f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_20 VPB N_VPWR_c_76_n 0.0444141f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.202
cc_21 VPB N_VPWR_c_77_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.202
cc_22 VPB N_VPWR_c_78_n 0.0432431f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_23 VPB N_VPWR_c_79_n 0.0163041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_24 VPB N_VPWR_c_74_n 0.0569095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_25 VPB N_VPWR_c_81_n 0.00497514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_26 VPB Y 0.00313618f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_27 VPB Y 2.54765e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 N_B_c_28_n N_A_c_52_n 0.0280333f $X=0.54 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_29 N_B_c_31_n N_A_c_53_n 0.00882543f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_30 N_B_c_30_n N_A_c_53_n 0.0280333f $X=0.515 $Y=1.202 $X2=0 $Y2=0
cc_31 N_B_c_31_n N_VPWR_c_76_n 0.00787079f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_32 B N_VPWR_c_76_n 0.0220525f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_33 N_B_c_30_n N_VPWR_c_76_n 0.00603357f $X=0.515 $Y=1.202 $X2=0 $Y2=0
cc_34 N_B_c_31_n N_VPWR_c_77_n 0.00597712f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_35 N_B_c_31_n N_VPWR_c_74_n 0.0109493f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_36 N_B_c_31_n Y 0.00180793f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_37 N_B_c_28_n Y 0.00882417f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_38 B Y 0.0166798f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_39 N_B_c_31_n Y 0.0120229f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_40 N_B_c_31_n Y 0.00662085f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_41 N_B_c_28_n N_VGND_c_127_n 0.00761923f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_42 B N_VGND_c_127_n 0.0244951f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_43 N_B_c_30_n N_VGND_c_127_n 0.00724028f $X=0.515 $Y=1.202 $X2=0 $Y2=0
cc_44 N_B_c_28_n N_VGND_c_128_n 0.00585385f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_45 N_B_c_28_n N_VGND_c_129_n 0.0117063f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_46 N_A_c_53_n N_VPWR_c_77_n 0.00673617f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_47 N_A_c_53_n N_VPWR_c_78_n 0.0141353f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_48 A N_VPWR_c_78_n 0.019414f $X=1.16 $Y=1.105 $X2=0 $Y2=0
cc_49 N_A_c_53_n N_VPWR_c_74_n 0.0131514f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_50 N_A_c_52_n Y 0.00857971f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_51 N_A_c_53_n Y 0.00173999f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_52 A Y 0.0189505f $X=1.16 $Y=1.105 $X2=0 $Y2=0
cc_53 N_A_c_53_n Y 0.00989133f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_54 N_A_c_53_n Y 0.00314168f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_55 N_A_c_52_n N_Y_c_99_n 0.0211053f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_56 N_A_c_53_n N_Y_c_99_n 0.00856845f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_57 A N_Y_c_99_n 0.0258904f $X=1.16 $Y=1.105 $X2=0 $Y2=0
cc_58 N_A_c_52_n N_VGND_c_128_n 0.00357877f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_59 N_A_c_52_n N_VGND_c_129_n 0.00657948f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_60 N_VPWR_c_74_n N_Y_M1000_d 0.00231261f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_61 N_VPWR_c_77_n Y 0.0223557f $X=1.135 $Y=2.72 $X2=0 $Y2=0
cc_62 N_VPWR_c_74_n Y 0.0140101f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_63 N_VPWR_c_76_n Y 0.0751091f $X=0.28 $Y=1.66 $X2=0 $Y2=0
cc_64 N_VPWR_c_78_n Y 0.0612532f $X=1.22 $Y=1.66 $X2=0 $Y2=0
cc_65 N_VPWR_c_78_n N_Y_c_99_n 7.22395e-19 $X=1.22 $Y=1.66 $X2=0 $Y2=0
cc_66 N_VPWR_c_76_n N_VGND_c_127_n 3.44647e-19 $X=0.28 $Y=1.66 $X2=0 $Y2=0
cc_67 N_Y_c_99_n N_VGND_c_128_n 0.0468195f $X=1.22 $Y=0.38 $X2=0 $Y2=0
cc_68 N_Y_M1001_d N_VGND_c_129_n 0.00250339f $X=1.035 $Y=0.235 $X2=0 $Y2=0
cc_69 N_Y_c_99_n N_VGND_c_129_n 0.0278594f $X=1.22 $Y=0.38 $X2=0 $Y2=0
cc_70 Y A_123_47# 4.34665e-19 $X=0.65 $Y=1.48 $X2=-0.19 $Y2=-0.24
cc_71 N_Y_c_99_n A_123_47# 0.00325659f $X=1.22 $Y=0.38 $X2=-0.19 $Y2=-0.24
cc_72 N_VGND_c_129_n A_123_47# 0.00338335f $X=1.61 $Y=0 $X2=-0.19 $Y2=-0.24
