* File: sky130_fd_sc_hdll__o221a_4.pex.spice
* Created: Thu Aug 27 19:20:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O221A_4%C1 1 3 4 6 7 9 10 12 13 20 23
c40 10 0 1.62953e-19 $X=0.99 $Y=0.995
r41 20 21 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r42 19 20 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.965 $Y2=1.202
r43 18 19 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r44 16 18 29.0521 $w=3.65e-07 $l=2.2e-07 $layer=POLY_cond $X=0.275 $Y=1.202
+ $X2=0.495 $Y2=1.202
r45 13 23 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.23 $Y2=1.175
r46 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r47 10 21 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r48 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r49 7 20 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r50 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r51 4 19 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r52 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r53 1 18 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r54 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_4%B1 1 3 4 6 7 9 10 12 13 16 21 32 34
c75 1 0 1.58247e-19 $X=1.435 $Y=1.41
r76 32 34 13.2011 $w=5.38e-07 $l=3.2e-07 $layer=LI1_cond $X=1.41 $Y=1.345
+ $X2=1.73 $Y2=1.345
r77 26 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.41
+ $Y=1.16 $X2=1.41 $Y2=1.16
r78 21 32 3.43319 $w=5.38e-07 $l=1.55e-07 $layer=LI1_cond $X=1.255 $Y=1.345
+ $X2=1.41 $Y2=1.345
r79 16 19 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.855 $Y=1.16
+ $X2=2.855 $Y2=1.53
r80 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.83
+ $Y=1.16 $X2=2.83 $Y2=1.16
r81 13 19 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.665 $Y=1.53
+ $X2=2.855 $Y2=1.53
r82 13 34 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=2.665 $Y=1.53 $X2=1.73
+ $Y2=1.53
r83 10 17 38.578 $w=2.95e-07 $l=1.72337e-07 $layer=POLY_cond $X=2.87 $Y=0.995
+ $X2=2.855 $Y2=1.16
r84 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.87 $Y=0.995
+ $X2=2.87 $Y2=0.56
r85 7 17 48.1208 $w=2.95e-07 $l=2.54951e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.855 $Y2=1.16
r86 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r87 4 26 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.435 $Y2=1.16
r88 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.46 $Y=0.995 $X2=1.46
+ $Y2=0.56
r89 1 26 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.16
r90 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_4%B2 1 3 4 6 7 9 10 12 13 20 23
c42 13 0 1.58247e-19 $X=2.19 $Y=1.105
r43 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.4 $Y2=1.202
r44 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=2.14 $Y=1.202
+ $X2=2.375 $Y2=1.202
r45 18 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.16 $X2=2.14 $Y2=1.16
r46 16 18 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=2.14 $Y2=1.202
r47 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.88 $Y=1.202
+ $X2=1.905 $Y2=1.202
r48 13 23 11.0909 $w=1.98e-07 $l=2e-07 $layer=LI1_cond $X=2.275 $Y=1.175
+ $X2=2.075 $Y2=1.175
r49 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.4 $Y=0.995
+ $X2=2.4 $Y2=1.202
r50 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.4 $Y=0.995 $X2=2.4
+ $Y2=0.56
r51 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r52 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r53 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r54 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r55 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.88 $Y=0.995
+ $X2=1.88 $Y2=1.202
r56 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.88 $Y=0.995 $X2=1.88
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_4%A1 1 3 4 6 7 9 10 12 13 16 21 22 32
c77 21 0 1.04028e-19 $X=5.1 $Y=1.445
c78 13 0 1.46864e-19 $X=4.975 $Y=1.53
c79 7 0 3.35826e-19 $X=5.245 $Y=1.41
r80 30 32 3.88182 $w=1.98e-07 $l=7e-08 $layer=LI1_cond $X=5.225 $Y=1.175
+ $X2=5.295 $Y2=1.175
r81 22 30 3.84807 $w=2e-07 $l=1.25e-07 $layer=LI1_cond $X=5.1 $Y=1.175 $X2=5.225
+ $Y2=1.175
r82 22 32 0.388182 $w=1.98e-07 $l=7e-09 $layer=LI1_cond $X=5.302 $Y=1.175
+ $X2=5.295 $Y2=1.175
r83 22 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.22
+ $Y=1.16 $X2=5.22 $Y2=1.16
r84 21 22 7.44331 $w=2.63e-07 $l=1.7e-07 $layer=LI1_cond $X=5.1 $Y=1.445 $X2=5.1
+ $Y2=1.275
r85 16 19 6.80845 $w=6.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.63 $Y=1.16
+ $X2=3.63 $Y2=1.53
r86 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.74
+ $Y=1.16 $X2=3.74 $Y2=1.16
r87 14 19 8.83581 $w=1.7e-07 $l=3.25e-07 $layer=LI1_cond $X=3.955 $Y=1.53
+ $X2=3.63 $Y2=1.53
r88 13 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.975 $Y=1.53
+ $X2=5.1 $Y2=1.445
r89 13 14 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=4.975 $Y=1.53
+ $X2=3.955 $Y2=1.53
r90 10 28 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=5.27 $Y=0.995
+ $X2=5.245 $Y2=1.16
r91 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.27 $Y=0.995
+ $X2=5.27 $Y2=0.56
r92 7 28 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.16
r93 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.985
r94 4 17 38.5416 $w=3.03e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.86 $Y=0.995
+ $X2=3.77 $Y2=1.16
r95 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.86 $Y=0.995 $X2=3.86
+ $Y2=0.56
r96 1 17 47.6478 $w=3.03e-07 $l=2.80624e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.77 $Y2=1.16
r97 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_4%A2 1 3 4 6 7 9 10 12 13 19 20 25
c50 19 0 1.69964e-19 $X=4.54 $Y=1.16
r51 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.775 $Y=1.202
+ $X2=4.8 $Y2=1.202
r52 19 25 11.0909 $w=1.98e-07 $l=2e-07 $layer=LI1_cond $X=4.54 $Y=1.175 $X2=4.34
+ $Y2=1.175
r53 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=4.54 $Y=1.202
+ $X2=4.775 $Y2=1.202
r54 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.54
+ $Y=1.16 $X2=4.54 $Y2=1.16
r55 16 18 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=4.305 $Y=1.202
+ $X2=4.54 $Y2=1.202
r56 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.28 $Y=1.202
+ $X2=4.305 $Y2=1.202
r57 13 25 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=4.325 $Y=1.175
+ $X2=4.34 $Y2=1.175
r58 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.8 $Y=0.995
+ $X2=4.8 $Y2=1.202
r59 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.8 $Y=0.995 $X2=4.8
+ $Y2=0.56
r60 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.202
r61 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
r62 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.202
r63 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.985
r64 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.28 $Y=0.995
+ $X2=4.28 $Y2=1.202
r65 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.28 $Y=0.995 $X2=4.28
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_4%A_117_297# 1 2 3 4 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 40 43 45 52 54 55 60 64 67 80
c151 55 0 1.65862e-19 $X=5.925 $Y=1.175
c152 16 0 2.50891e-19 $X=5.715 $Y=1.41
r153 80 81 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.125 $Y=1.202
+ $X2=7.15 $Y2=1.202
r154 77 78 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.63 $Y=1.202
+ $X2=6.655 $Y2=1.202
r155 76 77 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=6.185 $Y=1.202
+ $X2=6.63 $Y2=1.202
r156 75 76 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.16 $Y=1.202
+ $X2=6.185 $Y2=1.202
r157 72 73 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.69 $Y=1.202
+ $X2=5.715 $Y2=1.202
r158 64 66 4.9152 $w=3.78e-07 $l=1.35e-07 $layer=LI1_cond $X=0.705 $Y=0.73
+ $X2=0.705 $Y2=0.865
r159 61 80 30.4489 $w=3.72e-07 $l=2.35e-07 $layer=POLY_cond $X=6.89 $Y=1.202
+ $X2=7.125 $Y2=1.202
r160 61 78 30.4489 $w=3.72e-07 $l=2.35e-07 $layer=POLY_cond $X=6.89 $Y=1.202
+ $X2=6.655 $Y2=1.202
r161 60 61 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.89
+ $Y=1.16 $X2=6.89 $Y2=1.16
r162 58 75 27.2097 $w=3.72e-07 $l=2.1e-07 $layer=POLY_cond $X=5.95 $Y=1.202
+ $X2=6.16 $Y2=1.202
r163 58 73 30.4489 $w=3.72e-07 $l=2.35e-07 $layer=POLY_cond $X=5.95 $Y=1.202
+ $X2=5.715 $Y2=1.202
r164 57 60 52.1273 $w=1.98e-07 $l=9.4e-07 $layer=LI1_cond $X=5.95 $Y=1.175
+ $X2=6.89 $Y2=1.175
r165 57 58 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.95
+ $Y=1.16 $X2=5.95 $Y2=1.16
r166 55 57 1.38636 $w=1.98e-07 $l=2.5e-08 $layer=LI1_cond $X=5.925 $Y=1.175
+ $X2=5.95 $Y2=1.175
r167 54 68 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.815 $Y=1.53
+ $X2=5.56 $Y2=1.53
r168 53 55 6.83662 $w=2e-07 $l=1.51987e-07 $layer=LI1_cond $X=5.815 $Y=1.275
+ $X2=5.925 $Y2=1.175
r169 53 54 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=5.815 $Y=1.275
+ $X2=5.815 $Y2=1.445
r170 51 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.56 $Y=1.615
+ $X2=5.56 $Y2=1.53
r171 51 52 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.56 $Y=1.615
+ $X2=5.56 $Y2=1.785
r172 48 50 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.14 $Y=1.87
+ $X2=4.54 $Y2=1.87
r173 46 67 2.98021 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.895 $Y=1.87
+ $X2=0.755 $Y2=1.87
r174 46 48 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=0.895 $Y=1.87
+ $X2=2.14 $Y2=1.87
r175 45 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.475 $Y=1.87
+ $X2=5.56 $Y2=1.785
r176 45 50 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=5.475 $Y=1.87 $X2=4.54
+ $Y2=1.87
r177 41 67 3.52026 $w=2.65e-07 $l=9.21954e-08 $layer=LI1_cond $X=0.74 $Y=1.955
+ $X2=0.755 $Y2=1.87
r178 41 43 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.74 $Y=1.955
+ $X2=0.74 $Y2=1.96
r179 40 66 31.0748 $w=2.78e-07 $l=7.55e-07 $layer=LI1_cond $X=0.755 $Y=1.62
+ $X2=0.755 $Y2=0.865
r180 38 67 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=1.785
+ $X2=0.755 $Y2=1.87
r181 38 40 6.79118 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=0.755 $Y=1.785
+ $X2=0.755 $Y2=1.62
r182 34 81 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.15 $Y=0.995
+ $X2=7.15 $Y2=1.202
r183 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.15 $Y=0.995
+ $X2=7.15 $Y2=0.56
r184 31 80 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.202
r185 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.985
r186 28 78 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.202
r187 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.985
r188 25 77 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=1.202
r189 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=0.56
r190 22 76 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.202
r191 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.985
r192 19 75 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=1.202
r193 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=0.56
r194 16 73 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.202
r195 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.985
r196 13 72 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=1.202
r197 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=0.56
r198 4 50 600 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.485 $X2=4.54 $Y2=1.87
r199 3 48 600 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.87
r200 2 43 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.96
r201 2 40 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.62
r202 1 64 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_4%VPWR 1 2 3 4 5 6 19 21 25 29 33 37 41 44
+ 45 47 48 50 51 52 73 74 80 85 91
c110 5 0 1.27647e-19 $X=6.275 $Y=1.485
r111 90 91 9.97279 $w=6.78e-07 $l=1.25e-07 $layer=LI1_cond $X=3.6 $Y=2.465
+ $X2=3.725 $Y2=2.465
r112 87 90 2.63841 $w=6.78e-07 $l=1.5e-07 $layer=LI1_cond $X=3.45 $Y=2.465
+ $X2=3.6 $Y2=2.465
r113 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r114 84 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r115 83 87 8.09112 $w=6.78e-07 $l=4.6e-07 $layer=LI1_cond $X=2.99 $Y=2.465
+ $X2=3.45 $Y2=2.465
r116 83 85 8.21385 $w=6.78e-07 $l=2.5e-08 $layer=LI1_cond $X=2.99 $Y=2.465
+ $X2=2.965 $Y2=2.465
r117 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r118 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r119 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r120 71 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r121 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r122 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r123 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r124 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r125 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r126 62 65 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r127 62 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r128 61 64 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r129 61 91 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=3.725 $Y2=2.72
r130 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r131 58 84 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.99 $Y2=2.72
r132 58 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r133 57 85 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.965 $Y2=2.72
r134 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r135 55 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.21 $Y2=2.72
r136 55 57 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.61 $Y2=2.72
r137 52 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r138 52 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r139 50 70 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.235 $Y=2.72
+ $X2=7.13 $Y2=2.72
r140 50 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.235 $Y=2.72
+ $X2=7.36 $Y2=2.72
r141 49 73 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.485 $Y=2.72
+ $X2=7.59 $Y2=2.72
r142 49 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.485 $Y=2.72
+ $X2=7.36 $Y2=2.72
r143 47 67 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.295 $Y=2.72
+ $X2=6.21 $Y2=2.72
r144 47 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.295 $Y=2.72
+ $X2=6.42 $Y2=2.72
r145 46 70 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=6.545 $Y=2.72
+ $X2=7.13 $Y2=2.72
r146 46 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.545 $Y=2.72
+ $X2=6.42 $Y2=2.72
r147 44 64 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.355 $Y=2.72
+ $X2=5.29 $Y2=2.72
r148 44 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.355 $Y=2.72
+ $X2=5.48 $Y2=2.72
r149 43 67 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=5.605 $Y=2.72
+ $X2=6.21 $Y2=2.72
r150 43 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.605 $Y=2.72
+ $X2=5.48 $Y2=2.72
r151 39 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=2.635
+ $X2=7.36 $Y2=2.72
r152 39 41 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=7.36 $Y=2.635
+ $X2=7.36 $Y2=1.96
r153 35 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=2.72
r154 35 37 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=2.3
r155 31 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2.72
r156 31 33 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2.3
r157 27 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=2.635
+ $X2=1.21 $Y2=2.72
r158 27 29 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.21 $Y=2.635
+ $X2=1.21 $Y2=2.3
r159 26 77 3.97288 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r160 25 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.085 $Y=2.72
+ $X2=1.21 $Y2=2.72
r161 25 26 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.085 $Y=2.72
+ $X2=0.395 $Y2=2.72
r162 21 24 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.27 $Y=1.65
+ $X2=0.27 $Y2=2.33
r163 19 77 3.17028 $w=2.5e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.27 $Y=2.635
+ $X2=0.197 $Y2=2.72
r164 19 24 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.27 $Y=2.635
+ $X2=0.27 $Y2=2.33
r165 6 41 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=7.215
+ $Y=1.485 $X2=7.36 $Y2=1.96
r166 5 37 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=6.275
+ $Y=1.485 $X2=6.42 $Y2=2.3
r167 4 33 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=2.3
r168 3 90 300 $w=1.7e-07 $l=1.09827e-06 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.6 $Y2=2.3
r169 2 29 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.3
r170 1 24 400 $w=1.7e-07 $l=9.05345e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.33
r171 1 21 400 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.65
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_4%A_305_297# 1 2 7 10 15
r20 15 17 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.62 $Y=2.3 $X2=2.62
+ $Y2=2.38
r21 10 12 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=1.68 $Y=2.3 $X2=1.68
+ $Y2=2.38
r22 8 12 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.805 $Y=2.38
+ $X2=1.68 $Y2=2.38
r23 7 17 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.495 $Y=2.38
+ $X2=2.62 $Y2=2.38
r24 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.495 $Y=2.38 $X2=1.805
+ $Y2=2.38
r25 2 15 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.3
r26 1 10 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_4%A_785_297# 1 2 7 10 15
r18 15 17 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=5.01 $Y=2.3 $X2=5.01
+ $Y2=2.38
r19 10 12 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.07 $Y=2.3 $X2=4.07
+ $Y2=2.38
r20 8 12 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.195 $Y=2.38
+ $X2=4.07 $Y2=2.38
r21 7 17 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.885 $Y=2.38
+ $X2=5.01 $Y2=2.38
r22 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.885 $Y=2.38 $X2=4.195
+ $Y2=2.38
r23 2 15 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=2.3
r24 1 10 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_4%X 1 2 3 4 15 19 21 22 23 24 26 27 28 31 35
+ 39 41 43 44 46
c86 27 0 1.27647e-19 $X=6.765 $Y=1.53
r87 45 46 13.5704 $w=5.13e-07 $l=5.4e-07 $layer=LI1_cond $X=7.537 $Y=0.905
+ $X2=7.537 $Y2=1.445
r88 42 43 9.30075 $w=1.75e-07 $l=1.92484e-07 $layer=LI1_cond $X=7.055 $Y=0.82
+ $X2=6.865 $Y2=0.815
r89 41 45 7.89393 $w=1.7e-07 $l=2.10247e-07 $layer=LI1_cond $X=7.365 $Y=0.82
+ $X2=7.537 $Y2=0.905
r90 41 42 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=7.365 $Y=0.82
+ $X2=7.055 $Y2=0.82
r91 40 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.015 $Y=1.53
+ $X2=6.89 $Y2=1.53
r92 39 46 5.28309 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=7.365 $Y=1.53
+ $X2=7.537 $Y2=1.53
r93 39 40 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.365 $Y=1.53
+ $X2=7.015 $Y2=1.53
r94 35 37 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=6.89 $Y=1.62
+ $X2=6.89 $Y2=2.3
r95 33 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=1.615
+ $X2=6.89 $Y2=1.53
r96 33 35 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=6.89 $Y=1.615
+ $X2=6.89 $Y2=1.62
r97 29 43 1.23463 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=6.865 $Y=0.725
+ $X2=6.865 $Y2=0.815
r98 29 31 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.865 $Y=0.725
+ $X2=6.865 $Y2=0.39
r99 27 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.765 $Y=1.53
+ $X2=6.89 $Y2=1.53
r100 27 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.765 $Y=1.53
+ $X2=6.5 $Y2=1.53
r101 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.415 $Y=1.615
+ $X2=6.5 $Y2=1.53
r102 25 26 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.415 $Y=1.615
+ $X2=6.415 $Y2=1.785
r103 23 43 9.30075 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=6.675 $Y=0.815
+ $X2=6.865 $Y2=0.815
r104 23 24 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=6.675 $Y=0.815
+ $X2=6.115 $Y2=0.815
r105 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.33 $Y=1.87
+ $X2=6.415 $Y2=1.785
r106 21 22 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.33 $Y=1.87
+ $X2=6.075 $Y2=1.87
r107 17 22 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=5.97 $Y=1.955
+ $X2=6.075 $Y2=1.87
r108 17 19 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=5.97 $Y=1.955
+ $X2=5.97 $Y2=1.96
r109 13 24 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=5.925 $Y=0.725
+ $X2=6.115 $Y2=0.815
r110 13 15 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.925 $Y=0.725
+ $X2=5.925 $Y2=0.39
r111 4 37 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=2.3
r112 4 35 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=1.62
r113 3 19 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=1.96
r114 2 31 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=6.705
+ $Y=0.235 $X2=6.89 $Y2=0.39
r115 1 15 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=5.765
+ $Y=0.235 $X2=5.95 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_4%A_27_47# 1 2 3 4 13 15 17 21 27 32
c44 21 0 1.62953e-19 $X=1.2 $Y=0.73
r45 25 27 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=2.14 $Y=0.365
+ $X2=3.08 $Y2=0.365
r46 23 32 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=0.365
+ $X2=1.2 $Y2=0.365
r47 23 25 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=1.285 $Y=0.365
+ $X2=2.14 $Y2=0.365
r48 19 32 2.28545 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.2 $Y=0.475 $X2=1.2
+ $Y2=0.365
r49 19 21 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.2 $Y=0.475
+ $X2=1.2 $Y2=0.73
r50 18 30 3.72571 $w=2.2e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=0.365
+ $X2=0.215 $Y2=0.365
r51 17 32 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0.365
+ $X2=1.2 $Y2=0.365
r52 17 18 40.3355 $w=2.18e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=0.365
+ $X2=0.345 $Y2=0.365
r53 13 30 3.15253 $w=2.6e-07 $l=1.1e-07 $layer=LI1_cond $X=0.215 $Y=0.475
+ $X2=0.215 $Y2=0.365
r54 13 15 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.215 $Y=0.475
+ $X2=0.215 $Y2=0.73
r55 4 27 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.945
+ $Y=0.235 $X2=3.08 $Y2=0.38
r56 3 25 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.235 $X2=2.14 $Y2=0.39
r57 2 32 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.39
r58 2 21 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.73
r59 1 30 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
r60 1 15 182 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_4%A_307_47# 1 2 3 4 13 21 23 27 30
r61 25 27 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.985 $Y=0.725
+ $X2=4.985 $Y2=0.39
r62 24 30 5.73815 $w=2.2e-07 $l=1.43614e-07 $layer=LI1_cond $X=4.235 $Y=0.815
+ $X2=4.11 $Y2=0.775
r63 23 25 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=4.795 $Y=0.815
+ $X2=4.985 $Y2=0.725
r64 23 24 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.795 $Y=0.815
+ $X2=4.235 $Y2=0.815
r65 19 30 0.886536 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=4.11 $Y=0.645
+ $X2=4.11 $Y2=0.775
r66 19 21 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=4.11 $Y=0.645
+ $X2=4.11 $Y2=0.42
r67 15 18 41.6652 $w=2.58e-07 $l=9.4e-07 $layer=LI1_cond $X=1.67 $Y=0.775
+ $X2=2.61 $Y2=0.775
r68 13 30 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=3.985 $Y=0.775
+ $X2=4.11 $Y2=0.775
r69 13 18 60.9465 $w=2.58e-07 $l=1.375e-06 $layer=LI1_cond $X=3.985 $Y=0.775
+ $X2=2.61 $Y2=0.775
r70 4 27 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.875
+ $Y=0.235 $X2=5.01 $Y2=0.39
r71 3 30 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=3.935
+ $Y=0.235 $X2=4.07 $Y2=0.76
r72 3 21 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.935
+ $Y=0.235 $X2=4.07 $Y2=0.42
r73 2 18 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=2.61 $Y2=0.73
r74 1 15 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_4%VGND 1 2 3 4 5 18 22 26 30 34 37 38 40 41
+ 43 44 46 47 48 50 69 70 73
r110 73 74 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r111 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r112 67 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=7.59
+ $Y2=0
r113 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r114 64 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r115 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r116 61 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r117 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r118 58 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r119 58 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.45
+ $Y2=0
r120 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r121 55 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.765 $Y=0 $X2=3.6
+ $Y2=0
r122 55 57 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.765 $Y=0
+ $X2=4.37 $Y2=0
r123 50 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.6
+ $Y2=0
r124 50 52 209.096 $w=1.68e-07 $l=3.205e-06 $layer=LI1_cond $X=3.435 $Y=0
+ $X2=0.23 $Y2=0
r125 48 74 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=3.45 $Y2=0
r126 48 52 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r127 46 66 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.275 $Y=0
+ $X2=7.13 $Y2=0
r128 46 47 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=7.275 $Y=0
+ $X2=7.402 $Y2=0
r129 45 69 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=7.53 $Y=0 $X2=7.59
+ $Y2=0
r130 45 47 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=7.53 $Y=0 $X2=7.402
+ $Y2=0
r131 43 63 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.335 $Y=0
+ $X2=6.21 $Y2=0
r132 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.335 $Y=0 $X2=6.42
+ $Y2=0
r133 42 66 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=6.505 $Y=0
+ $X2=7.13 $Y2=0
r134 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.505 $Y=0 $X2=6.42
+ $Y2=0
r135 40 60 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=5.395 $Y=0
+ $X2=5.29 $Y2=0
r136 40 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=0 $X2=5.48
+ $Y2=0
r137 39 63 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=5.565 $Y=0
+ $X2=6.21 $Y2=0
r138 39 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=0 $X2=5.48
+ $Y2=0
r139 37 57 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=0 $X2=4.37
+ $Y2=0
r140 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=0 $X2=4.54
+ $Y2=0
r141 36 60 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.625 $Y=0 $X2=5.29
+ $Y2=0
r142 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=0 $X2=4.54
+ $Y2=0
r143 32 47 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=7.402 $Y=0.085
+ $X2=7.402 $Y2=0
r144 32 34 13.7841 $w=2.53e-07 $l=3.05e-07 $layer=LI1_cond $X=7.402 $Y=0.085
+ $X2=7.402 $Y2=0.39
r145 28 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0
r146 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0.39
r147 24 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0
r148 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.39
r149 20 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0
r150 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0.39
r151 16 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=0.085 $X2=3.6
+ $Y2=0
r152 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.6 $Y=0.085
+ $X2=3.6 $Y2=0.38
r153 5 34 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.225
+ $Y=0.235 $X2=7.36 $Y2=0.39
r154 4 30 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=6.235
+ $Y=0.235 $X2=6.42 $Y2=0.39
r155 3 26 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.345
+ $Y=0.235 $X2=5.48 $Y2=0.39
r156 2 22 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.355
+ $Y=0.235 $X2=4.54 $Y2=0.39
r157 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.475
+ $Y=0.235 $X2=3.6 $Y2=0.38
.ends

