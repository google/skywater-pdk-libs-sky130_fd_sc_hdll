# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__o2bb2ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o2bb2ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295000 1.075000 3.905000 1.285000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.075000 2.025000 1.285000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.845000 1.075000 10.940000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.065000 1.075000 8.675000 1.285000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.608500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.865000 0.645000 6.805000 0.905000 ;
        RECT 4.875000 1.455000 8.465000 1.625000 ;
        RECT 4.875000 1.625000 5.125000 2.465000 ;
        RECT 5.815000 1.625000 6.065000 2.465000 ;
        RECT 6.475000 0.905000 6.805000 1.455000 ;
        RECT 7.275000 1.625000 7.525000 2.125000 ;
        RECT 8.215000 1.625000 8.465000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.085000  0.645000  1.855000 0.905000 ;
      RECT  0.085000  0.905000  0.255000 1.455000 ;
      RECT  0.085000  1.455000  4.315000 1.625000 ;
      RECT  0.100000  0.255000  2.325000 0.475000 ;
      RECT  0.155000  1.795000  0.405000 2.635000 ;
      RECT  0.625000  1.625000  0.875000 2.465000 ;
      RECT  1.095000  1.795000  1.345000 2.635000 ;
      RECT  1.565000  1.625000  1.815000 2.465000 ;
      RECT  2.035000  1.795000  2.285000 2.635000 ;
      RECT  2.075000  0.475000  2.325000 0.725000 ;
      RECT  2.075000  0.725000  4.205000 0.905000 ;
      RECT  2.505000  1.625000  2.755000 2.465000 ;
      RECT  2.545000  0.085000  2.715000 0.555000 ;
      RECT  2.885000  0.255000  3.265000 0.725000 ;
      RECT  2.975000  1.795000  3.225000 2.635000 ;
      RECT  3.445000  1.625000  3.695000 2.465000 ;
      RECT  3.485000  0.085000  3.655000 0.555000 ;
      RECT  3.825000  0.255000  4.205000 0.725000 ;
      RECT  3.915000  1.795000  4.655000 2.635000 ;
      RECT  4.145000  1.075000  6.305000 1.285000 ;
      RECT  4.145000  1.285000  4.315000 1.455000 ;
      RECT  4.460000  0.255000  7.145000 0.475000 ;
      RECT  4.460000  0.475000  4.645000 0.835000 ;
      RECT  5.345000  1.795000  5.595000 2.635000 ;
      RECT  6.285000  1.795000  6.535000 2.635000 ;
      RECT  6.775000  1.795000  7.055000 2.295000 ;
      RECT  6.775000  2.295000  8.935000 2.465000 ;
      RECT  6.975000  0.475000  7.145000 0.735000 ;
      RECT  6.975000  0.735000 10.855000 0.905000 ;
      RECT  7.315000  0.085000  7.485000 0.555000 ;
      RECT  7.655000  0.255000  8.035000 0.725000 ;
      RECT  7.655000  0.725000 10.855000 0.735000 ;
      RECT  7.745000  1.795000  7.995000 2.295000 ;
      RECT  8.255000  0.085000  8.425000 0.555000 ;
      RECT  8.595000  0.255000  8.975000 0.725000 ;
      RECT  8.685000  1.455000 10.875000 1.625000 ;
      RECT  8.685000  1.625000  8.935000 2.295000 ;
      RECT  9.155000  1.795000  9.405000 2.635000 ;
      RECT  9.195000  0.085000  9.365000 0.555000 ;
      RECT  9.535000  0.255000  9.915000 0.725000 ;
      RECT  9.625000  1.625000  9.875000 2.465000 ;
      RECT 10.095000  1.795000 10.345000 2.635000 ;
      RECT 10.135000  0.085000 10.305000 0.555000 ;
      RECT 10.475000  0.255000 10.855000 0.725000 ;
      RECT 10.565000  1.625000 10.875000 2.465000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o2bb2ai_4
END LIBRARY
