* File: sky130_fd_sc_hdll__einvp_4.pex.spice
* Created: Thu Aug 27 19:08:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__EINVP_4%TE 1 3 4 6 7 9 11 12 14 16 17 19 21 22 24
+ 26 27 28 29 30 31
c82 29 0 1.15616e-19 $X=1.95 $Y=1.035
c83 28 0 1.15616e-19 $X=1.48 $Y=1.035
c84 22 0 4.65088e-19 $X=2.345 $Y=1.035
c85 12 0 1.96687e-19 $X=1.405 $Y=1.035
r86 34 36 14.7672 $w=4.08e-07 $l=1.25e-07 $layer=POLY_cond $X=0.35 $Y=1.035
+ $X2=0.35 $Y2=1.16
r87 30 31 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.207 $Y=1.16
+ $X2=0.207 $Y2=1.53
r88 30 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r89 24 26 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.42 $Y=0.96 $X2=2.42
+ $Y2=0.56
r90 23 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.025 $Y=1.035
+ $X2=1.95 $Y2=1.035
r91 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.345 $Y=1.035
+ $X2=2.42 $Y2=0.96
r92 22 23 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.345 $Y=1.035
+ $X2=2.025 $Y2=1.035
r93 19 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.95 $Y=0.96
+ $X2=1.95 $Y2=1.035
r94 19 21 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.95 $Y=0.96 $X2=1.95
+ $Y2=0.56
r95 18 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.555 $Y=1.035
+ $X2=1.48 $Y2=1.035
r96 17 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.875 $Y=1.035
+ $X2=1.95 $Y2=1.035
r97 17 18 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.875 $Y=1.035
+ $X2=1.555 $Y2=1.035
r98 14 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.48 $Y=0.96
+ $X2=1.48 $Y2=1.035
r99 14 16 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.48 $Y=0.96 $X2=1.48
+ $Y2=0.56
r100 13 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.065 $Y=1.035
+ $X2=0.99 $Y2=1.035
r101 12 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.405 $Y=1.035
+ $X2=1.48 $Y2=1.035
r102 12 13 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.405 $Y=1.035
+ $X2=1.065 $Y2=1.035
r103 9 27 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.99 $Y=0.96
+ $X2=0.99 $Y2=1.035
r104 9 11 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.99 $Y=0.96 $X2=0.99
+ $Y2=0.56
r105 8 34 26.3468 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=0.595 $Y=1.035
+ $X2=0.35 $Y2=1.035
r106 7 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.915 $Y=1.035
+ $X2=0.99 $Y2=1.035
r107 7 8 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.915 $Y=1.035
+ $X2=0.595 $Y2=1.035
r108 4 34 29.1132 $w=4.08e-07 $l=2.04083e-07 $layer=POLY_cond $X=0.52 $Y=0.96
+ $X2=0.35 $Y2=1.035
r109 4 6 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.52 $Y=0.96 $X2=0.52
+ $Y2=0.56
r110 1 36 44.8227 $w=4.08e-07 $l=3.14245e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.35 $Y2=1.16
r111 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_4%A_27_47# 1 2 7 9 10 11 12 14 15 17 19 20
+ 22 24 25 26 28 31 35 37 38 40 43 44 54
c115 54 0 1.9418e-19 $X=0.712 $Y=1.16
c116 28 0 1.46731e-19 $X=2.885 $Y=1.395
c117 25 0 9.78995e-20 $X=2.005 $Y=1.395
c118 22 0 1.9667e-19 $X=2.945 $Y=1.47
c119 15 0 1.40591e-19 $X=2.385 $Y=1.395
c120 10 0 7.37965e-20 $X=1.915 $Y=1.395
r121 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.86
+ $Y=1.16 $X2=2.86 $Y2=1.16
r122 41 54 1.39677 $w=3.3e-07 $l=2.13e-07 $layer=LI1_cond $X=0.925 $Y=1.16
+ $X2=0.712 $Y2=1.16
r123 41 43 67.5751 $w=3.28e-07 $l=1.935e-06 $layer=LI1_cond $X=0.925 $Y=1.16
+ $X2=2.86 $Y2=1.16
r124 39 54 5.10169 $w=3.35e-07 $l=1.65e-07 $layer=LI1_cond $X=0.712 $Y=1.325
+ $X2=0.712 $Y2=1.16
r125 39 40 12.4735 $w=4.23e-07 $l=4.6e-07 $layer=LI1_cond $X=0.712 $Y=1.325
+ $X2=0.712 $Y2=1.785
r126 38 54 5.10169 $w=3.35e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.622 $Y=0.995
+ $X2=0.712 $Y2=1.16
r127 37 38 7.99654 $w=2.43e-07 $l=1.7e-07 $layer=LI1_cond $X=0.622 $Y=0.825
+ $X2=0.622 $Y2=0.995
r128 33 40 32.4246 $w=1.68e-07 $l=4.97e-07 $layer=LI1_cond $X=0.215 $Y=1.87
+ $X2=0.712 $Y2=1.87
r129 33 35 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=1.955
+ $X2=0.215 $Y2=2.165
r130 29 37 26.5529 $w=1.68e-07 $l=4.07e-07 $layer=LI1_cond $X=0.215 $Y=0.74
+ $X2=0.622 $Y2=0.74
r131 29 31 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.215 $Y2=0.445
r132 27 44 28.8521 $w=3.2e-07 $l=1.6e-07 $layer=POLY_cond $X=2.885 $Y=1.32
+ $X2=2.885 $Y2=1.16
r133 27 28 13.0992 $w=2.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.885 $Y=1.32
+ $X2=2.885 $Y2=1.395
r134 22 28 13.0992 $w=2.5e-07 $l=1.00623e-07 $layer=POLY_cond $X=2.945 $Y=1.47
+ $X2=2.885 $Y2=1.395
r135 22 24 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.945 $Y=1.47
+ $X2=2.945 $Y2=2.015
r136 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.565 $Y=1.395
+ $X2=2.475 $Y2=1.395
r137 20 28 12.7694 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.725 $Y=1.395
+ $X2=2.885 $Y2=1.395
r138 20 21 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.725 $Y=1.395
+ $X2=2.565 $Y2=1.395
r139 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.475 $Y=1.47
+ $X2=2.475 $Y2=1.395
r140 17 19 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.475 $Y=1.47
+ $X2=2.475 $Y2=2.015
r141 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.095 $Y=1.395
+ $X2=2.005 $Y2=1.395
r142 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.385 $Y=1.395
+ $X2=2.475 $Y2=1.395
r143 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.385 $Y=1.395
+ $X2=2.095 $Y2=1.395
r144 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.005 $Y=1.47
+ $X2=2.005 $Y2=1.395
r145 12 14 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.005 $Y=1.47
+ $X2=2.005 $Y2=2.015
r146 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.915 $Y=1.395
+ $X2=2.005 $Y2=1.395
r147 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.915 $Y=1.395
+ $X2=1.625 $Y2=1.395
r148 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.535 $Y=1.47
+ $X2=1.625 $Y2=1.395
r149 7 9 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=1.535 $Y=1.47
+ $X2=1.535 $Y2=2.015
r150 2 35 600 $w=1.7e-07 $l=7.39865e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.165
r151 1 31 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_4%A 1 3 4 6 7 9 10 12 15 17 19 22 24 26 27
+ 28 29 46 56 60
r73 49 56 10.3946 $w=2.53e-07 $l=2.3e-07 $layer=LI1_cond $X=5.085 $Y=1.147
+ $X2=4.855 $Y2=1.147
r74 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.085
+ $Y=1.16 $X2=5.085 $Y2=1.16
r75 46 48 29.3205 $w=3.37e-07 $l=2.05e-07 $layer=POLY_cond $X=4.88 $Y=1.202
+ $X2=5.085 $Y2=1.202
r76 45 46 3.57567 $w=3.37e-07 $l=2.5e-08 $layer=POLY_cond $X=4.855 $Y=1.202
+ $X2=4.88 $Y2=1.202
r77 43 45 15.7329 $w=3.37e-07 $l=1.1e-07 $layer=POLY_cond $X=4.745 $Y=1.202
+ $X2=4.855 $Y2=1.202
r78 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.745
+ $Y=1.16 $X2=4.745 $Y2=1.16
r79 41 43 47.9139 $w=3.37e-07 $l=3.35e-07 $layer=POLY_cond $X=4.41 $Y=1.202
+ $X2=4.745 $Y2=1.202
r80 40 41 3.57567 $w=3.37e-07 $l=2.5e-08 $layer=POLY_cond $X=4.385 $Y=1.202
+ $X2=4.41 $Y2=1.202
r81 38 40 1.43027 $w=3.37e-07 $l=1e-08 $layer=POLY_cond $X=4.375 $Y=1.202
+ $X2=4.385 $Y2=1.202
r82 36 38 62.2166 $w=3.37e-07 $l=4.35e-07 $layer=POLY_cond $X=3.94 $Y=1.202
+ $X2=4.375 $Y2=1.202
r83 35 36 3.57567 $w=3.37e-07 $l=2.5e-08 $layer=POLY_cond $X=3.915 $Y=1.202
+ $X2=3.94 $Y2=1.202
r84 34 35 63.6469 $w=3.37e-07 $l=4.45e-07 $layer=POLY_cond $X=3.47 $Y=1.202
+ $X2=3.915 $Y2=1.202
r85 33 34 3.57567 $w=3.37e-07 $l=2.5e-08 $layer=POLY_cond $X=3.445 $Y=1.202
+ $X2=3.47 $Y2=1.202
r86 29 60 0.225969 $w=2.53e-07 $l=5e-09 $layer=LI1_cond $X=5.28 $Y=1.147
+ $X2=5.285 $Y2=1.147
r87 29 49 8.8128 $w=2.53e-07 $l=1.95e-07 $layer=LI1_cond $X=5.28 $Y=1.147
+ $X2=5.085 $Y2=1.147
r88 28 56 0.903877 $w=2.53e-07 $l=2e-08 $layer=LI1_cond $X=4.835 $Y=1.147
+ $X2=4.855 $Y2=1.147
r89 28 44 4.06745 $w=2.53e-07 $l=9e-08 $layer=LI1_cond $X=4.835 $Y=1.147
+ $X2=4.745 $Y2=1.147
r90 27 44 18.5295 $w=2.53e-07 $l=4.1e-07 $layer=LI1_cond $X=4.335 $Y=1.147
+ $X2=4.745 $Y2=1.147
r91 27 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.375
+ $Y=1.16 $X2=4.375 $Y2=1.16
r92 24 46 17.4215 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.88 $Y=1.41
+ $X2=4.88 $Y2=1.202
r93 24 26 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.88 $Y=1.41
+ $X2=4.88 $Y2=1.985
r94 20 45 21.7231 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=4.855 $Y=1.015
+ $X2=4.855 $Y2=1.202
r95 20 22 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.855 $Y=1.015
+ $X2=4.855 $Y2=0.56
r96 17 41 17.4215 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.41 $Y=1.41
+ $X2=4.41 $Y2=1.202
r97 17 19 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.41 $Y=1.41
+ $X2=4.41 $Y2=1.985
r98 13 40 21.7231 $w=1.5e-07 $l=1.77e-07 $layer=POLY_cond $X=4.385 $Y=1.025
+ $X2=4.385 $Y2=1.202
r99 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.385 $Y=1.025
+ $X2=4.385 $Y2=0.56
r100 10 36 17.4215 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.94 $Y=1.41
+ $X2=3.94 $Y2=1.202
r101 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.94 $Y=1.41
+ $X2=3.94 $Y2=1.985
r102 7 35 21.7231 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.915 $Y=0.995
+ $X2=3.915 $Y2=1.202
r103 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.915 $Y=0.995
+ $X2=3.915 $Y2=0.56
r104 4 34 17.4215 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.47 $Y=1.41
+ $X2=3.47 $Y2=1.202
r105 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.47 $Y=1.41
+ $X2=3.47 $Y2=1.985
r106 1 33 21.7231 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.445 $Y=0.995
+ $X2=3.445 $Y2=1.202
r107 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.445 $Y=0.995
+ $X2=3.445 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_4%VPWR 1 2 3 12 14 18 22 25 26 27 29 42 43
+ 46 49
r75 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r76 47 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r77 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r78 42 43 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r79 40 43 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=5.29 $Y2=2.72
r80 39 42 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=5.29 $Y2=2.72
r81 39 40 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r82 37 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r83 37 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r84 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r85 34 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=2.72
+ $X2=1.77 $Y2=2.72
r86 34 36 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=1.935 $Y=2.72
+ $X2=2.53 $Y2=2.72
r87 29 46 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.72 $Y2=2.72
r88 29 31 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r89 27 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r90 27 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r91 25 36 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.53 $Y2=2.72
r92 25 26 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.725 $Y2=2.72
r93 24 39 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.905 $Y=2.72
+ $X2=2.99 $Y2=2.72
r94 24 26 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.905 $Y=2.72
+ $X2=2.725 $Y2=2.72
r95 20 26 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=2.635
+ $X2=2.725 $Y2=2.72
r96 20 22 19.6876 $w=3.58e-07 $l=6.15e-07 $layer=LI1_cond $X=2.725 $Y=2.635
+ $X2=2.725 $Y2=2.02
r97 16 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.77 $Y=2.635
+ $X2=1.77 $Y2=2.72
r98 16 18 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.77 $Y=2.635
+ $X2=1.77 $Y2=2.02
r99 15 46 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=0.72 $Y2=2.72
r100 14 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=1.77 $Y2=2.72
r101 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=0.925 $Y2=2.72
r102 10 46 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=2.635
+ $X2=0.72 $Y2=2.72
r103 10 12 8.29197 $w=4.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.72 $Y=2.635
+ $X2=0.72 $Y2=2.34
r104 3 22 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.565
+ $Y=1.545 $X2=2.71 $Y2=2.02
r105 2 18 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.625
+ $Y=1.545 $X2=1.77 $Y2=2.02
r106 1 12 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_4%A_235_309# 1 2 3 4 5 18 20 21 24 26 31 32
+ 33 36 38 40 43 44
c72 43 0 1.97563e-19 $X=2.24 $Y=1.64
c73 26 0 7.0838e-20 $X=3.125 $Y=1.64
c74 20 0 2.31231e-19 $X=2.155 $Y=1.64
r75 40 42 10.7553 $w=3.8e-07 $l=3.35e-07 $layer=LI1_cond $X=5.22 $Y=2.295
+ $X2=5.22 $Y2=1.96
r76 39 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.26 $Y=2.38
+ $X2=4.175 $Y2=2.38
r77 38 40 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=5.03 $Y=2.38
+ $X2=5.22 $Y2=2.295
r78 38 39 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.03 $Y=2.38
+ $X2=4.26 $Y2=2.38
r79 34 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.175 $Y=2.295
+ $X2=4.175 $Y2=2.38
r80 34 36 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.175 $Y=2.295
+ $X2=4.175 $Y2=1.96
r81 32 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.09 $Y=2.38
+ $X2=4.175 $Y2=2.38
r82 32 33 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=4.09 $Y=2.38
+ $X2=3.295 $Y2=2.38
r83 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.21 $Y=2.295
+ $X2=3.295 $Y2=2.38
r84 29 31 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.21 $Y=2.295
+ $X2=3.21 $Y2=1.96
r85 28 31 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.21 $Y=1.725
+ $X2=3.21 $Y2=1.96
r86 27 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.325 $Y=1.64
+ $X2=2.24 $Y2=1.64
r87 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.125 $Y=1.64
+ $X2=3.21 $Y2=1.725
r88 26 27 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.125 $Y=1.64
+ $X2=2.325 $Y2=1.64
r89 22 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=1.725
+ $X2=2.24 $Y2=1.64
r90 22 24 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.24 $Y=1.725
+ $X2=2.24 $Y2=1.96
r91 20 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=1.64
+ $X2=2.24 $Y2=1.64
r92 20 21 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.155 $Y=1.64
+ $X2=1.385 $Y2=1.64
r93 16 21 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.28 $Y=1.725
+ $X2=1.385 $Y2=1.64
r94 16 18 27.1991 $w=2.08e-07 $l=5.15e-07 $layer=LI1_cond $X=1.28 $Y=1.725
+ $X2=1.28 $Y2=2.24
r95 5 42 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.97
+ $Y=1.485 $X2=5.115 $Y2=1.96
r96 4 36 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.03
+ $Y=1.485 $X2=4.175 $Y2=1.96
r97 3 31 300 $w=1.7e-07 $l=4.94823e-07 $layer=licon1_PDIFF $count=2 $X=3.035
+ $Y=1.545 $X2=3.21 $Y2=1.96
r98 2 24 300 $w=1.7e-07 $l=4.82079e-07 $layer=licon1_PDIFF $count=2 $X=2.095
+ $Y=1.545 $X2=2.24 $Y2=1.96
r99 1 18 600 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_PDIFF $count=1 $X=1.175
+ $Y=1.545 $X2=1.3 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_4%Z 1 2 3 4 15 19 21 22 23 24 25 44 48
c56 48 0 1.9667e-19 $X=3.805 $Y=1.87
c57 24 0 1.46731e-19 $X=3.825 $Y=1.53
r58 45 48 2.93156 $w=5.08e-07 $l=1.25e-07 $layer=LI1_cond $X=3.68 $Y=1.87
+ $X2=3.805 $Y2=1.87
r59 45 46 2.46227 $w=3.8e-07 $l=2.55e-07 $layer=LI1_cond $X=3.68 $Y=1.87
+ $X2=3.68 $Y2=1.615
r60 25 44 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.335 $Y=1.53
+ $X2=4.35 $Y2=1.53
r61 25 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.335 $Y=1.53
+ $X2=4.03 $Y2=1.53
r62 24 41 5.07913 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=3.76 $Y=1.53 $X2=4.03
+ $Y2=1.53
r63 24 46 2.1225 $w=4.6e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.76 $Y=1.53
+ $X2=3.68 $Y2=1.615
r64 24 48 9.00371 $w=1.3e-07 $l=2.55e-07 $layer=LI1_cond $X=3.805 $Y=1.615
+ $X2=3.805 $Y2=1.87
r65 23 24 5.01049 $w=7.08e-07 $l=2.55e-07 $layer=LI1_cond $X=3.76 $Y=1.19
+ $X2=3.76 $Y2=1.445
r66 22 23 6.60058 $w=5.38e-07 $l=2.98e-07 $layer=LI1_cond $X=3.76 $Y=0.892
+ $X2=3.76 $Y2=1.19
r67 19 44 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=4.43 $Y=1.53 $X2=4.35
+ $Y2=1.53
r68 19 21 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.43 $Y=1.53 $X2=4.62
+ $Y2=1.53
r69 13 22 6.14688 $w=2.15e-07 $l=2.7e-07 $layer=LI1_cond $X=4.03 $Y=0.742
+ $X2=3.76 $Y2=0.742
r70 13 15 32.9652 $w=2.13e-07 $l=6.15e-07 $layer=LI1_cond $X=4.03 $Y=0.742
+ $X2=4.645 $Y2=0.742
r71 4 21 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=4.5
+ $Y=1.485 $X2=4.645 $Y2=1.61
r72 3 24 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=3.56
+ $Y=1.485 $X2=3.705 $Y2=1.61
r73 2 15 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=4.46
+ $Y=0.235 $X2=4.645 $Y2=0.76
r74 1 22 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=3.52
+ $Y=0.235 $X2=3.705 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_4%VGND 1 2 3 12 16 20 22 24 29 34 44 45 48
+ 51 54
r77 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r78 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r79 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r80 44 45 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r81 42 45 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.99 $Y=0 $X2=5.29
+ $Y2=0
r82 42 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r83 41 44 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.99 $Y=0 $X2=5.29
+ $Y2=0
r84 41 42 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r85 39 54 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.805 $Y=0 $X2=2.61
+ $Y2=0
r86 39 41 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.805 $Y=0 $X2=2.99
+ $Y2=0
r87 38 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r88 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r89 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r90 35 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.665
+ $Y2=0
r91 35 37 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=2.07
+ $Y2=0
r92 34 54 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=2.61
+ $Y2=0
r93 34 37 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=2.07
+ $Y2=0
r94 33 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r95 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r96 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r97 30 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r98 30 32 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.15
+ $Y2=0
r99 29 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.665
+ $Y2=0
r100 29 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.475 $Y=0
+ $X2=1.15 $Y2=0
r101 24 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r102 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r103 22 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r104 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r105 18 54 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0
r106 18 20 8.1262 $w=3.88e-07 $l=2.75e-07 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0.36
r107 14 51 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=0.085
+ $X2=1.665 $Y2=0
r108 14 16 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=1.665 $Y=0.085
+ $X2=1.665 $Y2=0.36
r109 10 48 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r110 10 12 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.36
r111 3 20 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.495
+ $Y=0.235 $X2=2.63 $Y2=0.36
r112 2 16 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.235 $X2=1.69 $Y2=0.36
r113 1 12 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_4%A_213_47# 1 2 3 4 5 18 20 21 24 26 31 32
+ 36 38
c61 38 0 9.78995e-20 $X=2.16 $Y=0.74
c62 26 0 3.37278e-19 $X=2.985 $Y=0.74
c63 20 0 2.70484e-19 $X=2.075 $Y=0.74
r64 34 36 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=4.175 $Y=0.36
+ $X2=5.115 $Y2=0.36
r65 32 34 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=3.32 $Y=0.36
+ $X2=4.175 $Y2=0.36
r66 29 31 4.12815 $w=3.33e-07 $l=1.2e-07 $layer=LI1_cond $X=3.152 $Y=0.655
+ $X2=3.152 $Y2=0.535
r67 28 32 7.29352 $w=2.1e-07 $l=2.14159e-07 $layer=LI1_cond $X=3.152 $Y=0.465
+ $X2=3.32 $Y2=0.36
r68 28 31 2.40809 $w=3.33e-07 $l=7e-08 $layer=LI1_cond $X=3.152 $Y=0.465
+ $X2=3.152 $Y2=0.535
r69 27 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0.74
+ $X2=2.16 $Y2=0.74
r70 26 29 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=2.985 $Y=0.74
+ $X2=3.152 $Y2=0.655
r71 26 27 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.985 $Y=0.74
+ $X2=2.245 $Y2=0.74
r72 22 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.655
+ $X2=2.16 $Y2=0.74
r73 22 24 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.16 $Y=0.655
+ $X2=2.16 $Y2=0.535
r74 20 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0.74
+ $X2=2.16 $Y2=0.74
r75 20 21 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.075 $Y=0.74
+ $X2=1.305 $Y2=0.74
r76 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.22 $Y=0.655
+ $X2=1.305 $Y2=0.74
r77 16 18 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.22 $Y=0.655
+ $X2=1.22 $Y2=0.535
r78 5 36 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=4.93
+ $Y=0.235 $X2=5.115 $Y2=0.36
r79 4 34 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.235 $X2=4.175 $Y2=0.36
r80 3 31 182 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_NDIFF $count=1 $X=3.11
+ $Y=0.235 $X2=3.235 $Y2=0.535
r81 2 24 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.16 $Y2=0.535
r82 1 18 182 $w=1.7e-07 $l=3.69459e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.22 $Y2=0.535
.ends

