* File: sky130_fd_sc_hdll__clkmux2_2.pex.spice
* Created: Wed Sep  2 08:27:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_2%A_79_199# 1 2 7 9 12 16 18 20 23 26 27
+ 29 32 34 38 40 44
c98 40 0 1.9931e-19 $X=1.982 $Y=0.54
c99 38 0 1.80039e-19 $X=3.13 $Y=2.04
r100 43 44 4.53495 $w=3.72e-07 $l=3.5e-08 $layer=POLY_cond $X=0.93 $Y=1.202
+ $X2=0.965 $Y2=1.202
r101 42 43 54.4194 $w=3.72e-07 $l=4.2e-07 $layer=POLY_cond $X=0.51 $Y=1.202
+ $X2=0.93 $Y2=1.202
r102 41 42 1.94355 $w=3.72e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.51 $Y2=1.202
r103 36 38 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.415 $Y=2.04
+ $X2=3.13 $Y2=2.04
r104 34 36 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.07 $Y=2.04
+ $X2=2.415 $Y2=2.04
r105 30 40 3.49088 $w=2.67e-07 $l=1.4026e-07 $layer=LI1_cond $X=2.07 $Y=0.437
+ $X2=1.982 $Y2=0.54
r106 30 32 13.4189 $w=3.63e-07 $l=4.25e-07 $layer=LI1_cond $X=2.07 $Y=0.437
+ $X2=2.495 $Y2=0.437
r107 29 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.985 $Y=1.955
+ $X2=2.07 $Y2=2.04
r108 28 40 3.01551 $w=1.7e-07 $l=2.86496e-07 $layer=LI1_cond $X=1.985 $Y=0.825
+ $X2=1.982 $Y2=0.54
r109 28 29 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=1.985 $Y=0.825
+ $X2=1.985 $Y2=1.955
r110 26 40 3.49088 $w=2.67e-07 $l=2.39583e-07 $layer=LI1_cond $X=1.895 $Y=0.74
+ $X2=1.982 $Y2=0.54
r111 26 27 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.895 $Y=0.74
+ $X2=1.145 $Y2=0.74
r112 24 44 12.3091 $w=3.72e-07 $l=9.5e-08 $layer=POLY_cond $X=1.06 $Y=1.202
+ $X2=0.965 $Y2=1.202
r113 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.06
+ $Y=1.16 $X2=1.06 $Y2=1.16
r114 21 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.06 $Y=0.825
+ $X2=1.145 $Y2=0.74
r115 21 23 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.06 $Y=0.825
+ $X2=1.06 $Y2=1.16
r116 18 44 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r117 18 20 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r118 14 43 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.93 $Y=0.995
+ $X2=0.93 $Y2=1.202
r119 14 16 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.93 $Y=0.995
+ $X2=0.93 $Y2=0.495
r120 10 42 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.51 $Y=0.995
+ $X2=0.51 $Y2=1.202
r121 10 12 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.51 $Y=0.995
+ $X2=0.51 $Y2=0.495
r122 7 41 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r123 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r124 2 38 400 $w=1.7e-07 $l=1.07949e-06 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.545 $X2=3.13 $Y2=2.04
r125 2 36 400 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.545 $X2=2.415 $Y2=2.04
r126 1 32 182 $w=1.7e-07 $l=3.94968e-07 $layer=licon1_NDIFF $count=1 $X=2.195
+ $Y=0.235 $X2=2.495 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_2%S 1 3 6 8 10 13 16 17 18 19 20 21 23 27
+ 31 32
c95 16 0 1.20839e-19 $X=1.63 $Y=2.295
r96 31 32 13.2166 $w=3.58e-07 $l=3.33e-07 $layer=LI1_cond $X=3.932 $Y=1.535
+ $X2=4.265 $Y2=1.535
r97 27 30 7.79239 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.592 $Y=1.16
+ $X2=1.592 $Y2=1.325
r98 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.54
+ $Y=1.16 $X2=1.54 $Y2=1.16
r99 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.35
+ $Y=1.22 $X2=4.35 $Y2=1.22
r100 21 32 3.40825 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=4.36 $Y=1.44
+ $X2=4.36 $Y2=1.535
r101 21 23 12.8421 $w=1.88e-07 $l=2.2e-07 $layer=LI1_cond $X=4.36 $Y=1.44
+ $X2=4.36 $Y2=1.22
r102 19 31 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.79 $Y=1.63
+ $X2=3.79 $Y2=1.535
r103 19 20 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.79 $Y=1.63
+ $X2=3.79 $Y2=2.295
r104 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.705 $Y=2.38
+ $X2=3.79 $Y2=2.295
r105 17 18 128.85 $w=1.68e-07 $l=1.975e-06 $layer=LI1_cond $X=3.705 $Y=2.38
+ $X2=1.73 $Y2=2.38
r106 16 18 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.63 $Y=2.295
+ $X2=1.73 $Y2=2.38
r107 16 30 53.7909 $w=1.98e-07 $l=9.7e-07 $layer=LI1_cond $X=1.63 $Y=2.295
+ $X2=1.63 $Y2=1.325
r108 11 24 39.2931 $w=2.55e-07 $l=1.88348e-07 $layer=POLY_cond $X=4.4 $Y=1.055
+ $X2=4.35 $Y2=1.22
r109 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.4 $Y=1.055
+ $X2=4.4 $Y2=0.495
r110 8 24 51.486 $w=2.55e-07 $l=2.62202e-07 $layer=POLY_cond $X=4.375 $Y=1.47
+ $X2=4.35 $Y2=1.22
r111 8 10 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=4.375 $Y=1.47
+ $X2=4.375 $Y2=2.015
r112 4 28 39.2931 $w=2.55e-07 $l=1.94808e-07 $layer=POLY_cond $X=1.61 $Y=0.995
+ $X2=1.545 $Y2=1.16
r113 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.61 $Y=0.995
+ $X2=1.61 $Y2=0.445
r114 1 28 62.8272 $w=2.55e-07 $l=3.29393e-07 $layer=POLY_cond $X=1.585 $Y=1.47
+ $X2=1.545 $Y2=1.16
r115 1 3 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=1.585 $Y=1.47
+ $X2=1.585 $Y2=2.015
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_2%A1 3 5 7 10 11 13 14 16 17
c69 5 0 1.3232e-19 $X=3.365 $Y=1.47
r70 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.33
+ $Y=1.22 $X2=3.33 $Y2=1.22
r71 17 26 1.19218 $w=2.88e-07 $l=3e-08 $layer=LI1_cond $X=3.39 $Y=1.19 $X2=3.39
+ $Y2=1.22
r72 16 17 13.5114 $w=2.88e-07 $l=3.4e-07 $layer=LI1_cond $X=3.39 $Y=0.85
+ $X2=3.39 $Y2=1.19
r73 15 26 15.6971 $w=2.88e-07 $l=3.95e-07 $layer=LI1_cond $X=3.39 $Y=1.615
+ $X2=3.39 $Y2=1.22
r74 13 15 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=3.245 $Y=1.7
+ $X2=3.39 $Y2=1.615
r75 13 14 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=3.245 $Y=1.7
+ $X2=2.41 $Y2=1.7
r76 11 20 45.5456 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=2.325 $Y=0.975
+ $X2=2.12 $Y2=0.975
r77 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.325
+ $Y=0.975 $X2=2.325 $Y2=0.975
r78 8 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.325 $Y=1.615
+ $X2=2.41 $Y2=1.7
r79 8 10 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.325 $Y=1.615
+ $X2=2.325 $Y2=0.975
r80 5 25 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.365 $Y=1.47
+ $X2=3.33 $Y2=1.22
r81 5 7 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=3.365 $Y=1.47
+ $X2=3.365 $Y2=2.015
r82 1 20 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.12 $Y=0.84
+ $X2=2.12 $Y2=0.975
r83 1 3 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.12 $Y=0.84 $X2=2.12
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_2%A0 1 3 4 5 8 11 12 15 16
c50 1 0 1.20839e-19 $X=2.18 $Y=1.47
r51 15 18 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=0.98
+ $X2=2.835 $Y2=1.145
r52 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=0.98
+ $X2=2.835 $Y2=0.815
r53 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.835
+ $Y=0.98 $X2=2.835 $Y2=0.98
r54 12 16 7.44655 $w=3.23e-07 $l=2.1e-07 $layer=LI1_cond $X=2.912 $Y=1.19
+ $X2=2.912 $Y2=0.98
r55 11 18 58.026 $w=2e-07 $l=1.75e-07 $layer=POLY_cond $X=2.8 $Y=1.32 $X2=2.8
+ $Y2=1.145
r56 8 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.775 $Y=0.445
+ $X2=2.775 $Y2=0.815
r57 4 11 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=2.7 $Y=1.395
+ $X2=2.8 $Y2=1.32
r58 4 5 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.7 $Y=1.395 $X2=2.27
+ $Y2=1.395
r59 1 5 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.18 $Y=1.47
+ $X2=2.27 $Y2=1.395
r60 1 3 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.18 $Y=1.47 $X2=2.18
+ $Y2=2.015
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_2%A_741_21# 1 2 9 12 13 15 18 19 21 22 27
+ 32 33 34
c68 18 0 1.3232e-19 $X=3.87 $Y=1.02
c69 13 0 1.80039e-19 $X=3.805 $Y=1.47
c70 9 0 1.95128e-19 $X=3.78 $Y=0.445
r71 32 33 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=4.645 $Y=2
+ $X2=4.645 $Y2=1.835
r72 29 34 4.36305 $w=2.07e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.76 $Y=0.865
+ $X2=4.67 $Y2=0.78
r73 29 33 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=4.76 $Y=0.865
+ $X2=4.76 $Y2=1.835
r74 25 34 4.36305 $w=2.07e-07 $l=1.08305e-07 $layer=LI1_cond $X=4.617 $Y=0.695
+ $X2=4.67 $Y2=0.78
r75 25 27 11.2892 $w=2.43e-07 $l=2.4e-07 $layer=LI1_cond $X=4.617 $Y=0.695
+ $X2=4.617 $Y2=0.455
r76 21 34 2.06925 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=4.495 $Y=0.78
+ $X2=4.67 $Y2=0.78
r77 21 22 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.495 $Y=0.78
+ $X2=3.955 $Y2=0.78
r78 19 37 39.6736 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.855 $Y=1.02
+ $X2=3.855 $Y2=1.185
r79 19 36 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.855 $Y=1.02
+ $X2=3.855 $Y2=0.855
r80 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.87
+ $Y=1.02 $X2=3.87 $Y2=1.02
r81 16 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.87 $Y=0.865
+ $X2=3.955 $Y2=0.78
r82 16 18 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.87 $Y=0.865
+ $X2=3.87 $Y2=1.02
r83 13 15 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=3.805 $Y=1.47
+ $X2=3.805 $Y2=2.015
r84 12 13 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.805 $Y=1.37 $X2=3.805
+ $Y2=1.47
r85 12 37 61.3418 $w=2e-07 $l=1.85e-07 $layer=POLY_cond $X=3.805 $Y=1.37
+ $X2=3.805 $Y2=1.185
r86 9 36 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.78 $Y=0.445
+ $X2=3.78 $Y2=0.855
r87 2 32 300 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=2 $X=4.465
+ $Y=1.545 $X2=4.61 $Y2=2
r88 1 27 182 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_NDIFF $count=1 $X=4.475
+ $Y=0.235 $X2=4.61 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_2%VPWR 1 2 3 10 12 16 20 26 29 30 31 41 42
+ 48
r52 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r53 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r54 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r55 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r56 38 39 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r57 36 39 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=3.91 $Y2=2.72
r58 36 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r59 35 38 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=3.91 $Y2=2.72
r60 35 36 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r61 33 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.325 $Y=2.72
+ $X2=1.2 $Y2=2.72
r62 33 35 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.325 $Y=2.72
+ $X2=1.61 $Y2=2.72
r63 31 49 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.695 $Y=2.72
+ $X2=1.15 $Y2=2.72
r64 31 46 0.132312 $w=4.8e-07 $l=4.65e-07 $layer=MET1_cond $X=0.695 $Y=2.72
+ $X2=0.23 $Y2=2.72
r65 29 38 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.045 $Y=2.72
+ $X2=3.91 $Y2=2.72
r66 29 30 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.045 $Y=2.72
+ $X2=4.16 $Y2=2.72
r67 28 41 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=4.275 $Y=2.72
+ $X2=4.83 $Y2=2.72
r68 28 30 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.275 $Y=2.72
+ $X2=4.16 $Y2=2.72
r69 24 30 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.16 $Y=2.635
+ $X2=4.16 $Y2=2.72
r70 24 26 31.8174 $w=2.28e-07 $l=6.35e-07 $layer=LI1_cond $X=4.16 $Y=2.635
+ $X2=4.16 $Y2=2
r71 20 23 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=1.2 $Y=1.66 $X2=1.2
+ $Y2=2.34
r72 18 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.72
r73 18 23 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.34
r74 17 45 3.95006 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=2.72 $X2=0.19
+ $Y2=2.72
r75 16 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.075 $Y=2.72
+ $X2=1.2 $Y2=2.72
r76 16 17 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.075 $Y=2.72
+ $X2=0.38 $Y2=2.72
r77 12 15 31.9862 $w=2.43e-07 $l=6.8e-07 $layer=LI1_cond $X=0.257 $Y=1.66
+ $X2=0.257 $Y2=2.34
r78 10 45 3.16005 $w=2.45e-07 $l=1.13666e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.19 $Y2=2.72
r79 10 15 13.8764 $w=2.43e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.257 $Y2=2.34
r80 3 26 300 $w=1.7e-07 $l=5.60312e-07 $layer=licon1_PDIFF $count=2 $X=3.895
+ $Y=1.545 $X2=4.13 $Y2=2
r81 2 23 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.34
r82 2 20 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.66
r83 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r84 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_2%X 1 2 10 12 13 14
r20 14 27 4.4064 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=0.725 $Y=2.21
+ $X2=0.725 $Y2=2.34
r21 13 14 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.725 $Y=1.87
+ $X2=0.725 $Y2=2.21
r22 11 12 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=0.68 $Y=1.495
+ $X2=0.68 $Y2=0.475
r23 10 11 6.42278 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.66
+ $X2=0.725 $Y2=1.495
r24 8 13 6.94855 $w=3.38e-07 $l=2.05e-07 $layer=LI1_cond $X=0.725 $Y=1.665
+ $X2=0.725 $Y2=1.87
r25 8 10 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=1.665
+ $X2=0.725 $Y2=1.66
r26 2 27 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r27 2 10 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r28 1 12 182 $w=1.7e-07 $l=3e-07 $layer=licon1_NDIFF $count=1 $X=0.585 $Y=0.235
+ $X2=0.72 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_2%VGND 1 2 3 10 12 16 18 20 25 35 36 42
c62 25 0 1.95128e-19 $X=3.71 $Y=0
r63 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r64 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r65 36 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=3.91
+ $Y2=0
r66 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r67 33 35 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.225 $Y=0 $X2=4.83
+ $Y2=0
r68 32 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r69 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r70 29 32 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=3.45
+ $Y2=0
r71 29 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r72 28 31 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=3.45
+ $Y2=0
r73 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r74 26 42 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.165
+ $Y2=0
r75 26 28 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.61
+ $Y2=0
r76 25 49 8.36094 $w=5.13e-07 $l=3.6e-07 $layer=LI1_cond $X=3.967 $Y=0 $X2=3.967
+ $Y2=0.36
r77 25 33 7.34265 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=3.967 $Y=0 $X2=4.225
+ $Y2=0
r78 25 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r79 25 31 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.71 $Y=0 $X2=3.45
+ $Y2=0
r80 21 39 3.98448 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.192
+ $Y2=0
r81 21 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.69
+ $Y2=0
r82 20 42 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.165
+ $Y2=0
r83 20 23 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.69
+ $Y2=0
r84 18 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r85 18 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r86 18 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r87 14 42 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.165 $Y=0.085
+ $X2=1.165 $Y2=0
r88 14 16 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=1.165 $Y=0.085
+ $X2=1.165 $Y2=0.38
r89 10 39 3.15868 $w=2.5e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.192 $Y2=0
r90 10 12 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.49
r91 3 49 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=3.855
+ $Y=0.235 $X2=4.09 $Y2=0.36
r92 2 16 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.235 $X2=1.19 $Y2=0.38
r93 1 12 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.49
.ends

