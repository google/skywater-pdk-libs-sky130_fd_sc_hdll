* File: sky130_fd_sc_hdll__sdlclkp_4.spice
* Created: Wed Sep  2 08:52:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__sdlclkp_4.pex.spice"
.subckt sky130_fd_sc_hdll__sdlclkp_4  VNB VPB SCE GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1016 N_VGND_M1016_d N_SCE_M1016_g N_A_27_47#_M1016_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1001 N_A_27_47#_M1001_d N_GATE_M1001_g N_VGND_M1016_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0733385 AS=0.0672 PD=0.813077 PS=0.74 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1026 N_A_310_47#_M1026_d N_A_280_21#_M1026_g N_A_27_47#_M1001_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0765 AS=0.0628615 PD=0.785 PS=0.696923 NRD=31.656
+ NRS=19.992 M=1 R=2.4 SA=75001.2 SB=75002.1 A=0.054 P=1.02 MULT=1
MM1000 A_425_47# N_A_277_243#_M1000_g N_A_310_47#_M1026_d VNB NSHORT L=0.15
+ W=0.36 AD=0.101354 AS=0.0765 PD=0.904615 PS=0.785 NRD=75.504 NRS=16.656 M=1
+ R=2.4 SA=75001.8 SB=75001.5 A=0.054 P=1.02 MULT=1
MM1015 N_VGND_M1015_d N_A_505_315#_M1015_g A_425_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.120799 AS=0.118246 PD=0.902804 PS=1.05538 NRD=25.704 NRS=64.716 M=1 R=2.8
+ SA=75002.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1027 N_A_505_315#_M1027_d N_A_310_47#_M1027_g N_VGND_M1015_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.186951 PD=1.82 PS=1.3972 NRD=0 NRS=23.988 M=1 R=4.33333
+ SA=75001.9 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A_280_21#_M1008_g N_A_277_243#_M1008_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1006 N_A_280_21#_M1006_d N_CLK_M1006_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0672 PD=1.36 PS=0.74 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 A_1217_47# N_A_505_315#_M1018_g N_A_1125_47#_M1018_s VNB NSHORT L=0.15
+ W=0.65 AD=0.06825 AS=0.2015 PD=0.86 PS=1.92 NRD=9.228 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1021_d N_CLK_M1021_g A_1217_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.141375 AS=0.06825 PD=1.085 PS=0.86 NRD=14.76 NRS=9.228 M=1 R=4.33333
+ SA=75000.6 SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1004 N_GCLK_M1004_d N_A_1125_47#_M1004_g N_VGND_M1021_d VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.141375 PD=0.97 PS=1.085 NRD=8.304 NRS=13.836 M=1
+ R=4.33333 SA=75001.2 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1014 N_GCLK_M1004_d N_A_1125_47#_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.6 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1022 N_GCLK_M1022_d N_A_1125_47#_M1022_g N_VGND_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.164125 AS=0.104 PD=1.155 PS=0.97 NRD=33.228 NRS=0 M=1 R=4.33333
+ SA=75002.1 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1024 N_GCLK_M1022_d N_A_1125_47#_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15
+ W=0.65 AD=0.164125 AS=0.2405 PD=1.155 PS=2.04 NRD=8.304 NRS=15.684 M=1
+ R=4.33333 SA=75002.8 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1007 A_117_369# N_SCE_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0736 AS=0.1728 PD=0.87 PS=1.82 NRD=18.4589 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90002.2 A=0.1152 P=1.64 MULT=1
MM1002 N_A_27_47#_M1002_d N_GATE_M1002_g A_117_369# VPB PHIGHVT L=0.18 W=0.64
+ AD=0.143275 AS=0.0736 PD=1.25585 PS=0.87 NRD=18.4589 NRS=18.4589 M=1 R=3.55556
+ SA=90000.6 SB=90001.8 A=0.1152 P=1.64 MULT=1
MM1012 N_A_310_47#_M1012_d N_A_277_243#_M1012_g N_A_27_47#_M1002_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.0735 AS=0.0940245 PD=0.77 PS=0.824151 NRD=16.4101
+ NRS=28.1316 M=1 R=2.33333 SA=90001.2 SB=90002.1 A=0.0756 P=1.2 MULT=1
MM1005 A_421_413# N_A_280_21#_M1005_g N_A_310_47#_M1012_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0903 AS=0.0735 PD=0.85 PS=0.77 NRD=75.0373 NRS=16.4101 M=1
+ R=2.33333 SA=90001.7 SB=90001.5 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_A_505_315#_M1010_g A_421_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.116654 AS=0.0903 PD=0.934648 PS=0.85 NRD=89.1031 NRS=75.0373 M=1
+ R=2.33333 SA=90002.3 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1019 N_A_505_315#_M1019_d N_A_310_47#_M1019_g N_VPWR_M1010_d VPB PHIGHVT
+ L=0.18 W=1 AD=0.27 AS=0.277746 PD=2.54 PS=2.22535 NRD=0.9653 NRS=21.67 M=1
+ R=5.55556 SA=90001.4 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1013_d N_A_280_21#_M1013_g N_A_277_243#_M1013_s VPB PHIGHVT
+ L=0.18 W=0.64 AD=0.17565 AS=0.1728 PD=1.39 PS=1.82 NRD=67.5316 NRS=1.5366 M=1
+ R=3.55556 SA=90000.2 SB=90000.8 A=0.1152 P=1.64 MULT=1
MM1023 N_A_280_21#_M1023_d N_CLK_M1023_g N_VPWR_M1013_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.17565 PD=1.82 PS=1.39 NRD=1.5366 NRS=67.5316 M=1
+ R=3.55556 SA=90000.8 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1011 N_A_1125_47#_M1011_d N_A_505_315#_M1011_g N_VPWR_M1011_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.2 SB=90002.8 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_CLK_M1009_g N_A_1125_47#_M1011_d VPB PHIGHVT L=0.18 W=1
+ AD=0.1725 AS=0.145 PD=1.345 PS=1.29 NRD=6.8753 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90002.4 A=0.18 P=2.36 MULT=1
MM1003 N_GCLK_M1003_d N_A_1125_47#_M1003_g N_VPWR_M1009_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.1725 PD=1.29 PS=1.345 NRD=0.9653 NRS=5.8903 M=1 R=5.55556
+ SA=90001.2 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1017 N_GCLK_M1003_d N_A_1125_47#_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.7 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1020 N_GCLK_M1020_d N_A_1125_47#_M1020_g N_VPWR_M1017_s VPB PHIGHVT L=0.18 W=1
+ AD=0.2125 AS=0.145 PD=1.425 PS=1.29 NRD=27.5603 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1025 N_GCLK_M1020_d N_A_1125_47#_M1025_g N_VPWR_M1025_s VPB PHIGHVT L=0.18 W=1
+ AD=0.2125 AS=0.38 PD=1.425 PS=2.76 NRD=0.9653 NRS=18.715 M=1 R=5.55556
+ SA=90002.7 SB=90000.3 A=0.18 P=2.36 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.3759 P=22.37
c_83 VNB 0 2.53617e-19 $X=0.15 $Y=-0.085
c_156 VPB 0 1.12975e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__sdlclkp_4.pxi.spice"
*
.ends
*
*
