* File: sky130_fd_sc_hdll__inputiso0n_1.spice
* Created: Thu Aug 27 19:08:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__inputiso0n_1.pex.spice"
.subckt sky130_fd_sc_hdll__inputiso0n_1  VNB VPB A SLEEP_B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* SLEEP_B	SLEEP_B
* A	A
* VPB	VPB
* VNB	VNB
MM1005 A_123_75# N_A_M1005_g N_A_27_75#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1386 PD=0.69 PS=1.5 NRD=22.848 NRS=12.852 M=1 R=2.8 SA=75000.3
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_SLEEP_B_M1003_g A_123_75# VNB NSHORT L=0.15 W=0.42
+ AD=0.0960112 AS=0.0567 PD=0.855701 PS=0.69 NRD=48.564 NRS=22.848 M=1 R=2.8
+ SA=75000.7 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_27_75#_M1001_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.148589 PD=1.82 PS=1.3243 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_27_75#_M1002_d N_A_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0609 AS=0.1218 PD=0.71 PS=1.42 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1004 N_VPWR_M1004_d N_SLEEP_B_M1004_g N_A_27_75#_M1002_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.102723 AS=0.0609 PD=0.834085 PS=0.71 NRD=59.7895 NRS=2.3443 M=1
+ R=2.33333 SA=90000.7 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1000 N_X_M1000_d N_A_27_75#_M1000_g N_VPWR_M1004_d VPB PHIGHVT L=0.18 W=1
+ AD=0.37 AS=0.244577 PD=2.74 PS=1.98592 NRD=20.685 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90000.3 A=0.18 P=2.36 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
*
.include "sky130_fd_sc_hdll__inputiso0n_1.pxi.spice"
*
.ends
*
*
