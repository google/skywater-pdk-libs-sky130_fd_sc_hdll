* File: sky130_fd_sc_hdll__clkinv_16.spice
* Created: Thu Aug 27 19:02:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__clkinv_16.pex.spice"
.subckt sky130_fd_sc_hdll__clkinv_16  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.1113 PD=0.75 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75007.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_Y_M1000_d N_A_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0693 PD=0.75 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.7 SB=75007.1
+ A=0.063 P=1.14 MULT=1
MM1008 N_Y_M1008_d N_A_M1008_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.1 SB=75006.7
+ A=0.063 P=1.14 MULT=1
MM1010 N_Y_M1008_d N_A_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0693 PD=0.75 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.6 SB=75006.2
+ A=0.063 P=1.14 MULT=1
MM1011 N_Y_M1011_d N_A_M1011_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.1 SB=75005.7
+ A=0.063 P=1.14 MULT=1
MM1013 N_Y_M1011_d N_A_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.07665 PD=0.75 PS=0.785 NRD=0 NRS=21.42 M=1 R=2.8 SA=75002.6 SB=75005.2
+ A=0.063 P=1.14 MULT=1
MM1014 N_Y_M1014_d N_A_M1014_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.10185 AS=0.07665 PD=0.905 PS=0.785 NRD=22.848 NRS=2.856 M=1 R=2.8
+ SA=75003.1 SB=75004.7 A=0.063 P=1.14 MULT=1
MM1016 N_Y_M1014_d N_A_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.42
+ AD=0.10185 AS=0.0693 PD=0.905 PS=0.75 NRD=35.712 NRS=14.28 M=1 R=2.8
+ SA=75003.7 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1017 N_Y_M1017_d N_A_M1017_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75004.2 SB=75003.6
+ A=0.063 P=1.14 MULT=1
MM1028 N_Y_M1017_d N_A_M1028_g N_VGND_M1028_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0693 PD=0.75 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75004.7 SB=75003.1
+ A=0.063 P=1.14 MULT=1
MM1029 N_Y_M1029_d N_A_M1029_g N_VGND_M1028_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75005.2 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1031 N_Y_M1029_d N_A_M1031_g N_VGND_M1031_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0693 PD=0.75 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75005.7 SB=75002.2
+ A=0.063 P=1.14 MULT=1
MM1033 N_Y_M1033_d N_A_M1033_g N_VGND_M1031_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75006.1 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1035 N_Y_M1033_d N_A_M1035_g N_VGND_M1035_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0693 PD=0.75 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75006.6 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1036 N_Y_M1036_d N_A_M1036_g N_VGND_M1035_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75007.1 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1038 N_Y_M1036_d N_A_M1038_g N_VGND_M1038_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.1323 PD=0.75 PS=1.47 NRD=0 NRS=14.28 M=1 R=2.8 SA=75007.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1 AD=0.285
+ AS=0.15 PD=2.57 PS=1.3 NRD=0.9653 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90011.4 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90010.9 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1002_d N_A_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.2
+ SB=90010.5 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.6 SB=90010
+ A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1004_d N_A_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.1
+ SB=90009.5 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_Y_M1006_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.6 SB=90009
+ A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1007_d N_A_M1009_g N_Y_M1009_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90003.1
+ SB=90008.5 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_A_M1012_g N_Y_M1009_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90003.6
+ SB=90008.1 A=0.18 P=2.36 MULT=1
MM1015 N_VPWR_M1012_d N_A_M1015_g N_Y_M1015_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90004 SB=90007.6
+ A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1018_d N_A_M1018_g N_Y_M1015_s VPB PHIGHVT L=0.18 W=1 AD=0.1675
+ AS=0.15 PD=1.335 PS=1.3 NRD=5.8903 NRS=1.9503 M=1 R=5.55556 SA=90004.5
+ SB=90007.1 A=0.18 P=2.36 MULT=1
MM1019 N_VPWR_M1018_d N_A_M1019_g N_Y_M1019_s VPB PHIGHVT L=0.18 W=1 AD=0.1675
+ AS=0.2275 PD=1.335 PS=1.455 NRD=4.9053 NRS=27.5603 M=1 R=5.55556 SA=90005
+ SB=90006.6 A=0.18 P=2.36 MULT=1
MM1020 N_VPWR_M1020_d N_A_M1020_g N_Y_M1019_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.2275 PD=1.3 PS=1.455 NRD=0.9653 NRS=6.8753 M=1 R=5.55556 SA=90005.7
+ SB=90005.9 A=0.18 P=2.36 MULT=1
MM1021 N_VPWR_M1020_d N_A_M1021_g N_Y_M1021_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=2.9353 NRS=1.9503 M=1 R=5.55556 SA=90006.1
+ SB=90005.5 A=0.18 P=2.36 MULT=1
MM1022 N_VPWR_M1022_d N_A_M1022_g N_Y_M1021_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90006.6 SB=90005
+ A=0.18 P=2.36 MULT=1
MM1023 N_VPWR_M1022_d N_A_M1023_g N_Y_M1023_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90007.1
+ SB=90004.5 A=0.18 P=2.36 MULT=1
MM1024 N_VPWR_M1024_d N_A_M1024_g N_Y_M1023_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90007.6 SB=90004
+ A=0.18 P=2.36 MULT=1
MM1025 N_VPWR_M1024_d N_A_M1025_g N_Y_M1025_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90008.1
+ SB=90003.5 A=0.18 P=2.36 MULT=1
MM1026 N_VPWR_M1026_d N_A_M1026_g N_Y_M1025_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90008.5
+ SB=90003.1 A=0.18 P=2.36 MULT=1
MM1027 N_VPWR_M1026_d N_A_M1027_g N_Y_M1027_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90009 SB=90002.6
+ A=0.18 P=2.36 MULT=1
MM1030 N_VPWR_M1030_d N_A_M1030_g N_Y_M1027_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90009.5
+ SB=90002.1 A=0.18 P=2.36 MULT=1
MM1032 N_VPWR_M1030_d N_A_M1032_g N_Y_M1032_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90010 SB=90001.6
+ A=0.18 P=2.36 MULT=1
MM1034 N_VPWR_M1034_d N_A_M1034_g N_Y_M1032_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90010.5
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1037 N_VPWR_M1034_d N_A_M1037_g N_Y_M1037_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90010.9
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1039 N_VPWR_M1039_d N_A_M1039_g N_Y_M1037_s VPB PHIGHVT L=0.18 W=1 AD=0.275
+ AS=0.15 PD=2.55 PS=1.3 NRD=0.9653 NRS=1.9503 M=1 R=5.55556 SA=90011.4
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX40_noxref VNB VPB NWDIODE A=20.544 P=28.81
pX41_noxref noxref_7 Y Y PROBETYPE=1
c_152 VPB 0 8.51807e-20 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__clkinv_16.pxi.spice"
*
.ends
*
*
