* File: sky130_fd_sc_hdll__o211a_2.spice
* Created: Wed Sep  2 08:42:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o211a_2.pex.spice"
.subckt sky130_fd_sc_hdll__o211a_2  VNB VPB C1 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1001 A_120_47# N_C1_M1001_g N_A_27_47#_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.20475 PD=0.93 PS=1.93 NRD=15.684 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1004 N_A_206_47#_M1004_d N_B1_M1004_g A_120_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.091 PD=1.83 PS=0.93 NRD=0 NRS=15.684 M=1 R=4.33333 SA=75000.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_A_206_47#_M1005_d N_A2_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10075 AS=0.20475 PD=0.96 PS=1.93 NRD=5.532 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A1_M1009_g N_A_206_47#_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1105 AS=0.10075 PD=0.99 PS=0.96 NRD=3.684 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1006 N_X_M1006_d N_A_27_47#_M1006_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.117 AS=0.1105 PD=1.01 PS=0.99 NRD=5.532 NRS=7.38 M=1 R=4.33333 SA=75001.2
+ SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1007 N_X_M1006_d N_A_27_47#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.117 AS=0.3185 PD=1.01 PS=2.28 NRD=9.228 NRS=12.912 M=1 R=4.33333
+ SA=75001.7 SB=75000.4 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_C1_M1002_g N_A_27_47#_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90003.2 A=0.18 P=2.36 MULT=1
MM1008 N_A_27_47#_M1008_d N_B1_M1008_g N_VPWR_M1002_d VPB PHIGHVT L=0.18 W=1
+ AD=0.39 AS=0.15 PD=1.78 PS=1.3 NRD=15.7403 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90002.8 A=0.18 P=2.36 MULT=1
MM1010 A_406_297# N_A2_M1010_g N_A_27_47#_M1008_d VPB PHIGHVT L=0.18 W=1
+ AD=0.115 AS=0.39 PD=1.23 PS=1.78 NRD=11.8003 NRS=10.8153 M=1 R=5.55556
+ SA=90001.6 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_A1_M1011_g A_406_297# VPB PHIGHVT L=0.18 W=1 AD=0.205
+ AS=0.115 PD=1.41 PS=1.23 NRD=11.8003 NRS=11.8003 M=1 R=5.55556 SA=90002
+ SB=90001.4 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1011_d N_A_27_47#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.205 AS=0.15 PD=1.41 PS=1.3 NRD=13.7703 NRS=1.9503 M=1 R=5.55556
+ SA=90002.6 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_A_27_47#_M1003_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.41 AS=0.15 PD=2.82 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90003.1
+ SB=90000.3 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hdll__o211a_2.pxi.spice"
*
.ends
*
*
