* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__mux2_2 A0 A1 S VGND VNB VPB VPWR X
M1000 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=7.764e+11p pd=7.11e+06u as=2.9e+11p ps=2.58e+06u
M1001 a_280_21# S VPWR VPB phighvt w=640000u l=180000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1002 a_606_369# A0 a_79_21# VPB phighvt w=640000u l=180000u
+  ad=1.472e+11p pd=1.74e+06u as=1.92e+11p ps=1.88e+06u
M1003 VPWR S a_606_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_79_21# A0 a_310_47# VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=1.386e+11p ps=1.5e+06u
M1005 VGND S a_502_47# VNB nshort w=420000u l=150000u
+  ad=5.551e+11p pd=5.47e+06u as=3.108e+11p ps=2.32e+06u
M1006 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1007 a_502_47# A1 a_79_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_318_369# a_280_21# VPWR VPB phighvt w=640000u l=180000u
+  ad=4.992e+11p pd=2.84e+06u as=0p ps=0u
M1009 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_79_21# A1 a_318_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_310_47# a_280_21# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_280_21# S VGND VNB nshort w=420000u l=150000u
+  ad=1.155e+11p pd=1.39e+06u as=0p ps=0u
.ends
