* File: sky130_fd_sc_hdll__sdfxtp_4.pex.spice
* Created: Thu Aug 27 19:28:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_4%CLK 1 2 3 5 6 8 13
c38 1 0 2.71124e-20 $X=0.31 $Y=1.325
r39 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r40 6 9 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.5 $Y=1.665 $X2=0.31
+ $Y2=1.665
r41 6 8 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.5 $Y=1.74 $X2=0.5
+ $Y2=2.135
r42 3 16 89.156 $w=2.56e-07 $l=4.95076e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.33 $Y2=1.16
r43 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r44 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.31 $Y=1.59 $X2=0.31
+ $Y2=1.665
r45 1 16 39.2615 $w=2.56e-07 $l=1.74714e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.33 $Y2=1.16
r46 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.31 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_27_47# 1 2 9 12 13 15 18 20 21 23 24 26
+ 28 29 31 32 36 40 44 45 46 49 51 54 63 66 67 68 70 72 77 82 86
c238 66 0 1.55016e-19 $X=5.75 $Y=1.825
c239 46 0 1.76957e-19 $X=0.665 $Y=1.88
c240 36 0 7.21183e-20 $X=8.05 $Y=0.415
r241 85 87 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.275 $Y=1.41
+ $X2=7.275 $Y2=1.575
r242 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.25
+ $Y=1.41 $X2=7.25 $Y2=1.41
r243 82 85 16.2293 $w=3.2e-07 $l=9e-08 $layer=POLY_cond $X=7.275 $Y=1.32
+ $X2=7.275 $Y2=1.41
r244 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.55
+ $Y=1.74 $X2=5.55 $Y2=1.74
r245 76 77 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=0.94 $Y=1.235
+ $X2=0.97 $Y2=1.235
r246 71 86 19.9277 $w=2.38e-07 $l=4.15e-07 $layer=LI1_cond $X=7.285 $Y=1.825
+ $X2=7.285 $Y2=1.41
r247 70 72 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=7.31 $Y=1.825
+ $X2=7.115 $Y2=1.825
r248 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.31 $Y=1.825
+ $X2=7.31 $Y2=1.825
r249 68 72 1.5099 $w=1.4e-07 $l=1.22e-06 $layer=MET1_cond $X=5.895 $Y=1.87
+ $X2=7.115 $Y2=1.87
r250 66 81 6.49264 $w=3.53e-07 $l=2e-07 $layer=LI1_cond $X=5.75 $Y=1.832
+ $X2=5.55 $Y2=1.832
r251 65 68 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.75 $Y=1.825
+ $X2=5.895 $Y2=1.825
r252 65 67 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=5.75 $Y=1.825
+ $X2=5.555 $Y2=1.825
r253 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=1.825
+ $X2=5.75 $Y2=1.825
r254 63 67 5.76732 $w=1.4e-07 $l=4.66e-06 $layer=MET1_cond $X=0.895 $Y=1.87
+ $X2=5.555 $Y2=1.87
r255 60 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.75 $Y=1.825
+ $X2=0.895 $Y2=1.825
r256 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.75 $Y=1.825
+ $X2=0.75 $Y2=1.825
r257 52 76 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=0.81 $Y=1.235
+ $X2=0.94 $Y2=1.235
r258 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.81
+ $Y=1.235 $X2=0.81 $Y2=1.235
r259 49 61 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=1.795
+ $X2=0.78 $Y2=1.88
r260 49 51 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.78 $Y=1.795
+ $X2=0.78 $Y2=1.235
r261 48 51 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=0.805
+ $X2=0.78 $Y2=1.235
r262 47 54 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.35 $Y=1.88
+ $X2=0.265 $Y2=1.88
r263 46 61 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.665 $Y=1.88
+ $X2=0.78 $Y2=1.88
r264 46 47 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.665 $Y=1.88
+ $X2=0.35 $Y2=1.88
r265 44 48 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.665 $Y=0.72
+ $X2=0.78 $Y2=0.805
r266 44 45 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.665 $Y=0.72
+ $X2=0.345 $Y2=0.72
r267 38 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r268 38 40 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r269 34 36 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=8.05 $Y=1.245
+ $X2=8.05 $Y2=0.415
r270 33 82 20.4921 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=7.435 $Y=1.32
+ $X2=7.275 $Y2=1.32
r271 32 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.975 $Y=1.32
+ $X2=8.05 $Y2=1.245
r272 32 33 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=7.975 $Y=1.32
+ $X2=7.435 $Y2=1.32
r273 29 31 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.28 $Y=1.99
+ $X2=7.28 $Y2=2.275
r274 28 29 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.28 $Y=1.89 $X2=7.28
+ $Y2=1.99
r275 28 87 104.447 $w=2e-07 $l=3.15e-07 $layer=POLY_cond $X=7.28 $Y=1.89
+ $X2=7.28 $Y2=1.575
r276 24 80 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=5.515 $Y=1.99
+ $X2=5.575 $Y2=1.74
r277 24 26 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.515 $Y=1.99
+ $X2=5.515 $Y2=2.275
r278 23 80 31.9848 $w=2.95e-07 $l=1.92678e-07 $layer=POLY_cond $X=5.515 $Y=1.575
+ $X2=5.575 $Y2=1.74
r279 22 23 59.6839 $w=2e-07 $l=1.8e-07 $layer=POLY_cond $X=5.515 $Y=1.395
+ $X2=5.515 $Y2=1.575
r280 20 22 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=5.415 $Y=1.32
+ $X2=5.515 $Y2=1.395
r281 20 21 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=5.415 $Y=1.32
+ $X2=5.055 $Y2=1.32
r282 16 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.98 $Y=1.245
+ $X2=5.055 $Y2=1.32
r283 16 18 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=4.98 $Y=1.245
+ $X2=4.98 $Y2=0.415
r284 13 15 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.97 $Y=1.74
+ $X2=0.97 $Y2=2.135
r285 12 13 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.97 $Y=1.64 $X2=0.97
+ $Y2=1.74
r286 11 77 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=0.97 $Y=1.37
+ $X2=0.97 $Y2=1.235
r287 11 12 89.5258 $w=2e-07 $l=2.7e-07 $layer=POLY_cond $X=0.97 $Y=1.37 $X2=0.97
+ $Y2=1.64
r288 7 76 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.94 $Y=1.1
+ $X2=0.94 $Y2=1.235
r289 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.94 $Y=1.1 $X2=0.94
+ $Y2=0.445
r290 2 54 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.14
+ $Y=1.815 $X2=0.265 $Y2=1.96
r291 1 40 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_4%SCE 1 3 6 8 10 13 15 19 22 28 33 35 37
c100 35 0 4.47538e-20 $X=2.047 $Y=0.785
c101 28 0 7.84804e-20 $X=1.965 $Y=1.52
c102 15 0 1.59107e-19 $X=3.335 $Y=0.7
c103 6 0 1.4868e-19 $X=1.95 $Y=0.445
r104 35 37 1.89207 $w=3.33e-07 $l=5.5e-08 $layer=LI1_cond $X=2.047 $Y=0.785
+ $X2=2.047 $Y2=0.84
r105 28 30 81.5018 $w=2.75e-07 $l=4.65e-07 $layer=POLY_cond $X=1.965 $Y=1.577
+ $X2=2.43 $Y2=1.577
r106 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.965
+ $Y=1.52 $X2=1.965 $Y2=1.52
r107 26 28 0.876364 $w=2.75e-07 $l=5e-09 $layer=POLY_cond $X=1.96 $Y=1.577
+ $X2=1.965 $Y2=1.577
r108 25 26 1.75273 $w=2.75e-07 $l=1e-08 $layer=POLY_cond $X=1.95 $Y=1.577
+ $X2=1.96 $Y2=1.577
r109 22 35 2.62343 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.047 $Y=0.7
+ $X2=2.047 $Y2=0.785
r110 22 29 22.8081 $w=3.33e-07 $l=6.63e-07 $layer=LI1_cond $X=2.047 $Y=0.857
+ $X2=2.047 $Y2=1.52
r111 22 37 0.584822 $w=3.33e-07 $l=1.7e-08 $layer=LI1_cond $X=2.047 $Y=0.857
+ $X2=2.047 $Y2=0.84
r112 20 33 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=3.42 $Y=0.95
+ $X2=3.53 $Y2=0.95
r113 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.42
+ $Y=0.95 $X2=3.42 $Y2=0.95
r114 17 19 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.42 $Y=0.785
+ $X2=3.42 $Y2=0.95
r115 16 22 5.18513 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.215 $Y=0.7
+ $X2=2.047 $Y2=0.7
r116 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.335 $Y=0.7
+ $X2=3.42 $Y2=0.785
r117 15 16 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=3.335 $Y=0.7
+ $X2=2.215 $Y2=0.7
r118 11 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=0.785
+ $X2=3.53 $Y2=0.95
r119 11 13 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.53 $Y=0.785
+ $X2=3.53 $Y2=0.445
r120 8 30 12.7119 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.43 $Y=1.77
+ $X2=2.43 $Y2=1.577
r121 8 10 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.43 $Y=1.77
+ $X2=2.43 $Y2=2.165
r122 4 25 16.9318 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.95 $Y=1.385
+ $X2=1.95 $Y2=1.577
r123 4 6 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.95 $Y=1.385 $X2=1.95
+ $Y2=0.445
r124 1 26 12.7119 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.96 $Y=1.77
+ $X2=1.96 $Y2=1.577
r125 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.96 $Y=1.77
+ $X2=1.96 $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_319_47# 1 2 9 11 13 15 18 20 23 24 28
+ 34 36 39 40 42
c118 39 0 2.2716e-19 $X=2.55 $Y=1.04
c119 28 0 1.61748e-19 $X=3.44 $Y=1.52
r120 40 44 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.525 $Y=1.04
+ $X2=2.525 $Y2=0.875
r121 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.55
+ $Y=1.04 $X2=2.55 $Y2=1.04
r122 31 34 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.62 $Y=0.36
+ $X2=1.74 $Y2=0.36
r123 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.44
+ $Y=1.52 $X2=3.44 $Y2=1.52
r124 26 28 19.338 $w=1.93e-07 $l=3.4e-07 $layer=LI1_cond $X=3.427 $Y=1.86
+ $X2=3.427 $Y2=1.52
r125 25 42 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.555 $Y=1.967
+ $X2=2.47 $Y2=1.967
r126 24 26 6.83761 $w=2.15e-07 $l=1.47743e-07 $layer=LI1_cond $X=3.33 $Y=1.967
+ $X2=3.427 $Y2=1.86
r127 24 25 41.5415 $w=2.13e-07 $l=7.75e-07 $layer=LI1_cond $X=3.33 $Y=1.967
+ $X2=2.555 $Y2=1.967
r128 23 42 2.20034 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.47 $Y=1.86
+ $X2=2.47 $Y2=1.967
r129 22 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.47 $Y=1.125
+ $X2=2.47 $Y2=1.04
r130 22 23 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.47 $Y=1.125
+ $X2=2.47 $Y2=1.86
r131 21 36 1.46632 $w=2.15e-07 $l=1.38e-07 $layer=LI1_cond $X=1.81 $Y=1.967
+ $X2=1.672 $Y2=1.967
r132 20 42 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=1.967
+ $X2=2.47 $Y2=1.967
r133 20 21 30.8211 $w=2.13e-07 $l=5.75e-07 $layer=LI1_cond $X=2.385 $Y=1.967
+ $X2=1.81 $Y2=1.967
r134 16 36 5.02022 $w=2.22e-07 $l=1.08e-07 $layer=LI1_cond $X=1.672 $Y=2.075
+ $X2=1.672 $Y2=1.967
r135 16 18 4.1907 $w=2.73e-07 $l=1e-07 $layer=LI1_cond $X=1.672 $Y=2.075
+ $X2=1.672 $Y2=2.175
r136 15 36 5.02022 $w=2.22e-07 $l=1.30434e-07 $layer=LI1_cond $X=1.62 $Y=1.86
+ $X2=1.672 $Y2=1.967
r137 14 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.445
+ $X2=1.62 $Y2=0.36
r138 14 15 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=1.62 $Y=0.445
+ $X2=1.62 $Y2=1.86
r139 11 29 48.1208 $w=2.95e-07 $l=2.7157e-07 $layer=POLY_cond $X=3.42 $Y=1.77
+ $X2=3.465 $Y2=1.52
r140 11 13 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.42 $Y=1.77
+ $X2=3.42 $Y2=2.165
r141 9 44 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.51 $Y=0.445
+ $X2=2.51 $Y2=0.875
r142 2 18 600 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=1 $X=1.6
+ $Y=1.845 $X2=1.725 $Y2=2.175
r143 1 34 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.74 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_4%D 1 3 6 8 15
r39 11 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.91
+ $Y=1.52 $X2=2.91 $Y2=1.52
r40 8 15 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.99 $Y=1.52 $X2=2.91
+ $Y2=1.52
r41 4 11 38.535 $w=3.06e-07 $l=2.0106e-07 $layer=POLY_cond $X=3 $Y=1.355
+ $X2=2.92 $Y2=1.52
r42 4 6 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=3 $Y=1.355 $X2=3
+ $Y2=0.445
r43 1 11 47.4839 $w=3.06e-07 $l=2.64575e-07 $layer=POLY_cond $X=2.95 $Y=1.77
+ $X2=2.92 $Y2=1.52
r44 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.95 $Y=1.77 $X2=2.95
+ $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_4%SCD 3 6 7 9 10 13
c53 6 0 1.61748e-19 $X=3.935 $Y=1.67
c54 3 0 1.59107e-19 $X=3.91 $Y=0.445
r55 13 16 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.355
+ $X2=3.995 $Y2=1.52
r56 13 15 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.355
+ $X2=3.995 $Y2=1.19
r57 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.97
+ $Y=1.355 $X2=3.97 $Y2=1.355
r58 10 14 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.91 $Y=1.19
+ $X2=3.91 $Y2=1.355
r59 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.935 $Y=1.77
+ $X2=3.935 $Y2=2.165
r60 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.935 $Y=1.67 $X2=3.935
+ $Y2=1.77
r61 6 16 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=3.935 $Y=1.67 $X2=3.935
+ $Y2=1.52
r62 3 15 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.91 $Y=0.445
+ $X2=3.91 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_203_47# 1 2 7 9 10 12 13 15 16 18 21 25
+ 26 30 41 45 46 48 50 55 57 62 67
c205 48 0 7.21183e-20 $X=7.31 $Y=0.805
c206 46 0 1.7664e-19 $X=5.385 $Y=0.805
r207 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.53
+ $Y=0.87 $X2=7.53 $Y2=0.87
r208 59 62 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=7.385 $Y=0.87
+ $X2=7.53 $Y2=0.87
r209 54 57 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=5.45 $Y=0.87
+ $X2=5.56 $Y2=0.87
r210 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.45
+ $Y=0.87 $X2=5.45 $Y2=0.87
r211 49 63 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=7.31 $Y=0.87
+ $X2=7.53 $Y2=0.87
r212 48 50 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=7.31 $Y=0.805
+ $X2=7.115 $Y2=0.805
r213 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.31 $Y=0.805
+ $X2=7.31 $Y2=0.805
r214 46 50 2.14109 $w=1.4e-07 $l=1.73e-06 $layer=MET1_cond $X=5.385 $Y=0.85
+ $X2=7.115 $Y2=0.85
r215 44 55 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=5.24 $Y=0.87
+ $X2=5.45 $Y2=0.87
r216 44 76 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=5.24 $Y=0.87
+ $X2=5.05 $Y2=0.87
r217 43 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.24 $Y=0.805
+ $X2=5.385 $Y2=0.805
r218 43 45 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=5.24 $Y=0.805
+ $X2=5.045 $Y2=0.805
r219 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.24 $Y=0.805
+ $X2=5.24 $Y2=0.805
r220 41 45 4.52969 $w=1.4e-07 $l=3.66e-06 $layer=MET1_cond $X=1.385 $Y=0.85
+ $X2=5.045 $Y2=0.85
r221 39 71 57.8727 $w=2.28e-07 $l=1.155e-06 $layer=LI1_cond $X=1.23 $Y=0.805
+ $X2=1.23 $Y2=1.96
r222 39 67 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.23 $Y=0.805
+ $X2=1.23 $Y2=0.51
r223 38 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.24 $Y=0.805
+ $X2=1.385 $Y2=0.805
r224 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.24 $Y=0.805
+ $X2=1.24 $Y2=0.805
r225 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.81
+ $Y=1.74 $X2=7.81 $Y2=1.74
r226 27 30 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=7.67 $Y=1.74
+ $X2=7.81 $Y2=1.74
r227 26 63 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=7.575 $Y=0.87
+ $X2=7.53 $Y2=0.87
r228 25 27 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=7.67 $Y=1.575
+ $X2=7.67 $Y2=1.74
r229 24 26 7.47963 $w=3.3e-07 $l=2.07123e-07 $layer=LI1_cond $X=7.67 $Y=1.035
+ $X2=7.575 $Y2=0.87
r230 24 25 31.5215 $w=1.88e-07 $l=5.4e-07 $layer=LI1_cond $X=7.67 $Y=1.035
+ $X2=7.67 $Y2=1.575
r231 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.99
+ $Y=1.74 $X2=4.99 $Y2=1.74
r232 19 76 1.49285 $w=2.9e-07 $l=1.65e-07 $layer=LI1_cond $X=5.05 $Y=1.035
+ $X2=5.05 $Y2=0.87
r233 19 21 28.0163 $w=2.88e-07 $l=7.05e-07 $layer=LI1_cond $X=5.05 $Y=1.035
+ $X2=5.05 $Y2=1.74
r234 16 31 46.5577 $w=3.26e-07 $l=2.89396e-07 $layer=POLY_cond $X=7.75 $Y=1.99
+ $X2=7.835 $Y2=1.74
r235 16 18 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.75 $Y=1.99
+ $X2=7.75 $Y2=2.275
r236 13 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.385 $Y=0.705
+ $X2=7.385 $Y2=0.87
r237 13 15 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.385 $Y=0.705
+ $X2=7.385 $Y2=0.415
r238 10 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.56 $Y=0.705
+ $X2=5.56 $Y2=0.87
r239 10 12 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.56 $Y=0.705
+ $X2=5.56 $Y2=0.415
r240 7 22 46.5577 $w=3.26e-07 $l=2.57391e-07 $layer=POLY_cond $X=5 $Y=1.99
+ $X2=5.015 $Y2=1.74
r241 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5 $Y=1.99 $X2=5
+ $Y2=2.275
r242 2 71 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.06
+ $Y=1.815 $X2=1.205 $Y2=1.96
r243 1 67 182 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_1189_183# 1 2 8 9 11 14 16 22 25 27 29
+ 31 32 35
c98 9 0 1.55016e-19 $X=6.045 $Y=1.99
r99 34 35 10.6895 $w=2.48e-07 $l=5.5e-08 $layer=POLY_cond $X=6.045 $Y=0.93
+ $X2=6.1 $Y2=0.93
r100 31 32 7.18001 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=6.925 $Y=2.3
+ $X2=6.925 $Y2=2.135
r101 25 27 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.995 $Y=0.45
+ $X2=7.12 $Y2=0.45
r102 23 29 6.6318 $w=2.2e-07 $l=1.5e-07 $layer=LI1_cond $X=6.885 $Y=1.065
+ $X2=6.885 $Y2=0.915
r103 23 32 56.0506 $w=2.18e-07 $l=1.07e-06 $layer=LI1_cond $X=6.885 $Y=1.065
+ $X2=6.885 $Y2=2.135
r104 22 29 6.6318 $w=2.2e-07 $l=1.5e-07 $layer=LI1_cond $X=6.885 $Y=0.765
+ $X2=6.885 $Y2=0.915
r105 21 25 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=6.885 $Y=0.535
+ $X2=6.995 $Y2=0.45
r106 21 22 12.0483 $w=2.18e-07 $l=2.3e-07 $layer=LI1_cond $X=6.885 $Y=0.535
+ $X2=6.885 $Y2=0.765
r107 19 35 25.2661 $w=2.48e-07 $l=1.3e-07 $layer=POLY_cond $X=6.23 $Y=0.93
+ $X2=6.1 $Y2=0.93
r108 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.23
+ $Y=0.93 $X2=6.23 $Y2=0.93
r109 16 29 0.253446 $w=3e-07 $l=1.1e-07 $layer=LI1_cond $X=6.775 $Y=0.915
+ $X2=6.885 $Y2=0.915
r110 16 18 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=6.775 $Y=0.915
+ $X2=6.23 $Y2=0.915
r111 12 35 14.534 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.1 $Y=0.795
+ $X2=6.1 $Y2=0.93
r112 12 14 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.1 $Y=0.795
+ $X2=6.1 $Y2=0.445
r113 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.045 $Y=1.99
+ $X2=6.045 $Y2=2.275
r114 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=6.045 $Y=1.89 $X2=6.045
+ $Y2=1.99
r115 7 34 7.89931 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=6.045 $Y=1.065
+ $X2=6.045 $Y2=0.93
r116 7 8 273.551 $w=2e-07 $l=8.25e-07 $layer=POLY_cond $X=6.045 $Y=1.065
+ $X2=6.045 $Y2=1.89
r117 2 31 600 $w=1.7e-07 $l=6.33364e-07 $layer=licon1_PDIFF $count=1 $X=6.845
+ $Y=1.735 $X2=6.99 $Y2=2.3
r118 1 27 182 $w=1.7e-07 $l=2.85832e-07 $layer=licon1_NDIFF $count=1 $X=6.955
+ $Y=0.235 $X2=7.12 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_1011_47# 1 2 8 9 11 14 15 16 17 18 19
+ 23 28 30 31 33
r117 36 37 15.25 $w=2.76e-07 $l=3.45e-07 $layer=LI1_cond $X=5.81 $Y=1.41
+ $X2=6.155 $Y2=1.41
r118 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.52
+ $Y=1.41 $X2=6.52 $Y2=1.41
r119 31 37 4.4292 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=6.265 $Y=1.41
+ $X2=6.155 $Y2=1.41
r120 31 33 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=6.265 $Y=1.41
+ $X2=6.52 $Y2=1.41
r121 29 37 2.0678 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=6.155 $Y=1.575
+ $X2=6.155 $Y2=1.41
r122 29 30 32.216 $w=2.18e-07 $l=6.15e-07 $layer=LI1_cond $X=6.155 $Y=1.575
+ $X2=6.155 $Y2=2.19
r123 28 36 3.57235 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.81 $Y=1.245
+ $X2=5.81 $Y2=1.41
r124 27 28 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.81 $Y=0.535
+ $X2=5.81 $Y2=1.245
r125 23 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.725 $Y=0.45
+ $X2=5.81 $Y2=0.535
r126 23 25 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=5.725 $Y=0.45
+ $X2=5.3 $Y2=0.45
r127 19 30 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=6.045 $Y=2.275
+ $X2=6.155 $Y2=2.19
r128 19 21 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=6.045 $Y=2.275
+ $X2=5.26 $Y2=2.275
r129 17 34 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.52 $Y2=1.41
r130 17 18 0.448535 $w=2.7e-07 $l=1.253e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.755 $Y2=1.467
r131 15 16 54.0301 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=6.805 $Y=0.95
+ $X2=6.805 $Y2=1.1
r132 14 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.88 $Y=0.555
+ $X2=6.88 $Y2=0.95
r133 9 18 27.0491 $w=1.9e-07 $l=1.93e-07 $layer=POLY_cond $X=6.755 $Y=1.66
+ $X2=6.755 $Y2=1.467
r134 9 11 120.5 $w=1.8e-07 $l=4.5e-07 $layer=POLY_cond $X=6.755 $Y=1.66
+ $X2=6.755 $Y2=2.11
r135 8 18 27.0491 $w=1.9e-07 $l=1.92e-07 $layer=POLY_cond $X=6.755 $Y=1.275
+ $X2=6.755 $Y2=1.467
r136 8 16 58.026 $w=2e-07 $l=1.75e-07 $layer=POLY_cond $X=6.755 $Y=1.275
+ $X2=6.755 $Y2=1.1
r137 2 21 600 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_PDIFF $count=1 $X=5.09
+ $Y=2.065 $X2=5.26 $Y2=2.275
r138 1 25 182 $w=1.7e-07 $l=3.35708e-07 $layer=licon1_NDIFF $count=1 $X=5.055
+ $Y=0.235 $X2=5.3 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_1667_315# 1 2 7 9 12 14 16 17 19 20 22
+ 23 25 26 28 29 31 32 34 35 37 38 45 48 50 56 60 63 64 74
r139 74 75 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=11.43 $Y=1.202
+ $X2=11.455 $Y2=1.202
r140 71 72 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=10.935 $Y=1.202
+ $X2=10.96 $Y2=1.202
r141 70 71 59.1132 $w=3.71e-07 $l=4.55e-07 $layer=POLY_cond $X=10.48 $Y=1.202
+ $X2=10.935 $Y2=1.202
r142 69 70 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=10.455 $Y=1.202
+ $X2=10.48 $Y2=1.202
r143 66 67 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=9.985 $Y=1.202
+ $X2=10.01 $Y2=1.202
r144 60 62 16.9646 $w=3.58e-07 $l=4.4e-07 $layer=LI1_cond $X=9.32 $Y=0.385
+ $X2=9.32 $Y2=0.825
r145 57 74 27.9326 $w=3.71e-07 $l=2.15e-07 $layer=POLY_cond $X=11.215 $Y=1.202
+ $X2=11.43 $Y2=1.202
r146 57 72 33.1294 $w=3.71e-07 $l=2.55e-07 $layer=POLY_cond $X=11.215 $Y=1.202
+ $X2=10.96 $Y2=1.202
r147 56 57 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.215
+ $Y=1.16 $X2=11.215 $Y2=1.16
r148 54 69 53.2668 $w=3.71e-07 $l=4.1e-07 $layer=POLY_cond $X=10.045 $Y=1.202
+ $X2=10.455 $Y2=1.202
r149 54 67 4.54717 $w=3.71e-07 $l=3.5e-08 $layer=POLY_cond $X=10.045 $Y=1.202
+ $X2=10.01 $Y2=1.202
r150 53 56 53.9343 $w=2.48e-07 $l=1.17e-06 $layer=LI1_cond $X=10.045 $Y=1.2
+ $X2=11.215 $Y2=1.2
r151 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.045
+ $Y=1.16 $X2=10.045 $Y2=1.16
r152 51 64 0.237926 $w=2.5e-07 $l=9.3e-08 $layer=LI1_cond $X=9.505 $Y=1.2
+ $X2=9.412 $Y2=1.2
r153 51 53 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=9.505 $Y=1.2
+ $X2=10.045 $Y2=1.2
r154 50 63 6.7841 $w=2.35e-07 $l=1.88348e-07 $layer=LI1_cond $X=9.412 $Y=1.575
+ $X2=9.362 $Y2=1.74
r155 49 64 6.65529 $w=1.82e-07 $l=1.25e-07 $layer=LI1_cond $X=9.412 $Y=1.325
+ $X2=9.412 $Y2=1.2
r156 49 50 14.9877 $w=1.83e-07 $l=2.5e-07 $layer=LI1_cond $X=9.412 $Y=1.325
+ $X2=9.412 $Y2=1.575
r157 48 64 6.65529 $w=1.82e-07 $l=1.25996e-07 $layer=LI1_cond $X=9.41 $Y=1.075
+ $X2=9.412 $Y2=1.2
r158 48 62 15.404 $w=1.78e-07 $l=2.5e-07 $layer=LI1_cond $X=9.41 $Y=1.075
+ $X2=9.41 $Y2=0.825
r159 43 63 6.7841 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=9.362 $Y=1.905
+ $X2=9.362 $Y2=1.74
r160 43 45 1.81965 $w=2.83e-07 $l=4.5e-08 $layer=LI1_cond $X=9.362 $Y=1.905
+ $X2=9.362 $Y2=1.95
r161 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.64
+ $Y=1.74 $X2=8.64 $Y2=1.74
r162 38 63 0.153733 $w=3.3e-07 $l=1.42e-07 $layer=LI1_cond $X=9.22 $Y=1.74
+ $X2=9.362 $Y2=1.74
r163 38 40 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=9.22 $Y=1.74
+ $X2=8.64 $Y2=1.74
r164 35 75 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.455 $Y=0.995
+ $X2=11.455 $Y2=1.202
r165 35 37 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.455 $Y=0.995
+ $X2=11.455 $Y2=0.56
r166 32 74 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=11.43 $Y=1.41
+ $X2=11.43 $Y2=1.202
r167 32 34 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.43 $Y=1.41
+ $X2=11.43 $Y2=1.985
r168 29 72 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.96 $Y=1.41
+ $X2=10.96 $Y2=1.202
r169 29 31 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.96 $Y=1.41
+ $X2=10.96 $Y2=1.985
r170 26 71 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.935 $Y=0.995
+ $X2=10.935 $Y2=1.202
r171 26 28 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.935 $Y=0.995
+ $X2=10.935 $Y2=0.56
r172 23 70 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.48 $Y=1.41
+ $X2=10.48 $Y2=1.202
r173 23 25 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.48 $Y=1.41
+ $X2=10.48 $Y2=1.985
r174 20 69 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.455 $Y=0.995
+ $X2=10.455 $Y2=1.202
r175 20 22 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.455 $Y=0.995
+ $X2=10.455 $Y2=0.56
r176 17 67 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.01 $Y=1.41
+ $X2=10.01 $Y2=1.202
r177 17 19 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.01 $Y=1.41
+ $X2=10.01 $Y2=1.985
r178 14 66 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.985 $Y=0.995
+ $X2=9.985 $Y2=1.202
r179 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.985 $Y=0.995
+ $X2=9.985 $Y2=0.56
r180 10 41 39.3952 $w=3.9e-07 $l=1.79374e-07 $layer=POLY_cond $X=8.525 $Y=1.575
+ $X2=8.555 $Y2=1.74
r181 10 12 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=8.525 $Y=1.575
+ $X2=8.525 $Y2=0.445
r182 7 41 44.9977 $w=3.9e-07 $l=3.04138e-07 $layer=POLY_cond $X=8.435 $Y=1.99
+ $X2=8.555 $Y2=1.74
r183 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=8.435 $Y=1.99
+ $X2=8.435 $Y2=2.275
r184 2 45 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=9.18
+ $Y=1.485 $X2=9.305 $Y2=1.95
r185 1 60 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=9.18
+ $Y=0.235 $X2=9.305 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_1474_413# 1 2 7 9 10 12 13 14 15 19 26
+ 29 32 33
c89 10 0 1.67668e-19 $X=9.565 $Y=0.995
r90 32 34 11.1226 $w=3.48e-07 $l=2.45e-07 $layer=LI1_cond $X=8.16 $Y=1.16
+ $X2=8.16 $Y2=1.405
r91 32 33 7.01492 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.16 $Y=1.16
+ $X2=8.16 $Y2=0.995
r92 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.065
+ $Y=1.16 $X2=9.065 $Y2=1.16
r93 27 32 1.07274 $w=3.3e-07 $l=1.75e-07 $layer=LI1_cond $X=8.335 $Y=1.16
+ $X2=8.16 $Y2=1.16
r94 27 29 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=8.335 $Y=1.16
+ $X2=9.065 $Y2=1.16
r95 26 34 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=8.25 $Y=2.165
+ $X2=8.25 $Y2=1.405
r96 23 33 24.0965 $w=2.18e-07 $l=4.6e-07 $layer=LI1_cond $X=8.095 $Y=0.535
+ $X2=8.095 $Y2=0.995
r97 19 23 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=7.985 $Y=0.45
+ $X2=8.095 $Y2=0.535
r98 19 21 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.985 $Y=0.45
+ $X2=7.73 $Y2=0.45
r99 15 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.165 $Y=2.25
+ $X2=8.25 $Y2=2.165
r100 15 17 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=8.165 $Y=2.25
+ $X2=7.515 $Y2=2.25
r101 13 30 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=9.44 $Y=1.16
+ $X2=9.065 $Y2=1.16
r102 13 14 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=9.44 $Y=1.16
+ $X2=9.54 $Y2=1.202
r103 10 14 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=9.565 $Y=0.995
+ $X2=9.54 $Y2=1.202
r104 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.565 $Y=0.995
+ $X2=9.565 $Y2=0.56
r105 7 14 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=9.54 $Y=1.41
+ $X2=9.54 $Y2=1.202
r106 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.54 $Y=1.41
+ $X2=9.54 $Y2=1.985
r107 2 17 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=7.37
+ $Y=2.065 $X2=7.515 $Y2=2.25
r108 1 21 182 $w=1.7e-07 $l=3.6187e-07 $layer=licon1_NDIFF $count=1 $X=7.46
+ $Y=0.235 $X2=7.73 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_4%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51
+ 53 55 58 59 61 62 64 65 67 68 70 71 72 74 79 109 114 117 121
c175 8 0 1.26199e-19 $X=11.52 $Y=1.485
c176 1 0 1.76957e-19 $X=0.59 $Y=1.815
r177 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r178 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r179 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r180 112 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=11.73 $Y2=2.72
r181 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r182 109 120 3.40825 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.58 $Y=2.72
+ $X2=11.77 $Y2=2.72
r183 109 111 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=11.58 $Y=2.72
+ $X2=11.27 $Y2=2.72
r184 108 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=11.27 $Y2=2.72
r185 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r186 105 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=10.35 $Y2=2.72
r187 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r188 102 105 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r189 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r190 99 102 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=8.51 $Y2=2.72
r191 98 101 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=6.67 $Y=2.72
+ $X2=8.51 $Y2=2.72
r192 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r193 96 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r194 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r195 93 96 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=6.21 $Y2=2.72
r196 92 95 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=6.21 $Y2=2.72
r197 92 93 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r198 90 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r199 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r200 87 90 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r201 87 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r202 86 89 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r203 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r204 84 117 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.36 $Y=2.72
+ $X2=2.17 $Y2=2.72
r205 84 86 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.36 $Y=2.72
+ $X2=2.53 $Y2=2.72
r206 83 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r207 83 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r208 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r209 80 114 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.9 $Y=2.72
+ $X2=0.71 $Y2=2.72
r210 80 82 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.9 $Y=2.72
+ $X2=1.61 $Y2=2.72
r211 79 117 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.98 $Y=2.72
+ $X2=2.17 $Y2=2.72
r212 79 82 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.98 $Y=2.72
+ $X2=1.61 $Y2=2.72
r213 74 114 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.71 $Y2=2.72
r214 74 76 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.23 $Y2=2.72
r215 72 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r216 72 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r217 70 107 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=10.64 $Y=2.72
+ $X2=10.35 $Y2=2.72
r218 70 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.64 $Y=2.72
+ $X2=10.725 $Y2=2.72
r219 69 111 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=10.81 $Y=2.72
+ $X2=11.27 $Y2=2.72
r220 69 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.81 $Y=2.72
+ $X2=10.725 $Y2=2.72
r221 67 104 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=9.69 $Y=2.72
+ $X2=9.43 $Y2=2.72
r222 67 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.69 $Y=2.72
+ $X2=9.775 $Y2=2.72
r223 66 107 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=9.86 $Y=2.72
+ $X2=10.35 $Y2=2.72
r224 66 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.86 $Y=2.72
+ $X2=9.775 $Y2=2.72
r225 64 101 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=8.565 $Y=2.72
+ $X2=8.51 $Y2=2.72
r226 64 65 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=8.565 $Y=2.72
+ $X2=8.717 $Y2=2.72
r227 63 104 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.87 $Y=2.72
+ $X2=9.43 $Y2=2.72
r228 63 65 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.87 $Y=2.72
+ $X2=8.717 $Y2=2.72
r229 61 95 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.435 $Y=2.72
+ $X2=6.21 $Y2=2.72
r230 61 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=2.72
+ $X2=6.52 $Y2=2.72
r231 60 98 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.605 $Y=2.72
+ $X2=6.67 $Y2=2.72
r232 60 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.605 $Y=2.72
+ $X2=6.52 $Y2=2.72
r233 58 89 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.11 $Y=2.72 $X2=3.91
+ $Y2=2.72
r234 58 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=2.72
+ $X2=4.195 $Y2=2.72
r235 57 92 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.28 $Y=2.72 $X2=4.37
+ $Y2=2.72
r236 57 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.28 $Y=2.72
+ $X2=4.195 $Y2=2.72
r237 53 120 3.40825 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=11.665 $Y=2.635
+ $X2=11.77 $Y2=2.72
r238 53 55 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=11.665 $Y=2.635
+ $X2=11.665 $Y2=2.01
r239 49 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.725 $Y=2.635
+ $X2=10.725 $Y2=2.72
r240 49 51 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=10.725 $Y=2.635
+ $X2=10.725 $Y2=2.01
r241 45 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.775 $Y=2.635
+ $X2=9.775 $Y2=2.72
r242 45 47 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=9.775 $Y=2.635
+ $X2=9.775 $Y2=1.79
r243 41 65 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.717 $Y=2.635
+ $X2=8.717 $Y2=2.72
r244 41 43 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=8.717 $Y=2.635
+ $X2=8.717 $Y2=2.3
r245 37 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=2.635
+ $X2=6.52 $Y2=2.72
r246 37 39 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.52 $Y=2.635
+ $X2=6.52 $Y2=2
r247 33 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.195 $Y=2.635
+ $X2=4.195 $Y2=2.72
r248 33 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.195 $Y=2.635
+ $X2=4.195 $Y2=2.33
r249 29 117 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=2.635
+ $X2=2.17 $Y2=2.72
r250 29 31 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=2.17 $Y=2.635
+ $X2=2.17 $Y2=2.33
r251 25 114 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=2.635
+ $X2=0.71 $Y2=2.72
r252 25 27 12.5859 $w=3.78e-07 $l=4.15e-07 $layer=LI1_cond $X=0.71 $Y=2.635
+ $X2=0.71 $Y2=2.22
r253 8 55 300 $w=1.7e-07 $l=5.93085e-07 $layer=licon1_PDIFF $count=2 $X=11.52
+ $Y=1.485 $X2=11.665 $Y2=2.01
r254 7 51 300 $w=1.7e-07 $l=5.97495e-07 $layer=licon1_PDIFF $count=2 $X=10.57
+ $Y=1.485 $X2=10.725 $Y2=2.01
r255 6 47 300 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=2 $X=9.63
+ $Y=1.485 $X2=9.775 $Y2=1.79
r256 5 43 600 $w=1.7e-07 $l=3.53483e-07 $layer=licon1_PDIFF $count=1 $X=8.525
+ $Y=2.065 $X2=8.78 $Y2=2.3
r257 4 39 300 $w=1.7e-07 $l=4.16233e-07 $layer=licon1_PDIFF $count=2 $X=6.135
+ $Y=2.065 $X2=6.52 $Y2=2
r258 3 35 600 $w=1.7e-07 $l=5.63627e-07 $layer=licon1_PDIFF $count=1 $X=4.025
+ $Y=1.845 $X2=4.195 $Y2=2.33
r259 2 31 600 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=1.845 $X2=2.195 $Y2=2.33
r260 1 27 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.815 $X2=0.735 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_608_369# 1 2 3 4 13 17 22 24 25 26 27
+ 28 30 32 36 38 39
c113 30 0 1.7664e-19 $X=4.65 $Y=0.695
r114 39 41 21.3062 $w=2.09e-07 $l=3.65e-07 $layer=LI1_cond $X=4.682 $Y=1.91
+ $X2=4.682 $Y2=2.275
r115 33 36 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.65 $Y=0.45 $X2=4.75
+ $Y2=0.45
r116 32 39 5.42244 $w=2.09e-07 $l=9.97246e-08 $layer=LI1_cond $X=4.65 $Y=1.825
+ $X2=4.682 $Y2=1.91
r117 31 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.65 $Y=0.865
+ $X2=4.65 $Y2=0.78
r118 31 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.65 $Y=0.865
+ $X2=4.65 $Y2=1.825
r119 30 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.65 $Y=0.695
+ $X2=4.65 $Y2=0.78
r120 29 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.65 $Y=0.535
+ $X2=4.65 $Y2=0.45
r121 29 30 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.65 $Y=0.535
+ $X2=4.65 $Y2=0.695
r122 27 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=0.78
+ $X2=4.65 $Y2=0.78
r123 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.565 $Y=0.78
+ $X2=3.895 $Y2=0.78
r124 25 39 1.94907 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=4.565 $Y=1.91
+ $X2=4.682 $Y2=1.91
r125 25 26 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=4.565 $Y=1.91
+ $X2=3.89 $Y2=1.91
r126 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.81 $Y=0.695
+ $X2=3.895 $Y2=0.78
r127 23 24 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.81 $Y=0.445
+ $X2=3.81 $Y2=0.695
r128 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.805 $Y=1.995
+ $X2=3.89 $Y2=1.91
r129 21 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.805 $Y=1.995
+ $X2=3.805 $Y2=2.245
r130 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.725 $Y=0.36
+ $X2=3.81 $Y2=0.445
r131 17 19 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.725 $Y=0.36
+ $X2=3.265 $Y2=0.36
r132 13 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.72 $Y=2.33
+ $X2=3.805 $Y2=2.245
r133 13 15 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.72 $Y=2.33
+ $X2=3.185 $Y2=2.33
r134 4 41 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=4.59
+ $Y=2.065 $X2=4.715 $Y2=2.275
r135 3 15 600 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=1.845 $X2=3.185 $Y2=2.33
r136 2 36 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=4.625
+ $Y=0.235 $X2=4.75 $Y2=0.45
r137 1 19 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=3.075
+ $Y=0.235 $X2=3.265 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_4%Q 1 2 3 4 15 17 19 21 22 23 27 31 33 35
+ 39 41 44
c86 44 0 1.26199e-19 $X=11.715 $Y=1.19
c87 15 0 1.67668e-19 $X=10.245 $Y=0.395
r88 43 44 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=11.7 $Y=1.505
+ $X2=11.7 $Y2=1.19
r89 42 44 10.9482 $w=2.98e-07 $l=2.85e-07 $layer=LI1_cond $X=11.7 $Y=0.905
+ $X2=11.7 $Y2=1.19
r90 36 41 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.36 $Y=1.59
+ $X2=11.17 $Y2=1.59
r91 35 43 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=11.55 $Y=1.59
+ $X2=11.7 $Y2=1.505
r92 35 36 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=11.55 $Y=1.59
+ $X2=11.36 $Y2=1.59
r93 34 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.36 $Y=0.82
+ $X2=11.17 $Y2=0.82
r94 33 42 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=11.55 $Y=0.82
+ $X2=11.7 $Y2=0.905
r95 33 34 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=11.55 $Y=0.82
+ $X2=11.36 $Y2=0.82
r96 29 41 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=11.17 $Y=1.675
+ $X2=11.17 $Y2=1.59
r97 29 31 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=11.17 $Y=1.675
+ $X2=11.17 $Y2=2.31
r98 25 39 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=11.17 $Y=0.735
+ $X2=11.17 $Y2=0.82
r99 25 27 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=11.17 $Y=0.735
+ $X2=11.17 $Y2=0.395
r100 24 38 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.41 $Y=1.59
+ $X2=10.22 $Y2=1.59
r101 23 41 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.98 $Y=1.59
+ $X2=11.17 $Y2=1.59
r102 23 24 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=10.98 $Y=1.59
+ $X2=10.41 $Y2=1.59
r103 21 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.98 $Y=0.82
+ $X2=11.17 $Y2=0.82
r104 21 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=10.98 $Y=0.82
+ $X2=10.41 $Y2=0.82
r105 17 38 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=10.22 $Y=1.675
+ $X2=10.22 $Y2=1.59
r106 17 19 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=10.22 $Y=1.675
+ $X2=10.22 $Y2=2.31
r107 13 22 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=10.22 $Y=0.735
+ $X2=10.41 $Y2=0.82
r108 13 15 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=10.22 $Y=0.735
+ $X2=10.22 $Y2=0.395
r109 4 41 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=11.05
+ $Y=1.485 $X2=11.195 $Y2=1.63
r110 4 31 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=11.05
+ $Y=1.485 $X2=11.195 $Y2=2.31
r111 3 38 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.1
+ $Y=1.485 $X2=10.245 $Y2=1.63
r112 3 19 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=10.1
+ $Y=1.485 $X2=10.245 $Y2=2.31
r113 2 27 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=11.01
+ $Y=0.235 $X2=11.195 $Y2=0.395
r114 1 15 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=10.06
+ $Y=0.235 $X2=10.245 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_4%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 49
+ 51 54 55 57 58 60 61 63 64 66 67 68 70 94 105 111 117 121
c179 121 0 2.71124e-20 $X=11.73 $Y=0
r180 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r181 117 118 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r182 111 114 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.38
r183 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r184 108 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=11.73 $Y2=0
r185 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r186 105 120 3.40825 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.58 $Y=0
+ $X2=11.77 $Y2=0
r187 105 107 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=11.58 $Y=0
+ $X2=11.27 $Y2=0
r188 104 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=11.27 $Y2=0
r189 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r190 101 104 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.35 $Y2=0
r191 101 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=8.51 $Y2=0
r192 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r193 98 117 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=8.87 $Y=0 $X2=8.66
+ $Y2=0
r194 98 100 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.87 $Y=0 $X2=9.43
+ $Y2=0
r195 97 118 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=8.51 $Y2=0
r196 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r197 94 117 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=8.45 $Y=0 $X2=8.66
+ $Y2=0
r198 94 96 116.128 $w=1.68e-07 $l=1.78e-06 $layer=LI1_cond $X=8.45 $Y=0 $X2=6.67
+ $Y2=0
r199 93 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r200 92 93 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r201 90 93 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=6.21 $Y2=0
r202 89 92 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.37 $Y=0 $X2=6.21
+ $Y2=0
r203 89 90 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r204 87 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r205 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r206 84 87 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.91 $Y2=0
r207 83 86 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r208 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r209 81 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r210 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r211 78 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r212 78 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r213 77 80 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r214 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r215 75 111 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=0.705 $Y2=0
r216 75 77 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r217 70 111 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.705 $Y2=0
r218 70 72 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r219 68 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r220 68 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r221 66 103 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=10.64 $Y=0
+ $X2=10.35 $Y2=0
r222 66 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.64 $Y=0
+ $X2=10.725 $Y2=0
r223 65 107 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=10.81 $Y=0
+ $X2=11.27 $Y2=0
r224 65 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.81 $Y=0
+ $X2=10.725 $Y2=0
r225 63 100 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=9.69 $Y=0 $X2=9.43
+ $Y2=0
r226 63 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.69 $Y=0 $X2=9.775
+ $Y2=0
r227 62 103 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=9.86 $Y=0
+ $X2=10.35 $Y2=0
r228 62 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.86 $Y=0 $X2=9.775
+ $Y2=0
r229 60 92 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=6.225 $Y=0 $X2=6.21
+ $Y2=0
r230 60 61 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.225 $Y=0 $X2=6.41
+ $Y2=0
r231 59 96 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.595 $Y=0 $X2=6.67
+ $Y2=0
r232 59 61 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.595 $Y=0 $X2=6.41
+ $Y2=0
r233 57 86 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.115 $Y=0
+ $X2=3.91 $Y2=0
r234 57 58 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.115 $Y=0 $X2=4.215
+ $Y2=0
r235 56 89 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.315 $Y=0 $X2=4.37
+ $Y2=0
r236 56 58 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.315 $Y=0 $X2=4.215
+ $Y2=0
r237 54 80 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.125 $Y=0 $X2=2.07
+ $Y2=0
r238 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=2.29
+ $Y2=0
r239 53 83 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.53
+ $Y2=0
r240 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.29
+ $Y2=0
r241 49 120 3.40825 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=11.665 $Y=0.085
+ $X2=11.77 $Y2=0
r242 49 51 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=11.665 $Y=0.085
+ $X2=11.665 $Y2=0.395
r243 45 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.725 $Y=0.085
+ $X2=10.725 $Y2=0
r244 45 47 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.725 $Y=0.085
+ $X2=10.725 $Y2=0.395
r245 41 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.775 $Y=0.085
+ $X2=9.775 $Y2=0
r246 41 43 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=9.775 $Y=0.085
+ $X2=9.775 $Y2=0.53
r247 37 117 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.66 $Y=0.085
+ $X2=8.66 $Y2=0
r248 37 39 10.0153 $w=4.18e-07 $l=3.65e-07 $layer=LI1_cond $X=8.66 $Y=0.085
+ $X2=8.66 $Y2=0.45
r249 33 61 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.41 $Y=0.085
+ $X2=6.41 $Y2=0
r250 33 35 10.4343 $w=3.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.41 $Y=0.085
+ $X2=6.41 $Y2=0.42
r251 29 58 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.215 $Y=0.085
+ $X2=4.215 $Y2=0
r252 29 31 15.25 $w=1.98e-07 $l=2.75e-07 $layer=LI1_cond $X=4.215 $Y=0.085
+ $X2=4.215 $Y2=0.36
r253 25 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=0.085
+ $X2=2.29 $Y2=0
r254 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.29 $Y=0.085
+ $X2=2.29 $Y2=0.36
r255 8 51 182 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=1 $X=11.53
+ $Y=0.235 $X2=11.665 $Y2=0.395
r256 7 47 182 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_NDIFF $count=1 $X=10.53
+ $Y=0.235 $X2=10.725 $Y2=0.395
r257 6 43 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=9.64
+ $Y=0.235 $X2=9.775 $Y2=0.53
r258 5 39 182 $w=1.7e-07 $l=2.93258e-07 $layer=licon1_NDIFF $count=1 $X=8.6
+ $Y=0.235 $X2=8.785 $Y2=0.45
r259 4 35 182 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_NDIFF $count=1 $X=6.175
+ $Y=0.235 $X2=6.48 $Y2=0.42
r260 3 31 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=3.985
+ $Y=0.235 $X2=4.2 $Y2=0.36
r261 2 27 182 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.29 $Y2=0.36
r262 1 114 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

