* File: sky130_fd_sc_hdll__and4bb_4.pex.spice
* Created: Wed Sep  2 08:23:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND4BB_4%B_N 2 3 5 8 10 11 12 17
c39 8 0 1.38622e-19 $X=0.52 $Y=0.445
c40 2 0 1.7526e-19 $X=0.495 $Y=1.89
r41 17 20 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.16
+ $X2=0.54 $Y2=1.325
r42 17 19 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.16
+ $X2=0.54 $Y2=0.995
r43 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.16 $X2=0.515 $Y2=1.16
r44 11 12 9.79577 $w=3.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.63 $Y=1.19
+ $X2=0.63 $Y2=1.53
r45 11 18 0.864332 $w=3.98e-07 $l=3e-08 $layer=LI1_cond $X=0.63 $Y=1.19 $X2=0.63
+ $Y2=1.16
r46 10 18 8.93143 $w=3.98e-07 $l=3.1e-07 $layer=LI1_cond $X=0.63 $Y=0.85
+ $X2=0.63 $Y2=1.16
r47 8 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.445
+ $X2=0.52 $Y2=0.995
r48 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r49 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.89 $X2=0.495
+ $Y2=1.99
r50 2 20 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.495 $Y=1.89
+ $X2=0.495 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_4%A_184_21# 1 2 3 12 14 16 19 21 23 26 28
+ 30 33 35 37 38 44 46 47 48 49 53 56 57 58 59 62 71
c149 71 0 1.99894e-19 $X=2.405 $Y=1.217
r150 71 72 3.34722 $w=3.6e-07 $l=2.5e-08 $layer=POLY_cond $X=2.405 $Y=1.217
+ $X2=2.43 $Y2=1.217
r151 68 69 3.34722 $w=3.6e-07 $l=2.5e-08 $layer=POLY_cond $X=1.935 $Y=1.217
+ $X2=1.96 $Y2=1.217
r152 67 68 59.5806 $w=3.6e-07 $l=4.45e-07 $layer=POLY_cond $X=1.49 $Y=1.217
+ $X2=1.935 $Y2=1.217
r153 66 67 3.34722 $w=3.6e-07 $l=2.5e-08 $layer=POLY_cond $X=1.465 $Y=1.217
+ $X2=1.49 $Y2=1.217
r154 65 66 59.5806 $w=3.6e-07 $l=4.45e-07 $layer=POLY_cond $X=1.02 $Y=1.217
+ $X2=1.465 $Y2=1.217
r155 64 65 3.34722 $w=3.6e-07 $l=2.5e-08 $layer=POLY_cond $X=0.995 $Y=1.217
+ $X2=1.02 $Y2=1.217
r156 57 62 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=4.71 $Y=0.385
+ $X2=4.885 $Y2=0.385
r157 57 58 98.8396 $w=1.68e-07 $l=1.515e-06 $layer=LI1_cond $X=4.71 $Y=0.385
+ $X2=3.195 $Y2=0.385
r158 55 58 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.085 $Y=0.47
+ $X2=3.195 $Y2=0.385
r159 55 56 7.59565 $w=2.18e-07 $l=1.45e-07 $layer=LI1_cond $X=3.085 $Y=0.47
+ $X2=3.085 $Y2=0.615
r160 51 53 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=3.275 $Y=1.63
+ $X2=4.385 $Y2=1.63
r161 49 51 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.7 $Y=1.63
+ $X2=3.275 $Y2=1.63
r162 47 56 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.975 $Y=0.7
+ $X2=3.085 $Y2=0.615
r163 47 48 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.975 $Y=0.7
+ $X2=2.7 $Y2=0.7
r164 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.615 $Y=1.545
+ $X2=2.7 $Y2=1.63
r165 45 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=1.245
+ $X2=2.615 $Y2=1.16
r166 45 46 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.615 $Y=1.245
+ $X2=2.615 $Y2=1.545
r167 44 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=1.075
+ $X2=2.615 $Y2=1.16
r168 43 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.615 $Y=0.785
+ $X2=2.7 $Y2=0.7
r169 43 44 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.615 $Y=0.785
+ $X2=2.615 $Y2=1.075
r170 41 71 45.5222 $w=3.6e-07 $l=3.4e-07 $layer=POLY_cond $X=2.065 $Y=1.217
+ $X2=2.405 $Y2=1.217
r171 41 69 14.0583 $w=3.6e-07 $l=1.05e-07 $layer=POLY_cond $X=2.065 $Y=1.217
+ $X2=1.96 $Y2=1.217
r172 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.065
+ $Y=1.16 $X2=2.065 $Y2=1.16
r173 38 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=1.16
+ $X2=2.615 $Y2=1.16
r174 38 40 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.53 $Y=1.16
+ $X2=2.065 $Y2=1.16
r175 35 72 18.9685 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.43 $Y=1.41
+ $X2=2.43 $Y2=1.217
r176 35 37 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.43 $Y=1.41
+ $X2=2.43 $Y2=1.985
r177 31 71 23.3057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.405 $Y=1.025
+ $X2=2.405 $Y2=1.217
r178 31 33 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.405 $Y=1.025
+ $X2=2.405 $Y2=0.56
r179 28 69 18.9685 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.96 $Y=1.41
+ $X2=1.96 $Y2=1.217
r180 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.96 $Y=1.41
+ $X2=1.96 $Y2=1.985
r181 24 68 23.3057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.935 $Y=1.025
+ $X2=1.935 $Y2=1.217
r182 24 26 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.935 $Y=1.025
+ $X2=1.935 $Y2=0.56
r183 21 67 18.9685 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.49 $Y=1.41
+ $X2=1.49 $Y2=1.217
r184 21 23 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.49 $Y=1.41
+ $X2=1.49 $Y2=1.985
r185 17 66 23.3057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.465 $Y=1.025
+ $X2=1.465 $Y2=1.217
r186 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.465 $Y=1.025
+ $X2=1.465 $Y2=0.56
r187 14 65 18.9685 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.02 $Y=1.41
+ $X2=1.02 $Y2=1.217
r188 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.02 $Y=1.41
+ $X2=1.02 $Y2=1.985
r189 10 64 23.3057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.995 $Y=1.025
+ $X2=0.995 $Y2=1.217
r190 10 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.995 $Y=1.025
+ $X2=0.995 $Y2=0.56
r191 3 53 600 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=4.22
+ $Y=1.485 $X2=4.385 $Y2=1.63
r192 2 51 600 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=3.07
+ $Y=1.485 $X2=3.275 $Y2=1.63
r193 1 62 91 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_NDIFF $count=2 $X=4.71
+ $Y=0.235 $X2=4.895 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_4%D 1 3 4 6 7
c35 7 0 1.99894e-19 $X=2.995 $Y=1.19
c36 4 0 1.0531e-19 $X=2.98 $Y=1.41
r37 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.015
+ $Y=1.16 $X2=3.015 $Y2=1.16
r38 4 10 46.6797 $w=3.23e-07 $l=2.8592e-07 $layer=POLY_cond $X=2.98 $Y=1.41
+ $X2=3.057 $Y2=1.16
r39 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.98 $Y=1.41 $X2=2.98
+ $Y2=1.985
r40 1 10 38.5615 $w=3.23e-07 $l=2.09893e-07 $layer=POLY_cond $X=2.955 $Y=0.995
+ $X2=3.057 $Y2=1.16
r41 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.955 $Y=0.995
+ $X2=2.955 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_4%C 1 3 4 6 7 8 17
r33 13 17 7.80599 $w=4.73e-07 $l=3.1e-07 $layer=LI1_cond $X=3.602 $Y=1.16
+ $X2=3.602 $Y2=0.85
r34 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.635
+ $Y=1.16 $X2=3.635 $Y2=1.16
r35 8 13 0.755418 $w=4.73e-07 $l=3e-08 $layer=LI1_cond $X=3.602 $Y=1.19
+ $X2=3.602 $Y2=1.16
r36 7 17 1.51084 $w=4.73e-07 $l=6e-08 $layer=LI1_cond $X=3.602 $Y=0.79 $X2=3.602
+ $Y2=0.85
r37 4 12 46.0897 $w=3.39e-07 $l=2.90259e-07 $layer=POLY_cond $X=3.545 $Y=1.41
+ $X2=3.632 $Y2=1.16
r38 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.545 $Y=1.41
+ $X2=3.545 $Y2=1.985
r39 1 12 38.6704 $w=3.39e-07 $l=2.13787e-07 $layer=POLY_cond $X=3.52 $Y=0.995
+ $X2=3.632 $Y2=1.16
r40 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.52 $Y=0.995 $X2=3.52
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_4%A_27_47# 1 2 7 9 10 12 14 17 19 21 24 26
+ 29 31
c92 31 0 1.00528e-19 $X=4.165 $Y=1.16
r93 31 34 6.80989 $w=2.18e-07 $l=1.3e-07 $layer=LI1_cond $X=4.19 $Y=1.16
+ $X2=4.19 $Y2=1.29
r94 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.165
+ $Y=1.16 $X2=4.165 $Y2=1.16
r95 26 28 8.55024 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.215 $Y=0.42
+ $X2=0.215 $Y2=0.585
r96 23 24 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.855 $Y=1.375
+ $X2=4.855 $Y2=1.915
r97 22 34 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.3 $Y=1.29 $X2=4.19
+ $Y2=1.29
r98 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.77 $Y=1.29
+ $X2=4.855 $Y2=1.375
r99 21 22 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=4.77 $Y=1.29 $X2=4.3
+ $Y2=1.29
r100 20 29 2.24312 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=2 $X2=0.215
+ $Y2=2
r101 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.77 $Y=2
+ $X2=4.855 $Y2=1.915
r102 19 20 288.69 $w=1.68e-07 $l=4.425e-06 $layer=LI1_cond $X=4.77 $Y=2
+ $X2=0.345 $Y2=2
r103 15 29 4.18896 $w=2.17e-07 $l=8.5e-08 $layer=LI1_cond $X=0.215 $Y=2.085
+ $X2=0.215 $Y2=2
r104 15 17 9.52982 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=0.215 $Y=2.085
+ $X2=0.215 $Y2=2.3
r105 14 29 4.18896 $w=2.17e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.172 $Y=1.915
+ $X2=0.215 $Y2=2
r106 14 28 84.2909 $w=1.73e-07 $l=1.33e-06 $layer=LI1_cond $X=0.172 $Y=1.915
+ $X2=0.172 $Y2=0.585
r107 10 32 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=4.13 $Y=1.41
+ $X2=4.19 $Y2=1.16
r108 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.13 $Y=1.41
+ $X2=4.13 $Y2=1.985
r109 7 32 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=4.105 $Y=0.995
+ $X2=4.19 $Y2=1.16
r110 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.105 $Y=0.995
+ $X2=4.105 $Y2=0.56
r111 2 17 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
r112 1 26 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_4%A_912_21# 1 2 9 11 13 15 19 20 21 22 23
+ 24 27 31
c70 15 0 1.00528e-19 $X=4.66 $Y=1.217
r71 29 31 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.18 $Y=2.085
+ $X2=6.18 $Y2=2.3
r72 25 27 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.18 $Y=0.655
+ $X2=6.18 $Y2=0.42
r73 23 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.095 $Y=2
+ $X2=6.18 $Y2=2.085
r74 23 24 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=6.095 $Y=2 $X2=5.53
+ $Y2=2
r75 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.095 $Y=0.74
+ $X2=6.18 $Y2=0.655
r76 21 22 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=6.095 $Y=0.74
+ $X2=5.53 $Y2=0.74
r77 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.445
+ $Y=1.16 $X2=5.445 $Y2=1.16
r78 17 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.445 $Y=1.915
+ $X2=5.53 $Y2=2
r79 17 19 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=5.445 $Y=1.915
+ $X2=5.445 $Y2=1.16
r80 16 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.445 $Y=0.825
+ $X2=5.53 $Y2=0.74
r81 16 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.445 $Y=0.825
+ $X2=5.445 $Y2=1.16
r82 14 20 112.935 $w=3.5e-07 $l=6.85e-07 $layer=POLY_cond $X=4.76 $Y=1.2
+ $X2=5.445 $Y2=1.2
r83 14 15 4.60329 $w=3.5e-07 $l=1.08167e-07 $layer=POLY_cond $X=4.76 $Y=1.2
+ $X2=4.66 $Y2=1.217
r84 11 15 36.1676 $w=1.65e-07 $l=1.93e-07 $layer=POLY_cond $X=4.66 $Y=1.41
+ $X2=4.66 $Y2=1.217
r85 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.66 $Y=1.41
+ $X2=4.66 $Y2=1.985
r86 7 15 36.1676 $w=1.65e-07 $l=2.04118e-07 $layer=POLY_cond $X=4.635 $Y=1.025
+ $X2=4.66 $Y2=1.217
r87 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.635 $Y=1.025
+ $X2=4.635 $Y2=0.56
r88 2 31 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=6.035
+ $Y=2.065 $X2=6.18 $Y2=2.3
r89 1 27 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=5.995
+ $Y=0.235 $X2=6.18 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_4%A_N 3 6 7 9 10 11 15
r27 15 18 37.7576 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=6.025 $Y=1.16
+ $X2=6.025 $Y2=1.325
r28 15 17 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=6.025 $Y=1.16
+ $X2=6.025 $Y2=0.995
r29 10 11 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=6.14 $Y=1.16
+ $X2=6.14 $Y2=1.53
r30 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.02
+ $Y=1.16 $X2=6.02 $Y2=1.16
r31 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.945 $Y=1.99
+ $X2=5.945 $Y2=2.275
r32 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=5.945 $Y=1.89 $X2=5.945
+ $Y2=1.99
r33 6 18 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=5.945 $Y=1.89
+ $X2=5.945 $Y2=1.325
r34 3 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.92 $Y=0.445
+ $X2=5.92 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_4%VPWR 1 2 3 4 5 16 20 25 28 29 31 36 41 46
+ 51 52 55 62 69 76 81
r90 79 83 3.1533 $w=5.48e-07 $l=1.45e-07 $layer=LI1_cond $X=4.83 $Y=2.53
+ $X2=4.975 $Y2=2.53
r91 79 81 6.67868 $w=5.48e-07 $l=2e-08 $layer=LI1_cond $X=4.83 $Y=2.53 $X2=4.81
+ $Y2=2.53
r92 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r93 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r94 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r95 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r96 69 72 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=2.64 $Y=2.34
+ $X2=2.64 $Y2=2.72
r97 66 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r98 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r99 62 65 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=1.7 $Y=2.34 $X2=1.7
+ $Y2=2.72
r100 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r101 55 58 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=2.34
+ $X2=0.705 $Y2=2.72
r102 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r103 49 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r104 49 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r105 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r106 46 83 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=5.085 $Y=2.53
+ $X2=4.975 $Y2=2.53
r107 46 48 4.45811 $w=5.48e-07 $l=2.05e-07 $layer=LI1_cond $X=5.085 $Y=2.53
+ $X2=5.29 $Y2=2.53
r108 45 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r109 45 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r110 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r111 42 72 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.83 $Y=2.72
+ $X2=2.64 $Y2=2.72
r112 42 44 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.83 $Y=2.72
+ $X2=3.45 $Y2=2.72
r113 41 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.68 $Y=2.72
+ $X2=3.845 $Y2=2.72
r114 41 44 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.68 $Y=2.72
+ $X2=3.45 $Y2=2.72
r115 40 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r116 40 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r117 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r118 37 58 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r119 37 39 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r120 36 65 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.51 $Y=2.72 $X2=1.7
+ $Y2=2.72
r121 36 39 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.51 $Y=2.72
+ $X2=1.15 $Y2=2.72
r122 31 58 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r123 31 33 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r124 29 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r125 29 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r126 28 51 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=5.82 $Y=2.72
+ $X2=6.21 $Y2=2.72
r127 27 28 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.655 $Y=2.53
+ $X2=5.82 $Y2=2.53
r128 25 48 5.54545 $w=5.48e-07 $l=2.55e-07 $layer=LI1_cond $X=5.545 $Y=2.53
+ $X2=5.29 $Y2=2.53
r129 25 27 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=5.545 $Y=2.53
+ $X2=5.655 $Y2=2.53
r130 23 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.01 $Y=2.72
+ $X2=3.845 $Y2=2.72
r131 23 81 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=4.01 $Y=2.72 $X2=4.81
+ $Y2=2.72
r132 18 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.845 $Y=2.635
+ $X2=3.845 $Y2=2.72
r133 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.845 $Y=2.635
+ $X2=3.845 $Y2=2.34
r134 17 65 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.89 $Y=2.72 $X2=1.7
+ $Y2=2.72
r135 16 72 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.45 $Y=2.72
+ $X2=2.64 $Y2=2.72
r136 16 17 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.45 $Y=2.72
+ $X2=1.89 $Y2=2.72
r137 5 83 400 $w=1.7e-07 $l=9.60937e-07 $layer=licon1_PDIFF $count=1 $X=4.75
+ $Y=1.485 $X2=4.975 $Y2=2.34
r138 5 27 400 $w=1.7e-07 $l=1.26206e-06 $layer=licon1_PDIFF $count=1 $X=4.75
+ $Y=1.485 $X2=5.655 $Y2=2.34
r139 4 20 600 $w=1.7e-07 $l=9.54241e-07 $layer=licon1_PDIFF $count=1 $X=3.635
+ $Y=1.485 $X2=3.845 $Y2=2.34
r140 3 69 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.52
+ $Y=1.485 $X2=2.665 $Y2=2.34
r141 2 62 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.485 $X2=1.725 $Y2=2.34
r142 1 55 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.065 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_4%X 1 2 3 4 15 17 21 25 27 28 29 36 38 44
c49 38 0 3.13882e-19 $X=1.155 $Y=0.85
c50 21 0 1.0531e-19 $X=2.195 $Y=1.63
r51 36 44 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.175 $Y=1.545
+ $X2=1.175 $Y2=1.53
r52 35 38 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=1.175 $Y=0.82
+ $X2=1.175 $Y2=0.85
r53 29 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=0.735
+ $X2=1.175 $Y2=0.82
r54 29 38 0.942908 $w=3.28e-07 $l=2.7e-08 $layer=LI1_cond $X=1.175 $Y=0.877
+ $X2=1.175 $Y2=0.85
r55 28 36 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=1.63
+ $X2=1.175 $Y2=1.545
r56 28 44 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.175 $Y=1.495
+ $X2=1.175 $Y2=1.53
r57 27 28 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.175 $Y=1.19
+ $X2=1.175 $Y2=1.495
r58 27 29 10.9307 $w=3.28e-07 $l=3.13e-07 $layer=LI1_cond $X=1.175 $Y=1.19
+ $X2=1.175 $Y2=0.877
r59 23 25 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.195 $Y=0.65
+ $X2=2.195 $Y2=0.42
r60 19 28 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.34 $Y=1.63
+ $X2=1.175 $Y2=1.63
r61 19 21 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=1.34 $Y=1.63
+ $X2=2.195 $Y2=1.63
r62 18 29 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.34 $Y=0.735
+ $X2=1.175 $Y2=0.735
r63 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.11 $Y=0.735
+ $X2=2.195 $Y2=0.65
r64 17 18 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.11 $Y=0.735
+ $X2=1.34 $Y2=0.735
r65 13 29 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.255 $Y=0.65
+ $X2=1.175 $Y2=0.735
r66 13 15 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.255 $Y=0.65
+ $X2=1.255 $Y2=0.42
r67 4 21 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=1.485 $X2=2.195 $Y2=1.63
r68 3 28 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.11
+ $Y=1.485 $X2=1.255 $Y2=1.63
r69 2 25 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=2.01
+ $Y=0.235 $X2=2.195 $Y2=0.42
r70 1 15 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.235 $X2=1.255 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_4%VGND 1 2 3 4 17 21 23 27 31 34 35 36 38
+ 51 52 55 58 61 64
r100 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r101 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r102 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r103 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r104 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r105 49 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r106 48 49 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r107 46 49 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.99 $Y=0 $X2=5.29
+ $Y2=0
r108 46 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r109 45 48 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.99 $Y=0 $X2=5.29
+ $Y2=0
r110 45 46 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r111 43 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.635
+ $Y2=0
r112 43 45 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.99
+ $Y2=0
r113 42 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r114 42 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r115 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r116 39 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.785
+ $Y2=0
r117 39 41 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.15
+ $Y2=0
r118 38 58 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.51 $Y=0 $X2=1.7
+ $Y2=0
r119 38 41 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.51 $Y=0 $X2=1.15
+ $Y2=0
r120 36 56 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r121 36 64 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r122 34 48 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=5.385 $Y=0 $X2=5.29
+ $Y2=0
r123 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.385 $Y=0 $X2=5.55
+ $Y2=0
r124 33 51 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.715 $Y=0
+ $X2=6.21 $Y2=0
r125 33 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.715 $Y=0 $X2=5.55
+ $Y2=0
r126 29 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.55 $Y=0.085
+ $X2=5.55 $Y2=0
r127 29 31 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.55 $Y=0.085
+ $X2=5.55 $Y2=0.38
r128 25 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=0.085
+ $X2=2.635 $Y2=0
r129 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.635 $Y=0.085
+ $X2=2.635 $Y2=0.36
r130 24 58 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.7
+ $Y2=0
r131 23 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.635
+ $Y2=0
r132 23 24 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=1.89
+ $Y2=0
r133 19 58 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0
r134 19 21 9.09823 $w=3.78e-07 $l=3e-07 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0.385
r135 15 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0
r136 15 17 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0.38
r137 4 31 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=5.385
+ $Y=0.235 $X2=5.55 $Y2=0.38
r138 3 27 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.48
+ $Y=0.235 $X2=2.635 $Y2=0.36
r139 2 21 182 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_NDIFF $count=1 $X=1.54
+ $Y=0.235 $X2=1.725 $Y2=0.385
r140 1 17 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.785 $Y2=0.38
.ends

