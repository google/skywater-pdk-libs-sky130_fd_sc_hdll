* File: sky130_fd_sc_hdll__isobufsrc_2.pex.spice
* Created: Thu Aug 27 19:09:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%SLEEP 1 3 4 6 7 9 10 12 13 20 24
r36 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.01 $Y2=1.202
r37 18 20 43.1263 $w=3.8e-07 $l=3.4e-07 $layer=POLY_cond $X=0.645 $Y=1.202
+ $X2=0.985 $Y2=1.202
r38 18 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.645
+ $Y=1.16 $X2=0.645 $Y2=1.16
r39 16 18 16.4895 $w=3.8e-07 $l=1.3e-07 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.645 $Y2=1.202
r40 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.49 $Y=1.202
+ $X2=0.515 $Y2=1.202
r41 13 24 2.90476 $w=2.08e-07 $l=5.5e-08 $layer=LI1_cond $X=0.7 $Y=1.17
+ $X2=0.645 $Y2=1.17
r42 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=1.202
r43 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=0.56
r44 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r45 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r46 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r47 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r48 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.202
r49 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%A_271_21# 1 2 7 9 10 12 13 15 16 18 19
+ 24 27 30 32 33 38 42 44 47
c81 30 0 2.92282e-20 $X=2.522 $Y=1.075
c82 16 0 1.04966e-19 $X=1.95 $Y=0.995
r83 45 47 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.545 $Y=1.53
+ $X2=2.68 $Y2=1.53
r84 36 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=1.615
+ $X2=2.68 $Y2=1.53
r85 36 38 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.68 $Y=1.615
+ $X2=2.68 $Y2=2.28
r86 33 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=0.725
+ $X2=2.68 $Y2=0.81
r87 33 35 3.22941 $w=1.7e-07 $l=4.5e-08 $layer=LI1_cond $X=2.68 $Y=0.725
+ $X2=2.68 $Y2=0.68
r88 32 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=1.445
+ $X2=2.545 $Y2=1.53
r89 31 44 4.65272 $w=1.92e-07 $l=9.58123e-08 $layer=LI1_cond $X=2.545 $Y=1.245
+ $X2=2.522 $Y2=1.16
r90 31 32 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.545 $Y=1.245
+ $X2=2.545 $Y2=1.445
r91 30 44 4.65272 $w=1.92e-07 $l=8.5e-08 $layer=LI1_cond $X=2.522 $Y=1.075
+ $X2=2.522 $Y2=1.16
r92 29 42 10.308 $w=1.68e-07 $l=1.58e-07 $layer=LI1_cond $X=2.522 $Y=0.81
+ $X2=2.68 $Y2=0.81
r93 29 30 9.64836 $w=2.13e-07 $l=1.8e-07 $layer=LI1_cond $X=2.522 $Y=0.895
+ $X2=2.522 $Y2=1.075
r94 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.24
+ $Y=1.16 $X2=2.24 $Y2=1.16
r95 24 44 1.79375 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.415 $Y=1.16
+ $X2=2.522 $Y2=1.16
r96 24 26 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.415 $Y=1.16
+ $X2=2.24 $Y2=1.16
r97 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.925 $Y=1.202
+ $X2=1.95 $Y2=1.202
r98 21 22 59.6158 $w=3.8e-07 $l=4.7e-07 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.925 $Y2=1.202
r99 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.43 $Y=1.202
+ $X2=1.455 $Y2=1.202
r100 19 27 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=2.025 $Y=1.16
+ $X2=2.24 $Y2=1.16
r101 19 23 10.4773 $w=3.8e-07 $l=9.3675e-08 $layer=POLY_cond $X=2.025 $Y=1.16
+ $X2=1.95 $Y2=1.202
r102 16 23 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=1.202
r103 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=0.56
r104 13 22 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r105 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r106 10 21 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r107 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r108 7 20 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=1.202
r109 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=0.56
r110 2 38 600 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=2.555
+ $Y=2.065 $X2=2.68 $Y2=2.28
r111 1 35 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=2.555
+ $Y=0.465 $X2=2.68 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%A 3 5 6 8 9 10 11 18 20 30
c35 18 0 2.92282e-20 $X=2.965 $Y=1.16
r36 18 21 37.7183 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=2.982 $Y=1.16
+ $X2=2.982 $Y2=1.325
r37 18 20 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=2.982 $Y=1.16
+ $X2=2.982 $Y2=0.995
r38 18 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.965
+ $Y=1.16 $X2=2.965 $Y2=1.16
r39 10 11 18.2247 $w=2.13e-07 $l=3.4e-07 $layer=LI1_cond $X=3.447 $Y=1.53
+ $X2=3.447 $Y2=1.87
r40 9 30 13.6618 $w=3.78e-07 $l=3.75e-07 $layer=LI1_cond $X=3.34 $Y=1.17
+ $X2=2.965 $Y2=1.17
r41 9 10 9.86223 $w=3.83e-07 $l=2.55e-07 $layer=LI1_cond $X=3.447 $Y=1.275
+ $X2=3.447 $Y2=1.53
r42 6 8 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.915 $Y=1.99
+ $X2=2.915 $Y2=2.275
r43 5 6 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.915 $Y=1.89 $X2=2.915
+ $Y2=1.99
r44 5 21 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=2.915 $Y=1.89
+ $X2=2.915 $Y2=1.325
r45 3 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.89 $Y=0.675
+ $X2=2.89 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%A_27_297# 1 2 3 10 12 14 16 17 18 22
+ 24 25
r44 25 34 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=2.295
+ $X2=2.18 $Y2=2.38
r45 24 32 5.95937 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=2.18 $Y=2.035
+ $X2=2.18 $Y2=1.89
r46 24 25 10.3322 $w=2.88e-07 $l=2.6e-07 $layer=LI1_cond $X=2.18 $Y=2.035
+ $X2=2.18 $Y2=2.295
r47 22 32 11.7504 $w=2.53e-07 $l=2.6e-07 $layer=LI1_cond $X=2.162 $Y=1.63
+ $X2=2.162 $Y2=1.89
r48 19 31 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=2.38
+ $X2=1.22 $Y2=2.38
r49 18 34 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.035 $Y=2.38
+ $X2=2.18 $Y2=2.38
r50 18 19 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.035 $Y=2.38
+ $X2=1.345 $Y2=2.38
r51 17 31 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=2.295
+ $X2=1.22 $Y2=2.38
r52 16 29 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.22 $Y=1.655
+ $X2=1.22 $Y2=1.55
r53 16 17 29.5025 $w=2.48e-07 $l=6.4e-07 $layer=LI1_cond $X=1.22 $Y=1.655
+ $X2=1.22 $Y2=2.295
r54 15 27 4.35048 $w=2.1e-07 $l=1.6e-07 $layer=LI1_cond $X=0.405 $Y=1.55
+ $X2=0.245 $Y2=1.55
r55 14 29 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=1.55
+ $X2=1.22 $Y2=1.55
r56 14 15 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=1.55
+ $X2=0.405 $Y2=1.55
r57 10 27 2.855 $w=3.2e-07 $l=1.05e-07 $layer=LI1_cond $X=0.245 $Y=1.655
+ $X2=0.245 $Y2=1.55
r58 10 12 23.2289 $w=3.18e-07 $l=6.45e-07 $layer=LI1_cond $X=0.245 $Y=1.655
+ $X2=0.245 $Y2=2.3
r59 3 34 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=2.31
r60 3 22 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=1.63
r61 2 31 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.3
r62 2 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.62
r63 1 27 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r64 1 12 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%VPWR 1 2 11 15 18 19 20 30 31 34 37
r40 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r41 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r42 28 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r43 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r44 25 28 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 25 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r46 24 27 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r47 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r48 22 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=0.75 $Y2=2.72
r49 22 24 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=1.15 $Y2=2.72
r50 20 35 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r51 20 37 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r52 18 27 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.025 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 18 19 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.025 $Y=2.72
+ $X2=3.15 $Y2=2.72
r54 17 30 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.275 $Y=2.72
+ $X2=3.45 $Y2=2.72
r55 17 19 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.275 $Y=2.72
+ $X2=3.15 $Y2=2.72
r56 13 19 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.15 $Y=2.635
+ $X2=3.15 $Y2=2.72
r57 13 15 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=3.15 $Y=2.635
+ $X2=3.15 $Y2=2.31
r58 9 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r59 9 11 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2
r60 2 15 600 $w=1.7e-07 $l=3.09112e-07 $layer=licon1_PDIFF $count=1 $X=3.005
+ $Y=2.065 $X2=3.15 $Y2=2.31
r61 1 11 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%X 1 2 3 12 14 15 18 21 22 25
c46 21 0 1.04966e-19 $X=1.665 $Y=0.81
r47 22 25 3.63929 $w=3.78e-07 $l=1.2e-07 $layer=LI1_cond $X=1.665 $Y=0.51
+ $X2=1.665 $Y2=0.39
r48 20 22 6.5204 $w=3.78e-07 $l=2.15e-07 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.51
r49 20 21 2.84813 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.81
r50 16 21 2.84813 $w=3.35e-07 $l=8.74643e-08 $layer=LI1_cond $X=1.67 $Y=0.895
+ $X2=1.665 $Y2=0.81
r51 16 18 28.8111 $w=2.88e-07 $l=7.25e-07 $layer=LI1_cond $X=1.67 $Y=0.895
+ $X2=1.67 $Y2=1.62
r52 14 21 3.86674 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.475 $Y=0.81
+ $X2=1.665 $Y2=0.81
r53 14 15 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.475 $Y=0.81
+ $X2=0.915 $Y2=0.81
r54 10 15 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.915 $Y2=0.81
r55 10 12 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.725 $Y2=0.39
r56 3 18 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=1.62
r57 2 25 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.505
+ $Y=0.235 $X2=1.69 $Y2=0.39
r58 1 12 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%VGND 1 2 3 4 13 15 17 21 25 29 32 33
+ 35 36 37 47 48 54
r54 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r55 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r56 45 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r57 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r58 42 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r59 42 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r60 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r61 39 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.22
+ $Y2=0
r62 39 41 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=2.07
+ $Y2=0
r63 37 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r64 37 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r65 35 44 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.025 $Y=0 $X2=2.99
+ $Y2=0
r66 35 36 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=3.025 $Y=0 $X2=3.152
+ $Y2=0
r67 34 47 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.28 $Y=0 $X2=3.45
+ $Y2=0
r68 34 36 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=3.28 $Y=0 $X2=3.152
+ $Y2=0
r69 32 41 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.07
+ $Y2=0
r70 32 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.16
+ $Y2=0
r71 31 44 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.99
+ $Y2=0
r72 31 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.16
+ $Y2=0
r73 27 36 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=3.152 $Y=0.085
+ $X2=3.152 $Y2=0
r74 27 29 26.8903 $w=2.53e-07 $l=5.95e-07 $layer=LI1_cond $X=3.152 $Y=0.085
+ $X2=3.152 $Y2=0.68
r75 23 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0
r76 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0.39
r77 19 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r78 19 21 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.39
r79 18 51 4.33083 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r80 17 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.22
+ $Y2=0
r81 17 18 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=0 $X2=0.365
+ $Y2=0
r82 13 51 3.02922 $w=2.8e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.182 $Y2=0
r83 13 15 12.5534 $w=2.78e-07 $l=3.05e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.225 $Y2=0.39
r84 4 29 182 $w=1.7e-07 $l=2.93258e-07 $layer=licon1_NDIFF $count=1 $X=2.965
+ $Y=0.465 $X2=3.15 $Y2=0.68
r85 3 25 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.025
+ $Y=0.235 $X2=2.16 $Y2=0.39
r86 2 21 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.235 $X2=1.22 $Y2=0.39
r87 1 15 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

