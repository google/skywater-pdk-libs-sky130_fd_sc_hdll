* File: sky130_fd_sc_hdll__o2bb2a_2.spice
* Created: Wed Sep  2 08:46:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o2bb2a_2.pex.spice"
.subckt sky130_fd_sc_hdll__o2bb2a_2  VNB VPB A1_N A2_N B2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1003 N_X_M1003_d N_A_84_21#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.18525 PD=0.97 PS=1.87 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1011 N_X_M1003_d N_A_84_21#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.136196 PD=0.97 PS=1.24533 NRD=0 NRS=7.38 M=1 R=4.33333
+ SA=75000.7 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1012 A_313_47# N_A1_N_M1012_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.0880037 PD=0.8 PS=0.804673 NRD=38.568 NRS=15.708 M=1 R=2.8
+ SA=75001.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1000 N_A_321_369#_M1000_d N_A2_N_M1000_g A_313_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.126 AS=0.0798 PD=1.44 PS=0.8 NRD=9.996 NRS=38.568 M=1 R=2.8 SA=75001.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_627_47#_M1004_d N_A_321_369#_M1004_g N_A_84_21#_M1004_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0714 AS=0.1218 PD=0.76 PS=1.42 NRD=4.284 NRS=7.14 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_B2_M1010_g N_A_627_47#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.06825 AS=0.0714 PD=0.745 PS=0.76 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.7
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_627_47#_M1002_d N_B1_M1002_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.06825 PD=1.37 PS=0.745 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_84_21#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.295 AS=0.145 PD=2.59 PS=1.29 NRD=1.9503 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1013_d N_A_84_21#_M1013_g N_X_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.191707 AS=0.145 PD=1.64024 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1001 N_A_321_369#_M1001_d N_A1_N_M1001_g N_VPWR_M1013_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1826 AS=0.122693 PD=1.43 PS=1.04976 NRD=70.8806 NRS=18.4589 M=1
+ R=3.55556 SA=90001.2 SB=90002.7 A=0.1152 P=1.64 MULT=1
MM1008 N_VPWR_M1008_d N_A2_N_M1008_g N_A_321_369#_M1001_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.2336 AS=0.1826 PD=1.37 PS=1.43 NRD=64.6357 NRS=70.8806 M=1
+ R=3.55556 SA=90001.8 SB=90002.1 A=0.1152 P=1.64 MULT=1
MM1005 N_A_84_21#_M1005_d N_A_321_369#_M1005_g N_VPWR_M1008_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.0992 AS=0.2336 PD=0.95 PS=1.37 NRD=1.5366 NRS=73.8553 M=1
+ R=3.55556 SA=90002.7 SB=90001.2 A=0.1152 P=1.64 MULT=1
MM1009 A_723_369# N_B2_M1009_g N_A_84_21#_M1005_d VPB PHIGHVT L=0.18 W=0.64
+ AD=0.1104 AS=0.0992 PD=0.985 PS=0.95 NRD=36.1495 NRS=7.683 M=1 R=3.55556
+ SA=90003.2 SB=90000.7 A=0.1152 P=1.64 MULT=1
MM1006 N_VPWR_M1006_d N_B1_M1006_g A_723_369# VPB PHIGHVT L=0.18 W=0.64
+ AD=0.1792 AS=0.1104 PD=1.84 PS=0.985 NRD=4.6098 NRS=36.1495 M=1 R=3.55556
+ SA=90003.7 SB=90000.2 A=0.1152 P=1.64 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
*
.include "sky130_fd_sc_hdll__o2bb2a_2.pxi.spice"
*
.ends
*
*
