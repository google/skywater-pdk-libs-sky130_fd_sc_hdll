# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hdll__tap
  CLASS BLOCK ;
  FOREIGN sky130_fd_sc_hdll__tap ;
  ORIGIN  14.88000  15.82500 ;
  SIZE  2093.810 BY  34.45000 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 177.780000 4.880000 180.095000 5.595000 ;
        RECT 177.780000 5.895000 180.095000 6.610000 ;
        RECT 177.980000 5.595000 180.095000 5.895000 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 177.780000 1.550000 180.095000 2.265000 ;
        RECT 177.780000 2.565000 180.095000 3.280000 ;
        RECT 177.980000 2.265000 180.095000 2.565000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT    0.000000 -0.085000 2064.020000 0.085000 ;
      RECT    0.000000  2.635000 1944.615000 2.805000 ;
      RECT    0.000000  5.355000  234.600000 5.525000 ;
      RECT    0.090000  0.265000    0.425000 1.685000 ;
      RECT    0.090000  1.685000    0.355000 2.455000 ;
      RECT    0.095000  2.975000    0.425000 3.470000 ;
      RECT    0.095000  3.470000    2.275000 3.640000 ;
      RECT    0.095000  3.640000    0.355000 3.980000 ;
      RECT    0.095000  4.150000    0.695000 4.385000 ;
      RECT    0.205000  4.555000    0.535000 5.355000 ;
      RECT    0.525000  1.915000    0.905000 2.635000 ;
      RECT    0.525000  3.810000    1.875000 3.980000 ;
      RECT    0.525000  3.980000    0.695000 4.150000 ;
      RECT    0.595000  2.805000    0.865000 3.300000 ;
      RECT    0.605000  0.625000    3.535000 0.815000 ;
      RECT    0.605000  0.815000    0.845000 1.505000 ;
      RECT    0.605000  1.505000    3.545000 1.685000 ;
      RECT    0.655000  0.085000    1.400000 0.455000 ;
      RECT    0.865000  4.150000    1.535000 4.385000 ;
      RECT    1.015000  0.995000    1.695000 1.325000 ;
      RECT    1.035000  2.975000    1.365000 3.470000 ;
      RECT    1.035000  4.555000    3.735000 4.765000 ;
      RECT    1.035000  4.765000    1.365000 5.165000 ;
      RECT    1.095000  1.865000    2.565000 2.095000 ;
      RECT    1.095000  2.095000    1.355000 2.455000 ;
      RECT    1.525000  2.265000    2.085000 2.635000 ;
      RECT    1.535000  2.805000    1.805000 3.300000 ;
      RECT    1.705000  3.980000    1.875000 4.150000 ;
      RECT    1.705000  4.150000    2.045000 4.385000 ;
      RECT    1.865000  0.995000    2.390000 1.325000 ;
      RECT    1.945000  4.935000    2.275000 5.355000 ;
      RECT    1.975000  2.975000    3.245000 3.145000 ;
      RECT    1.975000  3.145000    2.275000 3.470000 ;
      RECT    2.045000  3.640000    2.275000 3.980000 ;
      RECT    2.195000  0.265000    2.520000 0.625000 ;
      RECT    2.305000  2.095000    2.565000 2.455000 ;
      RECT    2.445000  3.315000    2.745000 3.650000 ;
      RECT    2.445000  3.650000    2.695000 4.555000 ;
      RECT    2.445000  4.765000    2.745000 5.185000 ;
      RECT    2.590000  0.995000    3.075000 1.325000 ;
      RECT    2.700000  0.085000    3.080000 0.455000 ;
      RECT    2.865000  3.825000    3.195000 4.385000 ;
      RECT    2.915000  3.145000    3.245000 3.655000 ;
      RECT    2.915000  4.935000    3.735000 5.355000 ;
      RECT    3.205000  1.685000    3.545000 2.455000 ;
      RECT    3.305000  0.995000    3.585000 1.325000 ;
      RECT    3.310000  0.265000    3.535000 0.625000 ;
      RECT    3.485000  2.805000    3.735000 3.945000 ;
      RECT    3.565000  4.165000    5.455000 4.405000 ;
      RECT    3.565000  4.405000    3.735000 4.555000 ;
      RECT    3.765000  0.085000    4.055000 0.810000 ;
      RECT    3.765000  1.470000    4.055000 2.635000 ;
      RECT    3.905000  4.575000    6.115000 4.745000 ;
      RECT    3.905000  4.745000    4.235000 5.185000 ;
      RECT    3.935000  2.975000    4.205000 3.825000 ;
      RECT    3.935000  3.825000    6.085000 3.995000 ;
      RECT    4.230000  0.085000    4.525000 0.905000 ;
      RECT    4.230000  1.490000    4.525000 2.635000 ;
      RECT    4.375000  2.805000    4.705000 3.655000 ;
      RECT    4.405000  4.915000    4.675000 5.355000 ;
      RECT    4.745000  0.255000    4.975000 2.335000 ;
      RECT    4.845000  4.745000    5.175000 5.185000 ;
      RECT    4.875000  2.975000    5.145000 3.825000 ;
      RECT    5.145000  0.085000    5.910000 0.445000 ;
      RECT    5.240000  0.695000    8.075000 0.875000 ;
      RECT    5.240000  0.875000    5.495000 1.490000 ;
      RECT    5.240000  1.490000    8.075000 1.660000 ;
      RECT    5.240000  1.830000    5.495000 2.635000 ;
      RECT    5.315000  2.805000    5.645000 3.655000 ;
      RECT    5.345000  4.915000    5.615000 5.355000 ;
      RECT    5.625000  3.995000    5.875000 4.575000 ;
      RECT    5.665000  1.045000    6.100000 1.275000 ;
      RECT    5.695000  1.840000    7.185000 2.020000 ;
      RECT    5.695000  2.020000    6.075000 2.465000 ;
      RECT    5.785000  4.745000    6.115000 5.185000 ;
      RECT    5.815000  2.975000    6.085000 3.825000 ;
      RECT    6.265000  2.805000    6.595000 3.995000 ;
      RECT    6.285000  4.535000    6.535000 5.355000 ;
      RECT    6.295000  2.190000    6.570000 2.635000 ;
      RECT    6.430000  1.045000    6.835000 1.275000 ;
      RECT    6.615000  0.275000    6.995000 0.695000 ;
      RECT    6.855000  2.020000    7.185000 2.465000 ;
      RECT    6.985000  2.805000    7.275000 3.970000 ;
      RECT    6.985000  4.630000    7.275000 5.355000 ;
      RECT    7.005000  1.045000    7.335000 1.275000 ;
      RECT    7.250000  0.085000    7.525000 0.525000 ;
      RECT    7.455000  2.975000    7.785000 3.470000 ;
      RECT    7.455000  3.470000    9.635000 3.640000 ;
      RECT    7.455000  3.640000    7.715000 3.980000 ;
      RECT    7.455000  4.150000    8.055000 4.385000 ;
      RECT    7.505000  1.045000    7.875000 1.275000 ;
      RECT    7.565000  4.555000    7.895000 5.355000 ;
      RECT    7.695000  0.275000    8.075000 0.695000 ;
      RECT    7.695000  1.660000    8.075000 2.325000 ;
      RECT    7.885000  3.810000    9.235000 3.980000 ;
      RECT    7.885000  3.980000    8.055000 4.150000 ;
      RECT    7.955000  2.805000    8.225000 3.300000 ;
      RECT    8.225000  4.150000    8.895000 4.385000 ;
      RECT    8.365000  0.085000    8.655000 0.810000 ;
      RECT    8.365000  1.470000    8.655000 2.635000 ;
      RECT    8.395000  2.975000    8.725000 3.470000 ;
      RECT    8.395000  4.555000   11.095000 4.765000 ;
      RECT    8.395000  4.765000    8.725000 5.165000 ;
      RECT    8.825000  0.635000   10.965000 0.875000 ;
      RECT    8.825000  0.875000    9.080000 1.495000 ;
      RECT    8.825000  1.495000   10.530000 1.705000 ;
      RECT    8.830000  1.875000    9.165000 2.635000 ;
      RECT    8.895000  2.805000    9.165000 3.300000 ;
      RECT    9.065000  3.980000    9.235000 4.150000 ;
      RECT    9.065000  4.150000    9.405000 4.385000 ;
      RECT    9.225000  0.085000    9.605000 0.465000 ;
      RECT    9.265000  1.045000   11.360000 1.325000 ;
      RECT    9.305000  4.935000    9.635000 5.355000 ;
      RECT    9.335000  2.975000   10.605000 3.145000 ;
      RECT    9.335000  3.145000    9.635000 3.470000 ;
      RECT    9.385000  1.705000    9.570000 2.465000 ;
      RECT    9.405000  3.640000    9.635000 3.980000 ;
      RECT    9.790000  1.875000   10.120000 2.635000 ;
      RECT    9.805000  3.315000   10.105000 3.650000 ;
      RECT    9.805000  3.650000   10.055000 4.555000 ;
      RECT    9.805000  4.765000   10.105000 5.185000 ;
      RECT    9.825000  0.255000   10.015000 0.615000 ;
      RECT    9.825000  0.615000   10.965000 0.635000 ;
      RECT   10.185000  0.085000   10.565000 0.445000 ;
      RECT   10.225000  3.825000   10.555000 4.385000 ;
      RECT   10.275000  3.145000   10.605000 3.655000 ;
      RECT   10.275000  4.935000   11.095000 5.355000 ;
      RECT   10.340000  1.705000   10.530000 2.465000 ;
      RECT   10.750000  1.835000   11.000000 2.635000 ;
      RECT   10.785000  0.255000   10.965000 0.615000 ;
      RECT   10.845000  2.805000   11.095000 3.945000 ;
      RECT   10.925000  4.165000   13.495000 4.405000 ;
      RECT   10.925000  4.405000   11.095000 4.555000 ;
      RECT   11.125000  1.325000   11.360000 1.505000 ;
      RECT   11.125000  1.505000   11.445000 1.675000 ;
      RECT   11.135000  0.615000   14.780000 0.805000 ;
      RECT   11.135000  0.805000   11.360000 1.045000 ;
      RECT   11.160000  0.085000   11.545000 0.445000 ;
      RECT   11.265000  4.575000   14.415000 4.745000 ;
      RECT   11.265000  4.745000   11.595000 5.185000 ;
      RECT   11.270000  1.675000   11.445000 1.870000 ;
      RECT   11.270000  1.870000   12.600000 2.040000 ;
      RECT   11.295000  2.975000   11.565000 3.825000 ;
      RECT   11.295000  3.825000   14.385000 3.995000 ;
      RECT   11.310000  2.210000   13.640000 2.465000 ;
      RECT   11.530000  0.985000   11.845000 1.325000 ;
      RECT   11.615000  1.325000   11.845000 1.445000 ;
      RECT   11.615000  1.445000   13.365000 1.700000 ;
      RECT   11.735000  2.805000   12.065000 3.655000 ;
      RECT   11.765000  0.255000   12.010000 0.615000 ;
      RECT   11.765000  4.915000   12.035000 5.355000 ;
      RECT   12.015000  0.985000   12.785000 1.275000 ;
      RECT   12.180000  0.085000   12.560000 0.445000 ;
      RECT   12.205000  4.745000   12.535000 5.185000 ;
      RECT   12.235000  2.975000   12.505000 3.825000 ;
      RECT   12.675000  2.805000   13.005000 3.655000 ;
      RECT   12.705000  4.915000   12.975000 5.355000 ;
      RECT   12.780000  0.255000   13.160000 0.615000 ;
      RECT   12.985000  0.985000   13.365000 1.445000 ;
      RECT   13.145000  4.745000   13.475000 5.185000 ;
      RECT   13.175000  2.975000   13.445000 3.825000 ;
      RECT   13.310000  1.880000   15.735000 2.105000 ;
      RECT   13.310000  2.105000   13.640000 2.210000 ;
      RECT   13.380000  0.085000   13.750000 0.445000 ;
      RECT   13.615000  2.805000   13.945000 3.655000 ;
      RECT   13.645000  4.915000   13.915000 5.355000 ;
      RECT   13.685000  1.020000   14.065000 1.510000 ;
      RECT   13.685000  1.510000   15.185000 1.700000 ;
      RECT   13.810000  2.275000   14.190000 2.635000 ;
      RECT   13.905000  3.995000   14.155000 4.575000 ;
      RECT   14.085000  4.745000   14.415000 5.185000 ;
      RECT   14.115000  2.975000   14.385000 3.825000 ;
      RECT   14.275000  1.020000   14.670000 1.330000 ;
      RECT   14.400000  0.275000   14.780000 0.615000 ;
      RECT   14.400000  2.105000   14.710000 2.465000 ;
      RECT   14.575000  2.805000   14.885000 3.995000 ;
      RECT   14.585000  4.535000   14.835000 5.355000 ;
      RECT   14.865000  1.020000   15.615000 1.320000 ;
      RECT   14.865000  1.320000   15.185000 1.510000 ;
      RECT   14.880000  2.275000   15.260000 2.635000 ;
      RECT   15.265000  2.805000   15.555000 3.970000 ;
      RECT   15.265000  4.630000   15.555000 5.355000 ;
      RECT   15.355000  0.085000   15.735000 0.805000 ;
      RECT   15.355000  1.535000   15.735000 1.880000 ;
      RECT   15.480000  2.105000   15.735000 2.465000 ;
      RECT   15.725000  4.115000   16.255000 4.445000 ;
      RECT   15.735000  2.805000   16.035000 3.635000 ;
      RECT   15.735000  4.615000   16.065000 5.355000 ;
      RECT   16.075000  3.805000   17.525000 3.975000 ;
      RECT   16.075000  3.975000   16.255000 4.115000 ;
      RECT   16.185000  0.085000   16.475000 0.810000 ;
      RECT   16.185000  1.470000   16.475000 2.635000 ;
      RECT   16.205000  2.975000   16.505000 3.465000 ;
      RECT   16.205000  3.465000   17.945000 3.635000 ;
      RECT   16.505000  4.145000   17.175000 4.445000 ;
      RECT   16.645000  0.085000   16.985000 0.595000 ;
      RECT   16.655000  0.765000   16.995000 1.325000 ;
      RECT   16.655000  4.615000   17.945000 4.785000 ;
      RECT   16.655000  4.785000   16.985000 5.185000 ;
      RECT   16.675000  2.805000   17.005000 3.295000 ;
      RECT   16.685000  1.525000   17.890000 1.725000 ;
      RECT   16.685000  1.725000   16.935000 2.455000 ;
      RECT   17.105000  1.905000   17.485000 2.635000 ;
      RECT   17.165000  0.265000   17.465000 0.995000 ;
      RECT   17.165000  0.995000   17.840000 1.325000 ;
      RECT   17.175000  2.975000   17.445000 3.465000 ;
      RECT   17.345000  3.975000   17.525000 4.115000 ;
      RECT   17.345000  4.115000   17.605000 4.445000 ;
      RECT   17.580000  4.955000   17.910000 5.355000 ;
      RECT   17.615000  2.805000   17.945000 3.280000 ;
      RECT   17.705000  1.725000   17.890000 2.455000 ;
      RECT   17.715000  0.265000   17.900000 0.625000 ;
      RECT   17.715000  0.625000   19.210000 0.815000 ;
      RECT   17.775000  3.635000   17.945000 4.175000 ;
      RECT   17.775000  4.175000   19.945000 4.385000 ;
      RECT   17.775000  4.385000   17.945000 4.615000 ;
      RECT   18.060000  0.995000   18.355000 2.455000 ;
      RECT   18.110000  0.085000   18.490000 0.455000 ;
      RECT   18.115000  2.975000   18.385000 3.825000 ;
      RECT   18.115000  3.825000   20.615000 3.995000 ;
      RECT   18.115000  4.555000   20.615000 4.725000 ;
      RECT   18.115000  4.725000   18.385000 5.185000 ;
      RECT   18.525000  1.785000   19.210000 2.455000 ;
      RECT   18.540000  0.995000   18.825000 1.615000 ;
      RECT   18.555000  2.805000   18.885000 3.655000 ;
      RECT   18.555000  4.895000   18.885000 5.355000 ;
      RECT   18.815000  0.265000   19.040000 0.625000 ;
      RECT   18.995000  0.815000   19.210000 1.785000 ;
      RECT   19.055000  2.975000   19.325000 3.825000 ;
      RECT   19.055000  4.725000   19.325000 5.185000 ;
      RECT   19.405000  0.085000   19.695000 0.810000 ;
      RECT   19.405000  1.470000   19.695000 2.635000 ;
      RECT   19.495000  2.805000   19.825000 3.655000 ;
      RECT   19.495000  4.895000   19.825000 5.355000 ;
      RECT   19.880000  0.995000   20.185000 1.615000 ;
      RECT   19.925000  0.085000   20.175000 0.815000 ;
      RECT   19.925000  1.785000   20.185000 2.285000 ;
      RECT   19.925000  2.285000   22.195000 2.455000 ;
      RECT   19.995000  2.975000   20.265000 3.825000 ;
      RECT   19.995000  4.725000   20.265000 5.185000 ;
      RECT   20.115000  3.995000   20.615000 4.555000 ;
      RECT   20.355000  0.255000   20.665000 0.655000 ;
      RECT   20.355000  0.655000   23.175000 0.855000 ;
      RECT   20.355000  0.855000   20.675000 2.115000 ;
      RECT   20.435000  2.805000   20.765000 3.655000 ;
      RECT   20.435000  4.895000   20.765000 5.355000 ;
      RECT   20.835000  0.085000   21.215000 0.475000 ;
      RECT   20.845000  1.035000   21.715000 1.285000 ;
      RECT   20.845000  1.285000   21.065000 1.615000 ;
      RECT   20.955000  1.785000   21.145000 2.255000 ;
      RECT   20.955000  2.255000   22.195000 2.285000 ;
      RECT   21.245000  2.805000   21.535000 3.970000 ;
      RECT   21.245000  4.630000   21.535000 5.355000 ;
      RECT   21.315000  1.455000   24.105000 1.655000 ;
      RECT   21.315000  1.655000   21.695000 2.075000 ;
      RECT   21.705000  4.115000   22.235000 4.445000 ;
      RECT   21.715000  2.805000   22.015000 3.635000 ;
      RECT   21.715000  4.615000   22.045000 5.355000 ;
      RECT   21.795000  0.085000   22.175000 0.475000 ;
      RECT   21.915000  1.835000   22.195000 2.255000 ;
      RECT   22.055000  3.805000   23.505000 3.975000 ;
      RECT   22.055000  3.975000   22.235000 4.115000 ;
      RECT   22.185000  2.975000   22.485000 3.465000 ;
      RECT   22.185000  3.465000   23.925000 3.635000 ;
      RECT   22.365000  0.265000   23.575000 0.475000 ;
      RECT   22.415000  1.835000   22.645000 2.635000 ;
      RECT   22.485000  4.145000   23.155000 4.445000 ;
      RECT   22.590000  1.035000   23.350000 1.285000 ;
      RECT   22.635000  4.615000   23.925000 4.785000 ;
      RECT   22.635000  4.785000   22.965000 5.185000 ;
      RECT   22.655000  2.805000   22.985000 3.295000 ;
      RECT   22.875000  1.655000   23.145000 2.465000 ;
      RECT   23.155000  2.975000   23.425000 3.465000 ;
      RECT   23.325000  3.975000   23.505000 4.115000 ;
      RECT   23.325000  4.115000   23.585000 4.445000 ;
      RECT   23.375000  1.835000   23.605000 2.635000 ;
      RECT   23.405000  0.475000   23.575000 0.635000 ;
      RECT   23.405000  0.635000   24.615000 0.855000 ;
      RECT   23.560000  4.955000   23.890000 5.355000 ;
      RECT   23.595000  2.805000   23.925000 3.280000 ;
      RECT   23.670000  1.035000   24.695000 1.285000 ;
      RECT   23.755000  0.085000   24.135000 0.455000 ;
      RECT   23.755000  3.635000   23.925000 4.175000 ;
      RECT   23.755000  4.175000   26.945000 4.385000 ;
      RECT   23.755000  4.385000   23.925000 4.615000 ;
      RECT   23.835000  1.655000   24.105000 2.465000 ;
      RECT   24.095000  2.975000   24.365000 3.825000 ;
      RECT   24.095000  3.825000   27.535000 3.995000 ;
      RECT   24.095000  4.555000   27.535000 4.725000 ;
      RECT   24.095000  4.725000   24.365000 5.185000 ;
      RECT   24.335000  1.835000   24.565000 2.635000 ;
      RECT   24.365000  0.265000   24.615000 0.635000 ;
      RECT   24.465000  1.285000   24.695000 1.655000 ;
      RECT   24.535000  2.805000   24.865000 3.655000 ;
      RECT   24.535000  4.895000   24.865000 5.355000 ;
      RECT   24.925000  0.085000   25.215000 0.810000 ;
      RECT   24.925000  1.470000   25.215000 2.635000 ;
      RECT   25.035000  2.975000   25.305000 3.825000 ;
      RECT   25.035000  4.725000   25.305000 5.185000 ;
      RECT   25.395000  0.085000   25.695000 0.585000 ;
      RECT   25.395000  1.795000   29.405000 2.085000 ;
      RECT   25.395000  2.085000   25.645000 2.465000 ;
      RECT   25.400000  1.035000   26.835000 1.445000 ;
      RECT   25.400000  1.445000   29.275000 1.625000 ;
      RECT   25.475000  2.805000   25.805000 3.655000 ;
      RECT   25.475000  4.895000   25.805000 5.355000 ;
      RECT   25.815000  2.255000   26.195000 2.635000 ;
      RECT   25.915000  0.530000   26.125000 0.695000 ;
      RECT   25.915000  0.695000   27.055000 0.865000 ;
      RECT   25.975000  2.975000   26.245000 3.825000 ;
      RECT   25.975000  4.725000   26.245000 5.185000 ;
      RECT   26.300000  0.085000   26.585000 0.525000 ;
      RECT   26.415000  2.085000   29.405000 2.105000 ;
      RECT   26.415000  2.105000   26.585000 2.465000 ;
      RECT   26.415000  2.805000   26.745000 3.655000 ;
      RECT   26.415000  4.895000   26.745000 5.355000 ;
      RECT   26.755000  0.255000   29.015000 0.505000 ;
      RECT   26.755000  0.505000   27.055000 0.695000 ;
      RECT   26.755000  2.275000   27.135000 2.635000 ;
      RECT   26.915000  2.975000   27.185000 3.825000 ;
      RECT   26.915000  4.725000   27.185000 5.185000 ;
      RECT   27.105000  1.035000   28.605000 1.275000 ;
      RECT   27.115000  3.995000   27.535000 4.555000 ;
      RECT   27.225000  0.675000   28.980000 0.695000 ;
      RECT   27.225000  0.695000   33.460000 0.825000 ;
      RECT   27.225000  0.825000   32.355000 0.865000 ;
      RECT   27.355000  2.105000   27.525000 2.465000 ;
      RECT   27.355000  2.805000   27.685000 3.655000 ;
      RECT   27.355000  4.895000   27.685000 5.355000 ;
      RECT   27.695000  2.275000   28.075000 2.635000 ;
      RECT   28.145000  2.805000   28.435000 3.970000 ;
      RECT   28.145000  4.630000   28.435000 5.355000 ;
      RECT   28.295000  2.105000   28.465000 2.465000 ;
      RECT   28.605000  4.115000   28.915000 4.725000 ;
      RECT   28.615000  2.805000   28.915000 3.945000 ;
      RECT   28.635000  2.275000   29.015000 2.635000 ;
      RECT   28.665000  4.895000   28.915000 5.355000 ;
      RECT   28.895000  1.035000   29.275000 1.445000 ;
      RECT   29.085000  2.975000   29.415000 4.115000 ;
      RECT   29.085000  4.115000   31.910000 4.365000 ;
      RECT   29.085000  4.365000   29.415000 5.175000 ;
      RECT   29.235000  0.085000   29.405000 0.525000 ;
      RECT   29.235000  2.105000   29.405000 2.255000 ;
      RECT   29.235000  2.255000   33.370000 2.465000 ;
      RECT   29.445000  1.035000   30.605000 1.275000 ;
      RECT   29.445000  1.275000   30.260000 1.615000 ;
      RECT   29.575000  0.255000   29.945000 0.615000 ;
      RECT   29.575000  0.615000   30.895000 0.625000 ;
      RECT   29.575000  0.625000   33.460000 0.695000 ;
      RECT   29.575000  1.785000   30.760000 2.085000 ;
      RECT   29.585000  2.805000   29.855000 3.945000 ;
      RECT   29.585000  4.830000   29.855000 5.355000 ;
      RECT   30.025000  2.980000   30.355000 3.775000 ;
      RECT   30.025000  3.775000   32.595000 3.945000 ;
      RECT   30.025000  4.535000   32.595000 4.705000 ;
      RECT   30.025000  4.705000   30.355000 5.185000 ;
      RECT   30.165000  0.085000   30.495000 0.445000 ;
      RECT   30.430000  1.445000   31.910000 1.695000 ;
      RECT   30.430000  1.695000   30.760000 1.785000 ;
      RECT   30.525000  2.805000   30.795000 3.605000 ;
      RECT   30.525000  4.875000   30.795000 5.355000 ;
      RECT   30.725000  0.255000   30.895000 0.615000 ;
      RECT   30.850000  1.035000   32.350000 1.275000 ;
      RECT   30.965000  2.980000   31.295000 3.775000 ;
      RECT   30.965000  4.705000   31.295000 5.185000 ;
      RECT   31.020000  1.865000   33.460000 2.085000 ;
      RECT   31.115000  0.085000   31.445000 0.445000 ;
      RECT   31.465000  2.805000   31.735000 3.605000 ;
      RECT   31.465000  4.875000   31.735000 5.355000 ;
      RECT   31.665000  0.255000   31.835000 0.615000 ;
      RECT   31.665000  0.615000   33.460000 0.625000 ;
      RECT   31.905000  2.980000   32.235000 3.775000 ;
      RECT   31.905000  4.705000   32.235000 5.185000 ;
      RECT   32.055000  0.085000   32.385000 0.445000 ;
      RECT   32.130000  1.275000   32.350000 1.695000 ;
      RECT   32.265000  3.945000   32.595000 4.535000 ;
      RECT   32.405000  2.805000   32.675000 3.605000 ;
      RECT   32.405000  4.875000   32.675000 5.355000 ;
      RECT   32.600000  0.995000   33.035000 1.325000 ;
      RECT   32.600000  1.325000   32.810000 1.655000 ;
      RECT   32.965000  0.085000   33.370000 0.445000 ;
      RECT   32.980000  1.495000   33.460000 1.865000 ;
      RECT   33.205000  0.825000   33.460000 1.495000 ;
      RECT   33.205000  2.805000   33.495000 3.970000 ;
      RECT   33.205000  4.630000   33.495000 5.355000 ;
      RECT   33.665000  0.085000   33.955000 0.810000 ;
      RECT   33.665000  1.470000   33.955000 2.635000 ;
      RECT   33.675000  2.805000   33.975000 3.945000 ;
      RECT   33.675000  4.830000   34.005000 5.355000 ;
      RECT   34.105000  4.135000   34.900000 4.365000 ;
      RECT   34.145000  0.325000   34.375000 1.665000 ;
      RECT   34.145000  1.845000   35.005000 2.045000 ;
      RECT   34.145000  2.045000   34.385000 2.435000 ;
      RECT   34.145000  2.975000   34.475000 3.775000 ;
      RECT   34.145000  3.775000   35.385000 3.945000 ;
      RECT   34.150000  3.945000   35.385000 3.965000 ;
      RECT   34.175000  4.535000   35.385000 4.725000 ;
      RECT   34.175000  4.725000   34.445000 5.160000 ;
      RECT   34.555000  0.265000   34.835000 1.165000 ;
      RECT   34.555000  1.165000   35.005000 1.845000 ;
      RECT   34.555000  2.225000   34.955000 2.635000 ;
      RECT   34.615000  4.895000   34.945000 5.355000 ;
      RECT   34.645000  2.805000   34.915000 3.605000 ;
      RECT   35.085000  0.085000   35.330000 0.865000 ;
      RECT   35.115000  2.975000   35.385000 3.775000 ;
      RECT   35.115000  3.965000   35.385000 4.135000 ;
      RECT   35.115000  4.135000   40.265000 4.365000 ;
      RECT   35.115000  4.365000   35.385000 4.535000 ;
      RECT   35.115000  4.725000   35.385000 5.160000 ;
      RECT   35.175000  1.045000   35.770000 1.345000 ;
      RECT   35.175000  1.345000   35.505000 2.455000 ;
      RECT   35.500000  0.265000   35.980000 0.625000 ;
      RECT   35.500000  0.625000   37.585000 0.815000 ;
      RECT   35.500000  0.815000   35.770000 1.045000 ;
      RECT   35.555000  2.805000   35.855000 3.965000 ;
      RECT   35.555000  4.895000   35.885000 5.355000 ;
      RECT   35.725000  1.785000   36.850000 1.985000 ;
      RECT   35.725000  1.985000   35.905000 2.455000 ;
      RECT   35.940000  0.995000   36.315000 1.615000 ;
      RECT   36.025000  2.975000   36.325000 3.775000 ;
      RECT   36.025000  3.775000   41.025000 3.965000 ;
      RECT   36.055000  4.535000   41.025000 4.725000 ;
      RECT   36.055000  4.725000   36.325000 5.160000 ;
      RECT   36.075000  2.155000   36.455000 2.635000 ;
      RECT   36.485000  0.995000   36.745000 1.615000 ;
      RECT   36.495000  2.805000   36.825000 3.605000 ;
      RECT   36.495000  4.895000   36.825000 5.355000 ;
      RECT   36.660000  0.085000   37.390000 0.455000 ;
      RECT   36.680000  1.985000   36.850000 2.455000 ;
      RECT   36.995000  2.975000   37.265000 3.775000 ;
      RECT   36.995000  4.725000   37.265000 5.160000 ;
      RECT   37.115000  1.495000   37.400000 2.635000 ;
      RECT   37.325000  0.815000   37.585000 1.325000 ;
      RECT   37.435000  2.805000   37.765000 3.605000 ;
      RECT   37.435000  4.895000   37.765000 5.355000 ;
      RECT   37.755000  0.265000   38.035000 2.455000 ;
      RECT   37.935000  2.975000   38.205000 3.775000 ;
      RECT   37.935000  4.725000   38.205000 5.160000 ;
      RECT   38.265000  0.085000   38.555000 0.810000 ;
      RECT   38.265000  1.470000   38.555000 2.635000 ;
      RECT   38.375000  2.805000   38.705000 3.605000 ;
      RECT   38.375000  4.895000   38.705000 5.355000 ;
      RECT   38.730000  0.085000   38.985000 0.545000 ;
      RECT   38.730000  2.255000   39.065000 2.635000 ;
      RECT   38.750000  0.715000   39.540000 0.885000 ;
      RECT   38.750000  0.885000   39.020000 1.835000 ;
      RECT   38.750000  1.835000   39.540000 2.005000 ;
      RECT   38.875000  2.975000   39.145000 3.775000 ;
      RECT   38.875000  4.725000   39.145000 5.160000 ;
      RECT   39.160000  0.315000   39.540000 0.715000 ;
      RECT   39.260000  1.075000   39.590000 1.495000 ;
      RECT   39.260000  1.495000   40.025000 1.665000 ;
      RECT   39.285000  2.005000   39.540000 2.425000 ;
      RECT   39.315000  2.805000   39.645000 3.605000 ;
      RECT   39.315000  4.895000   39.645000 5.355000 ;
      RECT   39.710000  0.085000   40.040000 0.785000 ;
      RECT   39.780000  2.275000   40.110000 2.635000 ;
      RECT   39.815000  2.975000   40.085000 3.775000 ;
      RECT   39.815000  4.725000   40.085000 5.160000 ;
      RECT   39.855000  1.665000   40.025000 1.895000 ;
      RECT   39.855000  1.895000   41.015000 2.105000 ;
      RECT   39.865000  0.995000   40.335000 1.325000 ;
      RECT   40.195000  1.555000   40.675000 1.725000 ;
      RECT   40.245000  0.655000   40.675000 0.825000 ;
      RECT   40.255000  2.805000   40.585000 3.605000 ;
      RECT   40.255000  4.895000   40.585000 5.355000 ;
      RECT   40.505000  0.825000   40.675000 0.995000 ;
      RECT   40.505000  0.995000   40.965000 1.325000 ;
      RECT   40.505000  1.325000   40.675000 1.555000 ;
      RECT   40.540000  3.965000   41.025000 4.535000 ;
      RECT   40.755000  2.975000   41.025000 3.775000 ;
      RECT   40.755000  4.725000   41.025000 5.160000 ;
      RECT   40.765000  0.085000   41.095000 0.465000 ;
      RECT   40.765000  2.105000   41.015000 2.465000 ;
      RECT   40.845000  1.505000   41.355000 1.675000 ;
      RECT   40.845000  1.675000   41.015000 1.895000 ;
      RECT   41.135000  0.635000   41.580000 0.825000 ;
      RECT   41.135000  0.825000   41.355000 1.505000 ;
      RECT   41.185000  1.845000   42.515000 2.015000 ;
      RECT   41.185000  2.015000   41.565000 2.465000 ;
      RECT   41.195000  2.805000   41.525000 3.975000 ;
      RECT   41.195000  4.830000   41.525000 5.355000 ;
      RECT   41.525000  0.995000   41.725000 1.615000 ;
      RECT   41.795000  2.185000   41.965000 2.635000 ;
      RECT   41.945000  2.805000   42.235000 3.970000 ;
      RECT   41.945000  4.630000   42.235000 5.355000 ;
      RECT   42.015000  0.995000   42.305000 1.615000 ;
      RECT   42.135000  0.085000   42.515000 0.825000 ;
      RECT   42.135000  2.015000   42.515000 2.465000 ;
      RECT   42.415000  2.805000   42.745000 3.640000 ;
      RECT   42.435000  3.810000   50.975000 3.980000 ;
      RECT   42.435000  3.980000   42.605000 4.575000 ;
      RECT   42.435000  4.575000   50.975000 4.745000 ;
      RECT   42.775000  4.150000   50.245000 4.405000 ;
      RECT   42.865000  0.085000   43.155000 0.810000 ;
      RECT   42.865000  1.470000   43.155000 2.635000 ;
      RECT   42.915000  2.975000   43.185000 3.810000 ;
      RECT   43.345000  0.255000   43.750000 0.840000 ;
      RECT   43.345000  0.840000   43.540000 1.795000 ;
      RECT   43.345000  1.795000   43.775000 1.935000 ;
      RECT   43.345000  1.935000   46.330000 2.105000 ;
      RECT   43.345000  2.105000   43.760000 2.465000 ;
      RECT   43.355000  2.805000   43.685000 3.640000 ;
      RECT   43.485000  4.915000   44.155000 5.355000 ;
      RECT   43.710000  1.010000   44.090000 1.625000 ;
      RECT   43.855000  2.975000   44.125000 3.810000 ;
      RECT   43.920000  0.085000   44.310000 0.445000 ;
      RECT   43.930000  2.275000   44.310000 2.635000 ;
      RECT   44.290000  0.615000   45.750000 0.785000 ;
      RECT   44.290000  0.785000   44.780000 1.595000 ;
      RECT   44.290000  1.595000   45.820000 1.765000 ;
      RECT   44.295000  2.805000   44.625000 3.640000 ;
      RECT   44.325000  4.745000   44.595000 5.185000 ;
      RECT   44.765000  4.915000   45.095000 5.355000 ;
      RECT   44.795000  2.975000   45.065000 3.810000 ;
      RECT   44.890000  0.085000   45.270000 0.445000 ;
      RECT   44.890000  2.275000   45.270000 2.635000 ;
      RECT   44.950000  0.995000   46.270000 1.185000 ;
      RECT   44.950000  1.185000   45.990000 1.325000 ;
      RECT   45.235000  2.805000   45.565000 3.640000 ;
      RECT   45.265000  4.745000   45.535000 5.185000 ;
      RECT   45.705000  4.915000   46.035000 5.355000 ;
      RECT   45.735000  2.975000   46.005000 3.810000 ;
      RECT   45.845000  2.275000   46.230000 2.635000 ;
      RECT   45.975000  0.085000   46.745000 0.445000 ;
      RECT   46.100000  0.615000   47.155000 0.670000 ;
      RECT   46.100000  0.670000   48.625000 0.785000 ;
      RECT   46.100000  0.785000   46.270000 0.995000 ;
      RECT   46.160000  1.355000   46.765000 1.525000 ;
      RECT   46.160000  1.525000   46.330000 1.935000 ;
      RECT   46.175000  2.805000   46.505000 3.640000 ;
      RECT   46.205000  4.745000   46.475000 5.185000 ;
      RECT   46.455000  0.995000   46.765000 1.355000 ;
      RECT   46.515000  1.695000   46.685000 2.210000 ;
      RECT   46.515000  2.210000   47.625000 2.380000 ;
      RECT   46.645000  4.915000   46.975000 5.355000 ;
      RECT   46.675000  2.975000   46.945000 3.810000 ;
      RECT   46.985000  0.255000   47.155000 0.615000 ;
      RECT   46.985000  0.785000   48.625000 0.840000 ;
      RECT   46.985000  0.840000   47.155000 1.805000 ;
      RECT   47.115000  2.805000   47.445000 3.640000 ;
      RECT   47.145000  4.745000   47.415000 5.185000 ;
      RECT   47.415000  0.085000   47.745000 0.445000 ;
      RECT   47.445000  1.445000   47.625000 1.935000 ;
      RECT   47.445000  1.935000   49.585000 2.105000 ;
      RECT   47.445000  2.105000   47.625000 2.210000 ;
      RECT   47.585000  1.010000   48.030000 1.275000 ;
      RECT   47.585000  4.915000   47.915000 5.355000 ;
      RECT   47.615000  2.975000   47.885000 3.810000 ;
      RECT   47.795000  2.275000   48.175000 2.635000 ;
      RECT   47.805000  1.275000   48.030000 1.595000 ;
      RECT   47.805000  1.595000   49.100000 1.765000 ;
      RECT   48.055000  2.805000   48.385000 3.640000 ;
      RECT   48.085000  4.745000   48.355000 5.185000 ;
      RECT   48.200000  1.010000   48.615000 1.360000 ;
      RECT   48.345000  0.405000   48.625000 0.670000 ;
      RECT   48.525000  4.915000   48.855000 5.355000 ;
      RECT   48.555000  2.975000   48.825000 3.810000 ;
      RECT   48.735000  2.275000   49.115000 2.635000 ;
      RECT   48.870000  1.055000   49.460000 1.290000 ;
      RECT   48.870000  1.290000   49.100000 1.595000 ;
      RECT   48.995000  2.805000   49.325000 3.640000 ;
      RECT   49.025000  4.745000   49.295000 5.185000 ;
      RECT   49.305000  0.085000   49.585000 0.885000 ;
      RECT   49.330000  1.460000   49.585000 1.935000 ;
      RECT   49.465000  4.915000   50.135000 5.355000 ;
      RECT   49.495000  2.975000   49.765000 3.810000 ;
      RECT   49.765000  0.085000   50.055000 0.810000 ;
      RECT   49.765000  1.470000   50.055000 2.635000 ;
      RECT   49.935000  2.805000   50.265000 3.640000 ;
      RECT   50.235000  1.835000   50.995000 2.005000 ;
      RECT   50.235000  2.005000   50.495000 2.435000 ;
      RECT   50.245000  0.975000   50.475000 1.665000 ;
      RECT   50.420000  3.980000   50.975000 4.575000 ;
      RECT   50.435000  2.975000   50.705000 3.810000 ;
      RECT   50.505000  0.265000   50.995000 0.715000 ;
      RECT   50.655000  0.715000   50.995000 1.835000 ;
      RECT   50.665000  2.175000   51.035000 2.635000 ;
      RECT   50.875000  2.805000   51.205000 3.640000 ;
      RECT   51.165000  0.085000   51.395000 0.865000 ;
      RECT   51.205000  1.045000   51.920000 1.345000 ;
      RECT   51.205000  1.345000   51.665000 2.455000 ;
      RECT   51.580000  0.265000   51.920000 1.045000 ;
      RECT   51.605000  2.805000   51.895000 3.970000 ;
      RECT   51.605000  4.630000   51.895000 5.355000 ;
      RECT   51.885000  1.525000   53.145000 1.725000 ;
      RECT   51.885000  1.725000   52.075000 2.455000 ;
      RECT   52.075000  2.975000   54.285000 3.145000 ;
      RECT   52.075000  3.145000   52.375000 5.015000 ;
      RECT   52.075000  5.015000   54.285000 5.185000 ;
      RECT   52.125000  0.375000   52.380000 1.345000 ;
      RECT   52.245000  1.905000   52.625000 2.635000 ;
      RECT   52.545000  3.315000   52.875000 3.775000 ;
      RECT   52.545000  3.775000   53.815000 3.945000 ;
      RECT   52.545000  4.115000   53.895000 4.365000 ;
      RECT   52.545000  4.535000   56.215000 4.715000 ;
      RECT   52.545000  4.715000   52.875000 4.845000 ;
      RECT   52.790000  0.995000   53.265000 1.345000 ;
      RECT   52.855000  0.085000   53.215000 0.815000 ;
      RECT   52.975000  1.725000   53.145000 2.455000 ;
      RECT   53.045000  3.145000   53.315000 3.605000 ;
      RECT   53.045000  4.895000   53.315000 5.015000 ;
      RECT   53.445000  0.085000   53.735000 0.810000 ;
      RECT   53.445000  1.470000   53.735000 2.635000 ;
      RECT   53.485000  3.315000   53.815000 3.775000 ;
      RECT   53.485000  4.715000   53.815000 4.845000 ;
      RECT   53.915000  2.080000   54.245000 2.635000 ;
      RECT   53.940000  0.765000   54.245000 1.805000 ;
      RECT   53.985000  3.145000   54.285000 3.945000 ;
      RECT   53.985000  4.890000   54.285000 5.015000 ;
      RECT   54.085000  0.360000   54.645000 0.530000 ;
      RECT   54.465000  0.530000   54.645000 1.070000 ;
      RECT   54.465000  1.070000   55.175000 1.285000 ;
      RECT   54.465000  1.285000   54.645000 2.265000 ;
      RECT   54.505000  2.805000   54.775000 3.945000 ;
      RECT   54.505000  4.890000   54.775000 5.355000 ;
      RECT   54.905000  0.085000   55.145000 0.885000 ;
      RECT   54.905000  4.115000   56.255000 4.365000 ;
      RECT   54.920000  1.795000   55.170000 2.285000 ;
      RECT   54.920000  2.285000   56.235000 2.465000 ;
      RECT   54.945000  2.975000   55.275000 3.775000 ;
      RECT   54.945000  3.775000   56.215000 3.945000 ;
      RECT   54.945000  4.715000   55.275000 5.185000 ;
      RECT   55.345000  0.255000   55.690000 0.615000 ;
      RECT   55.345000  0.615000   57.180000 0.785000 ;
      RECT   55.345000  0.785000   55.685000 2.115000 ;
      RECT   55.445000  2.805000   55.715000 3.605000 ;
      RECT   55.445000  4.895000   55.715000 5.355000 ;
      RECT   55.855000  1.855000   58.140000 2.025000 ;
      RECT   55.855000  2.025000   56.235000 2.285000 ;
      RECT   55.885000  2.975000   56.215000 3.775000 ;
      RECT   55.885000  4.715000   56.215000 5.185000 ;
      RECT   55.960000  0.085000   56.290000 0.445000 ;
      RECT   56.115000  1.075000   56.495000 1.245000 ;
      RECT   56.120000  1.245000   56.495000 1.495000 ;
      RECT   56.120000  1.495000   57.905000 1.675000 ;
      RECT   56.385000  2.805000   56.655000 3.945000 ;
      RECT   56.385000  4.535000   56.655000 5.355000 ;
      RECT   56.455000  2.195000   56.625000 2.635000 ;
      RECT   56.675000  0.995000   57.385000 1.325000 ;
      RECT   56.800000  0.255000   57.180000 0.615000 ;
      RECT   56.825000  2.975000   57.155000 4.115000 ;
      RECT   56.825000  4.115000   59.075000 4.365000 ;
      RECT   56.825000  4.365000   57.155000 5.185000 ;
      RECT   56.930000  2.025000   58.140000 2.105000 ;
      RECT   56.930000  2.105000   57.100000 2.465000 ;
      RECT   57.280000  2.275000   57.660000 2.635000 ;
      RECT   57.325000  2.805000   57.595000 3.945000 ;
      RECT   57.325000  4.535000   57.595000 5.355000 ;
      RECT   57.555000  0.995000   57.905000 1.495000 ;
      RECT   57.765000  2.975000   58.095000 3.775000 ;
      RECT   57.765000  3.775000   59.035000 3.945000 ;
      RECT   57.765000  4.535000   61.435000 4.715000 ;
      RECT   57.765000  4.715000   58.095000 5.185000 ;
      RECT   57.810000  0.085000   58.150000 0.785000 ;
      RECT   57.880000  2.105000   58.140000 2.465000 ;
      RECT   58.265000  2.805000   58.535000 3.605000 ;
      RECT   58.265000  4.895000   58.535000 5.355000 ;
      RECT   58.505000  0.085000   58.795000 0.810000 ;
      RECT   58.505000  1.470000   58.795000 2.635000 ;
      RECT   58.705000  2.975000   59.035000 3.775000 ;
      RECT   58.705000  4.715000   59.035000 5.185000 ;
      RECT   58.970000  0.255000   59.325000 0.615000 ;
      RECT   58.970000  0.615000   60.035000 0.795000 ;
      RECT   58.975000  1.785000   59.890000 2.005000 ;
      RECT   58.975000  2.005000   59.305000 2.465000 ;
      RECT   58.995000  1.075000   59.550000 1.615000 ;
      RECT   59.205000  2.805000   59.475000 3.945000 ;
      RECT   59.205000  4.890000   59.475000 5.355000 ;
      RECT   59.330000  0.995000   59.550000 1.075000 ;
      RECT   59.525000  2.175000   59.785000 2.635000 ;
      RECT   59.650000  0.085000   60.035000 0.445000 ;
      RECT   59.695000  2.975000   61.905000 3.145000 ;
      RECT   59.695000  3.145000   59.995000 3.945000 ;
      RECT   59.695000  4.890000   59.995000 5.015000 ;
      RECT   59.695000  5.015000   61.905000 5.185000 ;
      RECT   59.720000  0.795000   60.035000 1.035000 ;
      RECT   59.720000  1.035000   61.500000 1.345000 ;
      RECT   59.720000  1.345000   59.890000 1.785000 ;
      RECT   60.060000  1.795000   60.305000 2.215000 ;
      RECT   60.060000  2.215000   62.245000 2.465000 ;
      RECT   60.085000  4.115000   61.435000 4.365000 ;
      RECT   60.165000  3.315000   60.495000 3.775000 ;
      RECT   60.165000  3.775000   61.435000 3.945000 ;
      RECT   60.165000  4.715000   60.495000 4.845000 ;
      RECT   60.255000  0.370000   60.445000 0.615000 ;
      RECT   60.255000  0.615000   61.405000 0.695000 ;
      RECT   60.255000  0.695000   64.265000 0.865000 ;
      RECT   60.560000  1.585000   62.010000 1.705000 ;
      RECT   60.560000  1.705000   61.825000 2.035000 ;
      RECT   60.665000  0.085000   61.045000 0.445000 ;
      RECT   60.665000  3.145000   60.935000 3.605000 ;
      RECT   60.665000  4.895000   60.935000 5.015000 ;
      RECT   60.935000  2.205000   62.245000 2.215000 ;
      RECT   61.105000  3.315000   61.435000 3.775000 ;
      RECT   61.105000  4.715000   61.435000 4.845000 ;
      RECT   61.215000  0.255000   61.405000 0.615000 ;
      RECT   61.605000  3.145000   61.905000 4.115000 ;
      RECT   61.605000  4.115000   66.805000 4.365000 ;
      RECT   61.605000  4.365000   61.905000 5.015000 ;
      RECT   61.625000  0.085000   62.265000 0.525000 ;
      RECT   61.700000  0.865000   64.265000 0.895000 ;
      RECT   61.700000  0.895000   62.010000 1.585000 ;
      RECT   62.045000  1.875000   66.120000 2.105000 ;
      RECT   62.045000  2.105000   62.245000 2.205000 ;
      RECT   62.125000  2.805000   62.395000 3.945000 ;
      RECT   62.125000  4.535000   62.395000 5.355000 ;
      RECT   62.180000  1.065000   62.575000 1.480000 ;
      RECT   62.180000  1.480000   66.000000 1.705000 ;
      RECT   62.415000  2.275000   62.795000 2.635000 ;
      RECT   62.435000  0.675000   64.265000 0.695000 ;
      RECT   62.445000  0.255000   64.745000 0.505000 ;
      RECT   62.565000  2.975000   62.895000 3.775000 ;
      RECT   62.565000  3.775000   67.595000 3.945000 ;
      RECT   62.565000  4.535000   67.595000 4.715000 ;
      RECT   62.565000  4.715000   62.895000 5.185000 ;
      RECT   62.745000  1.065000   64.320000 1.310000 ;
      RECT   63.065000  2.805000   63.335000 3.605000 ;
      RECT   63.065000  4.895000   63.335000 5.355000 ;
      RECT   63.375000  2.275000   63.755000 2.635000 ;
      RECT   63.505000  2.975000   63.835000 3.775000 ;
      RECT   63.505000  4.715000   63.835000 5.185000 ;
      RECT   63.975000  2.105000   64.165000 2.465000 ;
      RECT   64.005000  2.805000   64.275000 3.605000 ;
      RECT   64.005000  4.895000   64.275000 5.355000 ;
      RECT   64.335000  2.275000   64.715000 2.635000 ;
      RECT   64.445000  2.975000   64.775000 3.775000 ;
      RECT   64.445000  4.715000   64.775000 5.185000 ;
      RECT   64.485000  0.505000   64.745000 0.735000 ;
      RECT   64.485000  0.735000   65.705000 0.905000 ;
      RECT   64.605000  1.075000   66.000000 1.480000 ;
      RECT   64.930000  2.105000   65.115000 2.465000 ;
      RECT   64.945000  2.805000   65.215000 3.605000 ;
      RECT   64.945000  4.895000   65.215000 5.355000 ;
      RECT   64.965000  0.085000   65.155000 0.565000 ;
      RECT   65.295000  2.275000   65.675000 2.635000 ;
      RECT   65.325000  0.255000   65.705000 0.735000 ;
      RECT   65.385000  2.975000   65.715000 3.775000 ;
      RECT   65.385000  4.715000   65.715000 5.185000 ;
      RECT   65.870000  2.105000   66.120000 2.465000 ;
      RECT   65.880000  0.085000   66.120000 0.885000 ;
      RECT   65.885000  2.805000   66.155000 3.605000 ;
      RECT   65.885000  4.890000   66.155000 5.355000 ;
      RECT   66.325000  0.085000   66.615000 0.810000 ;
      RECT   66.325000  1.470000   66.615000 2.635000 ;
      RECT   66.325000  2.975000   66.655000 3.775000 ;
      RECT   66.325000  4.715000   66.655000 5.185000 ;
      RECT   66.795000  0.265000   67.055000 2.455000 ;
      RECT   66.825000  2.805000   67.095000 3.605000 ;
      RECT   66.825000  4.895000   67.095000 5.355000 ;
      RECT   67.225000  1.905000   67.615000 2.635000 ;
      RECT   67.245000  0.635000   68.515000 0.835000 ;
      RECT   67.245000  0.835000   67.585000 1.505000 ;
      RECT   67.245000  1.505000   68.065000 1.725000 ;
      RECT   67.265000  2.975000   67.595000 3.775000 ;
      RECT   67.265000  3.945000   67.595000 4.535000 ;
      RECT   67.265000  4.715000   67.595000 5.185000 ;
      RECT   67.365000  0.085000   68.035000 0.455000 ;
      RECT   67.765000  1.015000   68.310000 1.325000 ;
      RECT   67.765000  2.805000   68.035000 3.945000 ;
      RECT   67.765000  4.535000   68.035000 5.355000 ;
      RECT   67.795000  1.725000   68.065000 2.455000 ;
      RECT   68.215000  0.265000   68.515000 0.635000 ;
      RECT   68.295000  1.505000   69.565000 1.745000 ;
      RECT   68.295000  1.745000   68.525000 2.455000 ;
      RECT   68.480000  1.015000   68.915000 1.325000 ;
      RECT   68.625000  2.805000   68.915000 3.970000 ;
      RECT   68.625000  4.630000   68.915000 5.355000 ;
      RECT   68.685000  0.375000   68.915000 1.015000 ;
      RECT   68.705000  1.925000   69.085000 2.635000 ;
      RECT   69.095000  2.975000   71.305000 3.145000 ;
      RECT   69.095000  3.145000   69.395000 5.015000 ;
      RECT   69.095000  5.015000   71.305000 5.185000 ;
      RECT   69.110000  0.995000   69.360000 1.325000 ;
      RECT   69.275000  0.085000   69.565000 0.815000 ;
      RECT   69.305000  1.745000   69.565000 2.455000 ;
      RECT   69.565000  3.315000   69.895000 3.775000 ;
      RECT   69.565000  3.775000   70.835000 3.945000 ;
      RECT   69.565000  4.115000   70.915000 4.365000 ;
      RECT   69.565000  4.535000   73.235000 4.715000 ;
      RECT   69.565000  4.715000   69.895000 4.845000 ;
      RECT   70.005000  0.085000   70.295000 0.810000 ;
      RECT   70.005000  1.470000   70.295000 2.635000 ;
      RECT   70.065000  3.145000   70.335000 3.605000 ;
      RECT   70.065000  4.895000   70.335000 5.015000 ;
      RECT   70.475000  1.665000   70.755000 2.635000 ;
      RECT   70.505000  3.315000   70.835000 3.775000 ;
      RECT   70.505000  4.715000   70.835000 4.845000 ;
      RECT   70.555000  0.085000   70.725000 0.555000 ;
      RECT   70.925000  0.255000   71.205000 2.465000 ;
      RECT   71.005000  3.145000   71.305000 3.945000 ;
      RECT   71.005000  4.890000   71.305000 5.015000 ;
      RECT   71.375000  0.655000   72.620000 0.825000 ;
      RECT   71.375000  0.825000   71.810000 1.690000 ;
      RECT   71.375000  1.690000   72.420000 1.920000 ;
      RECT   71.435000  2.220000   71.865000 2.635000 ;
      RECT   71.525000  2.805000   71.795000 3.945000 ;
      RECT   71.525000  4.890000   71.795000 5.355000 ;
      RECT   71.655000  0.085000   72.035000 0.445000 ;
      RECT   71.925000  4.115000   73.275000 4.365000 ;
      RECT   71.965000  2.975000   72.295000 3.775000 ;
      RECT   71.965000  3.775000   73.235000 3.945000 ;
      RECT   71.965000  4.715000   72.295000 5.185000 ;
      RECT   72.055000  1.920000   72.420000 2.465000 ;
      RECT   72.245000  0.995000   72.620000 1.410000 ;
      RECT   72.430000  0.255000   72.620000 0.655000 ;
      RECT   72.465000  2.805000   72.735000 3.605000 ;
      RECT   72.465000  4.895000   72.735000 5.355000 ;
      RECT   72.640000  1.670000   73.855000 1.935000 ;
      RECT   72.640000  1.935000   72.865000 2.465000 ;
      RECT   72.790000  0.365000   73.110000 1.325000 ;
      RECT   72.905000  2.975000   73.235000 3.775000 ;
      RECT   72.905000  4.715000   73.235000 5.185000 ;
      RECT   73.085000  2.125000   73.415000 2.635000 ;
      RECT   73.405000  2.805000   73.675000 3.945000 ;
      RECT   73.405000  4.535000   73.675000 5.355000 ;
      RECT   73.535000  0.085000   73.915000 0.565000 ;
      RECT   73.540000  0.750000   73.915000 1.325000 ;
      RECT   73.635000  1.935000   73.855000 2.465000 ;
      RECT   73.845000  2.975000   74.175000 4.115000 ;
      RECT   73.845000  4.115000   76.095000 4.365000 ;
      RECT   73.845000  4.365000   74.175000 5.185000 ;
      RECT   74.145000  0.085000   74.435000 0.810000 ;
      RECT   74.145000  1.470000   74.435000 2.635000 ;
      RECT   74.345000  2.805000   74.615000 3.945000 ;
      RECT   74.345000  4.535000   74.615000 5.355000 ;
      RECT   74.625000  0.085000   74.965000 0.445000 ;
      RECT   74.635000  1.935000   74.965000 2.635000 ;
      RECT   74.665000  0.615000   76.405000 0.785000 ;
      RECT   74.665000  0.785000   75.200000 1.585000 ;
      RECT   74.665000  1.585000   76.405000 1.755000 ;
      RECT   74.785000  2.975000   75.115000 3.775000 ;
      RECT   74.785000  3.775000   76.055000 3.945000 ;
      RECT   74.785000  4.535000   78.455000 4.715000 ;
      RECT   74.785000  4.715000   75.115000 5.185000 ;
      RECT   75.195000  1.755000   75.365000 2.185000 ;
      RECT   75.285000  2.805000   75.555000 3.605000 ;
      RECT   75.285000  4.895000   75.555000 5.355000 ;
      RECT   75.370000  0.995000   76.820000 1.325000 ;
      RECT   75.545000  0.085000   75.925000 0.445000 ;
      RECT   75.545000  1.935000   75.925000 2.635000 ;
      RECT   75.725000  2.975000   76.055000 3.775000 ;
      RECT   75.725000  4.715000   76.055000 5.185000 ;
      RECT   76.155000  1.755000   76.405000 2.185000 ;
      RECT   76.225000  2.805000   76.495000 3.945000 ;
      RECT   76.225000  4.890000   76.495000 5.355000 ;
      RECT   76.585000  1.515000   76.835000 2.635000 ;
      RECT   76.630000  0.085000   77.405000 0.445000 ;
      RECT   76.650000  0.615000   77.815000 0.670000 ;
      RECT   76.650000  0.670000   79.285000 0.785000 ;
      RECT   76.650000  0.785000   76.820000 0.995000 ;
      RECT   76.715000  2.975000   78.925000 3.145000 ;
      RECT   76.715000  3.145000   77.015000 3.945000 ;
      RECT   76.715000  4.890000   77.015000 5.015000 ;
      RECT   76.715000  5.015000   78.925000 5.185000 ;
      RECT   77.020000  0.995000   77.425000 1.525000 ;
      RECT   77.105000  4.115000   78.455000 4.365000 ;
      RECT   77.175000  1.695000   77.345000 2.295000 ;
      RECT   77.175000  2.295000   78.285000 2.465000 ;
      RECT   77.185000  3.315000   77.515000 3.775000 ;
      RECT   77.185000  3.775000   78.455000 3.945000 ;
      RECT   77.185000  4.715000   77.515000 4.845000 ;
      RECT   77.645000  0.255000   77.815000 0.615000 ;
      RECT   77.645000  0.785000   79.285000 0.840000 ;
      RECT   77.645000  0.840000   77.815000 2.125000 ;
      RECT   77.685000  3.145000   77.955000 3.605000 ;
      RECT   77.685000  4.895000   77.955000 5.015000 ;
      RECT   78.075000  0.085000   78.405000 0.445000 ;
      RECT   78.105000  1.445000   78.285000 1.850000 ;
      RECT   78.105000  1.850000   80.380000 2.020000 ;
      RECT   78.105000  2.020000   78.285000 2.295000 ;
      RECT   78.125000  3.315000   78.455000 3.775000 ;
      RECT   78.125000  4.715000   78.455000 4.845000 ;
      RECT   78.245000  1.010000   78.690000 1.275000 ;
      RECT   78.455000  2.275000   78.835000 2.635000 ;
      RECT   78.465000  1.275000   78.690000 1.510000 ;
      RECT   78.465000  1.510000   79.955000 1.680000 ;
      RECT   78.625000  3.145000   78.925000 4.115000 ;
      RECT   78.625000  4.115000   85.865000 4.365000 ;
      RECT   78.625000  4.365000   78.925000 5.015000 ;
      RECT   78.860000  1.010000   79.485000 1.275000 ;
      RECT   79.005000  0.405000   79.285000 0.670000 ;
      RECT   79.055000  2.020000   79.225000 2.465000 ;
      RECT   79.145000  2.805000   79.415000 3.945000 ;
      RECT   79.145000  4.535000   79.415000 5.355000 ;
      RECT   79.395000  2.275000   79.775000 2.635000 ;
      RECT   79.585000  2.975000   79.915000 3.775000 ;
      RECT   79.585000  3.775000   86.495000 3.945000 ;
      RECT   79.585000  4.535000   86.495000 4.715000 ;
      RECT   79.585000  4.715000   79.915000 5.185000 ;
      RECT   79.655000  1.055000   80.120000 1.290000 ;
      RECT   79.655000  1.290000   79.955000 1.510000 ;
      RECT   79.965000  0.085000   80.245000 0.885000 ;
      RECT   80.050000  2.020000   80.380000 2.395000 ;
      RECT   80.085000  2.805000   80.355000 3.605000 ;
      RECT   80.085000  4.895000   80.355000 5.355000 ;
      RECT   80.125000  1.460000   80.380000 1.850000 ;
      RECT   80.525000  2.975000   80.855000 3.775000 ;
      RECT   80.525000  4.715000   80.855000 5.185000 ;
      RECT   80.585000  0.085000   80.875000 0.810000 ;
      RECT   80.585000  1.470000   80.875000 2.635000 ;
      RECT   81.025000  2.805000   81.295000 3.605000 ;
      RECT   81.025000  4.895000   81.295000 5.355000 ;
      RECT   81.055000  0.675000   81.295000 1.325000 ;
      RECT   81.055000  1.495000   81.690000 1.685000 ;
      RECT   81.055000  1.685000   81.330000 2.455000 ;
      RECT   81.070000  0.085000   81.400000 0.475000 ;
      RECT   81.465000  0.645000   81.845000 0.825000 ;
      RECT   81.465000  0.825000   81.690000 1.495000 ;
      RECT   81.465000  2.975000   81.795000 3.775000 ;
      RECT   81.465000  4.715000   81.795000 5.185000 ;
      RECT   81.500000  1.855000   82.855000 2.025000 ;
      RECT   81.500000  2.025000   81.880000 2.455000 ;
      RECT   81.620000  0.265000   81.845000 0.645000 ;
      RECT   81.860000  0.995000   82.255000 1.325000 ;
      RECT   81.860000  1.525000   82.855000 1.855000 ;
      RECT   81.965000  2.805000   82.235000 3.605000 ;
      RECT   81.965000  4.895000   82.235000 5.355000 ;
      RECT   82.025000  0.375000   82.255000 0.995000 ;
      RECT   82.100000  2.195000   82.295000 2.635000 ;
      RECT   82.405000  2.975000   82.735000 3.775000 ;
      RECT   82.405000  4.715000   82.735000 5.185000 ;
      RECT   82.475000  2.025000   82.855000 2.455000 ;
      RECT   82.485000  0.995000   82.780000 1.325000 ;
      RECT   82.555000  0.085000   82.855000 0.815000 ;
      RECT   82.905000  2.805000   83.175000 3.605000 ;
      RECT   82.905000  4.890000   83.175000 5.355000 ;
      RECT   83.345000  0.085000   83.635000 0.810000 ;
      RECT   83.345000  1.470000   83.635000 2.635000 ;
      RECT   83.345000  2.975000   83.675000 3.775000 ;
      RECT   83.345000  4.715000   83.675000 5.185000 ;
      RECT   83.820000  0.085000   84.115000 0.865000 ;
      RECT   83.830000  1.855000   86.065000 2.025000 ;
      RECT   83.830000  2.025000   85.040000 2.105000 ;
      RECT   83.830000  2.105000   84.090000 2.465000 ;
      RECT   83.845000  2.805000   84.115000 3.605000 ;
      RECT   83.845000  4.895000   84.115000 5.355000 ;
      RECT   83.865000  1.035000   84.415000 1.495000 ;
      RECT   83.865000  1.495000   85.850000 1.675000 ;
      RECT   84.260000  2.275000   84.640000 2.635000 ;
      RECT   84.285000  2.975000   84.615000 3.775000 ;
      RECT   84.285000  4.715000   84.615000 5.185000 ;
      RECT   84.615000  0.995000   85.295000 1.325000 ;
      RECT   84.725000  0.255000   85.120000 0.615000 ;
      RECT   84.725000  0.615000   86.585000 0.785000 ;
      RECT   84.785000  2.805000   85.055000 3.605000 ;
      RECT   84.785000  4.895000   85.055000 5.355000 ;
      RECT   84.870000  2.105000   85.040000 2.465000 ;
      RECT   85.225000  2.975000   85.555000 3.775000 ;
      RECT   85.225000  4.715000   85.555000 5.185000 ;
      RECT   85.345000  2.195000   85.515000 2.635000 ;
      RECT   85.475000  1.075000   85.850000 1.495000 ;
      RECT   85.630000  0.085000   86.010000 0.445000 ;
      RECT   85.725000  2.805000   85.995000 3.605000 ;
      RECT   85.725000  4.895000   85.995000 5.355000 ;
      RECT   85.735000  2.025000   86.065000 2.285000 ;
      RECT   85.735000  2.285000   87.110000 2.465000 ;
      RECT   86.085000  3.945000   86.495000 4.535000 ;
      RECT   86.130000  0.785000   86.585000 1.330000 ;
      RECT   86.165000  2.975000   86.495000 3.775000 ;
      RECT   86.165000  4.715000   86.495000 5.185000 ;
      RECT   86.235000  1.330000   86.585000 2.115000 ;
      RECT   86.265000  0.255000   86.585000 0.615000 ;
      RECT   86.665000  2.805000   86.935000 3.945000 ;
      RECT   86.665000  4.535000   86.935000 5.355000 ;
      RECT   86.755000  0.995000   87.255000 1.625000 ;
      RECT   86.805000  1.795000   87.110000 2.285000 ;
      RECT   86.815000  0.085000   87.145000 0.825000 ;
      RECT   87.485000  0.085000   87.775000 0.810000 ;
      RECT   87.485000  1.470000   87.775000 2.635000 ;
      RECT   87.485000  2.805000   87.775000 3.970000 ;
      RECT   87.485000  4.630000   87.775000 5.355000 ;
      RECT   87.950000  0.085000   88.285000 0.805000 ;
      RECT   87.950000  0.995000   88.260000 1.035000 ;
      RECT   87.950000  1.035000   89.440000 1.415000 ;
      RECT   87.950000  4.555000   91.025000 4.725000 ;
      RECT   87.950000  4.725000   88.285000 5.185000 ;
      RECT   87.985000  2.805000   88.255000 3.945000 ;
      RECT   88.040000  1.795000   88.235000 2.215000 ;
      RECT   88.040000  2.215000   90.175000 2.465000 ;
      RECT   88.255000  4.115000   90.625000 4.385000 ;
      RECT   88.425000  2.975000   88.755000 3.775000 ;
      RECT   88.425000  3.775000   93.455000 3.945000 ;
      RECT   88.455000  4.895000   88.725000 5.355000 ;
      RECT   88.490000  1.585000   89.940000 1.705000 ;
      RECT   88.490000  1.705000   89.755000 2.035000 ;
      RECT   88.505000  0.370000   88.695000 0.615000 ;
      RECT   88.505000  0.615000   89.655000 0.695000 ;
      RECT   88.505000  0.695000   92.165000 0.865000 ;
      RECT   88.865000  0.085000   89.245000 0.445000 ;
      RECT   88.865000  2.205000   90.175000 2.215000 ;
      RECT   88.895000  4.725000   89.225000 5.185000 ;
      RECT   88.925000  2.805000   89.195000 3.605000 ;
      RECT   89.365000  2.975000   89.695000 3.775000 ;
      RECT   89.395000  4.895000   89.665000 5.355000 ;
      RECT   89.465000  0.255000   89.655000 0.615000 ;
      RECT   89.610000  0.865000   92.165000 0.895000 ;
      RECT   89.610000  0.895000   89.940000 1.585000 ;
      RECT   89.835000  4.725000   90.165000 5.185000 ;
      RECT   89.845000  0.085000   90.175000 0.525000 ;
      RECT   89.865000  2.805000   90.135000 3.605000 ;
      RECT   89.975000  1.875000   94.085000 2.105000 ;
      RECT   89.975000  2.105000   90.175000 2.205000 ;
      RECT   90.110000  1.065000   90.505000 1.480000 ;
      RECT   90.110000  1.480000   93.930000 1.705000 ;
      RECT   90.305000  2.975000   90.635000 3.775000 ;
      RECT   90.335000  0.675000   92.165000 0.695000 ;
      RECT   90.335000  4.895000   90.605000 5.355000 ;
      RECT   90.345000  0.255000   92.645000 0.505000 ;
      RECT   90.345000  2.275000   90.725000 2.635000 ;
      RECT   90.675000  1.065000   92.260000 1.310000 ;
      RECT   90.775000  4.725000   91.025000 4.975000 ;
      RECT   90.775000  4.975000   93.925000 5.185000 ;
      RECT   90.805000  2.805000   91.075000 3.605000 ;
      RECT   90.945000  2.105000   91.135000 2.465000 ;
      RECT   91.195000  3.945000   91.495000 4.555000 ;
      RECT   91.195000  4.555000   93.455000 4.805000 ;
      RECT   91.245000  2.975000   91.575000 3.775000 ;
      RECT   91.305000  2.275000   91.685000 2.635000 ;
      RECT   91.665000  4.115000   93.015000 4.385000 ;
      RECT   91.745000  2.805000   92.015000 3.605000 ;
      RECT   91.905000  2.105000   92.095000 2.465000 ;
      RECT   92.185000  2.975000   92.515000 3.775000 ;
      RECT   92.265000  2.275000   92.645000 2.635000 ;
      RECT   92.385000  0.505000   92.645000 0.735000 ;
      RECT   92.385000  0.735000   93.605000 0.905000 ;
      RECT   92.535000  1.075000   93.930000 1.480000 ;
      RECT   92.685000  2.805000   92.955000 3.605000 ;
      RECT   92.865000  0.085000   93.055000 0.565000 ;
      RECT   92.865000  2.105000   93.045000 2.465000 ;
      RECT   93.125000  2.975000   93.455000 3.775000 ;
      RECT   93.185000  3.945000   93.455000 4.115000 ;
      RECT   93.185000  4.115000   93.775000 4.385000 ;
      RECT   93.185000  4.385000   93.455000 4.555000 ;
      RECT   93.225000  0.255000   93.605000 0.735000 ;
      RECT   93.225000  2.275000   93.605000 2.635000 ;
      RECT   93.625000  2.805000   93.895000 3.945000 ;
      RECT   93.625000  4.555000   93.925000 4.975000 ;
      RECT   93.825000  0.085000   94.085000 0.885000 ;
      RECT   93.825000  2.105000   94.085000 2.465000 ;
      RECT   94.385000  0.085000   94.675000 0.810000 ;
      RECT   94.385000  1.470000   94.675000 2.635000 ;
      RECT   94.385000  2.805000   94.675000 3.970000 ;
      RECT   94.385000  4.630000   94.675000 5.355000 ;
      RECT   94.845000  1.075000   95.195000 1.285000 ;
      RECT   94.850000  4.555000  100.745000 4.725000 ;
      RECT   94.850000  4.725000   95.185000 5.185000 ;
      RECT   94.885000  2.805000   95.155000 3.945000 ;
      RECT   94.930000  0.255000   95.105000 0.735000 ;
      RECT   94.930000  0.735000   96.095000 0.905000 ;
      RECT   94.935000  1.455000   97.210000 1.495000 ;
      RECT   94.935000  1.495000   98.295000 1.625000 ;
      RECT   94.935000  1.625000   95.105000 2.465000 ;
      RECT   95.095000  4.115000  100.525000 4.385000 ;
      RECT   95.275000  0.085000   95.655000 0.565000 ;
      RECT   95.275000  1.795000   95.575000 2.295000 ;
      RECT   95.275000  2.295000   96.595000 2.465000 ;
      RECT   95.325000  2.975000   95.655000 3.775000 ;
      RECT   95.325000  3.775000  105.995000 3.945000 ;
      RECT   95.355000  4.895000   95.625000 5.355000 ;
      RECT   95.365000  1.075000   95.915000 1.285000 ;
      RECT   95.795000  4.725000   96.125000 5.185000 ;
      RECT   95.825000  2.805000   96.095000 3.605000 ;
      RECT   95.875000  1.795000   96.935000 1.835000 ;
      RECT   95.875000  1.835000   97.585000 2.045000 ;
      RECT   95.875000  2.045000   96.100000 2.125000 ;
      RECT   95.925000  0.255000   97.540000 0.505000 ;
      RECT   95.925000  0.505000   96.095000 0.735000 ;
      RECT   96.085000  1.075000   96.575000 1.285000 ;
      RECT   96.215000  2.255000   96.595000 2.295000 ;
      RECT   96.265000  2.975000   96.595000 3.775000 ;
      RECT   96.285000  0.675000   96.575000 1.075000 ;
      RECT   96.295000  4.895000   96.565000 5.355000 ;
      RECT   96.735000  4.725000   97.065000 5.185000 ;
      RECT   96.745000  0.675000   97.110000 1.075000 ;
      RECT   96.745000  1.075000   97.185000 1.285000 ;
      RECT   96.765000  2.805000   97.035000 3.605000 ;
      RECT   96.785000  2.215000   97.115000 2.635000 ;
      RECT   97.060000  1.625000   98.295000 1.665000 ;
      RECT   97.205000  2.975000   97.535000 3.775000 ;
      RECT   97.235000  4.895000   97.505000 5.355000 ;
      RECT   97.335000  2.045000   97.585000 2.465000 ;
      RECT   97.340000  0.505000   97.540000 0.655000 ;
      RECT   97.340000  0.655000   98.295000 0.825000 ;
      RECT   97.430000  0.995000   97.835000 1.325000 ;
      RECT   97.675000  4.725000   98.005000 5.185000 ;
      RECT   97.705000  2.805000   97.975000 3.605000 ;
      RECT   97.790000  0.085000   98.120000 0.485000 ;
      RECT   97.805000  1.875000   98.135000 2.635000 ;
      RECT   98.015000  0.825000   98.295000 1.495000 ;
      RECT   98.145000  2.975000   98.475000 3.775000 ;
      RECT   98.175000  4.895000   98.445000 5.355000 ;
      RECT   98.525000  0.085000   98.815000 0.810000 ;
      RECT   98.525000  1.470000   98.815000 2.635000 ;
      RECT   98.615000  4.725000   98.945000 5.185000 ;
      RECT   98.645000  2.805000   98.915000 3.605000 ;
      RECT   98.990000  1.075000   99.320000 1.615000 ;
      RECT   98.990000  1.795000   99.335000 2.295000 ;
      RECT   98.990000  2.295000  100.275000 2.465000 ;
      RECT   99.005000  0.085000   99.255000 0.895000 ;
      RECT   99.085000  2.975000   99.415000 3.775000 ;
      RECT   99.115000  4.895000   99.385000 5.355000 ;
      RECT   99.425000  0.305000   99.805000 0.725000 ;
      RECT   99.425000  0.725000  103.695000 0.865000 ;
      RECT   99.505000  0.865000  103.695000 0.905000 ;
      RECT   99.505000  0.905000   99.805000 2.125000 ;
      RECT   99.555000  4.725000   99.885000 5.185000 ;
      RECT   99.585000  2.805000   99.855000 3.605000 ;
      RECT  100.025000  0.085000  100.715000 0.555000 ;
      RECT  100.025000  1.495000  100.275000 1.785000 ;
      RECT  100.025000  1.785000  102.165000 1.955000 ;
      RECT  100.025000  1.955000  100.275000 2.295000 ;
      RECT  100.025000  2.975000  100.355000 3.775000 ;
      RECT  100.055000  4.895000  100.325000 5.355000 ;
      RECT  100.495000  4.725000  100.745000 4.975000 ;
      RECT  100.495000  4.975000  106.465000 5.185000 ;
      RECT  100.505000  2.125000  100.755000 2.295000 ;
      RECT  100.505000  2.295000  102.675000 2.465000 ;
      RECT  100.525000  2.805000  100.795000 3.605000 ;
      RECT  100.630000  1.075000  101.090000 1.445000 ;
      RECT  100.630000  1.445000  102.465000 1.615000 ;
      RECT  100.805000  3.945000  101.215000 4.385000 ;
      RECT  100.885000  0.255000  102.205000 0.475000 ;
      RECT  100.915000  4.385000  101.215000 4.555000 ;
      RECT  100.915000  4.555000  105.995000 4.805000 ;
      RECT  100.965000  2.975000  101.295000 3.775000 ;
      RECT  100.975000  1.955000  101.225000 2.125000 ;
      RECT  101.260000  1.075000  101.915000 1.275000 ;
      RECT  101.335000  0.645000  101.735000 0.725000 ;
      RECT  101.385000  4.115000  105.455000 4.385000 ;
      RECT  101.445000  2.125000  101.695000 2.295000 ;
      RECT  101.465000  2.805000  101.735000 3.605000 ;
      RECT  101.905000  2.975000  102.235000 3.775000 ;
      RECT  101.915000  1.955000  102.165000 2.125000 ;
      RECT  102.085000  1.075000  102.465000 1.445000 ;
      RECT  102.405000  2.805000  102.675000 3.605000 ;
      RECT  102.425000  1.785000  104.595000 1.955000 ;
      RECT  102.425000  1.955000  102.675000 2.295000 ;
      RECT  102.470000  0.085000  102.640000 0.555000 ;
      RECT  102.635000  1.075000  102.965000 1.445000 ;
      RECT  102.635000  1.445000  104.170000 1.615000 ;
      RECT  102.845000  0.255000  104.165000 0.475000 ;
      RECT  102.845000  2.975000  103.175000 3.775000 ;
      RECT  102.935000  2.125000  103.185000 2.635000 ;
      RECT  103.135000  1.075000  103.815000 1.275000 ;
      RECT  103.315000  0.645000  103.695000 0.725000 ;
      RECT  103.345000  2.805000  103.615000 3.605000 ;
      RECT  103.405000  1.955000  103.655000 2.465000 ;
      RECT  103.785000  2.975000  104.115000 3.775000 ;
      RECT  103.875000  2.125000  104.125000 2.635000 ;
      RECT  103.915000  0.475000  104.165000 0.905000 ;
      RECT  104.000000  1.075000  104.785000 1.275000 ;
      RECT  104.000000  1.275000  104.170000 1.445000 ;
      RECT  104.285000  2.805000  104.555000 3.605000 ;
      RECT  104.385000  0.085000  104.555000 0.905000 ;
      RECT  104.390000  1.455000  104.595000 1.785000 ;
      RECT  104.390000  1.955000  104.595000 2.465000 ;
      RECT  104.725000  2.975000  105.055000 3.775000 ;
      RECT  104.965000  0.085000  105.255000 0.810000 ;
      RECT  104.965000  1.470000  105.255000 2.635000 ;
      RECT  105.225000  2.805000  105.495000 3.605000 ;
      RECT  105.430000  1.075000  106.775000 1.275000 ;
      RECT  105.430000  1.445000  105.745000 2.295000 ;
      RECT  105.430000  2.295000  107.665000 2.465000 ;
      RECT  105.455000  0.085000  105.705000 0.895000 ;
      RECT  105.665000  2.975000  105.995000 3.775000 ;
      RECT  105.725000  3.945000  105.995000 4.115000 ;
      RECT  105.725000  4.115000  106.195000 4.385000 ;
      RECT  105.725000  4.385000  105.995000 4.555000 ;
      RECT  105.875000  0.255000  106.255000 0.725000 ;
      RECT  105.875000  0.725000  107.195000 0.905000 ;
      RECT  105.965000  1.445000  107.195000 1.615000 ;
      RECT  105.965000  1.615000  106.215000 2.125000 ;
      RECT  106.165000  2.805000  106.435000 3.945000 ;
      RECT  106.215000  4.555000  106.465000 4.975000 ;
      RECT  106.435000  1.785000  106.685000 2.295000 ;
      RECT  106.475000  0.085000  106.645000 0.555000 ;
      RECT  106.805000  2.805000  107.095000 3.970000 ;
      RECT  106.805000  4.630000  107.095000 5.355000 ;
      RECT  106.815000  0.255000  107.195000 0.725000 ;
      RECT  106.905000  1.615000  107.155000 2.125000 ;
      RECT  106.995000  0.905000  107.195000 1.095000 ;
      RECT  106.995000  1.095000  108.935000 1.275000 ;
      RECT  106.995000  1.275000  107.195000 1.445000 ;
      RECT  107.275000  4.555000  115.045000 4.725000 ;
      RECT  107.275000  4.725000  107.605000 5.185000 ;
      RECT  107.305000  2.805000  107.575000 3.945000 ;
      RECT  107.415000  0.085000  107.585000 0.645000 ;
      RECT  107.415000  0.645000  108.545000 0.925000 ;
      RECT  107.415000  1.445000  108.670000 1.615000 ;
      RECT  107.415000  1.615000  107.665000 2.295000 ;
      RECT  107.575000  4.115000  114.705000 4.385000 ;
      RECT  107.745000  2.975000  108.075000 3.775000 ;
      RECT  107.745000  3.775000  122.175000 3.945000 ;
      RECT  107.775000  0.255000  111.525000 0.425000 ;
      RECT  107.775000  0.425000  108.200000 0.475000 ;
      RECT  107.775000  4.895000  108.045000 5.355000 ;
      RECT  107.905000  1.795000  108.155000 2.215000 ;
      RECT  107.905000  2.215000  111.995000 2.465000 ;
      RECT  108.215000  4.725000  108.545000 5.185000 ;
      RECT  108.245000  2.805000  108.515000 3.605000 ;
      RECT  108.375000  0.595000  108.545000 0.645000 ;
      RECT  108.375000  1.615000  108.670000 1.835000 ;
      RECT  108.375000  1.835000  111.525000 2.045000 ;
      RECT  108.675000  0.425000  111.525000 0.475000 ;
      RECT  108.685000  2.975000  109.015000 3.775000 ;
      RECT  108.715000  0.645000  111.620000 0.735000 ;
      RECT  108.715000  0.735000  113.925000 0.820000 ;
      RECT  108.715000  0.820000  108.935000 1.095000 ;
      RECT  108.715000  4.895000  108.985000 5.355000 ;
      RECT  109.105000  0.995000  109.505000 1.325000 ;
      RECT  109.155000  4.725000  109.485000 5.185000 ;
      RECT  109.185000  2.805000  109.455000 3.605000 ;
      RECT  109.285000  1.325000  109.505000 1.445000 ;
      RECT  109.285000  1.445000  111.750000 1.615000 ;
      RECT  109.625000  2.975000  109.955000 3.775000 ;
      RECT  109.655000  4.895000  109.925000 5.355000 ;
      RECT  109.675000  0.995000  111.225000 1.275000 ;
      RECT  110.095000  4.725000  110.425000 5.185000 ;
      RECT  110.125000  2.805000  110.395000 3.605000 ;
      RECT  110.565000  2.975000  110.895000 3.775000 ;
      RECT  110.595000  4.895000  110.865000 5.355000 ;
      RECT  111.035000  4.725000  111.365000 5.185000 ;
      RECT  111.065000  2.805000  111.335000 3.605000 ;
      RECT  111.405000  1.075000  111.750000 1.445000 ;
      RECT  111.450000  0.820000  112.470000 0.905000 ;
      RECT  111.505000  2.975000  111.835000 3.775000 ;
      RECT  111.535000  4.895000  111.805000 5.355000 ;
      RECT  111.745000  1.785000  114.865000 2.045000 ;
      RECT  111.745000  2.045000  111.995000 2.215000 ;
      RECT  111.795000  0.085000  111.965000 0.555000 ;
      RECT  111.925000  1.075000  112.305000 1.445000 ;
      RECT  111.925000  1.445000  114.475000 1.615000 ;
      RECT  111.975000  4.725000  112.305000 5.185000 ;
      RECT  112.005000  2.805000  112.275000 3.605000 ;
      RECT  112.135000  0.255000  114.395000 0.475000 ;
      RECT  112.165000  2.215000  114.425000 2.635000 ;
      RECT  112.300000  0.645000  113.925000 0.735000 ;
      RECT  112.445000  2.975000  112.775000 3.775000 ;
      RECT  112.475000  4.895000  112.745000 5.355000 ;
      RECT  112.485000  1.075000  114.095000 1.275000 ;
      RECT  112.915000  4.725000  113.245000 5.185000 ;
      RECT  112.945000  2.805000  113.215000 3.605000 ;
      RECT  113.385000  2.975000  113.715000 3.775000 ;
      RECT  113.415000  4.895000  113.685000 5.355000 ;
      RECT  113.855000  4.725000  114.185000 5.185000 ;
      RECT  113.885000  2.805000  114.155000 3.605000 ;
      RECT  114.145000  0.475000  114.395000 0.725000 ;
      RECT  114.145000  0.725000  115.335000 0.905000 ;
      RECT  114.305000  1.075000  115.740000 1.275000 ;
      RECT  114.305000  1.275000  114.475000 1.445000 ;
      RECT  114.325000  2.975000  114.655000 3.775000 ;
      RECT  114.355000  4.895000  114.625000 5.355000 ;
      RECT  114.615000  0.085000  114.785000 0.555000 ;
      RECT  114.615000  2.045000  114.785000 2.465000 ;
      RECT  114.695000  1.445000  115.765000 1.615000 ;
      RECT  114.695000  1.615000  114.865000 1.785000 ;
      RECT  114.795000  4.725000  115.045000 4.975000 ;
      RECT  114.795000  4.975000  122.645000 5.185000 ;
      RECT  114.825000  2.805000  115.095000 3.605000 ;
      RECT  114.955000  0.255000  115.335000 0.725000 ;
      RECT  115.085000  1.795000  115.255000 2.635000 ;
      RECT  115.105000  3.945000  115.515000 4.385000 ;
      RECT  115.215000  4.385000  115.515000 4.555000 ;
      RECT  115.215000  4.555000  122.175000 4.805000 ;
      RECT  115.265000  2.975000  115.595000 3.775000 ;
      RECT  115.505000  0.085000  115.675000 0.905000 ;
      RECT  115.515000  1.615000  115.765000 2.465000 ;
      RECT  115.685000  4.115000  121.455000 4.385000 ;
      RECT  115.765000  2.805000  116.035000 3.605000 ;
      RECT  116.005000  0.085000  116.295000 0.810000 ;
      RECT  116.005000  1.470000  116.295000 2.635000 ;
      RECT  116.205000  2.975000  116.535000 3.775000 ;
      RECT  116.465000  1.000000  116.975000 1.315000 ;
      RECT  116.475000  0.255000  116.805000 0.645000 ;
      RECT  116.475000  0.645000  119.355000 0.815000 ;
      RECT  116.475000  1.485000  118.035000 1.795000 ;
      RECT  116.475000  1.795000  116.725000 2.295000 ;
      RECT  116.705000  2.805000  116.975000 3.605000 ;
      RECT  116.945000  2.055000  117.275000 2.295000 ;
      RECT  116.945000  2.295000  118.845000 2.465000 ;
      RECT  117.145000  1.000000  117.615000 1.315000 ;
      RECT  117.145000  2.975000  117.475000 3.775000 ;
      RECT  117.305000  0.085000  118.085000 0.465000 ;
      RECT  117.645000  2.805000  117.915000 3.605000 ;
      RECT  117.785000  0.815000  118.035000 1.485000 ;
      RECT  118.085000  2.975000  118.415000 3.775000 ;
      RECT  118.205000  1.500000  120.405000 1.735000 ;
      RECT  118.205000  1.735000  119.315000 1.830000 ;
      RECT  118.265000  1.000000  118.625000 1.330000 ;
      RECT  118.550000  2.135000  118.845000 2.295000 ;
      RECT  118.585000  2.805000  118.855000 3.605000 ;
      RECT  118.790000  0.295000  119.355000 0.645000 ;
      RECT  118.795000  1.000000  119.115000 1.330000 ;
      RECT  119.025000  2.975000  119.355000 3.775000 ;
      RECT  119.065000  1.830000  119.315000 2.250000 ;
      RECT  119.285000  1.000000  119.685000 1.330000 ;
      RECT  119.525000  2.805000  119.795000 3.605000 ;
      RECT  119.535000  1.905000  119.865000 2.635000 ;
      RECT  119.855000  1.000000  120.375000 1.330000 ;
      RECT  119.935000  0.085000  120.345000 0.815000 ;
      RECT  119.965000  2.975000  120.295000 3.775000 ;
      RECT  120.145000  1.735000  120.405000 2.250000 ;
      RECT  120.465000  2.805000  120.735000 3.605000 ;
      RECT  120.605000  0.085000  120.895000 0.810000 ;
      RECT  120.605000  1.470000  120.895000 2.635000 ;
      RECT  120.905000  2.975000  121.235000 3.775000 ;
      RECT  121.065000  1.075000  121.605000 1.275000 ;
      RECT  121.070000  0.085000  121.575000 0.850000 ;
      RECT  121.070000  1.495000  124.015000 1.715000 ;
      RECT  121.070000  1.715000  121.325000 2.245000 ;
      RECT  121.070000  2.245000  121.405000 2.465000 ;
      RECT  121.405000  2.805000  121.675000 3.605000 ;
      RECT  121.545000  1.885000  123.375000 2.085000 ;
      RECT  121.795000  1.075000  122.265000 1.285000 ;
      RECT  121.845000  2.975000  122.175000 3.775000 ;
      RECT  121.850000  0.255000  123.260000 0.465000 ;
      RECT  121.905000  3.945000  122.175000 4.115000 ;
      RECT  121.905000  4.115000  122.295000 4.385000 ;
      RECT  121.905000  4.385000  122.175000 4.555000 ;
      RECT  122.045000  0.675000  122.265000 1.075000 ;
      RECT  122.345000  2.805000  122.615000 3.945000 ;
      RECT  122.395000  4.555000  122.645000 4.975000 ;
      RECT  122.505000  0.675000  122.725000 1.065000 ;
      RECT  122.505000  1.065000  123.065000 1.285000 ;
      RECT  122.520000  2.255000  122.875000 2.635000 ;
      RECT  122.905000  2.805000  123.195000 3.970000 ;
      RECT  122.905000  4.630000  123.195000 5.355000 ;
      RECT  123.045000  2.085000  123.375000 2.465000 ;
      RECT  123.090000  0.465000  123.260000 0.615000 ;
      RECT  123.090000  0.615000  124.015000 0.785000 ;
      RECT  123.255000  0.980000  123.605000 1.285000 ;
      RECT  123.395000  2.975000  123.685000 3.815000 ;
      RECT  123.395000  3.815000  126.505000 3.985000 ;
      RECT  123.395000  4.535000  123.695000 5.355000 ;
      RECT  123.565000  0.085000  123.895000 0.445000 ;
      RECT  123.565000  1.935000  123.895000 2.635000 ;
      RECT  123.785000  4.155000  126.155000 4.365000 ;
      RECT  123.845000  0.785000  124.015000 1.495000 ;
      RECT  123.865000  4.535000  135.115000 4.715000 ;
      RECT  123.865000  4.715000  124.195000 5.185000 ;
      RECT  123.905000  2.805000  124.155000 3.645000 ;
      RECT  124.255000  0.255000  124.515000 0.585000 ;
      RECT  124.255000  1.785000  124.515000 2.465000 ;
      RECT  124.345000  0.585000  124.515000 1.785000 ;
      RECT  124.365000  4.885000  124.635000 5.355000 ;
      RECT  124.375000  2.975000  124.625000 3.815000 ;
      RECT  124.745000  0.085000  125.035000 0.810000 ;
      RECT  124.745000  1.470000  125.035000 2.635000 ;
      RECT  124.805000  4.715000  125.135000 5.185000 ;
      RECT  124.845000  2.805000  125.095000 3.645000 ;
      RECT  125.210000  1.075000  125.745000 1.275000 ;
      RECT  125.215000  0.085000  125.715000 0.850000 ;
      RECT  125.215000  1.455000  128.135000 1.625000 ;
      RECT  125.215000  1.625000  125.545000 2.295000 ;
      RECT  125.215000  2.295000  126.485000 2.465000 ;
      RECT  125.305000  4.885000  125.575000 5.355000 ;
      RECT  125.315000  2.975000  125.565000 3.815000 ;
      RECT  125.745000  4.715000  126.075000 5.185000 ;
      RECT  125.765000  1.795000  127.500000 2.035000 ;
      RECT  125.765000  2.035000  125.995000 2.125000 ;
      RECT  125.785000  2.805000  126.035000 3.645000 ;
      RECT  125.935000  1.075000  126.460000 1.285000 ;
      RECT  125.990000  0.255000  127.415000 0.505000 ;
      RECT  126.155000  2.255000  126.485000 2.295000 ;
      RECT  126.185000  0.675000  126.460000 1.075000 ;
      RECT  126.245000  4.885000  126.515000 5.355000 ;
      RECT  126.255000  2.975000  129.365000 3.145000 ;
      RECT  126.255000  3.145000  126.505000 3.815000 ;
      RECT  126.605000  4.155000  128.975000 4.365000 ;
      RECT  126.645000  0.675000  126.940000 1.075000 ;
      RECT  126.645000  1.075000  127.060000 1.285000 ;
      RECT  126.675000  2.215000  127.030000 2.635000 ;
      RECT  126.685000  4.715000  127.015000 5.185000 ;
      RECT  126.725000  3.315000  126.975000 3.815000 ;
      RECT  126.725000  3.815000  132.195000 3.985000 ;
      RECT  127.185000  4.885000  127.455000 5.355000 ;
      RECT  127.195000  3.145000  127.445000 3.645000 ;
      RECT  127.245000  0.505000  127.415000 0.735000 ;
      RECT  127.245000  0.735000  128.135000 0.905000 ;
      RECT  127.250000  2.035000  127.500000 2.465000 ;
      RECT  127.280000  1.075000  127.735000 1.275000 ;
      RECT  127.625000  0.085000  128.005000 0.565000 ;
      RECT  127.625000  4.715000  127.955000 5.185000 ;
      RECT  127.665000  3.315000  127.915000 3.815000 ;
      RECT  127.720000  1.875000  128.050000 2.635000 ;
      RECT  127.965000  0.905000  128.135000 1.455000 ;
      RECT  128.125000  4.885000  128.395000 5.355000 ;
      RECT  128.135000  3.145000  128.385000 3.645000 ;
      RECT  128.270000  0.255000  128.680000 0.585000 ;
      RECT  128.270000  1.785000  128.680000 2.465000 ;
      RECT  128.360000  0.585000  128.680000 1.785000 ;
      RECT  128.565000  4.715000  128.895000 5.185000 ;
      RECT  128.605000  3.315000  128.855000 3.815000 ;
      RECT  128.875000  0.085000  129.045000 0.985000 ;
      RECT  128.875000  1.445000  129.045000 2.635000 ;
      RECT  129.065000  4.885000  129.855000 5.355000 ;
      RECT  129.075000  3.145000  129.365000 3.645000 ;
      RECT  129.345000  0.085000  129.635000 0.810000 ;
      RECT  129.345000  1.470000  129.635000 2.635000 ;
      RECT  129.555000  2.975000  135.535000 3.145000 ;
      RECT  129.555000  3.145000  129.845000 3.645000 ;
      RECT  129.805000  0.725000  131.640000 0.905000 ;
      RECT  129.805000  0.905000  130.090000 1.445000 ;
      RECT  129.805000  1.445000  131.600000 1.615000 ;
      RECT  129.940000  1.825000  130.190000 2.635000 ;
      RECT  129.945000  4.155000  132.315000 4.365000 ;
      RECT  129.980000  0.085000  130.150000 0.555000 ;
      RECT  130.025000  4.715000  130.355000 5.185000 ;
      RECT  130.065000  3.315000  130.315000 3.815000 ;
      RECT  130.260000  1.075000  132.150000 1.275000 ;
      RECT  130.320000  0.265000  130.700000 0.725000 ;
      RECT  130.410000  1.615000  130.660000 2.465000 ;
      RECT  130.525000  4.885000  130.795000 5.355000 ;
      RECT  130.535000  3.145000  130.785000 3.645000 ;
      RECT  130.880000  1.795000  131.130000 2.635000 ;
      RECT  130.920000  0.085000  131.090000 0.555000 ;
      RECT  130.965000  4.715000  131.295000 5.185000 ;
      RECT  131.005000  3.315000  131.255000 3.815000 ;
      RECT  131.260000  0.255000  131.640000 0.725000 ;
      RECT  131.350000  1.615000  131.600000 2.465000 ;
      RECT  131.465000  4.885000  131.735000 5.355000 ;
      RECT  131.475000  3.145000  131.725000 3.645000 ;
      RECT  131.820000  1.275000  132.150000 1.785000 ;
      RECT  131.820000  1.785000  134.000000 1.955000 ;
      RECT  131.820000  2.125000  132.070000 2.635000 ;
      RECT  131.860000  0.085000  132.550000 0.555000 ;
      RECT  131.860000  0.735000  135.530000 0.905000 ;
      RECT  131.860000  0.905000  132.150000 1.075000 ;
      RECT  131.905000  4.715000  132.235000 5.185000 ;
      RECT  131.945000  3.315000  132.195000 3.815000 ;
      RECT  132.340000  1.075000  132.925000 1.445000 ;
      RECT  132.340000  1.445000  134.300000 1.615000 ;
      RECT  132.340000  2.125000  132.590000 2.295000 ;
      RECT  132.340000  2.295000  134.550000 2.465000 ;
      RECT  132.405000  4.885000  132.675000 5.355000 ;
      RECT  132.415000  3.145000  132.665000 3.985000 ;
      RECT  132.675000  4.155000  134.365000 4.365000 ;
      RECT  132.720000  0.255000  134.040000 0.475000 ;
      RECT  132.810000  1.955000  133.060000 2.125000 ;
      RECT  132.845000  4.715000  133.175000 5.185000 ;
      RECT  132.885000  3.315000  133.135000 3.815000 ;
      RECT  132.885000  3.815000  135.115000 3.985000 ;
      RECT  133.095000  1.075000  133.750000 1.275000 ;
      RECT  133.140000  0.645000  133.625000 0.735000 ;
      RECT  133.280000  2.125000  133.530000 2.295000 ;
      RECT  133.345000  4.885000  133.615000 5.355000 ;
      RECT  133.355000  3.145000  133.605000 3.645000 ;
      RECT  133.750000  1.955000  134.000000 2.125000 ;
      RECT  133.785000  4.715000  134.115000 5.185000 ;
      RECT  133.825000  3.315000  134.075000 3.815000 ;
      RECT  133.920000  1.075000  134.300000 1.445000 ;
      RECT  134.220000  1.785000  136.430000 1.955000 ;
      RECT  134.220000  1.955000  134.550000 2.295000 ;
      RECT  134.285000  4.885000  134.555000 5.355000 ;
      RECT  134.295000  3.145000  134.545000 3.645000 ;
      RECT  134.305000  0.085000  134.475000 0.555000 ;
      RECT  134.470000  1.075000  134.850000 1.445000 ;
      RECT  134.470000  1.445000  136.005000 1.615000 ;
      RECT  134.680000  0.255000  136.000000 0.475000 ;
      RECT  134.725000  3.315000  135.115000 3.815000 ;
      RECT  134.725000  3.985000  135.115000 4.535000 ;
      RECT  134.725000  4.715000  135.115000 5.185000 ;
      RECT  134.770000  2.125000  135.020000 2.635000 ;
      RECT  135.070000  1.075000  135.615000 1.275000 ;
      RECT  135.105000  0.645000  135.530000 0.735000 ;
      RECT  135.240000  1.955000  135.490000 2.465000 ;
      RECT  135.285000  3.145000  135.535000 3.985000 ;
      RECT  135.285000  4.535000  135.535000 5.355000 ;
      RECT  135.710000  2.125000  135.960000 2.635000 ;
      RECT  135.750000  0.475000  136.000000 0.895000 ;
      RECT  135.785000  2.805000  136.075000 3.970000 ;
      RECT  135.785000  4.630000  136.075000 5.355000 ;
      RECT  135.835000  1.075000  136.535000 1.275000 ;
      RECT  135.835000  1.275000  136.005000 1.445000 ;
      RECT  136.220000  0.085000  136.390000 0.895000 ;
      RECT  136.225000  1.455000  136.430000 1.785000 ;
      RECT  136.225000  1.955000  136.430000 2.465000 ;
      RECT  136.255000  2.975000  136.585000 3.815000 ;
      RECT  136.255000  3.815000  140.305000 3.985000 ;
      RECT  136.295000  4.535000  136.555000 5.355000 ;
      RECT  136.565000  4.155000  139.955000 4.365000 ;
      RECT  136.705000  0.085000  136.995000 0.810000 ;
      RECT  136.705000  1.470000  136.995000 2.635000 ;
      RECT  136.725000  4.535000  151.675000 4.715000 ;
      RECT  136.725000  4.715000  137.055000 5.185000 ;
      RECT  136.765000  2.805000  137.015000 3.645000 ;
      RECT  137.175000  0.085000  137.675000 0.595000 ;
      RECT  137.175000  1.445000  140.215000 1.615000 ;
      RECT  137.175000  1.615000  137.505000 2.295000 ;
      RECT  137.175000  2.295000  138.455000 2.465000 ;
      RECT  137.205000  0.765000  137.705000 1.275000 ;
      RECT  137.225000  4.885000  137.495000 5.355000 ;
      RECT  137.235000  2.975000  137.485000 3.815000 ;
      RECT  137.665000  4.715000  137.995000 5.185000 ;
      RECT  137.705000  2.805000  137.955000 3.645000 ;
      RECT  137.725000  1.785000  139.355000 1.980000 ;
      RECT  137.725000  1.980000  137.895000 2.115000 ;
      RECT  137.895000  1.075000  138.395000 1.275000 ;
      RECT  137.950000  0.255000  139.355000 0.505000 ;
      RECT  138.115000  2.195000  138.455000 2.295000 ;
      RECT  138.145000  0.675000  138.395000 1.075000 ;
      RECT  138.165000  4.885000  138.435000 5.355000 ;
      RECT  138.175000  2.975000  138.425000 3.815000 ;
      RECT  138.605000  0.675000  138.815000 1.055000 ;
      RECT  138.605000  1.055000  139.165000 1.275000 ;
      RECT  138.605000  4.715000  138.935000 5.185000 ;
      RECT  138.635000  2.255000  138.990000 2.635000 ;
      RECT  138.645000  2.805000  138.895000 3.645000 ;
      RECT  139.105000  4.885000  139.375000 5.355000 ;
      RECT  139.115000  2.975000  139.365000 3.815000 ;
      RECT  139.175000  0.505000  139.355000 0.655000 ;
      RECT  139.175000  0.655000  140.215000 0.825000 ;
      RECT  139.185000  1.980000  139.355000 2.165000 ;
      RECT  139.345000  0.995000  139.705000 1.275000 ;
      RECT  139.545000  4.715000  139.875000 5.185000 ;
      RECT  139.585000  0.085000  139.915000 0.485000 ;
      RECT  139.585000  2.805000  139.835000 3.645000 ;
      RECT  139.640000  1.855000  139.905000 2.635000 ;
      RECT  139.875000  0.825000  140.215000 1.445000 ;
      RECT  140.045000  4.885000  140.315000 5.355000 ;
      RECT  140.055000  2.975000  144.105000 3.145000 ;
      RECT  140.055000  3.145000  140.305000 3.815000 ;
      RECT  140.385000  0.085000  140.675000 0.810000 ;
      RECT  140.385000  1.470000  140.675000 2.635000 ;
      RECT  140.405000  4.155000  143.795000 4.365000 ;
      RECT  140.485000  4.715000  140.815000 5.185000 ;
      RECT  140.525000  3.315000  140.775000 3.815000 ;
      RECT  140.525000  3.815000  147.875000 3.985000 ;
      RECT  140.855000  0.255000  141.105000 0.680000 ;
      RECT  140.855000  0.680000  142.045000 0.850000 ;
      RECT  140.855000  1.485000  143.120000 1.655000 ;
      RECT  140.855000  1.655000  141.105000 2.465000 ;
      RECT  140.910000  1.075000  141.590000 1.275000 ;
      RECT  140.985000  4.885000  141.255000 5.355000 ;
      RECT  140.995000  3.145000  141.245000 3.645000 ;
      RECT  141.275000  0.085000  141.655000 0.510000 ;
      RECT  141.275000  1.825000  141.575000 2.295000 ;
      RECT  141.275000  2.295000  143.585000 2.465000 ;
      RECT  141.425000  4.715000  141.755000 5.185000 ;
      RECT  141.465000  3.315000  141.715000 3.815000 ;
      RECT  141.745000  1.655000  142.125000 2.125000 ;
      RECT  141.790000  1.075000  142.505000 1.275000 ;
      RECT  141.875000  0.255000  143.065000 0.505000 ;
      RECT  141.875000  0.505000  142.045000 0.680000 ;
      RECT  141.925000  4.885000  142.195000 5.355000 ;
      RECT  141.935000  3.145000  142.185000 3.645000 ;
      RECT  142.215000  0.675000  144.055000 0.845000 ;
      RECT  142.345000  1.825000  142.515000 2.295000 ;
      RECT  142.365000  4.715000  142.695000 5.185000 ;
      RECT  142.405000  3.315000  142.655000 3.815000 ;
      RECT  142.685000  1.655000  143.120000 2.125000 ;
      RECT  142.690000  0.845000  143.120000 1.485000 ;
      RECT  142.865000  4.885000  143.135000 5.355000 ;
      RECT  142.875000  3.145000  143.125000 3.645000 ;
      RECT  143.255000  0.255000  144.545000 0.505000 ;
      RECT  143.305000  4.715000  143.635000 5.185000 ;
      RECT  143.335000  1.485000  145.565000 1.655000 ;
      RECT  143.335000  1.655000  143.585000 2.295000 ;
      RECT  143.345000  3.315000  143.595000 3.815000 ;
      RECT  143.405000  1.075000  144.295000 1.275000 ;
      RECT  143.805000  1.825000  143.975000 2.635000 ;
      RECT  143.805000  4.885000  144.595000 5.355000 ;
      RECT  143.815000  3.145000  144.105000 3.645000 ;
      RECT  144.145000  1.655000  144.625000 2.465000 ;
      RECT  144.295000  2.975000  152.155000 3.145000 ;
      RECT  144.295000  3.145000  144.585000 3.645000 ;
      RECT  144.375000  0.505000  144.545000 0.680000 ;
      RECT  144.375000  0.680000  145.635000 0.850000 ;
      RECT  144.530000  1.075000  145.380000 1.275000 ;
      RECT  144.605000  4.155000  147.995000 4.365000 ;
      RECT  144.740000  0.085000  145.120000 0.510000 ;
      RECT  144.765000  4.715000  145.095000 5.185000 ;
      RECT  144.805000  3.315000  145.055000 3.815000 ;
      RECT  144.845000  1.825000  145.015000 2.635000 ;
      RECT  145.185000  1.655000  145.565000 2.465000 ;
      RECT  145.235000  3.145000  145.525000 3.645000 ;
      RECT  145.265000  4.885000  145.535000 5.355000 ;
      RECT  145.315000  0.255000  145.635000 0.680000 ;
      RECT  145.705000  4.715000  146.035000 5.185000 ;
      RECT  145.745000  3.315000  145.995000 3.815000 ;
      RECT  145.905000  0.085000  146.195000 0.810000 ;
      RECT  145.905000  1.470000  146.195000 2.635000 ;
      RECT  146.205000  4.885000  146.475000 5.355000 ;
      RECT  146.215000  3.145000  146.465000 3.645000 ;
      RECT  146.370000  1.075000  148.375000 1.275000 ;
      RECT  146.370000  1.455000  146.705000 2.295000 ;
      RECT  146.370000  2.295000  150.945000 2.465000 ;
      RECT  146.375000  0.255000  146.705000 0.725000 ;
      RECT  146.375000  0.725000  148.505000 0.905000 ;
      RECT  146.645000  4.715000  146.975000 5.185000 ;
      RECT  146.685000  3.315000  146.935000 3.815000 ;
      RECT  146.925000  0.085000  147.095000 0.555000 ;
      RECT  146.925000  1.445000  149.955000 1.625000 ;
      RECT  146.925000  1.625000  147.135000 2.125000 ;
      RECT  147.145000  4.885000  147.415000 5.355000 ;
      RECT  147.155000  3.145000  147.405000 3.645000 ;
      RECT  147.265000  0.255000  147.645000 0.725000 ;
      RECT  147.355000  1.795000  147.605000 2.295000 ;
      RECT  147.585000  4.715000  147.915000 5.185000 ;
      RECT  147.625000  3.315000  147.875000 3.815000 ;
      RECT  147.825000  1.625000  148.075000 2.125000 ;
      RECT  147.865000  0.085000  148.035000 0.555000 ;
      RECT  148.085000  4.885000  148.355000 5.355000 ;
      RECT  148.095000  3.145000  148.345000 3.985000 ;
      RECT  148.205000  0.255000  150.465000 0.475000 ;
      RECT  148.205000  0.475000  148.505000 0.725000 ;
      RECT  148.295000  1.795000  148.545000 2.295000 ;
      RECT  148.525000  4.715000  148.855000 5.185000 ;
      RECT  148.565000  3.315000  148.815000 3.815000 ;
      RECT  148.565000  3.815000  151.635000 3.985000 ;
      RECT  148.565000  3.985000  148.975000 4.535000 ;
      RECT  148.675000  0.645000  152.395000 0.885000 ;
      RECT  148.675000  0.885000  148.975000 1.445000 ;
      RECT  148.765000  1.625000  149.015000 2.125000 ;
      RECT  149.025000  4.885000  149.295000 5.355000 ;
      RECT  149.035000  3.145000  149.285000 3.645000 ;
      RECT  149.145000  1.075000  150.720000 1.275000 ;
      RECT  149.145000  4.155000  151.515000 4.365000 ;
      RECT  149.235000  1.795000  149.485000 2.295000 ;
      RECT  149.465000  4.715000  149.795000 5.185000 ;
      RECT  149.505000  3.315000  149.755000 3.815000 ;
      RECT  149.705000  1.625000  149.955000 2.125000 ;
      RECT  149.965000  4.885000  150.235000 5.355000 ;
      RECT  149.975000  3.145000  150.225000 3.645000 ;
      RECT  150.175000  1.455000  154.705000 1.625000 ;
      RECT  150.175000  1.625000  150.945000 2.295000 ;
      RECT  150.405000  4.715000  150.735000 5.185000 ;
      RECT  150.445000  3.315000  150.695000 3.815000 ;
      RECT  150.655000  0.255000  152.865000 0.475000 ;
      RECT  150.905000  4.885000  151.175000 5.355000 ;
      RECT  150.915000  3.145000  151.165000 3.645000 ;
      RECT  150.955000  1.075000  152.565000 1.285000 ;
      RECT  151.165000  1.795000  151.415000 2.635000 ;
      RECT  151.345000  4.715000  151.675000 5.185000 ;
      RECT  151.385000  3.315000  151.635000 3.815000 ;
      RECT  151.635000  1.625000  151.885000 2.465000 ;
      RECT  151.845000  4.535000  152.125000 5.355000 ;
      RECT  151.855000  3.145000  152.155000 3.975000 ;
      RECT  152.105000  1.795000  152.355000 2.635000 ;
      RECT  152.345000  2.805000  152.635000 3.970000 ;
      RECT  152.345000  4.630000  152.635000 5.355000 ;
      RECT  152.575000  1.625000  152.825000 2.465000 ;
      RECT  152.615000  0.475000  152.865000 0.725000 ;
      RECT  152.615000  0.725000  154.745000 0.905000 ;
      RECT  152.790000  1.075000  154.815000 1.285000 ;
      RECT  152.815000  2.975000  153.145000 3.825000 ;
      RECT  152.815000  3.825000  154.315000 3.995000 ;
      RECT  152.860000  4.165000  153.960000 4.365000 ;
      RECT  152.865000  4.535000  154.315000 4.705000 ;
      RECT  152.865000  4.705000  153.165000 5.185000 ;
      RECT  153.045000  1.795000  153.295000 2.635000 ;
      RECT  153.085000  0.085000  153.255000 0.555000 ;
      RECT  153.315000  2.805000  153.585000 3.605000 ;
      RECT  153.335000  4.875000  153.615000 5.355000 ;
      RECT  153.425000  0.255000  153.805000 0.725000 ;
      RECT  153.515000  1.625000  153.765000 2.465000 ;
      RECT  153.755000  2.975000  154.085000 3.825000 ;
      RECT  153.785000  4.705000  154.055000 5.185000 ;
      RECT  153.985000  1.795000  154.235000 2.635000 ;
      RECT  154.025000  0.085000  154.195000 0.555000 ;
      RECT  154.140000  3.995000  154.315000 4.195000 ;
      RECT  154.140000  4.195000  156.765000 4.365000 ;
      RECT  154.140000  4.365000  154.315000 4.535000 ;
      RECT  154.225000  4.875000  154.525000 5.355000 ;
      RECT  154.255000  2.805000  154.525000 3.605000 ;
      RECT  154.365000  0.255000  154.745000 0.725000 ;
      RECT  154.455000  1.625000  154.705000 2.465000 ;
      RECT  154.695000  2.975000  155.025000 3.825000 ;
      RECT  154.695000  3.825000  157.845000 3.995000 ;
      RECT  154.695000  4.535000  157.845000 4.705000 ;
      RECT  154.695000  4.705000  155.025000 5.185000 ;
      RECT  155.105000  0.085000  155.395000 0.810000 ;
      RECT  155.105000  1.470000  155.395000 2.635000 ;
      RECT  155.195000  2.805000  155.465000 3.605000 ;
      RECT  155.195000  4.875000  155.465000 5.355000 ;
      RECT  155.565000  0.255000  155.825000 2.465000 ;
      RECT  155.635000  2.975000  155.965000 3.825000 ;
      RECT  155.635000  4.705000  155.965000 5.185000 ;
      RECT  155.995000  0.085000  156.475000 0.530000 ;
      RECT  155.995000  0.995000  156.165000 1.805000 ;
      RECT  155.995000  1.805000  156.855000 1.975000 ;
      RECT  155.995000  2.235000  156.375000 2.635000 ;
      RECT  156.135000  2.805000  156.405000 3.605000 ;
      RECT  156.135000  4.875000  156.405000 5.355000 ;
      RECT  156.425000  0.995000  156.805000 1.615000 ;
      RECT  156.575000  2.975000  156.905000 3.825000 ;
      RECT  156.575000  4.705000  156.905000 5.185000 ;
      RECT  156.635000  1.975000  156.855000 2.200000 ;
      RECT  156.635000  2.200000  157.865000 2.370000 ;
      RECT  156.745000  0.255000  156.915000 0.655000 ;
      RECT  156.745000  0.655000  157.690000 0.825000 ;
      RECT  156.975000  0.995000  157.210000 1.375000 ;
      RECT  157.010000  3.995000  157.845000 4.535000 ;
      RECT  157.075000  2.805000  157.345000 3.605000 ;
      RECT  157.075000  4.875000  157.345000 5.355000 ;
      RECT  157.150000  0.085000  157.870000 0.485000 ;
      RECT  157.170000  1.545000  157.690000 1.715000 ;
      RECT  157.170000  1.715000  157.340000 1.905000 ;
      RECT  157.515000  2.975000  157.845000 3.825000 ;
      RECT  157.515000  4.705000  157.845000 5.185000 ;
      RECT  157.520000  0.825000  157.690000 1.545000 ;
      RECT  157.610000  1.895000  158.080000 2.065000 ;
      RECT  157.610000  2.065000  157.865000 2.200000 ;
      RECT  157.610000  2.370000  157.865000 2.465000 ;
      RECT  157.860000  0.700000  158.335000 0.870000 ;
      RECT  157.860000  0.870000  158.080000 1.895000 ;
      RECT  158.015000  2.805000  158.315000 3.955000 ;
      RECT  158.015000  4.555000  158.265000 5.355000 ;
      RECT  158.085000  2.255000  158.425000 2.425000 ;
      RECT  158.165000  0.255000  158.335000 0.700000 ;
      RECT  158.255000  1.835000  159.295000 2.005000 ;
      RECT  158.255000  2.005000  158.425000 2.255000 ;
      RECT  158.375000  1.040000  158.635000 1.655000 ;
      RECT  158.635000  2.175000  158.895000 2.635000 ;
      RECT  158.785000  2.805000  159.075000 3.970000 ;
      RECT  158.785000  4.630000  159.075000 5.355000 ;
      RECT  158.845000  0.765000  159.105000 1.655000 ;
      RECT  158.970000  0.085000  159.420000 0.595000 ;
      RECT  159.115000  2.005000  159.295000 2.465000 ;
      RECT  159.250000  2.975000  159.575000 3.775000 ;
      RECT  159.250000  3.775000  160.515000 3.985000 ;
      RECT  159.305000  4.535000  159.575000 5.355000 ;
      RECT  159.575000  4.165000  160.245000 4.365000 ;
      RECT  159.705000  0.085000  159.995000 0.810000 ;
      RECT  159.705000  1.470000  159.995000 2.635000 ;
      RECT  159.745000  2.805000  160.075000 3.605000 ;
      RECT  159.745000  4.535000  161.535000 4.705000 ;
      RECT  159.745000  4.705000  161.015000 4.715000 ;
      RECT  159.745000  4.715000  160.075000 5.185000 ;
      RECT  160.245000  2.975000  161.485000 3.145000 ;
      RECT  160.245000  3.145000  160.515000 3.775000 ;
      RECT  160.245000  4.885000  160.515000 5.355000 ;
      RECT  160.265000  0.085000  160.435000 0.930000 ;
      RECT  160.265000  1.445000  160.435000 2.635000 ;
      RECT  160.515000  4.165000  161.185000 4.365000 ;
      RECT  160.605000  0.255000  160.910000 0.810000 ;
      RECT  160.605000  0.810000  160.825000 1.525000 ;
      RECT  160.605000  1.525000  160.910000 2.465000 ;
      RECT  160.685000  3.315000  161.015000 3.775000 ;
      RECT  160.685000  3.775000  161.535000 3.995000 ;
      RECT  160.685000  4.715000  161.015000 5.185000 ;
      RECT  160.995000  0.995000  161.300000 1.325000 ;
      RECT  161.080000  0.085000  161.560000 0.530000 ;
      RECT  161.080000  1.325000  161.300000 1.805000 ;
      RECT  161.080000  1.805000  161.940000 1.975000 ;
      RECT  161.080000  2.235000  161.460000 2.635000 ;
      RECT  161.185000  3.145000  161.485000 3.605000 ;
      RECT  161.185000  4.885000  161.975000 5.355000 ;
      RECT  161.355000  3.995000  161.535000 4.165000 ;
      RECT  161.355000  4.165000  164.685000 4.365000 ;
      RECT  161.355000  4.365000  161.535000 4.535000 ;
      RECT  161.525000  0.995000  161.895000 1.615000 ;
      RECT  161.705000  2.805000  161.975000 3.945000 ;
      RECT  161.705000  4.535000  161.975000 4.885000 ;
      RECT  161.720000  1.975000  161.940000 2.200000 ;
      RECT  161.720000  2.200000  162.950000 2.370000 ;
      RECT  161.845000  0.255000  162.015000 0.655000 ;
      RECT  161.845000  0.655000  162.790000 0.825000 ;
      RECT  162.065000  0.995000  162.415000 1.375000 ;
      RECT  162.145000  2.975000  162.475000 3.775000 ;
      RECT  162.145000  3.775000  165.495000 3.945000 ;
      RECT  162.145000  4.535000  165.495000 4.715000 ;
      RECT  162.145000  4.715000  162.445000 5.185000 ;
      RECT  162.235000  0.085000  162.970000 0.485000 ;
      RECT  162.255000  1.545000  162.790000 1.715000 ;
      RECT  162.255000  1.715000  162.425000 1.905000 ;
      RECT  162.615000  4.885000  162.945000 5.355000 ;
      RECT  162.620000  0.825000  162.790000 1.545000 ;
      RECT  162.645000  2.805000  162.915000 3.605000 ;
      RECT  162.720000  1.895000  163.180000 2.065000 ;
      RECT  162.720000  2.065000  162.950000 2.200000 ;
      RECT  162.780000  2.370000  162.950000 2.465000 ;
      RECT  162.960000  0.700000  163.360000 0.870000 ;
      RECT  162.960000  0.870000  163.180000 1.895000 ;
      RECT  163.085000  2.975000  163.415000 3.775000 ;
      RECT  163.115000  4.715000  163.385000 5.185000 ;
      RECT  163.190000  0.255000  163.360000 0.700000 ;
      RECT  163.205000  2.255000  163.535000 2.425000 ;
      RECT  163.365000  1.835000  164.395000 2.005000 ;
      RECT  163.365000  2.005000  163.535000 2.255000 ;
      RECT  163.380000  1.050000  163.840000 1.655000 ;
      RECT  163.555000  4.885000  163.885000 5.355000 ;
      RECT  163.585000  2.805000  163.855000 3.605000 ;
      RECT  163.755000  2.175000  164.005000 2.635000 ;
      RECT  163.985000  0.085000  164.435000 0.595000 ;
      RECT  164.025000  2.975000  164.355000 3.775000 ;
      RECT  164.055000  4.715000  164.325000 5.185000 ;
      RECT  164.160000  0.765000  164.535000 1.655000 ;
      RECT  164.225000  2.005000  164.395000 2.465000 ;
      RECT  164.495000  4.885000  164.825000 5.355000 ;
      RECT  164.525000  2.805000  164.795000 3.605000 ;
      RECT  164.765000  0.085000  165.055000 0.810000 ;
      RECT  164.765000  1.470000  165.055000 2.635000 ;
      RECT  164.965000  2.975000  165.295000 3.775000 ;
      RECT  164.995000  4.715000  165.265000 5.185000 ;
      RECT  165.095000  3.945000  165.495000 4.535000 ;
      RECT  165.225000  1.075000  165.765000 1.445000 ;
      RECT  165.225000  1.445000  166.975000 1.615000 ;
      RECT  165.275000  1.785000  167.405000 1.955000 ;
      RECT  165.275000  1.955000  165.525000 2.465000 ;
      RECT  165.315000  0.085000  165.485000 0.895000 ;
      RECT  165.435000  4.885000  165.765000 5.355000 ;
      RECT  165.465000  2.805000  165.735000 3.605000 ;
      RECT  165.655000  0.255000  166.975000 0.475000 ;
      RECT  165.655000  0.475000  165.955000 0.905000 ;
      RECT  165.745000  2.125000  165.995000 2.635000 ;
      RECT  165.995000  1.075000  166.585000 1.275000 ;
      RECT  166.125000  0.645000  166.510000 0.735000 ;
      RECT  166.125000  0.735000  167.915000 0.905000 ;
      RECT  166.145000  2.985000  166.435000 3.970000 ;
      RECT  166.145000  4.630000  166.435000 5.355000 ;
      RECT  166.215000  1.955000  166.465000 2.465000 ;
      RECT  166.605000  2.985000  166.895000 3.970000 ;
      RECT  166.605000  4.630000  166.895000 5.355000 ;
      RECT  166.685000  2.125000  166.935000 2.635000 ;
      RECT  166.805000  1.075000  167.235000 1.245000 ;
      RECT  166.805000  1.245000  166.975000 1.445000 ;
      RECT  167.070000  2.975000  167.395000 3.775000 ;
      RECT  167.070000  3.775000  168.335000 3.985000 ;
      RECT  167.125000  4.535000  167.395000 5.355000 ;
      RECT  167.155000  1.955000  167.405000 2.295000 ;
      RECT  167.155000  2.295000  168.345000 2.465000 ;
      RECT  167.195000  0.085000  167.365000 0.555000 ;
      RECT  167.195000  1.455000  167.405000 1.785000 ;
      RECT  167.395000  4.165000  168.065000 4.365000 ;
      RECT  167.535000  0.255000  167.915000 0.735000 ;
      RECT  167.565000  2.805000  167.895000 3.605000 ;
      RECT  167.565000  4.535000  169.355000 4.705000 ;
      RECT  167.565000  4.705000  168.835000 4.715000 ;
      RECT  167.565000  4.715000  167.895000 5.185000 ;
      RECT  167.625000  0.905000  167.835000 1.415000 ;
      RECT  167.625000  1.415000  168.010000 1.965000 ;
      RECT  167.625000  1.965000  167.875000 2.125000 ;
      RECT  168.005000  1.075000  168.585000 1.245000 ;
      RECT  168.065000  2.975000  169.305000 3.145000 ;
      RECT  168.065000  3.145000  168.335000 3.775000 ;
      RECT  168.065000  4.885000  168.335000 5.355000 ;
      RECT  168.095000  2.135000  168.345000 2.295000 ;
      RECT  168.135000  0.085000  168.825000 0.555000 ;
      RECT  168.335000  4.165000  169.005000 4.365000 ;
      RECT  168.395000  0.725000  170.315000 0.905000 ;
      RECT  168.395000  0.905000  168.585000 1.075000 ;
      RECT  168.395000  1.245000  168.585000 1.495000 ;
      RECT  168.395000  1.495000  168.745000 1.665000 ;
      RECT  168.505000  3.315000  168.835000 3.775000 ;
      RECT  168.505000  3.775000  169.355000 3.995000 ;
      RECT  168.505000  4.715000  168.835000 5.185000 ;
      RECT  168.575000  1.665000  168.745000 1.785000 ;
      RECT  168.575000  1.785000  169.805000 1.965000 ;
      RECT  168.615000  2.135000  168.865000 2.635000 ;
      RECT  168.755000  1.075000  169.145000 1.325000 ;
      RECT  168.915000  1.325000  169.145000 1.445000 ;
      RECT  168.915000  1.445000  170.605000 1.615000 ;
      RECT  168.995000  0.255000  169.375000 0.725000 ;
      RECT  169.005000  3.145000  169.305000 3.605000 ;
      RECT  169.005000  4.885000  169.795000 5.355000 ;
      RECT  169.085000  2.135000  169.335000 2.295000 ;
      RECT  169.085000  2.295000  170.275000 2.465000 ;
      RECT  169.175000  3.995000  169.355000 4.165000 ;
      RECT  169.175000  4.165000  171.825000 4.365000 ;
      RECT  169.175000  4.365000  169.355000 4.535000 ;
      RECT  169.345000  1.075000  170.055000 1.275000 ;
      RECT  169.525000  2.805000  169.795000 3.945000 ;
      RECT  169.525000  4.535000  169.795000 4.885000 ;
      RECT  169.555000  1.965000  169.805000 2.125000 ;
      RECT  169.595000  0.085000  169.765000 0.555000 ;
      RECT  169.935000  0.255000  170.315000 0.725000 ;
      RECT  169.965000  2.975000  170.295000 3.775000 ;
      RECT  169.965000  3.775000  172.395000 3.945000 ;
      RECT  169.965000  4.535000  172.395000 4.715000 ;
      RECT  169.965000  4.715000  170.265000 5.185000 ;
      RECT  170.025000  1.785000  170.275000 2.295000 ;
      RECT  170.225000  1.075000  170.605000 1.445000 ;
      RECT  170.435000  4.885000  170.765000 5.355000 ;
      RECT  170.465000  2.805000  170.735000 3.605000 ;
      RECT  170.495000  1.795000  170.745000 2.635000 ;
      RECT  170.535000  0.085000  170.705000 0.895000 ;
      RECT  170.775000  1.075000  172.230000 1.245000 ;
      RECT  170.775000  1.245000  171.150000 1.615000 ;
      RECT  170.875000  0.275000  171.255000 0.725000 ;
      RECT  170.875000  0.725000  172.815000 0.905000 ;
      RECT  170.905000  2.975000  171.235000 3.775000 ;
      RECT  170.935000  4.715000  171.205000 5.185000 ;
      RECT  170.965000  1.785000  172.155000 1.955000 ;
      RECT  170.965000  1.955000  171.215000 2.465000 ;
      RECT  171.375000  4.885000  171.705000 5.355000 ;
      RECT  171.405000  2.805000  171.675000 3.605000 ;
      RECT  171.435000  2.165000  171.685000 2.635000 ;
      RECT  171.475000  0.085000  171.645000 0.555000 ;
      RECT  171.815000  0.275000  172.195000 0.725000 ;
      RECT  171.845000  2.975000  172.175000 3.775000 ;
      RECT  171.875000  4.715000  172.145000 5.185000 ;
      RECT  171.905000  1.415000  172.815000 1.655000 ;
      RECT  171.905000  1.655000  172.155000 1.785000 ;
      RECT  171.905000  1.955000  172.155000 2.465000 ;
      RECT  171.995000  3.945000  172.395000 4.535000 ;
      RECT  172.315000  4.885000  172.645000 5.355000 ;
      RECT  172.345000  2.805000  172.615000 3.605000 ;
      RECT  172.375000  1.825000  172.625000 2.635000 ;
      RECT  172.415000  0.085000  172.585000 0.555000 ;
      RECT  172.450000  0.905000  172.815000 1.415000 ;
      RECT  173.045000  0.085000  173.335000 0.810000 ;
      RECT  173.045000  1.470000  173.335000 2.635000 ;
      RECT  173.045000  2.805000  173.335000 3.970000 ;
      RECT  173.045000  4.630000  173.335000 5.355000 ;
      RECT  173.515000  0.085000  173.845000 0.825000 ;
      RECT  173.515000  1.805000  173.845000 2.635000 ;
      RECT  173.515000  2.975000  173.845000 3.825000 ;
      RECT  173.515000  3.825000  175.015000 3.995000 ;
      RECT  173.560000  4.165000  174.660000 4.365000 ;
      RECT  173.565000  4.535000  175.015000 4.705000 ;
      RECT  173.565000  4.705000  173.865000 5.185000 ;
      RECT  173.570000  0.995000  173.940000 1.615000 ;
      RECT  174.015000  2.805000  174.285000 3.605000 ;
      RECT  174.035000  4.875000  174.315000 5.355000 ;
      RECT  174.065000  0.255000  174.235000 0.660000 ;
      RECT  174.065000  0.660000  175.235000 0.830000 ;
      RECT  174.195000  1.010000  174.760000 1.275000 ;
      RECT  174.345000  1.445000  175.235000 1.615000 ;
      RECT  174.345000  1.615000  174.725000 2.465000 ;
      RECT  174.455000  2.975000  174.785000 3.825000 ;
      RECT  174.465000  0.085000  175.135000 0.490000 ;
      RECT  174.485000  4.705000  174.755000 5.185000 ;
      RECT  174.840000  3.995000  175.015000 4.195000 ;
      RECT  174.840000  4.195000  177.465000 4.365000 ;
      RECT  174.840000  4.365000  175.015000 4.535000 ;
      RECT  174.925000  4.875000  175.225000 5.355000 ;
      RECT  174.940000  1.785000  175.575000 1.955000 ;
      RECT  174.940000  1.955000  175.305000 2.465000 ;
      RECT  174.955000  2.805000  175.225000 3.605000 ;
      RECT  175.065000  0.830000  175.235000 1.445000 ;
      RECT  175.395000  2.975000  175.725000 3.825000 ;
      RECT  175.395000  3.825000  178.545000 3.995000 ;
      RECT  175.395000  4.535000  178.545000 4.705000 ;
      RECT  175.395000  4.705000  175.725000 5.185000 ;
      RECT  175.405000  0.255000  175.695000 0.825000 ;
      RECT  175.405000  0.825000  175.575000 1.785000 ;
      RECT  175.475000  2.235000  175.915000 2.465000 ;
      RECT  175.745000  1.785000  176.810000 1.955000 ;
      RECT  175.745000  1.955000  175.915000 2.235000 ;
      RECT  175.805000  0.995000  176.035000 1.615000 ;
      RECT  175.865000  0.425000  176.035000 0.995000 ;
      RECT  175.895000  2.805000  176.165000 3.605000 ;
      RECT  175.895000  4.875000  176.165000 5.355000 ;
      RECT  176.085000  2.135000  176.335000 2.635000 ;
      RECT  176.305000  0.995000  176.645000 1.615000 ;
      RECT  176.335000  2.975000  176.665000 3.825000 ;
      RECT  176.335000  4.705000  176.665000 5.185000 ;
      RECT  176.425000  0.085000  176.805000 0.825000 ;
      RECT  176.555000  1.955000  176.810000 2.465000 ;
      RECT  176.835000  2.805000  177.105000 3.605000 ;
      RECT  176.835000  4.875000  177.105000 5.355000 ;
      RECT  177.185000  0.085000  177.475000 0.810000 ;
      RECT  177.185000  1.470000  177.475000 2.635000 ;
      RECT  177.275000  2.975000  177.605000 3.825000 ;
      RECT  177.275000  4.705000  177.605000 5.185000 ;
      RECT  177.670000  1.075000  178.200000 1.445000 ;
      RECT  177.670000  1.445000  179.655000 1.615000 ;
      RECT  177.695000  1.785000  179.825000 1.955000 ;
      RECT  177.695000  1.955000  177.945000 2.465000 ;
      RECT  177.710000  3.995000  178.545000 4.535000 ;
      RECT  177.735000  0.085000  177.905000 0.895000 ;
      RECT  177.775000  2.805000  178.045000 3.605000 ;
      RECT  177.775000  4.875000  178.045000 5.355000 ;
      RECT  178.075000  0.255000  179.395000 0.475000 ;
      RECT  178.075000  0.475000  178.375000 0.895000 ;
      RECT  178.165000  2.135000  178.415000 2.635000 ;
      RECT  178.215000  2.975000  178.545000 3.825000 ;
      RECT  178.215000  4.705000  178.545000 5.185000 ;
      RECT  178.415000  1.075000  179.005000 1.275000 ;
      RECT  178.545000  0.645000  178.925000 0.725000 ;
      RECT  178.545000  0.725000  180.335000 0.905000 ;
      RECT  178.635000  1.955000  178.885000 2.465000 ;
      RECT  178.715000  2.805000  179.015000 3.955000 ;
      RECT  178.715000  4.555000  178.965000 5.355000 ;
      RECT  179.105000  2.135000  179.355000 2.635000 ;
      RECT  179.275000  1.075000  179.655000 1.445000 ;
      RECT  179.485000  2.805000  179.775000 3.970000 ;
      RECT  179.485000  4.630000  179.775000 5.355000 ;
      RECT  179.575000  1.955000  179.825000 2.295000 ;
      RECT  179.575000  2.295000  180.765000 2.465000 ;
      RECT  179.615000  0.085000  179.785000 0.555000 ;
      RECT  179.945000  2.975000  180.255000 3.475000 ;
      RECT  179.945000  3.475000  180.755000 3.645000 ;
      RECT  179.945000  3.815000  180.295000 4.455000 ;
      RECT  179.955000  0.255000  180.335000 0.725000 ;
      RECT  180.005000  0.905000  180.335000 2.125000 ;
      RECT  180.085000  4.635000  180.635000 4.805000 ;
      RECT  180.085000  4.805000  180.255000 5.160000 ;
      RECT  180.425000  2.805000  180.755000 3.305000 ;
      RECT  180.425000  4.975000  180.755000 5.355000 ;
      RECT  180.465000  3.645000  180.755000 4.370000 ;
      RECT  180.465000  4.370000  180.635000 4.635000 ;
      RECT  180.515000  1.795000  180.765000 2.295000 ;
      RECT  180.555000  0.085000  181.245000 0.555000 ;
      RECT  180.555000  0.995000  180.845000 1.325000 ;
      RECT  180.675000  0.725000  182.735000 0.905000 ;
      RECT  180.675000  0.905000  180.845000 0.995000 ;
      RECT  180.675000  1.325000  180.845000 1.445000 ;
      RECT  180.675000  1.445000  182.695000 1.615000 ;
      RECT  180.925000  2.975000  181.195000 3.995000 ;
      RECT  180.925000  3.995000  181.095000 5.160000 ;
      RECT  181.035000  1.075000  182.030000 1.275000 ;
      RECT  181.035000  1.785000  182.225000 1.965000 ;
      RECT  181.035000  1.965000  181.285000 2.465000 ;
      RECT  181.295000  4.140000  181.625000 4.485000 ;
      RECT  181.415000  0.255000  181.795000 0.725000 ;
      RECT  181.415000  2.975000  181.745000 3.775000 ;
      RECT  181.415000  3.775000  181.975000 3.945000 ;
      RECT  181.505000  2.135000  181.755000 2.635000 ;
      RECT  181.520000  4.655000  182.395000 4.675000 ;
      RECT  181.520000  4.675000  181.975000 4.825000 ;
      RECT  181.520000  4.825000  181.715000 5.095000 ;
      RECT  181.805000  3.945000  181.975000 4.345000 ;
      RECT  181.805000  4.345000  182.395000 4.655000 ;
      RECT  181.885000  4.995000  182.215000 5.355000 ;
      RECT  181.915000  2.805000  182.185000 3.605000 ;
      RECT  181.975000  1.965000  182.225000 2.295000 ;
      RECT  181.975000  2.295000  183.165000 2.465000 ;
      RECT  182.015000  0.085000  182.185000 0.555000 ;
      RECT  182.280000  1.075000  182.995000 1.275000 ;
      RECT  182.305000  3.755000  182.815000 4.175000 ;
      RECT  182.355000  0.255000  182.735000 0.725000 ;
      RECT  182.445000  1.615000  182.695000 2.125000 ;
      RECT  182.640000  4.345000  183.155000 4.705000 ;
      RECT  182.880000  3.055000  183.710000 3.275000 ;
      RECT  182.900000  4.875000  183.520000 5.160000 ;
      RECT  182.915000  1.455000  183.165000 2.295000 ;
      RECT  182.955000  0.085000  183.125000 0.905000 ;
      RECT  182.985000  3.445000  183.370000 3.865000 ;
      RECT  182.985000  3.865000  183.155000 4.345000 ;
      RECT  183.350000  4.275000  184.240000 4.445000 ;
      RECT  183.350000  4.445000  183.520000 4.875000 ;
      RECT  183.540000  3.275000  183.710000 4.115000 ;
      RECT  183.540000  4.115000  184.240000 4.275000 ;
      RECT  183.625000  0.085000  183.915000 0.810000 ;
      RECT  183.625000  1.470000  183.915000 2.635000 ;
      RECT  183.730000  4.830000  184.060000 5.355000 ;
      RECT  183.880000  3.575000  185.030000 3.735000 ;
      RECT  183.880000  3.735000  185.585000 3.905000 ;
      RECT  183.910000  2.805000  184.495000 3.305000 ;
      RECT  184.085000  1.455000  185.315000 1.625000 ;
      RECT  184.085000  1.625000  184.425000 2.465000 ;
      RECT  184.100000  1.075000  185.705000 1.285000 ;
      RECT  184.175000  0.085000  184.345000 0.895000 ;
      RECT  184.315000  4.615000  184.645000 5.185000 ;
      RECT  184.410000  3.905000  184.580000 4.615000 ;
      RECT  184.515000  0.255000  184.895000 0.725000 ;
      RECT  184.515000  0.725000  185.755000 0.905000 ;
      RECT  184.645000  1.795000  184.855000 2.635000 ;
      RECT  184.745000  2.975000  185.030000 3.575000 ;
      RECT  184.750000  4.115000  185.245000 4.445000 ;
      RECT  185.075000  1.625000  185.315000 1.795000 ;
      RECT  185.075000  1.795000  188.145000 1.965000 ;
      RECT  185.075000  1.965000  185.315000 2.465000 ;
      RECT  185.115000  0.085000  185.285000 0.555000 ;
      RECT  185.180000  4.615000  185.510000 4.815000 ;
      RECT  185.180000  4.815000  185.455000 5.355000 ;
      RECT  185.205000  2.805000  185.505000 3.290000 ;
      RECT  185.205000  3.290000  185.535000 3.555000 ;
      RECT  185.415000  3.905000  185.585000 4.115000 ;
      RECT  185.415000  4.115000  185.755000 4.385000 ;
      RECT  185.455000  0.255000  187.715000 0.475000 ;
      RECT  185.455000  0.475000  185.755000 0.725000 ;
      RECT  185.535000  1.285000  185.705000 1.445000 ;
      RECT  185.535000  1.445000  187.975000 1.615000 ;
      RECT  185.545000  2.135000  185.795000 2.635000 ;
      RECT  185.625000  4.945000  186.155000 5.185000 ;
      RECT  185.675000  2.975000  186.155000 3.185000 ;
      RECT  185.680000  4.555000  186.155000 4.945000 ;
      RECT  185.755000  3.185000  186.155000 3.945000 ;
      RECT  185.875000  1.075000  187.425000 1.275000 ;
      RECT  185.925000  0.645000  187.295000 0.725000 ;
      RECT  185.925000  0.725000  189.595000 0.905000 ;
      RECT  185.925000  3.945000  186.155000 4.555000 ;
      RECT  186.015000  1.965000  186.265000 2.465000 ;
      RECT  186.385000  2.805000  186.675000 3.970000 ;
      RECT  186.385000  4.630000  186.675000 5.355000 ;
      RECT  186.485000  2.135000  186.735000 2.635000 ;
      RECT  186.845000  2.975000  187.155000 3.475000 ;
      RECT  186.845000  3.475000  187.535000 3.645000 ;
      RECT  186.845000  3.815000  187.195000 4.455000 ;
      RECT  186.955000  1.965000  187.205000 2.465000 ;
      RECT  186.985000  4.635000  187.535000 4.805000 ;
      RECT  186.985000  4.805000  187.155000 5.160000 ;
      RECT  187.325000  2.805000  187.655000 3.305000 ;
      RECT  187.325000  4.975000  187.655000 5.355000 ;
      RECT  187.365000  3.645000  187.535000 4.040000 ;
      RECT  187.365000  4.040000  187.655000 4.370000 ;
      RECT  187.365000  4.370000  187.535000 4.635000 ;
      RECT  187.425000  2.135000  187.675000 2.635000 ;
      RECT  187.595000  1.075000  187.975000 1.445000 ;
      RECT  187.825000  2.975000  188.095000 3.755000 ;
      RECT  187.825000  3.755000  187.995000 5.160000 ;
      RECT  187.895000  1.965000  188.145000 2.295000 ;
      RECT  187.895000  2.295000  190.065000 2.465000 ;
      RECT  187.935000  0.085000  188.105000 0.555000 ;
      RECT  188.145000  0.905000  188.365000 1.415000 ;
      RECT  188.145000  1.415000  189.515000 1.615000 ;
      RECT  188.195000  4.115000  188.525000 4.485000 ;
      RECT  188.275000  0.275000  188.655000 0.725000 ;
      RECT  188.315000  2.975000  188.645000 3.775000 ;
      RECT  188.315000  3.775000  188.875000 3.945000 ;
      RECT  188.365000  1.615000  188.615000 2.125000 ;
      RECT  188.420000  4.655000  189.295000 4.675000 ;
      RECT  188.420000  4.675000  188.875000 4.825000 ;
      RECT  188.420000  4.825000  188.615000 5.095000 ;
      RECT  188.535000  1.075000  190.325000 1.245000 ;
      RECT  188.705000  3.945000  188.875000 4.345000 ;
      RECT  188.705000  4.345000  189.295000 4.655000 ;
      RECT  188.785000  4.995000  189.115000 5.355000 ;
      RECT  188.815000  2.805000  189.085000 3.605000 ;
      RECT  188.835000  1.795000  189.075000 2.295000 ;
      RECT  188.875000  0.085000  189.045000 0.555000 ;
      RECT  189.205000  3.755000  189.715000 4.175000 ;
      RECT  189.215000  0.275000  189.595000 0.725000 ;
      RECT  189.245000  1.615000  189.515000 2.125000 ;
      RECT  189.540000  4.345000  190.055000 4.705000 ;
      RECT  189.685000  1.455000  190.065000 2.295000 ;
      RECT  189.780000  3.055000  190.610000 3.275000 ;
      RECT  189.800000  4.875000  190.420000 5.160000 ;
      RECT  189.815000  0.085000  190.505000 0.555000 ;
      RECT  189.885000  3.445000  190.270000 3.865000 ;
      RECT  189.885000  3.865000  190.055000 4.345000 ;
      RECT  190.155000  0.735000  194.460000 0.905000 ;
      RECT  190.155000  0.905000  190.325000 1.075000 ;
      RECT  190.250000  4.275000  191.140000 4.445000 ;
      RECT  190.250000  4.445000  190.420000 4.875000 ;
      RECT  190.255000  1.455000  192.425000 1.625000 ;
      RECT  190.255000  1.625000  190.585000 2.465000 ;
      RECT  190.440000  3.275000  190.610000 4.115000 ;
      RECT  190.440000  4.115000  191.140000 4.275000 ;
      RECT  190.545000  1.075000  192.070000 1.275000 ;
      RECT  190.630000  4.830000  190.960000 5.355000 ;
      RECT  190.675000  0.255000  191.055000 0.725000 ;
      RECT  190.675000  0.725000  193.875000 0.735000 ;
      RECT  190.780000  3.575000  191.930000 3.735000 ;
      RECT  190.780000  3.735000  192.485000 3.905000 ;
      RECT  190.805000  1.795000  191.015000 2.635000 ;
      RECT  190.810000  2.805000  191.395000 3.305000 ;
      RECT  191.215000  4.615000  191.545000 5.185000 ;
      RECT  191.240000  1.625000  191.480000 2.465000 ;
      RECT  191.275000  0.085000  191.445000 0.555000 ;
      RECT  191.310000  3.905000  191.480000 4.615000 ;
      RECT  191.615000  0.255000  191.995000 0.725000 ;
      RECT  191.645000  2.975000  191.930000 3.575000 ;
      RECT  191.650000  4.115000  192.145000 4.445000 ;
      RECT  191.705000  1.795000  191.955000 2.635000 ;
      RECT  192.080000  4.615000  192.410000 4.815000 ;
      RECT  192.080000  4.815000  192.355000 5.355000 ;
      RECT  192.105000  2.805000  192.405000 3.290000 ;
      RECT  192.105000  3.290000  192.435000 3.555000 ;
      RECT  192.175000  1.625000  192.425000 2.295000 ;
      RECT  192.175000  2.295000  194.310000 2.465000 ;
      RECT  192.215000  0.085000  192.385000 0.555000 ;
      RECT  192.315000  3.905000  192.485000 4.115000 ;
      RECT  192.315000  4.115000  192.655000 4.385000 ;
      RECT  192.440000  1.075000  193.965000 1.275000 ;
      RECT  192.525000  4.945000  193.055000 5.185000 ;
      RECT  192.555000  0.255000  192.935000 0.725000 ;
      RECT  192.575000  2.975000  193.055000 3.185000 ;
      RECT  192.580000  4.555000  193.055000 4.945000 ;
      RECT  192.645000  1.455000  194.460000 1.625000 ;
      RECT  192.645000  1.625000  192.895000 2.125000 ;
      RECT  192.655000  3.185000  193.055000 3.945000 ;
      RECT  192.825000  3.945000  193.055000 4.555000 ;
      RECT  193.115000  1.795000  193.365000 2.295000 ;
      RECT  193.155000  0.085000  193.325000 0.555000 ;
      RECT  193.285000  2.805000  193.575000 3.970000 ;
      RECT  193.285000  4.630000  193.575000 5.355000 ;
      RECT  193.495000  0.255000  193.875000 0.725000 ;
      RECT  193.585000  1.625000  193.835000 2.125000 ;
      RECT  193.745000  2.975000  194.055000 3.475000 ;
      RECT  193.745000  3.475000  194.555000 3.645000 ;
      RECT  193.745000  3.815000  194.095000 4.455000 ;
      RECT  193.885000  4.635000  194.435000 4.805000 ;
      RECT  193.885000  4.805000  194.055000 5.160000 ;
      RECT  194.060000  1.795000  194.310000 2.295000 ;
      RECT  194.095000  0.085000  194.265000 0.555000 ;
      RECT  194.135000  0.905000  194.460000 1.455000 ;
      RECT  194.225000  2.805000  194.555000 3.305000 ;
      RECT  194.225000  4.975000  194.555000 5.355000 ;
      RECT  194.265000  3.645000  194.555000 4.370000 ;
      RECT  194.265000  4.370000  194.435000 4.635000 ;
      RECT  194.665000  0.085000  194.955000 0.810000 ;
      RECT  194.665000  1.470000  194.955000 2.635000 ;
      RECT  194.725000  2.975000  194.995000 3.995000 ;
      RECT  194.725000  3.995000  194.895000 5.160000 ;
      RECT  195.095000  4.140000  195.425000 4.485000 ;
      RECT  195.135000  0.300000  195.465000 0.810000 ;
      RECT  195.135000  0.810000  195.325000 1.575000 ;
      RECT  195.135000  1.575000  195.465000 2.425000 ;
      RECT  195.215000  2.975000  195.545000 3.775000 ;
      RECT  195.215000  3.775000  195.775000 3.945000 ;
      RECT  195.320000  4.655000  196.195000 4.675000 ;
      RECT  195.320000  4.675000  195.775000 4.825000 ;
      RECT  195.320000  4.825000  195.515000 5.095000 ;
      RECT  195.495000  0.995000  195.855000 1.325000 ;
      RECT  195.605000  3.945000  195.775000 4.345000 ;
      RECT  195.605000  4.345000  196.195000 4.655000 ;
      RECT  195.645000  0.085000  195.975000 0.485000 ;
      RECT  195.685000  0.655000  198.125000 0.825000 ;
      RECT  195.685000  0.825000  195.855000 0.995000 ;
      RECT  195.685000  1.495000  195.935000 2.635000 ;
      RECT  195.685000  4.995000  196.015000 5.355000 ;
      RECT  195.715000  2.805000  195.985000 3.605000 ;
      RECT  196.025000  0.995000  196.380000 1.325000 ;
      RECT  196.105000  3.755000  196.615000 4.175000 ;
      RECT  196.115000  1.325000  196.380000 1.655000 ;
      RECT  196.125000  1.825000  197.565000 1.995000 ;
      RECT  196.125000  1.995000  196.425000 2.415000 ;
      RECT  196.440000  4.345000  196.955000 4.705000 ;
      RECT  196.555000  0.995000  196.855000 1.655000 ;
      RECT  196.680000  3.055000  197.510000 3.275000 ;
      RECT  196.700000  4.875000  197.320000 5.160000 ;
      RECT  196.705000  2.165000  197.035000 2.635000 ;
      RECT  196.785000  3.445000  197.170000 3.865000 ;
      RECT  196.785000  3.865000  196.955000 4.345000 ;
      RECT  197.025000  0.995000  197.315000 1.655000 ;
      RECT  197.150000  4.275000  198.040000 4.445000 ;
      RECT  197.150000  4.445000  197.320000 4.875000 ;
      RECT  197.165000  0.315000  197.545000 0.655000 ;
      RECT  197.315000  1.995000  197.565000 2.415000 ;
      RECT  197.340000  3.275000  197.510000 4.115000 ;
      RECT  197.340000  4.115000  198.040000 4.275000 ;
      RECT  197.485000  0.995000  197.785000 1.655000 ;
      RECT  197.530000  4.830000  197.860000 5.355000 ;
      RECT  197.680000  3.575000  198.830000 3.735000 ;
      RECT  197.680000  3.735000  199.385000 3.905000 ;
      RECT  197.710000  2.805000  198.295000 3.305000 ;
      RECT  197.765000  0.085000  198.095000 0.485000 ;
      RECT  197.795000  1.825000  198.125000 2.425000 ;
      RECT  197.955000  0.825000  198.125000 1.825000 ;
      RECT  198.115000  4.615000  198.445000 5.185000 ;
      RECT  198.210000  3.905000  198.380000 4.615000 ;
      RECT  198.345000  0.085000  198.635000 0.810000 ;
      RECT  198.345000  1.470000  198.635000 2.635000 ;
      RECT  198.545000  2.975000  198.830000 3.575000 ;
      RECT  198.550000  4.115000  199.045000 4.445000 ;
      RECT  198.810000  0.085000  199.145000 0.465000 ;
      RECT  198.810000  0.715000  199.535000 0.885000 ;
      RECT  198.810000  0.885000  199.065000 1.835000 ;
      RECT  198.810000  1.835000  199.535000 2.005000 ;
      RECT  198.855000  2.175000  199.105000 2.635000 ;
      RECT  198.975000  4.615000  199.305000 5.355000 ;
      RECT  199.005000  2.805000  199.305000 3.290000 ;
      RECT  199.005000  3.290000  199.335000 3.555000 ;
      RECT  199.215000  3.905000  199.385000 4.115000 ;
      RECT  199.215000  4.115000  199.525000 4.445000 ;
      RECT  199.235000  1.075000  199.565000 1.245000 ;
      RECT  199.235000  1.245000  199.405000 1.495000 ;
      RECT  199.235000  1.495000  202.065000 1.665000 ;
      RECT  199.365000  0.255000  199.535000 0.715000 ;
      RECT  199.365000  2.005000  199.535000 2.465000 ;
      RECT  199.475000  2.985000  199.865000 3.185000 ;
      RECT  199.475000  4.615000  199.865000 5.185000 ;
      RECT  199.555000  3.185000  199.865000 3.945000 ;
      RECT  199.695000  3.945000  199.865000 4.115000 ;
      RECT  199.695000  4.115000  200.095000 4.385000 ;
      RECT  199.695000  4.385000  199.865000 4.615000 ;
      RECT  199.705000  1.835000  200.005000 2.635000 ;
      RECT  199.725000  0.085000  200.105000 0.465000 ;
      RECT  199.750000  0.760000  200.090000 0.995000 ;
      RECT  199.750000  0.995000  200.265000 1.325000 ;
      RECT  200.035000  2.805000  200.240000 3.945000 ;
      RECT  200.035000  4.555000  200.245000 5.355000 ;
      RECT  200.175000  1.835000  201.615000 2.005000 ;
      RECT  200.175000  2.005000  200.475000 2.425000 ;
      RECT  200.625000  0.400000  200.875000 1.325000 ;
      RECT  200.645000  2.805000  200.935000 3.970000 ;
      RECT  200.645000  4.630000  200.935000 5.355000 ;
      RECT  200.735000  2.175000  201.065000 2.635000 ;
      RECT  201.105000  0.415000  201.335000 1.325000 ;
      RECT  201.105000  2.975000  201.415000 3.475000 ;
      RECT  201.105000  3.475000  201.795000 3.645000 ;
      RECT  201.105000  3.815000  201.455000 4.455000 ;
      RECT  201.245000  4.635000  201.795000 4.805000 ;
      RECT  201.245000  4.805000  201.415000 5.160000 ;
      RECT  201.305000  2.005000  201.615000 2.425000 ;
      RECT  201.505000  0.255000  201.675000 1.495000 ;
      RECT  201.585000  2.805000  201.915000 3.305000 ;
      RECT  201.585000  4.975000  201.915000 5.355000 ;
      RECT  201.625000  3.645000  201.795000 4.040000 ;
      RECT  201.625000  4.040000  201.915000 4.370000 ;
      RECT  201.625000  4.370000  201.795000 4.635000 ;
      RECT  201.895000  0.085000  202.185000 0.565000 ;
      RECT  201.895000  1.665000  202.065000 2.465000 ;
      RECT  201.915000  0.755000  202.255000 1.325000 ;
      RECT  202.085000  2.975000  202.355000 3.755000 ;
      RECT  202.085000  3.755000  202.255000 5.160000 ;
      RECT  202.455000  4.115000  202.785000 4.485000 ;
      RECT  202.485000  0.085000  202.775000 0.810000 ;
      RECT  202.485000  1.470000  202.775000 2.635000 ;
      RECT  202.575000  2.975000  202.905000 3.775000 ;
      RECT  202.575000  3.775000  203.135000 3.945000 ;
      RECT  202.680000  4.655000  203.555000 4.675000 ;
      RECT  202.680000  4.675000  203.135000 4.825000 ;
      RECT  202.680000  4.825000  202.875000 5.095000 ;
      RECT  202.965000  3.945000  203.135000 4.345000 ;
      RECT  202.965000  4.345000  203.555000 4.655000 ;
      RECT  203.005000  1.075000  203.385000 1.445000 ;
      RECT  203.005000  1.445000  206.015000 1.615000 ;
      RECT  203.035000  0.085000  203.205000 0.905000 ;
      RECT  203.035000  1.785000  206.145000 1.955000 ;
      RECT  203.035000  1.955000  203.205000 2.465000 ;
      RECT  203.045000  4.995000  203.375000 5.355000 ;
      RECT  203.075000  2.805000  203.345000 3.605000 ;
      RECT  203.375000  2.125000  203.755000 2.635000 ;
      RECT  203.465000  3.755000  203.975000 4.175000 ;
      RECT  203.635000  0.735000  205.230000 0.905000 ;
      RECT  203.635000  0.905000  204.115000 1.275000 ;
      RECT  203.800000  4.345000  204.315000 4.705000 ;
      RECT  203.975000  1.955000  204.145000 2.465000 ;
      RECT  204.040000  3.055000  204.870000 3.275000 ;
      RECT  204.060000  4.875000  204.680000 5.160000 ;
      RECT  204.145000  3.445000  204.530000 3.865000 ;
      RECT  204.145000  3.865000  204.315000 4.345000 ;
      RECT  204.315000  0.395000  205.630000 0.565000 ;
      RECT  204.315000  1.075000  204.715000 1.275000 ;
      RECT  204.315000  2.125000  204.695000 2.635000 ;
      RECT  204.510000  4.275000  205.400000 4.445000 ;
      RECT  204.510000  4.445000  204.680000 4.875000 ;
      RECT  204.700000  3.275000  204.870000 4.115000 ;
      RECT  204.700000  4.115000  205.400000 4.275000 ;
      RECT  204.890000  4.830000  205.220000 5.355000 ;
      RECT  204.915000  1.955000  205.085000 2.465000 ;
      RECT  205.040000  3.575000  206.190000 3.735000 ;
      RECT  205.040000  3.735000  206.745000 3.905000 ;
      RECT  205.045000  0.905000  205.230000 1.075000 ;
      RECT  205.045000  1.075000  205.425000 1.275000 ;
      RECT  205.070000  2.805000  205.655000 3.305000 ;
      RECT  205.255000  2.125000  205.635000 2.635000 ;
      RECT  205.460000  0.565000  205.630000 0.700000 ;
      RECT  205.460000  0.700000  206.695000 0.805000 ;
      RECT  205.460000  0.805000  206.555000 0.870000 ;
      RECT  205.475000  4.615000  205.805000 5.185000 ;
      RECT  205.570000  3.905000  205.740000 4.615000 ;
      RECT  205.635000  1.075000  206.015000 1.445000 ;
      RECT  205.810000  0.085000  206.145000 0.530000 ;
      RECT  205.905000  2.975000  206.190000 3.575000 ;
      RECT  205.910000  4.115000  206.405000 4.445000 ;
      RECT  205.975000  1.955000  206.145000 2.295000 ;
      RECT  205.975000  2.295000  207.085000 2.465000 ;
      RECT  206.315000  0.295000  206.695000 0.700000 ;
      RECT  206.315000  0.870000  206.555000 1.455000 ;
      RECT  206.315000  1.455000  207.680000 1.625000 ;
      RECT  206.315000  1.625000  206.695000 2.115000 ;
      RECT  206.335000  4.615000  206.665000 5.355000 ;
      RECT  206.365000  2.805000  206.665000 3.290000 ;
      RECT  206.365000  3.290000  206.695000 3.555000 ;
      RECT  206.575000  3.905000  206.745000 4.115000 ;
      RECT  206.575000  4.115000  206.885000 4.445000 ;
      RECT  206.785000  1.075000  207.315000 1.285000 ;
      RECT  206.835000  2.985000  207.225000 3.185000 ;
      RECT  206.835000  4.615000  207.225000 5.185000 ;
      RECT  206.915000  1.795000  207.085000 2.295000 ;
      RECT  206.915000  3.185000  207.225000 3.945000 ;
      RECT  206.995000  0.085000  207.525000 0.565000 ;
      RECT  207.055000  3.945000  207.225000 4.115000 ;
      RECT  207.055000  4.115000  207.455000 4.385000 ;
      RECT  207.055000  4.385000  207.225000 4.615000 ;
      RECT  207.075000  0.745000  207.315000 1.075000 ;
      RECT  207.355000  2.125000  207.685000 2.635000 ;
      RECT  207.395000  2.805000  207.600000 3.945000 ;
      RECT  207.395000  4.555000  207.605000 5.355000 ;
      RECT  207.510000  0.995000  209.215000 1.325000 ;
      RECT  207.510000  1.325000  207.680000 1.455000 ;
      RECT  207.765000  0.655000  209.640000 0.825000 ;
      RECT  207.795000  1.785000  209.640000 1.955000 ;
      RECT  207.905000  1.955000  208.075000 2.465000 ;
      RECT  208.005000  2.805000  208.295000 3.970000 ;
      RECT  208.005000  4.630000  208.295000 5.355000 ;
      RECT  208.245000  0.085000  208.625000 0.485000 ;
      RECT  208.245000  2.125000  208.625000 2.635000 ;
      RECT  208.465000  2.975000  208.775000 3.475000 ;
      RECT  208.465000  3.475000  209.275000 3.645000 ;
      RECT  208.465000  3.815000  208.815000 4.455000 ;
      RECT  208.605000  4.635000  209.155000 4.805000 ;
      RECT  208.605000  4.805000  208.775000 5.160000 ;
      RECT  208.845000  1.955000  209.015000 2.465000 ;
      RECT  208.945000  2.805000  209.275000 3.305000 ;
      RECT  208.945000  4.975000  209.275000 5.355000 ;
      RECT  208.985000  3.645000  209.275000 4.370000 ;
      RECT  208.985000  4.370000  209.155000 4.635000 ;
      RECT  209.185000  0.085000  209.565000 0.485000 ;
      RECT  209.185000  2.125000  209.565000 2.635000 ;
      RECT  209.445000  0.825000  209.640000 1.785000 ;
      RECT  209.445000  2.975000  209.715000 3.995000 ;
      RECT  209.445000  3.995000  209.615000 5.160000 ;
      RECT  209.815000  4.140000  210.145000 4.485000 ;
      RECT  209.845000  0.085000  210.135000 0.810000 ;
      RECT  209.845000  1.470000  210.135000 2.635000 ;
      RECT  209.935000  2.975000  210.265000 3.775000 ;
      RECT  209.935000  3.775000  210.495000 3.945000 ;
      RECT  210.040000  4.655000  210.915000 4.675000 ;
      RECT  210.040000  4.675000  210.495000 4.825000 ;
      RECT  210.040000  4.825000  210.235000 5.095000 ;
      RECT  210.305000  0.995000  210.655000 1.325000 ;
      RECT  210.310000  0.085000  210.650000 0.815000 ;
      RECT  210.310000  1.495000  210.640000 2.635000 ;
      RECT  210.325000  3.945000  210.495000 4.345000 ;
      RECT  210.325000  4.345000  210.915000 4.655000 ;
      RECT  210.405000  4.995000  210.735000 5.355000 ;
      RECT  210.435000  2.805000  210.705000 3.605000 ;
      RECT  210.825000  0.335000  211.385000 1.275000 ;
      RECT  210.825000  3.755000  211.335000 4.175000 ;
      RECT  210.860000  1.835000  212.035000 2.005000 ;
      RECT  210.860000  2.005000  211.035000 2.415000 ;
      RECT  211.160000  4.345000  211.675000 4.705000 ;
      RECT  211.255000  2.175000  211.585000 2.635000 ;
      RECT  211.285000  1.445000  211.915000 1.665000 ;
      RECT  211.400000  3.055000  212.230000 3.275000 ;
      RECT  211.420000  4.875000  212.040000 5.160000 ;
      RECT  211.505000  3.445000  211.890000 3.865000 ;
      RECT  211.505000  3.865000  211.675000 4.345000 ;
      RECT  211.590000  0.995000  211.915000 1.445000 ;
      RECT  211.700000  0.295000  212.375000 0.825000 ;
      RECT  211.840000  2.005000  212.035000 2.415000 ;
      RECT  211.870000  4.275000  212.760000 4.445000 ;
      RECT  211.870000  4.445000  212.040000 4.875000 ;
      RECT  212.060000  3.275000  212.230000 4.115000 ;
      RECT  212.060000  4.115000  212.760000 4.275000 ;
      RECT  212.205000  0.825000  212.375000 1.495000 ;
      RECT  212.205000  1.495000  212.630000 2.445000 ;
      RECT  212.250000  4.830000  212.580000 5.355000 ;
      RECT  212.400000  2.805000  213.085000 3.305000 ;
      RECT  212.400000  3.575000  213.555000 3.735000 ;
      RECT  212.400000  3.735000  214.105000 3.905000 ;
      RECT  212.545000  0.085000  212.805000 0.565000 ;
      RECT  212.545000  0.995000  212.870000 1.325000 ;
      RECT  212.835000  4.615000  213.165000 5.185000 ;
      RECT  212.930000  3.905000  213.100000 4.615000 ;
      RECT  213.065000  0.085000  213.355000 0.810000 ;
      RECT  213.065000  1.470000  213.355000 2.635000 ;
      RECT  213.255000  3.005000  213.555000 3.575000 ;
      RECT  213.270000  4.115000  213.765000 4.445000 ;
      RECT  213.535000  0.655000  215.745000 0.825000 ;
      RECT  213.585000  0.995000  214.310000 1.615000 ;
      RECT  213.615000  1.785000  217.295000 1.955000 ;
      RECT  213.615000  1.955000  213.785000 2.465000 ;
      RECT  213.695000  4.615000  214.025000 5.355000 ;
      RECT  213.725000  2.805000  214.025000 3.290000 ;
      RECT  213.725000  3.290000  214.055000 3.565000 ;
      RECT  213.935000  3.905000  214.105000 4.115000 ;
      RECT  213.935000  4.115000  214.615000 4.365000 ;
      RECT  213.955000  0.085000  214.335000 0.465000 ;
      RECT  213.955000  2.125000  214.335000 2.635000 ;
      RECT  214.195000  2.975000  214.525000 3.185000 ;
      RECT  214.195000  4.535000  215.465000 4.705000 ;
      RECT  214.195000  4.705000  214.575000 5.185000 ;
      RECT  214.225000  3.185000  214.525000 3.565000 ;
      RECT  214.275000  3.565000  214.525000 3.775000 ;
      RECT  214.275000  3.775000  215.465000 3.945000 ;
      RECT  214.555000  1.955000  214.725000 2.465000 ;
      RECT  214.590000  0.995000  215.345000 1.615000 ;
      RECT  214.695000  2.805000  214.965000 3.605000 ;
      RECT  214.755000  4.875000  214.965000 5.355000 ;
      RECT  214.785000  3.945000  215.465000 4.115000 ;
      RECT  214.785000  4.115000  215.645000 4.385000 ;
      RECT  214.785000  4.385000  215.465000 4.535000 ;
      RECT  214.895000  0.295000  216.815000 0.465000 ;
      RECT  214.895000  2.125000  215.275000 2.635000 ;
      RECT  215.135000  2.975000  215.465000 3.775000 ;
      RECT  215.135000  4.705000  215.465000 5.185000 ;
      RECT  215.495000  1.955000  215.665000 2.465000 ;
      RECT  215.635000  2.805000  215.890000 3.945000 ;
      RECT  215.635000  4.555000  215.845000 5.355000 ;
      RECT  215.770000  0.995000  216.530000 1.615000 ;
      RECT  215.985000  0.655000  218.395000 0.825000 ;
      RECT  216.000000  2.125000  216.720000 2.635000 ;
      RECT  216.285000  2.805000  216.575000 3.970000 ;
      RECT  216.285000  4.630000  216.575000 5.355000 ;
      RECT  216.745000  2.975000  217.055000 3.475000 ;
      RECT  216.745000  3.475000  217.435000 3.645000 ;
      RECT  216.745000  3.815000  217.095000 4.455000 ;
      RECT  216.770000  0.825000  218.395000 0.845000 ;
      RECT  216.770000  0.845000  217.085000 1.445000 ;
      RECT  216.770000  1.445000  217.925000 1.615000 ;
      RECT  216.885000  4.635000  217.435000 4.805000 ;
      RECT  216.885000  4.805000  217.055000 5.160000 ;
      RECT  217.045000  0.255000  217.215000 0.655000 ;
      RECT  217.125000  1.955000  217.295000 2.295000 ;
      RECT  217.125000  2.295000  218.315000 2.465000 ;
      RECT  217.225000  2.805000  217.555000 3.305000 ;
      RECT  217.225000  4.975000  217.555000 5.355000 ;
      RECT  217.265000  3.645000  217.435000 4.040000 ;
      RECT  217.265000  4.040000  217.555000 4.370000 ;
      RECT  217.265000  4.370000  217.435000 4.635000 ;
      RECT  217.465000  0.085000  217.845000 0.465000 ;
      RECT  217.595000  1.615000  217.925000 2.115000 ;
      RECT  217.660000  1.075000  218.380000 1.275000 ;
      RECT  217.725000  2.975000  217.995000 3.755000 ;
      RECT  217.725000  3.755000  217.895000 5.160000 ;
      RECT  218.015000  0.295000  218.395000 0.655000 ;
      RECT  218.095000  4.115000  218.425000 4.485000 ;
      RECT  218.145000  1.795000  218.315000 2.295000 ;
      RECT  218.155000  1.275000  218.380000 1.625000 ;
      RECT  218.215000  2.975000  218.545000 3.775000 ;
      RECT  218.215000  3.775000  218.775000 3.945000 ;
      RECT  218.320000  4.655000  219.195000 4.675000 ;
      RECT  218.320000  4.675000  218.775000 4.825000 ;
      RECT  218.320000  4.825000  218.515000 5.095000 ;
      RECT  218.585000  0.085000  218.875000 0.810000 ;
      RECT  218.585000  1.470000  218.875000 2.635000 ;
      RECT  218.605000  3.945000  218.775000 4.345000 ;
      RECT  218.605000  4.345000  219.195000 4.655000 ;
      RECT  218.685000  4.995000  219.015000 5.355000 ;
      RECT  218.715000  2.805000  218.985000 3.605000 ;
      RECT  219.080000  0.995000  220.845000 1.325000 ;
      RECT  219.105000  3.755000  219.615000 4.175000 ;
      RECT  219.135000  0.255000  219.305000 0.635000 ;
      RECT  219.135000  0.635000  223.145000 0.805000 ;
      RECT  219.135000  1.495000  224.965000 1.665000 ;
      RECT  219.135000  1.665000  219.305000 2.465000 ;
      RECT  219.440000  4.345000  219.955000 4.705000 ;
      RECT  219.475000  0.085000  219.855000 0.465000 ;
      RECT  219.475000  1.915000  219.855000 2.635000 ;
      RECT  219.680000  3.055000  220.510000 3.275000 ;
      RECT  219.700000  4.875000  220.320000 5.160000 ;
      RECT  219.785000  3.445000  220.170000 3.865000 ;
      RECT  219.785000  3.865000  219.955000 4.345000 ;
      RECT  220.075000  0.255000  220.245000 0.635000 ;
      RECT  220.075000  1.665000  220.245000 2.465000 ;
      RECT  220.150000  4.275000  221.040000 4.445000 ;
      RECT  220.150000  4.445000  220.320000 4.875000 ;
      RECT  220.340000  3.275000  220.510000 4.115000 ;
      RECT  220.340000  4.115000  221.040000 4.275000 ;
      RECT  220.415000  0.085000  220.795000 0.465000 ;
      RECT  220.415000  1.915000  220.795000 2.635000 ;
      RECT  220.530000  4.830000  220.860000 5.355000 ;
      RECT  220.680000  2.805000  221.365000 3.305000 ;
      RECT  220.680000  3.575000  221.835000 3.735000 ;
      RECT  220.680000  3.735000  222.385000 3.905000 ;
      RECT  221.015000  0.255000  221.185000 0.635000 ;
      RECT  221.015000  1.665000  221.185000 2.465000 ;
      RECT  221.095000  0.995000  222.910000 1.325000 ;
      RECT  221.115000  4.615000  221.445000 5.185000 ;
      RECT  221.210000  3.905000  221.380000 4.615000 ;
      RECT  221.355000  0.295000  225.125000 0.465000 ;
      RECT  221.355000  1.915000  221.735000 2.635000 ;
      RECT  221.535000  3.005000  221.835000 3.575000 ;
      RECT  221.550000  4.115000  222.045000 4.445000 ;
      RECT  221.955000  1.665000  222.125000 2.465000 ;
      RECT  221.975000  4.615000  222.305000 5.355000 ;
      RECT  222.005000  2.805000  222.305000 3.290000 ;
      RECT  222.005000  3.290000  222.335000 3.565000 ;
      RECT  222.215000  3.905000  222.385000 4.115000 ;
      RECT  222.215000  4.115000  222.895000 4.365000 ;
      RECT  222.295000  1.915000  222.675000 2.635000 ;
      RECT  222.475000  2.975000  222.805000 3.185000 ;
      RECT  222.475000  4.535000  223.745000 4.705000 ;
      RECT  222.475000  4.705000  222.855000 5.185000 ;
      RECT  222.505000  3.185000  222.805000 3.565000 ;
      RECT  222.555000  3.565000  222.805000 3.775000 ;
      RECT  222.555000  3.775000  223.745000 3.945000 ;
      RECT  222.895000  1.665000  223.065000 2.465000 ;
      RECT  222.975000  2.805000  223.245000 3.605000 ;
      RECT  223.035000  4.875000  223.245000 5.355000 ;
      RECT  223.065000  3.945000  223.745000 4.115000 ;
      RECT  223.065000  4.115000  223.925000 4.385000 ;
      RECT  223.065000  4.385000  223.745000 4.535000 ;
      RECT  223.185000  0.995000  224.980000 1.325000 ;
      RECT  223.255000  1.915000  223.635000 2.635000 ;
      RECT  223.385000  0.635000  227.395000 0.805000 ;
      RECT  223.415000  2.975000  223.745000 3.775000 ;
      RECT  223.415000  4.705000  223.745000 5.185000 ;
      RECT  223.855000  1.665000  224.025000 2.465000 ;
      RECT  223.915000  2.805000  224.170000 3.945000 ;
      RECT  223.915000  4.555000  224.125000 5.355000 ;
      RECT  224.195000  2.255000  224.575000 2.635000 ;
      RECT  224.565000  2.805000  224.855000 3.970000 ;
      RECT  224.565000  4.630000  224.855000 5.355000 ;
      RECT  224.795000  1.665000  224.965000 2.255000 ;
      RECT  224.795000  2.255000  227.475000 2.425000 ;
      RECT  224.795000  2.425000  224.965000 2.465000 ;
      RECT  225.025000  2.975000  225.775000 5.185000 ;
      RECT  225.230000  0.995000  226.565000 1.630000 ;
      RECT  225.685000  0.085000  226.065000 0.465000 ;
      RECT  225.685000  1.915000  227.045000 2.085000 ;
      RECT  225.945000  2.975000  227.615000 5.185000 ;
      RECT  226.285000  0.255000  226.455000 0.635000 ;
      RECT  226.625000  0.085000  227.005000 0.465000 ;
      RECT  226.805000  0.805000  227.045000 1.915000 ;
      RECT  227.225000  0.255000  227.395000 0.635000 ;
      RECT  227.225000  1.495000  227.475000 2.255000 ;
      RECT  227.785000  0.085000  228.075000 0.810000 ;
      RECT  227.785000  1.470000  228.075000 2.635000 ;
      RECT  227.785000  2.975000  230.375000 5.185000 ;
      RECT  228.250000  0.300000  228.585000 0.560000 ;
      RECT  228.250000  0.560000  228.505000 1.915000 ;
      RECT  228.250000  1.915000  228.585000 2.425000 ;
      RECT  228.730000  0.995000  229.005000 1.325000 ;
      RECT  228.755000  0.085000  229.135000 0.485000 ;
      RECT  228.835000  0.655000  229.475000 0.825000 ;
      RECT  228.835000  0.825000  229.005000 0.995000 ;
      RECT  228.835000  1.325000  229.005000 1.495000 ;
      RECT  228.835000  1.495000  231.485000 1.665000 ;
      RECT  228.885000  1.835000  229.215000 2.635000 ;
      RECT  229.175000  0.995000  229.515000 1.325000 ;
      RECT  229.305000  0.315000  231.070000 0.485000 ;
      RECT  229.305000  0.485000  229.475000 0.655000 ;
      RECT  229.510000  1.875000  231.035000 2.045000 ;
      RECT  229.510000  2.045000  229.795000 2.465000 ;
      RECT  229.685000  0.665000  230.110000 1.325000 ;
      RECT  230.100000  2.215000  230.430000 2.635000 ;
      RECT  230.420000  0.955000  230.825000 1.325000 ;
      RECT  230.540000  0.665000  230.825000 0.955000 ;
      RECT  230.545000  2.975000  234.055000 5.185000 ;
      RECT  230.705000  2.045000  231.035000 2.295000 ;
      RECT  230.705000  2.295000  232.055000 2.465000 ;
      RECT  230.995000  0.660000  231.295000 1.325000 ;
      RECT  231.315000  1.665000  231.485000 2.125000 ;
      RECT  231.590000  0.995000  232.190000 1.325000 ;
      RECT  231.665000  0.085000  232.045000 0.805000 ;
      RECT  231.795000  1.795000  232.055000 2.295000 ;
      RECT  231.950000  1.325000  232.190000 1.615000 ;
      RECT  232.385000  0.085000  232.675000 0.810000 ;
      RECT  232.385000  1.470000  232.675000 2.635000 ;
      RECT  232.850000  0.085000  233.185000 0.465000 ;
      RECT  232.895000  0.655000  233.655000 0.825000 ;
      RECT  232.895000  0.825000  233.105000 1.785000 ;
      RECT  232.895000  1.785000  234.045000 1.955000 ;
      RECT  232.895000  1.955000  233.105000 2.465000 ;
      RECT  233.275000  2.125000  233.655000 2.635000 ;
      RECT  233.295000  0.995000  233.515000 1.445000 ;
      RECT  233.295000  1.445000  235.035000 1.615000 ;
      RECT  233.745000  0.085000  234.500000 0.445000 ;
      RECT  233.825000  0.745000  234.390000 1.275000 ;
      RECT  233.875000  1.955000  234.045000 2.465000 ;
      RECT  234.225000  2.805000  234.515000 3.970000 ;
      RECT  234.225000  4.630000  234.515000 5.355000 ;
      RECT  234.395000  1.785000  234.565000 2.295000 ;
      RECT  234.395000  2.295000  235.505000 2.465000 ;
      RECT  234.560000  0.675000  235.465000 0.845000 ;
      RECT  234.560000  0.845000  234.800000 1.445000 ;
      RECT  234.785000  1.615000  235.035000 1.945000 ;
      RECT  234.785000  1.945000  235.115000 2.115000 ;
      RECT  234.995000  1.075000  235.430000 1.245000 ;
      RECT  235.165000  0.295000  235.465000 0.675000 ;
      RECT  235.205000  1.245000  235.430000 1.615000 ;
      RECT  235.335000  1.795000  236.605000 1.965000 ;
      RECT  235.335000  1.965000  235.505000 2.295000 ;
      RECT  235.635000  0.415000  235.905000 1.325000 ;
      RECT  235.675000  2.140000  236.055000 2.635000 ;
      RECT  236.075000  0.425000  236.410000 1.625000 ;
      RECT  236.435000  1.965000  236.605000 2.465000 ;
      RECT  236.775000  0.085000  237.160000 0.805000 ;
      RECT  236.775000  1.915000  237.160000 2.635000 ;
      RECT  236.925000  0.995000  237.265000 1.630000 ;
      RECT  237.445000  0.085000  237.735000 0.810000 ;
      RECT  237.445000  1.470000  237.735000 2.635000 ;
      RECT  237.915000  0.085000  238.245000 0.465000 ;
      RECT  237.915000  1.915000  238.245000 2.635000 ;
      RECT  237.940000  0.635000  239.575000 0.805000 ;
      RECT  237.940000  0.805000  238.160000 1.495000 ;
      RECT  237.940000  1.495000  239.575000 1.665000 ;
      RECT  238.440000  0.995000  239.990000 1.325000 ;
      RECT  238.465000  0.255000  238.635000 0.635000 ;
      RECT  238.465000  1.665000  238.635000 2.465000 ;
      RECT  238.805000  0.085000  239.185000 0.465000 ;
      RECT  238.805000  1.915000  239.185000 2.635000 ;
      RECT  239.405000  0.255000  239.575000 0.635000 ;
      RECT  239.405000  1.665000  239.575000 2.465000 ;
      RECT  239.745000  0.085000  240.125000 0.465000 ;
      RECT  239.745000  1.915000  240.125000 2.635000 ;
      RECT  239.770000  1.325000  239.990000 1.495000 ;
      RECT  239.770000  1.495000  243.770000 1.665000 ;
      RECT  240.230000  1.075000  241.225000 1.295000 ;
      RECT  240.345000  0.255000  240.515000 0.655000 ;
      RECT  240.345000  0.655000  242.055000 0.825000 ;
      RECT  240.345000  1.915000  243.385000 2.085000 ;
      RECT  240.345000  2.085000  240.515000 2.465000 ;
      RECT  240.685000  0.085000  241.065000 0.465000 ;
      RECT  240.685000  2.255000  241.065000 2.635000 ;
      RECT  241.255000  0.295000  243.465000 0.465000 ;
      RECT  241.335000  2.085000  241.505000 2.465000 ;
      RECT  241.455000  1.075000  242.250000 1.325000 ;
      RECT  241.675000  2.255000  242.055000 2.635000 ;
      RECT  242.275000  2.085000  242.445000 2.465000 ;
      RECT  242.500000  1.075000  243.395000 1.325000 ;
      RECT  242.615000  0.635000  244.555000 0.805000 ;
      RECT  242.615000  2.255000  242.995000 2.635000 ;
      RECT  243.215000  2.085000  243.385000 2.255000 ;
      RECT  243.215000  2.255000  246.005000 2.425000 ;
      RECT  243.600000  0.805000  243.770000 1.495000 ;
      RECT  243.600000  1.665000  243.770000 1.905000 ;
      RECT  243.600000  1.905000  244.330000 1.915000 ;
      RECT  243.600000  1.915000  245.535000 2.075000 ;
      RECT  243.750000  0.295000  244.985000 0.465000 ;
      RECT  243.940000  1.075000  244.960000 1.625000 ;
      RECT  244.265000  2.075000  245.535000 2.085000 ;
      RECT  244.815000  0.255000  244.985000 0.295000 ;
      RECT  244.815000  0.465000  244.985000 0.645000 ;
      RECT  244.815000  0.645000  245.925000 0.815000 ;
      RECT  245.155000  0.085000  245.535000 0.465000 ;
      RECT  245.260000  1.075000  245.990000 1.295000 ;
      RECT  245.260000  1.295000  245.455000 1.635000 ;
      RECT  245.755000  0.255000  245.925000 0.645000 ;
      RECT  245.755000  1.755000  246.005000 2.255000 ;
      RECT  246.185000  0.085000  246.475000 0.810000 ;
      RECT  246.185000  1.470000  246.475000 2.635000 ;
      RECT  246.645000  0.995000  246.905000 1.325000 ;
      RECT  246.645000  1.835000  246.905000 2.255000 ;
      RECT  246.645000  2.255000  248.005000 2.465000 ;
      RECT  246.670000  0.085000  247.000000 0.465000 ;
      RECT  247.075000  0.635000  247.825000 0.805000 ;
      RECT  247.075000  0.805000  247.335000 1.785000 ;
      RECT  247.075000  1.785000  247.475000 2.085000 ;
      RECT  247.505000  0.995000  247.795000 1.615000 ;
      RECT  247.525000  0.295000  247.825000 0.635000 ;
      RECT  247.755000  1.785000  248.945000 1.955000 ;
      RECT  247.755000  1.955000  248.005000 2.255000 ;
      RECT  248.035000  0.345000  248.255000 1.325000 ;
      RECT  248.265000  2.135000  248.515000 2.635000 ;
      RECT  248.545000  0.415000  248.745000 1.325000 ;
      RECT  248.775000  1.745000  248.945000 1.785000 ;
      RECT  248.775000  1.955000  248.945000 2.465000 ;
      RECT  248.950000  1.015000  249.415000 1.325000 ;
      RECT  249.115000  1.495000  249.505000 2.635000 ;
      RECT  249.130000  0.085000  249.520000 0.805000 ;
      RECT  249.865000  0.085000  250.155000 0.810000 ;
      RECT  249.865000  1.470000  250.155000 2.635000 ;
      RECT  250.335000  0.295000  250.665000 0.715000 ;
      RECT  250.335000  0.715000  251.525000 0.885000 ;
      RECT  250.385000  1.075000  251.115000 1.285000 ;
      RECT  250.385000  1.285000  250.565000 1.625000 ;
      RECT  250.415000  1.795000  250.585000 2.295000 ;
      RECT  250.415000  2.295000  252.465000 2.465000 ;
      RECT  250.805000  1.455000  252.435000 1.625000 ;
      RECT  250.805000  1.625000  251.135000 2.125000 ;
      RECT  250.885000  0.085000  251.055000 0.545000 ;
      RECT  251.275000  0.295000  252.545000 0.465000 ;
      RECT  251.275000  0.465000  251.525000 0.715000 ;
      RECT  251.305000  1.075000  252.035000 1.285000 ;
      RECT  251.355000  1.795000  251.525000 2.295000 ;
      RECT  251.695000  0.655000  253.485000 0.825000 ;
      RECT  251.825000  1.625000  251.995000 2.125000 ;
      RECT  252.205000  0.825000  252.435000 1.455000 ;
      RECT  252.295000  1.795000  256.505000 1.965000 ;
      RECT  252.295000  1.965000  252.465000 2.295000 ;
      RECT  252.615000  1.075000  253.495000 1.625000 ;
      RECT  252.685000  2.255000  253.405000 2.635000 ;
      RECT  252.735000  0.295000  254.845000 0.465000 ;
      RECT  253.655000  1.965000  253.825000 2.465000 ;
      RECT  253.960000  1.075000  254.815000 1.625000 ;
      RECT  253.995000  0.635000  256.040000 0.805000 ;
      RECT  254.010000  2.255000  254.765000 2.635000 ;
      RECT  254.935000  1.965000  255.105000 2.465000 ;
      RECT  255.105000  0.085000  255.490000 0.465000 ;
      RECT  255.265000  1.075000  256.560000 1.625000 ;
      RECT  255.365000  2.255000  256.085000 2.635000 ;
      RECT  255.660000  0.275000  256.040000 0.635000 ;
      RECT  256.335000  0.085000  256.505000 0.885000 ;
      RECT  256.335000  1.965000  256.505000 2.465000 ;
      RECT  256.765000  0.085000  257.055000 0.810000 ;
      RECT  256.765000  1.470000  257.055000 2.635000 ;
      RECT  257.235000  2.255000  261.245000 2.425000 ;
      RECT  257.250000  1.075000  259.040000 1.305000 ;
      RECT  257.250000  1.305000  257.470000 1.965000 ;
      RECT  257.315000  0.255000  257.485000 0.635000 ;
      RECT  257.315000  0.635000  259.365000 0.805000 ;
      RECT  257.655000  0.085000  258.035000 0.465000 ;
      RECT  257.655000  1.575000  260.855000 1.745000 ;
      RECT  257.655000  1.745000  258.035000 2.085000 ;
      RECT  258.255000  0.255000  258.425000 0.635000 ;
      RECT  258.595000  0.085000  258.975000 0.465000 ;
      RECT  258.595000  1.745000  258.975000 2.085000 ;
      RECT  259.195000  0.295000  261.325000 0.465000 ;
      RECT  259.195000  0.465000  259.365000 0.635000 ;
      RECT  259.315000  0.990000  259.755000 1.575000 ;
      RECT  259.315000  1.745000  259.915000 2.085000 ;
      RECT  259.535000  0.635000  263.305000 0.805000 ;
      RECT  259.535000  0.805000  259.755000 0.990000 ;
      RECT  259.975000  0.995000  261.095000 1.325000 ;
      RECT  260.475000  1.745000  260.855000 2.085000 ;
      RECT  261.075000  1.575000  268.115000 1.745000 ;
      RECT  261.075000  1.745000  261.245000 2.255000 ;
      RECT  261.315000  1.075000  263.205000 1.285000 ;
      RECT  261.435000  1.915000  261.815000 2.635000 ;
      RECT  261.565000  0.295000  265.795000 0.465000 ;
      RECT  262.035000  1.745000  262.205000 2.465000 ;
      RECT  262.460000  1.915000  263.180000 2.635000 ;
      RECT  263.430000  1.745000  263.600000 2.465000 ;
      RECT  263.885000  1.075000  265.685000 1.300000 ;
      RECT  264.005000  0.635000  267.645000 0.805000 ;
      RECT  264.005000  1.915000  264.385000 2.635000 ;
      RECT  264.605000  1.745000  264.775000 2.465000 ;
      RECT  264.945000  1.915000  265.325000 2.635000 ;
      RECT  265.545000  1.745000  265.715000 2.465000 ;
      RECT  265.985000  0.085000  266.315000 0.465000 ;
      RECT  266.285000  1.075000  268.175000 1.280000 ;
      RECT  266.405000  1.915000  266.785000 2.635000 ;
      RECT  266.535000  0.255000  266.705000 0.635000 ;
      RECT  266.875000  0.085000  267.255000 0.465000 ;
      RECT  267.005000  1.745000  267.175000 2.465000 ;
      RECT  267.345000  1.915000  267.725000 2.635000 ;
      RECT  267.475000  0.255000  267.645000 0.635000 ;
      RECT  267.825000  0.085000  268.215000 0.465000 ;
      RECT  267.895000  0.755000  268.175000 1.075000 ;
      RECT  267.945000  1.745000  268.115000 2.465000 ;
      RECT  268.725000  0.085000  269.015000 0.810000 ;
      RECT  268.725000  1.470000  269.015000 2.635000 ;
      RECT  269.200000  1.075000  269.765000 1.325000 ;
      RECT  269.200000  1.325000  269.555000 1.685000 ;
      RECT  269.225000  0.355000  269.555000 0.715000 ;
      RECT  269.225000  0.715000  270.675000 0.905000 ;
      RECT  269.225000  1.965000  269.505000 2.635000 ;
      RECT  269.725000  1.575000  270.675000 1.745000 ;
      RECT  269.725000  1.745000  270.025000 2.295000 ;
      RECT  269.985000  1.075000  270.335000 1.325000 ;
      RECT  270.195000  1.915000  270.525000 2.635000 ;
      RECT  270.205000  0.085000  270.455000 0.545000 ;
      RECT  270.505000  0.905000  270.675000 0.995000 ;
      RECT  270.505000  0.995000  270.760000 1.325000 ;
      RECT  270.505000  1.325000  270.675000 1.575000 ;
      RECT  270.625000  0.255000  271.255000 0.545000 ;
      RECT  270.830000  1.915000  271.255000 2.465000 ;
      RECT  270.960000  0.545000  271.255000 1.915000 ;
      RECT  271.485000  0.085000  271.775000 0.810000 ;
      RECT  271.485000  1.470000  271.775000 2.635000 ;
      RECT  271.955000  1.075000  272.575000 1.325000 ;
      RECT  271.955000  1.325000  272.210000 1.765000 ;
      RECT  271.975000  0.355000  272.305000 0.715000 ;
      RECT  271.975000  0.715000  273.465000 0.905000 ;
      RECT  271.975000  1.965000  272.255000 2.635000 ;
      RECT  272.475000  1.575000  273.465000 1.745000 ;
      RECT  272.475000  1.745000  272.775000 2.295000 ;
      RECT  272.745000  1.075000  273.125000 1.325000 ;
      RECT  273.025000  1.915000  273.365000 2.635000 ;
      RECT  273.035000  0.085000  273.285000 0.545000 ;
      RECT  273.295000  0.905000  273.465000 0.995000 ;
      RECT  273.295000  0.995000  273.625000 1.325000 ;
      RECT  273.295000  1.325000  273.465000 1.575000 ;
      RECT  273.455000  0.255000  274.065000 0.545000 ;
      RECT  273.605000  1.915000  274.065000 2.465000 ;
      RECT  273.795000  0.545000  274.065000 1.915000 ;
      RECT  274.235000  0.085000  274.525000 0.885000 ;
      RECT  274.235000  1.495000  274.525000 2.635000 ;
      RECT  274.705000  0.085000  274.995000 0.810000 ;
      RECT  274.705000  1.470000  274.995000 2.635000 ;
      RECT  275.175000  0.255000  275.505000 0.615000 ;
      RECT  275.175000  0.615000  276.540000 0.805000 ;
      RECT  275.175000  1.880000  275.505000 2.635000 ;
      RECT  275.205000  0.995000  275.515000 1.615000 ;
      RECT  275.685000  0.995000  276.160000 1.325000 ;
      RECT  275.735000  1.580000  276.540000 1.750000 ;
      RECT  275.735000  1.750000  275.915000 2.465000 ;
      RECT  276.135000  0.085000  276.465000 0.445000 ;
      RECT  276.170000  1.935000  276.500000 2.635000 ;
      RECT  276.330000  0.805000  276.540000 1.020000 ;
      RECT  276.330000  1.020000  278.015000 1.355000 ;
      RECT  276.330000  1.355000  276.540000 1.580000 ;
      RECT  276.760000  0.515000  276.950000 0.615000 ;
      RECT  276.760000  0.615000  278.650000 0.845000 ;
      RECT  276.760000  1.535000  278.650000 1.760000 ;
      RECT  276.760000  1.760000  276.950000 2.465000 ;
      RECT  277.120000  0.085000  277.500000 0.445000 ;
      RECT  277.120000  1.935000  277.500000 2.635000 ;
      RECT  277.720000  0.255000  277.910000 0.615000 ;
      RECT  277.720000  1.760000  278.650000 1.765000 ;
      RECT  277.720000  1.765000  277.910000 2.465000 ;
      RECT  278.080000  0.085000  278.460000 0.445000 ;
      RECT  278.080000  1.935000  278.460000 2.635000 ;
      RECT  278.370000  0.845000  278.650000 1.535000 ;
      RECT  278.845000  0.085000  279.135000 0.810000 ;
      RECT  278.845000  1.470000  279.135000 2.635000 ;
      RECT  279.310000  0.085000  279.645000 0.590000 ;
      RECT  279.365000  0.765000  279.665000 1.615000 ;
      RECT  279.395000  1.785000  280.120000 2.015000 ;
      RECT  279.395000  2.015000  279.565000 2.445000 ;
      RECT  279.735000  2.185000  280.115000 2.635000 ;
      RECT  279.865000  0.280000  280.105000 0.655000 ;
      RECT  279.885000  0.655000  280.105000 0.805000 ;
      RECT  279.885000  0.805000  280.470000 1.135000 ;
      RECT  279.885000  1.135000  280.120000 1.785000 ;
      RECT  280.290000  1.305000  281.725000 1.325000 ;
      RECT  280.290000  1.325000  281.300000 1.475000 ;
      RECT  280.290000  1.475000  280.625000 2.420000 ;
      RECT  280.435000  0.270000  280.605000 0.415000 ;
      RECT  280.435000  0.415000  280.860000 0.610000 ;
      RECT  280.640000  0.610000  280.860000 0.945000 ;
      RECT  280.640000  0.945000  281.725000 1.305000 ;
      RECT  280.850000  1.645000  281.495000 1.955000 ;
      RECT  280.855000  2.165000  281.495000 2.635000 ;
      RECT  281.220000  0.085000  281.665000 0.580000 ;
      RECT  281.665000  1.580000  282.300000 2.365000 ;
      RECT  281.925000  0.255000  282.300000 0.775000 ;
      RECT  281.990000  0.775000  282.300000 1.580000 ;
      RECT  282.525000  0.085000  282.815000 0.810000 ;
      RECT  282.525000  1.470000  282.815000 2.635000 ;
      RECT  282.995000  0.085000  283.325000 0.590000 ;
      RECT  283.045000  0.765000  283.350000 1.615000 ;
      RECT  283.075000  1.785000  283.805000 2.015000 ;
      RECT  283.075000  2.015000  283.245000 2.445000 ;
      RECT  283.415000  2.185000  283.795000 2.635000 ;
      RECT  283.545000  0.280000  283.785000 0.655000 ;
      RECT  283.570000  0.655000  283.785000 0.805000 ;
      RECT  283.570000  0.805000  284.175000 1.135000 ;
      RECT  283.570000  1.135000  283.805000 1.785000 ;
      RECT  283.995000  1.305000  285.435000 1.325000 ;
      RECT  283.995000  1.325000  285.005000 1.475000 ;
      RECT  283.995000  1.475000  284.330000 2.420000 ;
      RECT  284.115000  0.270000  284.285000 0.415000 ;
      RECT  284.115000  0.415000  284.565000 0.610000 ;
      RECT  284.345000  0.610000  284.565000 0.945000 ;
      RECT  284.345000  0.945000  285.435000 1.305000 ;
      RECT  284.555000  1.645000  285.300000 1.955000 ;
      RECT  284.560000  2.165000  285.295000 2.635000 ;
      RECT  285.005000  0.085000  285.375000 0.580000 ;
      RECT  285.475000  1.580000  285.990000 2.365000 ;
      RECT  285.595000  0.255000  285.990000 0.775000 ;
      RECT  285.655000  0.775000  285.990000 1.580000 ;
      RECT  286.225000  0.085000  286.495000 0.720000 ;
      RECT  286.225000  1.680000  286.495000 2.635000 ;
      RECT  286.665000  0.085000  286.955000 0.810000 ;
      RECT  286.665000  1.470000  286.955000 2.635000 ;
      RECT  287.130000  0.255000  287.465000 0.615000 ;
      RECT  287.130000  0.615000  288.495000 0.805000 ;
      RECT  287.130000  2.255000  287.465000 2.635000 ;
      RECT  287.205000  0.995000  287.465000 1.325000 ;
      RECT  287.205000  1.325000  287.375000 1.915000 ;
      RECT  287.205000  1.915000  290.980000 2.085000 ;
      RECT  287.555000  1.500000  288.455000 1.745000 ;
      RECT  287.645000  0.995000  288.115000 1.325000 ;
      RECT  288.095000  0.085000  288.425000 0.445000 ;
      RECT  288.130000  2.275000  288.460000 2.635000 ;
      RECT  288.285000  0.805000  288.495000 0.995000 ;
      RECT  288.285000  0.995000  289.215000 1.355000 ;
      RECT  288.285000  1.355000  288.460000 1.485000 ;
      RECT  288.285000  1.485000  288.455000 1.500000 ;
      RECT  288.675000  1.535000  290.020000 1.745000 ;
      RECT  288.715000  0.495000  288.905000 0.615000 ;
      RECT  288.715000  0.615000  290.020000 0.825000 ;
      RECT  289.075000  0.085000  289.455000 0.445000 ;
      RECT  289.095000  2.275000  289.475000 2.635000 ;
      RECT  289.485000  0.825000  290.020000 1.535000 ;
      RECT  290.035000  0.085000  290.415000 0.445000 ;
      RECT  290.035000  2.275000  290.415000 2.635000 ;
      RECT  290.240000  0.625000  290.585000 1.745000 ;
      RECT  290.765000  0.495000  290.980000 1.915000 ;
      RECT  291.265000  0.085000  291.555000 0.810000 ;
      RECT  291.265000  1.470000  291.555000 2.635000 ;
      RECT  291.725000  0.295000  292.715000 0.465000 ;
      RECT  291.725000  0.635000  292.325000 1.020000 ;
      RECT  291.725000  1.190000  292.715000 1.360000 ;
      RECT  291.725000  1.360000  291.985000 1.810000 ;
      RECT  291.725000  1.980000  292.390000 2.080000 ;
      RECT  291.725000  2.080000  292.380000 2.635000 ;
      RECT  292.155000  1.710000  292.535000 1.955000 ;
      RECT  292.155000  1.955000  292.390000 1.980000 ;
      RECT  292.495000  0.465000  292.715000 1.190000 ;
      RECT  292.535000  1.360000  292.715000 1.370000 ;
      RECT  292.535000  1.370000  293.910000 1.540000 ;
      RECT  292.555000  2.125000  293.135000 2.465000 ;
      RECT  292.800000  1.540000  293.910000 1.590000 ;
      RECT  292.800000  1.590000  293.805000 1.885000 ;
      RECT  293.030000  0.305000  293.400000 1.200000 ;
      RECT  293.550000  2.090000  293.805000 2.635000 ;
      RECT  293.570000  0.085000  293.740000 0.625000 ;
      RECT  293.680000  0.990000  293.910000 1.370000 ;
      RECT  294.025000  1.765000  294.300000 2.465000 ;
      RECT  294.040000  0.255000  294.300000 0.735000 ;
      RECT  294.130000  0.735000  294.300000 1.765000 ;
      RECT  294.485000  0.085000  294.775000 0.810000 ;
      RECT  294.485000  1.470000  294.775000 2.635000 ;
      RECT  294.945000  0.765000  295.330000 1.245000 ;
      RECT  294.945000  2.130000  295.625000 2.635000 ;
      RECT  294.960000  1.425000  296.900000 1.595000 ;
      RECT  294.960000  1.595000  295.215000 1.960000 ;
      RECT  294.965000  0.305000  295.755000 0.570000 ;
      RECT  295.385000  1.765000  295.765000 1.955000 ;
      RECT  295.385000  1.955000  295.625000 2.130000 ;
      RECT  295.550000  0.570000  295.755000 1.425000 ;
      RECT  295.805000  2.125000  296.380000 2.465000 ;
      RECT  295.925000  0.305000  296.175000 0.750000 ;
      RECT  295.925000  0.750000  296.485000 1.245000 ;
      RECT  296.040000  1.595000  296.340000 1.890000 ;
      RECT  296.345000  0.085000  296.675000 0.580000 ;
      RECT  296.565000  1.790000  296.780000 2.635000 ;
      RECT  296.670000  0.995000  296.900000 1.425000 ;
      RECT  296.845000  0.255000  297.290000 0.715000 ;
      RECT  297.030000  1.795000  297.480000 2.465000 ;
      RECT  297.120000  0.715000  297.290000 0.925000 ;
      RECT  297.120000  0.925000  297.785000 1.445000 ;
      RECT  297.120000  1.445000  297.480000 1.795000 ;
      RECT  297.555000  0.085000  297.830000 0.745000 ;
      RECT  297.650000  1.625000  297.910000 2.635000 ;
      RECT  298.165000  0.085000  298.455000 0.810000 ;
      RECT  298.165000  1.470000  298.455000 2.635000 ;
      RECT  298.655000  0.995000  299.415000 1.340000 ;
      RECT  298.655000  1.340000  298.870000 2.335000 ;
      RECT  299.005000  0.255000  300.365000 0.445000 ;
      RECT  299.005000  0.445000  299.340000 0.805000 ;
      RECT  299.040000  1.580000  300.970000 1.750000 ;
      RECT  299.040000  1.750000  299.220000 2.465000 ;
      RECT  299.435000  1.935000  299.935000 2.635000 ;
      RECT  299.585000  0.745000  299.895000 1.340000 ;
      RECT  300.065000  0.995000  300.590000 1.325000 ;
      RECT  300.160000  1.750000  300.340000 2.465000 ;
      RECT  300.175000  0.445000  300.365000 0.615000 ;
      RECT  300.175000  0.615000  300.970000 0.805000 ;
      RECT  300.595000  0.085000  300.925000 0.445000 ;
      RECT  300.600000  1.935000  300.930000 2.635000 ;
      RECT  300.760000  0.805000  300.970000 1.020000 ;
      RECT  300.760000  1.020000  302.445000 1.355000 ;
      RECT  300.760000  1.355000  300.970000 1.580000 ;
      RECT  301.190000  0.515000  301.380000 0.615000 ;
      RECT  301.190000  0.615000  303.030000 0.845000 ;
      RECT  301.190000  1.535000  303.030000 1.760000 ;
      RECT  301.190000  1.760000  301.380000 2.465000 ;
      RECT  301.550000  0.085000  301.930000 0.445000 ;
      RECT  301.550000  1.935000  301.930000 2.635000 ;
      RECT  302.150000  0.255000  302.340000 0.615000 ;
      RECT  302.150000  1.760000  303.030000 1.765000 ;
      RECT  302.150000  1.765000  302.340000 2.465000 ;
      RECT  302.510000  0.085000  302.890000 0.445000 ;
      RECT  302.510000  1.935000  302.890000 2.635000 ;
      RECT  302.750000  0.845000  303.030000 1.535000 ;
      RECT  303.225000  0.085000  303.515000 0.810000 ;
      RECT  303.225000  1.470000  303.515000 2.635000 ;
      RECT  303.685000  0.085000  303.945000 0.905000 ;
      RECT  303.685000  1.075000  304.025000 1.955000 ;
      RECT  303.685000  2.125000  303.945000 2.635000 ;
      RECT  304.115000  0.485000  304.495000 0.905000 ;
      RECT  304.245000  0.905000  304.495000 0.995000 ;
      RECT  304.245000  0.995000  305.120000 1.245000 ;
      RECT  304.245000  1.245000  304.415000 2.465000 ;
      RECT  304.685000  1.425000  306.785000 1.575000 ;
      RECT  304.685000  1.575000  306.650000 1.595000 ;
      RECT  304.685000  1.595000  304.935000 1.940000 ;
      RECT  304.685000  2.130000  305.350000 2.635000 ;
      RECT  304.705000  0.285000  305.545000 0.550000 ;
      RECT  305.105000  1.765000  305.485000 1.955000 ;
      RECT  305.105000  1.955000  305.350000 2.130000 ;
      RECT  305.290000  0.550000  305.545000 1.425000 ;
      RECT  305.520000  2.125000  306.095000 2.465000 ;
      RECT  305.755000  1.595000  306.650000 1.890000 ;
      RECT  305.880000  0.305000  306.245000 1.255000 ;
      RECT  306.395000  2.090000  306.610000 2.635000 ;
      RECT  306.415000  0.085000  306.705000 0.625000 ;
      RECT  306.565000  0.975000  306.785000 1.425000 ;
      RECT  306.870000  1.765000  307.135000 2.465000 ;
      RECT  306.875000  0.255000  307.135000 0.735000 ;
      RECT  306.965000  0.735000  307.135000 1.765000 ;
      RECT  307.365000  0.085000  307.655000 0.810000 ;
      RECT  307.365000  1.470000  307.655000 2.635000 ;
      RECT  307.825000  0.085000  308.095000 0.575000 ;
      RECT  307.825000  1.575000  308.140000 2.635000 ;
      RECT  307.885000  0.745000  308.150000 1.325000 ;
      RECT  308.370000  0.305000  308.645000 1.015000 ;
      RECT  308.370000  1.015000  309.205000 1.245000 ;
      RECT  308.370000  1.245000  308.645000 1.905000 ;
      RECT  308.820000  2.130000  309.485000 2.635000 ;
      RECT  308.840000  1.425000  310.760000 1.595000 ;
      RECT  308.840000  1.595000  309.075000 1.960000 ;
      RECT  308.845000  0.305000  309.555000 0.570000 ;
      RECT  309.245000  1.765000  309.625000 1.955000 ;
      RECT  309.245000  1.955000  309.485000 2.130000 ;
      RECT  309.385000  0.570000  309.555000 1.425000 ;
      RECT  309.655000  2.125000  310.230000 2.465000 ;
      RECT  309.725000  0.305000  310.110000 0.765000 ;
      RECT  309.725000  0.765000  310.360000 1.245000 ;
      RECT  309.900000  1.595000  310.090000 1.890000 ;
      RECT  310.350000  0.085000  310.680000 0.580000 ;
      RECT  310.400000  1.790000  310.615000 2.635000 ;
      RECT  310.530000  0.995000  310.760000 1.425000 ;
      RECT  310.865000  1.795000  311.330000 2.465000 ;
      RECT  310.905000  0.255000  311.310000 0.715000 ;
      RECT  310.980000  0.715000  311.310000 0.925000 ;
      RECT  310.980000  0.925000  311.780000 1.445000 ;
      RECT  310.980000  1.445000  311.330000 1.795000 ;
      RECT  311.500000  0.085000  311.765000 0.745000 ;
      RECT  311.500000  1.625000  311.765000 2.635000 ;
      RECT  311.965000  0.085000  312.255000 0.810000 ;
      RECT  311.965000  1.470000  312.255000 2.635000 ;
      RECT  312.490000  0.255000  312.975000 0.355000 ;
      RECT  312.490000  0.355000  314.040000 0.545000 ;
      RECT  312.490000  0.545000  312.975000 0.805000 ;
      RECT  312.490000  0.805000  312.710000 1.495000 ;
      RECT  312.490000  1.495000  312.850000 2.165000 ;
      RECT  312.880000  0.995000  313.205000 1.325000 ;
      RECT  313.020000  1.325000  313.205000 1.875000 ;
      RECT  313.020000  1.875000  317.245000 2.105000 ;
      RECT  313.070000  2.275000  313.570000 2.635000 ;
      RECT  313.375000  0.725000  313.625000 1.340000 ;
      RECT  313.670000  1.525000  314.545000 1.695000 ;
      RECT  313.830000  0.995000  314.205000 1.340000 ;
      RECT  313.860000  0.545000  314.040000 0.615000 ;
      RECT  313.860000  0.615000  314.605000 0.805000 ;
      RECT  314.235000  2.275000  314.565000 2.635000 ;
      RECT  314.270000  0.085000  314.600000 0.445000 ;
      RECT  314.375000  0.805000  314.605000 1.020000 ;
      RECT  314.375000  1.020000  315.740000 1.355000 ;
      RECT  314.375000  1.355000  314.545000 1.525000 ;
      RECT  314.715000  1.535000  316.335000 1.705000 ;
      RECT  314.825000  0.515000  315.015000 0.615000 ;
      RECT  314.825000  0.615000  316.335000 0.845000 ;
      RECT  315.185000  0.085000  315.535000 0.445000 ;
      RECT  315.185000  2.275000  315.570000 2.635000 ;
      RECT  315.705000  0.255000  315.975000 0.615000 ;
      RECT  315.910000  0.845000  316.335000 1.535000 ;
      RECT  316.145000  0.085000  316.525000 0.445000 ;
      RECT  316.145000  2.275000  316.525000 2.635000 ;
      RECT  316.505000  0.615000  316.795000 1.705000 ;
      RECT  316.965000  0.425000  317.245000 1.875000 ;
      RECT  317.485000  0.085000  317.775000 0.810000 ;
      RECT  317.485000  1.470000  317.775000 2.635000 ;
      RECT  317.945000  0.765000  318.185000 2.075000 ;
      RECT  317.950000  2.255000  318.285000 2.635000 ;
      RECT  318.030000  0.255000  318.545000 0.585000 ;
      RECT  318.355000  0.585000  318.545000 1.495000 ;
      RECT  318.355000  1.495000  320.395000 1.665000 ;
      RECT  318.465000  1.665000  318.715000 2.465000 ;
      RECT  318.715000  0.360000  319.095000 1.325000 ;
      RECT  318.895000  1.915000  319.225000 2.635000 ;
      RECT  319.265000  0.355000  319.555000 1.325000 ;
      RECT  319.420000  1.665000  319.670000 2.465000 ;
      RECT  319.745000  0.715000  320.025000 1.325000 ;
      RECT  319.865000  1.835000  320.235000 2.635000 ;
      RECT  319.925000  0.085000  320.195000 0.545000 ;
      RECT  320.195000  0.995000  320.395000 1.495000 ;
      RECT  320.555000  0.295000  320.945000 0.805000 ;
      RECT  320.555000  2.205000  320.945000 2.465000 ;
      RECT  320.685000  0.805000  320.945000 2.205000 ;
      RECT  321.165000  0.085000  321.455000 0.810000 ;
      RECT  321.165000  1.470000  321.455000 2.635000 ;
      RECT  321.635000  2.255000  321.965000 2.635000 ;
      RECT  321.665000  0.755000  321.870000 2.075000 ;
      RECT  321.715000  0.255000  322.210000 0.585000 ;
      RECT  322.040000  0.585000  322.210000 1.495000 ;
      RECT  322.040000  1.495000  324.205000 1.665000 ;
      RECT  322.185000  1.665000  322.355000 2.465000 ;
      RECT  322.395000  0.420000  322.775000 1.325000 ;
      RECT  322.575000  1.915000  322.905000 2.635000 ;
      RECT  322.945000  0.415000  323.245000 1.325000 ;
      RECT  323.110000  1.665000  323.360000 2.465000 ;
      RECT  323.425000  0.740000  323.695000 1.325000 ;
      RECT  323.705000  1.835000  323.955000 2.635000 ;
      RECT  323.825000  0.085000  323.995000 0.550000 ;
      RECT  324.035000  0.995000  324.205000 1.495000 ;
      RECT  324.165000  0.295000  324.615000 0.805000 ;
      RECT  324.165000  1.835000  324.615000 2.465000 ;
      RECT  324.375000  0.805000  324.615000 1.835000 ;
      RECT  324.785000  0.085000  325.115000 0.810000 ;
      RECT  324.785000  1.835000  325.105000 2.635000 ;
      RECT  325.305000  0.085000  325.595000 0.810000 ;
      RECT  325.305000  1.470000  325.595000 2.635000 ;
      RECT  325.785000  1.835000  326.065000 2.635000 ;
      RECT  325.805000  0.765000  326.010000 1.655000 ;
      RECT  325.855000  0.255000  326.400000 0.585000 ;
      RECT  326.180000  0.585000  326.400000 1.495000 ;
      RECT  326.180000  1.495000  328.295000 1.665000 ;
      RECT  326.285000  1.665000  326.495000 2.465000 ;
      RECT  326.570000  0.420000  327.025000 1.325000 ;
      RECT  326.735000  1.935000  327.065000 2.635000 ;
      RECT  327.195000  0.425000  327.460000 1.325000 ;
      RECT  327.285000  1.665000  327.475000 2.465000 ;
      RECT  327.665000  0.730000  327.955000 1.325000 ;
      RECT  327.905000  0.085000  328.215000 0.550000 ;
      RECT  327.905000  1.855000  328.235000 2.635000 ;
      RECT  328.125000  1.075000  329.615000 1.305000 ;
      RECT  328.125000  1.305000  328.295000 1.495000 ;
      RECT  328.465000  0.255000  328.635000 0.640000 ;
      RECT  328.465000  0.640000  330.135000 0.810000 ;
      RECT  328.465000  1.485000  330.135000 1.655000 ;
      RECT  328.465000  1.655000  328.715000 2.465000 ;
      RECT  328.805000  0.085000  329.185000 0.470000 ;
      RECT  328.935000  1.835000  329.185000 2.635000 ;
      RECT  329.405000  0.255000  329.575000 0.640000 ;
      RECT  329.405000  1.655000  330.135000 1.745000 ;
      RECT  329.405000  1.745000  329.575000 2.465000 ;
      RECT  329.745000  0.085000  330.125000 0.470000 ;
      RECT  329.745000  1.915000  330.125000 2.635000 ;
      RECT  329.880000  0.810000  330.135000 1.485000 ;
      RECT  330.365000  0.085000  330.655000 0.810000 ;
      RECT  330.365000  1.470000  330.655000 2.635000 ;
      RECT  330.825000  0.995000  331.190000 1.675000 ;
      RECT  330.910000  0.255000  331.085000 0.655000 ;
      RECT  330.910000  0.655000  331.590000 0.825000 ;
      RECT  330.910000  1.845000  331.590000 2.015000 ;
      RECT  330.910000  2.015000  331.085000 2.465000 ;
      RECT  331.255000  0.085000  331.635000 0.465000 ;
      RECT  331.255000  2.195000  331.635000 2.635000 ;
      RECT  331.420000  0.825000  331.590000 0.995000 ;
      RECT  331.420000  0.995000  331.765000 1.325000 ;
      RECT  331.420000  1.325000  331.590000 1.845000 ;
      RECT  331.880000  0.255000  332.110000 0.585000 ;
      RECT  331.940000  0.585000  332.110000 1.875000 ;
      RECT  331.940000  1.875000  334.155000 2.045000 ;
      RECT  331.940000  2.045000  332.110000 2.465000 ;
      RECT  332.395000  2.225000  333.115000 2.635000 ;
      RECT  332.415000  0.420000  332.895000 1.695000 ;
      RECT  333.065000  0.420000  333.355000 1.695000 ;
      RECT  333.370000  2.045000  333.540000 2.465000 ;
      RECT  333.525000  0.665000  333.815000 1.695000 ;
      RECT  333.695000  0.085000  334.090000 0.465000 ;
      RECT  333.800000  2.225000  334.130000 2.635000 ;
      RECT  333.985000  0.995000  334.275000 1.325000 ;
      RECT  333.985000  1.325000  334.155000 1.875000 ;
      RECT  334.260000  0.295000  334.735000 0.805000 ;
      RECT  334.375000  1.495000  334.735000 2.465000 ;
      RECT  334.465000  0.805000  334.735000 1.495000 ;
      RECT  334.965000  0.085000  335.255000 0.810000 ;
      RECT  334.965000  1.470000  335.255000 2.635000 ;
      RECT  335.435000  0.085000  335.765000 0.465000 ;
      RECT  335.475000  0.740000  335.675000 1.630000 ;
      RECT  335.515000  1.830000  336.195000 2.000000 ;
      RECT  335.515000  2.000000  335.685000 2.465000 ;
      RECT  335.855000  2.195000  336.235000 2.635000 ;
      RECT  335.985000  0.255000  336.195000 0.585000 ;
      RECT  336.025000  0.585000  336.195000 0.995000 ;
      RECT  336.025000  0.995000  336.415000 1.325000 ;
      RECT  336.025000  1.325000  336.195000 1.830000 ;
      RECT  336.455000  1.660000  336.755000 1.915000 ;
      RECT  336.455000  1.915000  338.805000 1.965000 ;
      RECT  336.455000  1.965000  338.200000 2.085000 ;
      RECT  336.455000  2.085000  336.625000 2.465000 ;
      RECT  336.535000  0.255000  336.755000 0.585000 ;
      RECT  336.585000  0.585000  336.755000 1.660000 ;
      RECT  337.045000  2.255000  337.765000 2.635000 ;
      RECT  337.235000  0.420000  337.495000 1.745000 ;
      RECT  337.715000  0.420000  337.955000 1.615000 ;
      RECT  338.010000  2.085000  338.200000 2.465000 ;
      RECT  338.030000  1.795000  338.805000 1.915000 ;
      RECT  338.125000  0.645000  338.455000 1.615000 ;
      RECT  338.350000  0.085000  338.730000 0.465000 ;
      RECT  338.480000  2.195000  338.810000 2.635000 ;
      RECT  338.635000  0.995000  338.895000 1.325000 ;
      RECT  338.635000  1.325000  338.805000 1.795000 ;
      RECT  338.900000  0.255000  339.235000 0.640000 ;
      RECT  338.900000  0.640000  339.795000 0.825000 ;
      RECT  339.030000  1.535000  339.795000 1.665000 ;
      RECT  339.030000  1.665000  339.335000 2.465000 ;
      RECT  339.115000  0.825000  339.795000 1.535000 ;
      RECT  339.405000  0.085000  339.790000 0.465000 ;
      RECT  339.535000  1.835000  339.790000 2.635000 ;
      RECT  340.025000  0.085000  340.315000 0.810000 ;
      RECT  340.025000  1.470000  340.315000 2.635000 ;
      RECT  340.485000  0.255000  340.745000 0.585000 ;
      RECT  340.485000  0.585000  340.660000 1.915000 ;
      RECT  340.485000  1.915000  345.285000 2.085000 ;
      RECT  340.485000  2.085000  340.745000 2.465000 ;
      RECT  340.840000  0.765000  341.240000 1.635000 ;
      RECT  340.915000  2.255000  341.295000 2.635000 ;
      RECT  340.965000  0.085000  341.215000 0.545000 ;
      RECT  341.430000  0.255000  341.740000 0.650000 ;
      RECT  341.430000  0.650000  342.680000 0.820000 ;
      RECT  341.430000  0.820000  341.760000 1.545000 ;
      RECT  341.430000  1.545000  342.760000 1.715000 ;
      RECT  341.910000  0.085000  342.290000 0.470000 ;
      RECT  341.910000  2.255000  342.290000 2.635000 ;
      RECT  341.930000  0.995000  343.100000 1.325000 ;
      RECT  342.510000  0.255000  342.680000 0.650000 ;
      RECT  342.850000  2.255000  343.230000 2.635000 ;
      RECT  342.930000  1.325000  343.100000 1.545000 ;
      RECT  342.930000  1.545000  344.930000 1.715000 ;
      RECT  342.935000  0.085000  343.265000 0.445000 ;
      RECT  343.270000  0.995000  343.520000 1.325000 ;
      RECT  343.730000  0.755000  344.040000 1.325000 ;
      RECT  343.910000  2.255000  344.290000 2.635000 ;
      RECT  344.210000  0.735000  344.590000 1.325000 ;
      RECT  344.760000  0.640000  345.300000 0.810000 ;
      RECT  344.760000  0.810000  344.930000 1.545000 ;
      RECT  344.970000  2.255000  345.350000 2.635000 ;
      RECT  345.115000  0.995000  345.285000 1.915000 ;
      RECT  345.545000  0.085000  345.835000 0.810000 ;
      RECT  345.545000  1.470000  345.835000 2.635000 ;
      RECT  346.005000  0.255000  346.265000 0.585000 ;
      RECT  346.005000  0.585000  346.175000 1.285000 ;
      RECT  346.005000  1.285000  347.155000 1.455000 ;
      RECT  346.005000  1.455000  346.175000 2.135000 ;
      RECT  346.005000  2.135000  346.265000 2.465000 ;
      RECT  346.345000  1.625000  346.735000 1.955000 ;
      RECT  346.445000  0.765000  346.705000 0.945000 ;
      RECT  346.445000  0.945000  347.085000 1.115000 ;
      RECT  346.495000  0.085000  346.875000 0.465000 ;
      RECT  346.495000  2.255000  346.875000 2.635000 ;
      RECT  346.935000  1.455000  347.155000 1.575000 ;
      RECT  346.935000  1.575000  347.565000 1.745000 ;
      RECT  347.085000  1.915000  347.905000 2.085000 ;
      RECT  347.085000  2.085000  347.295000 2.465000 ;
      RECT  347.105000  0.255000  348.585000 0.425000 ;
      RECT  347.105000  0.425000  347.505000 0.755000 ;
      RECT  347.335000  0.755000  347.505000 1.235000 ;
      RECT  347.335000  1.235000  347.905000 1.405000 ;
      RECT  347.545000  2.255000  347.875000 2.635000 ;
      RECT  347.675000  0.595000  348.245000 0.925000 ;
      RECT  347.735000  1.405000  347.905000 1.915000 ;
      RECT  348.075000  0.925000  348.245000 1.915000 ;
      RECT  348.075000  1.915000  349.900000 2.085000 ;
      RECT  348.105000  2.085000  348.275000 2.465000 ;
      RECT  348.415000  0.425000  348.585000 1.325000 ;
      RECT  348.470000  2.255000  348.850000 2.635000 ;
      RECT  348.795000  0.415000  349.095000 1.635000 ;
      RECT  349.130000  2.085000  349.300000 2.465000 ;
      RECT  349.265000  0.420000  349.560000 1.635000 ;
      RECT  349.620000  2.255000  349.950000 2.635000 ;
      RECT  349.730000  0.085000  349.900000 0.545000 ;
      RECT  349.730000  0.995000  350.035000 1.325000 ;
      RECT  349.730000  1.325000  349.900000 1.915000 ;
      RECT  350.170000  0.255000  350.430000 0.825000 ;
      RECT  350.170000  1.445000  350.430000 2.465000 ;
      RECT  350.205000  0.825000  350.430000 1.445000 ;
      RECT  350.605000  0.085000  350.895000 0.810000 ;
      RECT  350.605000  1.470000  350.895000 2.635000 ;
      RECT  351.130000  0.995000  351.310000 1.635000 ;
      RECT  351.155000  0.255000  351.325000 0.635000 ;
      RECT  351.155000  0.635000  351.700000 0.805000 ;
      RECT  351.155000  1.885000  353.055000 2.055000 ;
      RECT  351.155000  2.055000  351.325000 2.465000 ;
      RECT  351.480000  0.805000  351.700000 1.885000 ;
      RECT  351.495000  0.085000  351.875000 0.465000 ;
      RECT  351.495000  2.255000  351.875000 2.635000 ;
      RECT  352.045000  0.255000  352.320000 1.545000 ;
      RECT  352.045000  1.545000  352.400000 1.715000 ;
      RECT  352.490000  0.085000  352.870000 0.465000 ;
      RECT  352.495000  0.635000  353.585000 0.805000 ;
      RECT  352.495000  0.805000  352.715000 1.325000 ;
      RECT  352.620000  2.255000  353.290000 2.635000 ;
      RECT  352.885000  0.995000  353.195000 1.325000 ;
      RECT  352.885000  1.325000  353.055000 1.885000 ;
      RECT  353.125000  0.255000  353.295000 0.635000 ;
      RECT  353.365000  0.805000  353.585000 1.915000 ;
      RECT  353.365000  1.915000  354.695000 2.085000 ;
      RECT  353.575000  2.085000  353.745000 2.465000 ;
      RECT  353.775000  1.400000  353.995000 1.575000 ;
      RECT  353.775000  1.575000  355.085000 1.745000 ;
      RECT  353.915000  2.255000  354.305000 2.635000 ;
      RECT  354.250000  0.420000  354.515000 1.275000 ;
      RECT  354.525000  2.085000  354.695000 2.465000 ;
      RECT  354.685000  0.425000  354.985000 1.405000 ;
      RECT  354.865000  1.745000  355.085000 1.915000 ;
      RECT  354.865000  1.915000  355.895000 2.085000 ;
      RECT  355.085000  2.255000  355.415000 2.635000 ;
      RECT  355.155000  0.765000  355.505000 1.305000 ;
      RECT  355.165000  0.085000  355.415000 0.585000 ;
      RECT  355.635000  0.255000  355.895000 0.585000 ;
      RECT  355.635000  2.085000  355.895000 2.465000 ;
      RECT  355.725000  0.585000  355.895000 1.915000 ;
      RECT  356.125000  0.085000  356.415000 0.810000 ;
      RECT  356.125000  1.470000  356.415000 2.635000 ;
      RECT  356.585000  0.255000  356.845000 0.585000 ;
      RECT  356.585000  0.585000  356.760000 1.915000 ;
      RECT  356.585000  1.915000  361.440000 2.085000 ;
      RECT  356.585000  2.085000  356.845000 2.465000 ;
      RECT  356.930000  0.765000  357.330000 1.635000 ;
      RECT  357.015000  2.255000  357.395000 2.635000 ;
      RECT  357.120000  0.085000  357.450000 0.470000 ;
      RECT  357.510000  0.650000  358.780000 0.820000 ;
      RECT  357.510000  0.820000  357.840000 1.545000 ;
      RECT  357.510000  1.545000  358.860000 1.715000 ;
      RECT  357.670000  0.255000  357.840000 0.650000 ;
      RECT  358.010000  0.085000  358.390000 0.470000 ;
      RECT  358.010000  1.075000  359.200000 1.245000 ;
      RECT  358.010000  2.255000  358.390000 2.635000 ;
      RECT  358.610000  0.255000  358.780000 0.650000 ;
      RECT  358.950000  2.255000  359.330000 2.635000 ;
      RECT  358.970000  0.085000  359.300000 0.445000 ;
      RECT  359.030000  0.615000  359.695000 0.785000 ;
      RECT  359.030000  0.785000  359.200000 1.075000 ;
      RECT  359.030000  1.245000  359.200000 1.545000 ;
      RECT  359.030000  1.545000  361.050000 1.715000 ;
      RECT  359.405000  0.995000  359.695000 1.325000 ;
      RECT  359.475000  0.300000  361.560000 0.470000 ;
      RECT  359.475000  0.470000  359.695000 0.615000 ;
      RECT  359.865000  0.640000  360.340000 1.325000 ;
      RECT  360.180000  2.255000  360.510000 2.635000 ;
      RECT  360.580000  0.995000  360.800000 1.205000 ;
      RECT  360.580000  1.205000  361.440000 1.375000 ;
      RECT  361.210000  0.470000  361.560000 0.810000 ;
      RECT  361.270000  1.375000  361.440000 1.915000 ;
      RECT  361.310000  2.255000  362.320000 2.635000 ;
      RECT  361.860000  0.655000  362.765000 0.825000 ;
      RECT  361.860000  0.825000  362.030000 1.915000 ;
      RECT  361.860000  1.915000  362.765000 2.085000 ;
      RECT  361.885000  0.085000  362.215000 0.465000 ;
      RECT  362.435000  0.995000  362.845000 1.620000 ;
      RECT  362.595000  0.255000  362.765000 0.655000 ;
      RECT  362.595000  2.085000  362.765000 2.465000 ;
      RECT  363.025000  0.085000  363.315000 0.810000 ;
      RECT  363.025000  1.470000  363.315000 2.635000 ;
      RECT  363.505000  0.985000  363.945000 1.355000 ;
      RECT  363.565000  1.535000  364.290000 1.705000 ;
      RECT  363.565000  1.705000  363.745000 2.465000 ;
      RECT  363.575000  0.255000  363.745000 0.635000 ;
      RECT  363.575000  0.635000  364.290000 0.805000 ;
      RECT  363.925000  0.085000  364.295000 0.465000 ;
      RECT  363.925000  1.875000  364.295000 2.635000 ;
      RECT  364.120000  0.805000  364.290000 1.060000 ;
      RECT  364.120000  1.060000  364.435000 1.390000 ;
      RECT  364.120000  1.390000  364.290000 1.535000 ;
      RECT  364.465000  0.255000  364.795000 0.760000 ;
      RECT  364.465000  1.560000  364.795000 2.465000 ;
      RECT  364.615000  0.760000  364.795000 1.560000 ;
      RECT  365.325000  0.085000  365.615000 0.810000 ;
      RECT  365.325000  1.470000  365.615000 2.635000 ;
      RECT  365.795000  0.085000  366.125000 0.565000 ;
      RECT  365.835000  1.075000  367.510000 1.275000 ;
      RECT  365.875000  1.835000  366.045000 2.635000 ;
      RECT  366.215000  1.445000  367.915000 1.615000 ;
      RECT  366.215000  1.615000  366.595000 2.465000 ;
      RECT  366.345000  0.255000  366.515000 0.735000 ;
      RECT  366.345000  0.735000  367.915000 0.905000 ;
      RECT  366.685000  0.085000  367.065000 0.565000 ;
      RECT  366.815000  1.835000  366.985000 2.635000 ;
      RECT  367.155000  1.615000  367.535000 2.465000 ;
      RECT  367.285000  0.260000  367.455000 0.735000 ;
      RECT  367.625000  0.085000  368.005000 0.565000 ;
      RECT  367.740000  0.905000  367.915000 1.075000 ;
      RECT  367.740000  1.075000  370.665000 1.245000 ;
      RECT  367.740000  1.245000  367.915000 1.445000 ;
      RECT  367.755000  1.835000  367.925000 2.635000 ;
      RECT  368.225000  0.255000  368.395000 0.735000 ;
      RECT  368.225000  0.735000  373.095000 0.905000 ;
      RECT  368.225000  1.445000  373.095000 1.615000 ;
      RECT  368.225000  1.615000  368.395000 2.465000 ;
      RECT  368.565000  0.085000  368.945000 0.565000 ;
      RECT  368.565000  1.835000  368.945000 2.635000 ;
      RECT  369.165000  0.255000  369.335000 0.735000 ;
      RECT  369.165000  1.615000  369.335000 2.465000 ;
      RECT  369.505000  0.085000  369.885000 0.565000 ;
      RECT  369.505000  1.835000  369.885000 2.635000 ;
      RECT  370.105000  0.255000  370.275000 0.735000 ;
      RECT  370.105000  1.615000  370.275000 2.465000 ;
      RECT  370.445000  0.085000  370.825000 0.565000 ;
      RECT  370.445000  1.835000  370.825000 2.635000 ;
      RECT  370.910000  0.905000  373.095000 1.445000 ;
      RECT  371.045000  0.255000  371.215000 0.735000 ;
      RECT  371.045000  1.615000  371.215000 2.465000 ;
      RECT  371.385000  0.085000  371.765000 0.565000 ;
      RECT  371.385000  1.835000  371.765000 2.635000 ;
      RECT  371.985000  0.255000  372.155000 0.735000 ;
      RECT  371.985000  1.615000  372.155000 2.465000 ;
      RECT  372.325000  0.085000  372.705000 0.565000 ;
      RECT  372.325000  1.835000  372.705000 2.635000 ;
      RECT  372.925000  0.255000  373.095000 0.735000 ;
      RECT  372.925000  1.615000  373.095000 2.465000 ;
      RECT  373.265000  0.085000  373.645000 0.885000 ;
      RECT  373.265000  1.485000  373.645000 2.635000 ;
      RECT  374.065000  0.085000  374.355000 0.810000 ;
      RECT  374.065000  1.470000  374.355000 2.635000 ;
      RECT  374.525000  1.075000  377.175000 1.275000 ;
      RECT  374.615000  0.085000  374.785000 0.905000 ;
      RECT  374.615000  1.445000  374.785000 2.635000 ;
      RECT  374.955000  0.260000  375.335000 0.735000 ;
      RECT  374.955000  0.735000  377.605000 0.905000 ;
      RECT  374.955000  1.445000  377.605000 1.615000 ;
      RECT  374.955000  1.615000  375.335000 2.465000 ;
      RECT  375.555000  0.085000  375.725000 0.565000 ;
      RECT  375.555000  1.835000  375.725000 2.635000 ;
      RECT  375.895000  0.260000  376.275000 0.735000 ;
      RECT  375.895000  1.615000  376.275000 2.465000 ;
      RECT  376.495000  0.085000  376.665000 0.565000 ;
      RECT  376.495000  1.835000  376.665000 2.635000 ;
      RECT  376.835000  0.260000  377.215000 0.735000 ;
      RECT  376.835000  1.615000  377.215000 2.465000 ;
      RECT  377.430000  0.905000  377.605000 1.075000 ;
      RECT  377.430000  1.075000  384.615000 1.275000 ;
      RECT  377.430000  1.275000  377.605000 1.445000 ;
      RECT  377.435000  0.085000  377.605000 0.565000 ;
      RECT  377.435000  1.835000  377.605000 2.635000 ;
      RECT  377.775000  0.255000  378.075000 0.260000 ;
      RECT  377.775000  0.260000  378.155000 0.735000 ;
      RECT  377.775000  0.735000  385.575000 0.905000 ;
      RECT  377.775000  1.445000  385.575000 1.615000 ;
      RECT  377.775000  1.615000  378.155000 2.465000 ;
      RECT  378.375000  0.085000  378.545000 0.565000 ;
      RECT  378.375000  1.835000  378.545000 2.635000 ;
      RECT  378.715000  0.260000  379.095000 0.735000 ;
      RECT  378.715000  1.615000  379.095000 2.465000 ;
      RECT  378.845000  0.255000  379.015000 0.260000 ;
      RECT  379.315000  0.085000  379.485000 0.565000 ;
      RECT  379.315000  1.835000  379.485000 2.635000 ;
      RECT  379.655000  0.260000  380.035000 0.735000 ;
      RECT  379.655000  1.615000  380.035000 2.465000 ;
      RECT  379.785000  0.255000  379.955000 0.260000 ;
      RECT  380.255000  0.085000  380.425000 0.565000 ;
      RECT  380.255000  1.835000  380.425000 2.635000 ;
      RECT  380.595000  0.260000  380.975000 0.735000 ;
      RECT  380.595000  1.615000  380.975000 2.465000 ;
      RECT  381.195000  0.085000  381.365000 0.565000 ;
      RECT  381.195000  1.835000  381.365000 2.635000 ;
      RECT  381.535000  0.260000  381.915000 0.735000 ;
      RECT  381.535000  1.615000  381.915000 2.465000 ;
      RECT  382.135000  0.085000  382.305000 0.565000 ;
      RECT  382.135000  1.835000  382.305000 2.635000 ;
      RECT  382.475000  0.260000  382.855000 0.735000 ;
      RECT  382.475000  1.615000  382.855000 2.465000 ;
      RECT  383.075000  0.085000  383.245000 0.565000 ;
      RECT  383.075000  1.835000  383.245000 2.635000 ;
      RECT  383.415000  0.260000  383.795000 0.735000 ;
      RECT  383.415000  1.615000  383.795000 2.465000 ;
      RECT  384.015000  0.085000  384.185000 0.565000 ;
      RECT  384.015000  1.835000  384.185000 2.635000 ;
      RECT  384.355000  0.260000  384.735000 0.735000 ;
      RECT  384.355000  1.615000  384.735000 2.465000 ;
      RECT  384.955000  0.085000  385.125000 0.565000 ;
      RECT  384.955000  1.835000  385.125000 2.635000 ;
      RECT  385.075000  0.905000  385.575000 1.445000 ;
      RECT  385.300000  0.365000  385.575000 0.735000 ;
      RECT  385.300000  1.615000  385.575000 2.360000 ;
      RECT  386.025000  0.085000  386.315000 0.810000 ;
      RECT  386.025000  1.470000  386.315000 2.635000 ;
      RECT  386.485000  0.985000  386.840000 1.355000 ;
      RECT  386.575000  0.255000  386.745000 0.635000 ;
      RECT  386.575000  0.635000  387.340000 0.805000 ;
      RECT  386.575000  1.535000  387.295000 1.705000 ;
      RECT  386.575000  1.705000  386.745000 2.465000 ;
      RECT  387.000000  1.875000  387.330000 2.635000 ;
      RECT  387.010000  0.085000  387.340000 0.465000 ;
      RECT  387.125000  0.805000  387.340000 0.995000 ;
      RECT  387.125000  0.995000  387.425000 1.325000 ;
      RECT  387.125000  1.325000  387.295000 1.535000 ;
      RECT  387.670000  0.255000  388.095000 2.465000 ;
      RECT  388.265000  0.085000  388.525000 0.925000 ;
      RECT  388.265000  1.485000  388.525000 2.635000 ;
      RECT  388.785000  0.085000  389.075000 0.810000 ;
      RECT  388.785000  1.470000  389.075000 2.635000 ;
      RECT  389.250000  1.075000  389.630000 1.315000 ;
      RECT  389.255000  1.485000  390.020000 1.655000 ;
      RECT  389.255000  1.655000  389.585000 2.465000 ;
      RECT  389.335000  0.255000  389.505000 0.735000 ;
      RECT  389.335000  0.735000  390.020000 0.905000 ;
      RECT  389.685000  0.085000  389.975000 0.565000 ;
      RECT  389.805000  1.835000  390.045000 2.635000 ;
      RECT  389.850000  0.905000  390.020000 1.075000 ;
      RECT  389.850000  1.075000  390.400000 1.245000 ;
      RECT  389.850000  1.245000  390.020000 1.485000 ;
      RECT  390.275000  0.255000  390.445000 0.735000 ;
      RECT  390.275000  0.735000  391.385000 0.905000 ;
      RECT  390.275000  1.445000  391.385000 1.615000 ;
      RECT  390.275000  1.615000  390.445000 2.465000 ;
      RECT  390.615000  0.085000  390.995000 0.565000 ;
      RECT  390.615000  1.835000  390.995000 2.635000 ;
      RECT  391.080000  0.905000  391.385000 1.445000 ;
      RECT  391.215000  0.255000  391.385000 0.735000 ;
      RECT  391.215000  1.615000  391.385000 2.465000 ;
      RECT  391.555000  0.085000  391.935000 0.885000 ;
      RECT  391.555000  1.485000  391.935000 2.635000 ;
      RECT  392.465000  0.085000  392.755000 0.810000 ;
      RECT  392.465000  1.470000  392.755000 2.635000 ;
      RECT  393.120000  1.075000  394.105000 1.315000 ;
      RECT  393.275000  0.085000  393.445000 0.565000 ;
      RECT  393.275000  1.485000  393.445000 2.635000 ;
      RECT  393.615000  0.255000  393.995000 0.735000 ;
      RECT  393.615000  0.735000  394.465000 0.905000 ;
      RECT  393.615000  1.485000  394.465000 1.655000 ;
      RECT  393.615000  1.655000  393.995000 2.465000 ;
      RECT  394.215000  0.085000  394.385000 0.565000 ;
      RECT  394.215000  1.835000  394.455000 2.635000 ;
      RECT  394.295000  0.905000  394.465000 1.075000 ;
      RECT  394.295000  1.075000  394.815000 1.245000 ;
      RECT  394.295000  1.245000  394.465000 1.485000 ;
      RECT  394.685000  0.255000  394.855000 0.735000 ;
      RECT  394.685000  0.735000  396.735000 0.905000 ;
      RECT  394.685000  1.445000  396.735000 1.615000 ;
      RECT  394.685000  1.615000  394.855000 2.465000 ;
      RECT  395.025000  0.085000  395.405000 0.565000 ;
      RECT  395.025000  1.835000  395.405000 2.635000 ;
      RECT  395.250000  0.905000  396.735000 1.445000 ;
      RECT  395.625000  0.255000  395.795000 0.735000 ;
      RECT  395.625000  1.615000  395.795000 2.465000 ;
      RECT  395.965000  0.085000  396.345000 0.565000 ;
      RECT  395.965000  1.835000  396.345000 2.635000 ;
      RECT  396.565000  0.255000  396.735000 0.735000 ;
      RECT  396.565000  1.615000  396.735000 2.465000 ;
      RECT  396.905000  0.085000  397.285000 0.885000 ;
      RECT  396.905000  1.485000  397.285000 2.635000 ;
      RECT  397.525000  0.085000  397.815000 0.810000 ;
      RECT  397.525000  1.470000  397.815000 2.635000 ;
      RECT  397.995000  1.445000  399.645000 1.615000 ;
      RECT  397.995000  1.615000  398.325000 2.465000 ;
      RECT  398.040000  1.075000  399.240000 1.275000 ;
      RECT  398.075000  0.255000  398.245000 0.735000 ;
      RECT  398.075000  0.735000  399.645000 0.905000 ;
      RECT  398.415000  0.085000  398.795000 0.565000 ;
      RECT  398.545000  1.835000  398.715000 2.635000 ;
      RECT  398.885000  1.615000  399.265000 2.465000 ;
      RECT  399.015000  0.260000  399.185000 0.735000 ;
      RECT  399.355000  0.085000  399.735000 0.565000 ;
      RECT  399.470000  0.905000  399.645000 1.075000 ;
      RECT  399.470000  1.075000  402.395000 1.245000 ;
      RECT  399.470000  1.245000  399.645000 1.445000 ;
      RECT  399.485000  1.835000  399.655000 2.635000 ;
      RECT  399.955000  0.255000  400.125000 0.735000 ;
      RECT  399.955000  0.735000  402.945000 0.905000 ;
      RECT  399.955000  1.445000  402.945000 1.615000 ;
      RECT  399.955000  1.615000  400.125000 2.465000 ;
      RECT  400.295000  0.085000  400.675000 0.565000 ;
      RECT  400.295000  1.835000  400.675000 2.635000 ;
      RECT  400.895000  0.255000  401.065000 0.735000 ;
      RECT  400.895000  1.615000  401.065000 2.465000 ;
      RECT  401.235000  0.085000  401.615000 0.565000 ;
      RECT  401.235000  1.835000  401.615000 2.635000 ;
      RECT  401.835000  0.255000  402.005000 0.735000 ;
      RECT  401.835000  1.615000  402.005000 2.465000 ;
      RECT  402.175000  0.085000  402.555000 0.565000 ;
      RECT  402.175000  1.835000  402.555000 2.635000 ;
      RECT  402.590000  0.905000  402.945000 1.445000 ;
      RECT  402.775000  0.255000  402.945000 0.735000 ;
      RECT  402.775000  1.615000  402.945000 2.465000 ;
      RECT  403.115000  0.085000  403.495000 0.885000 ;
      RECT  403.115000  1.485000  403.495000 2.635000 ;
      RECT  403.965000  0.085000  404.255000 0.810000 ;
      RECT  403.965000  1.470000  404.255000 2.635000 ;
      RECT  404.450000  1.075000  404.780000 1.275000 ;
      RECT  404.515000  0.085000  404.685000 0.905000 ;
      RECT  404.515000  1.445000  404.685000 2.635000 ;
      RECT  404.855000  0.260000  405.235000 0.905000 ;
      RECT  404.855000  1.445000  405.235000 2.465000 ;
      RECT  405.000000  0.905000  405.235000 1.075000 ;
      RECT  405.000000  1.075000  406.695000 1.275000 ;
      RECT  405.000000  1.275000  405.235000 1.445000 ;
      RECT  405.425000  0.260000  405.755000 0.735000 ;
      RECT  405.425000  0.735000  407.085000 0.905000 ;
      RECT  405.425000  1.445000  407.085000 1.615000 ;
      RECT  405.425000  1.615000  405.755000 2.465000 ;
      RECT  405.975000  0.085000  406.145000 0.565000 ;
      RECT  405.975000  1.785000  406.145000 2.635000 ;
      RECT  406.315000  0.260000  406.695000 0.735000 ;
      RECT  406.315000  1.615000  406.695000 2.465000 ;
      RECT  406.915000  0.085000  407.085000 0.565000 ;
      RECT  406.915000  0.905000  407.085000 1.075000 ;
      RECT  406.915000  1.075000  409.475000 1.275000 ;
      RECT  406.915000  1.275000  407.085000 1.445000 ;
      RECT  406.915000  1.785000  407.085000 2.635000 ;
      RECT  407.255000  0.260000  407.635000 0.735000 ;
      RECT  407.255000  0.735000  409.905000 0.905000 ;
      RECT  407.255000  1.445000  409.905000 1.615000 ;
      RECT  407.255000  1.615000  407.635000 2.465000 ;
      RECT  407.855000  0.085000  408.025000 0.565000 ;
      RECT  407.855000  1.835000  408.025000 2.635000 ;
      RECT  408.195000  0.260000  408.575000 0.735000 ;
      RECT  408.195000  1.615000  408.575000 2.465000 ;
      RECT  408.795000  0.085000  408.965000 0.565000 ;
      RECT  408.795000  1.835000  408.965000 2.635000 ;
      RECT  409.135000  0.260000  409.515000 0.735000 ;
      RECT  409.135000  1.615000  409.515000 2.465000 ;
      RECT  409.730000  0.905000  409.905000 1.075000 ;
      RECT  409.730000  1.075000  417.040000 1.275000 ;
      RECT  409.730000  1.275000  409.905000 1.445000 ;
      RECT  409.735000  0.085000  409.905000 0.565000 ;
      RECT  409.735000  1.835000  409.905000 2.635000 ;
      RECT  410.075000  0.255000  410.375000 0.260000 ;
      RECT  410.075000  0.260000  410.455000 0.735000 ;
      RECT  410.075000  0.735000  417.560000 0.905000 ;
      RECT  410.075000  1.445000  417.560000 1.615000 ;
      RECT  410.075000  1.615000  410.455000 2.465000 ;
      RECT  410.675000  0.085000  410.845000 0.565000 ;
      RECT  410.675000  1.835000  410.845000 2.635000 ;
      RECT  411.015000  0.260000  411.395000 0.735000 ;
      RECT  411.015000  1.615000  411.395000 2.465000 ;
      RECT  411.145000  0.255000  411.315000 0.260000 ;
      RECT  411.615000  0.085000  411.785000 0.565000 ;
      RECT  411.615000  1.835000  411.785000 2.635000 ;
      RECT  411.955000  0.260000  412.335000 0.735000 ;
      RECT  411.955000  1.615000  412.335000 2.465000 ;
      RECT  412.085000  0.255000  412.255000 0.260000 ;
      RECT  412.555000  0.085000  412.725000 0.565000 ;
      RECT  412.555000  1.835000  412.725000 2.635000 ;
      RECT  412.895000  0.260000  413.275000 0.735000 ;
      RECT  412.895000  1.615000  413.275000 2.465000 ;
      RECT  413.495000  0.085000  413.665000 0.565000 ;
      RECT  413.495000  1.835000  413.665000 2.635000 ;
      RECT  413.835000  0.260000  414.215000 0.735000 ;
      RECT  413.835000  1.615000  414.215000 2.465000 ;
      RECT  414.435000  0.085000  414.605000 0.565000 ;
      RECT  414.435000  1.835000  414.605000 2.635000 ;
      RECT  414.775000  0.260000  415.155000 0.735000 ;
      RECT  414.775000  1.615000  415.155000 2.465000 ;
      RECT  415.375000  0.085000  415.545000 0.565000 ;
      RECT  415.375000  1.835000  415.545000 2.635000 ;
      RECT  415.715000  0.260000  416.095000 0.735000 ;
      RECT  415.715000  1.615000  416.095000 2.465000 ;
      RECT  416.315000  0.085000  416.485000 0.565000 ;
      RECT  416.315000  1.835000  416.485000 2.635000 ;
      RECT  416.655000  0.260000  417.035000 0.735000 ;
      RECT  416.655000  1.615000  417.035000 2.465000 ;
      RECT  417.255000  0.085000  417.425000 0.565000 ;
      RECT  417.255000  1.835000  417.425000 2.635000 ;
      RECT  417.260000  0.905000  417.560000 1.445000 ;
      RECT  417.765000  0.085000  418.055000 0.810000 ;
      RECT  417.765000  1.470000  418.055000 2.635000 ;
      RECT  418.235000  0.260000  418.565000 0.735000 ;
      RECT  418.235000  0.735000  418.970000 0.905000 ;
      RECT  418.235000  1.445000  418.970000 1.615000 ;
      RECT  418.235000  1.615000  418.565000 2.160000 ;
      RECT  418.250000  1.075000  418.580000 1.275000 ;
      RECT  418.785000  0.085000  418.955000 0.565000 ;
      RECT  418.785000  1.785000  418.955000 2.635000 ;
      RECT  418.800000  0.905000  418.970000 0.995000 ;
      RECT  418.800000  0.995000  419.280000 1.325000 ;
      RECT  418.800000  1.325000  418.970000 1.445000 ;
      RECT  419.190000  0.260000  419.620000 0.825000 ;
      RECT  419.190000  1.545000  419.620000 2.465000 ;
      RECT  419.450000  0.825000  419.620000 1.075000 ;
      RECT  419.450000  1.075000  421.060000 1.275000 ;
      RECT  419.450000  1.275000  419.620000 1.545000 ;
      RECT  419.790000  0.260000  420.120000 0.735000 ;
      RECT  419.790000  0.735000  421.450000 0.905000 ;
      RECT  419.790000  1.445000  421.450000 1.615000 ;
      RECT  419.790000  1.615000  420.120000 2.465000 ;
      RECT  420.340000  0.085000  420.510000 0.565000 ;
      RECT  420.340000  1.785000  420.510000 2.635000 ;
      RECT  420.680000  0.260000  421.060000 0.735000 ;
      RECT  420.680000  1.615000  421.060000 2.465000 ;
      RECT  421.280000  0.085000  421.450000 0.565000 ;
      RECT  421.280000  0.905000  421.450000 1.075000 ;
      RECT  421.280000  1.075000  424.050000 1.275000 ;
      RECT  421.280000  1.275000  421.450000 1.445000 ;
      RECT  421.280000  1.785000  421.450000 2.635000 ;
      RECT  421.620000  0.260000  422.000000 0.735000 ;
      RECT  421.620000  0.735000  425.380000 0.905000 ;
      RECT  421.620000  1.445000  425.380000 1.615000 ;
      RECT  421.620000  1.615000  422.000000 2.465000 ;
      RECT  422.220000  0.085000  422.390000 0.565000 ;
      RECT  422.220000  1.835000  422.390000 2.635000 ;
      RECT  422.560000  0.260000  422.940000 0.735000 ;
      RECT  422.560000  1.615000  422.940000 2.465000 ;
      RECT  423.160000  0.085000  423.330000 0.565000 ;
      RECT  423.160000  1.835000  423.330000 2.635000 ;
      RECT  423.500000  0.260000  423.880000 0.735000 ;
      RECT  423.500000  1.615000  423.880000 2.465000 ;
      RECT  424.100000  0.085000  424.270000 0.565000 ;
      RECT  424.100000  1.835000  424.270000 2.635000 ;
      RECT  424.440000  0.260000  424.820000 0.735000 ;
      RECT  424.440000  1.615000  424.820000 2.465000 ;
      RECT  425.000000  0.905000  425.380000 1.445000 ;
      RECT  425.040000  0.085000  425.210000 0.565000 ;
      RECT  425.040000  1.835000  425.210000 2.635000 ;
      RECT  425.585000  0.085000  425.875000 0.810000 ;
      RECT  425.585000  1.470000  425.875000 2.635000 ;
      RECT  426.050000  1.075000  427.325000 1.275000 ;
      RECT  426.055000  0.260000  426.385000 0.735000 ;
      RECT  426.055000  0.735000  427.715000 0.905000 ;
      RECT  426.055000  1.445000  427.715000 1.615000 ;
      RECT  426.055000  1.615000  426.385000 2.465000 ;
      RECT  426.605000  0.085000  426.775000 0.565000 ;
      RECT  426.605000  1.785000  426.775000 2.635000 ;
      RECT  426.945000  0.260000  427.325000 0.735000 ;
      RECT  426.945000  1.615000  427.325000 2.465000 ;
      RECT  427.545000  0.085000  427.715000 0.565000 ;
      RECT  427.545000  0.905000  427.715000 1.075000 ;
      RECT  427.545000  1.075000  430.105000 1.275000 ;
      RECT  427.545000  1.275000  427.715000 1.445000 ;
      RECT  427.545000  1.785000  427.715000 2.635000 ;
      RECT  427.885000  0.260000  428.265000 0.735000 ;
      RECT  427.885000  0.735000  430.535000 0.905000 ;
      RECT  427.885000  1.445000  430.535000 1.615000 ;
      RECT  427.885000  1.615000  428.265000 2.465000 ;
      RECT  428.485000  0.085000  428.655000 0.565000 ;
      RECT  428.485000  1.835000  428.655000 2.635000 ;
      RECT  428.825000  0.260000  429.205000 0.735000 ;
      RECT  428.825000  1.615000  429.205000 2.465000 ;
      RECT  429.425000  0.085000  429.595000 0.565000 ;
      RECT  429.425000  1.835000  429.595000 2.635000 ;
      RECT  429.765000  0.260000  430.145000 0.735000 ;
      RECT  429.765000  1.615000  430.145000 2.465000 ;
      RECT  430.360000  0.905000  430.535000 1.075000 ;
      RECT  430.360000  1.075000  437.670000 1.275000 ;
      RECT  430.360000  1.275000  430.535000 1.445000 ;
      RECT  430.365000  0.085000  430.535000 0.565000 ;
      RECT  430.365000  1.835000  430.535000 2.635000 ;
      RECT  430.705000  0.255000  431.005000 0.260000 ;
      RECT  430.705000  0.260000  431.085000 0.735000 ;
      RECT  430.705000  0.735000  438.165000 0.905000 ;
      RECT  430.705000  1.445000  438.165000 1.615000 ;
      RECT  430.705000  1.615000  431.085000 2.465000 ;
      RECT  431.305000  0.085000  431.475000 0.565000 ;
      RECT  431.305000  1.835000  431.475000 2.635000 ;
      RECT  431.645000  0.260000  432.025000 0.735000 ;
      RECT  431.645000  1.615000  432.025000 2.465000 ;
      RECT  431.775000  0.255000  431.945000 0.260000 ;
      RECT  432.245000  0.085000  432.415000 0.565000 ;
      RECT  432.245000  1.835000  432.415000 2.635000 ;
      RECT  432.585000  0.260000  432.965000 0.735000 ;
      RECT  432.585000  1.615000  432.965000 2.465000 ;
      RECT  432.715000  0.255000  432.885000 0.260000 ;
      RECT  433.185000  0.085000  433.355000 0.565000 ;
      RECT  433.185000  1.835000  433.355000 2.635000 ;
      RECT  433.525000  0.260000  433.905000 0.735000 ;
      RECT  433.525000  1.615000  433.905000 2.465000 ;
      RECT  434.125000  0.085000  434.295000 0.565000 ;
      RECT  434.125000  1.835000  434.295000 2.635000 ;
      RECT  434.465000  0.260000  434.845000 0.735000 ;
      RECT  434.465000  1.615000  434.845000 2.465000 ;
      RECT  435.065000  0.085000  435.235000 0.565000 ;
      RECT  435.065000  1.835000  435.235000 2.635000 ;
      RECT  435.405000  0.260000  435.785000 0.735000 ;
      RECT  435.405000  1.615000  435.785000 2.465000 ;
      RECT  436.005000  0.085000  436.175000 0.565000 ;
      RECT  436.005000  1.835000  436.175000 2.635000 ;
      RECT  436.345000  0.260000  436.725000 0.735000 ;
      RECT  436.345000  1.615000  436.725000 2.465000 ;
      RECT  436.945000  0.085000  437.115000 0.565000 ;
      RECT  436.945000  1.835000  437.115000 2.635000 ;
      RECT  437.285000  0.260000  437.665000 0.735000 ;
      RECT  437.285000  1.615000  437.665000 2.465000 ;
      RECT  437.885000  0.085000  438.055000 0.565000 ;
      RECT  437.885000  1.835000  438.055000 2.635000 ;
      RECT  437.890000  0.905000  438.165000 1.445000 ;
      RECT  438.465000  0.085000  438.755000 0.810000 ;
      RECT  438.465000  1.470000  438.755000 2.635000 ;
      RECT  438.925000  1.075000  439.345000 1.275000 ;
      RECT  439.015000  0.085000  439.185000 0.905000 ;
      RECT  439.015000  1.445000  439.185000 2.635000 ;
      RECT  439.355000  0.260000  439.735000 0.905000 ;
      RECT  439.355000  1.545000  439.735000 2.465000 ;
      RECT  439.565000  0.905000  439.735000 1.075000 ;
      RECT  439.565000  1.075000  441.195000 1.275000 ;
      RECT  439.565000  1.275000  439.735000 1.545000 ;
      RECT  439.925000  0.260000  440.255000 0.735000 ;
      RECT  439.925000  0.735000  441.585000 0.905000 ;
      RECT  439.925000  1.445000  441.585000 1.615000 ;
      RECT  439.925000  1.615000  440.255000 2.465000 ;
      RECT  440.475000  0.085000  440.645000 0.565000 ;
      RECT  440.475000  1.785000  440.645000 2.635000 ;
      RECT  440.815000  0.260000  441.195000 0.735000 ;
      RECT  440.815000  1.615000  441.195000 2.465000 ;
      RECT  441.415000  0.085000  441.585000 0.565000 ;
      RECT  441.415000  0.905000  441.585000 1.075000 ;
      RECT  441.415000  1.075000  445.085000 1.275000 ;
      RECT  441.415000  1.275000  441.585000 1.445000 ;
      RECT  441.415000  1.785000  441.585000 2.635000 ;
      RECT  441.755000  0.260000  442.135000 0.735000 ;
      RECT  441.755000  0.735000  445.645000 0.905000 ;
      RECT  441.755000  1.445000  445.645000 1.615000 ;
      RECT  441.755000  1.615000  442.135000 2.465000 ;
      RECT  442.355000  0.085000  442.525000 0.565000 ;
      RECT  442.355000  1.835000  442.525000 2.635000 ;
      RECT  442.695000  0.260000  443.075000 0.735000 ;
      RECT  442.695000  1.615000  443.075000 2.465000 ;
      RECT  443.295000  0.085000  443.465000 0.565000 ;
      RECT  443.295000  1.835000  443.465000 2.635000 ;
      RECT  443.635000  0.260000  444.015000 0.735000 ;
      RECT  443.635000  1.615000  444.015000 2.465000 ;
      RECT  444.235000  0.085000  444.405000 0.565000 ;
      RECT  444.235000  1.835000  444.405000 2.635000 ;
      RECT  444.575000  0.260000  444.955000 0.735000 ;
      RECT  444.575000  1.615000  444.955000 2.465000 ;
      RECT  445.175000  0.085000  445.345000 0.565000 ;
      RECT  445.175000  1.835000  445.345000 2.635000 ;
      RECT  445.255000  0.905000  445.645000 1.445000 ;
      RECT  445.825000  0.085000  446.115000 0.810000 ;
      RECT  445.825000  1.470000  446.115000 2.635000 ;
      RECT  446.285000  0.255000  446.545000 0.760000 ;
      RECT  446.285000  0.760000  446.455000 1.560000 ;
      RECT  446.285000  1.560000  446.555000 2.465000 ;
      RECT  446.625000  1.060000  446.960000 1.390000 ;
      RECT  446.725000  0.085000  447.475000 0.465000 ;
      RECT  446.725000  1.875000  447.475000 2.635000 ;
      RECT  446.740000  0.635000  447.825000 0.805000 ;
      RECT  446.740000  0.805000  446.960000 1.060000 ;
      RECT  446.740000  1.390000  446.960000 1.535000 ;
      RECT  446.740000  1.535000  447.865000 1.705000 ;
      RECT  447.565000  0.985000  447.945000 1.355000 ;
      RECT  447.655000  0.255000  447.825000 0.635000 ;
      RECT  447.695000  1.705000  447.865000 2.465000 ;
      RECT  448.125000  0.085000  448.415000 0.810000 ;
      RECT  448.125000  1.470000  448.415000 2.635000 ;
      RECT  448.585000  0.085000  448.890000 0.595000 ;
      RECT  448.585000  0.765000  448.900000 1.325000 ;
      RECT  448.595000  1.825000  448.890000 2.635000 ;
      RECT  449.120000  0.265000  449.370000 1.075000 ;
      RECT  449.120000  1.075000  457.040000 1.325000 ;
      RECT  449.120000  1.325000  449.365000 2.465000 ;
      RECT  449.590000  0.085000  449.850000 0.610000 ;
      RECT  449.590000  1.825000  449.850000 2.635000 ;
      RECT  450.080000  0.265000  450.330000 1.075000 ;
      RECT  450.080000  1.325000  450.330000 2.460000 ;
      RECT  450.550000  0.085000  450.810000 0.645000 ;
      RECT  450.550000  1.835000  450.810000 2.630000 ;
      RECT  450.550000  2.630000  457.525000 2.635000 ;
      RECT  451.030000  0.280000  451.290000 0.735000 ;
      RECT  451.030000  0.735000  458.525000 0.905000 ;
      RECT  451.030000  1.495000  458.525000 1.720000 ;
      RECT  451.030000  1.720000  457.035000 1.735000 ;
      RECT  451.030000  1.735000  451.290000 2.460000 ;
      RECT  451.510000  0.085000  451.770000 0.565000 ;
      RECT  451.510000  1.905000  451.770000 2.630000 ;
      RECT  451.990000  0.280000  452.250000 0.735000 ;
      RECT  451.990000  1.735000  452.250000 2.460000 ;
      RECT  452.470000  0.085000  452.730000 0.565000 ;
      RECT  452.470000  1.905000  452.730000 2.630000 ;
      RECT  452.950000  0.280000  453.210000 0.735000 ;
      RECT  452.950000  1.735000  453.210000 2.460000 ;
      RECT  453.430000  0.085000  453.675000 0.565000 ;
      RECT  453.430000  1.905000  453.690000 2.630000 ;
      RECT  453.845000  0.280000  454.170000 0.735000 ;
      RECT  453.910000  1.735000  454.170000 2.460000 ;
      RECT  454.390000  0.085000  454.635000 0.565000 ;
      RECT  454.390000  1.905000  454.635000 2.630000 ;
      RECT  454.855000  0.280000  455.115000 0.735000 ;
      RECT  454.855000  1.735000  455.115000 2.460000 ;
      RECT  455.345000  0.085000  455.595000 0.565000 ;
      RECT  455.350000  1.905000  455.595000 2.630000 ;
      RECT  455.815000  0.280000  456.075000 0.735000 ;
      RECT  455.815000  1.735000  456.075000 2.460000 ;
      RECT  456.305000  0.085000  456.555000 0.565000 ;
      RECT  456.310000  1.905000  456.555000 2.630000 ;
      RECT  456.775000  0.280000  457.035000 0.735000 ;
      RECT  456.775000  1.735000  457.035000 2.460000 ;
      RECT  457.260000  0.905000  458.525000 1.495000 ;
      RECT  457.265000  0.085000  457.525000 0.565000 ;
      RECT  457.270000  1.905000  457.525000 2.630000 ;
      RECT  457.745000  0.280000  458.005000 0.735000 ;
      RECT  457.745000  1.720000  458.035000 2.460000 ;
      RECT  458.225000  0.085000  458.525000 0.565000 ;
      RECT  458.255000  1.890000  458.525000 2.635000 ;
      RECT  458.705000  0.085000  458.995000 0.810000 ;
      RECT  458.705000  1.470000  458.995000 2.635000 ;
      RECT  459.165000  0.255000  459.425000 0.585000 ;
      RECT  459.165000  0.585000  459.335000 1.495000 ;
      RECT  459.165000  1.495000  460.395000 1.665000 ;
      RECT  459.165000  1.665000  459.435000 2.435000 ;
      RECT  459.505000  0.745000  459.915000 1.325000 ;
      RECT  459.605000  1.855000  459.985000 2.635000 ;
      RECT  459.685000  0.085000  459.960000 0.565000 ;
      RECT  460.095000  0.995000  460.395000 1.495000 ;
      RECT  460.220000  0.255000  460.425000 0.655000 ;
      RECT  460.220000  0.655000  460.955000 0.825000 ;
      RECT  460.240000  1.855000  460.955000 2.030000 ;
      RECT  460.240000  2.030000  460.425000 2.435000 ;
      RECT  460.565000  0.825000  460.955000 1.855000 ;
      RECT  460.595000  0.085000  460.980000 0.485000 ;
      RECT  460.595000  2.210000  460.980000 2.635000 ;
      RECT  461.465000  0.085000  461.755000 0.810000 ;
      RECT  461.465000  1.470000  461.755000 2.635000 ;
      RECT  461.925000  0.255000  462.225000 0.585000 ;
      RECT  461.925000  0.585000  462.095000 1.495000 ;
      RECT  461.925000  1.495000  463.055000 1.665000 ;
      RECT  461.925000  1.665000  462.235000 2.465000 ;
      RECT  462.265000  0.755000  462.665000 1.325000 ;
      RECT  462.445000  0.085000  462.720000 0.565000 ;
      RECT  462.455000  1.835000  462.765000 2.635000 ;
      RECT  462.835000  1.075000  464.080000 1.245000 ;
      RECT  462.835000  1.245000  463.055000 1.495000 ;
      RECT  462.890000  0.345000  463.245000 0.735000 ;
      RECT  462.890000  0.735000  464.750000 0.905000 ;
      RECT  462.985000  1.835000  464.205000 2.005000 ;
      RECT  462.985000  2.005000  463.245000 2.465000 ;
      RECT  463.465000  0.085000  463.720000 0.565000 ;
      RECT  463.465000  2.175000  463.720000 2.635000 ;
      RECT  463.945000  0.345000  464.205000 0.735000 ;
      RECT  463.945000  1.415000  464.750000 1.650000 ;
      RECT  463.945000  1.650000  464.205000 1.835000 ;
      RECT  463.945000  2.005000  464.205000 2.465000 ;
      RECT  464.250000  0.905000  464.750000 1.415000 ;
      RECT  464.385000  1.845000  464.715000 2.635000 ;
      RECT  464.425000  0.085000  464.705000 0.565000 ;
      RECT  465.145000  0.085000  465.435000 0.810000 ;
      RECT  465.145000  1.470000  465.435000 2.635000 ;
      RECT  465.605000  0.715000  465.920000 1.325000 ;
      RECT  465.615000  1.525000  465.910000 2.635000 ;
      RECT  465.665000  0.085000  465.910000 0.545000 ;
      RECT  466.140000  0.265000  466.390000 1.075000 ;
      RECT  466.140000  1.075000  469.510000 1.325000 ;
      RECT  466.140000  1.325000  466.390000 2.460000 ;
      RECT  466.610000  0.085000  466.870000 0.610000 ;
      RECT  466.610000  1.525000  466.870000 2.635000 ;
      RECT  467.090000  0.280000  467.350000 0.735000 ;
      RECT  467.090000  0.735000  470.750000 0.905000 ;
      RECT  467.090000  1.495000  470.750000 1.735000 ;
      RECT  467.090000  1.735000  467.350000 2.460000 ;
      RECT  467.570000  0.085000  467.830000 0.565000 ;
      RECT  467.570000  1.905000  467.830000 2.635000 ;
      RECT  468.050000  0.280000  468.310000 0.735000 ;
      RECT  468.050000  1.735000  468.310000 2.460000 ;
      RECT  468.530000  0.085000  468.790000 0.565000 ;
      RECT  468.530000  1.905000  468.790000 2.635000 ;
      RECT  469.010000  0.280000  469.270000 0.735000 ;
      RECT  469.010000  1.735000  469.270000 2.460000 ;
      RECT  469.490000  0.085000  469.750000 0.565000 ;
      RECT  469.490000  1.905000  469.750000 2.635000 ;
      RECT  469.680000  0.905000  470.750000 1.495000 ;
      RECT  469.970000  0.280000  470.230000 0.735000 ;
      RECT  469.970000  1.735000  470.230000 2.460000 ;
      RECT  470.450000  0.085000  470.750000 0.565000 ;
      RECT  470.450000  1.905000  470.745000 2.635000 ;
      RECT  471.125000  0.085000  471.415000 0.810000 ;
      RECT  471.125000  1.470000  471.415000 2.635000 ;
      RECT  471.585000  0.375000  471.825000 1.325000 ;
      RECT  471.585000  1.665000  471.845000 2.635000 ;
      RECT  472.015000  0.255000  472.390000 0.760000 ;
      RECT  472.015000  0.760000  472.895000 1.290000 ;
      RECT  472.015000  1.290000  472.395000 2.465000 ;
      RECT  472.615000  0.085000  472.895000 0.590000 ;
      RECT  472.615000  1.665000  472.895000 2.635000 ;
      RECT  473.425000  0.085000  473.715000 0.810000 ;
      RECT  473.425000  1.470000  473.715000 2.635000 ;
      RECT  473.940000  1.495000  474.205000 2.635000 ;
      RECT  474.145000  0.895000  476.155000 1.275000 ;
      RECT  474.425000  1.455000  485.430000 1.665000 ;
      RECT  474.425000  1.665000  474.680000 2.465000 ;
      RECT  474.900000  1.835000  475.160000 2.635000 ;
      RECT  475.385000  1.665000  475.640000 2.450000 ;
      RECT  475.855000  0.085000  476.125000 0.610000 ;
      RECT  475.865000  1.835000  476.120000 2.635000 ;
      RECT  476.375000  0.280000  476.600000 1.415000 ;
      RECT  476.375000  1.415000  483.505000 1.455000 ;
      RECT  476.375000  1.665000  476.600000 2.465000 ;
      RECT  476.820000  0.085000  477.085000 0.610000 ;
      RECT  476.820000  1.835000  477.080000 2.635000 ;
      RECT  477.305000  0.280000  477.560000 1.415000 ;
      RECT  477.305000  1.665000  477.560000 2.450000 ;
      RECT  477.780000  0.085000  478.045000 0.610000 ;
      RECT  477.785000  1.835000  478.040000 2.635000 ;
      RECT  478.265000  0.280000  478.505000 1.415000 ;
      RECT  478.265000  1.665000  478.505000 2.450000 ;
      RECT  478.765000  0.085000  479.030000 0.610000 ;
      RECT  478.765000  1.835000  479.020000 2.635000 ;
      RECT  479.255000  0.280000  479.605000 1.415000 ;
      RECT  479.255000  1.665000  479.630000 2.450000 ;
      RECT  479.890000  0.085000  480.155000 0.610000 ;
      RECT  479.890000  1.835000  480.145000 2.120000 ;
      RECT  479.890000  2.120000  480.150000 2.635000 ;
      RECT  480.375000  0.280000  480.625000 1.415000 ;
      RECT  480.375000  1.665000  480.625000 2.450000 ;
      RECT  480.850000  0.085000  481.075000 0.610000 ;
      RECT  480.855000  1.835000  481.110000 2.635000 ;
      RECT  481.335000  0.280000  481.585000 1.415000 ;
      RECT  481.335000  1.665000  481.585000 2.450000 ;
      RECT  481.810000  0.085000  482.075000 0.610000 ;
      RECT  481.815000  1.835000  482.070000 2.635000 ;
      RECT  482.295000  0.280000  482.545000 1.415000 ;
      RECT  482.295000  1.665000  482.545000 2.450000 ;
      RECT  482.770000  0.085000  483.035000 0.610000 ;
      RECT  482.775000  1.835000  483.030000 2.635000 ;
      RECT  483.255000  0.280000  483.505000 1.415000 ;
      RECT  483.255000  1.665000  483.505000 2.450000 ;
      RECT  483.730000  0.085000  483.995000 0.610000 ;
      RECT  483.730000  0.895000  485.710000 1.275000 ;
      RECT  483.735000  1.835000  483.990000 2.635000 ;
      RECT  484.215000  1.665000  484.455000 2.450000 ;
      RECT  484.695000  1.835000  484.950000 2.635000 ;
      RECT  485.175000  1.665000  485.430000 2.450000 ;
      RECT  485.650000  1.835000  485.910000 2.635000 ;
      RECT  486.305000  0.085000  486.595000 0.810000 ;
      RECT  486.305000  1.470000  486.595000 2.635000 ;
      RECT  486.765000  1.065000  488.015000 1.290000 ;
      RECT  486.835000  1.460000  488.835000 1.630000 ;
      RECT  486.835000  1.630000  487.090000 2.435000 ;
      RECT  487.240000  0.085000  487.585000 0.610000 ;
      RECT  487.310000  1.800000  487.570000 2.635000 ;
      RECT  487.790000  1.630000  488.050000 2.435000 ;
      RECT  487.805000  0.280000  488.030000 0.725000 ;
      RECT  487.805000  0.725000  488.835000 0.895000 ;
      RECT  488.200000  0.085000  488.580000 0.555000 ;
      RECT  488.200000  0.895000  488.835000 1.460000 ;
      RECT  488.285000  1.800000  488.540000 2.635000 ;
      RECT  489.065000  0.085000  489.355000 0.810000 ;
      RECT  489.065000  1.470000  489.355000 2.635000 ;
      RECT  489.525000  1.800000  489.870000 2.635000 ;
      RECT  489.545000  0.725000  493.010000 0.895000 ;
      RECT  489.545000  0.895000  489.715000 1.460000 ;
      RECT  489.545000  1.460000  493.010000 1.630000 ;
      RECT  489.885000  1.065000  492.350000 1.290000 ;
      RECT  490.005000  0.085000  490.350000 0.555000 ;
      RECT  490.095000  1.630000  490.350000 2.435000 ;
      RECT  490.570000  0.280000  490.830000 0.725000 ;
      RECT  490.570000  1.800000  490.830000 2.635000 ;
      RECT  491.050000  0.085000  491.310000 0.555000 ;
      RECT  491.055000  1.630000  491.310000 2.435000 ;
      RECT  491.530000  0.280000  491.785000 0.725000 ;
      RECT  491.530000  1.800000  491.790000 2.635000 ;
      RECT  492.005000  0.085000  492.305000 0.555000 ;
      RECT  492.010000  1.630000  492.270000 2.435000 ;
      RECT  492.490000  1.800000  492.875000 2.635000 ;
      RECT  492.710000  0.895000  493.010000 1.460000 ;
      RECT  493.205000  0.085000  493.495000 0.810000 ;
      RECT  493.205000  1.470000  493.495000 2.635000 ;
      RECT  493.695000  0.695000  499.910000 0.865000 ;
      RECT  493.695000  0.865000  493.865000 1.460000 ;
      RECT  493.695000  1.460000  499.910000 1.630000 ;
      RECT  493.715000  1.800000  493.975000 2.635000 ;
      RECT  494.035000  1.035000  499.145000 1.290000 ;
      RECT  494.195000  1.630000  494.435000 2.435000 ;
      RECT  494.655000  1.800000  494.915000 2.635000 ;
      RECT  494.715000  0.085000  495.045000 0.525000 ;
      RECT  495.135000  1.630000  495.375000 2.435000 ;
      RECT  495.265000  0.280000  495.455000 0.695000 ;
      RECT  495.595000  1.800000  495.855000 2.635000 ;
      RECT  495.675000  0.085000  496.005000 0.525000 ;
      RECT  496.075000  1.630000  496.325000 2.435000 ;
      RECT  496.225000  0.280000  496.415000 0.695000 ;
      RECT  496.545000  1.800000  496.790000 2.635000 ;
      RECT  496.635000  0.085000  497.015000 0.525000 ;
      RECT  497.010000  1.630000  497.255000 2.435000 ;
      RECT  497.185000  0.280000  497.375000 0.695000 ;
      RECT  497.475000  1.800000  497.780000 2.635000 ;
      RECT  497.595000  0.085000  498.025000 0.525000 ;
      RECT  498.000000  1.630000  498.305000 2.435000 ;
      RECT  498.245000  0.280000  498.435000 0.695000 ;
      RECT  498.525000  1.800000  498.825000 2.635000 ;
      RECT  498.655000  0.085000  499.085000 0.525000 ;
      RECT  499.045000  1.630000  499.285000 2.435000 ;
      RECT  499.505000  1.800000  499.760000 2.635000 ;
      RECT  499.640000  0.865000  499.910000 1.460000 ;
      RECT  500.105000  0.085000  500.395000 0.810000 ;
      RECT  500.105000  1.470000  500.395000 2.635000 ;
      RECT  500.625000  0.995000  501.080000 1.665000 ;
      RECT  500.705000  1.835000  501.035000 2.625000 ;
      RECT  500.705000  2.625000  502.145000 2.635000 ;
      RECT  500.775000  0.085000  501.095000 0.745000 ;
      RECT  501.265000  0.315000  502.025000 0.750000 ;
      RECT  501.265000  0.750000  501.715000 2.455000 ;
      RECT  501.885000  1.455000  502.145000 2.625000 ;
      RECT  502.405000  0.085000  502.695000 0.810000 ;
      RECT  502.405000  1.470000  502.695000 2.635000 ;
      RECT  502.865000  0.745000  503.205000 1.325000 ;
      RECT  502.875000  0.085000  503.205000 0.575000 ;
      RECT  502.875000  1.495000  503.200000 2.635000 ;
      RECT  503.385000  0.255000  503.945000 0.680000 ;
      RECT  503.385000  0.680000  503.735000 1.015000 ;
      RECT  503.385000  1.015000  504.765000 1.295000 ;
      RECT  503.385000  1.295000  503.725000 2.465000 ;
      RECT  503.965000  1.465000  504.240000 2.635000 ;
      RECT  504.435000  1.295000  504.765000 2.465000 ;
      RECT  504.455000  0.085000  504.780000 0.775000 ;
      RECT  505.005000  1.465000  505.285000 2.635000 ;
      RECT  505.625000  0.085000  505.915000 0.810000 ;
      RECT  505.625000  1.470000  505.915000 2.635000 ;
      RECT  506.085000  0.255000  506.605000 1.740000 ;
      RECT  506.275000  1.910000  506.605000 2.635000 ;
      RECT  506.775000  0.085000  507.115000 0.745000 ;
      RECT  506.775000  0.915000  507.295000 2.465000 ;
      RECT  507.465000  0.085000  507.755000 0.810000 ;
      RECT  507.465000  1.470000  507.755000 2.635000 ;
      RECT  507.930000  0.345000  508.185000 0.635000 ;
      RECT  507.930000  0.635000  508.730000 0.805000 ;
      RECT  507.930000  0.975000  508.280000 1.625000 ;
      RECT  507.930000  1.795000  508.730000 1.965000 ;
      RECT  507.930000  1.965000  508.185000 2.465000 ;
      RECT  508.355000  0.085000  508.735000 0.465000 ;
      RECT  508.355000  2.135000  508.735000 2.635000 ;
      RECT  508.500000  0.805000  508.730000 1.795000 ;
      RECT  508.955000  0.345000  509.125000 2.465000 ;
      RECT  509.295000  0.615000  509.745000 1.665000 ;
      RECT  509.295000  1.665000  509.610000 2.005000 ;
      RECT  509.415000  0.085000  509.745000 0.445000 ;
      RECT  509.610000  2.175000  509.780000 2.635000 ;
      RECT  509.915000  0.305000  510.335000 0.475000 ;
      RECT  509.915000  0.475000  510.085000 1.835000 ;
      RECT  509.915000  1.835000  510.180000 2.005000 ;
      RECT  510.010000  2.005000  510.180000 2.135000 ;
      RECT  510.010000  2.135000  510.260000 2.465000 ;
      RECT  510.265000  0.765000  510.525000 1.385000 ;
      RECT  510.350000  1.575000  510.865000 1.965000 ;
      RECT  510.525000  2.135000  511.205000 2.465000 ;
      RECT  510.535000  0.305000  511.440000 0.475000 ;
      RECT  510.695000  0.765000  511.050000 0.985000 ;
      RECT  510.695000  0.985000  510.865000 1.575000 ;
      RECT  511.035000  1.185000  512.825000 1.355000 ;
      RECT  511.035000  1.355000  511.205000 2.135000 ;
      RECT  511.270000  0.475000  511.440000 1.185000 ;
      RECT  511.375000  1.865000  512.550000 2.035000 ;
      RECT  511.375000  2.035000  511.545000 2.375000 ;
      RECT  511.565000  1.525000  513.165000 1.695000 ;
      RECT  511.645000  0.765000  512.485000 1.015000 ;
      RECT  511.830000  2.205000  512.160000 2.635000 ;
      RECT  512.365000  0.085000  512.695000 0.545000 ;
      RECT  512.380000  2.035000  512.550000 2.375000 ;
      RECT  512.655000  1.005000  512.825000 1.185000 ;
      RECT  512.845000  2.175000  513.265000 2.635000 ;
      RECT  512.905000  0.275000  513.305000 0.445000 ;
      RECT  512.905000  0.445000  513.165000 0.835000 ;
      RECT  512.995000  0.835000  513.165000 1.525000 ;
      RECT  512.995000  1.695000  513.165000 1.835000 ;
      RECT  512.995000  1.835000  513.655000 2.005000 ;
      RECT  513.445000  0.705000  513.615000 1.495000 ;
      RECT  513.445000  1.495000  514.155000 1.655000 ;
      RECT  513.445000  1.655000  514.500000 1.665000 ;
      RECT  513.485000  2.005000  513.655000 2.465000 ;
      RECT  513.575000  0.255000  514.495000 0.535000 ;
      RECT  513.785000  0.705000  514.155000 1.325000 ;
      RECT  513.890000  2.125000  514.845000 2.465000 ;
      RECT  513.985000  1.665000  514.500000 1.955000 ;
      RECT  514.325000  0.535000  514.495000 1.315000 ;
      RECT  514.325000  1.315000  514.895000 1.485000 ;
      RECT  514.665000  0.085000  514.835000 0.525000 ;
      RECT  514.675000  1.485000  514.895000 1.575000 ;
      RECT  514.675000  1.575000  516.110000 1.745000 ;
      RECT  514.675000  1.745000  514.845000 2.125000 ;
      RECT  514.795000  0.695000  515.175000 0.865000 ;
      RECT  514.795000  0.865000  515.065000 1.145000 ;
      RECT  515.005000  0.295000  516.475000 0.465000 ;
      RECT  515.005000  0.465000  515.175000 0.695000 ;
      RECT  515.180000  2.175000  515.430000 2.635000 ;
      RECT  515.345000  0.635000  515.745000 1.405000 ;
      RECT  515.650000  1.915000  516.450000 2.085000 ;
      RECT  515.650000  2.085000  515.820000 2.375000 ;
      RECT  516.000000  2.255000  516.380000 2.635000 ;
      RECT  516.130000  0.465000  516.475000 1.075000 ;
      RECT  516.130000  1.075000  516.910000 1.285000 ;
      RECT  516.130000  1.285000  516.450000 1.295000 ;
      RECT  516.280000  1.295000  516.450000 1.915000 ;
      RECT  516.650000  0.085000  516.820000 0.895000 ;
      RECT  516.650000  1.575000  516.820000 2.635000 ;
      RECT  517.080000  0.255000  517.415000 2.465000 ;
      RECT  517.585000  0.085000  517.875000 0.810000 ;
      RECT  517.585000  1.470000  517.875000 2.635000 ;
      RECT  518.050000  0.345000  518.305000 0.635000 ;
      RECT  518.050000  0.635000  518.850000 0.805000 ;
      RECT  518.050000  0.975000  518.400000 1.625000 ;
      RECT  518.050000  1.795000  518.850000 1.965000 ;
      RECT  518.050000  1.965000  518.305000 2.465000 ;
      RECT  518.475000  0.085000  518.855000 0.465000 ;
      RECT  518.475000  2.135000  518.855000 2.635000 ;
      RECT  518.620000  0.805000  518.850000 1.795000 ;
      RECT  519.075000  0.345000  519.245000 2.465000 ;
      RECT  519.415000  0.615000  519.865000 1.665000 ;
      RECT  519.415000  1.665000  519.730000 2.005000 ;
      RECT  519.535000  0.085000  519.865000 0.445000 ;
      RECT  519.730000  2.175000  519.900000 2.635000 ;
      RECT  520.035000  0.305000  520.455000 0.475000 ;
      RECT  520.035000  0.475000  520.205000 1.835000 ;
      RECT  520.035000  1.835000  520.300000 2.005000 ;
      RECT  520.130000  2.005000  520.300000 2.135000 ;
      RECT  520.130000  2.135000  520.380000 2.465000 ;
      RECT  520.385000  0.765000  520.645000 1.385000 ;
      RECT  520.470000  1.575000  520.985000 1.965000 ;
      RECT  520.645000  2.135000  521.325000 2.465000 ;
      RECT  520.655000  0.305000  521.560000 0.475000 ;
      RECT  520.815000  0.765000  521.170000 0.985000 ;
      RECT  520.815000  0.985000  520.985000 1.575000 ;
      RECT  521.155000  1.185000  522.945000 1.355000 ;
      RECT  521.155000  1.355000  521.325000 2.135000 ;
      RECT  521.390000  0.475000  521.560000 1.185000 ;
      RECT  521.495000  1.865000  522.670000 2.035000 ;
      RECT  521.495000  2.035000  521.665000 2.375000 ;
      RECT  521.685000  1.525000  523.285000 1.695000 ;
      RECT  521.765000  0.765000  522.605000 1.015000 ;
      RECT  521.950000  2.205000  522.280000 2.635000 ;
      RECT  522.485000  0.085000  522.815000 0.545000 ;
      RECT  522.500000  2.035000  522.670000 2.375000 ;
      RECT  522.775000  1.005000  522.945000 1.185000 ;
      RECT  522.965000  2.175000  523.385000 2.635000 ;
      RECT  523.025000  0.275000  523.425000 0.445000 ;
      RECT  523.025000  0.445000  523.285000 0.835000 ;
      RECT  523.115000  0.835000  523.285000 1.525000 ;
      RECT  523.115000  1.695000  523.285000 1.835000 ;
      RECT  523.115000  1.835000  523.775000 2.005000 ;
      RECT  523.565000  0.705000  523.735000 1.495000 ;
      RECT  523.565000  1.495000  524.275000 1.655000 ;
      RECT  523.565000  1.655000  524.620000 1.665000 ;
      RECT  523.605000  2.005000  523.775000 2.465000 ;
      RECT  523.695000  0.255000  524.615000 0.535000 ;
      RECT  523.905000  0.705000  524.275000 1.325000 ;
      RECT  524.010000  2.125000  524.965000 2.465000 ;
      RECT  524.105000  1.665000  524.620000 1.955000 ;
      RECT  524.445000  0.535000  524.615000 1.315000 ;
      RECT  524.445000  1.315000  525.015000 1.485000 ;
      RECT  524.785000  0.085000  524.955000 0.525000 ;
      RECT  524.795000  1.485000  525.015000 1.575000 ;
      RECT  524.795000  1.575000  526.230000 1.745000 ;
      RECT  524.795000  1.745000  524.965000 2.125000 ;
      RECT  524.915000  0.695000  525.295000 0.865000 ;
      RECT  524.915000  0.865000  525.185000 1.145000 ;
      RECT  525.125000  0.295000  526.595000 0.465000 ;
      RECT  525.125000  0.465000  525.295000 0.695000 ;
      RECT  525.300000  2.175000  525.550000 2.635000 ;
      RECT  525.465000  0.635000  525.865000 1.405000 ;
      RECT  525.770000  1.915000  526.570000 2.085000 ;
      RECT  525.770000  2.085000  525.940000 2.375000 ;
      RECT  526.120000  2.255000  526.500000 2.635000 ;
      RECT  526.250000  0.465000  526.595000 1.075000 ;
      RECT  526.250000  1.075000  527.295000 1.285000 ;
      RECT  526.250000  1.285000  526.570000 1.295000 ;
      RECT  526.400000  1.295000  526.570000 1.915000 ;
      RECT  526.770000  0.085000  526.940000 0.895000 ;
      RECT  526.770000  1.575000  526.940000 2.635000 ;
      RECT  527.110000  0.255000  527.490000 0.735000 ;
      RECT  527.110000  0.735000  527.970000 0.905000 ;
      RECT  527.200000  1.455000  527.970000 1.625000 ;
      RECT  527.200000  1.625000  527.490000 2.465000 ;
      RECT  527.585000  0.905000  527.970000 1.455000 ;
      RECT  527.710000  0.085000  527.880000 0.555000 ;
      RECT  527.710000  1.795000  527.880000 2.635000 ;
      RECT  528.165000  0.085000  528.455000 0.810000 ;
      RECT  528.165000  1.470000  528.455000 2.635000 ;
      RECT  528.630000  0.345000  528.885000 0.635000 ;
      RECT  528.630000  0.635000  529.430000 0.805000 ;
      RECT  528.630000  0.975000  528.980000 1.625000 ;
      RECT  528.630000  1.795000  529.430000 1.965000 ;
      RECT  528.630000  1.965000  528.885000 2.465000 ;
      RECT  529.055000  0.085000  529.435000 0.465000 ;
      RECT  529.055000  2.135000  529.435000 2.635000 ;
      RECT  529.200000  0.805000  529.430000 1.795000 ;
      RECT  529.655000  0.345000  529.825000 2.465000 ;
      RECT  529.995000  0.615000  530.515000 1.665000 ;
      RECT  529.995000  1.665000  530.320000 2.450000 ;
      RECT  530.185000  0.085000  530.515000 0.445000 ;
      RECT  530.490000  2.175000  530.740000 2.635000 ;
      RECT  530.685000  0.305000  531.230000 0.475000 ;
      RECT  530.685000  0.475000  530.855000 1.835000 ;
      RECT  530.685000  1.835000  531.130000 2.005000 ;
      RECT  530.960000  2.005000  531.130000 2.135000 ;
      RECT  530.960000  2.135000  531.210000 2.465000 ;
      RECT  531.075000  0.765000  531.475000 1.385000 ;
      RECT  531.300000  1.575000  531.815000 1.965000 ;
      RECT  531.475000  2.135000  532.205000 2.465000 ;
      RECT  531.485000  0.305000  532.390000 0.475000 ;
      RECT  531.645000  0.765000  532.050000 0.985000 ;
      RECT  531.645000  0.985000  531.815000 1.575000 ;
      RECT  532.035000  1.185000  533.825000 1.355000 ;
      RECT  532.035000  1.355000  532.205000 2.135000 ;
      RECT  532.220000  0.475000  532.390000 1.185000 ;
      RECT  532.375000  1.865000  533.550000 2.035000 ;
      RECT  532.375000  2.035000  532.545000 2.375000 ;
      RECT  532.565000  1.525000  534.215000 1.695000 ;
      RECT  532.715000  0.765000  533.485000 1.015000 ;
      RECT  532.830000  2.205000  533.160000 2.635000 ;
      RECT  533.365000  0.085000  533.695000 0.545000 ;
      RECT  533.380000  2.035000  533.550000 2.375000 ;
      RECT  533.655000  1.005000  533.825000 1.185000 ;
      RECT  533.845000  2.175000  534.265000 2.635000 ;
      RECT  533.905000  0.275000  534.305000 0.445000 ;
      RECT  533.905000  0.445000  534.215000 0.835000 ;
      RECT  534.045000  0.835000  534.215000 1.525000 ;
      RECT  534.045000  1.695000  534.215000 1.835000 ;
      RECT  534.045000  1.835000  534.655000 2.005000 ;
      RECT  534.455000  0.705000  534.665000 1.495000 ;
      RECT  534.455000  1.495000  535.230000 1.655000 ;
      RECT  534.455000  1.655000  535.570000 1.665000 ;
      RECT  534.485000  2.005000  534.655000 2.465000 ;
      RECT  534.575000  0.255000  535.675000 0.535000 ;
      RECT  534.835000  0.705000  535.285000 1.325000 ;
      RECT  534.890000  2.125000  536.010000 2.465000 ;
      RECT  535.010000  1.665000  535.570000 1.955000 ;
      RECT  535.505000  0.535000  535.675000 1.315000 ;
      RECT  535.505000  1.315000  536.010000 1.485000 ;
      RECT  535.790000  1.485000  536.010000 1.575000 ;
      RECT  535.790000  1.575000  537.160000 1.745000 ;
      RECT  535.790000  1.745000  536.010000 2.125000 ;
      RECT  535.895000  0.085000  536.135000 0.525000 ;
      RECT  535.895000  0.695000  536.475000 0.865000 ;
      RECT  535.895000  0.865000  536.165000 1.145000 ;
      RECT  536.180000  2.175000  536.430000 2.635000 ;
      RECT  536.305000  0.295000  537.475000 0.465000 ;
      RECT  536.305000  0.465000  536.475000 0.695000 ;
      RECT  536.345000  1.035000  536.935000 1.405000 ;
      RECT  536.650000  1.915000  537.500000 2.085000 ;
      RECT  536.650000  2.085000  536.820000 2.375000 ;
      RECT  536.695000  0.635000  536.935000 1.035000 ;
      RECT  537.000000  2.255000  537.380000 2.635000 ;
      RECT  537.155000  0.465000  537.475000 0.820000 ;
      RECT  537.155000  0.820000  537.480000 1.075000 ;
      RECT  537.155000  1.075000  539.335000 1.285000 ;
      RECT  537.155000  1.285000  537.500000 1.295000 ;
      RECT  537.330000  1.295000  537.500000 1.915000 ;
      RECT  537.675000  0.085000  537.845000 0.895000 ;
      RECT  537.675000  1.575000  537.845000 2.635000 ;
      RECT  538.015000  0.255000  538.395000 0.735000 ;
      RECT  538.015000  0.735000  539.945000 0.905000 ;
      RECT  538.105000  1.455000  539.945000 1.625000 ;
      RECT  538.105000  1.625000  538.395000 2.465000 ;
      RECT  538.615000  0.085000  538.785000 0.555000 ;
      RECT  538.615000  1.795000  538.785000 2.635000 ;
      RECT  538.955000  0.255000  539.335000 0.735000 ;
      RECT  539.045000  1.625000  539.295000 2.465000 ;
      RECT  539.535000  0.905000  539.945000 1.455000 ;
      RECT  539.555000  0.085000  539.725000 0.555000 ;
      RECT  539.555000  1.795000  539.725000 2.635000 ;
      RECT  540.125000  0.085000  540.415000 0.810000 ;
      RECT  540.125000  1.470000  540.415000 2.635000 ;
      RECT  540.590000  0.975000  540.940000 1.625000 ;
      RECT  540.675000  0.345000  540.845000 0.635000 ;
      RECT  540.675000  0.635000  541.390000 0.805000 ;
      RECT  540.675000  1.795000  541.390000 1.965000 ;
      RECT  540.675000  1.965000  540.845000 2.465000 ;
      RECT  541.015000  0.085000  541.395000 0.465000 ;
      RECT  541.015000  2.135000  541.395000 2.635000 ;
      RECT  541.160000  0.805000  541.390000 1.795000 ;
      RECT  541.615000  0.345000  541.840000 2.465000 ;
      RECT  542.030000  0.635000  542.775000 0.825000 ;
      RECT  542.030000  0.825000  542.200000 1.795000 ;
      RECT  542.030000  1.795000  542.775000 1.965000 ;
      RECT  542.055000  0.085000  542.385000 0.465000 ;
      RECT  542.055000  2.135000  542.385000 2.635000 ;
      RECT  542.370000  1.005000  542.830000 1.625000 ;
      RECT  542.605000  0.305000  542.775000 0.635000 ;
      RECT  542.605000  1.965000  542.775000 2.465000 ;
      RECT  543.000000  0.705000  543.270000 1.575000 ;
      RECT  543.000000  1.575000  543.600000 1.955000 ;
      RECT  543.010000  2.250000  543.940000 2.420000 ;
      RECT  543.125000  0.265000  544.240000 0.465000 ;
      RECT  543.450000  0.645000  543.850000 1.015000 ;
      RECT  543.770000  1.230000  544.240000 1.235000 ;
      RECT  543.770000  1.235000  545.270000 1.405000 ;
      RECT  543.770000  1.405000  543.940000 2.250000 ;
      RECT  544.020000  0.465000  544.240000 1.230000 ;
      RECT  544.110000  1.575000  544.410000 1.835000 ;
      RECT  544.110000  1.835000  545.610000 2.085000 ;
      RECT  544.230000  2.255000  544.610000 2.635000 ;
      RECT  544.410000  0.085000  544.870000 0.525000 ;
      RECT  544.410000  0.735000  545.010000 1.065000 ;
      RECT  544.840000  2.085000  545.010000 2.375000 ;
      RECT  544.970000  1.405000  545.270000 1.565000 ;
      RECT  545.180000  2.255000  545.560000 2.635000 ;
      RECT  545.290000  0.295000  545.460000 0.725000 ;
      RECT  545.290000  0.725000  545.610000 1.065000 ;
      RECT  545.440000  1.065000  545.610000 1.835000 ;
      RECT  545.640000  0.085000  546.030000 0.545000 ;
      RECT  545.830000  0.725000  547.250000 0.895000 ;
      RECT  545.830000  0.895000  546.000000 1.655000 ;
      RECT  545.830000  1.655000  546.400000 1.965000 ;
      RECT  546.060000  2.165000  546.790000 2.415000 ;
      RECT  546.220000  1.065000  546.400000 1.475000 ;
      RECT  546.570000  1.235000  548.670000 1.405000 ;
      RECT  546.570000  1.405000  546.790000 1.915000 ;
      RECT  546.570000  1.915000  547.880000 2.085000 ;
      RECT  546.570000  2.085000  546.790000 2.165000 ;
      RECT  546.690000  0.305000  547.590000 0.475000 ;
      RECT  546.870000  0.895000  547.250000 1.015000 ;
      RECT  546.960000  1.575000  549.050000 1.745000 ;
      RECT  546.970000  2.255000  547.440000 2.635000 ;
      RECT  547.420000  0.475000  547.590000 1.235000 ;
      RECT  547.640000  2.085000  547.880000 2.375000 ;
      RECT  547.760000  0.735000  548.280000 1.005000 ;
      RECT  547.760000  1.005000  548.140000 1.065000 ;
      RECT  547.820000  0.085000  548.530000 0.565000 ;
      RECT  548.210000  1.945000  548.540000 2.635000 ;
      RECT  548.290000  1.175000  548.670000 1.235000 ;
      RECT  548.710000  0.350000  549.050000 0.680000 ;
      RECT  548.710000  1.745000  549.050000 1.765000 ;
      RECT  548.710000  1.765000  548.880000 2.375000 ;
      RECT  548.840000  0.680000  549.050000 1.575000 ;
      RECT  549.150000  1.915000  549.480000 2.425000 ;
      RECT  549.230000  0.345000  549.480000 0.995000 ;
      RECT  549.230000  0.995000  550.080000 1.325000 ;
      RECT  549.230000  1.325000  549.480000 1.915000 ;
      RECT  549.650000  0.085000  550.085000 0.545000 ;
      RECT  549.650000  1.835000  550.070000 2.635000 ;
      RECT  550.240000  1.655000  550.525000 2.325000 ;
      RECT  550.255000  0.265000  550.525000 0.795000 ;
      RECT  550.300000  0.795000  550.525000 1.655000 ;
      RECT  550.705000  0.085000  550.995000 0.810000 ;
      RECT  550.705000  1.470000  550.995000 2.635000 ;
      RECT  551.170000  0.975000  551.520000 1.625000 ;
      RECT  551.255000  0.345000  551.425000 0.635000 ;
      RECT  551.255000  0.635000  551.970000 0.805000 ;
      RECT  551.255000  1.795000  551.970000 1.965000 ;
      RECT  551.255000  1.965000  551.425000 2.465000 ;
      RECT  551.595000  0.085000  551.975000 0.465000 ;
      RECT  551.595000  2.135000  551.975000 2.635000 ;
      RECT  551.740000  0.805000  551.970000 1.795000 ;
      RECT  552.195000  0.345000  552.420000 2.465000 ;
      RECT  552.610000  0.635000  553.355000 0.825000 ;
      RECT  552.610000  0.825000  552.780000 1.795000 ;
      RECT  552.610000  1.795000  553.355000 1.965000 ;
      RECT  552.635000  0.085000  552.965000 0.465000 ;
      RECT  552.635000  2.135000  552.965000 2.635000 ;
      RECT  552.950000  1.005000  553.410000 1.625000 ;
      RECT  553.185000  0.305000  553.355000 0.635000 ;
      RECT  553.185000  1.965000  553.355000 2.465000 ;
      RECT  553.580000  0.705000  553.850000 1.575000 ;
      RECT  553.580000  1.575000  554.180000 1.955000 ;
      RECT  553.590000  2.250000  554.520000 2.420000 ;
      RECT  553.705000  0.265000  554.820000 0.465000 ;
      RECT  554.030000  0.645000  554.430000 1.015000 ;
      RECT  554.350000  1.230000  554.820000 1.235000 ;
      RECT  554.350000  1.235000  555.850000 1.405000 ;
      RECT  554.350000  1.405000  554.520000 2.250000 ;
      RECT  554.600000  0.465000  554.820000 1.230000 ;
      RECT  554.690000  1.575000  554.990000 1.835000 ;
      RECT  554.690000  1.835000  556.190000 2.085000 ;
      RECT  554.810000  2.255000  555.190000 2.635000 ;
      RECT  554.990000  0.085000  555.450000 0.525000 ;
      RECT  554.990000  0.735000  555.590000 1.065000 ;
      RECT  555.420000  2.085000  555.590000 2.375000 ;
      RECT  555.550000  1.405000  555.850000 1.565000 ;
      RECT  555.760000  2.255000  556.140000 2.635000 ;
      RECT  555.870000  0.295000  556.040000 0.725000 ;
      RECT  555.870000  0.725000  556.190000 1.065000 ;
      RECT  556.020000  1.065000  556.190000 1.835000 ;
      RECT  556.220000  0.085000  556.610000 0.545000 ;
      RECT  556.410000  0.725000  557.830000 0.895000 ;
      RECT  556.410000  0.895000  556.580000 1.655000 ;
      RECT  556.410000  1.655000  556.980000 1.965000 ;
      RECT  556.640000  2.165000  557.370000 2.415000 ;
      RECT  556.800000  1.065000  556.980000 1.475000 ;
      RECT  557.150000  1.235000  559.250000 1.405000 ;
      RECT  557.150000  1.405000  557.370000 1.915000 ;
      RECT  557.150000  1.915000  558.460000 2.085000 ;
      RECT  557.150000  2.085000  557.370000 2.165000 ;
      RECT  557.270000  0.305000  558.170000 0.475000 ;
      RECT  557.450000  0.895000  557.830000 1.015000 ;
      RECT  557.540000  1.575000  559.630000 1.745000 ;
      RECT  557.550000  2.255000  558.020000 2.635000 ;
      RECT  558.000000  0.475000  558.170000 1.235000 ;
      RECT  558.220000  2.085000  558.460000 2.375000 ;
      RECT  558.340000  0.735000  558.860000 1.005000 ;
      RECT  558.340000  1.005000  558.720000 1.065000 ;
      RECT  558.400000  0.085000  559.110000 0.565000 ;
      RECT  558.790000  1.945000  559.120000 2.635000 ;
      RECT  558.870000  1.175000  559.250000 1.235000 ;
      RECT  559.290000  0.350000  559.630000 0.680000 ;
      RECT  559.290000  1.745000  559.630000 1.765000 ;
      RECT  559.290000  1.765000  559.460000 2.375000 ;
      RECT  559.420000  0.680000  559.630000 1.575000 ;
      RECT  559.730000  1.915000  560.060000 2.425000 ;
      RECT  559.810000  0.345000  559.980000 0.995000 ;
      RECT  559.810000  0.995000  560.660000 1.325000 ;
      RECT  559.810000  1.325000  560.060000 1.915000 ;
      RECT  560.150000  0.085000  560.530000 0.825000 ;
      RECT  560.280000  1.495000  560.450000 2.635000 ;
      RECT  560.620000  1.495000  561.565000 1.615000 ;
      RECT  560.620000  1.615000  561.095000 2.460000 ;
      RECT  560.765000  0.265000  561.095000 0.745000 ;
      RECT  560.765000  0.745000  561.565000 0.825000 ;
      RECT  560.830000  0.825000  561.565000 1.495000 ;
      RECT  561.265000  0.085000  561.530000 0.575000 ;
      RECT  561.265000  1.785000  561.530000 2.635000 ;
      RECT  561.745000  0.085000  562.035000 0.810000 ;
      RECT  561.745000  1.470000  562.035000 2.635000 ;
      RECT  562.210000  0.975000  562.560000 1.625000 ;
      RECT  562.295000  0.345000  562.465000 0.635000 ;
      RECT  562.295000  0.635000  563.010000 0.805000 ;
      RECT  562.295000  1.795000  563.010000 1.965000 ;
      RECT  562.295000  1.965000  562.465000 2.465000 ;
      RECT  562.635000  0.085000  563.015000 0.465000 ;
      RECT  562.635000  2.135000  563.015000 2.635000 ;
      RECT  562.780000  0.805000  563.010000 1.795000 ;
      RECT  563.235000  0.345000  563.460000 2.465000 ;
      RECT  563.650000  0.635000  564.395000 0.825000 ;
      RECT  563.650000  0.825000  563.820000 1.795000 ;
      RECT  563.650000  1.795000  564.395000 1.965000 ;
      RECT  563.675000  0.085000  564.005000 0.465000 ;
      RECT  563.675000  2.135000  564.005000 2.635000 ;
      RECT  563.990000  1.005000  564.450000 1.625000 ;
      RECT  564.225000  0.305000  564.395000 0.635000 ;
      RECT  564.225000  1.965000  564.395000 2.465000 ;
      RECT  564.620000  0.705000  564.890000 1.575000 ;
      RECT  564.620000  1.575000  565.220000 1.955000 ;
      RECT  564.630000  2.250000  565.560000 2.420000 ;
      RECT  564.745000  0.265000  565.860000 0.465000 ;
      RECT  565.070000  0.645000  565.470000 1.015000 ;
      RECT  565.390000  1.230000  565.860000 1.235000 ;
      RECT  565.390000  1.235000  566.890000 1.405000 ;
      RECT  565.390000  1.405000  565.560000 2.250000 ;
      RECT  565.640000  0.465000  565.860000 1.230000 ;
      RECT  565.730000  1.575000  566.030000 1.835000 ;
      RECT  565.730000  1.835000  567.230000 2.085000 ;
      RECT  565.850000  2.255000  566.230000 2.635000 ;
      RECT  566.030000  0.085000  566.490000 0.525000 ;
      RECT  566.030000  0.735000  566.630000 1.065000 ;
      RECT  566.460000  2.085000  566.630000 2.375000 ;
      RECT  566.590000  1.405000  566.890000 1.565000 ;
      RECT  566.800000  2.255000  567.180000 2.635000 ;
      RECT  566.910000  0.295000  567.080000 0.725000 ;
      RECT  566.910000  0.725000  567.230000 1.065000 ;
      RECT  567.060000  1.065000  567.230000 1.835000 ;
      RECT  567.260000  0.085000  567.650000 0.545000 ;
      RECT  567.450000  0.725000  568.870000 0.895000 ;
      RECT  567.450000  0.895000  567.620000 1.655000 ;
      RECT  567.450000  1.655000  568.020000 1.965000 ;
      RECT  567.680000  2.165000  568.410000 2.415000 ;
      RECT  567.840000  1.065000  568.020000 1.475000 ;
      RECT  568.190000  1.235000  570.290000 1.405000 ;
      RECT  568.190000  1.405000  568.410000 1.915000 ;
      RECT  568.190000  1.915000  569.500000 2.085000 ;
      RECT  568.190000  2.085000  568.410000 2.165000 ;
      RECT  568.310000  0.305000  569.210000 0.475000 ;
      RECT  568.490000  0.895000  568.870000 1.015000 ;
      RECT  568.580000  1.575000  570.670000 1.745000 ;
      RECT  568.590000  2.255000  569.060000 2.635000 ;
      RECT  569.040000  0.475000  569.210000 1.235000 ;
      RECT  569.260000  2.085000  569.500000 2.375000 ;
      RECT  569.380000  0.735000  569.900000 1.005000 ;
      RECT  569.380000  1.005000  569.760000 1.065000 ;
      RECT  569.440000  0.085000  570.150000 0.565000 ;
      RECT  569.830000  1.945000  570.160000 2.635000 ;
      RECT  569.910000  1.175000  570.290000 1.235000 ;
      RECT  570.330000  0.350000  570.670000 0.680000 ;
      RECT  570.330000  1.745000  570.670000 1.765000 ;
      RECT  570.330000  1.765000  570.500000 2.375000 ;
      RECT  570.460000  0.680000  570.670000 1.575000 ;
      RECT  570.770000  1.915000  571.100000 2.425000 ;
      RECT  570.850000  0.345000  571.100000 1.055000 ;
      RECT  570.850000  1.055000  573.560000 1.275000 ;
      RECT  570.850000  1.275000  571.100000 1.915000 ;
      RECT  571.310000  0.085000  571.595000 0.545000 ;
      RECT  571.310000  1.835000  571.665000 2.635000 ;
      RECT  571.845000  0.265000  572.145000 0.715000 ;
      RECT  571.845000  0.715000  573.980000 0.885000 ;
      RECT  571.845000  1.470000  573.980000 1.640000 ;
      RECT  571.845000  1.640000  572.115000 2.465000 ;
      RECT  572.285000  1.810000  572.540000 2.635000 ;
      RECT  572.315000  0.085000  572.615000 0.545000 ;
      RECT  572.785000  0.265000  572.955000 0.715000 ;
      RECT  572.785000  1.640000  572.955000 2.465000 ;
      RECT  573.175000  0.085000  573.555000 0.545000 ;
      RECT  573.175000  1.810000  573.555000 2.635000 ;
      RECT  573.725000  0.265000  573.980000 0.715000 ;
      RECT  573.725000  1.640000  573.980000 2.465000 ;
      RECT  573.730000  0.885000  573.980000 1.470000 ;
      RECT  574.165000  0.085000  574.455000 0.810000 ;
      RECT  574.165000  1.470000  574.455000 2.635000 ;
      RECT  574.625000  0.985000  574.870000 1.625000 ;
      RECT  574.715000  0.345000  574.885000 0.635000 ;
      RECT  574.715000  0.635000  575.370000 0.805000 ;
      RECT  574.715000  1.795000  575.370000 1.965000 ;
      RECT  574.715000  1.965000  574.885000 2.465000 ;
      RECT  575.055000  0.085000  575.435000 0.465000 ;
      RECT  575.055000  2.135000  575.435000 2.635000 ;
      RECT  575.200000  0.805000  575.370000 1.070000 ;
      RECT  575.200000  1.070000  575.430000 1.400000 ;
      RECT  575.200000  1.400000  575.370000 1.795000 ;
      RECT  575.655000  0.345000  575.825000 1.685000 ;
      RECT  575.655000  1.685000  575.880000 2.465000 ;
      RECT  576.005000  0.955000  576.430000 1.325000 ;
      RECT  576.095000  1.495000  576.830000 1.665000 ;
      RECT  576.095000  1.665000  576.425000 2.415000 ;
      RECT  576.175000  0.345000  576.345000 0.615000 ;
      RECT  576.175000  0.615000  576.830000 0.765000 ;
      RECT  576.175000  0.765000  577.080000 0.785000 ;
      RECT  576.515000  0.085000  576.895000 0.445000 ;
      RECT  576.645000  1.835000  576.960000 2.635000 ;
      RECT  576.660000  0.785000  577.080000 1.095000 ;
      RECT  576.660000  1.095000  576.830000 1.495000 ;
      RECT  577.210000  1.355000  577.495000 2.005000 ;
      RECT  577.425000  0.705000  577.880000 1.035000 ;
      RECT  577.545000  0.365000  578.390000 0.535000 ;
      RECT  577.560000  2.255000  578.390000 2.425000 ;
      RECT  577.710000  1.035000  577.880000 1.415000 ;
      RECT  577.710000  1.415000  578.050000 1.995000 ;
      RECT  578.220000  0.535000  578.390000 0.995000 ;
      RECT  578.220000  0.995000  578.970000 1.325000 ;
      RECT  578.220000  1.325000  578.390000 2.255000 ;
      RECT  578.560000  0.085000  578.840000 0.825000 ;
      RECT  578.590000  2.135000  578.890000 2.635000 ;
      RECT  578.610000  1.535000  579.330000 1.865000 ;
      RECT  579.110000  0.415000  579.330000 0.825000 ;
      RECT  579.110000  1.865000  579.330000 2.435000 ;
      RECT  579.160000  0.825000  579.330000 0.995000 ;
      RECT  579.160000  0.995000  579.960000 1.325000 ;
      RECT  579.160000  1.325000  579.330000 1.535000 ;
      RECT  579.560000  0.085000  579.830000 0.825000 ;
      RECT  579.560000  1.495000  579.830000 2.635000 ;
      RECT  580.130000  0.415000  580.415000 2.455000 ;
      RECT  580.605000  0.085000  580.895000 0.810000 ;
      RECT  580.605000  1.470000  580.895000 2.635000 ;
      RECT  581.065000  0.985000  581.310000 1.625000 ;
      RECT  581.155000  0.345000  581.325000 0.635000 ;
      RECT  581.155000  0.635000  581.810000 0.805000 ;
      RECT  581.155000  1.795000  581.810000 1.965000 ;
      RECT  581.155000  1.965000  581.325000 2.465000 ;
      RECT  581.495000  0.085000  581.875000 0.465000 ;
      RECT  581.495000  2.135000  581.875000 2.635000 ;
      RECT  581.640000  0.805000  581.810000 1.070000 ;
      RECT  581.640000  1.070000  581.870000 1.400000 ;
      RECT  581.640000  1.400000  581.810000 1.795000 ;
      RECT  582.095000  0.345000  582.265000 1.685000 ;
      RECT  582.095000  1.685000  582.320000 2.465000 ;
      RECT  582.445000  0.955000  582.870000 1.325000 ;
      RECT  582.535000  1.495000  583.270000 1.665000 ;
      RECT  582.535000  1.665000  582.865000 2.415000 ;
      RECT  582.615000  0.345000  582.785000 0.615000 ;
      RECT  582.615000  0.615000  583.270000 0.765000 ;
      RECT  582.615000  0.765000  583.520000 0.785000 ;
      RECT  582.955000  0.085000  583.335000 0.445000 ;
      RECT  583.085000  1.835000  583.400000 2.635000 ;
      RECT  583.100000  0.785000  583.520000 1.095000 ;
      RECT  583.100000  1.095000  583.270000 1.495000 ;
      RECT  583.650000  1.355000  583.935000 2.005000 ;
      RECT  583.895000  0.705000  584.320000 1.035000 ;
      RECT  584.065000  0.365000  584.775000 0.535000 ;
      RECT  584.125000  2.255000  584.925000 2.425000 ;
      RECT  584.150000  1.035000  584.320000 1.415000 ;
      RECT  584.150000  1.415000  584.490000 1.995000 ;
      RECT  584.605000  0.535000  584.775000 0.995000 ;
      RECT  584.605000  0.995000  585.525000 1.165000 ;
      RECT  584.755000  1.165000  585.525000 1.325000 ;
      RECT  584.755000  1.325000  584.925000 2.255000 ;
      RECT  585.015000  0.085000  585.395000 0.825000 ;
      RECT  585.145000  2.135000  585.445000 2.635000 ;
      RECT  585.165000  1.535000  585.885000 1.865000 ;
      RECT  585.665000  0.415000  585.885000 0.825000 ;
      RECT  585.665000  1.865000  585.885000 2.435000 ;
      RECT  585.715000  0.825000  585.885000 0.995000 ;
      RECT  585.715000  0.995000  586.515000 1.325000 ;
      RECT  585.715000  1.325000  585.885000 1.535000 ;
      RECT  586.115000  0.085000  586.385000 0.825000 ;
      RECT  586.115000  1.495000  586.385000 2.635000 ;
      RECT  586.605000  0.415000  586.890000 0.825000 ;
      RECT  586.605000  1.495000  586.890000 2.455000 ;
      RECT  586.720000  0.825000  586.890000 0.995000 ;
      RECT  586.720000  0.995000  587.325000 1.325000 ;
      RECT  586.720000  1.325000  586.890000 1.495000 ;
      RECT  587.075000  0.085000  587.335000 0.550000 ;
      RECT  587.075000  1.755000  587.325000 2.635000 ;
      RECT  587.505000  0.085000  587.795000 0.810000 ;
      RECT  587.505000  1.470000  587.795000 2.635000 ;
      RECT  587.965000  0.985000  588.210000 1.625000 ;
      RECT  588.055000  0.345000  588.225000 0.635000 ;
      RECT  588.055000  0.635000  588.770000 0.805000 ;
      RECT  588.055000  1.795000  588.770000 1.965000 ;
      RECT  588.055000  1.965000  588.225000 2.465000 ;
      RECT  588.395000  0.085000  588.775000 0.465000 ;
      RECT  588.395000  2.135000  588.775000 2.635000 ;
      RECT  588.540000  0.805000  588.770000 1.795000 ;
      RECT  588.995000  0.345000  589.165000 2.465000 ;
      RECT  589.355000  0.955000  589.770000 1.325000 ;
      RECT  589.435000  1.495000  590.170000 1.665000 ;
      RECT  589.435000  1.665000  589.765000 2.415000 ;
      RECT  589.515000  0.345000  589.685000 0.615000 ;
      RECT  589.515000  0.615000  590.170000 0.765000 ;
      RECT  589.515000  0.765000  590.420000 0.785000 ;
      RECT  589.855000  0.085000  590.235000 0.445000 ;
      RECT  589.985000  1.835000  590.300000 2.635000 ;
      RECT  590.000000  0.785000  590.420000 1.095000 ;
      RECT  590.000000  1.095000  590.170000 1.495000 ;
      RECT  590.550000  1.355000  590.835000 2.005000 ;
      RECT  590.795000  0.705000  591.225000 1.035000 ;
      RECT  590.905000  2.255000  591.830000 2.425000 ;
      RECT  590.970000  0.365000  591.830000 0.535000 ;
      RECT  591.055000  1.035000  591.225000 1.415000 ;
      RECT  591.055000  1.415000  591.445000 1.995000 ;
      RECT  591.660000  0.535000  591.830000 0.995000 ;
      RECT  591.660000  0.995000  592.380000 1.325000 ;
      RECT  591.660000  1.325000  591.830000 2.255000 ;
      RECT  592.000000  0.085000  592.170000 0.610000 ;
      RECT  592.000000  2.135000  592.170000 2.635000 ;
      RECT  592.020000  1.535000  592.740000 1.865000 ;
      RECT  592.520000  1.865000  592.740000 2.435000 ;
      RECT  592.550000  0.415000  592.740000 0.995000 ;
      RECT  592.550000  0.995000  593.370000 1.325000 ;
      RECT  592.550000  1.325000  592.740000 1.535000 ;
      RECT  592.970000  0.085000  593.255000 0.715000 ;
      RECT  592.970000  1.495000  593.255000 2.635000 ;
      RECT  593.475000  0.415000  593.775000 0.745000 ;
      RECT  593.475000  1.495000  593.775000 2.455000 ;
      RECT  593.590000  0.745000  593.775000 0.995000 ;
      RECT  593.590000  0.995000  595.115000 1.325000 ;
      RECT  593.590000  1.325000  593.775000 1.495000 ;
      RECT  593.945000  0.085000  594.195000 0.825000 ;
      RECT  593.945000  1.495000  594.195000 2.635000 ;
      RECT  594.415000  0.385000  594.685000 0.995000 ;
      RECT  594.415000  1.325000  594.685000 2.455000 ;
      RECT  594.885000  0.085000  595.055000 0.715000 ;
      RECT  594.885000  1.495000  595.055000 2.635000 ;
      RECT  595.325000  0.085000  595.615000 0.810000 ;
      RECT  595.325000  1.470000  595.615000 2.635000 ;
      RECT  595.785000  1.055000  596.305000 1.615000 ;
      RECT  595.785000  1.785000  596.645000 2.005000 ;
      RECT  595.785000  2.005000  596.080000 2.465000 ;
      RECT  595.795000  0.255000  596.080000 0.715000 ;
      RECT  595.795000  0.715000  596.645000 0.885000 ;
      RECT  596.300000  0.085000  596.515000 0.545000 ;
      RECT  596.300000  2.175000  596.515000 2.635000 ;
      RECT  596.475000  0.885000  596.645000 0.995000 ;
      RECT  596.475000  0.995000  596.780000 1.325000 ;
      RECT  596.475000  1.325000  596.645000 1.785000 ;
      RECT  596.685000  0.255000  597.120000 0.545000 ;
      RECT  596.685000  2.175000  597.120000 2.465000 ;
      RECT  596.950000  0.545000  597.120000 1.075000 ;
      RECT  596.950000  1.075000  597.700000 1.275000 ;
      RECT  596.950000  1.275000  597.120000 2.175000 ;
      RECT  597.315000  0.255000  597.540000 0.735000 ;
      RECT  597.315000  0.735000  598.310000 0.905000 ;
      RECT  597.315000  1.575000  598.310000 1.745000 ;
      RECT  597.315000  1.745000  597.540000 2.430000 ;
      RECT  597.845000  0.085000  598.255000 0.565000 ;
      RECT  597.845000  1.915000  598.215000 2.635000 ;
      RECT  598.100000  0.905000  598.310000 0.995000 ;
      RECT  598.100000  0.995000  598.430000 1.325000 ;
      RECT  598.100000  1.325000  598.310000 1.575000 ;
      RECT  598.530000  0.255000  598.820000 0.825000 ;
      RECT  598.560000  1.495000  598.820000 2.465000 ;
      RECT  598.650000  0.825000  598.820000 1.495000 ;
      RECT  599.005000  0.085000  599.295000 0.810000 ;
      RECT  599.005000  1.470000  599.295000 2.635000 ;
      RECT  599.465000  1.055000  599.985000 1.615000 ;
      RECT  599.465000  1.785000  600.325000 2.005000 ;
      RECT  599.465000  2.005000  599.760000 2.465000 ;
      RECT  599.475000  0.255000  599.760000 0.715000 ;
      RECT  599.475000  0.715000  600.325000 0.885000 ;
      RECT  599.980000  0.085000  600.195000 0.545000 ;
      RECT  599.980000  2.175000  600.195000 2.635000 ;
      RECT  600.155000  0.885000  600.325000 0.995000 ;
      RECT  600.155000  0.995000  600.460000 1.325000 ;
      RECT  600.155000  1.325000  600.325000 1.785000 ;
      RECT  600.365000  0.255000  600.800000 0.545000 ;
      RECT  600.365000  2.175000  600.800000 2.465000 ;
      RECT  600.630000  0.545000  600.800000 1.075000 ;
      RECT  600.630000  1.075000  601.475000 1.275000 ;
      RECT  600.630000  1.275000  600.800000 2.175000 ;
      RECT  600.995000  0.510000  601.220000 0.735000 ;
      RECT  600.995000  0.735000  601.990000 0.905000 ;
      RECT  600.995000  1.575000  601.990000 1.745000 ;
      RECT  600.995000  1.745000  601.220000 2.080000 ;
      RECT  601.525000  0.085000  601.935000 0.565000 ;
      RECT  601.525000  1.915000  601.895000 2.635000 ;
      RECT  601.780000  0.905000  601.990000 0.995000 ;
      RECT  601.780000  0.995000  602.070000 1.325000 ;
      RECT  601.780000  1.325000  601.990000 1.575000 ;
      RECT  602.160000  0.255000  602.490000 0.825000 ;
      RECT  602.160000  1.495000  602.490000 2.465000 ;
      RECT  602.240000  0.825000  602.490000 1.495000 ;
      RECT  602.685000  0.085000  602.975000 0.810000 ;
      RECT  602.685000  1.470000  602.975000 2.635000 ;
      RECT  603.145000  1.055000  603.665000 1.615000 ;
      RECT  603.145000  1.785000  604.005000 2.005000 ;
      RECT  603.145000  2.005000  603.440000 2.465000 ;
      RECT  603.155000  0.255000  603.440000 0.715000 ;
      RECT  603.155000  0.715000  604.005000 0.885000 ;
      RECT  603.660000  0.085000  603.875000 0.545000 ;
      RECT  603.665000  2.175000  603.915000 2.635000 ;
      RECT  603.835000  0.885000  604.005000 0.995000 ;
      RECT  603.835000  0.995000  604.460000 1.325000 ;
      RECT  603.835000  1.325000  604.005000 1.785000 ;
      RECT  604.365000  0.255000  604.800000 0.545000 ;
      RECT  604.365000  2.175000  604.800000 2.465000 ;
      RECT  604.630000  0.545000  604.800000 1.075000 ;
      RECT  604.630000  1.075000  605.535000 1.275000 ;
      RECT  604.630000  1.275000  604.800000 2.175000 ;
      RECT  604.970000  0.510000  605.200000 0.735000 ;
      RECT  604.970000  0.735000  606.080000 0.905000 ;
      RECT  604.970000  1.575000  606.080000 1.745000 ;
      RECT  604.970000  1.745000  605.190000 2.080000 ;
      RECT  605.750000  0.085000  606.080000 0.565000 ;
      RECT  605.750000  1.915000  606.080000 2.635000 ;
      RECT  605.870000  0.905000  606.080000 0.995000 ;
      RECT  605.870000  0.995000  606.215000 1.325000 ;
      RECT  605.870000  1.325000  606.080000 1.575000 ;
      RECT  606.250000  0.255000  606.655000 0.825000 ;
      RECT  606.250000  1.495000  606.655000 2.465000 ;
      RECT  606.385000  0.825000  606.655000 1.495000 ;
      RECT  606.825000  0.085000  607.115000 0.810000 ;
      RECT  606.825000  1.470000  607.115000 2.635000 ;
      RECT  607.285000  0.280000  607.545000 0.615000 ;
      RECT  607.285000  0.615000  608.435000 0.825000 ;
      RECT  607.285000  0.995000  607.555000 1.615000 ;
      RECT  607.285000  1.785000  607.990000 2.005000 ;
      RECT  607.285000  2.005000  607.545000 2.465000 ;
      RECT  607.715000  0.085000  608.095000 0.445000 ;
      RECT  607.715000  2.175000  608.090000 2.635000 ;
      RECT  607.725000  0.825000  607.990000 1.785000 ;
      RECT  608.160000  1.075000  608.490000 1.630000 ;
      RECT  608.265000  0.255000  609.375000 0.465000 ;
      RECT  608.265000  0.465000  608.435000 0.615000 ;
      RECT  608.315000  1.800000  609.105000 2.005000 ;
      RECT  608.315000  2.005000  608.570000 2.460000 ;
      RECT  608.660000  0.635000  608.990000 1.075000 ;
      RECT  608.660000  1.075000  609.945000 1.325000 ;
      RECT  608.660000  1.325000  609.105000 1.800000 ;
      RECT  608.740000  2.175000  609.100000 2.635000 ;
      RECT  609.160000  0.465000  609.375000 0.735000 ;
      RECT  609.160000  0.735000  610.285000 0.905000 ;
      RECT  609.325000  1.495000  610.785000 2.465000 ;
      RECT  609.545000  0.085000  610.285000 0.565000 ;
      RECT  610.115000  0.905000  610.285000 0.995000 ;
      RECT  610.115000  0.995000  610.345000 1.325000 ;
      RECT  610.455000  0.255000  610.785000 0.825000 ;
      RECT  610.515000  0.825000  610.785000 1.495000 ;
      RECT  610.965000  0.085000  611.255000 0.810000 ;
      RECT  610.965000  1.470000  611.255000 2.635000 ;
      RECT  611.425000  0.280000  611.685000 2.465000 ;
      RECT  611.855000  0.085000  612.240000 0.595000 ;
      RECT  611.855000  0.765000  612.115000 1.675000 ;
      RECT  611.855000  1.845000  612.340000 2.635000 ;
      RECT  612.285000  0.765000  612.640000 1.275000 ;
      RECT  612.410000  0.255000  613.170000 0.595000 ;
      RECT  612.560000  1.445000  613.155000 1.765000 ;
      RECT  612.560000  1.765000  612.850000 2.465000 ;
      RECT  612.890000  0.595000  613.170000 1.025000 ;
      RECT  612.890000  1.025000  614.555000 1.275000 ;
      RECT  612.890000  1.275000  613.155000 1.445000 ;
      RECT  613.040000  1.935000  614.715000 2.105000 ;
      RECT  613.040000  2.105000  613.250000 2.465000 ;
      RECT  613.325000  1.445000  615.800000 1.625000 ;
      RECT  613.325000  1.625000  615.335000 1.765000 ;
      RECT  613.340000  0.255000  613.660000 0.655000 ;
      RECT  613.340000  0.655000  614.715000 0.855000 ;
      RECT  613.420000  2.275000  613.800000 2.635000 ;
      RECT  613.830000  0.085000  614.210000 0.485000 ;
      RECT  614.020000  2.105000  614.715000 2.295000 ;
      RECT  614.020000  2.295000  615.765000 2.465000 ;
      RECT  614.430000  0.275000  615.740000 0.465000 ;
      RECT  614.430000  0.465000  614.715000 0.655000 ;
      RECT  614.835000  1.025000  615.295000 1.275000 ;
      RECT  614.885000  0.635000  615.800000 0.855000 ;
      RECT  614.935000  1.765000  615.335000 2.125000 ;
      RECT  615.505000  1.795000  615.765000 2.295000 ;
      RECT  615.570000  0.855000  615.800000 1.445000 ;
      RECT  616.025000  0.085000  616.315000 0.810000 ;
      RECT  616.025000  1.470000  616.315000 2.635000 ;
      RECT  616.485000  0.280000  616.745000 0.665000 ;
      RECT  616.485000  0.665000  616.720000 1.765000 ;
      RECT  616.485000  1.765000  616.745000 2.465000 ;
      RECT  616.890000  0.765000  617.230000 1.675000 ;
      RECT  616.915000  0.085000  617.380000 0.595000 ;
      RECT  616.915000  1.845000  617.380000 2.635000 ;
      RECT  617.400000  0.765000  617.780000 1.425000 ;
      RECT  617.600000  0.255000  618.225000 0.595000 ;
      RECT  617.600000  1.595000  618.225000 1.765000 ;
      RECT  617.600000  1.765000  617.855000 2.465000 ;
      RECT  617.950000  0.595000  618.225000 1.025000 ;
      RECT  617.950000  1.025000  620.560000 1.275000 ;
      RECT  617.950000  1.275000  618.225000 1.595000 ;
      RECT  618.065000  1.935000  622.685000 2.105000 ;
      RECT  618.065000  2.105000  618.310000 2.465000 ;
      RECT  618.395000  0.255000  618.725000 0.655000 ;
      RECT  618.395000  0.655000  620.725000 0.855000 ;
      RECT  618.395000  1.445000  622.735000 1.725000 ;
      RECT  618.395000  1.895000  622.685000 1.935000 ;
      RECT  618.480000  2.275000  618.860000 2.635000 ;
      RECT  618.895000  0.085000  619.275000 0.485000 ;
      RECT  619.080000  2.105000  619.250000 2.465000 ;
      RECT  619.470000  2.275000  619.800000 2.635000 ;
      RECT  619.495000  0.275000  619.665000 0.655000 ;
      RECT  619.835000  0.085000  620.215000 0.485000 ;
      RECT  620.020000  2.105000  622.685000 2.465000 ;
      RECT  620.435000  0.255000  622.685000 0.445000 ;
      RECT  620.435000  0.445000  620.725000 0.655000 ;
      RECT  620.730000  1.025000  622.335000 1.275000 ;
      RECT  620.895000  0.615000  622.735000 0.855000 ;
      RECT  622.505000  0.855000  622.735000 1.445000 ;
      RECT  622.925000  0.085000  623.215000 0.810000 ;
      RECT  622.925000  1.470000  623.215000 2.635000 ;
      RECT  623.385000  0.085000  623.745000 0.825000 ;
      RECT  623.385000  0.995000  623.730000 1.615000 ;
      RECT  623.385000  1.785000  623.745000 2.635000 ;
      RECT  623.950000  0.280000  624.150000 1.615000 ;
      RECT  623.965000  1.615000  624.150000 2.465000 ;
      RECT  624.320000  0.085000  624.705000 0.445000 ;
      RECT  624.320000  0.620000  624.705000 0.995000 ;
      RECT  624.320000  0.995000  624.830000 1.325000 ;
      RECT  624.320000  1.325000  624.705000 1.695000 ;
      RECT  624.320000  1.865000  624.705000 2.635000 ;
      RECT  624.875000  0.255000  625.435000 0.825000 ;
      RECT  624.875000  1.495000  625.275000 2.465000 ;
      RECT  625.050000  0.825000  625.435000 1.025000 ;
      RECT  625.050000  1.025000  630.175000 1.275000 ;
      RECT  625.050000  1.275000  625.275000 1.495000 ;
      RECT  625.445000  1.445000  634.225000 1.725000 ;
      RECT  625.445000  1.895000  634.225000 2.065000 ;
      RECT  625.445000  2.065000  625.695000 2.465000 ;
      RECT  625.605000  0.255000  625.985000 0.655000 ;
      RECT  625.605000  0.655000  630.355000 0.855000 ;
      RECT  625.865000  2.235000  626.295000 2.635000 ;
      RECT  626.155000  0.085000  626.585000 0.485000 ;
      RECT  626.515000  2.065000  626.685000 2.465000 ;
      RECT  626.805000  0.275000  627.025000 0.655000 ;
      RECT  626.905000  2.235000  627.335000 2.635000 ;
      RECT  627.195000  0.085000  627.625000 0.485000 ;
      RECT  627.555000  2.065000  627.725000 2.465000 ;
      RECT  627.845000  0.255000  628.065000 0.655000 ;
      RECT  627.945000  2.235000  628.375000 2.635000 ;
      RECT  628.235000  0.085000  628.665000 0.485000 ;
      RECT  628.595000  2.065000  628.765000 2.465000 ;
      RECT  628.885000  0.275000  629.105000 0.655000 ;
      RECT  628.985000  2.235000  629.415000 2.635000 ;
      RECT  629.275000  0.085000  629.705000 0.485000 ;
      RECT  629.635000  2.065000  634.225000 2.465000 ;
      RECT  629.925000  0.255000  634.225000 0.445000 ;
      RECT  629.925000  0.445000  630.355000 0.655000 ;
      RECT  630.425000  1.025000  633.755000 1.275000 ;
      RECT  630.525000  0.615000  634.225000 0.855000 ;
      RECT  633.975000  0.855000  634.225000 1.445000 ;
      RECT  634.425000  0.085000  634.715000 0.810000 ;
      RECT  634.425000  1.470000  634.715000 2.635000 ;
      RECT  634.885000  0.255000  635.170000 0.615000 ;
      RECT  634.885000  0.615000  636.400000 0.785000 ;
      RECT  634.885000  0.955000  635.310000 1.725000 ;
      RECT  634.885000  1.895000  635.720000 2.065000 ;
      RECT  634.885000  2.065000  635.170000 2.465000 ;
      RECT  635.340000  0.085000  636.390000 0.445000 ;
      RECT  635.340000  2.235000  635.720000 2.635000 ;
      RECT  635.535000  0.785000  636.400000 0.805000 ;
      RECT  635.535000  1.440000  636.400000 1.615000 ;
      RECT  635.535000  1.615000  635.720000 1.895000 ;
      RECT  635.920000  0.805000  636.400000 1.440000 ;
      RECT  636.200000  1.785000  637.475000 2.465000 ;
      RECT  636.770000  0.255000  637.475000 0.595000 ;
      RECT  636.770000  0.595000  637.010000 1.785000 ;
      RECT  637.230000  0.765000  637.475000 1.615000 ;
      RECT  637.645000  0.085000  637.935000 0.810000 ;
      RECT  637.645000  1.470000  637.935000 2.635000 ;
      RECT  638.105000  0.255000  638.365000 0.655000 ;
      RECT  638.105000  0.655000  638.910000 0.825000 ;
      RECT  638.105000  0.995000  638.345000 1.385000 ;
      RECT  638.105000  1.555000  638.965000 1.725000 ;
      RECT  638.105000  1.725000  638.365000 2.465000 ;
      RECT  638.515000  0.825000  638.910000 0.995000 ;
      RECT  638.515000  0.995000  640.200000 1.275000 ;
      RECT  638.515000  1.275000  638.965000 1.555000 ;
      RECT  638.535000  0.085000  638.915000 0.485000 ;
      RECT  638.535000  1.895000  638.965000 2.635000 ;
      RECT  639.085000  0.255000  639.400000 0.655000 ;
      RECT  639.085000  0.655000  640.290000 0.825000 ;
      RECT  639.190000  1.445000  639.945000 1.865000 ;
      RECT  639.190000  1.865000  640.885000 2.085000 ;
      RECT  639.190000  2.085000  639.360000 2.465000 ;
      RECT  639.530000  2.255000  640.495000 2.635000 ;
      RECT  639.620000  0.085000  639.950000 0.485000 ;
      RECT  640.120000  0.255000  641.455000 0.425000 ;
      RECT  640.120000  0.425000  640.290000 0.655000 ;
      RECT  640.165000  1.445000  641.555000 1.695000 ;
      RECT  640.465000  0.595000  640.835000 1.445000 ;
      RECT  640.715000  2.085000  640.885000 2.465000 ;
      RECT  641.005000  1.075000  641.555000 1.275000 ;
      RECT  641.055000  1.695000  641.555000 2.465000 ;
      RECT  641.185000  0.425000  641.455000 0.775000 ;
      RECT  641.785000  0.085000  642.075000 0.810000 ;
      RECT  641.785000  1.470000  642.075000 2.635000 ;
      RECT  642.245000  0.255000  642.505000 0.655000 ;
      RECT  642.245000  0.655000  643.055000 0.825000 ;
      RECT  642.245000  0.995000  642.505000 1.325000 ;
      RECT  642.245000  1.495000  643.055000 1.665000 ;
      RECT  642.245000  1.665000  642.505000 2.465000 ;
      RECT  642.675000  0.085000  643.055000 0.485000 ;
      RECT  642.675000  0.825000  643.055000 0.995000 ;
      RECT  642.675000  0.995000  645.480000 1.325000 ;
      RECT  642.675000  1.325000  643.055000 1.495000 ;
      RECT  642.675000  1.835000  643.055000 2.635000 ;
      RECT  643.225000  0.255000  643.545000 0.655000 ;
      RECT  643.225000  0.655000  645.455000 0.825000 ;
      RECT  643.225000  1.495000  645.480000 1.665000 ;
      RECT  643.225000  1.665000  643.500000 2.465000 ;
      RECT  643.670000  1.835000  644.050000 2.635000 ;
      RECT  643.765000  0.085000  644.095000 0.485000 ;
      RECT  644.270000  1.665000  644.440000 2.465000 ;
      RECT  644.315000  0.255000  644.485000 0.655000 ;
      RECT  644.610000  1.835000  645.050000 2.635000 ;
      RECT  644.705000  0.085000  645.035000 0.485000 ;
      RECT  645.270000  1.665000  645.480000 2.295000 ;
      RECT  645.270000  2.295000  647.360000 2.465000 ;
      RECT  645.285000  0.255000  647.595000 0.450000 ;
      RECT  645.285000  0.450000  645.455000 0.655000 ;
      RECT  645.650000  0.620000  646.970000 1.480000 ;
      RECT  645.650000  1.480000  646.030000 2.075000 ;
      RECT  646.250000  1.650000  646.420000 2.295000 ;
      RECT  646.590000  1.480000  646.970000 2.075000 ;
      RECT  647.140000  0.620000  647.575000 1.325000 ;
      RECT  647.190000  1.650000  647.360000 2.295000 ;
      RECT  647.765000  0.085000  648.055000 0.810000 ;
      RECT  647.765000  1.470000  648.055000 2.635000 ;
      RECT  648.230000  0.255000  648.485000 0.655000 ;
      RECT  648.230000  0.655000  649.035000 0.825000 ;
      RECT  648.230000  0.995000  648.485000 1.325000 ;
      RECT  648.230000  1.495000  649.035000 1.665000 ;
      RECT  648.230000  1.665000  648.485000 2.465000 ;
      RECT  648.655000  0.085000  649.035000 0.485000 ;
      RECT  648.655000  0.825000  649.035000 0.995000 ;
      RECT  648.655000  0.995000  653.115000 1.325000 ;
      RECT  648.655000  1.325000  649.035000 1.495000 ;
      RECT  648.655000  1.835000  649.035000 2.635000 ;
      RECT  649.205000  0.255000  649.525000 0.655000 ;
      RECT  649.205000  0.655000  653.340000 0.825000 ;
      RECT  649.205000  1.495000  653.340000 1.665000 ;
      RECT  649.205000  1.665000  649.480000 2.465000 ;
      RECT  649.650000  1.835000  650.030000 2.635000 ;
      RECT  649.745000  0.085000  650.075000 0.485000 ;
      RECT  650.250000  1.665000  650.420000 2.465000 ;
      RECT  650.295000  0.255000  650.465000 0.655000 ;
      RECT  650.590000  1.835000  650.970000 2.635000 ;
      RECT  650.685000  0.085000  651.015000 0.485000 ;
      RECT  651.190000  1.665000  651.360000 2.465000 ;
      RECT  651.235000  0.255000  651.405000 0.655000 ;
      RECT  651.530000  1.835000  651.910000 2.635000 ;
      RECT  651.625000  0.085000  651.955000 0.485000 ;
      RECT  652.130000  1.665000  652.300000 2.465000 ;
      RECT  652.175000  0.255000  652.345000 0.655000 ;
      RECT  652.470000  1.835000  652.870000 2.635000 ;
      RECT  652.565000  0.085000  652.905000 0.485000 ;
      RECT  653.090000  1.665000  653.340000 2.295000 ;
      RECT  653.090000  2.295000  657.235000 2.465000 ;
      RECT  653.125000  0.255000  657.235000 0.450000 ;
      RECT  653.125000  0.450000  653.340000 0.655000 ;
      RECT  653.285000  0.995000  656.790000 1.285000 ;
      RECT  653.510000  0.620000  657.235000 0.825000 ;
      RECT  653.510000  1.455000  657.235000 1.625000 ;
      RECT  653.510000  1.625000  653.890000 2.125000 ;
      RECT  654.110000  1.795000  654.280000 2.295000 ;
      RECT  654.450000  1.625000  654.830000 2.125000 ;
      RECT  655.050000  1.795000  655.220000 2.295000 ;
      RECT  655.390000  1.625000  655.770000 2.125000 ;
      RECT  655.990000  1.795000  656.160000 2.295000 ;
      RECT  656.330000  1.625000  656.710000 2.125000 ;
      RECT  656.930000  1.795000  657.235000 2.295000 ;
      RECT  657.010000  0.825000  657.235000 1.455000 ;
      RECT  657.425000  0.085000  657.715000 0.810000 ;
      RECT  657.425000  1.470000  657.715000 2.635000 ;
      RECT  657.885000  0.255000  658.145000 0.655000 ;
      RECT  657.885000  0.655000  659.490000 0.825000 ;
      RECT  657.885000  0.995000  658.395000 1.725000 ;
      RECT  657.885000  1.895000  659.490000 2.065000 ;
      RECT  657.885000  2.065000  658.145000 2.465000 ;
      RECT  658.315000  0.085000  659.300000 0.485000 ;
      RECT  658.315000  2.235000  659.540000 2.635000 ;
      RECT  658.565000  0.825000  659.490000 1.895000 ;
      RECT  659.780000  0.255000  660.425000 0.805000 ;
      RECT  659.780000  0.805000  659.955000 2.125000 ;
      RECT  659.780000  2.125000  660.425000 2.465000 ;
      RECT  660.185000  0.975000  660.425000 1.955000 ;
      RECT  660.645000  0.085000  660.935000 0.810000 ;
      RECT  660.645000  1.470000  660.935000 2.635000 ;
      RECT  661.105000  0.255000  661.365000 0.655000 ;
      RECT  661.105000  0.655000  661.945000 0.825000 ;
      RECT  661.105000  0.995000  661.350000 1.615000 ;
      RECT  661.105000  1.785000  661.945000 1.955000 ;
      RECT  661.105000  1.955000  661.365000 2.465000 ;
      RECT  661.520000  0.825000  661.945000 0.995000 ;
      RECT  661.520000  0.995000  663.125000 1.325000 ;
      RECT  661.520000  1.325000  661.945000 1.785000 ;
      RECT  661.535000  0.085000  661.945000 0.485000 ;
      RECT  661.535000  2.125000  661.945000 2.635000 ;
      RECT  662.165000  0.255000  662.360000 0.655000 ;
      RECT  662.165000  0.655000  663.495000 0.825000 ;
      RECT  662.165000  1.555000  663.375000 1.725000 ;
      RECT  662.165000  1.725000  662.405000 2.465000 ;
      RECT  662.530000  0.085000  662.900000 0.485000 ;
      RECT  662.625000  1.895000  662.955000 2.635000 ;
      RECT  663.160000  0.255000  664.550000 0.425000 ;
      RECT  663.160000  0.425000  663.495000 0.655000 ;
      RECT  663.205000  1.725000  663.375000 2.295000 ;
      RECT  663.205000  2.295000  664.550000 2.465000 ;
      RECT  663.665000  0.595000  664.095000 2.125000 ;
      RECT  664.265000  0.425000  664.550000 0.595000 ;
      RECT  664.265000  0.765000  664.555000 1.615000 ;
      RECT  664.265000  1.785000  664.550000 2.295000 ;
      RECT  664.785000  0.085000  665.075000 0.810000 ;
      RECT  664.785000  1.470000  665.075000 2.635000 ;
      RECT  665.245000  0.255000  665.505000 0.655000 ;
      RECT  665.245000  0.655000  665.905000 0.825000 ;
      RECT  665.245000  0.995000  665.490000 1.615000 ;
      RECT  665.245000  1.785000  666.085000 1.955000 ;
      RECT  665.245000  1.955000  665.505000 2.465000 ;
      RECT  665.660000  0.825000  665.905000 0.995000 ;
      RECT  665.660000  0.995000  668.480000 1.325000 ;
      RECT  665.660000  1.325000  666.085000 1.785000 ;
      RECT  665.675000  0.085000  666.055000 0.485000 ;
      RECT  665.675000  2.125000  666.085000 2.635000 ;
      RECT  666.295000  0.255000  666.465000 0.655000 ;
      RECT  666.295000  0.655000  668.480000 0.825000 ;
      RECT  666.335000  1.555000  668.455000 1.725000 ;
      RECT  666.335000  1.725000  666.545000 2.465000 ;
      RECT  666.635000  0.085000  667.015000 0.485000 ;
      RECT  666.765000  1.895000  667.095000 2.635000 ;
      RECT  667.235000  0.255000  667.405000 0.655000 ;
      RECT  667.315000  1.725000  667.485000 2.465000 ;
      RECT  667.575000  0.085000  667.965000 0.485000 ;
      RECT  667.705000  1.895000  668.065000 2.635000 ;
      RECT  668.145000  0.255000  670.570000 0.465000 ;
      RECT  668.145000  0.465000  668.480000 0.655000 ;
      RECT  668.285000  1.725000  668.455000 2.295000 ;
      RECT  668.285000  2.295000  670.570000 2.465000 ;
      RECT  668.650000  0.635000  670.570000 0.850000 ;
      RECT  668.650000  0.850000  669.190000 1.445000 ;
      RECT  668.650000  1.445000  669.970000 1.615000 ;
      RECT  668.650000  1.615000  669.030000 2.125000 ;
      RECT  669.250000  1.785000  669.420000 2.295000 ;
      RECT  669.370000  1.020000  670.570000 1.275000 ;
      RECT  669.590000  1.615000  669.970000 2.125000 ;
      RECT  670.190000  1.445000  670.570000 2.295000 ;
      RECT  670.765000  0.085000  671.055000 0.810000 ;
      RECT  670.765000  1.470000  671.055000 2.635000 ;
      RECT  671.225000  0.255000  671.485000 0.655000 ;
      RECT  671.225000  0.655000  671.885000 0.825000 ;
      RECT  671.225000  0.995000  671.470000 1.615000 ;
      RECT  671.225000  1.785000  672.065000 1.955000 ;
      RECT  671.225000  1.955000  671.485000 2.465000 ;
      RECT  671.640000  0.825000  671.885000 0.995000 ;
      RECT  671.640000  0.995000  676.340000 1.325000 ;
      RECT  671.640000  1.325000  672.065000 1.785000 ;
      RECT  671.655000  0.085000  672.035000 0.485000 ;
      RECT  671.655000  2.125000  672.065000 2.635000 ;
      RECT  672.275000  0.255000  672.445000 0.655000 ;
      RECT  672.275000  0.655000  676.340000 0.825000 ;
      RECT  672.315000  1.555000  676.340000 1.725000 ;
      RECT  672.315000  1.725000  672.525000 2.465000 ;
      RECT  672.615000  0.085000  672.995000 0.485000 ;
      RECT  672.745000  1.895000  673.075000 2.635000 ;
      RECT  673.215000  0.255000  673.385000 0.655000 ;
      RECT  673.295000  1.725000  673.465000 2.465000 ;
      RECT  673.555000  0.085000  673.935000 0.485000 ;
      RECT  673.685000  1.895000  674.015000 2.635000 ;
      RECT  674.155000  0.255000  674.325000 0.655000 ;
      RECT  674.235000  1.725000  674.405000 2.465000 ;
      RECT  674.495000  0.085000  674.875000 0.485000 ;
      RECT  674.625000  1.895000  674.955000 2.635000 ;
      RECT  675.095000  0.255000  675.265000 0.655000 ;
      RECT  675.175000  1.725000  675.345000 2.465000 ;
      RECT  675.435000  0.085000  675.825000 0.485000 ;
      RECT  675.565000  1.895000  675.895000 2.635000 ;
      RECT  675.995000  0.255000  680.235000 0.465000 ;
      RECT  675.995000  0.465000  676.340000 0.655000 ;
      RECT  676.115000  1.725000  676.340000 2.295000 ;
      RECT  676.115000  2.295000  680.235000 2.465000 ;
      RECT  676.510000  0.635000  680.235000 0.850000 ;
      RECT  676.510000  0.850000  676.940000 1.445000 ;
      RECT  676.510000  1.445000  679.710000 1.615000 ;
      RECT  676.510000  1.615000  676.890000 2.125000 ;
      RECT  677.110000  1.785000  677.280000 2.295000 ;
      RECT  677.160000  1.020000  680.190000 1.275000 ;
      RECT  677.450000  1.615000  677.830000 2.125000 ;
      RECT  678.050000  1.785000  678.220000 2.295000 ;
      RECT  678.390000  1.615000  678.770000 2.125000 ;
      RECT  678.990000  1.785000  679.160000 2.295000 ;
      RECT  679.330000  1.615000  679.710000 2.125000 ;
      RECT  679.930000  1.445000  680.235000 2.295000 ;
      RECT  680.425000  0.085000  680.715000 0.810000 ;
      RECT  680.425000  1.470000  680.715000 2.635000 ;
      RECT  680.895000  1.075000  681.450000 1.315000 ;
      RECT  681.120000  0.085000  681.350000 0.905000 ;
      RECT  681.140000  1.495000  681.350000 2.635000 ;
      RECT  681.570000  0.255000  682.085000 0.885000 ;
      RECT  681.570000  1.485000  682.085000 2.465000 ;
      RECT  681.795000  0.885000  682.085000 1.485000 ;
      RECT  682.265000  0.085000  682.555000 0.810000 ;
      RECT  682.265000  1.470000  682.555000 2.635000 ;
      RECT  682.725000  0.715000  688.960000 0.905000 ;
      RECT  682.725000  0.905000  683.150000 1.495000 ;
      RECT  682.725000  1.495000  688.960000 1.665000 ;
      RECT  682.895000  0.085000  683.150000 0.545000 ;
      RECT  682.895000  1.835000  683.150000 2.635000 ;
      RECT  683.320000  0.255000  683.700000 0.715000 ;
      RECT  683.320000  1.075000  688.440000 1.325000 ;
      RECT  683.320000  1.665000  683.700000 2.465000 ;
      RECT  683.920000  0.085000  684.090000 0.545000 ;
      RECT  683.920000  1.835000  684.090000 2.635000 ;
      RECT  684.260000  0.255000  684.640000 0.715000 ;
      RECT  684.260000  1.665000  684.640000 2.465000 ;
      RECT  684.860000  0.085000  685.030000 0.545000 ;
      RECT  684.860000  1.835000  685.030000 2.635000 ;
      RECT  685.200000  0.255000  685.580000 0.715000 ;
      RECT  685.200000  1.665000  685.580000 2.465000 ;
      RECT  685.800000  0.085000  685.970000 0.545000 ;
      RECT  685.800000  1.835000  685.970000 2.635000 ;
      RECT  686.140000  0.255000  686.520000 0.715000 ;
      RECT  686.140000  1.665000  686.520000 2.465000 ;
      RECT  686.740000  0.085000  686.910000 0.545000 ;
      RECT  686.740000  1.835000  686.910000 2.635000 ;
      RECT  687.080000  0.255000  687.460000 0.715000 ;
      RECT  687.080000  1.665000  687.460000 2.465000 ;
      RECT  687.680000  0.085000  687.850000 0.545000 ;
      RECT  687.680000  1.835000  687.850000 2.635000 ;
      RECT  688.020000  0.255000  688.400000 0.715000 ;
      RECT  688.020000  1.665000  688.400000 2.465000 ;
      RECT  688.600000  0.085000  688.870000 0.545000 ;
      RECT  688.610000  0.905000  688.960000 1.495000 ;
      RECT  688.615000  1.835000  688.870000 2.635000 ;
      RECT  689.165000  0.085000  689.455000 0.810000 ;
      RECT  689.165000  1.470000  689.455000 2.635000 ;
      RECT  689.625000  1.075000  695.665000 1.315000 ;
      RECT  689.720000  0.085000  689.950000 0.885000 ;
      RECT  689.740000  1.485000  689.950000 2.635000 ;
      RECT  690.120000  0.255000  690.500000 0.715000 ;
      RECT  690.120000  0.715000  697.080000 0.905000 ;
      RECT  690.120000  1.495000  697.080000 1.665000 ;
      RECT  690.120000  1.665000  690.500000 2.465000 ;
      RECT  690.720000  0.085000  690.890000 0.545000 ;
      RECT  690.720000  1.835000  690.890000 2.635000 ;
      RECT  691.060000  0.255000  691.440000 0.715000 ;
      RECT  691.060000  1.665000  691.440000 2.465000 ;
      RECT  691.660000  0.085000  691.830000 0.545000 ;
      RECT  691.660000  1.835000  691.830000 2.635000 ;
      RECT  692.000000  0.255000  692.380000 0.715000 ;
      RECT  692.000000  1.665000  692.380000 2.465000 ;
      RECT  692.600000  0.085000  692.770000 0.545000 ;
      RECT  692.600000  1.835000  692.770000 2.635000 ;
      RECT  692.940000  0.255000  693.320000 0.715000 ;
      RECT  692.940000  1.665000  693.320000 2.465000 ;
      RECT  693.540000  0.085000  693.710000 0.545000 ;
      RECT  693.540000  1.835000  693.710000 2.635000 ;
      RECT  693.880000  0.255000  694.260000 0.715000 ;
      RECT  693.880000  1.665000  694.260000 2.465000 ;
      RECT  694.480000  0.085000  694.650000 0.545000 ;
      RECT  694.480000  1.835000  694.650000 2.635000 ;
      RECT  694.820000  0.255000  695.200000 0.715000 ;
      RECT  694.820000  1.665000  695.200000 2.465000 ;
      RECT  695.420000  0.085000  695.590000 0.545000 ;
      RECT  695.420000  1.835000  695.590000 2.635000 ;
      RECT  695.760000  0.255000  696.140000 0.715000 ;
      RECT  695.760000  1.665000  696.140000 2.465000 ;
      RECT  696.360000  0.085000  696.530000 0.545000 ;
      RECT  696.360000  1.835000  696.530000 2.635000 ;
      RECT  696.555000  0.905000  697.080000 1.495000 ;
      RECT  696.700000  0.255000  697.080000 0.715000 ;
      RECT  696.700000  1.665000  697.080000 2.465000 ;
      RECT  697.300000  0.085000  697.510000 0.885000 ;
      RECT  697.300000  1.835000  697.510000 2.635000 ;
      RECT  697.905000  0.085000  698.195000 0.810000 ;
      RECT  697.905000  1.470000  698.195000 2.635000 ;
      RECT  698.385000  1.075000  698.715000 1.325000 ;
      RECT  698.405000  0.085000  698.635000 0.905000 ;
      RECT  698.405000  1.495000  698.635000 2.635000 ;
      RECT  698.805000  0.255000  699.185000 0.885000 ;
      RECT  698.805000  1.485000  699.185000 2.465000 ;
      RECT  698.885000  0.885000  699.185000 1.485000 ;
      RECT  699.405000  0.085000  699.615000 0.905000 ;
      RECT  699.405000  1.495000  699.615000 2.635000 ;
      RECT  700.205000  0.085000  700.495000 0.810000 ;
      RECT  700.205000  1.470000  700.495000 2.635000 ;
      RECT  700.685000  1.075000  702.465000 1.325000 ;
      RECT  700.710000  0.085000  700.975000 0.545000 ;
      RECT  700.710000  1.495000  700.975000 2.635000 ;
      RECT  701.145000  0.255000  701.525000 0.725000 ;
      RECT  701.145000  0.725000  703.245000 0.905000 ;
      RECT  701.145000  1.495000  703.245000 1.665000 ;
      RECT  701.145000  1.665000  701.525000 2.465000 ;
      RECT  701.745000  0.085000  701.915000 0.545000 ;
      RECT  701.745000  1.835000  701.915000 2.635000 ;
      RECT  702.085000  0.255000  702.465000 0.725000 ;
      RECT  702.085000  1.665000  703.245000 1.685000 ;
      RECT  702.085000  1.685000  702.465000 2.465000 ;
      RECT  702.685000  0.085000  702.935000 0.550000 ;
      RECT  702.685000  2.175000  702.895000 2.635000 ;
      RECT  702.975000  0.905000  703.245000 1.495000 ;
      RECT  703.425000  0.085000  703.715000 0.810000 ;
      RECT  703.425000  1.470000  703.715000 2.635000 ;
      RECT  703.930000  0.085000  704.195000 0.545000 ;
      RECT  703.975000  1.495000  704.145000 2.635000 ;
      RECT  704.085000  1.075000  706.495000 1.325000 ;
      RECT  704.315000  1.495000  707.065000 1.665000 ;
      RECT  704.315000  1.665000  704.695000 2.465000 ;
      RECT  704.445000  0.255000  704.615000 0.725000 ;
      RECT  704.445000  0.725000  707.065000 0.905000 ;
      RECT  704.915000  0.085000  705.085000 0.545000 ;
      RECT  704.915000  1.835000  705.085000 2.635000 ;
      RECT  705.255000  1.665000  705.635000 2.465000 ;
      RECT  705.385000  0.255000  705.555000 0.725000 ;
      RECT  705.855000  0.085000  706.025000 0.545000 ;
      RECT  705.855000  1.835000  706.025000 2.635000 ;
      RECT  706.195000  1.665000  707.065000 1.685000 ;
      RECT  706.195000  1.685000  706.575000 2.465000 ;
      RECT  706.325000  0.255000  706.495000 0.725000 ;
      RECT  706.665000  0.085000  706.965000 0.550000 ;
      RECT  706.665000  0.905000  707.065000 1.495000 ;
      RECT  706.795000  2.175000  706.965000 2.635000 ;
      RECT  707.565000  0.085000  707.855000 0.810000 ;
      RECT  707.565000  1.470000  707.855000 2.635000 ;
      RECT  708.025000  0.715000  712.445000 0.905000 ;
      RECT  708.025000  0.905000  708.370000 1.495000 ;
      RECT  708.025000  1.495000  712.445000 1.665000 ;
      RECT  708.195000  0.085000  708.450000 0.545000 ;
      RECT  708.195000  1.835000  708.450000 2.635000 ;
      RECT  708.620000  0.255000  709.000000 0.715000 ;
      RECT  708.620000  1.075000  711.825000 1.325000 ;
      RECT  708.620000  1.665000  709.000000 2.465000 ;
      RECT  709.220000  0.085000  709.390000 0.545000 ;
      RECT  709.220000  1.835000  709.390000 2.635000 ;
      RECT  709.560000  0.255000  709.940000 0.715000 ;
      RECT  709.560000  1.665000  709.940000 2.465000 ;
      RECT  710.160000  0.085000  710.330000 0.545000 ;
      RECT  710.160000  1.835000  710.330000 2.635000 ;
      RECT  710.500000  0.255000  710.880000 0.715000 ;
      RECT  710.500000  1.665000  710.880000 2.465000 ;
      RECT  711.100000  0.085000  711.270000 0.545000 ;
      RECT  711.100000  1.835000  711.270000 2.635000 ;
      RECT  711.440000  0.255000  711.820000 0.715000 ;
      RECT  711.440000  1.665000  711.820000 2.465000 ;
      RECT  712.040000  0.085000  712.345000 0.545000 ;
      RECT  712.040000  1.835000  712.340000 2.635000 ;
      RECT  712.125000  0.905000  712.445000 1.495000 ;
      RECT  712.625000  0.085000  712.915000 0.810000 ;
      RECT  712.625000  1.470000  712.915000 2.635000 ;
      RECT  713.090000  0.255000  713.345000 1.495000 ;
      RECT  713.090000  1.495000  713.425000 2.465000 ;
      RECT  713.515000  0.085000  713.895000 0.485000 ;
      RECT  713.515000  0.655000  714.610000 0.825000 ;
      RECT  713.515000  0.825000  713.685000 1.325000 ;
      RECT  713.645000  1.495000  713.815000 2.635000 ;
      RECT  713.995000  0.995000  714.270000 1.325000 ;
      RECT  714.070000  1.325000  714.270000 2.295000 ;
      RECT  714.070000  2.295000  716.415000 2.465000 ;
      RECT  714.435000  0.255000  714.955000 0.620000 ;
      RECT  714.435000  0.620000  714.610000 0.655000 ;
      RECT  714.440000  0.825000  714.610000 1.955000 ;
      RECT  714.440000  1.955000  715.750000 2.125000 ;
      RECT  714.780000  0.815000  714.950000 1.615000 ;
      RECT  714.780000  1.615000  716.075000 1.785000 ;
      RECT  715.290000  0.255000  715.615000 1.415000 ;
      RECT  715.855000  0.255000  716.075000 1.615000 ;
      RECT  716.245000  1.440000  717.045000 1.630000 ;
      RECT  716.245000  1.630000  716.415000 2.295000 ;
      RECT  716.250000  0.085000  716.765000 0.620000 ;
      RECT  716.285000  0.895000  717.500000 1.065000 ;
      RECT  716.585000  1.875000  716.755000 2.635000 ;
      RECT  717.035000  0.290000  717.280000 0.895000 ;
      RECT  717.040000  1.875000  717.500000 2.285000 ;
      RECT  717.215000  1.065000  717.500000 1.875000 ;
      RECT  717.685000  0.085000  717.975000 0.810000 ;
      RECT  717.685000  1.470000  717.975000 2.635000 ;
      RECT  718.150000  0.085000  718.405000 0.885000 ;
      RECT  718.150000  1.495000  718.405000 2.635000 ;
      RECT  718.575000  0.255000  718.860000 1.595000 ;
      RECT  718.575000  1.595000  718.935000 2.465000 ;
      RECT  719.030000  0.995000  719.325000 1.325000 ;
      RECT  719.045000  0.085000  719.425000 0.465000 ;
      RECT  719.155000  0.635000  719.765000 0.805000 ;
      RECT  719.155000  0.805000  719.325000 0.995000 ;
      RECT  719.155000  1.325000  719.325000 1.835000 ;
      RECT  719.155000  1.835000  719.685000 2.005000 ;
      RECT  719.175000  2.175000  719.345000 2.635000 ;
      RECT  719.495000  0.995000  719.715000 1.495000 ;
      RECT  719.495000  1.495000  720.025000 1.665000 ;
      RECT  719.515000  2.005000  719.685000 2.255000 ;
      RECT  719.515000  2.255000  720.920000 2.425000 ;
      RECT  719.595000  0.265000  720.310000 0.595000 ;
      RECT  719.595000  0.595000  719.765000 0.635000 ;
      RECT  719.855000  1.665000  720.025000 1.835000 ;
      RECT  719.855000  1.835000  722.295000 2.005000 ;
      RECT  719.980000  0.765000  720.355000 1.280000 ;
      RECT  719.980000  1.280000  721.135000 1.325000 ;
      RECT  720.185000  1.325000  721.135000 1.410000 ;
      RECT  720.195000  1.410000  721.135000 1.625000 ;
      RECT  720.590000  0.775000  721.135000 1.105000 ;
      RECT  720.930000  0.420000  721.135000 0.775000 ;
      RECT  721.415000  0.755000  721.605000 1.625000 ;
      RECT  721.520000  2.175000  721.740000 2.635000 ;
      RECT  721.545000  0.085000  721.745000 0.585000 ;
      RECT  721.910000  2.005000  722.295000 2.465000 ;
      RECT  722.045000  0.255000  722.295000 1.835000 ;
      RECT  722.745000  0.085000  723.035000 0.810000 ;
      RECT  722.745000  1.470000  723.035000 2.635000 ;
      RECT  723.210000  0.295000  723.465000 0.625000 ;
      RECT  723.210000  0.625000  723.380000 1.495000 ;
      RECT  723.210000  1.495000  724.300000 1.665000 ;
      RECT  723.210000  1.665000  723.465000 2.465000 ;
      RECT  723.550000  0.995000  723.910000 1.325000 ;
      RECT  723.635000  0.085000  724.015000 0.465000 ;
      RECT  723.635000  1.835000  723.990000 2.635000 ;
      RECT  723.740000  0.635000  726.170000 0.805000 ;
      RECT  723.740000  0.805000  723.910000 0.995000 ;
      RECT  724.080000  0.995000  724.300000 1.495000 ;
      RECT  724.160000  1.935000  724.560000 2.275000 ;
      RECT  724.160000  2.275000  726.090000 2.445000 ;
      RECT  724.570000  0.995000  724.915000 1.615000 ;
      RECT  724.750000  1.935000  726.565000 2.105000 ;
      RECT  725.085000  0.995000  725.705000 1.325000 ;
      RECT  725.195000  0.295000  726.550000 0.465000 ;
      RECT  725.250000  1.595000  727.105000 1.765000 ;
      RECT  726.000000  0.805000  726.170000 0.995000 ;
      RECT  726.000000  0.995000  726.715000 1.325000 ;
      RECT  726.380000  0.465000  726.550000 0.655000 ;
      RECT  726.380000  0.655000  727.105000 0.825000 ;
      RECT  726.395000  2.105000  726.565000 2.465000 ;
      RECT  726.735000  0.085000  727.115000 0.465000 ;
      RECT  726.735000  2.255000  727.115000 2.635000 ;
      RECT  726.935000  0.825000  727.105000 1.075000 ;
      RECT  726.935000  1.075000  728.550000 1.245000 ;
      RECT  726.935000  1.245000  727.105000 1.595000 ;
      RECT  727.335000  0.255000  727.505000 0.635000 ;
      RECT  727.335000  0.635000  729.000000 0.805000 ;
      RECT  727.335000  1.575000  729.000000 1.745000 ;
      RECT  727.335000  1.745000  727.505000 2.465000 ;
      RECT  727.675000  0.085000  728.055000 0.465000 ;
      RECT  727.675000  1.915000  728.055000 2.635000 ;
      RECT  728.275000  0.255000  728.445000 0.635000 ;
      RECT  728.275000  1.745000  728.445000 2.465000 ;
      RECT  728.615000  0.085000  728.995000 0.465000 ;
      RECT  728.615000  1.915000  728.995000 2.635000 ;
      RECT  728.770000  0.805000  729.000000 1.575000 ;
      RECT  729.185000  0.085000  729.475000 0.810000 ;
      RECT  729.185000  1.470000  729.475000 2.635000 ;
      RECT  729.650000  0.085000  729.985000 0.465000 ;
      RECT  729.650000  1.915000  729.985000 2.635000 ;
      RECT  730.165000  0.255000  730.375000 0.635000 ;
      RECT  730.165000  0.635000  733.195000 0.805000 ;
      RECT  730.165000  0.805000  730.425000 1.575000 ;
      RECT  730.165000  1.575000  733.195000 1.745000 ;
      RECT  730.165000  1.745000  730.375000 2.465000 ;
      RECT  730.545000  0.085000  730.925000 0.465000 ;
      RECT  730.545000  1.915000  730.925000 2.635000 ;
      RECT  730.645000  1.075000  733.535000 1.245000 ;
      RECT  731.145000  0.295000  731.315000 0.635000 ;
      RECT  731.145000  1.745000  731.315000 2.465000 ;
      RECT  731.485000  0.085000  731.865000 0.465000 ;
      RECT  731.485000  1.915000  731.865000 2.635000 ;
      RECT  732.085000  0.255000  732.255000 0.635000 ;
      RECT  732.085000  1.745000  732.255000 2.465000 ;
      RECT  732.425000  0.085000  732.805000 0.465000 ;
      RECT  732.425000  1.915000  732.805000 2.635000 ;
      RECT  733.025000  0.295000  733.195000 0.635000 ;
      RECT  733.025000  1.745000  733.195000 2.465000 ;
      RECT  733.365000  0.085000  733.745000 0.465000 ;
      RECT  733.365000  0.635000  734.900000 0.805000 ;
      RECT  733.365000  0.805000  733.535000 1.075000 ;
      RECT  733.365000  1.245000  733.535000 1.835000 ;
      RECT  733.365000  1.835000  738.535000 2.005000 ;
      RECT  733.365000  2.255000  733.745000 2.635000 ;
      RECT  733.705000  0.995000  733.925000 1.495000 ;
      RECT  733.705000  1.495000  736.145000 1.665000 ;
      RECT  733.915000  0.295000  735.085000 0.465000 ;
      RECT  734.190000  2.255000  735.965000 2.425000 ;
      RECT  734.250000  1.105000  734.485000 1.275000 ;
      RECT  734.265000  0.995000  734.485000 1.105000 ;
      RECT  734.265000  1.275000  734.485000 1.325000 ;
      RECT  734.730000  0.805000  734.900000 0.935000 ;
      RECT  735.140000  0.645000  737.055000 0.815000 ;
      RECT  735.140000  0.815000  735.360000 1.325000 ;
      RECT  735.315000  0.425000  735.950000 0.645000 ;
      RECT  735.730000  0.995000  736.145000 1.495000 ;
      RECT  736.220000  0.085000  736.550000 0.465000 ;
      RECT  736.235000  2.175000  736.405000 2.635000 ;
      RECT  736.455000  0.995000  736.675000 1.495000 ;
      RECT  736.455000  1.495000  739.195000 1.665000 ;
      RECT  736.590000  2.255000  739.005000 2.425000 ;
      RECT  736.735000  0.295000  738.125000 0.465000 ;
      RECT  736.885000  0.815000  737.055000 0.995000 ;
      RECT  736.885000  0.995000  737.405000 1.165000 ;
      RECT  737.185000  1.165000  737.405000 1.325000 ;
      RECT  737.275000  0.635000  737.930000 0.805000 ;
      RECT  737.710000  0.805000  737.930000 0.935000 ;
      RECT  738.445000  0.995000  738.730000 1.325000 ;
      RECT  738.975000  0.645000  739.945000 0.815000 ;
      RECT  738.975000  0.815000  739.195000 1.495000 ;
      RECT  738.975000  1.665000  739.195000 1.915000 ;
      RECT  738.975000  1.915000  739.945000 2.085000 ;
      RECT  739.225000  0.085000  739.605000 0.465000 ;
      RECT  739.225000  2.255000  739.605000 2.635000 ;
      RECT  739.365000  0.995000  739.795000 1.615000 ;
      RECT  739.775000  0.295000  739.945000 0.645000 ;
      RECT  739.775000  1.795000  739.945000 1.915000 ;
      RECT  739.775000  2.085000  739.945000 2.465000 ;
      RECT  740.225000  0.085000  740.515000 0.810000 ;
      RECT  740.225000  1.470000  740.515000 2.635000 ;
      RECT  740.685000  0.255000  742.455000 0.425000 ;
      RECT  740.685000  0.425000  741.040000 0.465000 ;
      RECT  740.685000  0.465000  740.945000 0.885000 ;
      RECT  740.685000  1.060000  741.020000 1.285000 ;
      RECT  740.720000  1.455000  741.020000 2.295000 ;
      RECT  740.720000  2.295000  742.325000 2.465000 ;
      RECT  741.205000  0.595000  741.435000 1.455000 ;
      RECT  741.205000  1.455000  741.490000 2.125000 ;
      RECT  741.605000  0.655000  742.350000 0.715000 ;
      RECT  741.605000  0.715000  743.300000 0.825000 ;
      RECT  741.605000  0.995000  741.865000 1.325000 ;
      RECT  741.665000  0.425000  742.455000 0.465000 ;
      RECT  741.665000  1.325000  741.865000 2.110000 ;
      RECT  742.085000  1.075000  743.795000 1.310000 ;
      RECT  742.105000  1.480000  743.345000 1.650000 ;
      RECT  742.105000  1.650000  742.325000 2.295000 ;
      RECT  742.175000  0.825000  743.300000 0.885000 ;
      RECT  742.495000  1.835000  742.775000 2.635000 ;
      RECT  742.625000  0.085000  742.795000 0.525000 ;
      RECT  742.965000  1.650000  743.345000 2.465000 ;
      RECT  743.065000  0.255000  743.300000 0.715000 ;
      RECT  743.530000  0.255000  743.795000 1.075000 ;
      RECT  743.570000  1.310000  743.795000 2.465000 ;
      RECT  743.965000  0.760000  744.350000 1.620000 ;
      RECT  744.075000  1.835000  744.370000 2.635000 ;
      RECT  744.115000  0.085000  744.335000 0.545000 ;
      RECT  744.825000  0.085000  745.115000 0.810000 ;
      RECT  744.825000  1.470000  745.115000 2.635000 ;
      RECT  745.285000  0.345000  745.545000 0.675000 ;
      RECT  745.285000  0.675000  745.460000 1.495000 ;
      RECT  745.285000  1.495000  746.745000 1.665000 ;
      RECT  745.285000  1.665000  745.460000 2.135000 ;
      RECT  745.285000  2.135000  745.545000 2.465000 ;
      RECT  745.630000  0.995000  746.030000 1.325000 ;
      RECT  745.715000  0.085000  746.085000 0.545000 ;
      RECT  745.715000  2.255000  746.095000 2.635000 ;
      RECT  745.830000  0.725000  746.030000 0.995000 ;
      RECT  746.185000  1.835000  747.085000 2.005000 ;
      RECT  746.315000  0.575000  746.555000 0.935000 ;
      RECT  746.525000  1.155000  747.385000 1.325000 ;
      RECT  746.525000  1.325000  746.745000 1.495000 ;
      RECT  746.655000  2.255000  747.035000 2.635000 ;
      RECT  746.785000  0.085000  747.035000 0.885000 ;
      RECT  746.915000  1.495000  748.965000 1.665000 ;
      RECT  746.915000  1.665000  747.085000 1.835000 ;
      RECT  747.005000  1.075000  747.385000 1.155000 ;
      RECT  747.255000  0.295000  747.425000 0.735000 ;
      RECT  747.255000  0.735000  748.965000 0.905000 ;
      RECT  747.255000  2.135000  747.480000 2.465000 ;
      RECT  747.310000  1.835000  748.335000 1.915000 ;
      RECT  747.310000  1.915000  749.950000 2.005000 ;
      RECT  747.310000  2.005000  747.480000 2.135000 ;
      RECT  747.725000  0.085000  747.895000 0.545000 ;
      RECT  747.725000  2.175000  747.975000 2.635000 ;
      RECT  747.920000  1.075000  749.225000 1.275000 ;
      RECT  748.165000  0.295000  750.625000 0.465000 ;
      RECT  748.165000  2.005000  749.950000 2.085000 ;
      RECT  748.165000  2.255000  750.625000 2.425000 ;
      RECT  748.585000  0.655000  748.965000 0.735000 ;
      RECT  748.585000  1.665000  748.965000 1.715000 ;
      RECT  749.400000  0.655000  749.945000 0.825000 ;
      RECT  749.400000  0.825000  749.705000 0.935000 ;
      RECT  749.910000  0.995000  750.285000 1.615000 ;
      RECT  750.400000  1.785000  750.625000 2.255000 ;
      RECT  750.455000  0.465000  750.625000 1.785000 ;
      RECT  750.805000  0.085000  751.095000 0.810000 ;
      RECT  750.805000  1.470000  751.095000 2.635000 ;
      RECT  751.275000  0.315000  755.365000 0.485000 ;
      RECT  751.275000  0.485000  751.500000 2.255000 ;
      RECT  751.275000  2.255000  755.365000 2.425000 ;
      RECT  751.695000  0.655000  753.030000 0.825000 ;
      RECT  751.695000  1.575000  757.310000 1.745000 ;
      RECT  751.770000  0.995000  752.415000 1.325000 ;
      RECT  752.635000  0.825000  753.030000 0.935000 ;
      RECT  753.535000  0.995000  755.230000 1.325000 ;
      RECT  753.575000  0.655000  757.215000 0.825000 ;
      RECT  753.575000  1.915000  759.095000 2.085000 ;
      RECT  755.425000  1.075000  757.710000 1.290000 ;
      RECT  755.555000  0.085000  755.885000 0.465000 ;
      RECT  755.555000  2.255000  755.885000 2.635000 ;
      RECT  756.105000  0.255000  756.275000 0.655000 ;
      RECT  756.445000  0.085000  756.825000 0.465000 ;
      RECT  756.445000  2.255000  756.825000 2.635000 ;
      RECT  757.045000  0.255000  757.215000 0.655000 ;
      RECT  757.385000  0.085000  757.760000 0.590000 ;
      RECT  757.385000  2.255000  757.765000 2.635000 ;
      RECT  757.540000  1.290000  757.710000 1.425000 ;
      RECT  757.540000  1.425000  759.830000 1.595000 ;
      RECT  757.980000  0.255000  758.155000 0.715000 ;
      RECT  757.980000  0.715000  759.095000 0.905000 ;
      RECT  757.980000  0.905000  758.280000 0.935000 ;
      RECT  757.985000  1.795000  758.155000 1.915000 ;
      RECT  757.985000  2.085000  758.155000 2.465000 ;
      RECT  758.325000  2.255000  758.705000 2.635000 ;
      RECT  758.425000  0.085000  758.675000 0.545000 ;
      RECT  758.610000  1.075000  759.490000 1.245000 ;
      RECT  758.925000  0.510000  759.095000 0.715000 ;
      RECT  758.925000  1.795000  759.095000 1.915000 ;
      RECT  758.925000  2.085000  759.095000 2.465000 ;
      RECT  759.270000  0.655000  760.225000 0.825000 ;
      RECT  759.270000  0.825000  759.490000 1.075000 ;
      RECT  759.415000  0.085000  759.745000 0.465000 ;
      RECT  759.415000  2.255000  759.745000 2.635000 ;
      RECT  759.660000  0.995000  759.830000 1.425000 ;
      RECT  759.965000  0.255000  760.225000 0.655000 ;
      RECT  759.965000  1.795000  760.225000 2.465000 ;
      RECT  760.050000  0.825000  760.225000 1.795000 ;
      RECT  760.465000  0.085000  760.755000 0.810000 ;
      RECT  760.465000  1.470000  760.755000 2.635000 ;
      RECT  760.925000  0.085000  761.235000 0.885000 ;
      RECT  760.925000  1.495000  761.205000 2.635000 ;
      RECT  760.935000  1.055000  761.270000 1.325000 ;
      RECT  761.375000  1.485000  761.755000 2.465000 ;
      RECT  761.490000  0.255000  762.235000 0.885000 ;
      RECT  761.490000  0.885000  761.660000 1.485000 ;
      RECT  761.830000  1.075000  762.215000 1.325000 ;
      RECT  761.975000  1.495000  762.235000 2.635000 ;
      RECT  762.765000  0.085000  763.055000 0.810000 ;
      RECT  762.765000  1.470000  763.055000 2.635000 ;
      RECT  763.225000  0.255000  763.565000 0.715000 ;
      RECT  763.225000  0.715000  764.425000 0.885000 ;
      RECT  763.225000  1.075000  764.035000 1.325000 ;
      RECT  763.225000  1.495000  763.485000 2.635000 ;
      RECT  763.655000  1.495000  765.370000 1.665000 ;
      RECT  763.655000  1.665000  764.035000 2.465000 ;
      RECT  763.785000  0.085000  763.955000 0.545000 ;
      RECT  764.125000  0.255000  765.445000 0.485000 ;
      RECT  764.125000  0.485000  764.425000 0.715000 ;
      RECT  764.205000  1.075000  764.920000 1.325000 ;
      RECT  764.255000  1.835000  764.425000 2.635000 ;
      RECT  764.595000  0.655000  765.370000 0.905000 ;
      RECT  764.595000  1.665000  764.975000 2.465000 ;
      RECT  765.090000  0.905000  765.370000 1.495000 ;
      RECT  765.195000  1.835000  765.450000 2.635000 ;
      RECT  765.985000  0.085000  766.275000 0.810000 ;
      RECT  765.985000  1.470000  766.275000 2.635000 ;
      RECT  766.450000  0.255000  766.785000 0.715000 ;
      RECT  766.450000  0.715000  768.585000 0.905000 ;
      RECT  766.450000  1.495000  766.705000 2.635000 ;
      RECT  766.470000  1.075000  768.240000 1.325000 ;
      RECT  766.875000  1.495000  770.075000 1.665000 ;
      RECT  766.875000  1.665000  767.255000 2.465000 ;
      RECT  767.005000  0.085000  767.175000 0.545000 ;
      RECT  767.345000  0.255000  767.725000 0.715000 ;
      RECT  767.475000  1.835000  767.645000 2.635000 ;
      RECT  767.815000  1.665000  768.195000 2.465000 ;
      RECT  767.945000  0.085000  768.115000 0.545000 ;
      RECT  768.285000  0.255000  770.545000 0.465000 ;
      RECT  768.285000  0.465000  768.585000 0.715000 ;
      RECT  768.415000  1.835000  768.585000 2.635000 ;
      RECT  768.755000  0.635000  770.075000 0.805000 ;
      RECT  768.755000  0.805000  769.055000 1.495000 ;
      RECT  768.755000  1.665000  769.135000 2.465000 ;
      RECT  769.225000  1.075000  770.475000 1.325000 ;
      RECT  769.355000  1.835000  769.525000 2.635000 ;
      RECT  769.695000  1.665000  770.075000 2.465000 ;
      RECT  770.295000  0.465000  770.545000 0.885000 ;
      RECT  770.295000  1.835000  770.545000 2.635000 ;
      RECT  771.045000  0.085000  771.335000 0.810000 ;
      RECT  771.045000  1.470000  771.335000 2.635000 ;
      RECT  771.510000  0.255000  771.845000 0.735000 ;
      RECT  771.510000  0.735000  775.525000 0.905000 ;
      RECT  771.510000  1.495000  771.765000 2.635000 ;
      RECT  771.930000  1.075000  775.135000 1.295000 ;
      RECT  771.935000  1.465000  778.895000 1.665000 ;
      RECT  771.935000  1.665000  772.315000 2.465000 ;
      RECT  772.065000  0.085000  772.235000 0.565000 ;
      RECT  772.405000  0.255000  772.785000 0.735000 ;
      RECT  772.535000  1.835000  772.705000 2.635000 ;
      RECT  772.875000  1.665000  773.255000 2.465000 ;
      RECT  773.005000  0.085000  773.175000 0.565000 ;
      RECT  773.345000  0.255000  773.725000 0.735000 ;
      RECT  773.475000  1.835000  773.645000 2.635000 ;
      RECT  773.815000  1.665000  774.195000 2.465000 ;
      RECT  773.945000  0.085000  774.115000 0.565000 ;
      RECT  774.285000  0.255000  774.665000 0.735000 ;
      RECT  774.415000  1.835000  774.585000 2.635000 ;
      RECT  774.755000  1.665000  775.135000 2.465000 ;
      RECT  774.885000  0.085000  775.055000 0.565000 ;
      RECT  775.225000  0.255000  779.490000 0.485000 ;
      RECT  775.225000  0.485000  775.525000 0.735000 ;
      RECT  775.355000  1.835000  775.525000 2.635000 ;
      RECT  775.460000  1.075000  775.990000 1.465000 ;
      RECT  775.695000  0.655000  778.895000 0.905000 ;
      RECT  775.695000  0.905000  775.990000 1.075000 ;
      RECT  775.695000  1.665000  776.075000 2.465000 ;
      RECT  776.160000  1.075000  778.425000 1.275000 ;
      RECT  776.295000  1.835000  776.465000 2.635000 ;
      RECT  776.635000  1.665000  777.015000 2.465000 ;
      RECT  777.235000  1.835000  777.405000 2.635000 ;
      RECT  777.575000  1.665000  777.955000 2.465000 ;
      RECT  778.175000  1.835000  778.345000 2.635000 ;
      RECT  778.515000  1.665000  778.895000 2.465000 ;
      RECT  778.645000  0.905000  778.895000 1.465000 ;
      RECT  779.115000  0.485000  779.490000 0.905000 ;
      RECT  779.135000  1.495000  779.490000 2.635000 ;
      RECT  779.785000  0.085000  780.075000 0.810000 ;
      RECT  779.785000  1.470000  780.075000 2.635000 ;
      RECT  780.250000  0.525000  780.520000 0.735000 ;
      RECT  780.250000  0.735000  781.780000 0.905000 ;
      RECT  780.250000  1.075000  780.580000 1.315000 ;
      RECT  780.250000  1.495000  781.780000 1.665000 ;
      RECT  780.250000  1.665000  780.530000 1.825000 ;
      RECT  780.750000  1.075000  781.345000 1.315000 ;
      RECT  780.790000  0.085000  781.120000 0.545000 ;
      RECT  780.790000  1.835000  781.040000 2.635000 ;
      RECT  781.210000  1.835000  782.350000 2.005000 ;
      RECT  781.210000  2.005000  781.590000 2.465000 ;
      RECT  781.520000  0.255000  782.350000 0.545000 ;
      RECT  781.610000  0.905000  781.780000 1.495000 ;
      RECT  781.810000  2.175000  782.025000 2.635000 ;
      RECT  781.980000  0.545000  782.350000 1.835000 ;
      RECT  782.545000  0.085000  782.835000 0.810000 ;
      RECT  782.545000  1.470000  782.835000 2.635000 ;
      RECT  783.030000  0.510000  783.265000 0.840000 ;
      RECT  783.030000  0.840000  783.200000 1.495000 ;
      RECT  783.030000  1.495000  784.110000 1.665000 ;
      RECT  783.030000  1.665000  783.330000 1.860000 ;
      RECT  783.375000  0.995000  783.770000 1.325000 ;
      RECT  783.515000  0.085000  783.685000 0.775000 ;
      RECT  783.550000  1.835000  783.805000 2.635000 ;
      RECT  783.940000  0.995000  784.110000 1.495000 ;
      RECT  783.955000  0.255000  785.125000 0.465000 ;
      RECT  784.055000  1.835000  785.535000 2.005000 ;
      RECT  784.055000  2.005000  784.385000 2.465000 ;
      RECT  784.375000  0.635000  784.705000 1.835000 ;
      RECT  784.645000  2.175000  785.020000 2.635000 ;
      RECT  784.875000  0.465000  785.125000 0.695000 ;
      RECT  784.875000  0.695000  786.015000 0.905000 ;
      RECT  785.030000  1.075000  786.015000 1.275000 ;
      RECT  785.205000  2.005000  785.535000 2.465000 ;
      RECT  785.260000  1.495000  785.535000 1.835000 ;
      RECT  785.345000  0.085000  785.515000 0.525000 ;
      RECT  785.685000  0.255000  786.015000 0.695000 ;
      RECT  785.765000  1.835000  785.935000 2.635000 ;
      RECT  785.825000  1.275000  786.015000 1.655000 ;
      RECT  786.225000  0.085000  786.515000 0.810000 ;
      RECT  786.225000  1.470000  786.515000 2.635000 ;
      RECT  786.690000  0.255000  787.025000 0.715000 ;
      RECT  786.690000  0.715000  787.430000 0.905000 ;
      RECT  786.690000  1.445000  787.430000 1.665000 ;
      RECT  786.690000  1.665000  787.025000 2.465000 ;
      RECT  786.710000  1.075000  787.040000 1.275000 ;
      RECT  787.245000  0.085000  787.440000 0.545000 ;
      RECT  787.245000  1.835000  787.935000 2.635000 ;
      RECT  787.260000  0.905000  787.430000 1.075000 ;
      RECT  787.260000  1.075000  788.955000 1.275000 ;
      RECT  787.260000  1.275000  787.430000 1.445000 ;
      RECT  787.620000  1.445000  787.935000 1.835000 ;
      RECT  787.685000  0.255000  789.910000 0.465000 ;
      RECT  787.685000  0.465000  787.935000 0.905000 ;
      RECT  788.105000  0.635000  789.440000 0.905000 ;
      RECT  788.105000  1.445000  791.320000 1.665000 ;
      RECT  788.105000  1.665000  788.485000 2.465000 ;
      RECT  788.705000  1.835000  788.875000 2.635000 ;
      RECT  789.045000  1.665000  789.440000 2.465000 ;
      RECT  789.175000  0.905000  789.440000 1.445000 ;
      RECT  789.660000  0.465000  789.910000 0.715000 ;
      RECT  789.660000  0.715000  791.900000 0.905000 ;
      RECT  789.660000  1.835000  789.830000 2.635000 ;
      RECT  790.000000  1.665000  790.380000 2.465000 ;
      RECT  790.005000  1.075000  791.990000 1.275000 ;
      RECT  790.130000  0.085000  790.300000 0.545000 ;
      RECT  790.470000  0.255000  790.850000 0.715000 ;
      RECT  790.600000  1.835000  790.770000 2.635000 ;
      RECT  790.940000  1.665000  791.320000 2.465000 ;
      RECT  791.070000  0.085000  791.310000 0.545000 ;
      RECT  791.570000  0.255000  791.900000 0.715000 ;
      RECT  791.570000  1.495000  791.900000 2.635000 ;
      RECT  792.205000  0.085000  792.495000 0.810000 ;
      RECT  792.205000  1.470000  792.495000 2.635000 ;
      RECT  792.670000  0.085000  792.925000 0.575000 ;
      RECT  792.670000  1.495000  792.925000 2.635000 ;
      RECT  792.690000  0.745000  792.910000 1.325000 ;
      RECT  793.095000  0.255000  794.475000 0.595000 ;
      RECT  793.095000  0.595000  793.325000 1.495000 ;
      RECT  793.095000  1.495000  794.475000 1.665000 ;
      RECT  793.095000  1.665000  793.475000 2.465000 ;
      RECT  793.495000  0.765000  793.865000 1.325000 ;
      RECT  793.695000  1.835000  793.925000 2.635000 ;
      RECT  794.055000  0.995000  794.485000 1.325000 ;
      RECT  794.095000  0.595000  794.475000 0.825000 ;
      RECT  794.095000  1.665000  794.475000 2.465000 ;
      RECT  794.965000  0.085000  795.255000 0.810000 ;
      RECT  794.965000  1.470000  795.255000 2.635000 ;
      RECT  795.430000  0.295000  797.645000 0.465000 ;
      RECT  795.430000  0.465000  795.685000 0.785000 ;
      RECT  795.430000  0.995000  795.670000 1.325000 ;
      RECT  795.430000  1.495000  795.685000 2.635000 ;
      RECT  795.855000  0.635000  796.235000 1.445000 ;
      RECT  795.855000  1.445000  798.635000 1.665000 ;
      RECT  795.855000  1.665000  796.235000 2.465000 ;
      RECT  796.455000  1.835000  796.625000 2.635000 ;
      RECT  796.510000  1.075000  797.955000 1.275000 ;
      RECT  796.795000  0.635000  798.635000 0.905000 ;
      RECT  796.795000  1.665000  797.175000 2.465000 ;
      RECT  797.395000  1.835000  798.085000 2.635000 ;
      RECT  797.835000  0.085000  798.165000 0.465000 ;
      RECT  798.125000  1.075000  799.340000 1.275000 ;
      RECT  798.255000  1.665000  798.635000 2.465000 ;
      RECT  798.855000  0.085000  799.235000 0.885000 ;
      RECT  798.855000  1.445000  799.235000 2.635000 ;
      RECT  799.565000  0.085000  799.855000 0.810000 ;
      RECT  799.565000  1.470000  799.855000 2.635000 ;
      RECT  800.030000  0.255000  800.365000 0.735000 ;
      RECT  800.030000  0.735000  804.125000 0.905000 ;
      RECT  800.030000  1.445000  800.285000 2.635000 ;
      RECT  800.050000  1.075000  801.790000 1.275000 ;
      RECT  800.455000  1.445000  806.725000 1.665000 ;
      RECT  800.455000  1.665000  800.835000 2.465000 ;
      RECT  800.585000  0.085000  800.755000 0.565000 ;
      RECT  800.925000  0.255000  801.305000 0.735000 ;
      RECT  801.055000  1.835000  801.225000 2.635000 ;
      RECT  801.395000  1.665000  801.775000 2.465000 ;
      RECT  801.525000  0.085000  801.695000 0.565000 ;
      RECT  801.865000  0.655000  802.245000 0.735000 ;
      RECT  801.995000  1.835000  802.165000 2.635000 ;
      RECT  802.215000  1.075000  803.965000 1.275000 ;
      RECT  802.335000  0.255000  806.540000 0.485000 ;
      RECT  802.335000  1.665000  802.715000 2.465000 ;
      RECT  802.805000  0.655000  803.185000 0.735000 ;
      RECT  802.935000  1.835000  803.105000 2.635000 ;
      RECT  803.275000  1.665000  803.655000 2.465000 ;
      RECT  803.745000  0.655000  804.125000 0.735000 ;
      RECT  803.875000  1.835000  804.565000 2.635000 ;
      RECT  804.190000  1.075000  806.310000 1.275000 ;
      RECT  804.735000  0.655000  806.725000 0.905000 ;
      RECT  804.735000  1.665000  805.115000 2.465000 ;
      RECT  805.335000  1.835000  805.505000 2.635000 ;
      RECT  805.675000  1.665000  806.055000 2.465000 ;
      RECT  806.275000  1.835000  806.540000 2.635000 ;
      RECT  806.495000  0.905000  806.725000 1.445000 ;
      RECT  806.925000  0.085000  807.215000 0.810000 ;
      RECT  806.925000  1.470000  807.215000 2.635000 ;
      RECT  807.385000  0.445000  807.810000 0.655000 ;
      RECT  807.385000  0.655000  809.520000 0.825000 ;
      RECT  807.385000  0.825000  807.555000 1.595000 ;
      RECT  807.385000  1.595000  807.810000 1.925000 ;
      RECT  807.725000  0.995000  808.125000 1.325000 ;
      RECT  808.060000  0.085000  808.390000 0.485000 ;
      RECT  808.060000  1.495000  808.310000 2.635000 ;
      RECT  808.315000  0.995000  808.635000 1.325000 ;
      RECT  808.480000  1.495000  809.975000 1.665000 ;
      RECT  808.480000  1.665000  808.860000 2.465000 ;
      RECT  808.820000  0.995000  809.095000 1.325000 ;
      RECT  809.090000  1.835000  809.260000 2.635000 ;
      RECT  809.300000  0.825000  809.520000 1.325000 ;
      RECT  809.430000  0.255000  809.975000 0.485000 ;
      RECT  809.430000  1.665000  809.975000 2.465000 ;
      RECT  809.710000  0.485000  809.975000 1.495000 ;
      RECT  810.145000  0.085000  810.435000 0.810000 ;
      RECT  810.145000  1.470000  810.435000 2.635000 ;
      RECT  810.610000  0.255000  810.930000 0.655000 ;
      RECT  810.610000  0.655000  810.780000 1.445000 ;
      RECT  810.610000  1.445000  814.520000 1.615000 ;
      RECT  810.610000  1.615000  810.780000 2.065000 ;
      RECT  810.610000  2.065000  810.930000 2.465000 ;
      RECT  810.950000  1.075000  811.350000 1.275000 ;
      RECT  811.150000  0.085000  811.460000 0.905000 ;
      RECT  811.150000  1.835000  811.460000 2.635000 ;
      RECT  811.585000  1.075000  812.410000 1.275000 ;
      RECT  811.630000  0.255000  812.010000 0.715000 ;
      RECT  811.630000  0.715000  813.520000 0.905000 ;
      RECT  811.630000  1.785000  815.010000 1.955000 ;
      RECT  811.630000  1.955000  812.950000 2.005000 ;
      RECT  811.630000  2.005000  812.010000 2.465000 ;
      RECT  812.230000  0.085000  812.480000 0.545000 ;
      RECT  812.230000  2.175000  812.400000 2.635000 ;
      RECT  812.570000  2.005000  812.950000 2.465000 ;
      RECT  812.670000  1.075000  813.960000 1.275000 ;
      RECT  812.720000  0.255000  814.970000 0.465000 ;
      RECT  812.720000  0.635000  813.520000 0.715000 ;
      RECT  813.170000  2.175000  813.420000 2.635000 ;
      RECT  813.610000  2.175000  813.910000 2.635000 ;
      RECT  813.740000  0.465000  813.910000 0.905000 ;
      RECT  814.080000  0.635000  815.010000 0.905000 ;
      RECT  814.080000  1.955000  815.010000 2.005000 ;
      RECT  814.080000  2.005000  814.380000 2.465000 ;
      RECT  814.190000  1.075000  814.520000 1.445000 ;
      RECT  814.680000  2.175000  814.970000 2.635000 ;
      RECT  814.770000  0.905000  815.010000 1.785000 ;
      RECT  815.205000  0.085000  815.495000 0.810000 ;
      RECT  815.205000  1.470000  815.495000 2.635000 ;
      RECT  815.665000  0.255000  816.005000 0.715000 ;
      RECT  815.665000  0.715000  816.915000 0.905000 ;
      RECT  815.665000  0.905000  815.840000 1.445000 ;
      RECT  815.665000  1.445000  816.005000 2.465000 ;
      RECT  816.010000  1.075000  816.410000 1.275000 ;
      RECT  816.225000  0.085000  816.475000 0.545000 ;
      RECT  816.225000  1.445000  816.915000 2.635000 ;
      RECT  816.635000  0.905000  816.915000 1.075000 ;
      RECT  816.635000  1.075000  818.405000 1.275000 ;
      RECT  816.665000  0.255000  820.755000 0.465000 ;
      RECT  817.085000  0.635000  818.795000 0.905000 ;
      RECT  817.085000  1.445000  822.685000 1.665000 ;
      RECT  817.085000  1.665000  817.465000 2.465000 ;
      RECT  817.685000  1.835000  817.855000 2.635000 ;
      RECT  818.025000  1.665000  819.345000 2.005000 ;
      RECT  818.025000  2.005000  818.405000 2.465000 ;
      RECT  818.625000  0.905000  818.795000 1.075000 ;
      RECT  818.625000  1.075000  819.135000 1.445000 ;
      RECT  818.625000  2.175000  818.795000 2.635000 ;
      RECT  818.965000  0.635000  820.755000 0.715000 ;
      RECT  818.965000  0.715000  822.685000 0.905000 ;
      RECT  818.965000  2.005000  819.345000 2.465000 ;
      RECT  819.305000  1.075000  820.510000 1.275000 ;
      RECT  819.565000  1.835000  819.735000 2.635000 ;
      RECT  819.905000  1.665000  820.285000 2.465000 ;
      RECT  820.505000  1.835000  821.195000 2.635000 ;
      RECT  820.765000  1.075000  822.680000 1.275000 ;
      RECT  820.945000  0.085000  821.195000 0.545000 ;
      RECT  821.365000  0.255000  821.745000 0.715000 ;
      RECT  821.365000  1.665000  821.745000 2.465000 ;
      RECT  821.965000  0.085000  822.135000 0.545000 ;
      RECT  821.965000  1.835000  822.135000 2.635000 ;
      RECT  822.305000  0.255000  822.685000 0.715000 ;
      RECT  822.305000  1.665000  822.685000 2.465000 ;
      RECT  822.905000  0.085000  823.235000 0.905000 ;
      RECT  822.905000  1.445000  823.235000 2.635000 ;
      RECT  823.485000  0.085000  823.775000 0.810000 ;
      RECT  823.485000  1.470000  823.775000 2.635000 ;
      RECT  823.945000  1.495000  824.205000 2.635000 ;
      RECT  823.950000  0.085000  824.285000 0.825000 ;
      RECT  823.970000  0.995000  824.255000 1.325000 ;
      RECT  824.375000  1.495000  825.805000 1.665000 ;
      RECT  824.375000  1.665000  824.755000 2.465000 ;
      RECT  824.455000  0.300000  824.720000 0.995000 ;
      RECT  824.455000  0.995000  824.935000 1.325000 ;
      RECT  824.890000  0.300000  825.275000 0.825000 ;
      RECT  824.975000  1.835000  825.145000 2.635000 ;
      RECT  825.105000  0.825000  825.275000 0.995000 ;
      RECT  825.105000  0.995000  825.465000 1.325000 ;
      RECT  825.395000  1.665000  825.725000 2.465000 ;
      RECT  825.530000  0.255000  826.275000 0.825000 ;
      RECT  825.635000  0.825000  825.805000 1.495000 ;
      RECT  825.975000  1.835000  826.255000 2.635000 ;
      RECT  826.035000  0.995000  826.500000 1.665000 ;
      RECT  826.705000  0.085000  826.995000 0.810000 ;
      RECT  826.705000  1.470000  826.995000 2.635000 ;
      RECT  827.170000  0.255000  827.505000 0.735000 ;
      RECT  827.170000  0.735000  828.365000 0.905000 ;
      RECT  827.170000  1.495000  827.425000 2.635000 ;
      RECT  827.190000  1.075000  827.975000 1.275000 ;
      RECT  827.595000  1.445000  831.405000 1.665000 ;
      RECT  827.595000  1.665000  827.975000 2.465000 ;
      RECT  827.725000  0.085000  827.895000 0.545000 ;
      RECT  828.065000  0.255000  829.405000 0.465000 ;
      RECT  828.065000  0.465000  828.365000 0.735000 ;
      RECT  828.145000  1.075000  828.930000 1.275000 ;
      RECT  828.195000  1.835000  828.365000 2.635000 ;
      RECT  828.535000  0.635000  830.465000 0.905000 ;
      RECT  828.535000  1.665000  828.915000 2.465000 ;
      RECT  829.135000  1.835000  829.465000 2.635000 ;
      RECT  829.515000  1.075000  830.460000 1.275000 ;
      RECT  829.595000  0.255000  831.955000 0.465000 ;
      RECT  829.635000  1.665000  830.015000 2.465000 ;
      RECT  830.375000  1.835000  830.755000 2.635000 ;
      RECT  830.685000  0.465000  830.855000 0.885000 ;
      RECT  830.800000  1.055000  831.405000 1.445000 ;
      RECT  831.025000  0.635000  831.405000 1.055000 ;
      RECT  831.025000  1.665000  831.405000 2.465000 ;
      RECT  831.625000  0.465000  831.955000 0.905000 ;
      RECT  831.625000  1.445000  831.955000 2.635000 ;
      RECT  831.695000  1.075000  832.025000 1.275000 ;
      RECT  832.225000  0.085000  832.515000 0.810000 ;
      RECT  832.225000  1.470000  832.515000 2.635000 ;
      RECT  832.690000  0.255000  832.945000 0.655000 ;
      RECT  832.690000  0.655000  834.825000 0.905000 ;
      RECT  832.690000  1.445000  832.945000 2.635000 ;
      RECT  832.705000  1.075000  834.435000 1.275000 ;
      RECT  833.115000  0.085000  833.495000 0.485000 ;
      RECT  833.115000  1.445000  840.655000 1.665000 ;
      RECT  833.115000  1.665000  833.495000 2.465000 ;
      RECT  833.715000  0.255000  833.885000 0.655000 ;
      RECT  833.715000  1.835000  833.885000 2.635000 ;
      RECT  834.055000  0.085000  834.435000 0.485000 ;
      RECT  834.055000  1.665000  834.435000 2.465000 ;
      RECT  834.655000  0.255000  836.785000 0.485000 ;
      RECT  834.655000  0.485000  834.825000 0.655000 ;
      RECT  834.655000  1.835000  834.825000 2.635000 ;
      RECT  834.790000  1.075000  836.625000 1.275000 ;
      RECT  834.995000  0.655000  838.715000 0.905000 ;
      RECT  834.995000  1.665000  835.375000 2.465000 ;
      RECT  835.595000  1.835000  835.765000 2.635000 ;
      RECT  835.935000  1.665000  836.315000 2.465000 ;
      RECT  836.535000  1.835000  837.225000 2.635000 ;
      RECT  836.850000  1.075000  838.715000 1.275000 ;
      RECT  836.975000  0.255000  841.130000 0.485000 ;
      RECT  837.395000  1.665000  837.775000 2.465000 ;
      RECT  837.995000  1.835000  838.165000 2.635000 ;
      RECT  838.335000  1.665000  838.715000 2.465000 ;
      RECT  838.970000  1.835000  839.140000 2.635000 ;
      RECT  839.145000  0.655000  840.655000 0.905000 ;
      RECT  839.145000  0.905000  839.425000 1.445000 ;
      RECT  839.335000  1.665000  839.715000 2.465000 ;
      RECT  839.715000  1.075000  841.110000 1.275000 ;
      RECT  839.935000  1.835000  840.105000 2.635000 ;
      RECT  840.275000  1.665000  840.655000 2.465000 ;
      RECT  840.875000  0.485000  841.130000 0.905000 ;
      RECT  840.875000  1.445000  841.135000 2.635000 ;
      RECT  841.425000  0.085000  841.715000 0.810000 ;
      RECT  841.425000  1.470000  841.715000 2.635000 ;
      RECT  841.885000  0.445000  842.270000 0.655000 ;
      RECT  841.885000  0.655000  843.170000 0.825000 ;
      RECT  841.885000  0.825000  842.055000 1.595000 ;
      RECT  841.885000  1.595000  842.305000 1.925000 ;
      RECT  842.225000  0.995000  842.620000 1.325000 ;
      RECT  842.465000  0.085000  842.830000 0.485000 ;
      RECT  842.555000  1.495000  842.805000 2.635000 ;
      RECT  842.810000  0.995000  843.130000 1.325000 ;
      RECT  842.975000  1.495000  844.935000 1.665000 ;
      RECT  842.975000  1.665000  843.355000 2.465000 ;
      RECT  843.000000  0.425000  844.400000 0.595000 ;
      RECT  843.000000  0.595000  843.170000 0.655000 ;
      RECT  843.300000  0.960000  843.560000 1.325000 ;
      RECT  843.340000  0.765000  843.560000 0.960000 ;
      RECT  843.525000  1.835000  843.800000 2.635000 ;
      RECT  843.730000  0.765000  844.025000 1.325000 ;
      RECT  843.975000  1.665000  844.305000 2.465000 ;
      RECT  844.195000  0.595000  844.400000 0.995000 ;
      RECT  844.195000  0.995000  844.505000 1.325000 ;
      RECT  844.575000  0.255000  844.935000 0.835000 ;
      RECT  844.675000  0.835000  844.935000 1.495000 ;
      RECT  844.675000  1.835000  844.890000 2.635000 ;
      RECT  845.105000  0.085000  845.395000 0.810000 ;
      RECT  845.105000  1.470000  845.395000 2.635000 ;
      RECT  845.570000  0.255000  845.825000 0.635000 ;
      RECT  845.570000  0.635000  846.200000 0.805000 ;
      RECT  845.570000  0.995000  845.810000 1.615000 ;
      RECT  845.570000  1.915000  846.200000 2.085000 ;
      RECT  845.570000  2.085000  845.825000 2.465000 ;
      RECT  845.980000  0.805000  846.200000 1.075000 ;
      RECT  845.980000  1.075000  846.815000 1.245000 ;
      RECT  845.980000  1.245000  846.200000 1.915000 ;
      RECT  845.995000  0.085000  846.375000 0.465000 ;
      RECT  845.995000  2.255000  846.815000 2.635000 ;
      RECT  846.565000  0.255000  847.755000 0.465000 ;
      RECT  846.565000  0.465000  846.815000 0.905000 ;
      RECT  846.565000  1.445000  846.815000 2.255000 ;
      RECT  846.985000  0.635000  847.365000 1.445000 ;
      RECT  846.985000  1.445000  850.745000 1.665000 ;
      RECT  846.985000  1.665000  847.365000 2.465000 ;
      RECT  847.585000  0.465000  847.755000 0.635000 ;
      RECT  847.585000  0.635000  848.775000 0.905000 ;
      RECT  847.585000  1.835000  847.755000 2.635000 ;
      RECT  847.640000  1.075000  848.830000 1.275000 ;
      RECT  847.925000  0.255000  849.765000 0.465000 ;
      RECT  847.925000  1.665000  848.305000 2.465000 ;
      RECT  848.525000  1.835000  849.165000 2.635000 ;
      RECT  848.965000  0.635000  850.285000 0.715000 ;
      RECT  848.965000  0.715000  851.270000 0.905000 ;
      RECT  849.090000  1.075000  850.165000 1.275000 ;
      RECT  849.335000  1.665000  849.715000 2.465000 ;
      RECT  849.935000  1.835000  850.195000 2.635000 ;
      RECT  849.985000  0.255000  850.245000 0.615000 ;
      RECT  849.985000  0.615000  850.285000 0.635000 ;
      RECT  850.365000  1.665000  850.745000 2.465000 ;
      RECT  850.500000  1.075000  851.365000 1.275000 ;
      RECT  850.545000  0.085000  850.715000 0.545000 ;
      RECT  850.935000  0.255000  851.270000 0.715000 ;
      RECT  850.965000  1.495000  851.360000 2.635000 ;
      RECT  851.545000  0.085000  851.835000 0.810000 ;
      RECT  851.545000  1.470000  851.835000 2.635000 ;
      RECT  852.010000  0.255000  852.345000 0.735000 ;
      RECT  852.010000  0.735000  852.775000 0.905000 ;
      RECT  852.010000  1.495000  852.775000 1.665000 ;
      RECT  852.010000  1.665000  852.345000 2.465000 ;
      RECT  852.030000  1.075000  852.360000 1.275000 ;
      RECT  852.565000  0.085000  852.815000 0.545000 ;
      RECT  852.565000  1.835000  853.255000 2.635000 ;
      RECT  852.580000  0.905000  852.775000 1.075000 ;
      RECT  852.580000  1.075000  853.895000 1.275000 ;
      RECT  852.580000  1.275000  852.775000 1.495000 ;
      RECT  852.965000  1.495000  853.255000 1.835000 ;
      RECT  853.005000  0.255000  857.095000 0.465000 ;
      RECT  853.005000  0.465000  853.255000 0.905000 ;
      RECT  853.425000  0.635000  854.760000 0.905000 ;
      RECT  853.425000  1.445000  860.905000 1.665000 ;
      RECT  853.425000  1.665000  853.805000 2.465000 ;
      RECT  854.025000  1.835000  854.195000 2.635000 ;
      RECT  854.330000  0.905000  854.760000 1.445000 ;
      RECT  854.365000  1.665000  854.745000 2.465000 ;
      RECT  854.965000  1.835000  855.135000 2.635000 ;
      RECT  855.100000  1.075000  856.960000 1.275000 ;
      RECT  855.305000  0.635000  859.025000 0.905000 ;
      RECT  855.305000  1.665000  855.685000 2.465000 ;
      RECT  855.905000  1.835000  856.075000 2.635000 ;
      RECT  856.245000  1.665000  856.625000 2.465000 ;
      RECT  856.845000  1.835000  857.535000 2.635000 ;
      RECT  857.160000  1.075000  859.030000 1.275000 ;
      RECT  857.285000  0.255000  859.495000 0.465000 ;
      RECT  857.705000  1.665000  858.085000 2.465000 ;
      RECT  858.305000  1.835000  858.475000 2.635000 ;
      RECT  858.645000  1.665000  859.025000 2.465000 ;
      RECT  859.245000  0.465000  859.495000 0.735000 ;
      RECT  859.245000  0.735000  861.380000 0.905000 ;
      RECT  859.245000  1.835000  859.415000 2.635000 ;
      RECT  859.585000  1.075000  861.425000 1.275000 ;
      RECT  859.585000  1.665000  859.965000 2.465000 ;
      RECT  859.715000  0.085000  859.885000 0.545000 ;
      RECT  860.055000  0.255000  860.435000 0.735000 ;
      RECT  860.185000  1.835000  860.355000 2.635000 ;
      RECT  860.525000  1.665000  860.905000 2.465000 ;
      RECT  860.655000  0.085000  860.825000 0.545000 ;
      RECT  860.995000  0.255000  861.380000 0.735000 ;
      RECT  861.125000  1.445000  861.380000 2.635000 ;
      RECT  861.665000  0.085000  861.955000 0.810000 ;
      RECT  861.665000  1.470000  861.955000 2.635000 ;
      RECT  862.125000  0.485000  862.465000 0.715000 ;
      RECT  862.125000  0.715000  863.260000 0.905000 ;
      RECT  862.125000  0.905000  862.300000 2.065000 ;
      RECT  862.125000  2.065000  862.465000 2.465000 ;
      RECT  862.470000  1.075000  862.865000 1.655000 ;
      RECT  862.685000  0.085000  862.920000 0.545000 ;
      RECT  862.685000  1.835000  863.015000 2.635000 ;
      RECT  863.035000  1.075000  863.365000 1.325000 ;
      RECT  863.090000  0.365000  864.280000 0.555000 ;
      RECT  863.090000  0.555000  863.260000 0.715000 ;
      RECT  863.195000  1.495000  864.720000 1.665000 ;
      RECT  863.195000  1.665000  863.525000 2.465000 ;
      RECT  863.535000  0.735000  863.800000 1.325000 ;
      RECT  863.735000  1.835000  864.055000 2.635000 ;
      RECT  864.030000  0.555000  864.280000 1.325000 ;
      RECT  864.230000  1.665000  864.720000 2.005000 ;
      RECT  864.230000  2.005000  864.620000 2.465000 ;
      RECT  864.450000  0.255000  865.040000 0.825000 ;
      RECT  864.450000  0.825000  864.720000 1.495000 ;
      RECT  864.790000  2.175000  865.560000 2.635000 ;
      RECT  864.890000  0.995000  865.165000 1.835000 ;
      RECT  864.890000  1.835000  866.095000 2.005000 ;
      RECT  865.230000  0.085000  865.580000 0.545000 ;
      RECT  865.340000  0.725000  865.750000 1.615000 ;
      RECT  865.750000  0.255000  866.095000 0.545000 ;
      RECT  865.780000  2.005000  866.095000 2.465000 ;
      RECT  865.925000  0.545000  866.095000 1.835000 ;
      RECT  866.265000  0.085000  866.555000 0.810000 ;
      RECT  866.265000  1.470000  866.555000 2.635000 ;
      RECT  866.725000  0.255000  866.985000 0.730000 ;
      RECT  866.725000  0.730000  867.970000 0.900000 ;
      RECT  866.725000  1.070000  866.970000 1.615000 ;
      RECT  866.725000  1.785000  867.970000 1.980000 ;
      RECT  866.725000  1.980000  867.010000 2.440000 ;
      RECT  867.155000  0.085000  867.455000 0.545000 ;
      RECT  867.180000  2.195000  867.455000 2.635000 ;
      RECT  867.200000  1.070000  867.580000 1.615000 ;
      RECT  867.625000  0.255000  868.315000 0.560000 ;
      RECT  867.625000  2.150000  868.315000 2.465000 ;
      RECT  867.800000  0.900000  867.970000 1.785000 ;
      RECT  868.140000  0.560000  868.315000 2.150000 ;
      RECT  868.485000  0.255000  870.615000 0.485000 ;
      RECT  868.485000  0.485000  868.655000 0.585000 ;
      RECT  868.485000  1.495000  868.655000 2.635000 ;
      RECT  868.825000  0.655000  869.270000 1.445000 ;
      RECT  868.825000  1.445000  872.515000 1.665000 ;
      RECT  868.825000  1.665000  869.125000 2.465000 ;
      RECT  869.295000  1.835000  869.595000 2.635000 ;
      RECT  869.585000  1.075000  869.965000 1.275000 ;
      RECT  869.765000  0.655000  871.575000 0.905000 ;
      RECT  869.765000  1.665000  870.145000 2.465000 ;
      RECT  870.135000  1.075000  870.685000 1.445000 ;
      RECT  870.365000  1.835000  871.025000 2.635000 ;
      RECT  870.805000  0.255000  872.045000 0.485000 ;
      RECT  870.880000  1.075000  871.590000 1.275000 ;
      RECT  871.195000  1.665000  871.575000 2.465000 ;
      RECT  871.795000  0.485000  872.045000 0.735000 ;
      RECT  871.795000  0.735000  872.985000 0.905000 ;
      RECT  871.795000  1.835000  871.965000 2.635000 ;
      RECT  871.955000  1.075000  872.935000 1.275000 ;
      RECT  872.135000  1.665000  872.515000 2.465000 ;
      RECT  872.265000  0.085000  872.435000 0.565000 ;
      RECT  872.605000  0.255000  872.985000 0.735000 ;
      RECT  872.735000  1.445000  872.985000 2.635000 ;
      RECT  873.165000  0.085000  873.455000 0.810000 ;
      RECT  873.165000  1.470000  873.455000 2.635000 ;
      RECT  873.625000  0.255000  873.885000 0.635000 ;
      RECT  873.625000  0.635000  875.045000 0.805000 ;
      RECT  873.625000  1.785000  875.045000 1.980000 ;
      RECT  873.625000  1.980000  873.910000 2.440000 ;
      RECT  873.640000  0.995000  873.870000 1.615000 ;
      RECT  874.055000  0.085000  874.435000 0.465000 ;
      RECT  874.080000  2.195000  874.355000 2.635000 ;
      RECT  874.125000  0.995000  874.565000 1.615000 ;
      RECT  874.525000  2.150000  875.385000 2.465000 ;
      RECT  874.655000  0.255000  875.385000 0.465000 ;
      RECT  874.735000  0.805000  875.045000 1.785000 ;
      RECT  875.215000  0.465000  875.385000 1.075000 ;
      RECT  875.215000  1.075000  875.565000 1.305000 ;
      RECT  875.215000  1.305000  875.385000 2.150000 ;
      RECT  875.555000  0.255000  879.565000 0.485000 ;
      RECT  875.555000  0.485000  875.725000 0.905000 ;
      RECT  875.555000  1.495000  875.725000 2.635000 ;
      RECT  875.895000  0.655000  877.555000 0.905000 ;
      RECT  875.895000  1.075000  876.740000 1.245000 ;
      RECT  875.895000  1.445000  883.405000 1.665000 ;
      RECT  875.895000  1.665000  876.195000 2.465000 ;
      RECT  876.365000  1.835000  876.665000 2.635000 ;
      RECT  876.835000  1.665000  877.215000 2.465000 ;
      RECT  877.205000  0.905000  877.555000 1.445000 ;
      RECT  877.435000  1.835000  877.605000 2.635000 ;
      RECT  877.725000  1.075000  879.095000 1.275000 ;
      RECT  877.775000  0.655000  881.550000 0.905000 ;
      RECT  877.775000  1.665000  878.155000 2.465000 ;
      RECT  878.375000  1.835000  878.545000 2.635000 ;
      RECT  878.715000  1.665000  879.095000 2.465000 ;
      RECT  879.365000  1.835000  880.005000 2.635000 ;
      RECT  879.585000  1.075000  881.525000 1.275000 ;
      RECT  879.805000  0.255000  881.915000 0.485000 ;
      RECT  880.205000  1.665000  880.585000 2.465000 ;
      RECT  880.805000  1.835000  880.975000 2.635000 ;
      RECT  881.145000  1.665000  881.525000 2.465000 ;
      RECT  881.745000  0.485000  881.915000 0.655000 ;
      RECT  881.745000  0.655000  883.825000 0.825000 ;
      RECT  881.745000  1.835000  881.915000 2.635000 ;
      RECT  881.935000  1.075000  883.880000 1.275000 ;
      RECT  882.085000  1.665000  882.465000 2.465000 ;
      RECT  882.135000  0.085000  882.465000 0.485000 ;
      RECT  882.685000  1.835000  882.855000 2.635000 ;
      RECT  883.025000  1.665000  883.405000 2.465000 ;
      RECT  883.075000  0.085000  883.405000 0.485000 ;
      RECT  883.625000  1.445000  883.900000 2.635000 ;
      RECT  884.205000  0.085000  884.495000 0.810000 ;
      RECT  884.205000  1.470000  884.495000 2.635000 ;
      RECT  884.665000  1.075000  885.015000 1.325000 ;
      RECT  884.675000  1.495000  885.355000 1.665000 ;
      RECT  884.675000  1.665000  885.005000 2.450000 ;
      RECT  884.685000  0.085000  884.925000 0.895000 ;
      RECT  885.095000  0.255000  885.475000 0.895000 ;
      RECT  885.185000  0.895000  885.355000 1.495000 ;
      RECT  885.625000  1.075000  885.975000 1.325000 ;
      RECT  885.645000  0.085000  886.155000 0.895000 ;
      RECT  885.695000  1.495000  886.205000 2.635000 ;
      RECT  886.505000  0.085000  886.795000 0.810000 ;
      RECT  886.505000  1.470000  886.795000 2.635000 ;
      RECT  886.970000  0.085000  887.245000 0.905000 ;
      RECT  886.970000  1.075000  887.740000 1.275000 ;
      RECT  886.970000  1.455000  888.185000 1.665000 ;
      RECT  886.970000  1.665000  887.245000 2.465000 ;
      RECT  887.415000  0.255000  887.795000 0.725000 ;
      RECT  887.415000  0.725000  888.735000 0.735000 ;
      RECT  887.415000  0.735000  889.190000 0.905000 ;
      RECT  887.415000  1.835000  887.795000 2.635000 ;
      RECT  887.910000  1.075000  888.780000 1.275000 ;
      RECT  888.015000  0.085000  888.185000 0.555000 ;
      RECT  888.015000  1.665000  888.185000 2.295000 ;
      RECT  888.015000  2.295000  889.255000 2.465000 ;
      RECT  888.355000  0.255000  888.735000 0.725000 ;
      RECT  888.355000  1.445000  889.190000 1.665000 ;
      RECT  888.355000  1.665000  888.735000 2.125000 ;
      RECT  888.955000  1.835000  889.255000 2.295000 ;
      RECT  888.975000  0.905000  889.190000 1.445000 ;
      RECT  889.020000  0.085000  889.360000 0.555000 ;
      RECT  889.725000  0.085000  890.015000 0.810000 ;
      RECT  889.725000  1.470000  890.015000 2.635000 ;
      RECT  890.190000  0.085000  890.465000 0.905000 ;
      RECT  890.190000  1.455000  892.425000 1.665000 ;
      RECT  890.190000  1.665000  890.465000 2.465000 ;
      RECT  890.240000  1.075000  892.050000 1.275000 ;
      RECT  890.635000  0.255000  891.015000 0.725000 ;
      RECT  890.635000  0.725000  894.590000 0.905000 ;
      RECT  890.635000  1.835000  891.015000 2.635000 ;
      RECT  891.235000  0.085000  891.405000 0.555000 ;
      RECT  891.235000  1.665000  891.405000 2.465000 ;
      RECT  891.575000  0.255000  891.955000 0.725000 ;
      RECT  891.575000  1.835000  891.875000 2.635000 ;
      RECT  892.045000  1.665000  892.425000 2.295000 ;
      RECT  892.045000  2.295000  894.390000 2.465000 ;
      RECT  892.175000  0.085000  892.345000 0.555000 ;
      RECT  892.420000  1.075000  893.935000 1.275000 ;
      RECT  892.515000  0.255000  892.895000 0.725000 ;
      RECT  892.645000  1.445000  894.590000 1.745000 ;
      RECT  892.645000  1.745000  892.815000 2.125000 ;
      RECT  892.985000  1.935000  893.365000 2.295000 ;
      RECT  893.115000  0.085000  893.285000 0.555000 ;
      RECT  893.455000  0.255000  893.835000 0.725000 ;
      RECT  893.585000  1.745000  893.755000 2.125000 ;
      RECT  893.925000  1.915000  894.390000 2.295000 ;
      RECT  894.055000  0.085000  894.340000 0.555000 ;
      RECT  894.195000  0.905000  894.590000 1.445000 ;
      RECT  894.785000  0.085000  895.075000 0.810000 ;
      RECT  894.785000  1.470000  895.075000 2.635000 ;
      RECT  895.250000  0.085000  895.525000 0.905000 ;
      RECT  895.250000  1.455000  899.325000 1.665000 ;
      RECT  895.250000  1.665000  895.565000 2.465000 ;
      RECT  895.520000  1.075000  899.090000 1.275000 ;
      RECT  895.695000  0.255000  896.075000 0.725000 ;
      RECT  895.695000  0.725000  903.185000 0.905000 ;
      RECT  895.785000  1.835000  896.035000 2.635000 ;
      RECT  896.255000  1.665000  896.505000 2.465000 ;
      RECT  896.295000  0.085000  896.465000 0.555000 ;
      RECT  896.635000  0.255000  897.015000 0.725000 ;
      RECT  896.725000  1.835000  896.975000 2.635000 ;
      RECT  897.195000  1.665000  897.445000 2.465000 ;
      RECT  897.235000  0.085000  897.405000 0.555000 ;
      RECT  897.575000  0.255000  897.955000 0.725000 ;
      RECT  897.665000  1.835000  897.915000 2.635000 ;
      RECT  898.135000  1.665000  898.385000 2.465000 ;
      RECT  898.175000  0.085000  898.345000 0.555000 ;
      RECT  898.515000  0.255000  898.895000 0.725000 ;
      RECT  898.605000  1.835000  898.855000 2.635000 ;
      RECT  899.075000  1.665000  899.325000 2.295000 ;
      RECT  899.075000  2.295000  903.085000 2.465000 ;
      RECT  899.115000  0.085000  899.285000 0.555000 ;
      RECT  899.360000  1.075000  902.450000 1.275000 ;
      RECT  899.455000  0.255000  899.835000 0.725000 ;
      RECT  899.545000  1.445000  903.185000 1.615000 ;
      RECT  899.545000  1.615000  899.795000 2.125000 ;
      RECT  900.015000  1.785000  900.265000 2.295000 ;
      RECT  900.055000  0.085000  900.225000 0.555000 ;
      RECT  900.395000  0.255000  900.775000 0.725000 ;
      RECT  900.485000  1.615000  900.735000 2.125000 ;
      RECT  900.955000  1.785000  901.205000 2.295000 ;
      RECT  900.995000  0.085000  901.165000 0.555000 ;
      RECT  901.335000  0.255000  901.715000 0.725000 ;
      RECT  901.425000  1.615000  901.675000 2.125000 ;
      RECT  901.895000  1.785000  902.145000 2.295000 ;
      RECT  901.935000  0.085000  902.105000 0.555000 ;
      RECT  902.275000  0.255000  902.655000 0.725000 ;
      RECT  902.365000  1.615000  902.615000 2.125000 ;
      RECT  902.620000  0.905000  903.185000 1.445000 ;
      RECT  902.835000  1.785000  903.085000 2.295000 ;
      RECT  902.875000  0.085000  903.165000 0.555000 ;
      RECT  903.525000  0.085000  903.815000 0.810000 ;
      RECT  903.525000  1.470000  903.815000 2.635000 ;
      RECT  903.995000  0.290000  904.245000 1.915000 ;
      RECT  903.995000  1.915000  905.385000 2.085000 ;
      RECT  904.415000  0.975000  904.685000 1.745000 ;
      RECT  904.575000  0.085000  904.865000 0.625000 ;
      RECT  904.675000  2.255000  905.005000 2.635000 ;
      RECT  904.855000  1.065000  905.185000 1.325000 ;
      RECT  905.035000  0.255000  905.415000 0.725000 ;
      RECT  905.035000  0.725000  906.115000 0.895000 ;
      RECT  905.215000  1.495000  905.555000 1.665000 ;
      RECT  905.215000  1.665000  905.385000 1.915000 ;
      RECT  905.385000  1.075000  905.765000 1.325000 ;
      RECT  905.385000  1.325000  905.555000 1.495000 ;
      RECT  905.555000  1.850000  906.115000 2.465000 ;
      RECT  905.635000  0.085000  906.020000 0.555000 ;
      RECT  905.935000  0.895000  906.115000 1.850000 ;
      RECT  906.285000  0.085000  906.575000 0.810000 ;
      RECT  906.285000  1.470000  906.575000 2.635000 ;
      RECT  906.745000  0.085000  907.025000 0.895000 ;
      RECT  906.745000  1.445000  908.005000 1.655000 ;
      RECT  906.745000  1.655000  907.065000 2.465000 ;
      RECT  907.140000  1.065000  907.920000 1.275000 ;
      RECT  907.195000  0.255000  907.595000 0.725000 ;
      RECT  907.195000  0.725000  908.515000 0.895000 ;
      RECT  907.285000  1.825000  907.535000 2.635000 ;
      RECT  907.755000  1.655000  908.005000 2.295000 ;
      RECT  907.755000  2.295000  908.985000 2.465000 ;
      RECT  907.795000  0.085000  907.965000 0.555000 ;
      RECT  908.135000  0.255000  908.515000 0.725000 ;
      RECT  908.225000  0.895000  908.475000 2.125000 ;
      RECT  908.695000  1.445000  908.985000 2.295000 ;
      RECT  908.735000  0.085000  908.905000 0.895000 ;
      RECT  908.735000  1.075000  909.425000 1.245000 ;
      RECT  909.255000  0.445000  909.425000 1.075000 ;
      RECT  909.255000  1.245000  909.425000 2.460000 ;
      RECT  909.620000  1.065000  910.195000 1.275000 ;
      RECT  909.845000  0.085000  910.100000 0.845000 ;
      RECT  909.845000  2.145000  910.095000 2.635000 ;
      RECT  909.930000  1.275000  910.195000 1.965000 ;
      RECT  910.425000  0.085000  910.715000 0.810000 ;
      RECT  910.425000  1.470000  910.715000 2.635000 ;
      RECT  910.885000  0.085000  911.165000 0.905000 ;
      RECT  910.885000  1.455000  913.125000 1.665000 ;
      RECT  910.885000  1.665000  911.165000 2.465000 ;
      RECT  911.160000  1.075000  912.750000 1.275000 ;
      RECT  911.335000  0.255000  911.715000 0.725000 ;
      RECT  911.335000  0.725000  914.535000 0.905000 ;
      RECT  911.335000  1.835000  911.715000 2.635000 ;
      RECT  911.935000  0.085000  912.105000 0.555000 ;
      RECT  911.935000  1.665000  912.105000 2.465000 ;
      RECT  912.275000  0.255000  912.655000 0.725000 ;
      RECT  912.275000  1.835000  912.575000 2.635000 ;
      RECT  912.745000  1.665000  913.125000 2.295000 ;
      RECT  912.745000  2.295000  915.025000 2.465000 ;
      RECT  912.875000  0.085000  913.045000 0.555000 ;
      RECT  913.215000  0.255000  913.595000 0.725000 ;
      RECT  913.345000  0.905000  913.675000 1.415000 ;
      RECT  913.345000  1.415000  914.455000 1.745000 ;
      RECT  913.345000  1.745000  913.515000 2.125000 ;
      RECT  913.685000  1.935000  914.065000 2.295000 ;
      RECT  913.815000  0.085000  913.985000 0.555000 ;
      RECT  913.865000  1.075000  915.555000 1.245000 ;
      RECT  914.155000  0.255000  914.535000 0.725000 ;
      RECT  914.285000  1.745000  914.455000 2.125000 ;
      RECT  914.625000  1.575000  915.025000 2.295000 ;
      RECT  914.755000  0.085000  914.925000 0.905000 ;
      RECT  915.195000  0.255000  915.555000 1.075000 ;
      RECT  915.195000  1.245000  915.555000 2.465000 ;
      RECT  915.725000  1.075000  916.225000 1.320000 ;
      RECT  915.775000  0.085000  916.065000 0.905000 ;
      RECT  915.775000  1.495000  916.180000 2.635000 ;
      RECT  916.405000  0.085000  916.695000 0.810000 ;
      RECT  916.405000  1.470000  916.695000 2.635000 ;
      RECT  916.870000  0.385000  917.125000 0.655000 ;
      RECT  916.870000  0.655000  918.195000 0.825000 ;
      RECT  916.870000  0.995000  917.205000 1.325000 ;
      RECT  916.870000  1.495000  917.205000 2.280000 ;
      RECT  916.870000  2.280000  918.195000 2.450000 ;
      RECT  917.295000  0.085000  917.675000 0.485000 ;
      RECT  917.375000  0.995000  917.855000 1.325000 ;
      RECT  917.375000  1.325000  917.660000 2.005000 ;
      RECT  917.895000  0.385000  918.065000 0.655000 ;
      RECT  918.025000  0.825000  918.195000 2.280000 ;
      RECT  918.235000  0.085000  918.955000 0.485000 ;
      RECT  918.365000  1.835000  918.955000 2.635000 ;
      RECT  918.520000  0.655000  918.985000 1.665000 ;
      RECT  919.165000  0.085000  919.455000 0.810000 ;
      RECT  919.165000  1.470000  919.455000 2.635000 ;
      RECT  919.630000  0.085000  919.905000 0.905000 ;
      RECT  919.675000  1.075000  920.555000 1.285000 ;
      RECT  919.690000  1.455000  921.815000 1.625000 ;
      RECT  919.690000  1.625000  919.945000 2.465000 ;
      RECT  920.075000  0.255000  920.455000 0.725000 ;
      RECT  920.075000  0.725000  923.535000 0.905000 ;
      RECT  920.165000  1.795000  920.415000 2.635000 ;
      RECT  920.635000  1.625000  920.885000 2.465000 ;
      RECT  920.675000  0.085000  920.845000 0.555000 ;
      RECT  920.775000  1.075000  921.815000 1.285000 ;
      RECT  921.015000  0.255000  921.395000 0.725000 ;
      RECT  921.105000  1.795000  921.355000 2.295000 ;
      RECT  921.105000  2.295000  923.400000 2.465000 ;
      RECT  921.575000  1.625000  921.815000 2.125000 ;
      RECT  921.615000  0.085000  922.420000 0.555000 ;
      RECT  921.985000  1.075000  922.850000 1.285000 ;
      RECT  921.985000  1.285000  922.475000 1.625000 ;
      RECT  922.250000  1.795000  922.460000 2.295000 ;
      RECT  922.590000  0.255000  922.970000 0.725000 ;
      RECT  922.720000  1.455000  923.535000 1.625000 ;
      RECT  922.720000  1.625000  922.930000 2.125000 ;
      RECT  923.020000  0.905000  923.535000 1.455000 ;
      RECT  923.150000  1.795000  923.400000 2.295000 ;
      RECT  923.190000  0.085000  923.480000 0.555000 ;
      RECT  923.765000  0.085000  924.055000 0.810000 ;
      RECT  923.765000  1.470000  924.055000 2.635000 ;
      RECT  924.230000  0.085000  924.505000 0.905000 ;
      RECT  924.230000  1.075000  926.165000 1.285000 ;
      RECT  924.290000  1.455000  926.425000 1.625000 ;
      RECT  924.290000  1.625000  924.545000 2.465000 ;
      RECT  924.675000  0.255000  925.055000 0.725000 ;
      RECT  924.675000  0.725000  930.485000 0.905000 ;
      RECT  924.765000  1.795000  925.015000 2.635000 ;
      RECT  925.235000  1.625000  925.485000 2.465000 ;
      RECT  925.275000  0.085000  925.445000 0.555000 ;
      RECT  925.615000  0.255000  925.995000 0.725000 ;
      RECT  925.705000  1.795000  925.955000 2.635000 ;
      RECT  926.175000  1.625000  926.425000 2.085000 ;
      RECT  926.175000  2.085000  927.365000 2.465000 ;
      RECT  926.215000  0.085000  926.385000 0.555000 ;
      RECT  926.435000  1.075000  928.225000 1.285000 ;
      RECT  926.555000  0.255000  926.935000 0.725000 ;
      RECT  926.645000  1.455000  927.835000 1.625000 ;
      RECT  926.645000  1.625000  926.895000 1.915000 ;
      RECT  927.115000  1.795000  927.365000 2.085000 ;
      RECT  927.155000  0.085000  927.325000 0.555000 ;
      RECT  927.495000  0.255000  927.875000 0.725000 ;
      RECT  927.585000  1.625000  927.835000 2.295000 ;
      RECT  927.585000  2.295000  929.715000 2.465000 ;
      RECT  928.055000  1.285000  928.225000 1.445000 ;
      RECT  928.055000  1.445000  929.855000 1.615000 ;
      RECT  928.055000  1.785000  930.485000 1.955000 ;
      RECT  928.055000  1.955000  929.245000 1.965000 ;
      RECT  928.055000  1.965000  928.305000 2.125000 ;
      RECT  928.095000  0.085000  928.265000 0.555000 ;
      RECT  928.395000  1.075000  929.455000 1.275000 ;
      RECT  928.435000  0.255000  928.815000 0.725000 ;
      RECT  928.525000  2.135000  928.775000 2.295000 ;
      RECT  928.995000  1.965000  929.245000 2.125000 ;
      RECT  929.035000  0.085000  929.205000 0.555000 ;
      RECT  929.375000  0.255000  929.755000 0.725000 ;
      RECT  929.465000  2.135000  929.715000 2.295000 ;
      RECT  929.685000  1.075000  930.025000 1.285000 ;
      RECT  929.685000  1.285000  929.855000 1.445000 ;
      RECT  929.935000  2.125000  930.185000 2.465000 ;
      RECT  929.975000  0.085000  930.145000 0.555000 ;
      RECT  930.195000  0.905000  930.485000 1.785000 ;
      RECT  930.665000  0.085000  930.955000 0.810000 ;
      RECT  930.665000  1.470000  930.955000 2.635000 ;
      RECT  931.125000  0.255000  931.645000 0.655000 ;
      RECT  931.125000  0.655000  932.585000 0.825000 ;
      RECT  931.125000  0.825000  931.295000 1.445000 ;
      RECT  931.125000  1.445000  931.585000 2.455000 ;
      RECT  931.465000  1.075000  931.925000 1.245000 ;
      RECT  931.755000  1.245000  931.925000 1.785000 ;
      RECT  931.755000  1.785000  933.715000 1.955000 ;
      RECT  931.815000  0.085000  932.195000 0.485000 ;
      RECT  932.095000  0.995000  932.345000 1.615000 ;
      RECT  932.415000  0.310000  932.585000 0.655000 ;
      RECT  932.515000  0.995000  932.855000 1.615000 ;
      RECT  932.755000  0.085000  933.135000 0.825000 ;
      RECT  932.755000  2.125000  933.135000 2.635000 ;
      RECT  933.025000  0.995000  933.375000 1.615000 ;
      RECT  933.420000  0.405000  933.590000 0.655000 ;
      RECT  933.420000  0.655000  933.715000 0.825000 ;
      RECT  933.545000  0.825000  933.715000 1.785000 ;
      RECT  933.885000  0.085000  934.175000 0.810000 ;
      RECT  933.885000  1.470000  934.175000 2.635000 ;
      RECT  934.350000  0.085000  934.625000 0.905000 ;
      RECT  934.350000  1.455000  936.585000 1.625000 ;
      RECT  934.350000  1.625000  934.665000 2.465000 ;
      RECT  934.370000  1.075000  935.275000 1.285000 ;
      RECT  934.795000  0.255000  935.175000 0.725000 ;
      RECT  934.795000  0.725000  937.615000 0.905000 ;
      RECT  934.885000  1.795000  935.135000 2.635000 ;
      RECT  935.355000  1.625000  935.605000 2.465000 ;
      RECT  935.395000  0.085000  935.565000 0.555000 ;
      RECT  935.495000  1.075000  936.460000 1.285000 ;
      RECT  935.735000  0.255000  936.115000 0.725000 ;
      RECT  935.825000  1.795000  936.075000 2.275000 ;
      RECT  935.825000  2.275000  938.040000 2.465000 ;
      RECT  936.255000  1.625000  936.585000 2.035000 ;
      RECT  936.335000  0.085000  937.025000 0.555000 ;
      RECT  937.130000  0.905000  937.615000 2.045000 ;
      RECT  937.195000  0.255000  937.615000 0.725000 ;
      RECT  937.795000  1.075000  938.420000 1.285000 ;
      RECT  937.795000  1.455000  938.040000 2.275000 ;
      RECT  937.835000  0.085000  938.040000 0.895000 ;
      RECT  938.250000  0.380000  938.605000 0.905000 ;
      RECT  938.250000  0.905000  938.420000 1.075000 ;
      RECT  938.250000  1.285000  938.420000 1.455000 ;
      RECT  938.250000  1.455000  938.605000 1.870000 ;
      RECT  938.590000  1.075000  939.175000 1.285000 ;
      RECT  938.825000  0.085000  939.115000 0.825000 ;
      RECT  938.825000  1.540000  939.075000 2.635000 ;
      RECT  939.405000  0.085000  939.695000 0.810000 ;
      RECT  939.405000  1.470000  939.695000 2.635000 ;
      RECT  939.890000  0.255000  940.225000 0.735000 ;
      RECT  939.890000  0.735000  940.615000 0.905000 ;
      RECT  939.890000  1.075000  940.225000 1.285000 ;
      RECT  939.890000  1.455000  944.935000 1.625000 ;
      RECT  939.890000  1.625000  940.185000 2.465000 ;
      RECT  940.405000  1.795000  940.655000 2.635000 ;
      RECT  940.445000  0.085000  940.615000 0.555000 ;
      RECT  940.445000  0.905000  940.615000 1.455000 ;
      RECT  940.785000  0.255000  941.165000 0.725000 ;
      RECT  940.785000  0.725000  947.025000 0.905000 ;
      RECT  940.875000  1.795000  944.465000 1.965000 ;
      RECT  940.875000  1.965000  941.125000 2.465000 ;
      RECT  940.990000  1.075000  942.550000 1.285000 ;
      RECT  941.345000  2.135000  941.595000 2.635000 ;
      RECT  941.385000  0.085000  941.555000 0.555000 ;
      RECT  941.725000  0.255000  942.105000 0.725000 ;
      RECT  941.815000  1.965000  942.065000 2.465000 ;
      RECT  942.285000  2.135000  942.535000 2.635000 ;
      RECT  942.325000  0.085000  943.015000 0.555000 ;
      RECT  942.805000  2.135000  943.055000 2.295000 ;
      RECT  942.805000  2.295000  946.815000 2.465000 ;
      RECT  943.065000  1.075000  944.480000 1.285000 ;
      RECT  943.185000  0.255000  943.565000 0.725000 ;
      RECT  943.275000  1.965000  943.525000 2.125000 ;
      RECT  943.745000  2.135000  943.995000 2.295000 ;
      RECT  943.785000  0.085000  943.955000 0.555000 ;
      RECT  944.125000  0.255000  944.505000 0.725000 ;
      RECT  944.215000  1.965000  944.465000 2.125000 ;
      RECT  944.685000  1.795000  944.935000 2.295000 ;
      RECT  944.725000  0.085000  944.895000 0.555000 ;
      RECT  944.765000  1.075000  946.500000 1.285000 ;
      RECT  944.765000  1.285000  944.935000 1.455000 ;
      RECT  945.065000  0.255000  945.445000 0.725000 ;
      RECT  945.155000  1.455000  947.025000 1.625000 ;
      RECT  945.155000  1.625000  945.405000 2.125000 ;
      RECT  945.625000  1.795000  945.875000 2.295000 ;
      RECT  945.665000  0.085000  945.835000 0.555000 ;
      RECT  946.005000  0.255000  946.385000 0.725000 ;
      RECT  946.095000  1.625000  946.345000 2.125000 ;
      RECT  946.565000  1.795000  946.815000 2.295000 ;
      RECT  946.605000  0.085000  946.775000 0.555000 ;
      RECT  946.685000  0.905000  947.025000 1.455000 ;
      RECT  947.225000  0.085000  947.515000 0.810000 ;
      RECT  947.225000  1.470000  947.515000 2.635000 ;
      RECT  947.685000  0.085000  947.945000 0.575000 ;
      RECT  947.685000  0.745000  947.935000 1.325000 ;
      RECT  947.690000  1.495000  948.375000 1.665000 ;
      RECT  947.690000  1.665000  948.025000 2.450000 ;
      RECT  948.115000  0.385000  948.415000 0.655000 ;
      RECT  948.115000  0.655000  949.365000 0.825000 ;
      RECT  948.115000  0.825000  948.375000 1.495000 ;
      RECT  948.565000  0.995000  948.885000 2.450000 ;
      RECT  948.635000  0.085000  948.965000 0.485000 ;
      RECT  949.055000  0.995000  949.345000 2.450000 ;
      RECT  949.195000  0.385000  949.365000 0.655000 ;
      RECT  949.535000  0.655000  949.805000 1.665000 ;
      RECT  949.605000  0.085000  950.120000 0.485000 ;
      RECT  949.735000  1.835000  950.135000 2.635000 ;
      RECT  950.445000  0.085000  950.735000 0.810000 ;
      RECT  950.445000  1.470000  950.735000 2.635000 ;
      RECT  950.910000  0.085000  951.185000 0.905000 ;
      RECT  950.970000  1.455000  953.105000 1.625000 ;
      RECT  950.970000  1.625000  951.225000 2.465000 ;
      RECT  951.020000  1.075000  951.835000 1.285000 ;
      RECT  951.390000  0.255000  951.770000 0.725000 ;
      RECT  951.390000  0.725000  955.770000 0.905000 ;
      RECT  951.445000  1.795000  951.695000 2.635000 ;
      RECT  951.915000  1.625000  952.165000 2.465000 ;
      RECT  951.955000  0.085000  952.125000 0.555000 ;
      RECT  952.055000  1.075000  952.960000 1.285000 ;
      RECT  952.330000  0.255000  952.710000 0.725000 ;
      RECT  952.385000  1.795000  952.635000 2.295000 ;
      RECT  952.385000  2.295000  954.135000 2.465000 ;
      RECT  952.855000  1.625000  953.105000 2.125000 ;
      RECT  952.895000  0.085000  953.625000 0.555000 ;
      RECT  953.230000  1.075000  954.175000 1.285000 ;
      RECT  953.415000  1.455000  954.605000 1.625000 ;
      RECT  953.415000  1.625000  953.665000 2.125000 ;
      RECT  953.830000  0.255000  954.210000 0.725000 ;
      RECT  953.885000  1.795000  954.135000 2.295000 ;
      RECT  954.355000  1.625000  954.605000 2.295000 ;
      RECT  954.355000  2.295000  955.545000 2.465000 ;
      RECT  954.395000  0.085000  954.565000 0.555000 ;
      RECT  954.460000  1.075000  955.095000 1.285000 ;
      RECT  954.770000  0.255000  955.150000 0.725000 ;
      RECT  954.860000  1.455000  955.770000 1.625000 ;
      RECT  954.860000  1.625000  955.110000 2.125000 ;
      RECT  955.295000  1.795000  955.545000 2.295000 ;
      RECT  955.335000  0.085000  955.625000 0.555000 ;
      RECT  955.435000  0.905000  955.770000 1.455000 ;
      RECT  955.965000  0.085000  956.255000 0.810000 ;
      RECT  955.965000  1.470000  956.255000 2.635000 ;
      RECT  956.430000  0.085000  956.705000 0.905000 ;
      RECT  956.430000  1.455000  958.625000 1.625000 ;
      RECT  956.430000  1.625000  956.745000 2.465000 ;
      RECT  956.520000  1.075000  958.365000 1.285000 ;
      RECT  956.875000  0.255000  957.255000 0.725000 ;
      RECT  956.875000  0.725000  964.970000 0.905000 ;
      RECT  956.965000  1.795000  957.215000 2.635000 ;
      RECT  957.435000  1.625000  957.685000 2.465000 ;
      RECT  957.475000  0.085000  957.645000 0.555000 ;
      RECT  957.815000  0.255000  958.195000 0.725000 ;
      RECT  957.905000  1.795000  958.155000 2.635000 ;
      RECT  958.375000  1.625000  958.625000 2.295000 ;
      RECT  958.375000  2.295000  960.560000 2.465000 ;
      RECT  958.415000  0.085000  958.585000 0.555000 ;
      RECT  958.635000  1.075000  960.810000 1.285000 ;
      RECT  958.755000  0.255000  959.135000 0.725000 ;
      RECT  958.845000  1.455000  962.435000 1.625000 ;
      RECT  958.845000  1.625000  959.095000 2.125000 ;
      RECT  959.315000  1.795000  959.565000 2.295000 ;
      RECT  959.355000  0.085000  959.525000 0.555000 ;
      RECT  959.695000  0.255000  960.075000 0.725000 ;
      RECT  959.785000  1.625000  960.035000 2.125000 ;
      RECT  960.255000  1.795000  960.560000 2.295000 ;
      RECT  960.295000  0.085000  960.985000 0.555000 ;
      RECT  960.745000  1.795000  961.025000 2.295000 ;
      RECT  960.745000  2.295000  964.785000 2.465000 ;
      RECT  961.035000  1.075000  962.645000 1.285000 ;
      RECT  961.155000  0.255000  961.535000 0.725000 ;
      RECT  961.245000  1.625000  961.495000 2.125000 ;
      RECT  961.715000  1.795000  961.965000 2.295000 ;
      RECT  961.755000  0.085000  961.925000 0.555000 ;
      RECT  962.095000  0.255000  962.475000 0.725000 ;
      RECT  962.185000  1.625000  962.435000 2.125000 ;
      RECT  962.655000  1.795000  962.905000 2.295000 ;
      RECT  962.695000  0.085000  962.865000 0.555000 ;
      RECT  962.815000  1.075000  964.385000 1.285000 ;
      RECT  963.035000  0.255000  963.415000 0.725000 ;
      RECT  963.125000  1.455000  964.970000 1.625000 ;
      RECT  963.125000  1.625000  963.375000 2.125000 ;
      RECT  963.595000  1.795000  963.845000 2.295000 ;
      RECT  963.635000  0.085000  963.805000 0.555000 ;
      RECT  963.975000  0.255000  964.355000 0.725000 ;
      RECT  964.065000  1.625000  964.315000 2.125000 ;
      RECT  964.535000  1.795000  964.785000 2.295000 ;
      RECT  964.575000  0.085000  964.745000 0.555000 ;
      RECT  964.700000  0.905000  964.970000 1.455000 ;
      RECT  965.165000  0.085000  965.455000 0.810000 ;
      RECT  965.165000  1.470000  965.455000 2.635000 ;
      RECT  965.625000  0.655000  967.615000 0.825000 ;
      RECT  965.625000  0.825000  965.885000 2.450000 ;
      RECT  965.895000  0.085000  966.225000 0.480000 ;
      RECT  966.065000  0.995000  966.285000 1.795000 ;
      RECT  966.065000  1.795000  969.105000 2.005000 ;
      RECT  966.445000  0.300000  966.645000 0.655000 ;
      RECT  966.475000  0.995000  966.825000 1.615000 ;
      RECT  966.865000  0.085000  967.195000 0.485000 ;
      RECT  967.015000  0.995000  967.475000 1.615000 ;
      RECT  967.415000  0.310000  967.615000 0.655000 ;
      RECT  967.715000  0.995000  968.195000 1.615000 ;
      RECT  967.785000  0.085000  968.275000 0.825000 ;
      RECT  967.865000  2.185000  968.245000 2.635000 ;
      RECT  968.365000  0.995000  968.765000 1.615000 ;
      RECT  968.630000  0.405000  968.800000 0.655000 ;
      RECT  968.630000  0.655000  969.105000 0.825000 ;
      RECT  968.935000  0.825000  969.105000 1.795000 ;
      RECT  969.305000  0.085000  969.595000 0.810000 ;
      RECT  969.305000  1.470000  969.595000 2.635000 ;
      RECT  969.765000  0.085000  970.025000 0.905000 ;
      RECT  969.765000  1.455000  971.985000 1.625000 ;
      RECT  969.765000  1.625000  970.105000 2.465000 ;
      RECT  969.780000  1.075000  971.020000 1.285000 ;
      RECT  970.195000  0.255000  970.575000 0.725000 ;
      RECT  970.195000  0.725000  973.950000 0.905000 ;
      RECT  970.325000  1.795000  970.535000 2.635000 ;
      RECT  970.755000  1.625000  971.005000 2.465000 ;
      RECT  970.795000  0.085000  970.965000 0.555000 ;
      RECT  971.135000  0.255000  971.515000 0.725000 ;
      RECT  971.205000  1.075000  972.330000 1.285000 ;
      RECT  971.225000  1.795000  971.435000 2.295000 ;
      RECT  971.225000  2.295000  972.970000 2.465000 ;
      RECT  971.605000  1.625000  971.985000 2.125000 ;
      RECT  971.735000  0.085000  972.460000 0.555000 ;
      RECT  972.155000  1.455000  973.440000 1.625000 ;
      RECT  972.155000  1.625000  972.540000 2.125000 ;
      RECT  972.540000  1.075000  973.340000 1.285000 ;
      RECT  972.630000  0.255000  973.010000 0.725000 ;
      RECT  972.760000  1.795000  972.970000 2.295000 ;
      RECT  973.190000  1.625000  973.440000 2.295000 ;
      RECT  973.190000  2.295000  974.375000 2.465000 ;
      RECT  973.230000  0.085000  973.400000 0.555000 ;
      RECT  973.570000  0.255000  973.950000 0.725000 ;
      RECT  973.660000  1.455000  974.170000 1.625000 ;
      RECT  973.660000  1.625000  973.910000 2.125000 ;
      RECT  973.745000  0.905000  973.950000 1.075000 ;
      RECT  973.745000  1.075000  974.170000 1.455000 ;
      RECT  974.130000  1.795000  974.375000 2.295000 ;
      RECT  974.170000  0.085000  974.375000 0.895000 ;
      RECT  974.400000  1.075000  974.715000 1.245000 ;
      RECT  974.545000  0.380000  974.900000 0.905000 ;
      RECT  974.545000  0.905000  974.715000 1.075000 ;
      RECT  974.545000  1.245000  974.715000 2.035000 ;
      RECT  974.545000  2.035000  974.900000 2.450000 ;
      RECT  974.885000  1.075000  975.565000 1.285000 ;
      RECT  975.120000  0.085000  975.370000 0.825000 ;
      RECT  975.120000  2.135000  975.370000 2.635000 ;
      RECT  975.295000  1.285000  975.565000 1.955000 ;
      RECT  975.745000  0.085000  976.035000 0.810000 ;
      RECT  975.745000  1.470000  976.035000 2.635000 ;
      RECT  976.215000  1.455000  978.385000 1.625000 ;
      RECT  976.215000  1.625000  976.545000 2.465000 ;
      RECT  976.295000  0.085000  976.465000 0.895000 ;
      RECT  976.515000  1.075000  978.125000 1.285000 ;
      RECT  976.635000  0.255000  977.015000 0.725000 ;
      RECT  976.635000  0.725000  984.115000 0.905000 ;
      RECT  976.765000  1.795000  976.975000 2.635000 ;
      RECT  977.195000  1.625000  977.445000 2.465000 ;
      RECT  977.235000  0.085000  977.405000 0.555000 ;
      RECT  977.575000  0.255000  977.955000 0.725000 ;
      RECT  977.665000  1.795000  977.915000 2.635000 ;
      RECT  978.135000  1.625000  978.385000 2.295000 ;
      RECT  978.135000  2.295000  980.265000 2.465000 ;
      RECT  978.175000  0.085000  978.345000 0.555000 ;
      RECT  978.395000  1.075000  980.270000 1.285000 ;
      RECT  978.515000  0.255000  978.895000 0.725000 ;
      RECT  978.605000  1.455000  982.195000 1.625000 ;
      RECT  978.605000  1.625000  978.855000 2.125000 ;
      RECT  979.075000  1.795000  979.325000 2.295000 ;
      RECT  979.115000  0.085000  979.285000 0.555000 ;
      RECT  979.455000  0.255000  979.835000 0.725000 ;
      RECT  979.545000  1.625000  979.795000 2.125000 ;
      RECT  980.015000  1.795000  980.265000 2.295000 ;
      RECT  980.055000  0.085000  980.745000 0.555000 ;
      RECT  980.505000  1.075000  982.405000 1.285000 ;
      RECT  980.535000  1.795000  980.785000 2.295000 ;
      RECT  980.535000  2.295000  984.545000 2.465000 ;
      RECT  980.915000  0.255000  981.295000 0.725000 ;
      RECT  981.005000  1.625000  981.255000 2.125000 ;
      RECT  981.475000  1.795000  981.725000 2.295000 ;
      RECT  981.515000  0.085000  981.685000 0.555000 ;
      RECT  981.855000  0.255000  982.235000 0.725000 ;
      RECT  981.945000  1.625000  982.195000 2.125000 ;
      RECT  982.415000  1.455000  982.665000 2.295000 ;
      RECT  982.455000  0.085000  982.625000 0.555000 ;
      RECT  982.795000  0.255000  983.175000 0.725000 ;
      RECT  982.885000  0.905000  983.370000 1.455000 ;
      RECT  982.885000  1.455000  984.075000 1.625000 ;
      RECT  982.885000  1.625000  983.135000 2.125000 ;
      RECT  983.355000  1.795000  983.605000 2.295000 ;
      RECT  983.395000  0.085000  983.565000 0.555000 ;
      RECT  983.540000  1.075000  984.560000 1.285000 ;
      RECT  983.735000  0.255000  984.115000 0.725000 ;
      RECT  983.825000  1.625000  984.075000 2.125000 ;
      RECT  984.295000  1.795000  984.545000 2.295000 ;
      RECT  984.335000  0.085000  984.505000 0.555000 ;
      RECT  984.390000  0.735000  985.105000 0.905000 ;
      RECT  984.390000  0.905000  984.560000 1.075000 ;
      RECT  984.390000  1.285000  984.560000 1.455000 ;
      RECT  984.390000  1.455000  985.105000 1.625000 ;
      RECT  984.730000  0.255000  985.105000 0.735000 ;
      RECT  984.770000  1.625000  985.105000 2.465000 ;
      RECT  984.975000  1.075000  985.670000 1.285000 ;
      RECT  985.325000  0.085000  985.555000 0.905000 ;
      RECT  985.325000  1.455000  985.555000 2.635000 ;
      RECT  985.865000  0.085000  986.155000 0.810000 ;
      RECT  985.865000  1.470000  986.155000 2.635000 ;
      RECT  986.325000  0.450000  986.645000 0.825000 ;
      RECT  986.325000  0.825000  986.500000 1.885000 ;
      RECT  986.325000  1.885000  987.545000 2.070000 ;
      RECT  986.325000  2.070000  986.585000 2.455000 ;
      RECT  986.670000  0.995000  987.070000 1.695000 ;
      RECT  986.755000  2.240000  987.135000 2.635000 ;
      RECT  986.945000  0.085000  987.115000 0.825000 ;
      RECT  987.240000  0.995000  987.580000 1.325000 ;
      RECT  987.340000  1.525000  988.030000 1.715000 ;
      RECT  987.375000  2.070000  987.545000 2.295000 ;
      RECT  987.375000  2.295000  988.855000 2.465000 ;
      RECT  987.415000  0.450000  987.585000 0.655000 ;
      RECT  987.415000  0.655000  988.030000 0.825000 ;
      RECT  987.815000  1.955000  988.450000 2.125000 ;
      RECT  987.860000  0.085000  988.190000 0.480000 ;
      RECT  987.860000  0.825000  988.030000 1.525000 ;
      RECT  988.200000  0.655000  989.580000 0.825000 ;
      RECT  988.200000  0.825000  988.450000 1.955000 ;
      RECT  988.410000  0.300000  988.610000 0.655000 ;
      RECT  988.620000  0.995000  988.855000 2.295000 ;
      RECT  988.830000  0.085000  989.160000 0.485000 ;
      RECT  989.060000  0.995000  989.370000 2.410000 ;
      RECT  989.380000  0.310000  989.580000 0.655000 ;
      RECT  989.600000  0.995000  989.905000 1.705000 ;
      RECT  989.750000  0.085000  990.230000 0.825000 ;
      RECT  989.750000  1.875000  990.230000 2.635000 ;
      RECT  990.465000  0.085000  990.755000 0.810000 ;
      RECT  990.465000  1.470000  990.755000 2.635000 ;
      RECT  990.925000  0.450000  991.305000 0.825000 ;
      RECT  990.925000  0.825000  991.095000 1.885000 ;
      RECT  990.925000  1.885000  992.790000 2.055000 ;
      RECT  990.925000  2.055000  991.185000 2.455000 ;
      RECT  991.265000  0.995000  991.670000 1.695000 ;
      RECT  991.355000  2.240000  991.735000 2.635000 ;
      RECT  991.525000  0.085000  991.695000 0.825000 ;
      RECT  991.840000  0.995000  992.110000 1.325000 ;
      RECT  991.885000  1.525000  992.450000 1.715000 ;
      RECT  991.995000  0.450000  992.190000 0.655000 ;
      RECT  991.995000  0.655000  992.450000 0.825000 ;
      RECT  992.280000  0.825000  992.450000 1.075000 ;
      RECT  992.280000  1.075000  993.315000 1.245000 ;
      RECT  992.280000  1.245000  992.450000 1.525000 ;
      RECT  992.435000  0.085000  992.765000 0.480000 ;
      RECT  992.515000  2.225000  994.725000 2.465000 ;
      RECT  992.620000  1.415000  993.705000 1.585000 ;
      RECT  992.620000  1.585000  992.790000 1.885000 ;
      RECT  992.935000  0.255000  993.315000 0.725000 ;
      RECT  992.935000  0.725000  996.675000 0.905000 ;
      RECT  992.985000  1.875000  995.735000 2.045000 ;
      RECT  993.535000  0.085000  993.705000 0.555000 ;
      RECT  993.535000  1.075000  994.480000 1.275000 ;
      RECT  993.535000  1.275000  993.705000 1.415000 ;
      RECT  993.875000  0.255000  994.255000 0.725000 ;
      RECT  993.875000  1.445000  995.070000 1.705000 ;
      RECT  994.475000  0.085000  995.185000 0.555000 ;
      RECT  994.650000  0.905000  995.070000 1.445000 ;
      RECT  994.935000  2.215000  996.165000 2.465000 ;
      RECT  995.240000  1.075000  996.135000 1.275000 ;
      RECT  995.355000  0.255000  995.735000 0.725000 ;
      RECT  995.445000  1.455000  995.735000 1.875000 ;
      RECT  995.955000  0.085000  996.125000 0.555000 ;
      RECT  995.955000  1.455000  997.145000 1.625000 ;
      RECT  995.955000  1.625000  996.165000 2.215000 ;
      RECT  996.295000  0.255000  996.675000 0.725000 ;
      RECT  996.305000  1.075000  997.170000 1.275000 ;
      RECT  996.385000  1.795000  996.595000 2.635000 ;
      RECT  996.765000  1.625000  997.145000 2.465000 ;
      RECT  996.895000  0.085000  997.170000 0.905000 ;
      RECT  997.365000  0.085000  997.655000 0.810000 ;
      RECT  997.365000  1.470000  997.655000 2.635000 ;
      RECT  997.825000  0.255000  998.185000 0.725000 ;
      RECT  997.825000  0.725000  998.575000 0.895000 ;
      RECT  997.825000  1.535000  998.575000 1.875000 ;
      RECT  997.825000  1.875000 1001.565000 2.045000 ;
      RECT  997.825000  2.045000  998.105000 2.465000 ;
      RECT  997.850000  1.075000  998.185000 1.365000 ;
      RECT  998.275000  2.215000  998.655000 2.635000 ;
      RECT  998.405000  0.085000  998.575000 0.555000 ;
      RECT  998.405000  0.895000  998.575000 1.535000 ;
      RECT  998.745000  0.255000  999.125000 0.735000 ;
      RECT  998.745000  0.735000  999.475000 0.905000 ;
      RECT  998.745000  1.075000  999.135000 1.325000 ;
      RECT  998.745000  1.535000  999.475000 1.705000 ;
      RECT  999.305000  0.905000  999.475000 1.075000 ;
      RECT  999.305000  1.075000 1000.835000 1.245000 ;
      RECT  999.305000  1.245000  999.475000 1.535000 ;
      RECT  999.355000  2.215000 1001.565000 2.295000 ;
      RECT  999.355000  2.295000 1003.435000 2.465000 ;
      RECT  999.435000  0.085000  999.605000 0.555000 ;
      RECT  999.680000  1.415000 1001.175000 1.705000 ;
      RECT  999.775000  0.255000 1000.155000 0.725000 ;
      RECT  999.775000  0.725000 1007.255000 0.905000 ;
      RECT 1000.375000  0.085000 1000.545000 0.555000 ;
      RECT 1000.715000  0.255000 1001.095000 0.725000 ;
      RECT 1001.005000  0.905000 1001.175000 1.415000 ;
      RECT 1001.315000  0.085000 1001.485000 0.555000 ;
      RECT 1001.395000  1.075000 1003.145000 1.285000 ;
      RECT 1001.395000  1.285000 1001.565000 1.875000 ;
      RECT 1001.655000  0.255000 1002.035000 0.725000 ;
      RECT 1001.785000  1.455000 1005.335000 1.625000 ;
      RECT 1001.785000  1.625000 1001.995000 2.125000 ;
      RECT 1002.215000  1.795000 1002.465000 2.295000 ;
      RECT 1002.255000  0.085000 1002.425000 0.555000 ;
      RECT 1002.595000  0.255000 1002.975000 0.725000 ;
      RECT 1002.685000  1.625000 1002.935000 2.125000 ;
      RECT 1003.155000  1.795000 1003.435000 2.295000 ;
      RECT 1003.195000  0.085000 1003.885000 0.555000 ;
      RECT 1003.390000  1.075000 1005.545000 1.285000 ;
      RECT 1003.620000  1.795000 1003.925000 2.295000 ;
      RECT 1003.620000  2.295000 1005.805000 2.465000 ;
      RECT 1004.055000  0.255000 1004.435000 0.725000 ;
      RECT 1004.145000  1.625000 1004.395000 2.125000 ;
      RECT 1004.615000  1.795000 1004.865000 2.295000 ;
      RECT 1004.655000  0.085000 1004.825000 0.555000 ;
      RECT 1004.995000  0.255000 1005.375000 0.725000 ;
      RECT 1005.085000  1.625000 1005.335000 2.125000 ;
      RECT 1005.555000  1.455000 1007.750000 1.625000 ;
      RECT 1005.555000  1.625000 1005.805000 2.295000 ;
      RECT 1005.595000  0.085000 1005.765000 0.555000 ;
      RECT 1005.815000  1.075000 1007.750000 1.285000 ;
      RECT 1005.935000  0.255000 1006.315000 0.725000 ;
      RECT 1006.025000  1.795000 1006.275000 2.635000 ;
      RECT 1006.495000  1.625000 1006.745000 2.465000 ;
      RECT 1006.535000  0.085000 1006.705000 0.555000 ;
      RECT 1006.875000  0.255000 1007.255000 0.725000 ;
      RECT 1006.965000  1.795000 1007.215000 2.635000 ;
      RECT 1007.435000  1.625000 1007.750000 2.465000 ;
      RECT 1007.475000  0.085000 1007.750000 0.905000 ;
      RECT 1007.945000  0.085000 1008.235000 0.810000 ;
      RECT 1007.945000  1.470000 1008.235000 2.635000 ;
      RECT 1008.405000  0.255000 1008.745000 0.885000 ;
      RECT 1008.405000  0.885000 1008.580000 1.495000 ;
      RECT 1008.405000  1.495000 1008.745000 2.465000 ;
      RECT 1008.750000  1.075000 1009.495000 1.245000 ;
      RECT 1008.965000  0.085000 1009.215000 0.885000 ;
      RECT 1008.965000  1.495000 1009.135000 2.635000 ;
      RECT 1009.325000  1.245000 1009.495000 1.495000 ;
      RECT 1009.325000  1.495000 1012.120000 1.665000 ;
      RECT 1009.405000  0.255000 1009.735000 0.735000 ;
      RECT 1009.405000  0.735000 1010.730000 0.905000 ;
      RECT 1009.405000  1.835000 1009.655000 2.635000 ;
      RECT 1009.670000  1.075000 1010.135000 1.275000 ;
      RECT 1009.955000  0.085000 1010.180000 0.545000 ;
      RECT 1010.305000  1.075000 1010.690000 1.275000 ;
      RECT 1010.350000  0.255000 1010.730000 0.735000 ;
      RECT 1010.405000  1.665000 1010.785000 2.465000 ;
      RECT 1010.860000  1.075000 1011.400000 1.275000 ;
      RECT 1011.080000  1.835000 1011.410000 2.635000 ;
      RECT 1011.135000  0.435000 1011.400000 1.075000 ;
      RECT 1011.570000  0.255000 1012.120000 0.865000 ;
      RECT 1011.570000  0.865000 1011.790000 1.495000 ;
      RECT 1011.790000  1.665000 1012.120000 2.465000 ;
      RECT 1011.960000  1.075000 1012.325000 1.325000 ;
      RECT 1012.545000  0.085000 1012.835000 0.810000 ;
      RECT 1012.545000  1.470000 1012.835000 2.635000 ;
      RECT 1013.005000  0.995000 1013.280000 1.325000 ;
      RECT 1013.010000  1.510000 1015.945000 1.735000 ;
      RECT 1013.010000  1.735000 1014.740000 1.765000 ;
      RECT 1013.010000  1.765000 1013.275000 2.465000 ;
      RECT 1013.015000  0.255000 1013.350000 0.425000 ;
      RECT 1013.015000  0.425000 1013.680000 0.825000 ;
      RECT 1013.445000  1.935000 1013.825000 2.635000 ;
      RECT 1013.450000  0.825000 1013.680000 1.510000 ;
      RECT 1013.850000  0.635000 1015.295000 0.825000 ;
      RECT 1013.850000  0.995000 1014.230000 1.325000 ;
      RECT 1014.045000  1.765000 1014.740000 2.465000 ;
      RECT 1014.425000  0.995000 1014.865000 1.325000 ;
      RECT 1014.455000  0.085000 1014.790000 0.465000 ;
      RECT 1015.085000  0.995000 1015.595000 1.325000 ;
      RECT 1015.295000  1.935000 1015.775000 2.635000 ;
      RECT 1015.460000  0.085000 1015.695000 0.525000 ;
      RECT 1015.775000  0.995000 1016.485000 1.325000 ;
      RECT 1015.775000  1.325000 1015.945000 1.510000 ;
      RECT 1015.865000  0.255000 1016.245000 0.615000 ;
      RECT 1015.865000  0.615000 1016.955000 0.785000 ;
      RECT 1016.005000  1.905000 1016.955000 2.075000 ;
      RECT 1016.005000  2.075000 1016.195000 2.465000 ;
      RECT 1016.365000  2.255000 1016.745000 2.635000 ;
      RECT 1016.465000  0.085000 1016.795000 0.445000 ;
      RECT 1016.685000  0.785000 1016.955000 1.905000 ;
      RECT 1017.145000  0.085000 1017.435000 0.810000 ;
      RECT 1017.145000  1.470000 1017.435000 2.635000 ;
      RECT 1017.605000  0.635000 1019.275000 0.805000 ;
      RECT 1017.605000  0.805000 1017.885000 1.435000 ;
      RECT 1017.605000  1.435000 1019.750000 1.700000 ;
      RECT 1017.615000  0.085000 1017.945000 0.465000 ;
      RECT 1018.000000  1.870000 1018.380000 2.635000 ;
      RECT 1018.055000  1.065000 1020.140000 1.265000 ;
      RECT 1018.165000  0.255000 1018.335000 0.615000 ;
      RECT 1018.165000  0.615000 1019.275000 0.635000 ;
      RECT 1018.555000  0.085000 1018.885000 0.445000 ;
      RECT 1018.600000  1.700000 1018.780000 2.465000 ;
      RECT 1018.960000  1.870000 1019.340000 2.635000 ;
      RECT 1019.105000  0.255000 1019.275000 0.615000 ;
      RECT 1019.445000  0.085000 1019.860000 0.465000 ;
      RECT 1019.560000  1.700000 1019.750000 2.465000 ;
      RECT 1019.920000  0.635000 1021.340000 0.815000 ;
      RECT 1019.920000  0.815000 1020.140000 1.065000 ;
      RECT 1019.920000  1.265000 1020.140000 1.855000 ;
      RECT 1019.920000  1.855000 1023.365000 2.025000 ;
      RECT 1019.920000  2.200000 1020.300000 2.635000 ;
      RECT 1020.100000  0.255000 1022.325000 0.465000 ;
      RECT 1020.310000  0.995000 1020.605000 1.445000 ;
      RECT 1020.310000  1.445000 1022.120000 1.685000 ;
      RECT 1020.520000  2.025000 1020.880000 2.465000 ;
      RECT 1020.775000  1.035000 1021.610000 1.275000 ;
      RECT 1021.055000  2.195000 1021.435000 2.635000 ;
      RECT 1021.605000  2.025000 1021.935000 2.465000 ;
      RECT 1021.790000  1.035000 1022.120000 1.445000 ;
      RECT 1021.995000  0.465000 1022.325000 0.695000 ;
      RECT 1021.995000  0.695000 1024.325000 0.865000 ;
      RECT 1022.115000  2.195000 1022.380000 2.635000 ;
      RECT 1022.345000  1.035000 1022.675000 1.495000 ;
      RECT 1022.345000  1.495000 1024.335000 1.685000 ;
      RECT 1022.500000  0.085000 1022.815000 0.525000 ;
      RECT 1022.860000  1.035000 1023.635000 1.325000 ;
      RECT 1022.985000  0.255000 1023.365000 0.695000 ;
      RECT 1022.985000  2.025000 1023.365000 2.465000 ;
      RECT 1023.585000  0.085000 1023.775000 0.525000 ;
      RECT 1023.820000  1.035000 1024.335000 1.495000 ;
      RECT 1023.945000  0.255000 1024.325000 0.695000 ;
      RECT 1023.945000  1.915000 1024.325000 2.635000 ;
      RECT 1024.505000  0.085000 1024.795000 0.810000 ;
      RECT 1024.505000  1.470000 1024.795000 2.635000 ;
      RECT 1024.965000  0.995000 1025.275000 1.325000 ;
      RECT 1024.975000  0.255000 1025.280000 0.615000 ;
      RECT 1024.975000  0.615000 1026.330000 0.825000 ;
      RECT 1024.975000  1.495000 1025.275000 2.635000 ;
      RECT 1025.445000  0.995000 1025.960000 1.325000 ;
      RECT 1025.445000  1.325000 1025.705000 2.250000 ;
      RECT 1025.450000  0.085000 1025.780000 0.445000 ;
      RECT 1025.875000  1.595000 1026.205000 1.815000 ;
      RECT 1025.875000  1.815000 1027.555000 2.045000 ;
      RECT 1025.875000  2.045000 1026.205000 2.445000 ;
      RECT 1025.950000  0.255000 1026.330000 0.615000 ;
      RECT 1026.300000  0.995000 1026.625000 1.345000 ;
      RECT 1026.375000  1.345000 1026.625000 1.615000 ;
      RECT 1026.420000  2.275000 1026.750000 2.635000 ;
      RECT 1026.605000  0.255000 1027.555000 0.825000 ;
      RECT 1026.795000  1.020000 1027.150000 1.615000 ;
      RECT 1026.955000  2.045000 1027.555000 2.465000 ;
      RECT 1027.320000  0.825000 1027.555000 1.815000 ;
      RECT 1027.725000  0.085000 1028.015000 0.810000 ;
      RECT 1027.725000  1.470000 1028.015000 2.635000 ;
      RECT 1028.185000  0.995000 1028.475000 1.970000 ;
      RECT 1028.195000  0.255000 1030.465000 0.445000 ;
      RECT 1028.215000  2.175000 1028.475000 2.635000 ;
      RECT 1028.645000  0.670000 1029.025000 1.540000 ;
      RECT 1028.645000  1.540000 1031.505000 1.710000 ;
      RECT 1028.645000  1.710000 1028.955000 2.465000 ;
      RECT 1029.125000  1.915000 1029.505000 2.635000 ;
      RECT 1029.245000  0.445000 1030.465000 0.465000 ;
      RECT 1029.245000  0.465000 1029.435000 0.890000 ;
      RECT 1029.315000  1.075000 1030.310000 1.365000 ;
      RECT 1029.605000  0.635000 1032.395000 0.845000 ;
      RECT 1029.725000  1.710000 1029.915000 2.465000 ;
      RECT 1030.085000  1.915000 1030.465000 2.635000 ;
      RECT 1030.695000  0.085000 1031.025000 0.445000 ;
      RECT 1030.695000  2.100000 1030.955000 2.295000 ;
      RECT 1030.695000  2.295000 1031.915000 2.465000 ;
      RECT 1030.770000  1.075000 1031.735000 1.355000 ;
      RECT 1031.125000  1.710000 1031.505000 2.125000 ;
      RECT 1031.625000  0.085000 1032.005000 0.445000 ;
      RECT 1031.725000  1.525000 1032.945000 1.695000 ;
      RECT 1031.725000  1.695000 1031.915000 2.295000 ;
      RECT 1031.905000  1.075000 1033.015000 1.295000 ;
      RECT 1032.085000  1.865000 1032.465000 2.635000 ;
      RECT 1032.205000  0.515000 1032.395000 0.635000 ;
      RECT 1032.565000  0.085000 1032.970000 0.445000 ;
      RECT 1032.565000  0.765000 1033.015000 1.075000 ;
      RECT 1032.685000  1.695000 1032.945000 2.465000 ;
      RECT 1033.245000  0.085000 1033.535000 0.810000 ;
      RECT 1033.245000  1.470000 1033.535000 2.635000 ;
      RECT 1033.710000  1.665000 1034.005000 2.635000 ;
      RECT 1033.775000  0.535000 1033.975000 0.625000 ;
      RECT 1033.775000  0.625000 1037.855000 0.795000 ;
      RECT 1033.775000  0.795000 1037.100000 0.905000 ;
      RECT 1034.020000  1.075000 1035.180000 1.330000 ;
      RECT 1034.145000  0.085000 1034.525000 0.445000 ;
      RECT 1034.225000  1.860000 1034.445000 1.935000 ;
      RECT 1034.225000  1.935000 1035.405000 2.105000 ;
      RECT 1034.225000  2.105000 1034.445000 2.190000 ;
      RECT 1034.625000  2.275000 1035.005000 2.635000 ;
      RECT 1034.635000  1.330000 1035.180000 1.515000 ;
      RECT 1034.635000  1.515000 1037.650000 1.685000 ;
      RECT 1034.745000  0.425000 1034.960000 0.625000 ;
      RECT 1035.155000  0.085000 1035.485000 0.455000 ;
      RECT 1035.225000  2.105000 1035.405000 2.275000 ;
      RECT 1035.225000  2.275000 1037.405000 2.465000 ;
      RECT 1035.475000  1.075000 1037.150000 1.345000 ;
      RECT 1035.575000  1.855000 1042.100000 2.025000 ;
      RECT 1035.575000  2.025000 1037.440000 2.105000 ;
      RECT 1036.065000  0.085000 1036.445000 0.445000 ;
      RECT 1037.025000  0.085000 1037.405000 0.445000 ;
      RECT 1037.320000  0.995000 1037.650000 1.515000 ;
      RECT 1037.625000  0.255000 1039.090000 0.455000 ;
      RECT 1037.625000  0.455000 1037.855000 0.625000 ;
      RECT 1037.635000  2.195000 1037.905000 2.635000 ;
      RECT 1037.820000  0.995000 1039.145000 1.410000 ;
      RECT 1038.025000  0.635000 1040.490000 0.815000 ;
      RECT 1038.115000  2.025000 1042.100000 2.105000 ;
      RECT 1038.330000  1.410000 1039.145000 1.515000 ;
      RECT 1038.330000  1.515000 1041.420000 1.685000 ;
      RECT 1038.505000  2.275000 1038.885000 2.635000 ;
      RECT 1039.450000  0.270000 1041.105000 0.450000 ;
      RECT 1039.450000  2.275000 1039.830000 2.635000 ;
      RECT 1039.590000  1.075000 1040.760000 1.345000 ;
      RECT 1040.390000  2.275000 1040.775000 2.635000 ;
      RECT 1040.885000  0.450000 1041.105000 0.655000 ;
      RECT 1040.885000  0.655000 1041.780000 0.825000 ;
      RECT 1041.200000  0.995000 1041.420000 1.515000 ;
      RECT 1041.350000  0.310000 1042.110000 0.480000 ;
      RECT 1041.600000  0.825000 1041.780000 1.340000 ;
      RECT 1041.600000  1.340000 1042.100000 1.855000 ;
      RECT 1041.775000  2.275000 1042.105000 2.635000 ;
      RECT 1041.940000  0.480000 1042.110000 0.595000 ;
      RECT 1042.445000  0.085000 1042.735000 0.810000 ;
      RECT 1042.445000  1.470000 1042.735000 2.635000 ;
      RECT 1042.905000  0.255000 1043.245000 1.030000 ;
      RECT 1042.905000  1.030000 1043.185000 2.465000 ;
      RECT 1043.355000  1.860000 1044.085000 2.635000 ;
      RECT 1043.420000  0.715000 1044.205000 0.905000 ;
      RECT 1043.420000  0.905000 1043.705000 1.475000 ;
      RECT 1043.420000  1.475000 1044.630000 1.690000 ;
      RECT 1043.435000  0.085000 1043.605000 0.545000 ;
      RECT 1043.845000  0.255000 1044.205000 0.715000 ;
      RECT 1043.875000  1.075000 1044.375000 1.305000 ;
      RECT 1044.300000  1.690000 1044.630000 2.465000 ;
      RECT 1044.375000  0.555000 1044.585000 0.715000 ;
      RECT 1044.375000  0.715000 1045.530000 0.905000 ;
      RECT 1044.545000  1.075000 1044.975000 1.275000 ;
      RECT 1044.800000  0.085000 1044.970000 0.545000 ;
      RECT 1044.805000  1.275000 1044.975000 2.390000 ;
      RECT 1045.145000  1.075000 1045.495000 1.615000 ;
      RECT 1045.200000  0.255000 1045.530000 0.715000 ;
      RECT 1045.200000  1.915000 1045.920000 2.635000 ;
      RECT 1046.125000  0.085000 1046.415000 0.810000 ;
      RECT 1046.125000  1.470000 1046.415000 2.635000 ;
      RECT 1046.590000  1.635000 1046.845000 2.635000 ;
      RECT 1046.605000  0.085000 1046.845000 0.885000 ;
      RECT 1047.030000  0.255000 1047.325000 2.465000 ;
      RECT 1047.495000  0.085000 1047.875000 0.465000 ;
      RECT 1047.495000  0.635000 1048.395000 0.840000 ;
      RECT 1047.495000  0.840000 1047.855000 1.330000 ;
      RECT 1047.495000  2.185000 1048.395000 2.635000 ;
      RECT 1047.685000  1.330000 1047.855000 1.785000 ;
      RECT 1047.685000  1.785000 1048.875000 2.005000 ;
      RECT 1048.025000  1.010000 1048.455000 1.615000 ;
      RECT 1048.065000  0.255000 1048.395000 0.635000 ;
      RECT 1048.615000  0.465000 1048.825000 0.635000 ;
      RECT 1048.615000  0.635000 1050.030000 0.825000 ;
      RECT 1048.615000  2.005000 1048.875000 2.465000 ;
      RECT 1048.820000  1.025000 1049.575000 1.400000 ;
      RECT 1048.995000  0.085000 1049.535000 0.465000 ;
      RECT 1049.300000  1.400000 1049.575000 1.985000 ;
      RECT 1049.745000  1.650000 1050.030000 2.635000 ;
      RECT 1049.755000  0.495000 1050.030000 0.635000 ;
      RECT 1049.775000  0.995000 1050.035000 1.450000 ;
      RECT 1050.265000  0.085000 1050.555000 0.810000 ;
      RECT 1050.265000  1.470000 1050.555000 2.635000 ;
      RECT 1050.730000  0.635000 1052.505000 0.805000 ;
      RECT 1050.730000  0.805000 1050.990000 1.530000 ;
      RECT 1050.730000  1.530000 1052.795000 1.700000 ;
      RECT 1050.735000  0.085000 1051.065000 0.465000 ;
      RECT 1051.055000  1.870000 1051.435000 2.635000 ;
      RECT 1051.160000  0.995000 1053.205000 1.335000 ;
      RECT 1051.285000  0.615000 1052.505000 0.635000 ;
      RECT 1051.655000  1.700000 1051.845000 2.465000 ;
      RECT 1051.695000  0.085000 1052.025000 0.445000 ;
      RECT 1052.015000  1.870000 1052.395000 2.635000 ;
      RECT 1052.615000  1.700000 1052.795000 2.465000 ;
      RECT 1052.655000  0.085000 1052.985000 0.465000 ;
      RECT 1052.955000  0.655000 1054.025000 0.870000 ;
      RECT 1052.955000  0.870000 1053.205000 0.995000 ;
      RECT 1052.965000  1.335000 1053.205000 1.830000 ;
      RECT 1052.965000  1.830000 1053.835000 1.875000 ;
      RECT 1052.965000  1.875000 1055.515000 2.085000 ;
      RECT 1052.975000  2.255000 1053.375000 2.635000 ;
      RECT 1053.225000  0.255000 1054.525000 0.485000 ;
      RECT 1053.375000  1.075000 1054.125000 1.615000 ;
      RECT 1053.595000  2.085000 1055.515000 2.105000 ;
      RECT 1053.595000  2.105000 1053.835000 2.465000 ;
      RECT 1054.155000  2.275000 1054.485000 2.635000 ;
      RECT 1054.195000  0.485000 1054.525000 0.615000 ;
      RECT 1054.195000  0.615000 1056.475000 0.785000 ;
      RECT 1054.400000  0.990000 1054.755000 1.495000 ;
      RECT 1054.400000  1.495000 1056.520000 1.705000 ;
      RECT 1054.695000  0.085000 1055.035000 0.445000 ;
      RECT 1055.060000  0.995000 1055.710000 1.325000 ;
      RECT 1055.135000  2.105000 1055.515000 2.445000 ;
      RECT 1055.615000  0.085000 1055.995000 0.445000 ;
      RECT 1056.050000  0.995000 1056.520000 1.495000 ;
      RECT 1056.095000  1.935000 1056.505000 2.635000 ;
      RECT 1056.705000  0.085000 1056.995000 0.810000 ;
      RECT 1056.705000  1.470000 1056.995000 2.635000 ;
      RECT 1057.170000  0.265000 1057.460000 0.615000 ;
      RECT 1057.170000  0.615000 1058.485000 0.785000 ;
      RECT 1057.170000  1.495000 1057.490000 2.635000 ;
      RECT 1057.225000  0.995000 1057.490000 1.325000 ;
      RECT 1057.660000  0.995000 1058.155000 1.325000 ;
      RECT 1057.660000  1.325000 1057.915000 2.375000 ;
      RECT 1057.705000  0.085000 1058.085000 0.445000 ;
      RECT 1058.085000  1.505000 1058.495000 2.465000 ;
      RECT 1058.255000  0.310000 1058.485000 0.615000 ;
      RECT 1058.325000  0.955000 1059.190000 1.125000 ;
      RECT 1058.325000  1.125000 1058.495000 1.505000 ;
      RECT 1058.725000  0.275000 1059.190000 0.955000 ;
      RECT 1058.725000  1.835000 1059.190000 2.635000 ;
      RECT 1058.735000  1.295000 1059.295000 1.655000 ;
      RECT 1059.465000  0.085000 1059.755000 0.810000 ;
      RECT 1059.465000  1.470000 1059.755000 2.635000 ;
      RECT 1059.945000  0.255000 1060.275000 0.715000 ;
      RECT 1059.945000  0.715000 1062.305000 0.885000 ;
      RECT 1059.945000  1.785000 1060.275000 2.635000 ;
      RECT 1059.960000  1.055000 1060.290000 1.445000 ;
      RECT 1059.960000  1.445000 1062.135000 1.615000 ;
      RECT 1060.495000  1.785000 1060.715000 2.295000 ;
      RECT 1060.495000  2.295000 1061.705000 2.465000 ;
      RECT 1060.505000  0.085000 1060.675000 0.545000 ;
      RECT 1060.510000  1.075000 1061.410000 1.275000 ;
      RECT 1060.855000  0.255000 1061.235000 0.715000 ;
      RECT 1060.935000  1.785000 1062.950000 1.965000 ;
      RECT 1060.935000  1.965000 1061.235000 2.125000 ;
      RECT 1061.515000  0.085000 1061.685000 0.545000 ;
      RECT 1061.515000  2.135000 1061.705000 2.295000 ;
      RECT 1061.590000  1.075000 1062.135000 1.445000 ;
      RECT 1061.900000  2.175000 1062.280000 2.635000 ;
      RECT 1061.975000  0.255000 1063.370000 0.425000 ;
      RECT 1061.975000  0.425000 1062.305000 0.715000 ;
      RECT 1062.535000  0.595000 1062.950000 1.785000 ;
      RECT 1062.535000  1.965000 1062.950000 2.465000 ;
      RECT 1063.120000  0.425000 1063.370000 0.595000 ;
      RECT 1063.120000  0.765000 1063.410000 1.400000 ;
      RECT 1063.120000  1.570000 1063.370000 2.635000 ;
      RECT 1063.605000  0.085000 1063.895000 0.810000 ;
      RECT 1063.605000  1.470000 1063.895000 2.635000 ;
      RECT 1064.100000  0.615000 1068.240000 0.820000 ;
      RECT 1064.100000  1.820000 1064.385000 2.635000 ;
      RECT 1064.105000  1.015000 1065.605000 1.320000 ;
      RECT 1064.530000  0.085000 1064.910000 0.445000 ;
      RECT 1064.605000  1.320000 1065.605000 1.515000 ;
      RECT 1064.605000  1.515000 1068.075000 1.685000 ;
      RECT 1064.605000  1.915000 1065.800000 2.085000 ;
      RECT 1064.605000  2.085000 1064.840000 2.465000 ;
      RECT 1065.010000  2.255000 1065.390000 2.635000 ;
      RECT 1065.490000  0.085000 1065.870000 0.445000 ;
      RECT 1065.610000  2.085000 1065.800000 2.275000 ;
      RECT 1065.610000  2.275000 1067.790000 2.465000 ;
      RECT 1065.970000  1.855000 1069.680000 2.025000 ;
      RECT 1066.165000  1.070000 1067.605000 1.345000 ;
      RECT 1066.450000  0.085000 1066.830000 0.445000 ;
      RECT 1067.410000  0.085000 1067.790000 0.445000 ;
      RECT 1067.775000  0.990000 1068.075000 1.515000 ;
      RECT 1068.010000  0.255000 1070.230000 0.445000 ;
      RECT 1068.010000  0.445000 1068.240000 0.615000 ;
      RECT 1068.010000  2.195000 1068.290000 2.635000 ;
      RECT 1068.285000  1.015000 1069.580000 1.275000 ;
      RECT 1068.315000  1.445000 1070.310000 1.700000 ;
      RECT 1068.315000  1.700000 1069.680000 1.855000 ;
      RECT 1068.410000  0.615000 1070.310000 0.845000 ;
      RECT 1068.510000  2.025000 1069.680000 2.085000 ;
      RECT 1068.510000  2.085000 1068.720000 2.465000 ;
      RECT 1068.890000  2.255000 1069.270000 2.635000 ;
      RECT 1069.490000  2.085000 1069.680000 2.465000 ;
      RECT 1069.850000  1.880000 1070.230000 2.635000 ;
      RECT 1069.900000  0.845000 1070.310000 1.445000 ;
      RECT 1070.505000  0.085000 1070.795000 0.810000 ;
      RECT 1070.505000  1.470000 1070.795000 2.635000 ;
      RECT 1070.965000  0.450000 1071.325000 0.825000 ;
      RECT 1070.965000  0.825000 1071.220000 1.480000 ;
      RECT 1070.965000  1.480000 1071.305000 2.465000 ;
      RECT 1071.390000  0.995000 1071.740000 1.325000 ;
      RECT 1071.475000  2.205000 1071.885000 2.635000 ;
      RECT 1071.525000  1.325000 1071.740000 1.865000 ;
      RECT 1071.525000  1.865000 1073.465000 2.035000 ;
      RECT 1071.555000  0.085000 1071.725000 0.825000 ;
      RECT 1071.910000  0.995000 1072.260000 1.325000 ;
      RECT 1071.955000  1.525000 1072.600000 1.695000 ;
      RECT 1072.090000  0.450000 1072.260000 0.655000 ;
      RECT 1072.090000  0.655000 1072.600000 0.825000 ;
      RECT 1072.430000  0.825000 1072.600000 1.525000 ;
      RECT 1072.650000  2.215000 1072.980000 2.635000 ;
      RECT 1072.770000  0.255000 1072.940000 1.455000 ;
      RECT 1072.770000  1.455000 1073.465000 1.865000 ;
      RECT 1073.110000  1.075000 1073.730000 1.285000 ;
      RECT 1073.160000  0.255000 1073.490000 0.735000 ;
      RECT 1073.160000  0.735000 1074.445000 0.905000 ;
      RECT 1073.160000  2.035000 1073.465000 2.465000 ;
      RECT 1073.710000  0.085000 1073.880000 0.555000 ;
      RECT 1073.900000  1.075000 1074.450000 1.285000 ;
      RECT 1074.050000  1.535000 1074.430000 2.635000 ;
      RECT 1074.115000  0.270000 1074.445000 0.735000 ;
      RECT 1074.645000  0.085000 1074.935000 0.810000 ;
      RECT 1074.645000  1.470000 1074.935000 2.635000 ;
      RECT 1075.105000  0.430000 1075.365000 0.825000 ;
      RECT 1075.105000  0.825000 1075.275000 1.495000 ;
      RECT 1075.105000  1.495000 1075.415000 1.865000 ;
      RECT 1075.105000  1.865000 1077.105000 2.035000 ;
      RECT 1075.445000  0.995000 1075.845000 1.325000 ;
      RECT 1075.540000  2.205000 1075.980000 2.635000 ;
      RECT 1075.625000  1.325000 1075.845000 1.695000 ;
      RECT 1075.665000  0.085000 1075.845000 0.825000 ;
      RECT 1076.015000  0.295000 1076.400000 0.465000 ;
      RECT 1076.015000  0.465000 1076.255000 1.495000 ;
      RECT 1076.015000  1.495000 1076.475000 1.695000 ;
      RECT 1076.425000  0.655000 1077.490000 0.825000 ;
      RECT 1076.425000  0.825000 1076.595000 1.325000 ;
      RECT 1076.540000  2.205000 1077.400000 2.635000 ;
      RECT 1076.580000  0.085000 1076.945000 0.465000 ;
      RECT 1076.935000  0.995000 1077.105000 1.865000 ;
      RECT 1077.160000  0.255000 1077.490000 0.655000 ;
      RECT 1077.275000  0.825000 1077.490000 1.455000 ;
      RECT 1077.275000  1.455000 1077.945000 2.035000 ;
      RECT 1077.620000  2.035000 1077.945000 2.465000 ;
      RECT 1077.665000  1.075000 1078.200000 1.285000 ;
      RECT 1077.715000  0.365000 1077.965000 0.735000 ;
      RECT 1077.715000  0.735000 1078.910000 0.905000 ;
      RECT 1078.185000  0.085000 1078.355000 0.555000 ;
      RECT 1078.370000  1.075000 1078.915000 1.625000 ;
      RECT 1078.470000  1.875000 1078.850000 2.635000 ;
      RECT 1078.575000  0.270000 1078.910000 0.735000 ;
      RECT 1079.245000  0.085000 1079.535000 0.810000 ;
      RECT 1079.245000  1.470000 1079.535000 2.635000 ;
      RECT 1079.705000  0.265000 1080.165000 0.855000 ;
      RECT 1079.705000  0.855000 1079.875000 1.455000 ;
      RECT 1079.705000  1.455000 1080.055000 1.875000 ;
      RECT 1079.705000  1.875000 1082.435000 2.045000 ;
      RECT 1079.705000  2.045000 1080.055000 2.465000 ;
      RECT 1080.045000  1.075000 1080.555000 1.285000 ;
      RECT 1080.225000  1.285000 1080.555000 1.705000 ;
      RECT 1080.255000  2.215000 1080.635000 2.635000 ;
      RECT 1080.385000  0.085000 1080.555000 0.905000 ;
      RECT 1080.775000  0.255000 1081.105000 0.725000 ;
      RECT 1080.775000  0.725000 1081.995000 0.910000 ;
      RECT 1080.775000  0.910000 1081.325000 1.445000 ;
      RECT 1080.775000  1.445000 1082.045000 1.705000 ;
      RECT 1081.195000  2.215000 1081.575000 2.635000 ;
      RECT 1081.325000  0.085000 1081.495000 0.555000 ;
      RECT 1081.495000  1.080000 1082.435000 1.250000 ;
      RECT 1081.665000  0.255000 1081.995000 0.725000 ;
      RECT 1082.135000  2.215000 1082.515000 2.635000 ;
      RECT 1082.185000  0.085000 1082.515000 0.475000 ;
      RECT 1082.265000  0.645000 1083.555000 0.895000 ;
      RECT 1082.265000  0.895000 1082.435000 1.080000 ;
      RECT 1082.265000  1.445000 1082.825000 1.615000 ;
      RECT 1082.265000  1.615000 1082.435000 1.875000 ;
      RECT 1082.605000  1.075000 1083.055000 1.245000 ;
      RECT 1082.605000  1.245000 1082.825000 1.445000 ;
      RECT 1082.725000  0.255000 1084.025000 0.475000 ;
      RECT 1082.735000  1.795000 1084.450000 1.965000 ;
      RECT 1082.735000  1.965000 1082.905000 2.465000 ;
      RECT 1083.170000  2.135000 1083.420000 2.635000 ;
      RECT 1083.365000  0.895000 1083.555000 1.795000 ;
      RECT 1083.655000  2.135000 1083.945000 2.295000 ;
      RECT 1083.655000  2.295000 1084.885000 2.465000 ;
      RECT 1083.775000  0.475000 1084.025000 0.725000 ;
      RECT 1083.775000  0.725000 1085.930000 0.905000 ;
      RECT 1083.800000  1.075000 1084.940000 1.275000 ;
      RECT 1084.205000  1.445000 1084.450000 1.795000 ;
      RECT 1084.205000  1.965000 1084.450000 2.125000 ;
      RECT 1084.245000  0.085000 1084.415000 0.555000 ;
      RECT 1084.585000  0.255000 1084.965000 0.725000 ;
      RECT 1084.715000  1.455000 1085.930000 1.665000 ;
      RECT 1084.715000  1.665000 1084.885000 2.295000 ;
      RECT 1085.055000  1.835000 1085.435000 2.635000 ;
      RECT 1085.160000  1.075000 1085.975000 1.275000 ;
      RECT 1085.185000  0.085000 1085.355000 0.555000 ;
      RECT 1085.525000  0.265000 1085.930000 0.725000 ;
      RECT 1085.655000  1.665000 1085.930000 2.465000 ;
      RECT 1086.145000  0.085000 1086.435000 0.810000 ;
      RECT 1086.145000  1.470000 1086.435000 2.635000 ;
      RECT 1086.605000  0.085000 1086.880000 0.825000 ;
      RECT 1086.605000  0.995000 1087.055000 1.345000 ;
      RECT 1086.605000  1.345000 1086.875000 2.445000 ;
      RECT 1087.045000  1.535000 1087.585000 1.705000 ;
      RECT 1087.045000  1.705000 1087.370000 2.210000 ;
      RECT 1087.195000  0.495000 1087.460000 0.825000 ;
      RECT 1087.290000  0.825000 1087.460000 0.995000 ;
      RECT 1087.290000  0.995000 1087.585000 1.535000 ;
      RECT 1087.590000  1.875000 1087.920000 2.635000 ;
      RECT 1087.755000  0.255000 1087.975000 1.445000 ;
      RECT 1087.755000  1.445000 1088.675000 1.625000 ;
      RECT 1088.155000  1.625000 1088.675000 2.465000 ;
      RECT 1088.160000  0.255000 1088.490000 0.735000 ;
      RECT 1088.160000  0.735000 1089.435000 0.905000 ;
      RECT 1088.195000  1.075000 1088.715000 1.275000 ;
      RECT 1088.715000  0.085000 1088.885000 0.555000 ;
      RECT 1088.885000  1.075000 1089.445000 1.285000 ;
      RECT 1088.990000  1.535000 1089.580000 2.635000 ;
      RECT 1089.055000  0.270000 1089.435000 0.735000 ;
      RECT 1089.825000  0.085000 1090.115000 0.810000 ;
      RECT 1089.825000  1.470000 1090.115000 2.635000 ;
      RECT 1090.285000  0.995000 1090.680000 1.325000 ;
      RECT 1090.380000  0.085000 1090.550000 0.825000 ;
      RECT 1090.380000  1.495000 1091.115000 1.665000 ;
      RECT 1090.380000  1.665000 1090.550000 1.915000 ;
      RECT 1090.835000  1.875000 1091.165000 2.635000 ;
      RECT 1090.850000  0.445000 1091.020000 1.075000 ;
      RECT 1090.850000  1.075000 1091.540000 1.245000 ;
      RECT 1090.850000  1.245000 1091.115000 1.495000 ;
      RECT 1091.260000  0.255000 1092.675000 0.475000 ;
      RECT 1091.260000  0.475000 1091.540000 0.905000 ;
      RECT 1091.385000  1.445000 1093.100000 1.615000 ;
      RECT 1091.385000  1.615000 1091.555000 2.465000 ;
      RECT 1091.710000  0.645000 1092.205000 1.445000 ;
      RECT 1091.820000  1.795000 1092.070000 2.635000 ;
      RECT 1092.305000  1.795000 1092.635000 2.295000 ;
      RECT 1092.305000  2.295000 1093.535000 2.465000 ;
      RECT 1092.375000  1.075000 1093.590000 1.275000 ;
      RECT 1092.425000  0.475000 1092.675000 0.725000 ;
      RECT 1092.425000  0.725000 1094.580000 0.905000 ;
      RECT 1092.855000  1.615000 1093.100000 2.125000 ;
      RECT 1092.895000  0.085000 1093.065000 0.555000 ;
      RECT 1093.235000  0.255000 1093.615000 0.725000 ;
      RECT 1093.365000  1.455000 1094.580000 1.665000 ;
      RECT 1093.365000  1.665000 1093.535000 2.295000 ;
      RECT 1093.705000  1.835000 1094.085000 2.635000 ;
      RECT 1093.810000  1.075000 1094.655000 1.275000 ;
      RECT 1093.835000  0.085000 1094.005000 0.555000 ;
      RECT 1094.175000  0.265000 1094.580000 0.725000 ;
      RECT 1094.305000  1.665000 1094.580000 2.465000 ;
      RECT 1094.885000  0.085000 1095.175000 0.810000 ;
      RECT 1094.885000  1.470000 1095.175000 2.635000 ;
      RECT 1095.345000  1.075000 1095.770000 1.285000 ;
      RECT 1095.405000  1.455000 1096.110000 1.625000 ;
      RECT 1095.405000  1.625000 1095.735000 2.435000 ;
      RECT 1095.485000  0.085000 1095.655000 0.895000 ;
      RECT 1095.825000  0.290000 1096.205000 0.895000 ;
      RECT 1095.940000  0.895000 1096.205000 1.075000 ;
      RECT 1095.940000  1.075000 1097.785000 1.285000 ;
      RECT 1095.940000  1.285000 1096.110000 1.455000 ;
      RECT 1095.955000  1.795000 1096.125000 2.635000 ;
      RECT 1096.295000  1.455000 1100.025000 1.625000 ;
      RECT 1096.295000  1.625000 1096.635000 2.465000 ;
      RECT 1096.440000  0.305000 1098.655000 0.475000 ;
      RECT 1096.780000  0.645000 1098.185000 0.815000 ;
      RECT 1096.855000  1.795000 1097.105000 2.635000 ;
      RECT 1097.325000  1.625000 1097.575000 2.465000 ;
      RECT 1097.795000  1.795000 1098.045000 2.635000 ;
      RECT 1097.955000  0.815000 1098.185000 1.075000 ;
      RECT 1097.955000  1.075000 1098.455000 1.445000 ;
      RECT 1097.955000  1.445000 1100.025000 1.455000 ;
      RECT 1098.285000  1.795000 1098.615000 2.295000 ;
      RECT 1098.285000  2.295000 1100.495000 2.465000 ;
      RECT 1098.405000  0.475000 1098.655000 0.725000 ;
      RECT 1098.405000  0.725000 1102.415000 0.905000 ;
      RECT 1098.625000  1.075000 1100.235000 1.275000 ;
      RECT 1098.835000  1.625000 1099.085000 2.125000 ;
      RECT 1098.875000  0.085000 1099.045000 0.555000 ;
      RECT 1099.215000  0.255000 1099.595000 0.725000 ;
      RECT 1099.305000  1.795000 1099.555000 2.295000 ;
      RECT 1099.775000  1.625000 1100.025000 2.125000 ;
      RECT 1099.815000  0.085000 1099.985000 0.555000 ;
      RECT 1100.155000  0.255000 1100.535000 0.725000 ;
      RECT 1100.245000  1.455000 1102.375000 1.625000 ;
      RECT 1100.245000  1.625000 1100.495000 2.295000 ;
      RECT 1100.405000  1.075000 1102.510000 1.285000 ;
      RECT 1100.715000  1.795000 1100.965000 2.635000 ;
      RECT 1100.755000  0.085000 1100.925000 0.555000 ;
      RECT 1101.095000  0.255000 1101.475000 0.725000 ;
      RECT 1101.185000  1.625000 1101.435000 2.465000 ;
      RECT 1101.655000  1.795000 1101.905000 2.635000 ;
      RECT 1101.695000  0.085000 1101.865000 0.555000 ;
      RECT 1102.035000  0.255000 1102.415000 0.725000 ;
      RECT 1102.125000  1.625000 1102.375000 2.465000 ;
      RECT 1102.705000  0.085000 1102.995000 0.810000 ;
      RECT 1102.705000  1.470000 1102.995000 2.635000 ;
      RECT 1103.165000  0.995000 1103.495000 1.285000 ;
      RECT 1103.165000  1.455000 1103.835000 1.495000 ;
      RECT 1103.165000  1.495000 1104.315000 1.720000 ;
      RECT 1103.165000  1.720000 1103.445000 2.465000 ;
      RECT 1103.250000  0.255000 1103.580000 0.645000 ;
      RECT 1103.250000  0.645000 1103.835000 0.825000 ;
      RECT 1103.640000  2.085000 1103.940000 2.635000 ;
      RECT 1103.665000  0.825000 1103.835000 1.455000 ;
      RECT 1103.780000  0.305000 1104.985000 0.475000 ;
      RECT 1104.005000  0.985000 1104.315000 1.325000 ;
      RECT 1104.110000  1.720000 1104.315000 1.875000 ;
      RECT 1104.110000  1.875000 1105.825000 2.045000 ;
      RECT 1104.115000  0.645000 1106.015000 0.815000 ;
      RECT 1104.485000  0.985000 1104.870000 1.705000 ;
      RECT 1104.580000  2.045000 1105.435000 2.465000 ;
      RECT 1105.060000  0.985000 1105.695000 1.255000 ;
      RECT 1105.060000  1.255000 1105.395000 1.705000 ;
      RECT 1105.165000  0.085000 1105.505000 0.475000 ;
      RECT 1105.655000  1.455000 1106.625000 1.625000 ;
      RECT 1105.655000  1.625000 1105.825000 1.875000 ;
      RECT 1105.685000  0.270000 1106.015000 0.645000 ;
      RECT 1105.895000  1.075000 1106.225000 1.285000 ;
      RECT 1105.995000  1.795000 1106.375000 2.635000 ;
      RECT 1106.185000  0.085000 1106.355000 0.640000 ;
      RECT 1106.455000  0.995000 1106.625000 1.455000 ;
      RECT 1106.525000  0.265000 1107.110000 0.825000 ;
      RECT 1106.545000  1.875000 1107.110000 2.465000 ;
      RECT 1106.795000  0.825000 1107.110000 1.875000 ;
      RECT 1107.305000  0.085000 1107.595000 0.810000 ;
      RECT 1107.305000  1.470000 1107.595000 2.635000 ;
      RECT 1107.765000  0.975000 1108.025000 1.325000 ;
      RECT 1107.850000  0.255000 1108.180000 0.635000 ;
      RECT 1107.850000  0.635000 1108.445000 0.805000 ;
      RECT 1107.930000  1.495000 1109.030000 1.670000 ;
      RECT 1107.930000  1.670000 1108.260000 2.465000 ;
      RECT 1108.225000  0.805000 1108.445000 1.445000 ;
      RECT 1108.225000  1.445000 1109.030000 1.495000 ;
      RECT 1108.350000  0.295000 1109.685000 0.465000 ;
      RECT 1108.480000  1.850000 1108.690000 2.635000 ;
      RECT 1108.615000  1.075000 1109.010000 1.275000 ;
      RECT 1108.815000  0.645000 1109.250000 0.735000 ;
      RECT 1108.815000  0.735000 1110.665000 0.905000 ;
      RECT 1108.860000  1.670000 1109.030000 1.875000 ;
      RECT 1108.860000  1.875000 1110.645000 2.045000 ;
      RECT 1109.200000  1.075000 1109.585000 1.705000 ;
      RECT 1109.380000  2.045000 1110.135000 2.465000 ;
      RECT 1109.915000  1.075000 1110.295000 1.705000 ;
      RECT 1109.945000  0.085000 1110.115000 0.555000 ;
      RECT 1110.285000  0.270000 1110.665000 0.735000 ;
      RECT 1110.475000  1.455000 1111.395000 1.625000 ;
      RECT 1110.475000  1.625000 1110.645000 1.875000 ;
      RECT 1110.515000  1.075000 1111.005000 1.285000 ;
      RECT 1110.825000  1.795000 1111.055000 2.635000 ;
      RECT 1110.885000  0.085000 1111.055000 0.905000 ;
      RECT 1111.175000  1.075000 1111.555000 1.285000 ;
      RECT 1111.175000  1.285000 1111.395000 1.455000 ;
      RECT 1111.225000  0.265000 1111.605000 0.735000 ;
      RECT 1111.225000  0.735000 1112.170000 0.905000 ;
      RECT 1111.225000  1.875000 1112.170000 2.045000 ;
      RECT 1111.225000  2.045000 1111.525000 2.465000 ;
      RECT 1111.695000  2.215000 1112.085000 2.635000 ;
      RECT 1111.825000  0.085000 1111.995000 0.565000 ;
      RECT 1111.860000  0.905000 1112.170000 1.875000 ;
      RECT 1112.365000  0.085000 1112.655000 0.810000 ;
      RECT 1112.365000  1.470000 1112.655000 2.635000 ;
      RECT 1112.825000  0.255000 1115.995000 0.475000 ;
      RECT 1112.825000  0.475000 1113.085000 0.895000 ;
      RECT 1112.830000  1.075000 1113.180000 1.275000 ;
      RECT 1112.885000  1.455000 1113.135000 2.635000 ;
      RECT 1113.255000  0.645000 1113.635000 0.865000 ;
      RECT 1113.355000  0.865000 1113.635000 1.785000 ;
      RECT 1113.355000  1.785000 1118.385000 1.955000 ;
      RECT 1113.355000  1.955000 1113.605000 2.465000 ;
      RECT 1113.805000  1.075000 1114.470000 1.445000 ;
      RECT 1113.805000  1.445000 1115.785000 1.615000 ;
      RECT 1113.825000  2.125000 1114.075000 2.635000 ;
      RECT 1113.855000  0.475000 1114.025000 0.905000 ;
      RECT 1114.195000  0.645000 1116.975000 0.725000 ;
      RECT 1114.195000  0.725000 1117.915000 0.905000 ;
      RECT 1114.295000  2.125000 1114.545000 2.295000 ;
      RECT 1114.295000  2.295000 1115.485000 2.465000 ;
      RECT 1114.690000  1.075000 1115.235000 1.275000 ;
      RECT 1115.235000  2.125000 1115.485000 2.295000 ;
      RECT 1115.405000  1.075000 1115.785000 1.445000 ;
      RECT 1115.705000  2.125000 1116.465000 2.635000 ;
      RECT 1116.045000  1.075000 1116.695000 1.445000 ;
      RECT 1116.045000  1.445000 1117.965000 1.615000 ;
      RECT 1116.175000  0.085000 1116.505000 0.465000 ;
      RECT 1116.685000  2.125000 1116.935000 2.295000 ;
      RECT 1116.685000  2.295000 1117.875000 2.465000 ;
      RECT 1116.725000  0.255000 1116.975000 0.645000 ;
      RECT 1116.865000  1.075000 1117.495000 1.275000 ;
      RECT 1117.195000  0.085000 1117.365000 0.555000 ;
      RECT 1117.535000  0.255000 1117.915000 0.725000 ;
      RECT 1117.625000  2.125000 1117.875000 2.295000 ;
      RECT 1117.715000  1.075000 1118.275000 1.275000 ;
      RECT 1117.715000  1.275000 1117.965000 1.445000 ;
      RECT 1118.095000  2.125000 1118.345000 2.635000 ;
      RECT 1118.135000  0.085000 1118.305000 0.905000 ;
      RECT 1118.215000  1.445000 1118.665000 1.615000 ;
      RECT 1118.215000  1.615000 1118.385000 1.785000 ;
      RECT 1118.445000  1.075000 1119.795000 1.275000 ;
      RECT 1118.445000  1.275000 1118.665000 1.445000 ;
      RECT 1118.475000  0.255000 1118.855000 0.725000 ;
      RECT 1118.475000  0.725000 1119.795000 0.735000 ;
      RECT 1118.475000  0.735000 1120.450000 0.905000 ;
      RECT 1118.605000  1.785000 1119.240000 1.955000 ;
      RECT 1118.605000  1.955000 1118.815000 2.465000 ;
      RECT 1119.035000  2.125000 1119.285000 2.635000 ;
      RECT 1119.070000  1.445000 1120.450000 1.615000 ;
      RECT 1119.070000  1.615000 1119.240000 1.785000 ;
      RECT 1119.075000  0.085000 1119.245000 0.555000 ;
      RECT 1119.415000  0.255000 1119.795000 0.725000 ;
      RECT 1119.505000  1.615000 1119.755000 2.465000 ;
      RECT 1119.975000  1.795000 1120.225000 2.635000 ;
      RECT 1120.015000  0.085000 1120.270000 0.565000 ;
      RECT 1120.105000  0.905000 1120.450000 1.445000 ;
      RECT 1120.645000  0.085000 1120.935000 0.810000 ;
      RECT 1120.645000  1.470000 1120.935000 2.635000 ;
      RECT 1121.105000  0.365000 1121.365000 0.645000 ;
      RECT 1121.105000  0.645000 1121.865000 0.825000 ;
      RECT 1121.105000  0.995000 1121.485000 1.325000 ;
      RECT 1121.105000  1.495000 1123.485000 1.705000 ;
      RECT 1121.105000  1.705000 1121.385000 2.465000 ;
      RECT 1121.535000  0.305000 1123.085000 0.475000 ;
      RECT 1121.620000  1.875000 1122.600000 2.635000 ;
      RECT 1121.695000  0.825000 1121.865000 1.495000 ;
      RECT 1122.035000  0.995000 1122.615000 1.325000 ;
      RECT 1122.270000  0.645000 1123.580000 0.695000 ;
      RECT 1122.270000  0.695000 1124.595000 0.825000 ;
      RECT 1122.835000  0.995000 1123.345000 1.325000 ;
      RECT 1122.920000  1.705000 1123.485000 2.180000 ;
      RECT 1122.920000  2.180000 1123.525000 2.465000 ;
      RECT 1123.305000  0.280000 1123.580000 0.645000 ;
      RECT 1123.465000  0.825000 1124.595000 0.865000 ;
      RECT 1123.525000  1.075000 1123.915000 1.245000 ;
      RECT 1123.655000  1.245000 1123.915000 1.445000 ;
      RECT 1123.655000  1.445000 1124.145000 1.615000 ;
      RECT 1123.865000  0.085000 1124.035000 0.525000 ;
      RECT 1123.875000  1.615000 1124.145000 2.405000 ;
      RECT 1124.085000  1.075000 1124.595000 1.275000 ;
      RECT 1124.205000  0.280000 1124.595000 0.695000 ;
      RECT 1124.335000  1.455000 1124.595000 2.635000 ;
      RECT 1124.785000  0.085000 1125.075000 0.810000 ;
      RECT 1124.785000  1.470000 1125.075000 2.635000 ;
      RECT 1125.245000  1.075000 1125.595000 1.275000 ;
      RECT 1125.260000  0.255000 1126.530000 0.475000 ;
      RECT 1125.260000  0.475000 1125.510000 0.895000 ;
      RECT 1125.300000  1.455000 1125.550000 2.635000 ;
      RECT 1125.680000  0.645000 1126.060000 0.865000 ;
      RECT 1125.770000  1.445000 1126.060000 1.785000 ;
      RECT 1125.770000  1.785000 1129.910000 1.955000 ;
      RECT 1125.770000  1.955000 1126.020000 2.465000 ;
      RECT 1125.815000  0.865000 1126.060000 1.445000 ;
      RECT 1126.240000  2.125000 1127.010000 2.635000 ;
      RECT 1126.280000  0.475000 1126.530000 0.645000 ;
      RECT 1126.280000  0.645000 1128.460000 0.905000 ;
      RECT 1126.280000  1.075000 1127.345000 1.445000 ;
      RECT 1126.280000  1.445000 1128.720000 1.615000 ;
      RECT 1126.720000  0.255000 1129.010000 0.475000 ;
      RECT 1127.230000  2.125000 1127.480000 2.295000 ;
      RECT 1127.230000  2.295000 1128.420000 2.465000 ;
      RECT 1127.515000  1.075000 1128.170000 1.275000 ;
      RECT 1127.700000  1.955000 1127.950000 2.125000 ;
      RECT 1128.170000  2.125000 1128.420000 2.295000 ;
      RECT 1128.340000  1.075000 1128.720000 1.445000 ;
      RECT 1128.640000  2.125000 1128.970000 2.635000 ;
      RECT 1128.680000  0.475000 1129.010000 0.735000 ;
      RECT 1128.680000  0.735000 1130.890000 0.905000 ;
      RECT 1128.890000  1.075000 1129.270000 1.445000 ;
      RECT 1128.890000  1.445000 1130.425000 1.615000 ;
      RECT 1129.190000  2.125000 1129.440000 2.295000 ;
      RECT 1129.190000  2.295000 1130.380000 2.465000 ;
      RECT 1129.230000  0.085000 1129.400000 0.555000 ;
      RECT 1129.440000  1.075000 1130.035000 1.275000 ;
      RECT 1129.570000  0.255000 1129.950000 0.725000 ;
      RECT 1129.570000  0.725000 1130.890000 0.735000 ;
      RECT 1129.660000  1.955000 1129.910000 2.125000 ;
      RECT 1130.130000  1.785000 1130.380000 2.295000 ;
      RECT 1130.170000  0.085000 1130.340000 0.555000 ;
      RECT 1130.255000  1.075000 1130.995000 1.275000 ;
      RECT 1130.255000  1.275000 1130.425000 1.445000 ;
      RECT 1130.510000  0.255000 1130.890000 0.725000 ;
      RECT 1130.645000  1.455000 1130.850000 2.635000 ;
      RECT 1131.225000  0.085000 1131.515000 0.810000 ;
      RECT 1131.225000  1.470000 1131.515000 2.635000 ;
      RECT 1131.690000  1.075000 1133.500000 1.275000 ;
      RECT 1131.715000  0.255000 1137.735000 0.475000 ;
      RECT 1131.715000  0.475000 1131.965000 0.895000 ;
      RECT 1131.755000  1.485000 1132.005000 2.635000 ;
      RECT 1132.135000  0.645000 1133.925000 0.865000 ;
      RECT 1132.225000  1.445000 1136.165000 1.615000 ;
      RECT 1132.225000  1.615000 1132.475000 2.465000 ;
      RECT 1132.695000  1.825000 1132.945000 2.635000 ;
      RECT 1133.165000  1.615000 1133.925000 1.955000 ;
      RECT 1133.165000  1.955000 1133.415000 2.465000 ;
      RECT 1133.635000  2.125000 1134.405000 2.635000 ;
      RECT 1133.720000  0.865000 1133.925000 1.445000 ;
      RECT 1134.115000  0.645000 1138.285000 0.735000 ;
      RECT 1134.115000  0.735000 1142.045000 0.820000 ;
      RECT 1134.160000  1.075000 1136.525000 1.275000 ;
      RECT 1134.625000  1.785000 1135.775000 1.955000 ;
      RECT 1134.625000  1.955000 1134.875000 2.465000 ;
      RECT 1135.095000  2.125000 1135.345000 2.635000 ;
      RECT 1135.565000  1.955000 1135.775000 2.265000 ;
      RECT 1135.565000  2.265000 1137.735000 2.465000 ;
      RECT 1135.945000  1.615000 1136.165000 1.785000 ;
      RECT 1135.945000  1.785000 1140.165000 2.005000 ;
      RECT 1136.335000  1.275000 1136.525000 1.445000 ;
      RECT 1136.335000  1.445000 1137.995000 1.615000 ;
      RECT 1136.695000  0.995000 1137.435000 1.275000 ;
      RECT 1137.615000  0.820000 1142.045000 0.905000 ;
      RECT 1137.615000  1.075000 1137.995000 1.445000 ;
      RECT 1137.955000  0.255000 1138.285000 0.645000 ;
      RECT 1137.955000  2.175000 1138.205000 2.635000 ;
      RECT 1138.165000  1.075000 1138.545000 1.445000 ;
      RECT 1138.165000  1.445000 1140.920000 1.615000 ;
      RECT 1138.375000  2.265000 1140.595000 2.465000 ;
      RECT 1138.505000  0.085000 1138.675000 0.555000 ;
      RECT 1138.725000  1.075000 1140.335000 1.275000 ;
      RECT 1138.845000  0.255000 1139.225000 0.725000 ;
      RECT 1138.845000  0.725000 1140.165000 0.735000 ;
      RECT 1139.445000  0.085000 1139.615000 0.555000 ;
      RECT 1139.785000  0.255000 1140.165000 0.725000 ;
      RECT 1140.385000  0.085000 1140.555000 0.555000 ;
      RECT 1140.385000  1.785000 1141.535000 1.955000 ;
      RECT 1140.385000  1.955000 1140.595000 2.265000 ;
      RECT 1140.605000  1.075000 1141.735000 1.275000 ;
      RECT 1140.605000  1.275000 1140.920000 1.445000 ;
      RECT 1140.725000  0.255000 1141.105000 0.725000 ;
      RECT 1140.725000  0.725000 1142.045000 0.735000 ;
      RECT 1140.815000  2.125000 1141.065000 2.635000 ;
      RECT 1141.285000  1.445000 1141.535000 1.785000 ;
      RECT 1141.285000  1.955000 1141.535000 2.465000 ;
      RECT 1141.325000  0.085000 1141.495000 0.555000 ;
      RECT 1141.665000  0.255000 1142.045000 0.725000 ;
      RECT 1141.755000  1.445000 1142.005000 2.635000 ;
      RECT 1142.265000  0.085000 1142.555000 0.810000 ;
      RECT 1142.265000  1.470000 1142.555000 2.635000 ;
      RECT 1142.725000  0.365000 1143.005000 2.465000 ;
      RECT 1143.175000  0.715000 1144.445000 0.895000 ;
      RECT 1143.175000  0.895000 1143.500000 1.495000 ;
      RECT 1143.175000  1.495000 1144.915000 1.705000 ;
      RECT 1143.245000  1.875000 1144.000000 2.635000 ;
      RECT 1143.255000  0.085000 1143.425000 0.545000 ;
      RECT 1143.695000  0.295000 1145.035000 0.475000 ;
      RECT 1143.705000  1.075000 1144.175000 1.325000 ;
      RECT 1144.080000  0.645000 1144.445000 0.715000 ;
      RECT 1144.370000  1.075000 1144.795000 1.325000 ;
      RECT 1144.445000  1.705000 1144.915000 2.465000 ;
      RECT 1144.705000  0.475000 1145.035000 0.695000 ;
      RECT 1144.705000  0.695000 1145.995000 0.865000 ;
      RECT 1144.975000  1.075000 1145.305000 1.325000 ;
      RECT 1145.085000  1.325000 1145.305000 2.405000 ;
      RECT 1145.265000  0.085000 1145.435000 0.525000 ;
      RECT 1145.475000  1.075000 1145.950000 1.275000 ;
      RECT 1145.605000  0.280000 1145.995000 0.695000 ;
      RECT 1145.625000  1.455000 1146.180000 2.635000 ;
      RECT 1146.405000  0.085000 1146.695000 0.810000 ;
      RECT 1146.405000  1.470000 1146.695000 2.635000 ;
      RECT 1146.895000  1.445000 1147.145000 2.635000 ;
      RECT 1146.965000  0.085000 1147.135000 0.885000 ;
      RECT 1147.385000  0.365000 1147.635000 2.465000 ;
      RECT 1147.855000  0.715000 1149.145000 0.895000 ;
      RECT 1147.855000  0.895000 1148.135000 1.455000 ;
      RECT 1147.855000  1.455000 1149.475000 1.705000 ;
      RECT 1147.875000  1.875000 1148.675000 2.635000 ;
      RECT 1147.905000  0.085000 1148.085000 0.545000 ;
      RECT 1148.305000  1.075000 1148.670000 1.275000 ;
      RECT 1148.345000  0.295000 1149.710000 0.475000 ;
      RECT 1148.730000  0.645000 1149.145000 0.715000 ;
      RECT 1148.890000  1.075000 1149.405000 1.275000 ;
      RECT 1149.120000  1.705000 1149.475000 2.465000 ;
      RECT 1149.370000  0.475000 1149.710000 0.695000 ;
      RECT 1149.370000  0.695000 1150.670000 0.865000 ;
      RECT 1149.575000  1.075000 1149.955000 1.275000 ;
      RECT 1149.685000  1.275000 1149.955000 2.405000 ;
      RECT 1149.975000  0.085000 1150.145000 0.525000 ;
      RECT 1150.125000  1.075000 1150.485000 1.615000 ;
      RECT 1150.335000  0.280000 1150.670000 0.695000 ;
      RECT 1150.350000  1.795000 1150.670000 2.635000 ;
      RECT 1151.005000  0.085000 1151.295000 0.810000 ;
      RECT 1151.005000  1.470000 1151.295000 2.635000 ;
      RECT 1151.465000  0.725000 1153.300000 0.905000 ;
      RECT 1151.465000  0.905000 1151.750000 1.445000 ;
      RECT 1151.465000  1.445000 1153.260000 1.615000 ;
      RECT 1151.600000  1.825000 1151.850000 2.635000 ;
      RECT 1151.640000  0.085000 1151.810000 0.555000 ;
      RECT 1151.920000  1.075000 1153.810000 1.275000 ;
      RECT 1151.980000  0.265000 1152.360000 0.725000 ;
      RECT 1152.070000  1.615000 1152.320000 2.465000 ;
      RECT 1152.540000  1.795000 1152.790000 2.635000 ;
      RECT 1152.580000  0.085000 1152.750000 0.555000 ;
      RECT 1152.920000  0.255000 1153.300000 0.725000 ;
      RECT 1153.010000  1.615000 1153.260000 2.465000 ;
      RECT 1153.480000  1.275000 1153.810000 1.785000 ;
      RECT 1153.480000  1.785000 1157.150000 1.955000 ;
      RECT 1153.480000  2.125000 1154.250000 2.635000 ;
      RECT 1153.520000  0.085000 1153.690000 0.555000 ;
      RECT 1153.520000  0.735000 1155.700000 0.905000 ;
      RECT 1153.520000  0.905000 1153.810000 1.075000 ;
      RECT 1153.960000  0.255000 1156.250000 0.475000 ;
      RECT 1153.995000  0.645000 1155.700000 0.735000 ;
      RECT 1154.000000  1.075000 1154.560000 1.445000 ;
      RECT 1154.000000  1.445000 1155.920000 1.615000 ;
      RECT 1154.470000  2.125000 1154.720000 2.295000 ;
      RECT 1154.470000  2.295000 1155.660000 2.465000 ;
      RECT 1154.730000  1.075000 1155.410000 1.275000 ;
      RECT 1154.940000  1.955000 1155.190000 2.125000 ;
      RECT 1155.410000  2.125000 1155.660000 2.295000 ;
      RECT 1155.580000  1.075000 1155.920000 1.445000 ;
      RECT 1155.880000  2.125000 1156.210000 2.635000 ;
      RECT 1155.920000  0.475000 1156.250000 0.735000 ;
      RECT 1155.920000  0.735000 1158.130000 0.905000 ;
      RECT 1156.090000  1.075000 1156.510000 1.445000 ;
      RECT 1156.090000  1.445000 1157.665000 1.615000 ;
      RECT 1156.430000  2.125000 1156.680000 2.295000 ;
      RECT 1156.430000  2.295000 1157.620000 2.465000 ;
      RECT 1156.470000  0.085000 1156.640000 0.555000 ;
      RECT 1156.730000  1.075000 1157.285000 1.275000 ;
      RECT 1156.810000  0.255000 1157.190000 0.725000 ;
      RECT 1156.810000  0.725000 1158.130000 0.735000 ;
      RECT 1156.900000  1.955000 1157.150000 2.125000 ;
      RECT 1157.370000  1.785000 1157.620000 2.295000 ;
      RECT 1157.410000  0.085000 1157.580000 0.555000 ;
      RECT 1157.455000  1.075000 1158.195000 1.275000 ;
      RECT 1157.455000  1.275000 1157.665000 1.445000 ;
      RECT 1157.750000  0.255000 1158.130000 0.725000 ;
      RECT 1157.885000  1.455000 1158.090000 2.635000 ;
      RECT 1158.365000  0.085000 1158.655000 0.810000 ;
      RECT 1158.365000  1.470000 1158.655000 2.635000 ;
      RECT 1158.825000  0.295000 1160.360000 0.475000 ;
      RECT 1158.825000  0.665000 1159.065000 1.990000 ;
      RECT 1158.875000  2.175000 1159.085000 2.635000 ;
      RECT 1159.235000  0.645000 1159.635000 0.825000 ;
      RECT 1159.235000  0.825000 1159.530000 1.835000 ;
      RECT 1159.235000  1.835000 1160.420000 2.045000 ;
      RECT 1159.790000  0.995000 1160.090000 1.665000 ;
      RECT 1159.870000  2.045000 1160.420000 2.465000 ;
      RECT 1160.030000  0.475000 1160.360000 0.695000 ;
      RECT 1160.030000  0.695000 1161.400000 0.825000 ;
      RECT 1160.200000  0.825000 1161.400000 0.865000 ;
      RECT 1160.305000  1.075000 1160.720000 1.245000 ;
      RECT 1160.490000  1.245000 1160.720000 1.445000 ;
      RECT 1160.490000  1.445000 1160.910000 1.615000 ;
      RECT 1160.630000  0.085000 1160.800000 0.525000 ;
      RECT 1160.660000  1.615000 1160.910000 2.405000 ;
      RECT 1160.890000  1.075000 1161.400000 1.275000 ;
      RECT 1161.010000  0.280000 1161.400000 0.695000 ;
      RECT 1161.080000  1.455000 1161.400000 2.635000 ;
      RECT 1161.585000  0.085000 1161.875000 0.810000 ;
      RECT 1161.585000  1.470000 1161.875000 2.635000 ;
      RECT 1162.050000  0.305000 1164.945000 0.475000 ;
      RECT 1162.050000  0.475000 1162.325000 0.905000 ;
      RECT 1162.110000  1.455000 1163.305000 1.625000 ;
      RECT 1162.110000  1.625000 1162.365000 2.465000 ;
      RECT 1162.160000  1.075000 1163.075000 1.285000 ;
      RECT 1162.495000  0.645000 1164.605000 0.905000 ;
      RECT 1162.585000  1.795000 1162.835000 2.635000 ;
      RECT 1163.055000  1.625000 1163.305000 2.295000 ;
      RECT 1163.055000  2.295000 1164.245000 2.465000 ;
      RECT 1163.285000  1.075000 1164.085000 1.275000 ;
      RECT 1163.525000  1.445000 1165.275000 1.625000 ;
      RECT 1163.525000  1.625000 1163.775000 2.125000 ;
      RECT 1163.995000  1.795000 1164.245000 2.295000 ;
      RECT 1164.365000  0.905000 1164.605000 1.445000 ;
      RECT 1164.555000  1.795000 1164.805000 2.295000 ;
      RECT 1164.555000  2.295000 1165.745000 2.465000 ;
      RECT 1164.775000  0.475000 1164.945000 0.725000 ;
      RECT 1164.775000  0.725000 1166.725000 0.905000 ;
      RECT 1164.795000  1.075000 1165.515000 1.275000 ;
      RECT 1165.025000  1.625000 1165.275000 2.125000 ;
      RECT 1165.115000  0.085000 1165.285000 0.555000 ;
      RECT 1165.455000  0.255000 1165.785000 0.725000 ;
      RECT 1165.495000  1.455000 1166.690000 1.625000 ;
      RECT 1165.495000  1.625000 1165.745000 2.295000 ;
      RECT 1165.725000  1.075000 1166.525000 1.285000 ;
      RECT 1165.965000  1.795000 1166.215000 2.635000 ;
      RECT 1166.005000  0.085000 1166.175000 0.555000 ;
      RECT 1166.345000  0.255000 1166.725000 0.725000 ;
      RECT 1166.435000  1.625000 1166.690000 2.465000 ;
      RECT 1167.105000  0.085000 1167.395000 0.810000 ;
      RECT 1167.105000  1.470000 1167.395000 2.635000 ;
      RECT 1167.565000  1.075000 1169.045000 1.275000 ;
      RECT 1167.605000  0.255000 1167.935000 0.725000 ;
      RECT 1167.605000  0.725000 1168.875000 0.735000 ;
      RECT 1167.605000  0.735000 1171.665000 0.905000 ;
      RECT 1167.645000  1.445000 1167.895000 2.635000 ;
      RECT 1168.115000  1.445000 1168.365000 1.785000 ;
      RECT 1168.115000  1.785000 1169.265000 1.955000 ;
      RECT 1168.115000  1.955000 1168.365000 2.465000 ;
      RECT 1168.155000  0.085000 1168.325000 0.555000 ;
      RECT 1168.495000  0.255000 1168.875000 0.725000 ;
      RECT 1168.585000  2.125000 1168.835000 2.635000 ;
      RECT 1168.730000  1.275000 1169.045000 1.445000 ;
      RECT 1168.730000  1.445000 1171.510000 1.615000 ;
      RECT 1169.055000  1.955000 1169.265000 2.295000 ;
      RECT 1169.055000  2.295000 1171.225000 2.465000 ;
      RECT 1169.095000  0.085000 1169.265000 0.555000 ;
      RECT 1169.315000  1.075000 1170.925000 1.275000 ;
      RECT 1169.435000  0.255000 1169.815000 0.725000 ;
      RECT 1169.435000  0.725000 1170.755000 0.735000 ;
      RECT 1169.435000  1.785000 1171.850000 1.955000 ;
      RECT 1169.435000  1.955000 1169.775000 2.125000 ;
      RECT 1169.995000  2.125000 1170.245000 2.295000 ;
      RECT 1170.035000  0.085000 1170.205000 0.555000 ;
      RECT 1170.375000  0.255000 1170.755000 0.725000 ;
      RECT 1170.465000  1.955000 1170.715000 2.125000 ;
      RECT 1170.935000  2.125000 1171.225000 2.295000 ;
      RECT 1170.975000  0.085000 1171.145000 0.555000 ;
      RECT 1171.105000  1.075000 1171.510000 1.445000 ;
      RECT 1171.315000  0.255000 1175.525000 0.475000 ;
      RECT 1171.315000  0.475000 1171.665000 0.735000 ;
      RECT 1171.445000  2.125000 1171.665000 2.635000 ;
      RECT 1171.680000  1.445000 1172.055000 1.615000 ;
      RECT 1171.680000  1.615000 1171.850000 1.785000 ;
      RECT 1171.835000  0.645000 1175.650000 0.820000 ;
      RECT 1171.835000  0.820000 1172.055000 1.445000 ;
      RECT 1171.835000  2.125000 1172.190000 2.465000 ;
      RECT 1172.020000  1.785000 1173.115000 1.955000 ;
      RECT 1172.020000  1.955000 1172.190000 2.125000 ;
      RECT 1172.225000  0.995000 1172.970000 1.445000 ;
      RECT 1172.225000  1.445000 1175.215000 1.615000 ;
      RECT 1172.405000  2.125000 1172.645000 2.635000 ;
      RECT 1172.865000  1.955000 1173.115000 2.295000 ;
      RECT 1172.865000  2.295000 1174.995000 2.465000 ;
      RECT 1173.140000  1.075000 1174.640000 1.275000 ;
      RECT 1173.335000  1.785000 1175.650000 1.955000 ;
      RECT 1173.335000  1.955000 1173.585000 2.125000 ;
      RECT 1173.805000  2.125000 1174.055000 2.295000 ;
      RECT 1174.275000  1.955000 1174.525000 2.125000 ;
      RECT 1174.745000  2.135000 1174.995000 2.295000 ;
      RECT 1174.945000  0.995000 1175.215000 1.445000 ;
      RECT 1175.215000  2.125000 1175.495000 2.635000 ;
      RECT 1175.385000  0.820000 1175.650000 1.785000 ;
      RECT 1175.845000  0.085000 1176.135000 0.810000 ;
      RECT 1175.845000  1.470000 1176.135000 2.635000 ;
      RECT 1176.305000  0.255000 1176.645000 0.825000 ;
      RECT 1176.305000  0.825000 1176.480000 1.795000 ;
      RECT 1176.305000  1.795000 1176.565000 2.465000 ;
      RECT 1176.650000  0.995000 1176.870000 1.445000 ;
      RECT 1176.650000  1.445000 1177.095000 1.615000 ;
      RECT 1176.735000  2.235000 1177.115000 2.635000 ;
      RECT 1176.890000  0.085000 1177.060000 0.750000 ;
      RECT 1176.925000  1.615000 1177.095000 1.885000 ;
      RECT 1176.925000  1.885000 1179.155000 2.055000 ;
      RECT 1177.040000  1.075000 1177.540000 1.275000 ;
      RECT 1177.235000  0.380000 1177.520000 0.735000 ;
      RECT 1177.235000  0.735000 1177.935000 0.905000 ;
      RECT 1177.265000  1.495000 1178.380000 1.715000 ;
      RECT 1177.710000  0.905000 1177.935000 1.100000 ;
      RECT 1177.780000  0.395000 1178.275000 0.565000 ;
      RECT 1178.085000  2.235000 1178.485000 2.635000 ;
      RECT 1178.105000  0.565000 1178.275000 1.355000 ;
      RECT 1178.105000  1.355000 1178.380000 1.495000 ;
      RECT 1178.445000  0.320000 1178.695000 0.690000 ;
      RECT 1178.525000  0.690000 1178.695000 1.075000 ;
      RECT 1178.525000  1.075000 1178.720000 1.245000 ;
      RECT 1178.550000  1.245000 1178.720000 1.495000 ;
      RECT 1178.550000  1.495000 1179.155000 1.885000 ;
      RECT 1178.775000  2.055000 1179.155000 2.290000 ;
      RECT 1178.915000  0.320000 1179.165000 0.725000 ;
      RECT 1178.915000  0.725000 1180.275000 0.905000 ;
      RECT 1178.940000  1.075000 1179.755000 1.325000 ;
      RECT 1179.355000  0.085000 1179.705000 0.555000 ;
      RECT 1179.555000  1.325000 1179.755000 2.425000 ;
      RECT 1179.885000  0.320000 1180.275000 0.725000 ;
      RECT 1179.925000  1.075000 1180.275000 1.645000 ;
      RECT 1179.925000  1.815000 1180.275000 2.635000 ;
      RECT 1180.445000  0.085000 1180.735000 0.810000 ;
      RECT 1180.445000  1.470000 1180.735000 2.635000 ;
      RECT 1180.930000  0.085000 1181.185000 0.910000 ;
      RECT 1180.930000  1.410000 1181.185000 2.635000 ;
      RECT 1181.355000  0.255000 1181.740000 0.825000 ;
      RECT 1181.355000  0.825000 1181.575000 1.795000 ;
      RECT 1181.355000  1.795000 1181.660000 2.465000 ;
      RECT 1181.745000  0.995000 1181.965000 1.445000 ;
      RECT 1181.745000  1.445000 1182.190000 1.615000 ;
      RECT 1181.830000  2.235000 1182.210000 2.635000 ;
      RECT 1181.955000  0.085000 1182.125000 0.750000 ;
      RECT 1182.020000  1.615000 1182.190000 1.885000 ;
      RECT 1182.020000  1.885000 1184.255000 2.055000 ;
      RECT 1182.135000  1.075000 1182.655000 1.275000 ;
      RECT 1182.340000  0.380000 1182.705000 0.735000 ;
      RECT 1182.340000  0.735000 1183.045000 0.905000 ;
      RECT 1182.360000  1.495000 1183.480000 1.715000 ;
      RECT 1182.825000  0.905000 1183.045000 1.100000 ;
      RECT 1182.875000  0.395000 1183.385000 0.565000 ;
      RECT 1183.180000  2.235000 1183.585000 2.635000 ;
      RECT 1183.215000  0.565000 1183.385000 1.355000 ;
      RECT 1183.215000  1.355000 1183.480000 1.495000 ;
      RECT 1183.555000  0.320000 1183.800000 0.690000 ;
      RECT 1183.630000  0.690000 1183.800000 1.075000 ;
      RECT 1183.630000  1.075000 1183.820000 1.245000 ;
      RECT 1183.650000  1.245000 1183.820000 1.495000 ;
      RECT 1183.650000  1.495000 1184.255000 1.885000 ;
      RECT 1183.855000  2.055000 1184.255000 2.425000 ;
      RECT 1184.025000  0.320000 1184.255000 0.725000 ;
      RECT 1184.025000  0.725000 1185.225000 0.905000 ;
      RECT 1184.040000  1.075000 1184.645000 1.325000 ;
      RECT 1184.475000  1.325000 1184.645000 1.915000 ;
      RECT 1184.475000  1.915000 1184.815000 2.425000 ;
      RECT 1184.495000  0.085000 1184.665000 0.555000 ;
      RECT 1184.820000  1.075000 1185.285000 1.645000 ;
      RECT 1184.835000  0.320000 1185.225000 0.725000 ;
      RECT 1184.985000  1.815000 1185.300000 2.635000 ;
      RECT 1185.505000  0.085000 1185.795000 0.810000 ;
      RECT 1185.505000  1.470000 1185.795000 2.635000 ;
      RECT 1185.965000  1.075000 1186.505000 1.445000 ;
      RECT 1185.965000  1.445000 1187.975000 1.615000 ;
      RECT 1185.975000  0.255000 1186.305000 0.725000 ;
      RECT 1185.975000  0.725000 1187.245000 0.735000 ;
      RECT 1185.975000  0.735000 1188.105000 0.905000 ;
      RECT 1186.020000  1.795000 1186.225000 2.635000 ;
      RECT 1186.485000  1.785000 1186.735000 2.295000 ;
      RECT 1186.485000  2.295000 1187.675000 2.465000 ;
      RECT 1186.525000  0.085000 1186.695000 0.555000 ;
      RECT 1186.735000  1.075000 1187.325000 1.275000 ;
      RECT 1186.865000  0.255000 1187.245000 0.725000 ;
      RECT 1186.955000  1.785000 1188.745000 1.955000 ;
      RECT 1186.955000  1.955000 1187.205000 2.125000 ;
      RECT 1187.425000  2.125000 1187.675000 2.295000 ;
      RECT 1187.465000  0.085000 1187.635000 0.555000 ;
      RECT 1187.595000  1.075000 1187.975000 1.445000 ;
      RECT 1187.805000  0.255000 1189.125000 0.475000 ;
      RECT 1187.805000  0.475000 1188.105000 0.735000 ;
      RECT 1187.895000  2.125000 1188.145000 2.635000 ;
      RECT 1188.145000  1.075000 1188.575000 1.415000 ;
      RECT 1188.145000  1.415000 1188.745000 1.785000 ;
      RECT 1188.275000  0.645000 1188.655000 0.815000 ;
      RECT 1188.275000  0.815000 1188.575000 1.075000 ;
      RECT 1188.365000  1.955000 1188.745000 1.965000 ;
      RECT 1188.365000  1.965000 1188.655000 2.465000 ;
      RECT 1188.745000  1.075000 1189.325000 1.245000 ;
      RECT 1188.875000  2.135000 1189.605000 2.635000 ;
      RECT 1189.135000  0.725000 1190.585000 0.905000 ;
      RECT 1189.135000  0.905000 1189.325000 1.075000 ;
      RECT 1189.135000  1.245000 1189.325000 1.785000 ;
      RECT 1189.135000  1.785000 1191.015000 1.965000 ;
      RECT 1189.395000  0.085000 1189.565000 0.555000 ;
      RECT 1189.495000  1.075000 1189.875000 1.445000 ;
      RECT 1189.495000  1.445000 1191.345000 1.615000 ;
      RECT 1189.735000  0.305000 1191.055000 0.475000 ;
      RECT 1189.825000  1.965000 1190.075000 2.125000 ;
      RECT 1190.045000  1.075000 1190.765000 1.275000 ;
      RECT 1190.205000  0.645000 1190.585000 0.725000 ;
      RECT 1190.295000  2.135000 1190.545000 2.635000 ;
      RECT 1190.765000  1.965000 1191.015000 2.465000 ;
      RECT 1190.805000  0.475000 1191.055000 0.895000 ;
      RECT 1190.935000  1.075000 1191.345000 1.445000 ;
      RECT 1191.235000  1.795000 1191.485000 2.635000 ;
      RECT 1191.275000  0.085000 1191.445000 0.895000 ;
      RECT 1191.545000  1.075000 1192.965000 1.245000 ;
      RECT 1191.545000  1.245000 1191.885000 1.615000 ;
      RECT 1191.615000  0.275000 1191.995000 0.725000 ;
      RECT 1191.615000  0.725000 1193.590000 0.905000 ;
      RECT 1191.705000  1.785000 1192.895000 1.955000 ;
      RECT 1191.705000  1.955000 1191.955000 2.465000 ;
      RECT 1192.175000  2.165000 1192.425000 2.635000 ;
      RECT 1192.215000  0.085000 1192.385000 0.555000 ;
      RECT 1192.555000  0.275000 1192.935000 0.725000 ;
      RECT 1192.645000  1.415000 1193.590000 1.655000 ;
      RECT 1192.645000  1.655000 1192.895000 1.785000 ;
      RECT 1192.645000  1.955000 1192.895000 2.465000 ;
      RECT 1193.115000  1.825000 1193.365000 2.635000 ;
      RECT 1193.155000  0.085000 1193.325000 0.555000 ;
      RECT 1193.285000  0.905000 1193.590000 1.415000 ;
      RECT 1193.785000  0.085000 1194.075000 0.810000 ;
      RECT 1193.785000  1.470000 1194.075000 2.635000 ;
      RECT 1194.245000  0.985000 1194.595000 1.285000 ;
      RECT 1194.250000  0.085000 1194.585000 0.815000 ;
      RECT 1194.310000  1.455000 1194.560000 2.635000 ;
      RECT 1194.765000  0.280000 1194.985000 0.995000 ;
      RECT 1194.765000  0.995000 1195.260000 1.325000 ;
      RECT 1194.780000  1.495000 1195.600000 1.665000 ;
      RECT 1194.780000  1.665000 1195.030000 2.465000 ;
      RECT 1195.160000  0.280000 1195.600000 0.825000 ;
      RECT 1195.250000  1.835000 1195.940000 2.635000 ;
      RECT 1195.430000  0.825000 1195.600000 0.995000 ;
      RECT 1195.430000  0.995000 1195.740000 1.325000 ;
      RECT 1195.430000  1.325000 1195.600000 1.495000 ;
      RECT 1195.770000  0.430000 1196.090000 0.790000 ;
      RECT 1195.920000  0.790000 1196.090000 1.445000 ;
      RECT 1195.920000  1.445000 1196.435000 1.665000 ;
      RECT 1196.110000  1.665000 1196.435000 2.465000 ;
      RECT 1196.260000  0.425000 1196.510000 0.725000 ;
      RECT 1196.260000  0.725000 1197.400000 0.905000 ;
      RECT 1196.310000  1.075000 1196.775000 1.275000 ;
      RECT 1196.605000  1.275000 1196.775000 2.425000 ;
      RECT 1196.680000  0.085000 1196.850000 0.555000 ;
      RECT 1197.020000  0.275000 1197.400000 0.725000 ;
      RECT 1197.025000  1.075000 1197.405000 1.285000 ;
      RECT 1197.110000  1.455000 1197.360000 2.635000 ;
      RECT 1197.925000  0.085000 1198.215000 0.810000 ;
      RECT 1197.925000  1.470000 1198.215000 2.635000 ;
      RECT 1198.390000  1.075000 1198.975000 1.445000 ;
      RECT 1198.390000  1.445000 1200.445000 1.615000 ;
      RECT 1198.450000  1.795000 1198.700000 2.635000 ;
      RECT 1198.495000  0.085000 1198.665000 0.895000 ;
      RECT 1198.835000  0.305000 1200.155000 0.475000 ;
      RECT 1198.835000  0.475000 1199.135000 0.895000 ;
      RECT 1198.925000  1.785000 1200.785000 1.965000 ;
      RECT 1198.925000  1.965000 1199.175000 2.465000 ;
      RECT 1199.145000  1.075000 1199.800000 1.275000 ;
      RECT 1199.305000  0.645000 1199.685000 0.725000 ;
      RECT 1199.305000  0.725000 1200.785000 0.905000 ;
      RECT 1199.395000  2.135000 1199.645000 2.635000 ;
      RECT 1200.065000  1.075000 1200.445000 1.445000 ;
      RECT 1200.335000  0.085000 1200.505000 0.555000 ;
      RECT 1200.335000  2.135000 1201.025000 2.635000 ;
      RECT 1200.615000  0.905000 1200.785000 0.995000 ;
      RECT 1200.615000  0.995000 1201.025000 1.325000 ;
      RECT 1200.615000  1.325000 1200.785000 1.785000 ;
      RECT 1200.775000  0.255000 1202.080000 0.475000 ;
      RECT 1200.775000  0.475000 1201.025000 0.555000 ;
      RECT 1201.195000  0.645000 1201.575000 1.075000 ;
      RECT 1201.195000  1.075000 1201.765000 1.785000 ;
      RECT 1201.195000  1.785000 1202.980000 1.955000 ;
      RECT 1201.195000  1.955000 1201.535000 2.465000 ;
      RECT 1201.755000  2.125000 1202.040000 2.635000 ;
      RECT 1201.795000  0.475000 1202.080000 0.735000 ;
      RECT 1201.795000  0.735000 1203.960000 0.905000 ;
      RECT 1201.950000  1.075000 1202.340000 1.445000 ;
      RECT 1201.950000  1.445000 1203.760000 1.615000 ;
      RECT 1202.260000  2.125000 1202.510000 2.295000 ;
      RECT 1202.260000  2.295000 1203.450000 2.465000 ;
      RECT 1202.300000  0.085000 1202.470000 0.555000 ;
      RECT 1202.560000  1.075000 1203.200000 1.275000 ;
      RECT 1202.640000  0.255000 1203.020000 0.725000 ;
      RECT 1202.640000  0.725000 1203.960000 0.735000 ;
      RECT 1202.730000  1.955000 1202.980000 2.125000 ;
      RECT 1203.200000  1.785000 1203.450000 2.295000 ;
      RECT 1203.240000  0.085000 1203.410000 0.555000 ;
      RECT 1203.430000  1.075000 1203.760000 1.445000 ;
      RECT 1203.580000  0.255000 1203.960000 0.725000 ;
      RECT 1203.715000  1.795000 1203.920000 2.635000 ;
      RECT 1204.365000  0.085000 1204.655000 0.810000 ;
      RECT 1204.365000  1.470000 1204.655000 2.635000 ;
      RECT 1204.825000  0.645000 1206.595000 0.905000 ;
      RECT 1204.825000  0.905000 1204.995000 1.455000 ;
      RECT 1204.825000  1.455000 1209.055000 1.625000 ;
      RECT 1204.840000  0.255000 1207.065000 0.475000 ;
      RECT 1204.895000  1.795000 1205.145000 2.635000 ;
      RECT 1205.165000  1.075000 1206.765000 1.285000 ;
      RECT 1205.365000  1.625000 1205.615000 2.465000 ;
      RECT 1205.835000  1.795000 1206.085000 2.635000 ;
      RECT 1206.305000  1.625000 1206.555000 2.465000 ;
      RECT 1206.775000  1.795000 1207.025000 2.635000 ;
      RECT 1206.815000  0.475000 1207.065000 0.725000 ;
      RECT 1206.815000  0.725000 1208.945000 0.905000 ;
      RECT 1207.035000  1.075000 1208.645000 1.285000 ;
      RECT 1207.245000  1.625000 1207.495000 2.465000 ;
      RECT 1207.285000  0.085000 1207.455000 0.555000 ;
      RECT 1207.625000  0.255000 1208.005000 0.725000 ;
      RECT 1207.715000  1.795000 1207.965000 2.635000 ;
      RECT 1208.185000  1.625000 1208.435000 2.465000 ;
      RECT 1208.225000  0.085000 1208.395000 0.555000 ;
      RECT 1208.565000  0.255000 1208.945000 0.725000 ;
      RECT 1208.655000  1.795000 1209.395000 2.635000 ;
      RECT 1208.885000  1.075000 1211.045000 1.285000 ;
      RECT 1208.885000  1.285000 1209.055000 1.455000 ;
      RECT 1209.200000  0.255000 1211.885000 0.475000 ;
      RECT 1209.200000  0.475000 1209.385000 0.835000 ;
      RECT 1209.605000  0.645000 1211.545000 0.905000 ;
      RECT 1209.615000  1.455000 1213.205000 1.625000 ;
      RECT 1209.615000  1.625000 1209.865000 2.465000 ;
      RECT 1210.085000  1.795000 1210.335000 2.635000 ;
      RECT 1210.555000  1.625000 1210.805000 2.465000 ;
      RECT 1211.025000  1.795000 1211.275000 2.635000 ;
      RECT 1211.215000  0.905000 1211.545000 1.455000 ;
      RECT 1211.515000  1.795000 1211.795000 2.295000 ;
      RECT 1211.515000  2.295000 1213.675000 2.465000 ;
      RECT 1211.715000  0.475000 1211.885000 0.735000 ;
      RECT 1211.715000  0.735000 1215.595000 0.905000 ;
      RECT 1211.805000  1.075000 1213.415000 1.285000 ;
      RECT 1212.015000  1.625000 1212.265000 2.125000 ;
      RECT 1212.055000  0.085000 1212.225000 0.555000 ;
      RECT 1212.395000  0.255000 1212.775000 0.725000 ;
      RECT 1212.395000  0.725000 1215.595000 0.735000 ;
      RECT 1212.485000  1.795000 1212.735000 2.295000 ;
      RECT 1212.955000  1.625000 1213.205000 2.125000 ;
      RECT 1212.995000  0.085000 1213.165000 0.555000 ;
      RECT 1213.335000  0.255000 1213.715000 0.725000 ;
      RECT 1213.425000  1.455000 1215.615000 1.625000 ;
      RECT 1213.425000  1.625000 1213.675000 2.295000 ;
      RECT 1213.585000  1.075000 1215.680000 1.285000 ;
      RECT 1213.895000  1.795000 1214.145000 2.635000 ;
      RECT 1213.935000  0.085000 1214.105000 0.555000 ;
      RECT 1214.275000  0.255000 1214.655000 0.725000 ;
      RECT 1214.365000  1.625000 1214.615000 2.465000 ;
      RECT 1214.835000  1.795000 1215.085000 2.635000 ;
      RECT 1214.875000  0.085000 1215.045000 0.555000 ;
      RECT 1215.215000  0.255000 1215.595000 0.725000 ;
      RECT 1215.305000  1.625000 1215.615000 2.465000 ;
      RECT 1215.865000  0.085000 1216.155000 0.810000 ;
      RECT 1215.865000  1.470000 1216.155000 2.635000 ;
      RECT 1216.325000  1.495000 1216.660000 2.635000 ;
      RECT 1216.330000  1.075000 1216.675000 1.325000 ;
      RECT 1216.415000  0.085000 1216.585000 0.905000 ;
      RECT 1216.755000  0.255000 1217.135000 0.735000 ;
      RECT 1216.755000  0.735000 1217.955000 0.905000 ;
      RECT 1216.845000  1.075000 1217.345000 2.465000 ;
      RECT 1217.365000  0.085000 1217.535000 0.565000 ;
      RECT 1217.555000  1.075000 1217.935000 1.325000 ;
      RECT 1217.695000  1.325000 1217.935000 2.405000 ;
      RECT 1217.705000  0.460000 1217.955000 0.735000 ;
      RECT 1218.125000  0.260000 1218.735000 0.825000 ;
      RECT 1218.125000  0.825000 1218.395000 2.465000 ;
      RECT 1218.565000  0.995000 1218.890000 1.325000 ;
      RECT 1218.595000  1.495000 1218.765000 2.635000 ;
      RECT 1219.085000  0.085000 1219.375000 0.810000 ;
      RECT 1219.085000  1.470000 1219.375000 2.635000 ;
      RECT 1219.550000  0.255000 1219.905000 0.715000 ;
      RECT 1219.550000  0.715000 1223.315000 0.885000 ;
      RECT 1219.550000  1.055000 1220.770000 1.325000 ;
      RECT 1219.550000  1.495000 1221.785000 1.665000 ;
      RECT 1219.550000  1.665000 1219.905000 2.465000 ;
      RECT 1220.125000  0.085000 1220.295000 0.545000 ;
      RECT 1220.125000  1.835000 1220.295000 2.635000 ;
      RECT 1220.465000  0.255000 1220.845000 0.715000 ;
      RECT 1220.465000  1.665000 1220.845000 2.465000 ;
      RECT 1220.960000  1.055000 1221.880000 1.325000 ;
      RECT 1221.065000  0.085000 1221.625000 0.545000 ;
      RECT 1221.065000  1.835000 1221.235000 2.295000 ;
      RECT 1221.065000  2.295000 1222.765000 2.465000 ;
      RECT 1221.405000  1.665000 1221.785000 2.125000 ;
      RECT 1221.885000  0.255000 1222.215000 0.715000 ;
      RECT 1222.045000  1.495000 1224.425000 1.665000 ;
      RECT 1222.045000  1.665000 1222.375000 2.125000 ;
      RECT 1222.160000  1.055000 1223.015000 1.325000 ;
      RECT 1222.385000  0.085000 1222.765000 0.545000 ;
      RECT 1222.595000  1.835000 1222.765000 2.295000 ;
      RECT 1222.935000  0.255000 1224.425000 0.425000 ;
      RECT 1222.935000  0.425000 1223.315000 0.715000 ;
      RECT 1222.935000  1.665000 1223.315000 2.465000 ;
      RECT 1223.535000  0.595000 1223.915000 1.495000 ;
      RECT 1223.535000  1.835000 1223.865000 2.635000 ;
      RECT 1224.085000  1.665000 1224.425000 2.465000 ;
      RECT 1224.090000  0.425000 1224.425000 0.585000 ;
      RECT 1224.090000  0.755000 1224.430000 1.325000 ;
      RECT 1224.605000  0.085000 1224.895000 0.810000 ;
      RECT 1224.605000  1.470000 1224.895000 2.635000 ;
      RECT 1225.070000  0.255000 1225.425000 0.715000 ;
      RECT 1225.070000  0.715000 1231.570000 0.885000 ;
      RECT 1225.070000  1.055000 1226.910000 1.425000 ;
      RECT 1225.070000  1.595000 1227.305000 1.895000 ;
      RECT 1225.070000  1.895000 1225.425000 2.465000 ;
      RECT 1225.645000  0.085000 1225.815000 0.545000 ;
      RECT 1225.645000  2.065000 1225.815000 2.635000 ;
      RECT 1225.985000  0.255000 1226.365000 0.715000 ;
      RECT 1225.985000  1.895000 1226.365000 2.465000 ;
      RECT 1226.585000  0.085000 1226.755000 0.545000 ;
      RECT 1226.585000  2.065000 1226.755000 2.635000 ;
      RECT 1226.925000  0.255000 1227.305000 0.715000 ;
      RECT 1226.925000  1.895000 1227.305000 2.205000 ;
      RECT 1226.925000  2.205000 1229.265000 2.465000 ;
      RECT 1227.130000  1.055000 1228.985000 1.425000 ;
      RECT 1227.525000  0.085000 1227.695000 0.545000 ;
      RECT 1227.525000  1.595000 1228.985000 1.765000 ;
      RECT 1227.525000  1.765000 1227.695000 2.035000 ;
      RECT 1227.865000  0.255000 1228.245000 0.715000 ;
      RECT 1227.865000  1.935000 1228.245000 2.205000 ;
      RECT 1228.465000  0.085000 1228.635000 0.545000 ;
      RECT 1228.465000  1.765000 1228.985000 1.865000 ;
      RECT 1228.465000  1.865000 1231.180000 2.035000 ;
      RECT 1228.805000  0.255000 1229.185000 0.715000 ;
      RECT 1229.155000  1.055000 1231.570000 1.275000 ;
      RECT 1229.155000  1.445000 1233.605000 1.695000 ;
      RECT 1229.425000  0.085000 1230.120000 0.545000 ;
      RECT 1229.510000  2.035000 1231.180000 2.465000 ;
      RECT 1230.340000  0.395000 1230.510000 0.715000 ;
      RECT 1230.770000  0.085000 1231.140000 0.545000 ;
      RECT 1231.400000  0.255000 1233.565000 0.475000 ;
      RECT 1231.400000  0.475000 1231.570000 0.715000 ;
      RECT 1231.400000  1.695000 1231.570000 2.465000 ;
      RECT 1231.740000  0.645000 1233.060000 0.885000 ;
      RECT 1231.740000  0.885000 1231.975000 1.445000 ;
      RECT 1231.740000  1.890000 1232.120000 2.635000 ;
      RECT 1232.145000  1.055000 1233.565000 1.275000 ;
      RECT 1232.340000  1.695000 1232.510000 2.465000 ;
      RECT 1232.680000  1.890000 1233.060000 2.635000 ;
      RECT 1233.280000  0.475000 1233.565000 0.885000 ;
      RECT 1233.280000  1.695000 1233.605000 2.465000 ;
      RECT 1233.805000  0.085000 1234.095000 0.810000 ;
      RECT 1233.805000  1.470000 1234.095000 2.635000 ;
      RECT 1234.265000  0.255000 1235.620000 0.485000 ;
      RECT 1234.270000  0.685000 1234.540000 1.325000 ;
      RECT 1234.270000  1.495000 1234.540000 2.635000 ;
      RECT 1234.710000  0.655000 1235.075000 0.825000 ;
      RECT 1234.710000  0.825000 1234.930000 1.785000 ;
      RECT 1234.710000  1.785000 1235.710000 2.465000 ;
      RECT 1235.100000  0.995000 1235.485000 1.615000 ;
      RECT 1235.245000  0.485000 1235.620000 0.655000 ;
      RECT 1235.245000  0.655000 1236.735000 0.825000 ;
      RECT 1235.655000  0.995000 1235.925000 1.615000 ;
      RECT 1235.825000  0.085000 1236.155000 0.485000 ;
      RECT 1236.095000  0.995000 1236.385000 2.465000 ;
      RECT 1236.565000  0.375000 1236.735000 0.655000 ;
      RECT 1236.575000  0.995000 1237.170000 1.325000 ;
      RECT 1236.905000  0.085000 1237.275000 0.825000 ;
      RECT 1236.965000  1.495000 1237.315000 2.635000 ;
      RECT 1237.485000  0.085000 1237.775000 0.810000 ;
      RECT 1237.485000  1.470000 1237.775000 2.635000 ;
      RECT 1237.950000  0.255000 1240.515000 0.485000 ;
      RECT 1237.950000  0.485000 1238.205000 0.905000 ;
      RECT 1237.950000  1.075000 1238.755000 1.325000 ;
      RECT 1237.950000  1.495000 1238.205000 2.295000 ;
      RECT 1237.950000  2.295000 1239.225000 2.465000 ;
      RECT 1238.375000  0.655000 1240.105000 0.905000 ;
      RECT 1238.375000  1.495000 1241.265000 1.665000 ;
      RECT 1238.375000  1.665000 1238.755000 2.095000 ;
      RECT 1238.925000  1.075000 1239.675000 1.325000 ;
      RECT 1238.975000  1.835000 1240.165000 2.005000 ;
      RECT 1238.975000  2.005000 1239.225000 2.295000 ;
      RECT 1239.445000  2.175000 1239.615000 2.635000 ;
      RECT 1239.785000  2.005000 1240.165000 2.455000 ;
      RECT 1239.845000  0.905000 1240.105000 1.105000 ;
      RECT 1239.845000  1.105000 1240.230000 1.495000 ;
      RECT 1240.345000  0.485000 1240.515000 0.715000 ;
      RECT 1240.345000  0.715000 1244.165000 0.905000 ;
      RECT 1240.445000  1.835000 1240.695000 2.255000 ;
      RECT 1240.445000  2.255000 1242.695000 2.445000 ;
      RECT 1240.515000  1.075000 1241.225000 1.325000 ;
      RECT 1240.730000  0.085000 1241.110000 0.545000 ;
      RECT 1240.885000  1.665000 1241.265000 2.085000 ;
      RECT 1241.295000  0.255000 1241.675000 0.715000 ;
      RECT 1241.485000  1.495000 1241.655000 2.255000 ;
      RECT 1241.580000  1.075000 1242.790000 1.325000 ;
      RECT 1241.875000  1.495000 1243.685000 1.665000 ;
      RECT 1241.875000  1.665000 1242.205000 2.085000 ;
      RECT 1241.895000  0.085000 1242.065000 0.545000 ;
      RECT 1242.365000  0.255000 1243.035000 0.715000 ;
      RECT 1242.445000  1.835000 1242.695000 2.255000 ;
      RECT 1242.930000  1.835000 1243.135000 2.635000 ;
      RECT 1243.060000  1.075000 1244.155000 1.325000 ;
      RECT 1243.215000  0.085000 1243.595000 0.545000 ;
      RECT 1243.355000  1.665000 1243.685000 2.460000 ;
      RECT 1243.835000  0.255000 1244.165000 0.715000 ;
      RECT 1243.905000  1.495000 1244.125000 2.635000 ;
      RECT 1244.385000  0.085000 1244.675000 0.810000 ;
      RECT 1244.385000  1.470000 1244.675000 2.635000 ;
      RECT 1244.850000  0.255000 1248.960000 0.465000 ;
      RECT 1244.850000  0.465000 1245.105000 0.905000 ;
      RECT 1244.850000  1.495000 1245.105000 2.255000 ;
      RECT 1244.850000  2.255000 1247.000000 2.465000 ;
      RECT 1244.870000  1.075000 1246.595000 1.275000 ;
      RECT 1245.275000  0.655000 1248.490000 0.905000 ;
      RECT 1245.275000  1.495000 1250.890000 1.665000 ;
      RECT 1245.275000  1.665000 1245.655000 2.085000 ;
      RECT 1245.875000  1.835000 1246.045000 2.255000 ;
      RECT 1246.215000  1.665000 1246.610000 2.085000 ;
      RECT 1246.815000  0.905000 1246.995000 1.495000 ;
      RECT 1246.830000  1.835000 1248.960000 2.005000 ;
      RECT 1246.830000  2.005000 1247.000000 2.255000 ;
      RECT 1247.165000  1.075000 1248.700000 1.275000 ;
      RECT 1247.170000  2.175000 1247.550000 2.635000 ;
      RECT 1247.770000  2.005000 1247.940000 2.425000 ;
      RECT 1248.110000  2.175000 1248.490000 2.635000 ;
      RECT 1248.710000  0.465000 1248.960000 0.735000 ;
      RECT 1248.710000  0.735000 1255.685000 0.905000 ;
      RECT 1248.710000  2.005000 1248.960000 2.465000 ;
      RECT 1248.930000  1.075000 1250.740000 1.275000 ;
      RECT 1249.150000  1.835000 1249.400000 2.255000 ;
      RECT 1249.150000  2.255000 1253.240000 2.465000 ;
      RECT 1249.180000  0.085000 1249.350000 0.545000 ;
      RECT 1249.520000  0.255000 1249.900000 0.735000 ;
      RECT 1249.620000  1.665000 1249.950000 2.085000 ;
      RECT 1250.120000  0.085000 1250.450000 0.545000 ;
      RECT 1250.170000  1.835000 1250.340000 2.255000 ;
      RECT 1250.510000  1.665000 1250.890000 2.085000 ;
      RECT 1250.670000  0.255000 1251.340000 0.735000 ;
      RECT 1251.110000  1.835000 1251.280000 2.255000 ;
      RECT 1251.280000  1.075000 1252.770000 1.275000 ;
      RECT 1251.450000  1.495000 1255.170000 1.665000 ;
      RECT 1251.450000  1.665000 1251.830000 2.085000 ;
      RECT 1251.580000  0.085000 1251.750000 0.545000 ;
      RECT 1251.920000  0.255000 1252.300000 0.735000 ;
      RECT 1252.050000  1.835000 1252.220000 2.255000 ;
      RECT 1252.390000  1.665000 1252.770000 2.085000 ;
      RECT 1252.520000  0.085000 1252.690000 0.545000 ;
      RECT 1252.860000  0.255000 1253.600000 0.735000 ;
      RECT 1252.990000  1.835000 1253.240000 2.255000 ;
      RECT 1253.430000  1.835000 1253.680000 2.635000 ;
      RECT 1253.850000  1.075000 1255.685000 1.275000 ;
      RECT 1253.850000  1.665000 1254.230000 2.465000 ;
      RECT 1253.980000  0.085000 1254.150000 0.545000 ;
      RECT 1254.320000  0.255000 1254.700000 0.735000 ;
      RECT 1254.450000  1.835000 1254.620000 2.635000 ;
      RECT 1254.790000  1.665000 1255.170000 2.465000 ;
      RECT 1254.920000  0.085000 1255.135000 0.545000 ;
      RECT 1255.305000  0.255000 1255.685000 0.735000 ;
      RECT 1255.435000  1.495000 1255.685000 2.635000 ;
      RECT 1255.885000  0.085000 1256.175000 0.810000 ;
      RECT 1255.885000  1.470000 1256.175000 2.635000 ;
      RECT 1256.345000  0.765000 1256.700000 1.325000 ;
      RECT 1256.370000  0.085000 1256.610000 0.595000 ;
      RECT 1256.380000  1.495000 1258.005000 1.665000 ;
      RECT 1256.380000  1.665000 1256.770000 1.840000 ;
      RECT 1256.870000  0.265000 1257.110000 0.595000 ;
      RECT 1256.870000  0.595000 1257.040000 1.495000 ;
      RECT 1257.210000  0.765000 1257.545000 1.325000 ;
      RECT 1257.355000  1.835000 1257.685000 2.635000 ;
      RECT 1257.390000  0.085000 1257.605000 0.595000 ;
      RECT 1257.775000  0.255000 1258.475000 0.825000 ;
      RECT 1257.785000  0.995000 1258.005000 1.495000 ;
      RECT 1257.905000  1.845000 1258.475000 2.465000 ;
      RECT 1258.175000  0.825000 1258.475000 1.845000 ;
      RECT 1258.645000  0.085000 1258.935000 0.810000 ;
      RECT 1258.645000  1.470000 1258.935000 2.635000 ;
      RECT 1259.125000  0.085000 1259.365000 0.595000 ;
      RECT 1259.145000  0.765000 1259.365000 1.325000 ;
      RECT 1259.175000  1.495000 1260.785000 1.665000 ;
      RECT 1259.175000  1.665000 1259.535000 1.840000 ;
      RECT 1259.535000  0.255000 1259.875000 0.595000 ;
      RECT 1259.535000  0.595000 1259.765000 1.495000 ;
      RECT 1259.935000  0.765000 1260.395000 1.325000 ;
      RECT 1260.155000  0.085000 1260.470000 0.595000 ;
      RECT 1260.220000  1.835000 1260.390000 2.635000 ;
      RECT 1260.560000  1.835000 1261.435000 2.005000 ;
      RECT 1260.560000  2.005000 1260.940000 2.465000 ;
      RECT 1260.565000  0.995000 1260.785000 1.495000 ;
      RECT 1260.690000  0.385000 1260.860000 0.655000 ;
      RECT 1260.690000  0.655000 1261.435000 0.825000 ;
      RECT 1260.955000  0.825000 1261.435000 1.835000 ;
      RECT 1261.030000  0.085000 1261.410000 0.485000 ;
      RECT 1261.160000  2.175000 1261.330000 2.635000 ;
      RECT 1261.865000  0.085000 1262.155000 0.810000 ;
      RECT 1261.865000  1.470000 1262.155000 2.635000 ;
      RECT 1262.330000  0.765000 1262.585000 1.325000 ;
      RECT 1262.345000  0.085000 1262.585000 0.595000 ;
      RECT 1262.395000  1.495000 1264.005000 1.665000 ;
      RECT 1262.395000  1.665000 1262.755000 2.465000 ;
      RECT 1262.755000  0.290000 1263.135000 0.825000 ;
      RECT 1262.755000  0.825000 1262.985000 1.495000 ;
      RECT 1263.155000  0.995000 1263.580000 1.325000 ;
      RECT 1263.400000  0.085000 1263.570000 0.825000 ;
      RECT 1263.400000  1.835000 1263.570000 2.635000 ;
      RECT 1263.750000  1.075000 1264.860000 1.245000 ;
      RECT 1263.750000  1.245000 1264.005000 1.495000 ;
      RECT 1263.830000  0.265000 1264.210000 0.735000 ;
      RECT 1263.830000  0.735000 1265.410000 0.905000 ;
      RECT 1263.830000  1.835000 1265.150000 2.005000 ;
      RECT 1263.830000  2.005000 1264.210000 2.465000 ;
      RECT 1264.380000  0.085000 1264.550000 0.565000 ;
      RECT 1264.380000  2.175000 1264.550000 2.635000 ;
      RECT 1264.770000  0.265000 1265.150000 0.735000 ;
      RECT 1264.770000  1.495000 1265.410000 1.665000 ;
      RECT 1264.770000  1.665000 1265.150000 1.835000 ;
      RECT 1264.770000  2.005000 1265.150000 2.465000 ;
      RECT 1265.065000  0.905000 1265.410000 1.495000 ;
      RECT 1265.320000  0.085000 1265.490000 0.565000 ;
      RECT 1265.320000  1.835000 1265.490000 2.635000 ;
      RECT 1266.005000  0.085000 1266.295000 0.810000 ;
      RECT 1266.005000  1.470000 1266.295000 2.635000 ;
      RECT 1266.470000  1.075000 1266.805000 1.325000 ;
      RECT 1266.470000  1.495000 1266.725000 2.635000 ;
      RECT 1266.490000  0.265000 1266.800000 0.735000 ;
      RECT 1266.490000  0.735000 1267.275000 0.905000 ;
      RECT 1266.920000  2.085000 1268.215000 2.415000 ;
      RECT 1267.020000  0.085000 1267.755000 0.565000 ;
      RECT 1267.025000  0.905000 1267.275000 0.995000 ;
      RECT 1267.025000  0.995000 1267.765000 1.325000 ;
      RECT 1267.025000  1.325000 1267.195000 1.885000 ;
      RECT 1267.420000  1.495000 1268.765000 1.665000 ;
      RECT 1267.420000  1.665000 1267.840000 1.915000 ;
      RECT 1267.975000  0.305000 1268.145000 0.655000 ;
      RECT 1267.975000  0.655000 1268.765000 0.825000 ;
      RECT 1268.315000  0.085000 1268.745000 0.485000 ;
      RECT 1268.445000  1.835000 1268.725000 2.635000 ;
      RECT 1268.595000  0.825000 1268.765000 0.995000 ;
      RECT 1268.595000  0.995000 1268.825000 1.325000 ;
      RECT 1268.595000  1.325000 1268.765000 1.495000 ;
      RECT 1268.985000  0.415000 1269.470000 0.760000 ;
      RECT 1268.985000  1.495000 1269.470000 2.465000 ;
      RECT 1269.085000  0.760000 1269.470000 1.495000 ;
      RECT 1269.685000  0.085000 1269.975000 0.810000 ;
      RECT 1269.685000  1.470000 1269.975000 2.635000 ;
      RECT 1270.145000  1.075000 1270.485000 1.325000 ;
      RECT 1270.145000  1.495000 1270.405000 2.635000 ;
      RECT 1270.165000  0.265000 1270.480000 0.735000 ;
      RECT 1270.165000  0.735000 1270.950000 0.905000 ;
      RECT 1270.600000  2.085000 1271.890000 2.415000 ;
      RECT 1270.700000  0.085000 1271.430000 0.565000 ;
      RECT 1270.705000  0.905000 1270.950000 0.995000 ;
      RECT 1270.705000  0.995000 1271.440000 1.325000 ;
      RECT 1270.705000  1.325000 1270.875000 1.885000 ;
      RECT 1271.095000  1.495000 1272.500000 1.665000 ;
      RECT 1271.095000  1.665000 1271.515000 1.915000 ;
      RECT 1271.650000  0.305000 1271.820000 0.655000 ;
      RECT 1271.650000  0.655000 1272.500000 0.825000 ;
      RECT 1272.090000  0.085000 1272.420000 0.485000 ;
      RECT 1272.120000  1.835000 1272.400000 2.635000 ;
      RECT 1272.330000  0.825000 1272.500000 1.495000 ;
      RECT 1272.850000  0.415000 1273.170000 2.465000 ;
      RECT 1273.345000  0.085000 1273.580000 0.925000 ;
      RECT 1273.345000  1.460000 1273.580000 2.635000 ;
      RECT 1273.825000  0.085000 1274.115000 0.810000 ;
      RECT 1273.825000  1.470000 1274.115000 2.635000 ;
      RECT 1274.290000  1.075000 1274.625000 1.955000 ;
      RECT 1274.290000  2.125000 1274.545000 2.635000 ;
      RECT 1274.310000  0.265000 1274.620000 0.735000 ;
      RECT 1274.310000  0.735000 1275.095000 0.905000 ;
      RECT 1274.840000  0.085000 1275.495000 0.565000 ;
      RECT 1274.845000  0.905000 1275.095000 0.995000 ;
      RECT 1274.845000  0.995000 1275.370000 1.325000 ;
      RECT 1274.845000  1.325000 1275.015000 2.465000 ;
      RECT 1275.240000  1.495000 1277.060000 1.615000 ;
      RECT 1275.240000  1.615000 1275.760000 2.465000 ;
      RECT 1275.540000  0.735000 1276.045000 0.905000 ;
      RECT 1275.540000  0.905000 1275.760000 1.445000 ;
      RECT 1275.540000  1.445000 1277.060000 1.495000 ;
      RECT 1275.665000  0.305000 1276.045000 0.735000 ;
      RECT 1275.930000  1.075000 1276.670000 1.275000 ;
      RECT 1276.265000  1.835000 1276.545000 2.635000 ;
      RECT 1276.330000  0.085000 1276.505000 0.905000 ;
      RECT 1276.675000  0.290000 1277.055000 0.735000 ;
      RECT 1276.675000  0.735000 1278.690000 0.905000 ;
      RECT 1276.765000  1.785000 1277.955000 1.955000 ;
      RECT 1276.765000  1.955000 1277.015000 2.465000 ;
      RECT 1276.890000  1.075000 1278.000000 1.245000 ;
      RECT 1276.890000  1.245000 1277.060000 1.445000 ;
      RECT 1277.235000  2.135000 1277.485000 2.635000 ;
      RECT 1277.275000  0.085000 1277.445000 0.550000 ;
      RECT 1277.280000  1.445000 1278.690000 1.615000 ;
      RECT 1277.280000  1.615000 1277.955000 1.785000 ;
      RECT 1277.615000  0.290000 1277.995000 0.735000 ;
      RECT 1277.705000  1.955000 1277.955000 2.465000 ;
      RECT 1278.175000  1.795000 1278.425000 2.635000 ;
      RECT 1278.215000  0.085000 1278.385000 0.550000 ;
      RECT 1278.305000  0.905000 1278.690000 1.445000 ;
      RECT 1278.885000  0.085000 1279.175000 0.810000 ;
      RECT 1278.885000  1.470000 1279.175000 2.635000 ;
      RECT 1279.345000  0.995000 1279.690000 1.325000 ;
      RECT 1279.345000  2.125000 1280.635000 2.415000 ;
      RECT 1279.360000  0.305000 1279.615000 0.655000 ;
      RECT 1279.360000  0.655000 1281.235000 0.825000 ;
      RECT 1279.365000  1.495000 1279.690000 1.785000 ;
      RECT 1279.365000  1.785000 1280.635000 1.955000 ;
      RECT 1279.785000  0.085000 1280.165000 0.485000 ;
      RECT 1279.865000  0.995000 1280.750000 1.325000 ;
      RECT 1279.865000  1.325000 1280.105000 1.615000 ;
      RECT 1280.385000  0.305000 1280.555000 0.655000 ;
      RECT 1280.465000  1.495000 1281.235000 1.665000 ;
      RECT 1280.465000  1.665000 1280.635000 1.785000 ;
      RECT 1280.725000  0.085000 1281.155000 0.485000 ;
      RECT 1280.855000  1.835000 1281.135000 2.635000 ;
      RECT 1281.065000  0.825000 1281.235000 1.495000 ;
      RECT 1281.600000  0.415000 1281.875000 0.760000 ;
      RECT 1281.600000  1.495000 1281.875000 2.465000 ;
      RECT 1281.705000  0.760000 1281.875000 1.495000 ;
      RECT 1282.105000  0.085000 1282.395000 0.810000 ;
      RECT 1282.105000  1.470000 1282.395000 2.635000 ;
      RECT 1282.565000  0.995000 1282.865000 1.325000 ;
      RECT 1282.565000  2.125000 1283.860000 2.415000 ;
      RECT 1282.585000  0.305000 1282.840000 0.655000 ;
      RECT 1282.585000  0.655000 1284.590000 0.825000 ;
      RECT 1282.585000  1.495000 1282.865000 1.785000 ;
      RECT 1282.585000  1.785000 1283.850000 1.955000 ;
      RECT 1283.010000  0.085000 1283.390000 0.485000 ;
      RECT 1283.035000  0.995000 1284.060000 1.325000 ;
      RECT 1283.035000  1.325000 1283.360000 1.615000 ;
      RECT 1283.610000  0.305000 1283.780000 0.655000 ;
      RECT 1283.680000  1.495000 1284.590000 1.665000 ;
      RECT 1283.680000  1.665000 1283.850000 1.785000 ;
      RECT 1283.950000  0.085000 1284.570000 0.485000 ;
      RECT 1284.080000  1.835000 1284.550000 2.635000 ;
      RECT 1284.370000  0.825000 1284.590000 0.995000 ;
      RECT 1284.370000  0.995000 1284.780000 1.325000 ;
      RECT 1284.370000  1.325000 1284.590000 1.495000 ;
      RECT 1284.810000  0.415000 1285.135000 0.760000 ;
      RECT 1284.810000  1.495000 1285.135000 2.465000 ;
      RECT 1284.950000  0.760000 1285.135000 1.495000 ;
      RECT 1285.305000  0.085000 1285.595000 0.915000 ;
      RECT 1285.305000  1.430000 1285.595000 2.635000 ;
      RECT 1285.785000  0.085000 1286.075000 0.810000 ;
      RECT 1285.785000  1.470000 1286.075000 2.635000 ;
      RECT 1286.245000  0.255000 1286.585000 0.725000 ;
      RECT 1286.245000  0.725000 1288.400000 0.905000 ;
      RECT 1286.245000  1.075000 1286.585000 1.325000 ;
      RECT 1286.245000  1.495000 1286.585000 2.295000 ;
      RECT 1286.245000  2.295000 1287.525000 2.465000 ;
      RECT 1286.755000  1.075000 1287.315000 1.325000 ;
      RECT 1286.755000  1.325000 1286.990000 2.050000 ;
      RECT 1286.805000  0.085000 1286.975000 0.555000 ;
      RECT 1287.145000  0.255000 1287.525000 0.725000 ;
      RECT 1287.260000  1.495000 1288.400000 1.665000 ;
      RECT 1287.260000  1.665000 1287.525000 2.295000 ;
      RECT 1287.485000  1.075000 1288.010000 1.325000 ;
      RECT 1287.745000  0.085000 1288.445000 0.555000 ;
      RECT 1287.745000  1.835000 1288.445000 2.635000 ;
      RECT 1288.180000  0.905000 1288.400000 1.075000 ;
      RECT 1288.180000  1.075000 1290.105000 1.245000 ;
      RECT 1288.180000  1.245000 1288.400000 1.495000 ;
      RECT 1288.615000  0.265000 1288.995000 0.735000 ;
      RECT 1288.615000  0.735000 1290.615000 0.905000 ;
      RECT 1288.705000  1.445000 1290.615000 1.615000 ;
      RECT 1288.705000  1.615000 1288.955000 2.465000 ;
      RECT 1289.175000  1.795000 1289.425000 2.635000 ;
      RECT 1289.215000  0.085000 1289.385000 0.555000 ;
      RECT 1289.555000  0.265000 1289.935000 0.735000 ;
      RECT 1289.645000  1.615000 1289.895000 2.465000 ;
      RECT 1290.115000  1.795000 1290.365000 2.635000 ;
      RECT 1290.155000  0.085000 1290.325000 0.555000 ;
      RECT 1290.275000  0.905000 1290.615000 1.445000 ;
      RECT 1290.845000  0.085000 1291.135000 0.810000 ;
      RECT 1290.845000  1.470000 1291.135000 2.635000 ;
      RECT 1291.305000  0.085000 1291.565000 0.905000 ;
      RECT 1291.305000  1.495000 1291.565000 2.635000 ;
      RECT 1291.310000  1.075000 1291.645000 1.325000 ;
      RECT 1291.735000  0.485000 1292.115000 0.905000 ;
      RECT 1291.855000  2.125000 1293.570000 2.455000 ;
      RECT 1291.865000  0.905000 1292.115000 0.995000 ;
      RECT 1291.865000  0.995000 1292.490000 1.325000 ;
      RECT 1291.865000  1.325000 1292.035000 1.885000 ;
      RECT 1292.295000  0.255000 1292.555000 0.655000 ;
      RECT 1292.295000  0.655000 1294.110000 0.825000 ;
      RECT 1292.295000  1.495000 1292.555000 1.785000 ;
      RECT 1292.295000  1.785000 1293.570000 1.955000 ;
      RECT 1292.725000  0.085000 1293.105000 0.485000 ;
      RECT 1292.745000  0.995000 1293.685000 1.325000 ;
      RECT 1292.745000  1.325000 1292.990000 1.615000 ;
      RECT 1293.325000  0.305000 1293.495000 0.655000 ;
      RECT 1293.400000  1.495000 1294.110000 1.665000 ;
      RECT 1293.400000  1.665000 1293.570000 1.785000 ;
      RECT 1293.665000  0.085000 1294.090000 0.485000 ;
      RECT 1293.790000  1.835000 1294.070000 2.635000 ;
      RECT 1293.940000  0.825000 1294.110000 0.995000 ;
      RECT 1293.940000  0.995000 1294.215000 1.325000 ;
      RECT 1293.940000  1.325000 1294.110000 1.495000 ;
      RECT 1294.330000  0.415000 1294.755000 0.760000 ;
      RECT 1294.330000  1.495000 1294.755000 2.465000 ;
      RECT 1294.435000  0.760000 1294.755000 1.495000 ;
      RECT 1294.985000  0.085000 1295.275000 0.810000 ;
      RECT 1294.985000  1.470000 1295.275000 2.635000 ;
      RECT 1295.445000  0.290000 1295.705000 0.735000 ;
      RECT 1295.445000  0.735000 1296.175000 0.905000 ;
      RECT 1295.445000  1.075000 1295.785000 1.640000 ;
      RECT 1295.445000  1.810000 1296.175000 1.870000 ;
      RECT 1295.445000  1.870000 1298.380000 1.955000 ;
      RECT 1295.445000  1.955000 1297.340000 2.040000 ;
      RECT 1295.445000  2.040000 1295.705000 2.220000 ;
      RECT 1295.960000  2.210000 1296.320000 2.635000 ;
      RECT 1296.005000  0.085000 1296.175000 0.565000 ;
      RECT 1296.005000  0.905000 1296.175000 1.810000 ;
      RECT 1296.345000  0.265000 1296.745000 0.595000 ;
      RECT 1296.345000  0.595000 1296.595000 1.495000 ;
      RECT 1296.345000  1.495000 1296.790000 1.700000 ;
      RECT 1296.845000  0.735000 1298.905000 0.825000 ;
      RECT 1296.845000  0.825000 1297.895000 0.905000 ;
      RECT 1296.845000  0.905000 1297.015000 1.325000 ;
      RECT 1297.045000  2.210000 1297.375000 2.635000 ;
      RECT 1297.170000  1.785000 1298.380000 1.870000 ;
      RECT 1297.225000  0.085000 1297.395000 0.565000 ;
      RECT 1297.315000  1.075000 1297.900000 1.615000 ;
      RECT 1297.555000  2.125000 1298.905000 2.365000 ;
      RECT 1297.725000  0.305000 1297.895000 0.655000 ;
      RECT 1297.725000  0.655000 1298.905000 0.735000 ;
      RECT 1298.100000  0.085000 1298.430000 0.485000 ;
      RECT 1298.210000  0.995000 1298.560000 1.325000 ;
      RECT 1298.210000  1.325000 1298.380000 1.785000 ;
      RECT 1298.600000  0.305000 1298.905000 0.655000 ;
      RECT 1298.600000  1.495000 1298.905000 1.925000 ;
      RECT 1298.735000  0.825000 1298.905000 1.495000 ;
      RECT 1299.125000  0.085000 1299.415000 0.810000 ;
      RECT 1299.125000  1.470000 1299.415000 2.635000 ;
      RECT 1299.585000  0.290000 1299.845000 0.735000 ;
      RECT 1299.585000  0.735000 1300.315000 0.905000 ;
      RECT 1299.585000  1.075000 1299.925000 1.640000 ;
      RECT 1299.585000  1.810000 1300.315000 1.870000 ;
      RECT 1299.585000  1.870000 1303.530000 2.040000 ;
      RECT 1299.585000  2.040000 1299.845000 2.220000 ;
      RECT 1300.100000  2.210000 1300.460000 2.635000 ;
      RECT 1300.145000  0.905000 1300.315000 1.810000 ;
      RECT 1300.170000  0.085000 1300.340000 0.565000 ;
      RECT 1300.510000  0.285000 1300.930000 0.735000 ;
      RECT 1300.510000  0.735000 1301.740000 0.905000 ;
      RECT 1300.510000  0.905000 1300.770000 1.415000 ;
      RECT 1300.510000  1.415000 1301.920000 1.700000 ;
      RECT 1300.940000  1.075000 1302.115000 1.245000 ;
      RECT 1301.020000  2.210000 1301.400000 2.635000 ;
      RECT 1301.150000  0.085000 1301.320000 0.565000 ;
      RECT 1301.505000  0.255000 1301.740000 0.735000 ;
      RECT 1301.945000  0.655000 1303.955000 0.825000 ;
      RECT 1301.945000  0.825000 1302.115000 1.075000 ;
      RECT 1301.955000  2.210000 1302.345000 2.635000 ;
      RECT 1301.960000  0.085000 1302.340000 0.485000 ;
      RECT 1302.300000  0.995000 1302.610000 1.700000 ;
      RECT 1302.830000  0.995000 1303.070000 1.700000 ;
      RECT 1302.900000  0.085000 1303.340000 0.485000 ;
      RECT 1303.360000  0.995000 1303.530000 1.870000 ;
      RECT 1303.370000  2.210000 1303.955000 2.425000 ;
      RECT 1303.750000  0.825000 1303.955000 2.210000 ;
      RECT 1304.185000  0.085000 1304.475000 0.810000 ;
      RECT 1304.185000  1.470000 1304.475000 2.635000 ;
      RECT 1304.650000  0.755000 1305.000000 1.325000 ;
      RECT 1304.650000  1.495000 1304.970000 1.785000 ;
      RECT 1304.650000  1.785000 1306.390000 1.955000 ;
      RECT 1304.650000  2.125000 1306.455000 2.415000 ;
      RECT 1304.655000  0.085000 1304.985000 0.585000 ;
      RECT 1305.220000  0.995000 1305.915000 1.615000 ;
      RECT 1305.235000  0.305000 1305.405000 0.655000 ;
      RECT 1305.235000  0.655000 1306.995000 0.825000 ;
      RECT 1305.605000  0.085000 1305.985000 0.485000 ;
      RECT 1306.085000  0.995000 1306.655000 1.325000 ;
      RECT 1306.205000  0.305000 1306.375000 0.655000 ;
      RECT 1306.220000  1.495000 1306.995000 1.665000 ;
      RECT 1306.220000  1.665000 1306.390000 1.785000 ;
      RECT 1306.545000  0.085000 1306.975000 0.485000 ;
      RECT 1306.675000  1.835000 1306.955000 2.635000 ;
      RECT 1306.825000  0.825000 1306.995000 0.995000 ;
      RECT 1306.825000  0.995000 1307.115000 1.325000 ;
      RECT 1306.825000  1.325000 1306.995000 1.495000 ;
      RECT 1307.365000  0.415000 1307.635000 0.760000 ;
      RECT 1307.365000  1.495000 1307.635000 2.465000 ;
      RECT 1307.465000  0.760000 1307.635000 1.495000 ;
      RECT 1307.865000  0.085000 1308.155000 0.810000 ;
      RECT 1307.865000  1.470000 1308.155000 2.635000 ;
      RECT 1308.325000  0.755000 1308.675000 1.325000 ;
      RECT 1308.325000  1.495000 1308.650000 1.785000 ;
      RECT 1308.325000  1.785000 1310.070000 1.955000 ;
      RECT 1308.325000  2.125000 1310.135000 2.415000 ;
      RECT 1308.330000  0.085000 1308.665000 0.585000 ;
      RECT 1308.845000  0.995000 1309.545000 1.615000 ;
      RECT 1308.915000  0.305000 1309.085000 0.655000 ;
      RECT 1308.915000  0.655000 1310.675000 0.825000 ;
      RECT 1309.285000  0.085000 1309.665000 0.485000 ;
      RECT 1309.715000  0.995000 1310.335000 1.325000 ;
      RECT 1309.885000  0.305000 1310.055000 0.655000 ;
      RECT 1309.900000  1.495000 1310.675000 1.665000 ;
      RECT 1309.900000  1.665000 1310.070000 1.785000 ;
      RECT 1310.225000  0.085000 1310.655000 0.485000 ;
      RECT 1310.355000  1.835000 1310.635000 2.635000 ;
      RECT 1310.505000  0.825000 1310.675000 0.995000 ;
      RECT 1310.505000  0.995000 1310.940000 1.325000 ;
      RECT 1310.505000  1.325000 1310.675000 1.495000 ;
      RECT 1311.060000  0.415000 1311.365000 0.760000 ;
      RECT 1311.060000  1.495000 1311.365000 2.465000 ;
      RECT 1311.130000  0.760000 1311.365000 1.495000 ;
      RECT 1311.555000  0.085000 1311.775000 1.000000 ;
      RECT 1311.555000  1.455000 1311.775000 2.635000 ;
      RECT 1312.005000  0.085000 1312.295000 0.810000 ;
      RECT 1312.005000  1.470000 1312.295000 2.635000 ;
      RECT 1312.465000  0.755000 1312.750000 1.325000 ;
      RECT 1312.495000  1.495000 1313.140000 1.665000 ;
      RECT 1312.495000  1.665000 1312.830000 2.450000 ;
      RECT 1312.500000  0.085000 1312.750000 0.585000 ;
      RECT 1312.920000  0.655000 1314.930000 0.825000 ;
      RECT 1312.920000  0.825000 1313.140000 1.495000 ;
      RECT 1313.130000  0.305000 1313.300000 0.655000 ;
      RECT 1313.310000  0.995000 1313.480000 1.620000 ;
      RECT 1313.310000  1.620000 1313.710000 2.375000 ;
      RECT 1313.500000  0.085000 1313.880000 0.485000 ;
      RECT 1313.760000  0.995000 1314.140000 1.450000 ;
      RECT 1313.880000  1.450000 1314.140000 1.785000 ;
      RECT 1313.880000  1.785000 1314.250000 2.375000 ;
      RECT 1314.100000  0.305000 1314.270000 0.655000 ;
      RECT 1314.320000  0.995000 1314.590000 1.445000 ;
      RECT 1314.320000  1.445000 1314.855000 1.615000 ;
      RECT 1314.540000  0.085000 1314.920000 0.485000 ;
      RECT 1314.585000  1.795000 1314.835000 2.635000 ;
      RECT 1314.760000  0.825000 1314.930000 1.075000 ;
      RECT 1314.760000  1.075000 1316.370000 1.245000 ;
      RECT 1315.110000  1.455000 1316.865000 1.625000 ;
      RECT 1315.110000  1.625000 1315.360000 2.465000 ;
      RECT 1315.150000  0.255000 1315.400000 0.725000 ;
      RECT 1315.150000  0.725000 1316.865000 0.905000 ;
      RECT 1315.580000  1.795000 1315.830000 2.635000 ;
      RECT 1315.620000  0.085000 1315.790000 0.555000 ;
      RECT 1315.960000  0.255000 1316.340000 0.725000 ;
      RECT 1316.050000  1.625000 1316.300000 2.465000 ;
      RECT 1316.520000  1.795000 1316.770000 2.635000 ;
      RECT 1316.560000  0.085000 1316.730000 0.555000 ;
      RECT 1316.590000  0.905000 1316.865000 1.455000 ;
      RECT 1317.065000  0.085000 1317.355000 0.810000 ;
      RECT 1317.065000  1.470000 1317.355000 2.635000 ;
      RECT 1317.525000  0.085000 1317.865000 0.585000 ;
      RECT 1317.525000  0.755000 1317.865000 1.325000 ;
      RECT 1317.525000  1.560000 1317.865000 2.635000 ;
      RECT 1318.085000  0.305000 1318.330000 0.995000 ;
      RECT 1318.085000  0.995000 1318.740000 1.325000 ;
      RECT 1318.085000  1.325000 1318.325000 1.920000 ;
      RECT 1318.100000  2.125000 1320.300000 2.415000 ;
      RECT 1318.520000  1.495000 1318.840000 1.785000 ;
      RECT 1318.520000  1.785000 1320.300000 1.955000 ;
      RECT 1318.525000  0.085000 1318.855000 0.585000 ;
      RECT 1319.060000  0.995000 1319.850000 1.615000 ;
      RECT 1319.105000  0.305000 1319.275000 0.655000 ;
      RECT 1319.105000  0.655000 1320.855000 0.825000 ;
      RECT 1319.450000  0.085000 1319.830000 0.485000 ;
      RECT 1320.050000  0.305000 1320.220000 0.655000 ;
      RECT 1320.070000  0.995000 1320.515000 1.325000 ;
      RECT 1320.130000  1.495000 1320.855000 1.665000 ;
      RECT 1320.130000  1.665000 1320.300000 1.785000 ;
      RECT 1320.390000  0.085000 1320.820000 0.485000 ;
      RECT 1320.520000  1.835000 1320.800000 2.635000 ;
      RECT 1320.685000  0.825000 1320.855000 0.995000 ;
      RECT 1320.685000  0.995000 1320.945000 1.325000 ;
      RECT 1320.685000  1.325000 1320.855000 1.495000 ;
      RECT 1321.060000  0.415000 1321.435000 0.760000 ;
      RECT 1321.060000  1.495000 1321.435000 2.465000 ;
      RECT 1321.165000  0.760000 1321.435000 1.495000 ;
      RECT 1321.665000  0.085000 1321.955000 0.810000 ;
      RECT 1321.665000  1.470000 1321.955000 2.635000 ;
      RECT 1322.125000  0.325000 1322.390000 0.735000 ;
      RECT 1322.125000  0.735000 1322.855000 0.905000 ;
      RECT 1322.125000  1.075000 1322.465000 1.435000 ;
      RECT 1322.125000  1.605000 1322.855000 1.890000 ;
      RECT 1322.550000  1.890000 1322.855000 1.995000 ;
      RECT 1322.550000  1.995000 1323.905000 2.165000 ;
      RECT 1322.555000  2.335000 1322.935000 2.635000 ;
      RECT 1322.685000  0.905000 1322.855000 1.605000 ;
      RECT 1322.720000  0.085000 1322.890000 0.565000 ;
      RECT 1323.060000  0.260000 1323.390000 0.790000 ;
      RECT 1323.060000  0.790000 1323.275000 1.495000 ;
      RECT 1323.060000  1.495000 1323.390000 1.825000 ;
      RECT 1323.445000  0.960000 1323.775000 1.325000 ;
      RECT 1323.560000  1.325000 1323.775000 1.445000 ;
      RECT 1323.560000  1.445000 1325.950000 1.615000 ;
      RECT 1323.575000  0.085000 1324.005000 0.485000 ;
      RECT 1323.580000  1.785000 1325.370000 1.955000 ;
      RECT 1323.580000  1.955000 1323.905000 1.995000 ;
      RECT 1323.605000  0.700000 1325.345000 0.870000 ;
      RECT 1323.605000  0.870000 1323.775000 0.960000 ;
      RECT 1323.670000  2.335000 1324.005000 2.635000 ;
      RECT 1323.945000  1.075000 1324.560000 1.275000 ;
      RECT 1324.225000  0.270000 1324.395000 0.700000 ;
      RECT 1324.225000  2.125000 1324.960000 2.415000 ;
      RECT 1324.625000  0.085000 1324.955000 0.485000 ;
      RECT 1324.840000  1.075000 1325.940000 1.275000 ;
      RECT 1325.175000  0.270000 1325.345000 0.700000 ;
      RECT 1325.200000  1.955000 1325.370000 2.215000 ;
      RECT 1325.200000  2.215000 1325.735000 2.385000 ;
      RECT 1325.565000  0.085000 1325.945000 0.585000 ;
      RECT 1325.565000  1.615000 1325.950000 1.780000 ;
      RECT 1326.265000  0.085000 1326.555000 0.810000 ;
      RECT 1326.265000  1.470000 1326.555000 2.635000 ;
      RECT 1326.725000  0.085000 1326.985000 0.825000 ;
      RECT 1326.725000  2.135000 1327.005000 2.635000 ;
      RECT 1326.745000  0.995000 1327.085000 1.955000 ;
      RECT 1327.285000  0.435000 1327.475000 0.995000 ;
      RECT 1327.285000  0.995000 1327.905000 1.325000 ;
      RECT 1327.285000  1.325000 1327.475000 2.455000 ;
      RECT 1327.725000  0.085000 1327.975000 0.585000 ;
      RECT 1327.725000  1.575000 1328.365000 1.745000 ;
      RECT 1327.725000  1.745000 1328.055000 2.450000 ;
      RECT 1328.145000  0.655000 1330.155000 0.825000 ;
      RECT 1328.145000  0.825000 1328.365000 1.575000 ;
      RECT 1328.355000  0.305000 1328.525000 0.655000 ;
      RECT 1328.535000  0.995000 1328.825000 2.375000 ;
      RECT 1328.725000  0.085000 1329.105000 0.485000 ;
      RECT 1329.015000  0.995000 1329.345000 2.375000 ;
      RECT 1329.325000  0.305000 1329.495000 0.655000 ;
      RECT 1329.515000  0.995000 1329.815000 1.445000 ;
      RECT 1329.515000  1.445000 1330.080000 1.615000 ;
      RECT 1329.765000  0.085000 1330.145000 0.485000 ;
      RECT 1329.810000  1.795000 1330.060000 2.635000 ;
      RECT 1329.985000  0.825000 1330.155000 1.075000 ;
      RECT 1329.985000  1.075000 1331.595000 1.245000 ;
      RECT 1330.335000  1.455000 1332.055000 1.625000 ;
      RECT 1330.335000  1.625000 1330.585000 2.465000 ;
      RECT 1330.375000  0.255000 1330.625000 0.725000 ;
      RECT 1330.375000  0.725000 1332.055000 0.905000 ;
      RECT 1330.805000  1.795000 1331.055000 2.635000 ;
      RECT 1330.845000  0.085000 1331.015000 0.555000 ;
      RECT 1331.185000  0.255000 1331.565000 0.725000 ;
      RECT 1331.275000  1.625000 1331.525000 2.465000 ;
      RECT 1331.745000  1.795000 1331.995000 2.635000 ;
      RECT 1331.785000  0.085000 1331.955000 0.555000 ;
      RECT 1331.815000  0.905000 1332.055000 1.455000 ;
      RECT 1332.245000  0.085000 1332.535000 0.810000 ;
      RECT 1332.245000  1.470000 1332.535000 2.635000 ;
      RECT 1332.705000  0.450000 1333.020000 0.825000 ;
      RECT 1332.705000  0.825000 1332.875000 1.865000 ;
      RECT 1332.705000  1.865000 1334.635000 2.035000 ;
      RECT 1332.705000  2.035000 1332.965000 2.455000 ;
      RECT 1333.045000  0.995000 1333.430000 1.695000 ;
      RECT 1333.135000  2.205000 1333.515000 2.635000 ;
      RECT 1333.325000  0.085000 1333.495000 0.825000 ;
      RECT 1333.600000  0.995000 1333.955000 1.325000 ;
      RECT 1333.660000  1.525000 1334.295000 1.695000 ;
      RECT 1333.795000  0.450000 1333.965000 0.655000 ;
      RECT 1333.795000  0.655000 1334.295000 0.825000 ;
      RECT 1334.125000  0.825000 1334.295000 1.075000 ;
      RECT 1334.125000  1.075000 1334.775000 1.245000 ;
      RECT 1334.125000  1.245000 1334.295000 1.525000 ;
      RECT 1334.190000  0.085000 1334.565000 0.485000 ;
      RECT 1334.230000  2.205000 1335.025000 2.375000 ;
      RECT 1334.465000  1.415000 1335.165000 1.585000 ;
      RECT 1334.465000  1.585000 1334.635000 1.865000 ;
      RECT 1334.785000  0.305000 1334.955000 0.655000 ;
      RECT 1334.785000  0.655000 1336.530000 0.825000 ;
      RECT 1334.855000  1.785000 1335.990000 1.955000 ;
      RECT 1334.855000  1.955000 1335.025000 2.205000 ;
      RECT 1334.995000  0.995000 1335.165000 1.415000 ;
      RECT 1335.140000  0.085000 1335.520000 0.485000 ;
      RECT 1335.300000  2.125000 1335.990000 2.455000 ;
      RECT 1335.435000  0.995000 1336.190000 1.325000 ;
      RECT 1335.740000  0.305000 1335.910000 0.655000 ;
      RECT 1335.820000  1.495000 1336.530000 1.665000 ;
      RECT 1335.820000  1.665000 1335.990000 1.785000 ;
      RECT 1336.080000  0.085000 1336.510000 0.485000 ;
      RECT 1336.210000  1.835000 1336.490000 2.635000 ;
      RECT 1336.360000  0.825000 1336.530000 0.995000 ;
      RECT 1336.360000  0.995000 1336.650000 1.325000 ;
      RECT 1336.360000  1.325000 1336.530000 1.495000 ;
      RECT 1336.750000  0.415000 1337.075000 0.760000 ;
      RECT 1336.750000  1.495000 1337.075000 2.465000 ;
      RECT 1336.855000  0.760000 1337.075000 1.495000 ;
      RECT 1337.305000  0.085000 1337.595000 0.810000 ;
      RECT 1337.305000  1.470000 1337.595000 2.635000 ;
      RECT 1337.765000  0.450000 1338.085000 0.825000 ;
      RECT 1337.765000  0.825000 1337.940000 1.865000 ;
      RECT 1337.765000  1.865000 1339.720000 2.035000 ;
      RECT 1337.765000  2.035000 1338.025000 2.455000 ;
      RECT 1338.110000  0.995000 1338.510000 1.695000 ;
      RECT 1338.195000  2.205000 1338.575000 2.635000 ;
      RECT 1338.390000  0.085000 1338.560000 0.825000 ;
      RECT 1338.680000  0.995000 1339.020000 1.325000 ;
      RECT 1338.725000  1.525000 1339.380000 1.695000 ;
      RECT 1338.860000  0.450000 1339.030000 0.655000 ;
      RECT 1338.860000  0.655000 1339.380000 0.825000 ;
      RECT 1339.190000  0.825000 1339.380000 1.075000 ;
      RECT 1339.190000  1.075000 1339.635000 1.245000 ;
      RECT 1339.190000  1.245000 1339.380000 1.525000 ;
      RECT 1339.275000  0.085000 1339.650000 0.485000 ;
      RECT 1339.315000  2.205000 1340.110000 2.375000 ;
      RECT 1339.550000  1.415000 1340.250000 1.585000 ;
      RECT 1339.550000  1.585000 1339.720000 1.865000 ;
      RECT 1339.870000  0.305000 1340.040000 0.655000 ;
      RECT 1339.870000  0.655000 1341.615000 0.825000 ;
      RECT 1339.940000  1.785000 1341.075000 1.955000 ;
      RECT 1339.940000  1.955000 1340.110000 2.205000 ;
      RECT 1340.080000  0.995000 1340.250000 1.415000 ;
      RECT 1340.225000  0.085000 1340.605000 0.485000 ;
      RECT 1340.385000  2.125000 1341.075000 2.455000 ;
      RECT 1340.520000  0.995000 1341.275000 1.325000 ;
      RECT 1340.825000  0.305000 1340.995000 0.655000 ;
      RECT 1340.905000  1.495000 1341.615000 1.665000 ;
      RECT 1340.905000  1.665000 1341.075000 1.785000 ;
      RECT 1341.165000  0.085000 1341.595000 0.485000 ;
      RECT 1341.295000  1.835000 1341.575000 2.635000 ;
      RECT 1341.445000  0.825000 1341.615000 0.995000 ;
      RECT 1341.445000  0.995000 1341.720000 1.325000 ;
      RECT 1341.445000  1.325000 1341.615000 1.495000 ;
      RECT 1341.835000  0.415000 1342.135000 0.760000 ;
      RECT 1341.835000  1.495000 1342.135000 2.465000 ;
      RECT 1341.940000  0.760000 1342.135000 1.495000 ;
      RECT 1342.330000  0.085000 1342.500000 0.915000 ;
      RECT 1342.330000  1.440000 1342.500000 2.635000 ;
      RECT 1342.825000  0.085000 1343.115000 0.810000 ;
      RECT 1342.825000  1.470000 1343.115000 2.635000 ;
      RECT 1343.295000  0.450000 1343.600000 0.825000 ;
      RECT 1343.295000  0.825000 1343.465000 1.900000 ;
      RECT 1343.295000  1.900000 1344.595000 2.070000 ;
      RECT 1343.295000  2.070000 1343.545000 2.455000 ;
      RECT 1343.635000  0.995000 1344.025000 1.695000 ;
      RECT 1343.715000  2.240000 1344.095000 2.635000 ;
      RECT 1343.905000  0.085000 1344.075000 0.825000 ;
      RECT 1344.195000  0.995000 1344.535000 1.325000 ;
      RECT 1344.240000  1.560000 1344.895000 1.730000 ;
      RECT 1344.375000  0.450000 1344.545000 0.655000 ;
      RECT 1344.375000  0.655000 1344.895000 0.825000 ;
      RECT 1344.425000  2.070000 1344.595000 2.295000 ;
      RECT 1344.425000  2.295000 1345.765000 2.465000 ;
      RECT 1344.705000  0.825000 1344.895000 0.995000 ;
      RECT 1344.705000  0.995000 1344.995000 1.325000 ;
      RECT 1344.705000  1.325000 1344.895000 1.560000 ;
      RECT 1344.810000  1.955000 1345.425000 2.125000 ;
      RECT 1344.815000  0.085000 1345.145000 0.480000 ;
      RECT 1345.235000  0.655000 1347.215000 0.825000 ;
      RECT 1345.235000  0.825000 1345.425000 1.955000 ;
      RECT 1345.445000  0.305000 1345.615000 0.655000 ;
      RECT 1345.595000  0.995000 1345.765000 2.295000 ;
      RECT 1345.785000  0.085000 1346.165000 0.485000 ;
      RECT 1346.045000  0.995000 1346.345000 2.375000 ;
      RECT 1346.385000  0.305000 1346.555000 0.655000 ;
      RECT 1346.515000  1.400000 1346.875000 1.615000 ;
      RECT 1346.655000  0.995000 1346.875000 1.400000 ;
      RECT 1346.815000  0.085000 1347.195000 0.485000 ;
      RECT 1346.860000  1.795000 1347.110000 2.635000 ;
      RECT 1347.045000  0.825000 1347.215000 1.075000 ;
      RECT 1347.045000  1.075000 1348.645000 1.245000 ;
      RECT 1347.385000  1.455000 1349.055000 1.625000 ;
      RECT 1347.385000  1.625000 1347.635000 2.465000 ;
      RECT 1347.425000  0.255000 1347.675000 0.725000 ;
      RECT 1347.425000  0.725000 1349.055000 0.905000 ;
      RECT 1347.855000  1.795000 1348.105000 2.635000 ;
      RECT 1347.895000  0.085000 1348.065000 0.555000 ;
      RECT 1348.235000  0.255000 1348.615000 0.725000 ;
      RECT 1348.325000  1.625000 1348.575000 2.465000 ;
      RECT 1348.795000  1.795000 1349.045000 2.635000 ;
      RECT 1348.825000  0.905000 1349.055000 1.455000 ;
      RECT 1348.835000  0.085000 1349.005000 0.555000 ;
      RECT 1349.265000  0.085000 1349.555000 0.810000 ;
      RECT 1349.265000  1.470000 1349.555000 2.635000 ;
      RECT 1349.725000  0.975000 1350.075000 1.625000 ;
      RECT 1349.810000  0.345000 1349.985000 0.635000 ;
      RECT 1349.810000  0.635000 1350.525000 0.805000 ;
      RECT 1349.810000  1.795000 1350.525000 1.965000 ;
      RECT 1349.810000  1.965000 1349.985000 2.465000 ;
      RECT 1350.155000  0.085000 1350.535000 0.465000 ;
      RECT 1350.155000  2.135000 1350.535000 2.635000 ;
      RECT 1350.295000  0.805000 1350.525000 1.795000 ;
      RECT 1350.755000  0.345000 1350.960000 2.465000 ;
      RECT 1351.130000  1.025000 1351.405000 1.685000 ;
      RECT 1351.195000  0.085000 1351.445000 0.635000 ;
      RECT 1351.195000  1.885000 1351.525000 2.635000 ;
      RECT 1351.575000  0.760000 1351.895000 0.765000 ;
      RECT 1351.575000  0.765000 1352.245000 1.015000 ;
      RECT 1351.575000  1.015000 1351.895000 1.695000 ;
      RECT 1351.615000  0.345000 1351.895000 0.760000 ;
      RECT 1352.025000  1.875000 1352.405000 2.385000 ;
      RECT 1352.190000  0.265000 1352.595000 0.595000 ;
      RECT 1352.190000  1.185000 1352.915000 1.365000 ;
      RECT 1352.190000  1.365000 1352.405000 1.875000 ;
      RECT 1352.425000  0.595000 1352.595000 1.075000 ;
      RECT 1352.425000  1.075000 1352.915000 1.185000 ;
      RECT 1352.585000  1.575000 1353.535000 1.745000 ;
      RECT 1352.585000  1.745000 1352.905000 1.905000 ;
      RECT 1352.735000  1.905000 1352.905000 2.465000 ;
      RECT 1352.765000  0.305000 1352.965000 0.625000 ;
      RECT 1352.765000  0.625000 1353.535000 0.765000 ;
      RECT 1352.765000  0.765000 1353.710000 0.795000 ;
      RECT 1353.150000  2.215000 1353.530000 2.635000 ;
      RECT 1353.260000  0.085000 1353.590000 0.445000 ;
      RECT 1353.365000  0.795000 1353.710000 1.095000 ;
      RECT 1353.365000  1.095000 1353.535000 1.575000 ;
      RECT 1353.795000  1.325000 1354.115000 2.375000 ;
      RECT 1354.285000  0.305000 1354.455000 2.465000 ;
      RECT 1354.625000  0.705000 1354.885000 1.575000 ;
      RECT 1354.625000  1.575000 1355.215000 1.955000 ;
      RECT 1354.675000  2.250000 1355.555000 2.420000 ;
      RECT 1354.740000  0.265000 1355.855000 0.465000 ;
      RECT 1355.065000  0.645000 1355.465000 1.015000 ;
      RECT 1355.385000  1.195000 1355.855000 1.235000 ;
      RECT 1355.385000  1.235000 1356.835000 1.405000 ;
      RECT 1355.385000  1.405000 1355.555000 2.250000 ;
      RECT 1355.635000  0.465000 1355.855000 1.195000 ;
      RECT 1355.725000  1.575000 1356.025000 1.785000 ;
      RECT 1355.725000  1.785000 1357.225000 2.035000 ;
      RECT 1355.845000  2.205000 1356.225000 2.635000 ;
      RECT 1356.025000  0.085000 1356.195000 0.525000 ;
      RECT 1356.025000  0.735000 1356.435000 1.065000 ;
      RECT 1356.415000  0.255000 1357.685000 0.425000 ;
      RECT 1356.415000  0.425000 1356.745000 0.465000 ;
      RECT 1356.575000  2.035000 1356.745000 2.375000 ;
      RECT 1356.585000  1.405000 1356.835000 1.485000 ;
      RECT 1356.615000  1.155000 1356.835000 1.235000 ;
      RECT 1356.915000  0.595000 1357.295000 0.765000 ;
      RECT 1357.055000  0.765000 1357.295000 0.895000 ;
      RECT 1357.055000  0.895000 1358.515000 1.065000 ;
      RECT 1357.055000  1.065000 1357.225000 1.785000 ;
      RECT 1357.445000  1.235000 1357.775000 1.415000 ;
      RECT 1357.445000  1.415000 1358.550000 1.655000 ;
      RECT 1357.465000  1.915000 1357.795000 2.635000 ;
      RECT 1357.490000  0.425000 1357.685000 0.715000 ;
      RECT 1357.930000  0.085000 1358.315000 0.465000 ;
      RECT 1358.085000  1.065000 1358.515000 1.235000 ;
      RECT 1358.750000  1.575000 1358.985000 1.985000 ;
      RECT 1358.810000  0.705000 1359.150000 1.125000 ;
      RECT 1358.810000  1.125000 1359.530000 1.305000 ;
      RECT 1358.940000  2.250000 1359.870000 2.420000 ;
      RECT 1359.055000  0.265000 1359.870000 0.465000 ;
      RECT 1359.275000  1.305000 1359.530000 1.905000 ;
      RECT 1359.700000  0.465000 1359.870000 1.235000 ;
      RECT 1359.700000  1.235000 1361.150000 1.405000 ;
      RECT 1359.700000  1.405000 1359.870000 2.250000 ;
      RECT 1360.040000  1.575000 1360.340000 1.915000 ;
      RECT 1360.040000  1.915000 1363.070000 2.085000 ;
      RECT 1360.050000  0.085000 1360.360000 0.525000 ;
      RECT 1360.160000  2.255000 1360.540000 2.635000 ;
      RECT 1360.295000  0.735000 1360.720000 1.065000 ;
      RECT 1360.620000  0.255000 1361.940000 0.425000 ;
      RECT 1360.620000  0.425000 1361.020000 0.465000 ;
      RECT 1360.830000  2.085000 1361.000000 2.375000 ;
      RECT 1360.930000  1.075000 1361.150000 1.235000 ;
      RECT 1361.175000  0.645000 1361.555000 0.815000 ;
      RECT 1361.370000  0.815000 1361.555000 1.915000 ;
      RECT 1361.580000  2.255000 1363.070000 2.635000 ;
      RECT 1361.765000  0.425000 1361.940000 0.585000 ;
      RECT 1361.770000  0.755000 1362.455000 0.925000 ;
      RECT 1361.770000  0.925000 1361.985000 1.575000 ;
      RECT 1361.770000  1.575000 1362.545000 1.745000 ;
      RECT 1362.155000  1.095000 1362.730000 1.325000 ;
      RECT 1362.255000  0.265000 1362.455000 0.755000 ;
      RECT 1362.740000  0.085000 1363.070000 0.805000 ;
      RECT 1362.900000  0.995000 1363.165000 1.325000 ;
      RECT 1362.900000  1.325000 1363.070000 1.915000 ;
      RECT 1363.355000  0.255000 1363.755000 0.715000 ;
      RECT 1363.355000  1.630000 1363.735000 2.465000 ;
      RECT 1363.460000  0.715000 1363.755000 1.520000 ;
      RECT 1363.460000  1.520000 1363.735000 1.630000 ;
      RECT 1363.905000  1.725000 1364.160000 2.415000 ;
      RECT 1363.955000  0.255000 1364.160000 0.995000 ;
      RECT 1363.955000  0.995000 1364.730000 1.325000 ;
      RECT 1363.955000  1.325000 1364.160000 1.725000 ;
      RECT 1364.385000  1.765000 1364.680000 2.635000 ;
      RECT 1364.390000  0.085000 1364.680000 0.545000 ;
      RECT 1364.900000  0.255000 1365.185000 0.825000 ;
      RECT 1364.900000  1.605000 1365.185000 2.465000 ;
      RECT 1364.950000  0.825000 1365.185000 1.605000 ;
      RECT 1365.365000  0.085000 1365.655000 0.810000 ;
      RECT 1365.365000  1.470000 1365.655000 2.635000 ;
      RECT 1365.830000  1.795000 1366.655000 1.965000 ;
      RECT 1365.830000  1.965000 1366.085000 2.465000 ;
      RECT 1365.835000  0.345000 1366.085000 0.635000 ;
      RECT 1365.835000  0.635000 1366.625000 0.805000 ;
      RECT 1365.880000  0.975000 1366.230000 1.625000 ;
      RECT 1366.255000  0.085000 1366.635000 0.465000 ;
      RECT 1366.270000  2.135000 1366.650000 2.635000 ;
      RECT 1366.450000  0.805000 1366.625000 0.995000 ;
      RECT 1366.450000  0.995000 1366.765000 1.325000 ;
      RECT 1366.450000  1.325000 1366.655000 1.795000 ;
      RECT 1366.855000  0.345000 1367.105000 0.675000 ;
      RECT 1366.875000  1.730000 1367.105000 2.465000 ;
      RECT 1366.935000  0.675000 1367.105000 1.730000 ;
      RECT 1367.325000  1.070000 1367.730000 1.335000 ;
      RECT 1367.325000  1.335000 1367.960000 1.745000 ;
      RECT 1367.435000  0.395000 1367.605000 0.730000 ;
      RECT 1367.435000  0.730000 1368.175000 0.900000 ;
      RECT 1367.775000  0.085000 1368.155000 0.560000 ;
      RECT 1367.850000  1.915000 1368.470000 2.085000 ;
      RECT 1367.850000  2.085000 1368.120000 2.400000 ;
      RECT 1368.005000  0.900000 1368.175000 0.995000 ;
      RECT 1368.005000  0.995000 1369.185000 1.165000 ;
      RECT 1368.215000  1.165000 1369.185000 1.185000 ;
      RECT 1368.215000  1.185000 1368.470000 1.915000 ;
      RECT 1368.340000  2.255000 1368.670000 2.635000 ;
      RECT 1368.395000  0.085000 1368.775000 0.825000 ;
      RECT 1368.860000  1.355000 1369.395000 2.465000 ;
      RECT 1369.015000  0.255000 1370.175000 0.425000 ;
      RECT 1369.015000  0.425000 1369.185000 0.995000 ;
      RECT 1369.405000  0.675000 1369.785000 1.075000 ;
      RECT 1369.610000  1.075000 1369.785000 1.935000 ;
      RECT 1369.610000  1.935000 1371.390000 2.105000 ;
      RECT 1369.610000  2.105000 1369.780000 2.465000 ;
      RECT 1370.005000  0.425000 1370.175000 1.685000 ;
      RECT 1370.350000  0.710000 1370.695000 1.700000 ;
      RECT 1370.595000  2.275000 1370.945000 2.635000 ;
      RECT 1370.745000  0.085000 1371.090000 0.540000 ;
      RECT 1370.880000  0.715000 1371.460000 0.895000 ;
      RECT 1370.880000  0.895000 1371.050000 1.935000 ;
      RECT 1371.220000  1.065000 1371.390000 1.395000 ;
      RECT 1371.220000  2.105000 1371.390000 2.185000 ;
      RECT 1371.220000  2.185000 1371.590000 2.435000 ;
      RECT 1371.290000  0.335000 1371.630000 0.505000 ;
      RECT 1371.290000  0.505000 1371.460000 0.715000 ;
      RECT 1371.560000  1.575000 1371.860000 1.955000 ;
      RECT 1371.640000  0.705000 1372.390000 1.035000 ;
      RECT 1371.640000  1.035000 1371.860000 1.575000 ;
      RECT 1371.835000  2.135000 1372.200000 2.465000 ;
      RECT 1371.850000  0.305000 1372.750000 0.475000 ;
      RECT 1372.030000  1.215000 1373.890000 1.385000 ;
      RECT 1372.030000  1.385000 1372.200000 2.135000 ;
      RECT 1372.420000  1.935000 1373.680000 2.105000 ;
      RECT 1372.420000  2.105000 1372.590000 2.375000 ;
      RECT 1372.580000  0.475000 1372.750000 1.215000 ;
      RECT 1372.700000  1.595000 1374.280000 1.765000 ;
      RECT 1372.875000  2.355000 1373.205000 2.635000 ;
      RECT 1372.970000  0.765000 1373.550000 1.045000 ;
      RECT 1373.430000  0.085000 1373.760000 0.545000 ;
      RECT 1373.510000  2.105000 1373.680000 2.375000 ;
      RECT 1373.720000  1.005000 1373.890000 1.215000 ;
      RECT 1373.890000  2.175000 1374.310000 2.635000 ;
      RECT 1373.970000  0.275000 1374.350000 0.445000 ;
      RECT 1373.970000  0.445000 1374.280000 0.835000 ;
      RECT 1373.970000  1.765000 1374.280000 1.835000 ;
      RECT 1373.970000  1.835000 1374.725000 2.005000 ;
      RECT 1374.110000  0.835000 1374.280000 1.595000 ;
      RECT 1374.450000  0.705000 1374.710000 1.495000 ;
      RECT 1374.450000  1.495000 1375.185000 1.660000 ;
      RECT 1374.450000  1.660000 1375.585000 1.665000 ;
      RECT 1374.520000  0.255000 1375.630000 0.535000 ;
      RECT 1374.555000  2.005000 1374.725000 2.465000 ;
      RECT 1374.925000  1.665000 1375.585000 1.955000 ;
      RECT 1374.935000  2.125000 1375.955000 2.465000 ;
      RECT 1374.975000  0.920000 1375.145000 1.325000 ;
      RECT 1375.410000  0.535000 1375.630000 1.315000 ;
      RECT 1375.410000  1.315000 1376.025000 1.485000 ;
      RECT 1375.780000  1.485000 1376.025000 1.575000 ;
      RECT 1375.780000  1.575000 1377.110000 1.745000 ;
      RECT 1375.780000  1.745000 1375.955000 2.125000 ;
      RECT 1375.850000  0.085000 1376.070000 0.525000 ;
      RECT 1375.890000  0.695000 1376.470000 0.865000 ;
      RECT 1375.890000  0.865000 1376.110000 1.145000 ;
      RECT 1376.155000  2.195000 1376.405000 2.635000 ;
      RECT 1376.300000  0.295000 1377.475000 0.465000 ;
      RECT 1376.300000  0.465000 1376.470000 0.695000 ;
      RECT 1376.340000  1.065000 1377.110000 1.275000 ;
      RECT 1376.650000  1.915000 1377.470000 2.085000 ;
      RECT 1376.650000  2.085000 1376.820000 2.375000 ;
      RECT 1376.805000  0.635000 1377.110000 1.065000 ;
      RECT 1376.995000  2.255000 1377.375000 2.635000 ;
      RECT 1377.300000  0.465000 1377.475000 0.995000 ;
      RECT 1377.300000  0.995000 1377.945000 1.325000 ;
      RECT 1377.300000  1.325000 1377.470000 1.915000 ;
      RECT 1377.645000  0.085000 1377.930000 0.710000 ;
      RECT 1377.645000  1.495000 1377.930000 2.635000 ;
      RECT 1378.160000  0.265000 1378.510000 2.395000 ;
      RECT 1378.680000  0.255000 1378.850000 0.635000 ;
      RECT 1378.680000  0.635000 1379.345000 0.805000 ;
      RECT 1378.680000  1.535000 1379.345000 1.705000 ;
      RECT 1378.680000  1.705000 1378.850000 2.465000 ;
      RECT 1379.025000  0.085000 1379.435000 0.465000 ;
      RECT 1379.025000  1.875000 1379.435000 2.635000 ;
      RECT 1379.175000  0.805000 1379.345000 0.995000 ;
      RECT 1379.175000  0.995000 1379.505000 1.325000 ;
      RECT 1379.175000  1.325000 1379.345000 1.535000 ;
      RECT 1379.625000  0.255000 1379.905000 0.870000 ;
      RECT 1379.625000  1.475000 1379.905000 2.465000 ;
      RECT 1379.675000  0.870000 1379.905000 1.475000 ;
      RECT 1380.085000  0.085000 1380.375000 0.810000 ;
      RECT 1380.085000  1.470000 1380.375000 2.635000 ;
      RECT 1380.550000  1.795000 1381.375000 1.965000 ;
      RECT 1380.550000  1.965000 1380.805000 2.465000 ;
      RECT 1380.555000  0.345000 1380.805000 0.635000 ;
      RECT 1380.555000  0.635000 1381.345000 0.805000 ;
      RECT 1380.600000  0.975000 1380.950000 1.625000 ;
      RECT 1380.975000  0.085000 1381.355000 0.465000 ;
      RECT 1380.990000  2.135000 1381.370000 2.635000 ;
      RECT 1381.170000  0.805000 1381.345000 0.995000 ;
      RECT 1381.170000  0.995000 1381.485000 1.325000 ;
      RECT 1381.170000  1.325000 1381.375000 1.795000 ;
      RECT 1381.575000  0.345000 1381.825000 0.675000 ;
      RECT 1381.595000  1.730000 1381.825000 2.465000 ;
      RECT 1381.655000  0.675000 1381.825000 1.730000 ;
      RECT 1382.045000  1.070000 1382.450000 1.335000 ;
      RECT 1382.045000  1.335000 1382.680000 1.745000 ;
      RECT 1382.155000  0.395000 1382.325000 0.730000 ;
      RECT 1382.155000  0.730000 1382.895000 0.900000 ;
      RECT 1382.495000  0.085000 1382.875000 0.560000 ;
      RECT 1382.570000  1.915000 1383.190000 2.085000 ;
      RECT 1382.570000  2.085000 1382.840000 2.400000 ;
      RECT 1382.725000  0.900000 1382.895000 0.995000 ;
      RECT 1382.725000  0.995000 1383.905000 1.165000 ;
      RECT 1382.935000  1.165000 1383.905000 1.185000 ;
      RECT 1382.935000  1.185000 1383.190000 1.915000 ;
      RECT 1383.060000  2.255000 1383.390000 2.635000 ;
      RECT 1383.115000  0.085000 1383.495000 0.825000 ;
      RECT 1383.580000  1.355000 1384.115000 2.465000 ;
      RECT 1383.735000  0.255000 1384.895000 0.425000 ;
      RECT 1383.735000  0.425000 1383.905000 0.995000 ;
      RECT 1384.125000  0.675000 1384.505000 1.075000 ;
      RECT 1384.330000  1.075000 1384.505000 1.935000 ;
      RECT 1384.330000  1.935000 1386.110000 2.105000 ;
      RECT 1384.330000  2.105000 1384.500000 2.465000 ;
      RECT 1384.725000  0.425000 1384.895000 1.685000 ;
      RECT 1385.070000  0.710000 1385.415000 1.700000 ;
      RECT 1385.315000  2.275000 1385.665000 2.635000 ;
      RECT 1385.465000  0.085000 1385.810000 0.540000 ;
      RECT 1385.600000  0.715000 1386.180000 0.895000 ;
      RECT 1385.600000  0.895000 1385.770000 1.935000 ;
      RECT 1385.940000  1.065000 1386.110000 1.395000 ;
      RECT 1385.940000  2.105000 1386.110000 2.185000 ;
      RECT 1385.940000  2.185000 1386.310000 2.435000 ;
      RECT 1386.010000  0.335000 1386.350000 0.505000 ;
      RECT 1386.010000  0.505000 1386.180000 0.715000 ;
      RECT 1386.280000  1.575000 1386.580000 1.955000 ;
      RECT 1386.360000  0.705000 1387.110000 1.035000 ;
      RECT 1386.360000  1.035000 1386.580000 1.575000 ;
      RECT 1386.555000  2.135000 1386.920000 2.465000 ;
      RECT 1386.570000  0.305000 1387.470000 0.475000 ;
      RECT 1386.750000  1.215000 1388.610000 1.385000 ;
      RECT 1386.750000  1.385000 1386.920000 2.135000 ;
      RECT 1387.140000  1.935000 1388.400000 2.105000 ;
      RECT 1387.140000  2.105000 1387.310000 2.375000 ;
      RECT 1387.300000  0.475000 1387.470000 1.215000 ;
      RECT 1387.420000  1.595000 1389.000000 1.765000 ;
      RECT 1387.595000  2.355000 1387.925000 2.635000 ;
      RECT 1387.690000  0.765000 1388.270000 1.045000 ;
      RECT 1388.150000  0.085000 1388.480000 0.545000 ;
      RECT 1388.230000  2.105000 1388.400000 2.375000 ;
      RECT 1388.440000  1.005000 1388.610000 1.215000 ;
      RECT 1388.610000  2.175000 1389.030000 2.635000 ;
      RECT 1388.690000  0.275000 1389.070000 0.445000 ;
      RECT 1388.690000  0.445000 1389.000000 0.835000 ;
      RECT 1388.690000  1.765000 1389.000000 1.835000 ;
      RECT 1388.690000  1.835000 1389.445000 2.005000 ;
      RECT 1388.830000  0.835000 1389.000000 1.595000 ;
      RECT 1389.170000  0.705000 1389.430000 1.495000 ;
      RECT 1389.170000  1.495000 1389.905000 1.660000 ;
      RECT 1389.170000  1.660000 1390.305000 1.665000 ;
      RECT 1389.240000  0.255000 1390.350000 0.535000 ;
      RECT 1389.275000  2.005000 1389.445000 2.465000 ;
      RECT 1389.645000  1.665000 1390.305000 1.955000 ;
      RECT 1389.655000  2.125000 1390.675000 2.465000 ;
      RECT 1389.695000  0.920000 1389.865000 1.325000 ;
      RECT 1390.130000  0.535000 1390.350000 1.315000 ;
      RECT 1390.130000  1.315000 1390.745000 1.485000 ;
      RECT 1390.500000  1.485000 1390.745000 1.575000 ;
      RECT 1390.500000  1.575000 1391.830000 1.745000 ;
      RECT 1390.500000  1.745000 1390.675000 2.125000 ;
      RECT 1390.570000  0.085000 1390.790000 0.525000 ;
      RECT 1390.610000  0.695000 1391.190000 0.865000 ;
      RECT 1390.610000  0.865000 1390.830000 1.145000 ;
      RECT 1390.875000  2.195000 1391.125000 2.635000 ;
      RECT 1391.020000  0.295000 1392.190000 0.465000 ;
      RECT 1391.020000  0.465000 1391.190000 0.695000 ;
      RECT 1391.060000  1.065000 1391.830000 1.275000 ;
      RECT 1391.370000  1.915000 1392.190000 2.085000 ;
      RECT 1391.370000  2.085000 1391.540000 2.375000 ;
      RECT 1391.525000  0.635000 1391.830000 1.065000 ;
      RECT 1391.715000  2.255000 1392.095000 2.635000 ;
      RECT 1392.020000  0.465000 1392.190000 0.995000 ;
      RECT 1392.020000  0.995000 1392.665000 1.325000 ;
      RECT 1392.020000  1.325000 1392.190000 1.915000 ;
      RECT 1392.360000  0.345000 1392.530000 0.655000 ;
      RECT 1392.360000  0.655000 1393.100000 0.825000 ;
      RECT 1392.360000  1.795000 1393.100000 1.865000 ;
      RECT 1392.360000  1.865000 1394.060000 2.035000 ;
      RECT 1392.360000  2.035000 1392.535000 2.465000 ;
      RECT 1392.715000  2.205000 1393.175000 2.635000 ;
      RECT 1392.785000  0.085000 1393.115000 0.485000 ;
      RECT 1392.925000  0.825000 1393.100000 1.795000 ;
      RECT 1393.320000  0.265000 1393.720000 1.695000 ;
      RECT 1393.730000  2.255000 1394.185000 2.635000 ;
      RECT 1393.890000  0.995000 1394.325000 1.325000 ;
      RECT 1393.890000  1.325000 1394.060000 1.865000 ;
      RECT 1393.900000  0.085000 1394.070000 0.825000 ;
      RECT 1394.230000  1.535000 1394.665000 2.080000 ;
      RECT 1394.240000  0.310000 1394.665000 0.825000 ;
      RECT 1394.495000  0.825000 1394.665000 1.535000 ;
      RECT 1394.835000  0.085000 1395.005000 0.930000 ;
      RECT 1394.835000  1.495000 1395.085000 2.635000 ;
      RECT 1395.265000  0.085000 1395.555000 0.810000 ;
      RECT 1395.265000  1.470000 1395.555000 2.635000 ;
      RECT 1395.730000  1.795000 1396.555000 1.965000 ;
      RECT 1395.730000  1.965000 1395.985000 2.465000 ;
      RECT 1395.735000  0.345000 1395.985000 0.635000 ;
      RECT 1395.735000  0.635000 1396.525000 0.805000 ;
      RECT 1395.780000  0.975000 1396.130000 1.625000 ;
      RECT 1396.155000  0.085000 1396.535000 0.465000 ;
      RECT 1396.170000  2.135000 1396.550000 2.635000 ;
      RECT 1396.350000  0.805000 1396.525000 0.995000 ;
      RECT 1396.350000  0.995000 1396.665000 1.325000 ;
      RECT 1396.350000  1.325000 1396.555000 1.795000 ;
      RECT 1396.755000  0.345000 1397.005000 0.675000 ;
      RECT 1396.775000  1.730000 1397.005000 2.465000 ;
      RECT 1396.835000  0.675000 1397.005000 1.730000 ;
      RECT 1397.225000  1.070000 1397.630000 1.335000 ;
      RECT 1397.225000  1.335000 1397.860000 1.745000 ;
      RECT 1397.335000  0.395000 1397.505000 0.730000 ;
      RECT 1397.335000  0.730000 1398.075000 0.900000 ;
      RECT 1397.675000  0.085000 1398.055000 0.560000 ;
      RECT 1397.750000  1.915000 1398.370000 2.085000 ;
      RECT 1397.750000  2.085000 1398.020000 2.400000 ;
      RECT 1397.905000  0.900000 1398.075000 0.995000 ;
      RECT 1397.905000  0.995000 1399.085000 1.165000 ;
      RECT 1398.115000  1.165000 1399.085000 1.185000 ;
      RECT 1398.115000  1.185000 1398.370000 1.915000 ;
      RECT 1398.240000  2.255000 1398.570000 2.635000 ;
      RECT 1398.295000  0.085000 1398.675000 0.825000 ;
      RECT 1398.760000  1.355000 1399.295000 2.465000 ;
      RECT 1398.915000  0.255000 1400.075000 0.425000 ;
      RECT 1398.915000  0.425000 1399.085000 0.995000 ;
      RECT 1399.305000  0.675000 1399.685000 1.075000 ;
      RECT 1399.510000  1.075000 1399.685000 1.935000 ;
      RECT 1399.510000  1.935000 1401.290000 2.105000 ;
      RECT 1399.510000  2.105000 1399.680000 2.465000 ;
      RECT 1399.905000  0.425000 1400.075000 1.685000 ;
      RECT 1400.250000  0.710000 1400.595000 1.700000 ;
      RECT 1400.495000  2.275000 1400.845000 2.635000 ;
      RECT 1400.645000  0.085000 1400.990000 0.540000 ;
      RECT 1400.780000  0.715000 1401.360000 0.895000 ;
      RECT 1400.780000  0.895000 1400.950000 1.935000 ;
      RECT 1401.120000  1.065000 1401.290000 1.395000 ;
      RECT 1401.120000  2.105000 1401.290000 2.185000 ;
      RECT 1401.120000  2.185000 1401.490000 2.435000 ;
      RECT 1401.190000  0.335000 1401.530000 0.505000 ;
      RECT 1401.190000  0.505000 1401.360000 0.715000 ;
      RECT 1401.460000  1.575000 1401.760000 1.955000 ;
      RECT 1401.540000  0.705000 1402.290000 1.035000 ;
      RECT 1401.540000  1.035000 1401.760000 1.575000 ;
      RECT 1401.735000  2.135000 1402.100000 2.465000 ;
      RECT 1401.750000  0.305000 1402.650000 0.475000 ;
      RECT 1401.930000  1.215000 1403.790000 1.385000 ;
      RECT 1401.930000  1.385000 1402.100000 2.135000 ;
      RECT 1402.320000  1.935000 1403.580000 2.105000 ;
      RECT 1402.320000  2.105000 1402.490000 2.375000 ;
      RECT 1402.480000  0.475000 1402.650000 1.215000 ;
      RECT 1402.600000  1.595000 1404.180000 1.765000 ;
      RECT 1402.775000  2.355000 1403.105000 2.635000 ;
      RECT 1402.870000  0.765000 1403.450000 1.045000 ;
      RECT 1403.330000  0.085000 1403.660000 0.545000 ;
      RECT 1403.410000  2.105000 1403.580000 2.375000 ;
      RECT 1403.620000  1.005000 1403.790000 1.215000 ;
      RECT 1403.790000  2.175000 1404.210000 2.635000 ;
      RECT 1403.870000  0.275000 1404.250000 0.445000 ;
      RECT 1403.870000  0.445000 1404.180000 0.835000 ;
      RECT 1403.870000  1.765000 1404.180000 1.835000 ;
      RECT 1403.870000  1.835000 1404.625000 2.005000 ;
      RECT 1404.010000  0.835000 1404.180000 1.595000 ;
      RECT 1404.350000  0.705000 1404.610000 1.495000 ;
      RECT 1404.350000  1.495000 1405.085000 1.660000 ;
      RECT 1404.350000  1.660000 1405.485000 1.665000 ;
      RECT 1404.420000  0.255000 1405.530000 0.535000 ;
      RECT 1404.455000  2.005000 1404.625000 2.465000 ;
      RECT 1404.825000  1.665000 1405.485000 1.955000 ;
      RECT 1404.835000  2.125000 1405.855000 2.465000 ;
      RECT 1404.875000  0.920000 1405.045000 1.325000 ;
      RECT 1405.310000  0.535000 1405.530000 1.315000 ;
      RECT 1405.310000  1.315000 1405.925000 1.485000 ;
      RECT 1405.680000  1.485000 1405.925000 1.575000 ;
      RECT 1405.680000  1.575000 1407.010000 1.745000 ;
      RECT 1405.680000  1.745000 1405.855000 2.125000 ;
      RECT 1405.750000  0.085000 1405.970000 0.525000 ;
      RECT 1405.790000  0.695000 1406.370000 0.865000 ;
      RECT 1405.790000  0.865000 1406.010000 1.145000 ;
      RECT 1406.055000  2.195000 1406.305000 2.635000 ;
      RECT 1406.200000  0.295000 1407.375000 0.465000 ;
      RECT 1406.200000  0.465000 1406.370000 0.695000 ;
      RECT 1406.240000  1.065000 1407.010000 1.275000 ;
      RECT 1406.550000  1.915000 1407.370000 2.085000 ;
      RECT 1406.550000  2.085000 1406.720000 2.375000 ;
      RECT 1406.705000  0.635000 1407.010000 1.065000 ;
      RECT 1406.895000  2.255000 1407.275000 2.635000 ;
      RECT 1407.200000  0.465000 1407.375000 0.995000 ;
      RECT 1407.200000  0.995000 1407.845000 1.325000 ;
      RECT 1407.200000  1.325000 1407.370000 1.915000 ;
      RECT 1407.545000  0.085000 1407.830000 0.710000 ;
      RECT 1407.545000  1.495000 1407.830000 2.635000 ;
      RECT 1408.060000  0.265000 1408.425000 2.325000 ;
      RECT 1408.605000  0.085000 1408.895000 0.810000 ;
      RECT 1408.605000  1.470000 1408.895000 2.635000 ;
      RECT 1409.070000  1.795000 1409.895000 1.965000 ;
      RECT 1409.070000  1.965000 1409.325000 2.465000 ;
      RECT 1409.075000  0.345000 1409.325000 0.635000 ;
      RECT 1409.075000  0.635000 1409.865000 0.805000 ;
      RECT 1409.120000  0.975000 1409.470000 1.625000 ;
      RECT 1409.495000  0.085000 1409.875000 0.465000 ;
      RECT 1409.510000  2.135000 1409.890000 2.635000 ;
      RECT 1409.690000  0.805000 1409.865000 0.995000 ;
      RECT 1409.690000  0.995000 1410.005000 1.325000 ;
      RECT 1409.690000  1.325000 1409.895000 1.795000 ;
      RECT 1410.095000  0.345000 1410.345000 0.675000 ;
      RECT 1410.115000  1.730000 1410.345000 2.465000 ;
      RECT 1410.175000  0.675000 1410.345000 1.730000 ;
      RECT 1410.565000  1.070000 1410.970000 1.335000 ;
      RECT 1410.565000  1.335000 1411.200000 1.745000 ;
      RECT 1410.675000  0.395000 1410.845000 0.730000 ;
      RECT 1410.675000  0.730000 1411.415000 0.900000 ;
      RECT 1411.015000  0.085000 1411.395000 0.560000 ;
      RECT 1411.090000  1.915000 1411.710000 2.085000 ;
      RECT 1411.090000  2.085000 1411.360000 2.400000 ;
      RECT 1411.245000  0.900000 1411.415000 0.995000 ;
      RECT 1411.245000  0.995000 1412.425000 1.165000 ;
      RECT 1411.455000  1.165000 1412.425000 1.185000 ;
      RECT 1411.455000  1.185000 1411.710000 1.915000 ;
      RECT 1411.580000  2.255000 1411.910000 2.635000 ;
      RECT 1411.635000  0.085000 1412.015000 0.825000 ;
      RECT 1412.100000  1.355000 1412.635000 2.465000 ;
      RECT 1412.255000  0.255000 1413.415000 0.425000 ;
      RECT 1412.255000  0.425000 1412.425000 0.995000 ;
      RECT 1412.645000  0.675000 1413.025000 1.075000 ;
      RECT 1412.850000  1.075000 1413.025000 1.935000 ;
      RECT 1412.850000  1.935000 1414.630000 2.105000 ;
      RECT 1412.850000  2.105000 1413.020000 2.465000 ;
      RECT 1413.245000  0.425000 1413.415000 1.685000 ;
      RECT 1413.590000  0.710000 1413.935000 1.700000 ;
      RECT 1413.835000  2.275000 1414.185000 2.635000 ;
      RECT 1413.985000  0.085000 1414.330000 0.540000 ;
      RECT 1414.120000  0.715000 1414.700000 0.895000 ;
      RECT 1414.120000  0.895000 1414.290000 1.935000 ;
      RECT 1414.460000  1.065000 1414.630000 1.395000 ;
      RECT 1414.460000  2.105000 1414.630000 2.185000 ;
      RECT 1414.460000  2.185000 1414.830000 2.435000 ;
      RECT 1414.530000  0.335000 1414.870000 0.505000 ;
      RECT 1414.530000  0.505000 1414.700000 0.715000 ;
      RECT 1414.800000  1.575000 1415.100000 1.955000 ;
      RECT 1414.880000  0.705000 1415.630000 1.035000 ;
      RECT 1414.880000  1.035000 1415.100000 1.575000 ;
      RECT 1415.075000  2.135000 1415.440000 2.465000 ;
      RECT 1415.090000  0.305000 1415.990000 0.475000 ;
      RECT 1415.270000  1.215000 1417.130000 1.385000 ;
      RECT 1415.270000  1.385000 1415.440000 2.135000 ;
      RECT 1415.660000  1.935000 1416.920000 2.105000 ;
      RECT 1415.660000  2.105000 1415.830000 2.375000 ;
      RECT 1415.820000  0.475000 1415.990000 1.215000 ;
      RECT 1415.940000  1.595000 1417.520000 1.765000 ;
      RECT 1416.115000  2.355000 1416.445000 2.635000 ;
      RECT 1416.210000  0.765000 1416.790000 1.045000 ;
      RECT 1416.670000  0.085000 1417.000000 0.545000 ;
      RECT 1416.750000  2.105000 1416.920000 2.375000 ;
      RECT 1416.960000  1.005000 1417.130000 1.215000 ;
      RECT 1417.130000  2.175000 1417.550000 2.635000 ;
      RECT 1417.210000  0.275000 1417.590000 0.445000 ;
      RECT 1417.210000  0.445000 1417.520000 0.835000 ;
      RECT 1417.210000  1.765000 1417.520000 1.835000 ;
      RECT 1417.210000  1.835000 1417.965000 2.005000 ;
      RECT 1417.350000  0.835000 1417.520000 1.595000 ;
      RECT 1417.690000  0.705000 1417.950000 1.495000 ;
      RECT 1417.690000  1.495000 1418.425000 1.660000 ;
      RECT 1417.690000  1.660000 1418.825000 1.665000 ;
      RECT 1417.760000  0.255000 1418.870000 0.535000 ;
      RECT 1417.795000  2.005000 1417.965000 2.465000 ;
      RECT 1418.165000  1.665000 1418.825000 1.955000 ;
      RECT 1418.175000  2.125000 1419.195000 2.465000 ;
      RECT 1418.215000  0.920000 1418.385000 1.325000 ;
      RECT 1418.650000  0.535000 1418.870000 1.315000 ;
      RECT 1418.650000  1.315000 1419.265000 1.485000 ;
      RECT 1419.020000  1.485000 1419.265000 1.575000 ;
      RECT 1419.020000  1.575000 1420.350000 1.745000 ;
      RECT 1419.020000  1.745000 1419.195000 2.125000 ;
      RECT 1419.090000  0.085000 1419.310000 0.525000 ;
      RECT 1419.130000  0.695000 1419.710000 0.865000 ;
      RECT 1419.130000  0.865000 1419.350000 1.145000 ;
      RECT 1419.395000  2.195000 1419.645000 2.635000 ;
      RECT 1419.540000  0.295000 1420.715000 0.465000 ;
      RECT 1419.540000  0.465000 1419.710000 0.695000 ;
      RECT 1419.580000  1.065000 1420.350000 1.275000 ;
      RECT 1419.890000  1.915000 1420.710000 2.085000 ;
      RECT 1419.890000  2.085000 1420.060000 2.375000 ;
      RECT 1420.045000  0.635000 1420.350000 1.065000 ;
      RECT 1420.235000  2.255000 1420.615000 2.635000 ;
      RECT 1420.540000  0.465000 1420.715000 0.995000 ;
      RECT 1420.540000  0.995000 1421.185000 1.325000 ;
      RECT 1420.540000  1.325000 1420.710000 1.915000 ;
      RECT 1420.885000  0.085000 1421.170000 0.710000 ;
      RECT 1420.885000  1.495000 1421.170000 2.635000 ;
      RECT 1421.400000  0.265000 1421.765000 2.325000 ;
      RECT 1421.945000  0.085000 1422.235000 0.810000 ;
      RECT 1421.945000  1.470000 1422.235000 2.635000 ;
      RECT 1422.410000  1.795000 1423.235000 1.965000 ;
      RECT 1422.410000  1.965000 1422.665000 2.465000 ;
      RECT 1422.415000  0.345000 1422.665000 0.635000 ;
      RECT 1422.415000  0.635000 1423.205000 0.805000 ;
      RECT 1422.460000  0.975000 1422.810000 1.625000 ;
      RECT 1422.835000  0.085000 1423.215000 0.465000 ;
      RECT 1422.850000  2.135000 1423.230000 2.635000 ;
      RECT 1423.030000  0.805000 1423.205000 0.995000 ;
      RECT 1423.030000  0.995000 1423.345000 1.325000 ;
      RECT 1423.030000  1.325000 1423.235000 1.795000 ;
      RECT 1423.435000  0.345000 1423.685000 0.675000 ;
      RECT 1423.455000  1.730000 1423.685000 2.465000 ;
      RECT 1423.515000  0.675000 1423.685000 1.730000 ;
      RECT 1423.905000  1.070000 1424.310000 1.335000 ;
      RECT 1423.905000  1.335000 1424.540000 1.745000 ;
      RECT 1424.015000  0.395000 1424.185000 0.730000 ;
      RECT 1424.015000  0.730000 1424.755000 0.900000 ;
      RECT 1424.355000  0.085000 1424.735000 0.560000 ;
      RECT 1424.430000  1.915000 1425.050000 2.085000 ;
      RECT 1424.430000  2.085000 1424.700000 2.400000 ;
      RECT 1424.585000  0.900000 1424.755000 0.995000 ;
      RECT 1424.585000  0.995000 1425.765000 1.165000 ;
      RECT 1424.795000  1.165000 1425.765000 1.185000 ;
      RECT 1424.795000  1.185000 1425.050000 1.915000 ;
      RECT 1424.920000  2.255000 1425.250000 2.635000 ;
      RECT 1424.975000  0.085000 1425.355000 0.825000 ;
      RECT 1425.440000  1.355000 1425.975000 2.465000 ;
      RECT 1425.595000  0.255000 1426.755000 0.425000 ;
      RECT 1425.595000  0.425000 1425.765000 0.995000 ;
      RECT 1425.985000  0.675000 1426.365000 1.075000 ;
      RECT 1426.190000  1.075000 1426.365000 1.935000 ;
      RECT 1426.190000  1.935000 1427.970000 2.105000 ;
      RECT 1426.190000  2.105000 1426.360000 2.465000 ;
      RECT 1426.585000  0.425000 1426.755000 1.685000 ;
      RECT 1426.930000  0.710000 1427.275000 1.700000 ;
      RECT 1427.175000  2.275000 1427.525000 2.635000 ;
      RECT 1427.325000  0.085000 1427.670000 0.540000 ;
      RECT 1427.460000  0.715000 1428.040000 0.895000 ;
      RECT 1427.460000  0.895000 1427.630000 1.935000 ;
      RECT 1427.800000  1.065000 1427.970000 1.395000 ;
      RECT 1427.800000  2.105000 1427.970000 2.185000 ;
      RECT 1427.800000  2.185000 1428.170000 2.435000 ;
      RECT 1427.870000  0.335000 1428.210000 0.505000 ;
      RECT 1427.870000  0.505000 1428.040000 0.715000 ;
      RECT 1428.140000  1.575000 1428.440000 1.955000 ;
      RECT 1428.220000  0.705000 1428.970000 1.035000 ;
      RECT 1428.220000  1.035000 1428.440000 1.575000 ;
      RECT 1428.415000  2.135000 1428.780000 2.465000 ;
      RECT 1428.430000  0.305000 1429.330000 0.475000 ;
      RECT 1428.610000  1.215000 1430.470000 1.385000 ;
      RECT 1428.610000  1.385000 1428.780000 2.135000 ;
      RECT 1429.000000  1.935000 1430.260000 2.105000 ;
      RECT 1429.000000  2.105000 1429.170000 2.375000 ;
      RECT 1429.160000  0.475000 1429.330000 1.215000 ;
      RECT 1429.280000  1.595000 1430.860000 1.765000 ;
      RECT 1429.455000  2.355000 1429.785000 2.635000 ;
      RECT 1429.550000  0.765000 1430.130000 1.045000 ;
      RECT 1430.010000  0.085000 1430.340000 0.545000 ;
      RECT 1430.090000  2.105000 1430.260000 2.375000 ;
      RECT 1430.300000  1.005000 1430.470000 1.215000 ;
      RECT 1430.470000  2.175000 1430.890000 2.635000 ;
      RECT 1430.550000  0.275000 1430.930000 0.445000 ;
      RECT 1430.550000  0.445000 1430.860000 0.835000 ;
      RECT 1430.550000  1.765000 1430.860000 1.835000 ;
      RECT 1430.550000  1.835000 1431.305000 2.005000 ;
      RECT 1430.690000  0.835000 1430.860000 1.595000 ;
      RECT 1431.030000  0.705000 1431.290000 1.495000 ;
      RECT 1431.030000  1.495000 1431.765000 1.660000 ;
      RECT 1431.030000  1.660000 1432.165000 1.665000 ;
      RECT 1431.100000  0.255000 1432.210000 0.535000 ;
      RECT 1431.135000  2.005000 1431.305000 2.465000 ;
      RECT 1431.505000  1.665000 1432.165000 1.955000 ;
      RECT 1431.515000  2.125000 1432.535000 2.465000 ;
      RECT 1431.555000  0.920000 1431.725000 1.325000 ;
      RECT 1431.990000  0.535000 1432.210000 1.315000 ;
      RECT 1431.990000  1.315000 1432.605000 1.485000 ;
      RECT 1432.360000  1.485000 1432.605000 1.575000 ;
      RECT 1432.360000  1.575000 1433.690000 1.745000 ;
      RECT 1432.360000  1.745000 1432.535000 2.125000 ;
      RECT 1432.430000  0.085000 1432.650000 0.525000 ;
      RECT 1432.470000  0.695000 1433.050000 0.865000 ;
      RECT 1432.470000  0.865000 1432.690000 1.145000 ;
      RECT 1432.735000  2.195000 1432.985000 2.635000 ;
      RECT 1432.880000  0.295000 1434.055000 0.465000 ;
      RECT 1432.880000  0.465000 1433.050000 0.695000 ;
      RECT 1432.920000  1.065000 1433.690000 1.275000 ;
      RECT 1433.230000  1.915000 1434.050000 2.085000 ;
      RECT 1433.230000  2.085000 1433.400000 2.375000 ;
      RECT 1433.385000  0.635000 1433.690000 1.065000 ;
      RECT 1433.575000  2.255000 1433.955000 2.635000 ;
      RECT 1433.880000  0.465000 1434.055000 0.995000 ;
      RECT 1433.880000  0.995000 1434.555000 1.325000 ;
      RECT 1433.880000  1.325000 1434.050000 1.915000 ;
      RECT 1434.225000  0.085000 1434.645000 0.670000 ;
      RECT 1434.225000  1.495000 1434.650000 2.635000 ;
      RECT 1434.820000  0.265000 1435.105000 2.325000 ;
      RECT 1435.315000  0.085000 1435.485000 0.545000 ;
      RECT 1435.315000  1.495000 1435.565000 2.635000 ;
      RECT 1435.745000  0.085000 1436.035000 0.810000 ;
      RECT 1435.745000  1.470000 1436.035000 2.635000 ;
      RECT 1436.205000  0.085000 1436.550000 0.595000 ;
      RECT 1436.205000  0.765000 1436.485000 1.675000 ;
      RECT 1436.205000  1.845000 1437.325000 2.025000 ;
      RECT 1436.205000  2.025000 1436.465000 2.465000 ;
      RECT 1436.635000  2.195000 1436.935000 2.635000 ;
      RECT 1436.670000  0.765000 1436.980000 1.675000 ;
      RECT 1437.095000  0.280000 1437.965000 0.560000 ;
      RECT 1437.150000  0.765000 1437.545000 1.675000 ;
      RECT 1437.155000  2.025000 1437.325000 2.255000 ;
      RECT 1437.155000  2.255000 1438.365000 2.465000 ;
      RECT 1437.515000  1.870000 1437.965000 2.075000 ;
      RECT 1437.775000  0.560000 1437.965000 1.870000 ;
      RECT 1438.145000  0.085000 1438.325000 0.545000 ;
      RECT 1438.185000  0.715000 1438.835000 0.905000 ;
      RECT 1438.185000  0.905000 1438.520000 1.770000 ;
      RECT 1438.185000  1.770000 1438.805000 2.085000 ;
      RECT 1438.580000  0.255000 1438.835000 0.715000 ;
      RECT 1438.590000  2.085000 1438.805000 2.465000 ;
      RECT 1438.690000  1.075000 1439.070000 1.550000 ;
      RECT 1438.975000  1.720000 1439.455000 1.970000 ;
      RECT 1439.060000  0.085000 1439.400000 0.555000 ;
      RECT 1439.060000  2.140000 1439.400000 2.635000 ;
      RECT 1439.275000  1.055000 1439.935000 1.590000 ;
      RECT 1439.275000  1.590000 1439.455000 1.720000 ;
      RECT 1439.625000  1.775000 1440.415000 1.955000 ;
      RECT 1439.625000  1.955000 1439.795000 2.325000 ;
      RECT 1439.640000  0.255000 1439.825000 0.715000 ;
      RECT 1439.640000  0.715000 1440.415000 0.885000 ;
      RECT 1439.965000  2.275000 1440.345000 2.635000 ;
      RECT 1440.050000  0.085000 1440.360000 0.545000 ;
      RECT 1440.155000  0.885000 1440.415000 1.775000 ;
      RECT 1440.565000  2.135000 1440.910000 2.465000 ;
      RECT 1440.580000  0.255000 1440.805000 0.585000 ;
      RECT 1440.635000  0.585000 1440.805000 1.090000 ;
      RECT 1440.635000  1.090000 1440.960000 1.420000 ;
      RECT 1440.635000  1.420000 1440.910000 2.135000 ;
      RECT 1440.975000  0.255000 1441.300000 0.920000 ;
      RECT 1441.080000  1.590000 1441.300000 2.465000 ;
      RECT 1441.130000  0.920000 1441.300000 1.590000 ;
      RECT 1441.520000  0.255000 1442.010000 1.225000 ;
      RECT 1441.520000  1.225000 1444.480000 1.275000 ;
      RECT 1441.550000  2.135000 1442.325000 2.465000 ;
      RECT 1441.605000  1.275000 1443.055000 1.395000 ;
      RECT 1441.725000  1.575000 1441.985000 1.955000 ;
      RECT 1442.155000  1.395000 1442.325000 2.135000 ;
      RECT 1442.180000  0.085000 1442.715000 0.465000 ;
      RECT 1442.180000  0.635000 1443.205000 0.805000 ;
      RECT 1442.180000  0.805000 1442.595000 1.015000 ;
      RECT 1442.545000  1.575000 1442.715000 1.935000 ;
      RECT 1442.545000  1.935000 1443.485000 2.105000 ;
      RECT 1442.565000  2.275000 1442.895000 2.635000 ;
      RECT 1442.870000  0.975000 1444.480000 1.225000 ;
      RECT 1442.895000  0.255000 1443.205000 0.635000 ;
      RECT 1443.220000  2.105000 1443.485000 2.450000 ;
      RECT 1443.310000  1.445000 1443.845000 1.765000 ;
      RECT 1443.660000  0.085000 1444.395000 0.690000 ;
      RECT 1443.775000  2.125000 1444.830000 2.635000 ;
      RECT 1444.030000  1.495000 1444.875000 1.955000 ;
      RECT 1444.070000  1.275000 1444.480000 1.325000 ;
      RECT 1444.655000  0.695000 1446.010000 0.895000 ;
      RECT 1444.655000  0.895000 1444.875000 1.495000 ;
      RECT 1445.000000  2.125000 1445.855000 2.460000 ;
      RECT 1445.235000  1.075000 1445.515000 1.905000 ;
      RECT 1445.280000  0.275000 1446.895000 0.445000 ;
      RECT 1445.685000  1.895000 1447.585000 2.065000 ;
      RECT 1445.685000  2.065000 1445.855000 2.125000 ;
      RECT 1445.730000  0.895000 1446.010000 1.245000 ;
      RECT 1445.805000  1.415000 1446.080000 1.525000 ;
      RECT 1445.805000  1.525000 1447.195000 1.725000 ;
      RECT 1446.165000  2.235000 1446.545000 2.635000 ;
      RECT 1446.260000  0.855000 1446.485000 1.185000 ;
      RECT 1446.260000  1.185000 1448.065000 1.355000 ;
      RECT 1446.725000  0.445000 1446.895000 0.845000 ;
      RECT 1446.725000  0.845000 1447.665000 1.015000 ;
      RECT 1446.765000  2.065000 1446.980000 2.450000 ;
      RECT 1447.255000  2.235000 1447.585000 2.635000 ;
      RECT 1447.340000  0.085000 1447.510000 0.545000 ;
      RECT 1447.365000  1.525000 1447.585000 1.895000 ;
      RECT 1447.680000  0.255000 1448.065000 0.540000 ;
      RECT 1447.805000  1.355000 1448.065000 2.465000 ;
      RECT 1447.885000  0.540000 1448.065000 1.185000 ;
      RECT 1448.290000  0.085000 1448.500000 0.885000 ;
      RECT 1448.290000  1.485000 1448.500000 2.635000 ;
      RECT 1448.670000  0.255000 1449.050000 2.465000 ;
      RECT 1449.280000  0.255000 1449.490000 0.995000 ;
      RECT 1449.280000  0.995000 1450.170000 1.325000 ;
      RECT 1449.280000  1.325000 1449.490000 2.465000 ;
      RECT 1449.810000  0.085000 1450.015000 0.825000 ;
      RECT 1449.845000  1.575000 1450.015000 2.635000 ;
      RECT 1450.185000  0.275000 1450.745000 0.825000 ;
      RECT 1450.185000  1.495000 1450.745000 2.450000 ;
      RECT 1450.390000  0.825000 1450.745000 1.495000 ;
      RECT 1450.925000  0.085000 1451.215000 0.810000 ;
      RECT 1450.925000  1.470000 1451.215000 2.635000 ;
      RECT 1451.385000  0.085000 1451.730000 0.595000 ;
      RECT 1451.385000  0.765000 1451.665000 1.675000 ;
      RECT 1451.385000  1.845000 1452.505000 2.025000 ;
      RECT 1451.385000  2.025000 1451.645000 2.465000 ;
      RECT 1451.815000  2.195000 1452.115000 2.635000 ;
      RECT 1451.850000  0.765000 1452.160000 1.675000 ;
      RECT 1452.275000  0.280000 1453.145000 0.560000 ;
      RECT 1452.330000  0.765000 1452.725000 1.675000 ;
      RECT 1452.335000  2.025000 1452.505000 2.255000 ;
      RECT 1452.335000  2.255000 1453.545000 2.465000 ;
      RECT 1452.695000  1.870000 1453.145000 2.075000 ;
      RECT 1452.955000  0.560000 1453.145000 1.870000 ;
      RECT 1453.325000  0.085000 1453.505000 0.545000 ;
      RECT 1453.365000  0.715000 1454.015000 0.905000 ;
      RECT 1453.365000  0.905000 1453.700000 1.770000 ;
      RECT 1453.365000  1.770000 1453.985000 2.085000 ;
      RECT 1453.760000  0.255000 1454.015000 0.715000 ;
      RECT 1453.770000  2.085000 1453.985000 2.465000 ;
      RECT 1453.870000  1.075000 1454.250000 1.550000 ;
      RECT 1454.155000  1.720000 1454.635000 1.970000 ;
      RECT 1454.240000  0.085000 1454.580000 0.555000 ;
      RECT 1454.240000  2.140000 1454.580000 2.635000 ;
      RECT 1454.455000  1.055000 1455.115000 1.590000 ;
      RECT 1454.455000  1.590000 1454.635000 1.720000 ;
      RECT 1454.805000  1.775000 1455.595000 1.955000 ;
      RECT 1454.805000  1.955000 1454.975000 2.325000 ;
      RECT 1454.820000  0.255000 1455.005000 0.715000 ;
      RECT 1454.820000  0.715000 1455.595000 0.885000 ;
      RECT 1455.145000  2.275000 1455.525000 2.635000 ;
      RECT 1455.230000  0.085000 1455.540000 0.545000 ;
      RECT 1455.335000  0.885000 1455.595000 1.775000 ;
      RECT 1455.745000  2.135000 1456.090000 2.465000 ;
      RECT 1455.760000  0.255000 1455.985000 0.585000 ;
      RECT 1455.815000  0.585000 1455.985000 1.090000 ;
      RECT 1455.815000  1.090000 1456.140000 1.420000 ;
      RECT 1455.815000  1.420000 1456.090000 2.135000 ;
      RECT 1456.155000  0.255000 1456.480000 0.920000 ;
      RECT 1456.260000  1.590000 1456.480000 2.465000 ;
      RECT 1456.310000  0.920000 1456.480000 1.590000 ;
      RECT 1456.700000  0.255000 1457.190000 1.225000 ;
      RECT 1456.700000  1.225000 1459.660000 1.275000 ;
      RECT 1456.730000  2.135000 1457.505000 2.465000 ;
      RECT 1456.785000  1.275000 1458.235000 1.395000 ;
      RECT 1456.905000  1.575000 1457.165000 1.955000 ;
      RECT 1457.335000  1.395000 1457.505000 2.135000 ;
      RECT 1457.360000  0.085000 1457.895000 0.465000 ;
      RECT 1457.360000  0.635000 1458.385000 0.805000 ;
      RECT 1457.360000  0.805000 1457.775000 1.015000 ;
      RECT 1457.725000  1.575000 1457.895000 1.935000 ;
      RECT 1457.725000  1.935000 1458.665000 2.105000 ;
      RECT 1457.745000  2.275000 1458.075000 2.635000 ;
      RECT 1458.050000  0.975000 1459.660000 1.225000 ;
      RECT 1458.075000  0.255000 1458.385000 0.635000 ;
      RECT 1458.400000  2.105000 1458.665000 2.450000 ;
      RECT 1458.490000  1.445000 1459.025000 1.765000 ;
      RECT 1458.840000  0.085000 1459.575000 0.690000 ;
      RECT 1458.955000  2.125000 1460.010000 2.635000 ;
      RECT 1459.210000  1.495000 1460.055000 1.955000 ;
      RECT 1459.250000  1.275000 1459.660000 1.325000 ;
      RECT 1459.835000  0.695000 1461.190000 0.895000 ;
      RECT 1459.835000  0.895000 1460.055000 1.495000 ;
      RECT 1460.180000  2.125000 1461.035000 2.460000 ;
      RECT 1460.415000  1.075000 1460.695000 1.905000 ;
      RECT 1460.460000  0.275000 1462.075000 0.445000 ;
      RECT 1460.865000  1.895000 1462.765000 2.065000 ;
      RECT 1460.865000  2.065000 1461.035000 2.125000 ;
      RECT 1460.910000  0.895000 1461.190000 1.245000 ;
      RECT 1460.985000  1.415000 1461.260000 1.525000 ;
      RECT 1460.985000  1.525000 1462.375000 1.725000 ;
      RECT 1461.345000  2.235000 1461.725000 2.635000 ;
      RECT 1461.440000  0.855000 1461.665000 1.185000 ;
      RECT 1461.440000  1.185000 1463.245000 1.355000 ;
      RECT 1461.905000  0.445000 1462.075000 0.845000 ;
      RECT 1461.905000  0.845000 1462.845000 1.015000 ;
      RECT 1461.945000  2.065000 1462.160000 2.450000 ;
      RECT 1462.435000  2.235000 1462.765000 2.635000 ;
      RECT 1462.520000  0.085000 1462.690000 0.545000 ;
      RECT 1462.545000  1.525000 1462.765000 1.895000 ;
      RECT 1462.860000  0.255000 1463.245000 0.540000 ;
      RECT 1462.985000  1.355000 1463.245000 2.465000 ;
      RECT 1463.065000  0.540000 1463.245000 1.185000 ;
      RECT 1463.470000  0.085000 1463.680000 0.885000 ;
      RECT 1463.470000  1.485000 1463.680000 2.635000 ;
      RECT 1463.855000  0.255000 1464.300000 2.465000 ;
      RECT 1464.515000  0.085000 1464.805000 0.885000 ;
      RECT 1464.515000  1.485000 1464.805000 2.635000 ;
      RECT 1465.020000  0.255000 1465.205000 0.995000 ;
      RECT 1465.020000  0.995000 1465.885000 1.325000 ;
      RECT 1465.020000  1.325000 1465.205000 2.465000 ;
      RECT 1465.375000  0.085000 1465.780000 0.825000 ;
      RECT 1465.375000  1.635000 1465.780000 2.635000 ;
      RECT 1466.000000  0.275000 1466.380000 0.825000 ;
      RECT 1466.000000  1.495000 1466.380000 2.450000 ;
      RECT 1466.105000  0.825000 1466.380000 1.495000 ;
      RECT 1466.550000  0.085000 1466.815000 0.885000 ;
      RECT 1466.550000  1.485000 1466.815000 2.635000 ;
      RECT 1467.025000  0.085000 1467.315000 0.810000 ;
      RECT 1467.025000  1.470000 1467.315000 2.635000 ;
      RECT 1467.485000  0.085000 1468.150000 0.595000 ;
      RECT 1467.485000  0.765000 1467.740000 1.675000 ;
      RECT 1467.485000  1.845000 1468.625000 2.025000 ;
      RECT 1467.485000  2.025000 1467.745000 2.465000 ;
      RECT 1467.915000  2.195000 1468.235000 2.635000 ;
      RECT 1467.940000  0.765000 1468.270000 1.675000 ;
      RECT 1468.320000  0.255000 1469.245000 0.595000 ;
      RECT 1468.440000  0.765000 1468.885000 1.675000 ;
      RECT 1468.455000  2.025000 1468.625000 2.255000 ;
      RECT 1468.455000  2.255000 1469.645000 2.465000 ;
      RECT 1468.795000  1.845000 1469.245000 2.085000 ;
      RECT 1469.055000  0.595000 1469.245000 1.845000 ;
      RECT 1469.425000  0.085000 1469.690000 0.545000 ;
      RECT 1469.465000  0.715000 1470.120000 0.905000 ;
      RECT 1469.465000  0.905000 1469.800000 1.770000 ;
      RECT 1469.465000  1.770000 1470.120000 2.085000 ;
      RECT 1469.860000  0.255000 1470.120000 0.715000 ;
      RECT 1469.870000  2.085000 1470.120000 2.465000 ;
      RECT 1469.970000  1.075000 1470.350000 1.600000 ;
      RECT 1470.340000  0.085000 1470.750000 0.555000 ;
      RECT 1470.340000  2.140000 1470.635000 2.635000 ;
      RECT 1470.555000  1.055000 1471.215000 1.650000 ;
      RECT 1470.905000  1.830000 1471.695000 2.000000 ;
      RECT 1470.905000  2.000000 1471.075000 2.325000 ;
      RECT 1470.920000  0.255000 1471.105000 0.715000 ;
      RECT 1470.920000  0.715000 1471.695000 0.885000 ;
      RECT 1471.245000  2.275000 1471.625000 2.635000 ;
      RECT 1471.325000  0.085000 1471.655000 0.545000 ;
      RECT 1471.435000  0.885000 1471.695000 1.830000 ;
      RECT 1471.845000  2.135000 1472.190000 2.465000 ;
      RECT 1471.875000  0.255000 1472.085000 1.085000 ;
      RECT 1471.875000  1.085000 1472.240000 1.420000 ;
      RECT 1471.875000  1.420000 1472.190000 2.135000 ;
      RECT 1472.255000  0.255000 1472.580000 0.780000 ;
      RECT 1472.365000  1.590000 1472.580000 2.465000 ;
      RECT 1472.410000  0.780000 1472.580000 1.590000 ;
      RECT 1472.835000  2.135000 1473.605000 2.465000 ;
      RECT 1472.865000  0.255000 1473.290000 1.225000 ;
      RECT 1472.865000  1.225000 1475.715000 1.275000 ;
      RECT 1472.865000  1.275000 1474.375000 1.395000 ;
      RECT 1473.005000  1.575000 1473.265000 1.955000 ;
      RECT 1473.435000  1.395000 1473.605000 2.135000 ;
      RECT 1473.460000  0.085000 1473.995000 0.465000 ;
      RECT 1473.495000  0.635000 1474.435000 0.805000 ;
      RECT 1473.495000  0.805000 1473.875000 1.015000 ;
      RECT 1473.825000  1.575000 1473.995000 1.935000 ;
      RECT 1473.825000  1.935000 1474.820000 2.105000 ;
      RECT 1473.845000  2.275000 1474.230000 2.635000 ;
      RECT 1474.185000  0.255000 1474.435000 0.635000 ;
      RECT 1474.205000  0.975000 1475.715000 1.225000 ;
      RECT 1474.555000  2.105000 1474.820000 2.450000 ;
      RECT 1474.590000  1.445000 1475.115000 1.765000 ;
      RECT 1474.655000  0.085000 1475.715000 0.805000 ;
      RECT 1475.110000  2.125000 1476.025000 2.635000 ;
      RECT 1475.285000  1.670000 1476.185000 1.955000 ;
      RECT 1475.305000  1.275000 1475.715000 1.325000 ;
      RECT 1475.885000  0.720000 1477.250000 0.905000 ;
      RECT 1475.885000  0.905000 1476.185000 1.670000 ;
      RECT 1476.195000  2.125000 1477.090000 2.460000 ;
      RECT 1476.355000  1.075000 1476.690000 1.905000 ;
      RECT 1476.425000  0.275000 1478.050000 0.545000 ;
      RECT 1476.920000  0.905000 1477.250000 1.255000 ;
      RECT 1476.920000  1.895000 1478.655000 2.065000 ;
      RECT 1476.920000  2.065000 1477.090000 2.125000 ;
      RECT 1476.980000  1.425000 1477.260000 1.545000 ;
      RECT 1476.980000  1.545000 1478.095000 1.725000 ;
      RECT 1477.260000  2.235000 1477.590000 2.635000 ;
      RECT 1477.435000  0.855000 1477.680000 1.195000 ;
      RECT 1477.435000  1.195000 1479.085000 1.365000 ;
      RECT 1477.795000  2.065000 1477.995000 2.450000 ;
      RECT 1477.850000  0.545000 1478.050000 0.785000 ;
      RECT 1477.850000  0.785000 1478.685000 1.015000 ;
      RECT 1478.235000  0.085000 1478.485000 0.545000 ;
      RECT 1478.275000  1.605000 1478.655000 1.895000 ;
      RECT 1478.275000  2.235000 1478.655000 2.635000 ;
      RECT 1478.745000  0.255000 1479.085000 0.585000 ;
      RECT 1478.825000  1.365000 1479.085000 2.465000 ;
      RECT 1478.855000  0.585000 1479.085000 1.195000 ;
      RECT 1479.255000  0.255000 1479.515000 0.995000 ;
      RECT 1479.255000  0.995000 1480.145000 1.325000 ;
      RECT 1479.255000  1.325000 1479.595000 2.465000 ;
      RECT 1479.685000  0.085000 1480.090000 0.550000 ;
      RECT 1479.835000  1.845000 1480.090000 2.635000 ;
      RECT 1480.315000  0.275000 1480.640000 2.450000 ;
      RECT 1480.825000  0.085000 1481.115000 0.810000 ;
      RECT 1480.825000  1.470000 1481.115000 2.635000 ;
      RECT 1481.285000  0.085000 1481.950000 0.595000 ;
      RECT 1481.285000  0.765000 1481.540000 1.675000 ;
      RECT 1481.285000  1.845000 1482.425000 2.025000 ;
      RECT 1481.285000  2.025000 1481.545000 2.465000 ;
      RECT 1481.715000  2.195000 1482.035000 2.635000 ;
      RECT 1481.740000  0.765000 1482.070000 1.675000 ;
      RECT 1482.120000  0.255000 1483.045000 0.595000 ;
      RECT 1482.240000  0.765000 1482.685000 1.675000 ;
      RECT 1482.255000  2.025000 1482.425000 2.255000 ;
      RECT 1482.255000  2.255000 1483.445000 2.465000 ;
      RECT 1482.595000  1.845000 1483.045000 2.085000 ;
      RECT 1482.855000  0.595000 1483.045000 1.845000 ;
      RECT 1483.225000  0.085000 1483.490000 0.545000 ;
      RECT 1483.265000  0.715000 1483.920000 0.905000 ;
      RECT 1483.265000  0.905000 1483.600000 1.770000 ;
      RECT 1483.265000  1.770000 1483.920000 2.085000 ;
      RECT 1483.660000  0.255000 1483.920000 0.715000 ;
      RECT 1483.670000  2.085000 1483.920000 2.465000 ;
      RECT 1483.770000  1.075000 1484.150000 1.600000 ;
      RECT 1484.140000  0.085000 1484.550000 0.555000 ;
      RECT 1484.140000  2.140000 1484.435000 2.635000 ;
      RECT 1484.355000  1.055000 1485.015000 1.650000 ;
      RECT 1484.705000  1.830000 1485.495000 2.000000 ;
      RECT 1484.705000  2.000000 1484.875000 2.325000 ;
      RECT 1484.720000  0.255000 1484.905000 0.715000 ;
      RECT 1484.720000  0.715000 1485.495000 0.885000 ;
      RECT 1485.045000  2.275000 1485.425000 2.635000 ;
      RECT 1485.125000  0.085000 1485.455000 0.545000 ;
      RECT 1485.235000  0.885000 1485.495000 1.830000 ;
      RECT 1485.645000  2.135000 1485.990000 2.465000 ;
      RECT 1485.675000  0.255000 1485.885000 1.085000 ;
      RECT 1485.675000  1.085000 1486.040000 1.420000 ;
      RECT 1485.675000  1.420000 1485.990000 2.135000 ;
      RECT 1486.055000  0.255000 1486.380000 0.780000 ;
      RECT 1486.165000  1.590000 1486.380000 2.465000 ;
      RECT 1486.210000  0.780000 1486.380000 1.590000 ;
      RECT 1486.635000  2.135000 1487.405000 2.465000 ;
      RECT 1486.665000  0.255000 1487.090000 1.225000 ;
      RECT 1486.665000  1.225000 1489.615000 1.275000 ;
      RECT 1486.665000  1.275000 1488.175000 1.395000 ;
      RECT 1486.805000  1.575000 1487.065000 1.955000 ;
      RECT 1487.235000  1.395000 1487.405000 2.135000 ;
      RECT 1487.260000  0.085000 1487.795000 0.465000 ;
      RECT 1487.295000  0.635000 1488.235000 0.805000 ;
      RECT 1487.295000  0.805000 1487.675000 1.015000 ;
      RECT 1487.625000  1.575000 1487.795000 1.935000 ;
      RECT 1487.625000  1.935000 1488.620000 2.105000 ;
      RECT 1487.645000  2.275000 1488.030000 2.635000 ;
      RECT 1487.985000  0.255000 1488.235000 0.635000 ;
      RECT 1488.005000  0.975000 1489.615000 1.225000 ;
      RECT 1488.355000  2.105000 1488.620000 2.450000 ;
      RECT 1488.390000  1.445000 1488.915000 1.765000 ;
      RECT 1488.455000  0.085000 1489.615000 0.805000 ;
      RECT 1488.910000  2.125000 1489.965000 2.635000 ;
      RECT 1489.085000  1.670000 1490.085000 1.955000 ;
      RECT 1489.205000  1.275000 1489.615000 1.325000 ;
      RECT 1489.785000  0.720000 1491.205000 0.905000 ;
      RECT 1489.785000  0.905000 1490.085000 1.670000 ;
      RECT 1490.135000  2.125000 1491.040000 2.460000 ;
      RECT 1490.375000  1.075000 1490.700000 1.905000 ;
      RECT 1490.465000  0.275000 1492.110000 0.545000 ;
      RECT 1490.870000  0.905000 1491.205000 1.255000 ;
      RECT 1490.870000  1.895000 1492.785000 2.065000 ;
      RECT 1490.870000  2.065000 1491.040000 2.125000 ;
      RECT 1490.930000  1.425000 1491.235000 1.545000 ;
      RECT 1490.930000  1.545000 1492.195000 1.725000 ;
      RECT 1491.260000  2.235000 1491.640000 2.635000 ;
      RECT 1491.420000  0.855000 1491.680000 1.195000 ;
      RECT 1491.420000  1.195000 1493.215000 1.365000 ;
      RECT 1491.810000  2.065000 1492.215000 2.450000 ;
      RECT 1491.910000  0.545000 1492.110000 0.785000 ;
      RECT 1491.910000  0.785000 1492.815000 1.015000 ;
      RECT 1492.365000  0.085000 1492.615000 0.545000 ;
      RECT 1492.405000  1.605000 1492.785000 1.895000 ;
      RECT 1492.405000  2.235000 1492.785000 2.635000 ;
      RECT 1492.875000  0.255000 1493.215000 0.585000 ;
      RECT 1492.955000  1.365000 1493.215000 2.465000 ;
      RECT 1492.985000  0.585000 1493.215000 1.195000 ;
      RECT 1493.385000  0.255000 1493.645000 0.995000 ;
      RECT 1493.385000  0.995000 1494.325000 1.325000 ;
      RECT 1493.385000  1.325000 1493.725000 2.465000 ;
      RECT 1493.815000  0.085000 1494.220000 0.550000 ;
      RECT 1493.965000  1.845000 1494.220000 2.635000 ;
      RECT 1494.445000  0.275000 1494.855000 0.825000 ;
      RECT 1494.445000  1.495000 1494.855000 2.450000 ;
      RECT 1494.550000  0.825000 1494.855000 1.495000 ;
      RECT 1495.025000  0.085000 1495.195000 0.885000 ;
      RECT 1495.025000  1.495000 1495.195000 2.635000 ;
      RECT 1495.545000  0.085000 1495.835000 0.810000 ;
      RECT 1495.545000  1.470000 1495.835000 2.635000 ;
      RECT 1496.005000  0.085000 1496.670000 0.595000 ;
      RECT 1496.005000  0.765000 1496.260000 1.675000 ;
      RECT 1496.005000  1.845000 1497.145000 2.025000 ;
      RECT 1496.005000  2.025000 1496.265000 2.465000 ;
      RECT 1496.435000  2.195000 1496.755000 2.635000 ;
      RECT 1496.460000  0.765000 1496.790000 1.675000 ;
      RECT 1496.840000  0.255000 1497.765000 0.595000 ;
      RECT 1496.960000  0.765000 1497.405000 1.675000 ;
      RECT 1496.975000  2.025000 1497.145000 2.255000 ;
      RECT 1496.975000  2.255000 1498.165000 2.465000 ;
      RECT 1497.315000  1.845000 1497.765000 2.085000 ;
      RECT 1497.575000  0.595000 1497.765000 1.845000 ;
      RECT 1497.945000  0.085000 1498.210000 0.545000 ;
      RECT 1497.985000  0.715000 1498.640000 0.905000 ;
      RECT 1497.985000  0.905000 1498.320000 1.770000 ;
      RECT 1497.985000  1.770000 1498.640000 2.085000 ;
      RECT 1498.380000  0.255000 1498.640000 0.715000 ;
      RECT 1498.390000  2.085000 1498.640000 2.465000 ;
      RECT 1498.490000  1.075000 1498.870000 1.600000 ;
      RECT 1498.860000  0.085000 1499.270000 0.555000 ;
      RECT 1498.860000  2.140000 1499.155000 2.635000 ;
      RECT 1499.075000  1.055000 1499.735000 1.650000 ;
      RECT 1499.425000  1.830000 1500.215000 2.000000 ;
      RECT 1499.425000  2.000000 1499.595000 2.325000 ;
      RECT 1499.440000  0.255000 1499.625000 0.715000 ;
      RECT 1499.440000  0.715000 1500.215000 0.885000 ;
      RECT 1499.765000  2.275000 1500.145000 2.635000 ;
      RECT 1499.845000  0.085000 1500.175000 0.545000 ;
      RECT 1499.955000  0.885000 1500.215000 1.830000 ;
      RECT 1500.365000  2.135000 1500.710000 2.465000 ;
      RECT 1500.395000  0.255000 1500.605000 1.085000 ;
      RECT 1500.395000  1.085000 1500.760000 1.420000 ;
      RECT 1500.395000  1.420000 1500.710000 2.135000 ;
      RECT 1500.775000  0.255000 1501.100000 0.780000 ;
      RECT 1500.885000  1.590000 1501.100000 2.465000 ;
      RECT 1500.930000  0.780000 1501.100000 1.590000 ;
      RECT 1501.355000  2.135000 1502.125000 2.465000 ;
      RECT 1501.385000  0.255000 1501.810000 1.225000 ;
      RECT 1501.385000  1.225000 1504.335000 1.275000 ;
      RECT 1501.385000  1.275000 1502.895000 1.395000 ;
      RECT 1501.525000  1.575000 1501.785000 1.955000 ;
      RECT 1501.955000  1.395000 1502.125000 2.135000 ;
      RECT 1501.980000  0.085000 1502.515000 0.465000 ;
      RECT 1502.015000  0.635000 1502.955000 0.805000 ;
      RECT 1502.015000  0.805000 1502.395000 1.015000 ;
      RECT 1502.345000  1.575000 1502.515000 1.935000 ;
      RECT 1502.345000  1.935000 1503.340000 2.105000 ;
      RECT 1502.365000  2.275000 1502.750000 2.635000 ;
      RECT 1502.705000  0.255000 1502.955000 0.635000 ;
      RECT 1502.725000  0.975000 1504.335000 1.225000 ;
      RECT 1503.075000  2.105000 1503.340000 2.450000 ;
      RECT 1503.110000  1.445000 1503.635000 1.765000 ;
      RECT 1503.175000  0.085000 1504.335000 0.805000 ;
      RECT 1503.630000  2.125000 1504.685000 2.635000 ;
      RECT 1503.805000  1.670000 1504.805000 1.955000 ;
      RECT 1503.925000  1.275000 1504.335000 1.325000 ;
      RECT 1504.505000  0.720000 1505.925000 0.905000 ;
      RECT 1504.505000  0.905000 1504.805000 1.670000 ;
      RECT 1504.855000  2.125000 1505.760000 2.460000 ;
      RECT 1505.095000  1.075000 1505.420000 1.905000 ;
      RECT 1505.185000  0.275000 1506.830000 0.545000 ;
      RECT 1505.590000  0.905000 1505.925000 1.255000 ;
      RECT 1505.590000  1.895000 1507.505000 2.065000 ;
      RECT 1505.590000  2.065000 1505.760000 2.125000 ;
      RECT 1505.650000  1.425000 1505.955000 1.545000 ;
      RECT 1505.650000  1.545000 1506.915000 1.725000 ;
      RECT 1505.980000  2.235000 1506.360000 2.635000 ;
      RECT 1506.140000  0.855000 1506.400000 1.195000 ;
      RECT 1506.140000  1.195000 1507.935000 1.365000 ;
      RECT 1506.530000  2.065000 1506.935000 2.450000 ;
      RECT 1506.630000  0.545000 1506.830000 0.785000 ;
      RECT 1506.630000  0.785000 1507.535000 1.015000 ;
      RECT 1507.085000  0.085000 1507.335000 0.545000 ;
      RECT 1507.125000  1.605000 1507.505000 1.895000 ;
      RECT 1507.125000  2.235000 1507.505000 2.635000 ;
      RECT 1507.595000  0.255000 1507.935000 0.585000 ;
      RECT 1507.675000  1.365000 1507.935000 2.465000 ;
      RECT 1507.705000  0.585000 1507.935000 1.195000 ;
      RECT 1508.105000  0.255000 1508.365000 0.995000 ;
      RECT 1508.105000  0.995000 1509.045000 1.325000 ;
      RECT 1508.105000  1.325000 1508.365000 2.465000 ;
      RECT 1508.535000  0.085000 1508.940000 0.825000 ;
      RECT 1508.535000  1.495000 1508.940000 2.635000 ;
      RECT 1509.160000  0.275000 1509.490000 0.825000 ;
      RECT 1509.160000  1.495000 1509.490000 2.450000 ;
      RECT 1509.265000  0.825000 1509.490000 1.055000 ;
      RECT 1509.265000  1.055000 1510.530000 1.325000 ;
      RECT 1509.265000  1.325000 1509.490000 1.495000 ;
      RECT 1509.710000  0.085000 1509.880000 0.885000 ;
      RECT 1509.710000  1.495000 1509.880000 2.635000 ;
      RECT 1510.050000  0.255000 1510.530000 1.055000 ;
      RECT 1510.050000  1.325000 1510.530000 2.465000 ;
      RECT 1510.700000  0.085000 1510.985000 0.885000 ;
      RECT 1510.700000  1.495000 1510.985000 2.635000 ;
      RECT 1511.185000  0.085000 1511.475000 0.810000 ;
      RECT 1511.185000  1.470000 1511.475000 2.635000 ;
      RECT 1511.655000  0.975000 1512.005000 1.625000 ;
      RECT 1511.735000  0.345000 1511.905000 0.635000 ;
      RECT 1511.735000  0.635000 1512.420000 0.805000 ;
      RECT 1511.735000  1.795000 1512.455000 1.965000 ;
      RECT 1511.735000  1.965000 1511.905000 2.465000 ;
      RECT 1512.075000  0.085000 1512.455000 0.465000 ;
      RECT 1512.075000  2.135000 1512.455000 2.635000 ;
      RECT 1512.225000  0.805000 1512.420000 0.970000 ;
      RECT 1512.225000  0.970000 1512.455000 1.795000 ;
      RECT 1512.675000  0.345000 1512.845000 2.465000 ;
      RECT 1513.080000  0.255000 1513.465000 0.445000 ;
      RECT 1513.080000  0.445000 1513.250000 1.860000 ;
      RECT 1513.080000  1.860000 1515.090000 2.075000 ;
      RECT 1513.080000  2.075000 1513.365000 2.445000 ;
      RECT 1513.420000  0.615000 1515.095000 0.785000 ;
      RECT 1513.420000  0.785000 1513.590000 1.685000 ;
      RECT 1513.535000  2.245000 1513.915000 2.635000 ;
      RECT 1513.705000  0.085000 1514.035000 0.445000 ;
      RECT 1513.810000  0.955000 1514.255000 1.125000 ;
      RECT 1513.810000  1.125000 1513.980000 1.860000 ;
      RECT 1514.315000  1.355000 1514.685000 1.685000 ;
      RECT 1514.435000  2.245000 1515.430000 2.415000 ;
      RECT 1514.610000  0.275000 1515.435000 0.445000 ;
      RECT 1514.875000  0.785000 1515.095000 1.115000 ;
      RECT 1514.895000  1.355000 1515.115000 1.685000 ;
      RECT 1514.895000  1.685000 1515.090000 1.860000 ;
      RECT 1515.260000  1.825000 1516.245000 1.995000 ;
      RECT 1515.260000  1.995000 1515.430000 2.245000 ;
      RECT 1515.265000  0.445000 1515.435000 0.715000 ;
      RECT 1515.265000  0.715000 1516.245000 0.885000 ;
      RECT 1515.375000  1.055000 1515.905000 1.655000 ;
      RECT 1515.650000  2.165000 1515.820000 2.635000 ;
      RECT 1515.655000  0.085000 1515.855000 0.545000 ;
      RECT 1516.075000  0.365000 1516.425000 0.535000 ;
      RECT 1516.075000  0.535000 1516.245000 0.715000 ;
      RECT 1516.075000  0.885000 1516.245000 1.825000 ;
      RECT 1516.075000  1.995000 1516.245000 2.070000 ;
      RECT 1516.075000  2.070000 1516.360000 2.440000 ;
      RECT 1516.415000  0.705000 1517.045000 1.035000 ;
      RECT 1516.415000  1.035000 1516.705000 1.905000 ;
      RECT 1516.555000  2.190000 1517.775000 2.360000 ;
      RECT 1516.645000  0.365000 1517.435000 0.535000 ;
      RECT 1516.895000  1.655000 1517.385000 2.010000 ;
      RECT 1517.265000  0.535000 1517.435000 1.315000 ;
      RECT 1517.265000  1.315000 1518.115000 1.485000 ;
      RECT 1517.555000  1.485000 1518.115000 1.575000 ;
      RECT 1517.555000  1.575000 1517.775000 2.190000 ;
      RECT 1517.655000  0.765000 1518.505000 1.065000 ;
      RECT 1517.655000  1.065000 1517.825000 1.095000 ;
      RECT 1517.735000  0.085000 1518.105000 0.585000 ;
      RECT 1517.945000  1.245000 1518.115000 1.315000 ;
      RECT 1517.945000  1.835000 1518.115000 2.635000 ;
      RECT 1518.285000  0.365000 1518.795000 0.535000 ;
      RECT 1518.285000  0.535000 1518.505000 0.765000 ;
      RECT 1518.285000  1.065000 1518.505000 2.135000 ;
      RECT 1518.285000  2.135000 1518.585000 2.465000 ;
      RECT 1518.675000  0.705000 1519.275000 1.035000 ;
      RECT 1518.675000  1.245000 1518.915000 1.965000 ;
      RECT 1518.810000  2.165000 1519.845000 2.335000 ;
      RECT 1519.075000  0.365000 1519.715000 0.535000 ;
      RECT 1519.085000  1.035000 1519.275000 1.575000 ;
      RECT 1519.085000  1.575000 1519.455000 1.905000 ;
      RECT 1519.495000  0.535000 1519.715000 0.995000 ;
      RECT 1519.495000  0.995000 1520.605000 1.325000 ;
      RECT 1519.495000  1.325000 1519.845000 1.405000 ;
      RECT 1519.675000  1.405000 1519.845000 2.165000 ;
      RECT 1519.940000  0.085000 1520.360000 0.615000 ;
      RECT 1520.045000  1.575000 1520.960000 1.905000 ;
      RECT 1520.075000  2.135000 1520.380000 2.635000 ;
      RECT 1520.630000  0.300000 1520.960000 0.825000 ;
      RECT 1520.670000  1.905000 1520.960000 2.455000 ;
      RECT 1520.775000  0.825000 1520.960000 0.995000 ;
      RECT 1520.775000  0.995000 1521.610000 1.325000 ;
      RECT 1520.775000  1.325000 1520.960000 1.575000 ;
      RECT 1521.180000  0.085000 1521.350000 0.695000 ;
      RECT 1521.180000  1.625000 1521.350000 2.635000 ;
      RECT 1521.520000  0.305000 1522.000000 0.825000 ;
      RECT 1521.540000  1.505000 1522.000000 2.465000 ;
      RECT 1521.780000  0.825000 1522.000000 1.505000 ;
      RECT 1522.170000  0.345000 1522.420000 0.995000 ;
      RECT 1522.170000  0.995000 1523.000000 1.325000 ;
      RECT 1522.170000  1.325000 1522.420000 2.425000 ;
      RECT 1522.625000  0.085000 1522.955000 0.805000 ;
      RECT 1522.650000  1.495000 1522.955000 2.635000 ;
      RECT 1523.175000  0.265000 1523.430000 2.325000 ;
      RECT 1523.605000  0.085000 1523.895000 0.810000 ;
      RECT 1523.605000  1.470000 1523.895000 2.635000 ;
      RECT 1524.075000  0.975000 1524.425000 1.625000 ;
      RECT 1524.155000  0.345000 1524.325000 0.635000 ;
      RECT 1524.155000  0.635000 1524.840000 0.805000 ;
      RECT 1524.155000  1.795000 1524.875000 1.965000 ;
      RECT 1524.155000  1.965000 1524.325000 2.465000 ;
      RECT 1524.495000  0.085000 1524.875000 0.465000 ;
      RECT 1524.495000  2.135000 1524.875000 2.635000 ;
      RECT 1524.645000  0.805000 1524.840000 0.970000 ;
      RECT 1524.645000  0.970000 1524.875000 1.795000 ;
      RECT 1525.095000  0.345000 1525.265000 2.465000 ;
      RECT 1525.500000  0.255000 1525.885000 0.445000 ;
      RECT 1525.500000  0.445000 1525.670000 1.860000 ;
      RECT 1525.500000  1.860000 1527.510000 2.075000 ;
      RECT 1525.500000  2.075000 1525.785000 2.445000 ;
      RECT 1525.840000  0.615000 1527.515000 0.785000 ;
      RECT 1525.840000  0.785000 1526.010000 1.685000 ;
      RECT 1525.955000  2.245000 1526.335000 2.635000 ;
      RECT 1526.125000  0.085000 1526.455000 0.445000 ;
      RECT 1526.230000  0.955000 1526.675000 1.125000 ;
      RECT 1526.230000  1.125000 1526.400000 1.860000 ;
      RECT 1526.735000  1.355000 1527.105000 1.685000 ;
      RECT 1526.855000  2.245000 1527.850000 2.415000 ;
      RECT 1527.030000  0.275000 1527.855000 0.445000 ;
      RECT 1527.295000  0.785000 1527.515000 1.115000 ;
      RECT 1527.315000  1.355000 1527.535000 1.685000 ;
      RECT 1527.315000  1.685000 1527.510000 1.860000 ;
      RECT 1527.680000  1.825000 1528.665000 1.995000 ;
      RECT 1527.680000  1.995000 1527.850000 2.245000 ;
      RECT 1527.685000  0.445000 1527.855000 0.715000 ;
      RECT 1527.685000  0.715000 1528.665000 0.885000 ;
      RECT 1527.795000  1.055000 1528.325000 1.655000 ;
      RECT 1528.070000  2.165000 1528.240000 2.635000 ;
      RECT 1528.075000  0.085000 1528.275000 0.545000 ;
      RECT 1528.495000  0.365000 1528.845000 0.535000 ;
      RECT 1528.495000  0.535000 1528.665000 0.715000 ;
      RECT 1528.495000  0.885000 1528.665000 1.825000 ;
      RECT 1528.495000  1.995000 1528.665000 2.070000 ;
      RECT 1528.495000  2.070000 1528.780000 2.440000 ;
      RECT 1528.835000  0.705000 1529.465000 1.035000 ;
      RECT 1528.835000  1.035000 1529.125000 1.905000 ;
      RECT 1528.975000  2.190000 1530.195000 2.360000 ;
      RECT 1529.065000  0.365000 1529.855000 0.535000 ;
      RECT 1529.315000  1.655000 1529.805000 2.010000 ;
      RECT 1529.685000  0.535000 1529.855000 1.315000 ;
      RECT 1529.685000  1.315000 1530.535000 1.485000 ;
      RECT 1529.975000  1.485000 1530.535000 1.575000 ;
      RECT 1529.975000  1.575000 1530.195000 2.190000 ;
      RECT 1530.075000  0.765000 1530.925000 1.065000 ;
      RECT 1530.075000  1.065000 1530.245000 1.095000 ;
      RECT 1530.155000  0.085000 1530.525000 0.585000 ;
      RECT 1530.365000  1.245000 1530.535000 1.315000 ;
      RECT 1530.365000  1.835000 1530.535000 2.635000 ;
      RECT 1530.705000  0.365000 1531.215000 0.535000 ;
      RECT 1530.705000  0.535000 1530.925000 0.765000 ;
      RECT 1530.705000  1.065000 1530.925000 2.135000 ;
      RECT 1530.705000  2.135000 1531.005000 2.465000 ;
      RECT 1531.095000  0.705000 1531.695000 1.035000 ;
      RECT 1531.095000  1.245000 1531.335000 1.965000 ;
      RECT 1531.230000  2.165000 1532.265000 2.335000 ;
      RECT 1531.495000  0.365000 1532.135000 0.535000 ;
      RECT 1531.505000  1.035000 1531.695000 1.575000 ;
      RECT 1531.505000  1.575000 1531.875000 1.905000 ;
      RECT 1531.915000  0.535000 1532.135000 0.995000 ;
      RECT 1531.915000  0.995000 1533.025000 1.325000 ;
      RECT 1531.915000  1.325000 1532.265000 1.405000 ;
      RECT 1532.095000  1.405000 1532.265000 2.165000 ;
      RECT 1532.360000  0.085000 1532.780000 0.615000 ;
      RECT 1532.465000  1.575000 1533.380000 1.905000 ;
      RECT 1532.495000  2.135000 1532.800000 2.635000 ;
      RECT 1533.015000  0.300000 1533.380000 0.825000 ;
      RECT 1533.050000  1.905000 1533.380000 2.455000 ;
      RECT 1533.195000  0.825000 1533.380000 0.995000 ;
      RECT 1533.195000  0.995000 1533.980000 1.325000 ;
      RECT 1533.195000  1.325000 1533.380000 1.575000 ;
      RECT 1533.550000  0.085000 1533.970000 0.695000 ;
      RECT 1533.550000  1.625000 1533.970000 2.635000 ;
      RECT 1534.190000  0.255000 1534.470000 2.455000 ;
      RECT 1534.660000  0.085000 1534.890000 0.690000 ;
      RECT 1534.670000  1.615000 1534.840000 2.635000 ;
      RECT 1535.110000  0.345000 1535.360000 0.995000 ;
      RECT 1535.110000  0.995000 1536.320000 1.325000 ;
      RECT 1535.110000  1.325000 1535.440000 2.425000 ;
      RECT 1535.645000  0.085000 1536.275000 0.805000 ;
      RECT 1535.670000  1.495000 1536.275000 2.635000 ;
      RECT 1536.495000  0.265000 1536.765000 2.325000 ;
      RECT 1536.965000  0.085000 1537.135000 0.955000 ;
      RECT 1536.965000  1.395000 1537.135000 2.635000 ;
      RECT 1537.405000  0.085000 1537.695000 0.810000 ;
      RECT 1537.405000  1.470000 1537.695000 2.635000 ;
      RECT 1537.875000  0.975000 1538.225000 1.625000 ;
      RECT 1537.955000  0.345000 1538.125000 0.635000 ;
      RECT 1537.955000  0.635000 1538.675000 0.805000 ;
      RECT 1537.960000  1.795000 1538.675000 1.965000 ;
      RECT 1537.960000  1.965000 1538.130000 2.465000 ;
      RECT 1538.295000  0.085000 1538.675000 0.465000 ;
      RECT 1538.300000  2.135000 1538.680000 2.635000 ;
      RECT 1538.445000  0.805000 1538.675000 1.795000 ;
      RECT 1538.895000  0.345000 1539.125000 2.465000 ;
      RECT 1539.315000  0.275000 1539.685000 0.445000 ;
      RECT 1539.315000  0.445000 1539.485000 1.860000 ;
      RECT 1539.315000  1.860000 1541.320000 2.075000 ;
      RECT 1539.315000  2.075000 1539.590000 2.445000 ;
      RECT 1539.660000  0.615000 1541.285000 0.785000 ;
      RECT 1539.660000  0.785000 1539.995000 1.685000 ;
      RECT 1539.760000  2.245000 1540.140000 2.635000 ;
      RECT 1539.855000  0.085000 1540.185000 0.445000 ;
      RECT 1540.165000  0.955000 1540.495000 1.125000 ;
      RECT 1540.165000  1.125000 1540.335000 1.860000 ;
      RECT 1540.525000  1.355000 1540.930000 1.685000 ;
      RECT 1540.675000  2.245000 1541.670000 2.415000 ;
      RECT 1540.850000  0.275000 1541.675000 0.445000 ;
      RECT 1541.110000  1.355000 1541.320000 1.860000 ;
      RECT 1541.115000  0.785000 1541.285000 1.115000 ;
      RECT 1541.500000  1.825000 1542.515000 1.995000 ;
      RECT 1541.500000  1.995000 1541.670000 2.245000 ;
      RECT 1541.505000  0.445000 1541.675000 0.695000 ;
      RECT 1541.505000  0.695000 1542.515000 0.865000 ;
      RECT 1541.505000  1.035000 1541.875000 1.655000 ;
      RECT 1541.890000  2.165000 1542.060000 2.635000 ;
      RECT 1541.895000  0.085000 1542.095000 0.525000 ;
      RECT 1542.345000  0.365000 1542.695000 0.535000 ;
      RECT 1542.345000  0.535000 1542.515000 0.695000 ;
      RECT 1542.345000  0.865000 1542.515000 1.825000 ;
      RECT 1542.345000  1.995000 1542.515000 2.065000 ;
      RECT 1542.345000  2.065000 1542.580000 2.440000 ;
      RECT 1542.685000  0.705000 1543.315000 1.035000 ;
      RECT 1542.685000  1.035000 1542.975000 1.905000 ;
      RECT 1542.825000  2.190000 1544.010000 2.360000 ;
      RECT 1542.915000  0.365000 1543.655000 0.535000 ;
      RECT 1543.165000  1.655000 1543.655000 2.010000 ;
      RECT 1543.485000  0.535000 1543.655000 1.315000 ;
      RECT 1543.485000  1.315000 1544.465000 1.485000 ;
      RECT 1543.825000  0.765000 1544.840000 1.095000 ;
      RECT 1543.825000  1.485000 1544.465000 1.575000 ;
      RECT 1543.825000  1.575000 1544.010000 2.190000 ;
      RECT 1544.005000  0.085000 1544.375000 0.585000 ;
      RECT 1544.180000  1.835000 1544.350000 2.635000 ;
      RECT 1544.555000  0.365000 1545.040000 0.535000 ;
      RECT 1544.555000  0.535000 1544.840000 0.765000 ;
      RECT 1544.635000  1.095000 1544.840000 2.465000 ;
      RECT 1545.010000  1.245000 1545.250000 1.965000 ;
      RECT 1545.030000  0.705000 1545.725000 1.035000 ;
      RECT 1545.030000  2.165000 1546.065000 2.335000 ;
      RECT 1545.235000  0.365000 1546.065000 0.535000 ;
      RECT 1545.515000  1.035000 1545.725000 1.905000 ;
      RECT 1545.895000  0.535000 1546.065000 0.995000 ;
      RECT 1545.895000  0.995000 1546.830000 1.325000 ;
      RECT 1545.895000  1.325000 1546.065000 2.165000 ;
      RECT 1546.235000  0.085000 1546.550000 0.615000 ;
      RECT 1546.235000  1.575000 1547.185000 1.905000 ;
      RECT 1546.245000  2.135000 1546.550000 2.635000 ;
      RECT 1546.820000  0.300000 1547.180000 0.825000 ;
      RECT 1546.900000  1.905000 1547.185000 2.455000 ;
      RECT 1547.000000  0.825000 1547.180000 0.995000 ;
      RECT 1547.000000  0.995000 1547.810000 1.325000 ;
      RECT 1547.000000  1.325000 1547.185000 1.575000 ;
      RECT 1547.370000  0.085000 1547.540000 0.695000 ;
      RECT 1547.370000  1.625000 1547.540000 2.635000 ;
      RECT 1547.710000  0.305000 1548.250000 0.820000 ;
      RECT 1547.710000  1.545000 1548.250000 2.395000 ;
      RECT 1548.010000  0.820000 1548.250000 1.545000 ;
      RECT 1548.445000  0.085000 1548.735000 0.810000 ;
      RECT 1548.445000  1.470000 1548.735000 2.635000 ;
      RECT 1548.915000  0.975000 1549.265000 1.625000 ;
      RECT 1548.995000  0.345000 1549.165000 0.635000 ;
      RECT 1548.995000  0.635000 1549.715000 0.805000 ;
      RECT 1549.000000  1.795000 1549.715000 1.965000 ;
      RECT 1549.000000  1.965000 1549.170000 2.465000 ;
      RECT 1549.335000  0.085000 1549.715000 0.465000 ;
      RECT 1549.340000  2.135000 1549.720000 2.635000 ;
      RECT 1549.485000  0.805000 1549.715000 1.795000 ;
      RECT 1549.935000  0.345000 1550.165000 2.465000 ;
      RECT 1550.355000  0.275000 1550.725000 0.445000 ;
      RECT 1550.355000  0.445000 1550.525000 1.860000 ;
      RECT 1550.355000  1.860000 1552.345000 2.075000 ;
      RECT 1550.355000  2.075000 1550.630000 2.445000 ;
      RECT 1550.700000  0.615000 1552.325000 0.785000 ;
      RECT 1550.700000  0.785000 1551.035000 1.685000 ;
      RECT 1550.800000  2.245000 1551.180000 2.635000 ;
      RECT 1550.945000  0.085000 1551.275000 0.445000 ;
      RECT 1551.205000  0.955000 1551.535000 1.125000 ;
      RECT 1551.205000  1.125000 1551.375000 1.860000 ;
      RECT 1551.565000  1.355000 1551.970000 1.685000 ;
      RECT 1551.715000  2.245000 1552.710000 2.415000 ;
      RECT 1551.890000  0.275000 1552.715000 0.445000 ;
      RECT 1552.150000  1.355000 1552.345000 1.860000 ;
      RECT 1552.155000  0.785000 1552.325000 1.115000 ;
      RECT 1552.540000  1.825000 1553.555000 1.995000 ;
      RECT 1552.540000  1.995000 1552.710000 2.245000 ;
      RECT 1552.545000  0.445000 1552.715000 0.695000 ;
      RECT 1552.545000  0.695000 1553.555000 0.865000 ;
      RECT 1552.545000  1.035000 1552.915000 1.655000 ;
      RECT 1552.930000  2.165000 1553.100000 2.635000 ;
      RECT 1552.935000  0.085000 1553.135000 0.525000 ;
      RECT 1553.385000  0.365000 1553.735000 0.535000 ;
      RECT 1553.385000  0.535000 1553.555000 0.695000 ;
      RECT 1553.385000  0.865000 1553.555000 1.825000 ;
      RECT 1553.385000  1.995000 1553.555000 2.065000 ;
      RECT 1553.385000  2.065000 1553.620000 2.440000 ;
      RECT 1553.725000  0.705000 1554.355000 1.035000 ;
      RECT 1553.725000  1.035000 1554.015000 1.905000 ;
      RECT 1553.865000  2.190000 1555.085000 2.360000 ;
      RECT 1553.955000  0.365000 1554.715000 0.535000 ;
      RECT 1554.205000  1.655000 1554.695000 2.010000 ;
      RECT 1554.545000  0.535000 1554.715000 1.245000 ;
      RECT 1554.545000  1.245000 1555.425000 1.485000 ;
      RECT 1554.865000  1.485000 1555.425000 1.575000 ;
      RECT 1554.865000  1.575000 1555.085000 2.190000 ;
      RECT 1554.885000  0.765000 1555.815000 1.065000 ;
      RECT 1555.045000  0.085000 1555.415000 0.585000 ;
      RECT 1555.255000  1.835000 1555.425000 2.635000 ;
      RECT 1555.595000  0.365000 1556.105000 0.535000 ;
      RECT 1555.595000  0.535000 1555.815000 0.765000 ;
      RECT 1555.595000  1.065000 1555.815000 2.135000 ;
      RECT 1555.595000  2.135000 1555.895000 2.465000 ;
      RECT 1555.985000  0.705000 1556.585000 1.035000 ;
      RECT 1555.985000  1.245000 1556.225000 1.965000 ;
      RECT 1556.120000  2.165000 1557.155000 2.335000 ;
      RECT 1556.385000  0.365000 1557.025000 0.535000 ;
      RECT 1556.395000  1.035000 1556.585000 1.575000 ;
      RECT 1556.395000  1.575000 1556.765000 1.905000 ;
      RECT 1556.805000  0.535000 1557.025000 0.995000 ;
      RECT 1556.805000  0.995000 1557.970000 1.325000 ;
      RECT 1556.805000  1.325000 1557.155000 1.405000 ;
      RECT 1556.985000  1.405000 1557.155000 2.165000 ;
      RECT 1557.270000  0.085000 1557.690000 0.615000 ;
      RECT 1557.375000  1.575000 1558.325000 1.905000 ;
      RECT 1557.385000  2.135000 1557.690000 2.635000 ;
      RECT 1557.960000  0.300000 1558.320000 0.825000 ;
      RECT 1558.040000  1.905000 1558.325000 2.455000 ;
      RECT 1558.140000  0.825000 1558.320000 0.995000 ;
      RECT 1558.140000  0.995000 1558.950000 1.325000 ;
      RECT 1558.140000  1.325000 1558.325000 1.575000 ;
      RECT 1558.510000  0.085000 1558.680000 0.695000 ;
      RECT 1558.510000  1.625000 1558.680000 2.635000 ;
      RECT 1558.850000  0.305000 1559.320000 0.820000 ;
      RECT 1558.850000  1.545000 1559.320000 2.395000 ;
      RECT 1559.150000  0.820000 1559.320000 1.545000 ;
      RECT 1559.490000  0.085000 1559.660000 0.565000 ;
      RECT 1559.490000  1.845000 1559.660000 2.635000 ;
      RECT 1559.945000  0.085000 1560.235000 0.810000 ;
      RECT 1559.945000  1.470000 1560.235000 2.635000 ;
      RECT 1560.415000  0.975000 1560.765000 1.625000 ;
      RECT 1560.495000  0.345000 1560.665000 0.635000 ;
      RECT 1560.495000  0.635000 1561.215000 0.805000 ;
      RECT 1560.500000  1.795000 1561.215000 1.965000 ;
      RECT 1560.500000  1.965000 1560.670000 2.465000 ;
      RECT 1560.835000  0.085000 1561.215000 0.465000 ;
      RECT 1560.840000  2.135000 1561.220000 2.635000 ;
      RECT 1560.985000  0.805000 1561.215000 1.795000 ;
      RECT 1561.435000  0.345000 1561.665000 2.465000 ;
      RECT 1561.855000  0.275000 1562.225000 0.445000 ;
      RECT 1561.855000  0.445000 1562.025000 1.860000 ;
      RECT 1561.855000  1.860000 1563.845000 2.075000 ;
      RECT 1561.855000  2.075000 1562.130000 2.445000 ;
      RECT 1562.200000  0.615000 1563.825000 0.785000 ;
      RECT 1562.200000  0.785000 1562.535000 1.685000 ;
      RECT 1562.300000  2.245000 1562.680000 2.635000 ;
      RECT 1562.445000  0.085000 1562.775000 0.445000 ;
      RECT 1562.705000  0.955000 1563.035000 1.125000 ;
      RECT 1562.705000  1.125000 1562.875000 1.860000 ;
      RECT 1563.065000  1.355000 1563.470000 1.685000 ;
      RECT 1563.215000  2.245000 1564.210000 2.415000 ;
      RECT 1563.390000  0.275000 1564.215000 0.445000 ;
      RECT 1563.650000  1.355000 1563.845000 1.860000 ;
      RECT 1563.655000  0.785000 1563.825000 1.115000 ;
      RECT 1564.040000  1.825000 1565.055000 1.995000 ;
      RECT 1564.040000  1.995000 1564.210000 2.245000 ;
      RECT 1564.045000  0.445000 1564.215000 0.695000 ;
      RECT 1564.045000  0.695000 1565.055000 0.865000 ;
      RECT 1564.045000  1.035000 1564.415000 1.655000 ;
      RECT 1564.430000  2.165000 1564.600000 2.635000 ;
      RECT 1564.435000  0.085000 1564.635000 0.525000 ;
      RECT 1564.885000  0.365000 1565.235000 0.535000 ;
      RECT 1564.885000  0.535000 1565.055000 0.695000 ;
      RECT 1564.885000  0.865000 1565.055000 1.825000 ;
      RECT 1564.885000  1.995000 1565.055000 2.065000 ;
      RECT 1564.885000  2.065000 1565.120000 2.440000 ;
      RECT 1565.225000  0.705000 1565.855000 1.035000 ;
      RECT 1565.225000  1.035000 1565.515000 1.905000 ;
      RECT 1565.365000  2.190000 1566.585000 2.360000 ;
      RECT 1565.455000  0.365000 1566.215000 0.535000 ;
      RECT 1565.705000  1.655000 1566.195000 2.010000 ;
      RECT 1566.045000  0.535000 1566.215000 1.245000 ;
      RECT 1566.045000  1.245000 1566.925000 1.485000 ;
      RECT 1566.365000  1.485000 1566.925000 1.575000 ;
      RECT 1566.365000  1.575000 1566.585000 2.190000 ;
      RECT 1566.385000  0.765000 1567.315000 1.065000 ;
      RECT 1566.545000  0.085000 1566.915000 0.585000 ;
      RECT 1566.755000  1.835000 1566.925000 2.635000 ;
      RECT 1567.095000  0.365000 1567.605000 0.535000 ;
      RECT 1567.095000  0.535000 1567.315000 0.765000 ;
      RECT 1567.095000  1.065000 1567.315000 2.135000 ;
      RECT 1567.095000  2.135000 1567.395000 2.465000 ;
      RECT 1567.485000  0.705000 1568.085000 1.035000 ;
      RECT 1567.485000  1.245000 1567.725000 1.965000 ;
      RECT 1567.620000  2.165000 1568.655000 2.335000 ;
      RECT 1567.885000  0.365000 1568.525000 0.535000 ;
      RECT 1567.895000  1.035000 1568.085000 1.575000 ;
      RECT 1567.895000  1.575000 1568.265000 1.905000 ;
      RECT 1568.305000  0.535000 1568.525000 0.995000 ;
      RECT 1568.305000  0.995000 1569.470000 1.325000 ;
      RECT 1568.305000  1.325000 1568.655000 1.405000 ;
      RECT 1568.485000  1.405000 1568.655000 2.165000 ;
      RECT 1568.770000  0.085000 1569.190000 0.615000 ;
      RECT 1568.875000  1.575000 1569.825000 1.905000 ;
      RECT 1568.885000  2.135000 1569.190000 2.635000 ;
      RECT 1569.460000  0.300000 1569.820000 0.825000 ;
      RECT 1569.540000  1.905000 1569.825000 2.455000 ;
      RECT 1569.640000  0.825000 1569.820000 1.075000 ;
      RECT 1569.640000  1.075000 1571.700000 1.325000 ;
      RECT 1569.640000  1.325000 1569.825000 1.575000 ;
      RECT 1570.010000  0.085000 1570.180000 0.695000 ;
      RECT 1570.010000  1.625000 1570.180000 2.635000 ;
      RECT 1570.350000  0.305000 1570.730000 0.735000 ;
      RECT 1570.350000  0.735000 1572.170000 0.905000 ;
      RECT 1570.350000  1.505000 1572.170000 1.675000 ;
      RECT 1570.350000  1.675000 1570.730000 2.395000 ;
      RECT 1570.960000  0.085000 1571.130000 0.565000 ;
      RECT 1570.960000  1.845000 1571.130000 2.635000 ;
      RECT 1571.300000  0.305000 1571.680000 0.735000 ;
      RECT 1571.300000  1.675000 1571.680000 2.395000 ;
      RECT 1571.870000  0.905000 1572.170000 1.505000 ;
      RECT 1571.900000  0.085000 1572.070000 0.565000 ;
      RECT 1571.900000  1.845000 1572.070000 2.635000 ;
      RECT 1572.365000  0.085000 1572.655000 0.810000 ;
      RECT 1572.365000  1.470000 1572.655000 2.635000 ;
      RECT 1572.825000  0.255000 1573.085000 0.615000 ;
      RECT 1572.825000  0.615000 1574.035000 0.785000 ;
      RECT 1572.825000  0.955000 1573.070000 1.665000 ;
      RECT 1572.825000  1.835000 1573.085000 2.635000 ;
      RECT 1573.255000  0.085000 1573.635000 0.445000 ;
      RECT 1573.255000  0.785000 1573.425000 2.125000 ;
      RECT 1573.255000  2.125000 1574.020000 2.465000 ;
      RECT 1573.595000  0.955000 1573.975000 1.955000 ;
      RECT 1573.855000  0.255000 1574.035000 0.615000 ;
      RECT 1574.205000  0.255000 1575.385000 0.535000 ;
      RECT 1574.205000  0.705000 1574.540000 1.205000 ;
      RECT 1574.205000  1.205000 1574.700000 1.955000 ;
      RECT 1574.350000  2.125000 1575.040000 2.465000 ;
      RECT 1574.710000  0.705000 1575.045000 1.035000 ;
      RECT 1574.870000  1.205000 1575.945000 1.375000 ;
      RECT 1574.870000  1.375000 1575.040000 2.125000 ;
      RECT 1575.210000  1.575000 1575.405000 1.635000 ;
      RECT 1575.210000  1.635000 1576.285000 1.905000 ;
      RECT 1575.215000  0.535000 1575.385000 0.995000 ;
      RECT 1575.215000  0.995000 1575.945000 1.205000 ;
      RECT 1575.260000  2.075000 1575.845000 2.635000 ;
      RECT 1575.650000  0.085000 1575.820000 0.825000 ;
      RECT 1576.065000  1.905000 1576.285000 1.915000 ;
      RECT 1576.065000  1.915000 1578.475000 2.085000 ;
      RECT 1576.065000  2.085000 1576.285000 2.465000 ;
      RECT 1576.115000  0.255000 1576.285000 1.635000 ;
      RECT 1576.475000  0.255000 1576.805000 0.935000 ;
      RECT 1576.475000  0.935000 1576.645000 1.575000 ;
      RECT 1576.475000  1.575000 1576.885000 1.745000 ;
      RECT 1576.625000  2.255000 1578.475000 2.635000 ;
      RECT 1576.815000  1.105000 1577.290000 1.275000 ;
      RECT 1577.025000  0.085000 1577.355000 0.445000 ;
      RECT 1577.105000  1.275000 1577.290000 1.495000 ;
      RECT 1577.105000  1.495000 1577.955000 1.745000 ;
      RECT 1577.120000  0.615000 1577.955000 0.785000 ;
      RECT 1577.120000  0.785000 1577.290000 1.105000 ;
      RECT 1577.485000  0.995000 1577.800000 1.325000 ;
      RECT 1577.705000  0.255000 1577.955000 0.615000 ;
      RECT 1578.125000  0.995000 1578.475000 1.915000 ;
      RECT 1578.275000  0.255000 1578.445000 0.615000 ;
      RECT 1578.275000  0.615000 1579.555000 0.785000 ;
      RECT 1578.695000  0.995000 1579.135000 1.325000 ;
      RECT 1578.695000  1.495000 1579.555000 2.085000 ;
      RECT 1578.695000  2.085000 1578.865000 2.465000 ;
      RECT 1579.065000  0.085000 1579.425000 0.445000 ;
      RECT 1579.125000  2.255000 1579.455000 2.635000 ;
      RECT 1579.385000  0.785000 1579.555000 1.495000 ;
      RECT 1579.725000  0.255000 1579.975000 2.465000 ;
      RECT 1580.185000  0.085000 1580.475000 0.810000 ;
      RECT 1580.185000  1.470000 1580.475000 2.635000 ;
      RECT 1580.645000  0.255000 1580.905000 0.615000 ;
      RECT 1580.645000  0.615000 1581.855000 0.785000 ;
      RECT 1580.645000  0.955000 1580.890000 1.665000 ;
      RECT 1580.645000  1.835000 1580.905000 2.635000 ;
      RECT 1581.075000  0.085000 1581.455000 0.445000 ;
      RECT 1581.075000  0.785000 1581.280000 2.125000 ;
      RECT 1581.075000  2.125000 1581.840000 2.465000 ;
      RECT 1581.450000  0.955000 1581.855000 1.955000 ;
      RECT 1581.675000  0.255000 1581.855000 0.615000 ;
      RECT 1582.025000  0.255000 1583.205000 0.535000 ;
      RECT 1582.025000  0.705000 1582.360000 1.205000 ;
      RECT 1582.025000  1.205000 1582.520000 1.955000 ;
      RECT 1582.170000  2.125000 1582.860000 2.465000 ;
      RECT 1582.530000  0.705000 1582.865000 1.035000 ;
      RECT 1582.690000  1.205000 1583.765000 1.375000 ;
      RECT 1582.690000  1.375000 1582.860000 2.125000 ;
      RECT 1583.030000  1.575000 1583.225000 1.635000 ;
      RECT 1583.030000  1.635000 1584.105000 1.905000 ;
      RECT 1583.035000  0.535000 1583.205000 0.995000 ;
      RECT 1583.035000  0.995000 1583.765000 1.205000 ;
      RECT 1583.080000  2.075000 1583.665000 2.635000 ;
      RECT 1583.470000  0.085000 1583.640000 0.825000 ;
      RECT 1583.885000  1.905000 1584.105000 1.915000 ;
      RECT 1583.885000  1.915000 1586.315000 2.085000 ;
      RECT 1583.885000  2.085000 1584.105000 2.465000 ;
      RECT 1583.935000  0.255000 1584.105000 1.635000 ;
      RECT 1584.295000  0.255000 1584.625000 0.765000 ;
      RECT 1584.295000  0.765000 1584.720000 0.935000 ;
      RECT 1584.295000  0.935000 1584.465000 1.575000 ;
      RECT 1584.295000  1.575000 1584.705000 1.745000 ;
      RECT 1584.445000  2.255000 1586.315000 2.635000 ;
      RECT 1584.635000  1.105000 1585.230000 1.275000 ;
      RECT 1584.845000  0.085000 1585.175000 0.445000 ;
      RECT 1584.925000  1.275000 1585.230000 1.495000 ;
      RECT 1584.925000  1.495000 1585.775000 1.745000 ;
      RECT 1584.940000  0.615000 1585.645000 0.785000 ;
      RECT 1584.940000  0.785000 1585.230000 1.105000 ;
      RECT 1585.395000  0.255000 1585.645000 0.615000 ;
      RECT 1585.525000  0.995000 1585.745000 1.325000 ;
      RECT 1585.965000  0.995000 1586.315000 1.915000 ;
      RECT 1586.065000  0.255000 1586.235000 0.615000 ;
      RECT 1586.065000  0.615000 1587.310000 0.785000 ;
      RECT 1586.535000  0.995000 1586.965000 1.325000 ;
      RECT 1586.535000  1.495000 1587.310000 2.085000 ;
      RECT 1586.535000  2.085000 1586.705000 2.465000 ;
      RECT 1586.895000  0.085000 1587.230000 0.445000 ;
      RECT 1586.955000  2.255000 1587.285000 2.635000 ;
      RECT 1587.140000  0.785000 1587.310000 1.055000 ;
      RECT 1587.140000  1.055000 1587.830000 1.315000 ;
      RECT 1587.140000  1.315000 1587.310000 1.495000 ;
      RECT 1587.400000  0.255000 1587.730000 0.445000 ;
      RECT 1587.530000  0.445000 1587.730000 0.715000 ;
      RECT 1587.530000  0.715000 1588.235000 0.885000 ;
      RECT 1587.530000  1.485000 1588.235000 1.655000 ;
      RECT 1587.530000  1.655000 1587.780000 2.465000 ;
      RECT 1587.950000  0.085000 1588.120000 0.545000 ;
      RECT 1588.000000  1.825000 1588.250000 2.635000 ;
      RECT 1588.050000  0.885000 1588.235000 1.485000 ;
      RECT 1588.465000  0.085000 1588.755000 0.810000 ;
      RECT 1588.465000  1.470000 1588.755000 2.635000 ;
      RECT 1588.925000  0.255000 1589.185000 0.615000 ;
      RECT 1588.925000  0.615000 1590.135000 0.785000 ;
      RECT 1588.925000  0.955000 1589.185000 1.665000 ;
      RECT 1588.925000  1.835000 1589.185000 2.635000 ;
      RECT 1589.355000  0.085000 1589.735000 0.445000 ;
      RECT 1589.355000  0.785000 1589.575000 2.125000 ;
      RECT 1589.355000  2.125000 1590.200000 2.465000 ;
      RECT 1589.745000  0.955000 1590.135000 1.445000 ;
      RECT 1589.745000  1.445000 1590.180000 1.955000 ;
      RECT 1589.955000  0.255000 1590.135000 0.615000 ;
      RECT 1590.305000  0.255000 1591.540000 0.535000 ;
      RECT 1590.305000  0.705000 1590.695000 1.205000 ;
      RECT 1590.305000  1.205000 1590.855000 1.325000 ;
      RECT 1590.350000  1.325000 1590.855000 1.955000 ;
      RECT 1590.370000  2.125000 1591.245000 2.465000 ;
      RECT 1590.865000  0.705000 1591.200000 1.035000 ;
      RECT 1591.075000  1.205000 1592.105000 1.375000 ;
      RECT 1591.075000  1.375000 1591.245000 2.125000 ;
      RECT 1591.370000  0.535000 1591.540000 0.995000 ;
      RECT 1591.370000  0.995000 1592.105000 1.205000 ;
      RECT 1591.415000  1.575000 1591.635000 1.635000 ;
      RECT 1591.415000  1.635000 1592.545000 1.905000 ;
      RECT 1591.415000  2.075000 1592.105000 2.635000 ;
      RECT 1591.760000  0.085000 1592.105000 0.825000 ;
      RECT 1592.325000  0.255000 1592.545000 1.635000 ;
      RECT 1592.325000  1.905000 1592.545000 1.915000 ;
      RECT 1592.325000  1.915000 1594.755000 2.085000 ;
      RECT 1592.325000  2.085000 1592.545000 2.465000 ;
      RECT 1592.735000  0.255000 1593.065000 0.765000 ;
      RECT 1592.735000  0.765000 1593.160000 0.935000 ;
      RECT 1592.735000  0.935000 1592.905000 1.575000 ;
      RECT 1592.735000  1.575000 1593.145000 1.745000 ;
      RECT 1592.735000  2.255000 1594.755000 2.635000 ;
      RECT 1593.075000  1.105000 1593.670000 1.275000 ;
      RECT 1593.235000  0.085000 1593.615000 0.445000 ;
      RECT 1593.365000  1.275000 1593.670000 1.495000 ;
      RECT 1593.365000  1.495000 1594.215000 1.745000 ;
      RECT 1593.380000  0.615000 1594.085000 0.785000 ;
      RECT 1593.380000  0.785000 1593.670000 1.105000 ;
      RECT 1593.835000  0.255000 1594.085000 0.615000 ;
      RECT 1593.895000  0.995000 1594.185000 1.325000 ;
      RECT 1594.255000  0.255000 1594.675000 0.615000 ;
      RECT 1594.255000  0.615000 1595.750000 0.785000 ;
      RECT 1594.405000  0.995000 1594.755000 1.915000 ;
      RECT 1594.845000  0.085000 1595.670000 0.445000 ;
      RECT 1594.975000  0.995000 1595.405000 1.325000 ;
      RECT 1594.975000  1.495000 1595.750000 2.085000 ;
      RECT 1594.975000  2.085000 1595.145000 2.465000 ;
      RECT 1595.395000  2.255000 1595.725000 2.635000 ;
      RECT 1595.580000  0.785000 1595.750000 1.055000 ;
      RECT 1595.580000  1.055000 1596.270000 1.315000 ;
      RECT 1595.580000  1.315000 1595.750000 1.495000 ;
      RECT 1595.840000  0.255000 1596.220000 0.445000 ;
      RECT 1595.970000  0.445000 1596.220000 0.715000 ;
      RECT 1595.970000  0.715000 1596.660000 0.885000 ;
      RECT 1595.970000  1.485000 1596.660000 1.655000 ;
      RECT 1595.970000  1.655000 1596.220000 2.465000 ;
      RECT 1596.440000  0.085000 1596.690000 0.545000 ;
      RECT 1596.440000  1.825000 1596.690000 2.635000 ;
      RECT 1596.490000  0.885000 1596.660000 1.055000 ;
      RECT 1596.490000  1.055000 1597.895000 1.315000 ;
      RECT 1596.490000  1.315000 1596.660000 1.485000 ;
      RECT 1597.045000  0.255000 1597.435000 1.055000 ;
      RECT 1597.045000  1.315000 1597.435000 2.465000 ;
      RECT 1597.605000  0.085000 1597.875000 0.885000 ;
      RECT 1597.605000  1.485000 1597.875000 2.635000 ;
      RECT 1598.125000  0.085000 1598.415000 0.810000 ;
      RECT 1598.125000  1.470000 1598.415000 2.635000 ;
      RECT 1598.595000  0.975000 1598.945000 1.625000 ;
      RECT 1598.675000  0.345000 1598.845000 0.635000 ;
      RECT 1598.675000  0.635000 1599.395000 0.805000 ;
      RECT 1598.675000  1.795000 1599.395000 1.965000 ;
      RECT 1598.675000  1.965000 1598.845000 2.465000 ;
      RECT 1599.015000  0.085000 1599.395000 0.465000 ;
      RECT 1599.015000  2.135000 1599.395000 2.635000 ;
      RECT 1599.165000  0.805000 1599.395000 1.795000 ;
      RECT 1599.615000  0.345000 1599.785000 2.465000 ;
      RECT 1599.955000  0.255000 1600.385000 0.515000 ;
      RECT 1599.955000  0.515000 1600.125000 1.890000 ;
      RECT 1599.955000  1.890000 1600.385000 2.465000 ;
      RECT 1600.295000  0.765000 1600.655000 1.720000 ;
      RECT 1600.825000  0.765000 1601.265000 1.185000 ;
      RECT 1600.825000  1.185000 1601.025000 1.370000 ;
      RECT 1600.885000  0.085000 1601.265000 0.515000 ;
      RECT 1600.885000  1.890000 1601.265000 2.635000 ;
      RECT 1601.195000  1.355000 1601.785000 1.720000 ;
      RECT 1601.455000  1.720000 1601.785000 2.425000 ;
      RECT 1601.480000  0.255000 1601.705000 0.845000 ;
      RECT 1601.480000  0.845000 1602.385000 1.175000 ;
      RECT 1601.480000  1.175000 1601.785000 1.355000 ;
      RECT 1601.885000  0.085000 1602.265000 0.610000 ;
      RECT 1602.015000  1.825000 1602.210000 2.635000 ;
      RECT 1602.605000  0.685000 1602.775000 1.320000 ;
      RECT 1602.605000  1.320000 1603.025000 1.650000 ;
      RECT 1602.925000  1.820000 1603.365000 2.020000 ;
      RECT 1602.925000  2.020000 1603.305000 2.465000 ;
      RECT 1602.945000  0.255000 1603.265000 0.980000 ;
      RECT 1602.945000  0.980000 1603.365000 1.150000 ;
      RECT 1603.195000  1.150000 1603.365000 1.820000 ;
      RECT 1603.495000  0.255000 1603.695000 0.645000 ;
      RECT 1603.495000  0.645000 1603.755000 0.825000 ;
      RECT 1603.535000  2.210000 1603.865000 2.465000 ;
      RECT 1603.585000  0.825000 1603.755000 1.785000 ;
      RECT 1603.585000  1.785000 1603.865000 2.210000 ;
      RECT 1603.865000  0.255000 1604.725000 0.515000 ;
      RECT 1604.105000  1.105000 1604.385000 1.615000 ;
      RECT 1604.290000  1.835000 1605.870000 2.005000 ;
      RECT 1604.290000  2.005000 1604.630000 2.465000 ;
      RECT 1604.395000  0.515000 1604.725000 0.935000 ;
      RECT 1604.555000  0.935000 1604.725000 1.835000 ;
      RECT 1604.850000  2.175000 1605.195000 2.635000 ;
      RECT 1604.945000  0.085000 1605.195000 0.905000 ;
      RECT 1604.945000  1.105000 1605.450000 1.665000 ;
      RECT 1605.620000  1.355000 1605.870000 1.835000 ;
      RECT 1605.800000  0.255000 1606.420000 0.565000 ;
      RECT 1605.800000  0.565000 1606.210000 1.185000 ;
      RECT 1605.960000  2.150000 1606.290000 2.465000 ;
      RECT 1606.040000  1.185000 1606.210000 1.865000 ;
      RECT 1606.040000  1.865000 1606.290000 2.150000 ;
      RECT 1606.380000  1.125000 1606.615000 1.720000 ;
      RECT 1606.400000  0.735000 1606.955000 0.955000 ;
      RECT 1606.500000  2.175000 1607.690000 2.375000 ;
      RECT 1606.640000  0.255000 1607.365000 0.565000 ;
      RECT 1606.785000  0.955000 1606.955000 1.655000 ;
      RECT 1606.785000  1.655000 1607.300000 2.005000 ;
      RECT 1607.195000  0.565000 1607.365000 1.315000 ;
      RECT 1607.195000  1.315000 1608.095000 1.485000 ;
      RECT 1607.470000  1.485000 1608.095000 1.575000 ;
      RECT 1607.470000  1.575000 1607.690000 2.175000 ;
      RECT 1607.555000  0.765000 1608.720000 1.045000 ;
      RECT 1607.555000  1.045000 1609.230000 1.065000 ;
      RECT 1607.555000  1.065000 1607.805000 1.095000 ;
      RECT 1607.680000  0.085000 1608.075000 0.560000 ;
      RECT 1607.860000  1.835000 1608.095000 2.635000 ;
      RECT 1607.925000  1.245000 1608.095000 1.315000 ;
      RECT 1608.265000  0.255000 1608.720000 0.765000 ;
      RECT 1608.265000  1.065000 1609.230000 1.375000 ;
      RECT 1608.265000  1.375000 1608.645000 2.465000 ;
      RECT 1608.855000  2.105000 1609.145000 2.635000 ;
      RECT 1608.950000  0.085000 1609.225000 0.615000 ;
      RECT 1609.625000  1.245000 1609.865000 1.965000 ;
      RECT 1609.760000  2.165000 1610.875000 2.355000 ;
      RECT 1609.875000  0.705000 1610.405000 1.035000 ;
      RECT 1609.910000  0.330000 1610.875000 0.535000 ;
      RECT 1610.035000  1.035000 1610.405000 1.995000 ;
      RECT 1610.625000  0.535000 1610.875000 2.165000 ;
      RECT 1611.045000  0.085000 1611.290000 0.900000 ;
      RECT 1611.095000  1.495000 1611.265000 2.635000 ;
      RECT 1611.460000  0.255000 1611.815000 2.465000 ;
      RECT 1611.985000  0.890000 1612.445000 1.220000 ;
      RECT 1612.105000  0.255000 1612.445000 0.890000 ;
      RECT 1612.105000  1.220000 1612.445000 2.465000 ;
      RECT 1612.615000  1.070000 1612.945000 1.295000 ;
      RECT 1612.665000  0.085000 1612.900000 0.900000 ;
      RECT 1612.665000  1.465000 1612.900000 2.635000 ;
      RECT 1613.155000  0.255000 1613.570000 2.420000 ;
      RECT 1613.765000  0.085000 1614.055000 0.810000 ;
      RECT 1613.765000  1.470000 1614.055000 2.635000 ;
      RECT 1614.235000  0.975000 1614.585000 1.625000 ;
      RECT 1614.315000  0.345000 1614.485000 0.635000 ;
      RECT 1614.315000  0.635000 1615.035000 0.805000 ;
      RECT 1614.315000  1.795000 1615.035000 1.965000 ;
      RECT 1614.315000  1.965000 1614.485000 2.465000 ;
      RECT 1614.655000  0.085000 1615.035000 0.465000 ;
      RECT 1614.655000  2.135000 1615.035000 2.635000 ;
      RECT 1614.805000  0.805000 1615.035000 1.795000 ;
      RECT 1615.255000  0.345000 1615.425000 2.465000 ;
      RECT 1615.595000  0.255000 1616.025000 0.515000 ;
      RECT 1615.595000  0.515000 1615.765000 1.890000 ;
      RECT 1615.595000  1.890000 1616.025000 2.465000 ;
      RECT 1615.935000  0.765000 1616.295000 1.720000 ;
      RECT 1616.465000  0.765000 1616.905000 1.185000 ;
      RECT 1616.465000  1.185000 1616.665000 1.370000 ;
      RECT 1616.525000  0.085000 1616.905000 0.515000 ;
      RECT 1616.525000  1.890000 1616.905000 2.635000 ;
      RECT 1616.835000  1.355000 1617.425000 1.720000 ;
      RECT 1617.095000  1.720000 1617.425000 2.425000 ;
      RECT 1617.120000  0.255000 1617.345000 0.845000 ;
      RECT 1617.120000  0.845000 1618.025000 1.175000 ;
      RECT 1617.120000  1.175000 1617.425000 1.355000 ;
      RECT 1617.525000  0.085000 1617.905000 0.610000 ;
      RECT 1617.655000  1.825000 1617.850000 2.635000 ;
      RECT 1618.245000  0.685000 1618.415000 1.320000 ;
      RECT 1618.245000  1.320000 1618.665000 1.650000 ;
      RECT 1618.565000  1.820000 1619.005000 2.020000 ;
      RECT 1618.565000  2.020000 1618.945000 2.465000 ;
      RECT 1618.585000  0.255000 1618.905000 0.980000 ;
      RECT 1618.585000  0.980000 1619.005000 1.150000 ;
      RECT 1618.835000  1.150000 1619.005000 1.820000 ;
      RECT 1619.135000  0.255000 1619.335000 0.645000 ;
      RECT 1619.135000  0.645000 1619.395000 0.825000 ;
      RECT 1619.175000  2.210000 1619.505000 2.465000 ;
      RECT 1619.225000  0.825000 1619.395000 1.785000 ;
      RECT 1619.225000  1.785000 1619.505000 2.210000 ;
      RECT 1619.505000  0.255000 1620.365000 0.515000 ;
      RECT 1619.745000  1.105000 1620.025000 1.615000 ;
      RECT 1619.930000  1.835000 1621.510000 2.005000 ;
      RECT 1619.930000  2.005000 1620.270000 2.465000 ;
      RECT 1620.035000  0.515000 1620.365000 0.935000 ;
      RECT 1620.195000  0.935000 1620.365000 1.835000 ;
      RECT 1620.490000  2.175000 1620.835000 2.635000 ;
      RECT 1620.585000  0.085000 1620.835000 0.905000 ;
      RECT 1620.585000  1.105000 1621.090000 1.665000 ;
      RECT 1621.260000  1.355000 1621.510000 1.835000 ;
      RECT 1621.440000  0.255000 1622.060000 0.565000 ;
      RECT 1621.440000  0.565000 1621.850000 1.185000 ;
      RECT 1621.600000  2.150000 1621.930000 2.465000 ;
      RECT 1621.680000  1.185000 1621.850000 1.865000 ;
      RECT 1621.680000  1.865000 1621.930000 2.150000 ;
      RECT 1622.020000  1.125000 1622.255000 1.720000 ;
      RECT 1622.040000  0.735000 1622.595000 0.955000 ;
      RECT 1622.140000  2.175000 1623.330000 2.375000 ;
      RECT 1622.280000  0.255000 1623.005000 0.565000 ;
      RECT 1622.425000  0.955000 1622.595000 1.655000 ;
      RECT 1622.425000  1.655000 1622.940000 2.005000 ;
      RECT 1622.835000  0.565000 1623.005000 1.315000 ;
      RECT 1622.835000  1.315000 1623.735000 1.485000 ;
      RECT 1623.110000  1.485000 1623.735000 1.575000 ;
      RECT 1623.110000  1.575000 1623.330000 2.175000 ;
      RECT 1623.195000  0.765000 1624.360000 1.045000 ;
      RECT 1623.195000  1.045000 1624.870000 1.065000 ;
      RECT 1623.195000  1.065000 1623.445000 1.095000 ;
      RECT 1623.320000  0.085000 1623.715000 0.560000 ;
      RECT 1623.500000  1.835000 1623.735000 2.635000 ;
      RECT 1623.565000  1.245000 1623.735000 1.315000 ;
      RECT 1623.905000  0.255000 1624.360000 0.765000 ;
      RECT 1623.905000  1.065000 1624.870000 1.375000 ;
      RECT 1623.905000  1.375000 1624.285000 2.465000 ;
      RECT 1624.495000  2.105000 1624.785000 2.635000 ;
      RECT 1624.590000  0.085000 1624.865000 0.615000 ;
      RECT 1625.265000  1.245000 1625.505000 1.965000 ;
      RECT 1625.400000  2.165000 1626.515000 2.355000 ;
      RECT 1625.530000  0.705000 1626.045000 1.035000 ;
      RECT 1625.550000  0.330000 1626.515000 0.535000 ;
      RECT 1625.675000  1.035000 1626.045000 1.995000 ;
      RECT 1626.265000  0.535000 1626.515000 2.165000 ;
      RECT 1626.735000  1.495000 1626.905000 2.635000 ;
      RECT 1626.770000  0.085000 1627.020000 0.900000 ;
      RECT 1627.075000  1.065000 1627.570000 1.300000 ;
      RECT 1627.075000  1.300000 1627.455000 2.465000 ;
      RECT 1627.240000  0.255000 1627.570000 1.065000 ;
      RECT 1627.675000  1.465000 1627.925000 2.635000 ;
      RECT 1627.790000  0.085000 1628.040000 0.900000 ;
      RECT 1628.095000  1.575000 1628.325000 2.010000 ;
      RECT 1628.210000  0.890000 1628.835000 1.220000 ;
      RECT 1628.495000  0.255000 1628.835000 0.890000 ;
      RECT 1628.495000  1.220000 1628.835000 2.465000 ;
      RECT 1629.055000  0.085000 1629.290000 0.900000 ;
      RECT 1629.055000  1.465000 1629.290000 2.635000 ;
      RECT 1629.460000  0.255000 1629.840000 2.420000 ;
      RECT 1630.060000  0.085000 1630.320000 0.900000 ;
      RECT 1630.060000  1.465000 1630.320000 2.635000 ;
      RECT 1630.785000  0.085000 1631.075000 0.810000 ;
      RECT 1630.785000  1.470000 1631.075000 2.635000 ;
      RECT 1631.245000  0.280000 1631.710000 0.825000 ;
      RECT 1631.245000  0.825000 1631.415000 1.785000 ;
      RECT 1631.245000  1.785000 1633.715000 1.955000 ;
      RECT 1631.245000  2.125000 1631.545000 2.635000 ;
      RECT 1631.585000  0.995000 1631.970000 1.445000 ;
      RECT 1631.585000  1.445000 1633.325000 1.615000 ;
      RECT 1631.715000  1.955000 1632.095000 2.465000 ;
      RECT 1632.140000  1.075000 1632.935000 1.275000 ;
      RECT 1632.315000  0.085000 1632.485000 0.905000 ;
      RECT 1632.315000  2.125000 1632.995000 2.635000 ;
      RECT 1632.655000  0.255000 1633.035000 0.655000 ;
      RECT 1632.655000  0.655000 1634.055000 0.825000 ;
      RECT 1633.105000  1.075000 1633.805000 1.245000 ;
      RECT 1633.105000  1.245000 1633.325000 1.445000 ;
      RECT 1633.255000  0.085000 1633.655000 0.475000 ;
      RECT 1633.495000  1.415000 1634.255000 1.585000 ;
      RECT 1633.495000  1.585000 1633.715000 1.785000 ;
      RECT 1633.675000  2.125000 1634.055000 2.295000 ;
      RECT 1633.825000  0.255000 1634.055000 0.655000 ;
      RECT 1633.885000  1.755000 1634.755000 1.955000 ;
      RECT 1633.885000  1.955000 1634.055000 2.125000 ;
      RECT 1634.035000  0.995000 1634.255000 1.415000 ;
      RECT 1634.275000  2.125000 1634.575000 2.635000 ;
      RECT 1634.335000  0.345000 1634.755000 0.825000 ;
      RECT 1634.515000  0.825000 1634.755000 1.755000 ;
      RECT 1634.925000  0.085000 1635.215000 0.810000 ;
      RECT 1634.925000  1.470000 1635.215000 2.635000 ;
      RECT 1635.385000  0.645000 1636.210000 0.895000 ;
      RECT 1635.385000  0.895000 1635.615000 1.785000 ;
      RECT 1635.385000  1.785000 1639.080000 1.955000 ;
      RECT 1635.385000  1.955000 1637.580000 1.965000 ;
      RECT 1635.385000  1.965000 1635.700000 2.465000 ;
      RECT 1635.405000  0.255000 1636.680000 0.475000 ;
      RECT 1635.785000  1.075000 1636.310000 1.285000 ;
      RECT 1635.920000  2.135000 1636.170000 2.635000 ;
      RECT 1636.140000  1.285000 1636.310000 1.445000 ;
      RECT 1636.140000  1.445000 1638.650000 1.615000 ;
      RECT 1636.390000  1.965000 1636.640000 2.465000 ;
      RECT 1636.430000  0.475000 1636.680000 0.725000 ;
      RECT 1636.430000  0.725000 1637.620000 0.905000 ;
      RECT 1636.655000  1.075000 1638.205000 1.275000 ;
      RECT 1636.860000  2.135000 1637.110000 2.635000 ;
      RECT 1636.900000  0.085000 1637.070000 0.555000 ;
      RECT 1637.240000  0.255000 1637.620000 0.725000 ;
      RECT 1637.330000  1.965000 1637.580000 2.465000 ;
      RECT 1637.890000  2.125000 1638.140000 2.465000 ;
      RECT 1637.930000  0.085000 1638.100000 0.905000 ;
      RECT 1638.270000  0.255000 1638.650000 0.725000 ;
      RECT 1638.270000  0.725000 1641.055000 0.905000 ;
      RECT 1638.360000  2.135000 1638.610000 2.635000 ;
      RECT 1638.480000  1.075000 1639.605000 1.285000 ;
      RECT 1638.480000  1.285000 1638.650000 1.445000 ;
      RECT 1638.830000  2.125000 1639.155000 2.295000 ;
      RECT 1638.830000  2.295000 1640.055000 2.465000 ;
      RECT 1638.870000  0.085000 1639.040000 0.555000 ;
      RECT 1638.910000  1.455000 1640.505000 1.625000 ;
      RECT 1638.910000  1.625000 1639.080000 1.785000 ;
      RECT 1639.210000  0.255000 1639.625000 0.725000 ;
      RECT 1639.375000  1.795000 1641.045000 1.965000 ;
      RECT 1639.375000  1.965000 1639.585000 2.125000 ;
      RECT 1639.805000  2.135000 1640.055000 2.295000 ;
      RECT 1639.845000  0.085000 1640.015000 0.555000 ;
      RECT 1640.285000  0.305000 1641.640000 0.475000 ;
      RECT 1640.325000  2.135000 1640.575000 2.635000 ;
      RECT 1640.335000  1.075000 1641.045000 1.245000 ;
      RECT 1640.335000  1.245000 1640.505000 1.455000 ;
      RECT 1640.705000  0.645000 1641.055000 0.725000 ;
      RECT 1640.795000  1.415000 1641.640000 1.625000 ;
      RECT 1640.795000  1.625000 1641.045000 1.795000 ;
      RECT 1640.795000  1.965000 1641.045000 2.125000 ;
      RECT 1641.250000  0.475000 1641.640000 1.415000 ;
      RECT 1641.265000  1.795000 1641.640000 2.635000 ;
      RECT 1641.825000  0.085000 1642.115000 0.810000 ;
      RECT 1641.825000  1.470000 1642.115000 2.635000 ;
      RECT 1642.285000  0.645000 1644.110000 0.905000 ;
      RECT 1642.285000  0.905000 1642.520000 1.445000 ;
      RECT 1642.285000  1.445000 1643.600000 1.615000 ;
      RECT 1642.285000  1.615000 1642.660000 2.465000 ;
      RECT 1642.370000  0.255000 1644.580000 0.475000 ;
      RECT 1642.690000  1.075000 1644.205000 1.275000 ;
      RECT 1642.880000  1.835000 1643.130000 2.635000 ;
      RECT 1643.350000  1.615000 1643.600000 1.785000 ;
      RECT 1643.350000  1.785000 1646.420000 2.005000 ;
      RECT 1643.350000  2.005000 1643.600000 2.465000 ;
      RECT 1643.820000  2.175000 1644.070000 2.635000 ;
      RECT 1644.035000  1.275000 1644.205000 1.445000 ;
      RECT 1644.035000  1.445000 1648.470000 1.615000 ;
      RECT 1644.290000  2.005000 1644.540000 2.465000 ;
      RECT 1644.330000  0.475000 1644.580000 0.725000 ;
      RECT 1644.330000  0.725000 1646.460000 0.905000 ;
      RECT 1644.575000  1.075000 1648.130000 1.275000 ;
      RECT 1644.760000  2.175000 1645.010000 2.635000 ;
      RECT 1644.800000  0.085000 1644.970000 0.555000 ;
      RECT 1645.140000  0.255000 1645.520000 0.725000 ;
      RECT 1645.230000  2.005000 1645.480000 2.465000 ;
      RECT 1645.700000  2.175000 1645.950000 2.635000 ;
      RECT 1645.740000  0.085000 1645.910000 0.555000 ;
      RECT 1646.080000  0.255000 1646.460000 0.725000 ;
      RECT 1646.170000  2.005000 1646.420000 2.465000 ;
      RECT 1646.625000  1.785000 1648.780000 2.005000 ;
      RECT 1646.625000  2.005000 1646.940000 2.465000 ;
      RECT 1646.630000  0.085000 1646.900000 0.905000 ;
      RECT 1647.070000  0.255000 1647.450000 0.725000 ;
      RECT 1647.070000  0.725000 1650.370000 0.735000 ;
      RECT 1647.070000  0.735000 1651.180000 0.905000 ;
      RECT 1647.160000  2.175000 1647.410000 2.635000 ;
      RECT 1647.630000  2.005000 1647.880000 2.465000 ;
      RECT 1647.670000  0.085000 1647.840000 0.555000 ;
      RECT 1648.010000  0.255000 1648.390000 0.725000 ;
      RECT 1648.100000  2.175000 1648.350000 2.635000 ;
      RECT 1648.300000  1.075000 1650.370000 1.275000 ;
      RECT 1648.300000  1.275000 1648.470000 1.445000 ;
      RECT 1648.570000  2.005000 1648.780000 2.215000 ;
      RECT 1648.570000  2.215000 1650.740000 2.465000 ;
      RECT 1648.610000  0.085000 1648.780000 0.555000 ;
      RECT 1648.690000  1.445000 1650.760000 1.615000 ;
      RECT 1648.950000  0.255000 1649.330000 0.725000 ;
      RECT 1648.950000  1.785000 1651.260000 2.045000 ;
      RECT 1649.550000  0.085000 1649.720000 0.555000 ;
      RECT 1649.890000  0.255000 1650.270000 0.725000 ;
      RECT 1650.490000  0.085000 1650.660000 0.555000 ;
      RECT 1650.590000  1.075000 1652.735000 1.275000 ;
      RECT 1650.590000  1.275000 1650.760000 1.445000 ;
      RECT 1650.930000  0.305000 1653.140000 0.475000 ;
      RECT 1650.930000  0.475000 1651.180000 0.735000 ;
      RECT 1650.930000  1.445000 1653.140000 1.665000 ;
      RECT 1650.930000  1.665000 1651.260000 1.785000 ;
      RECT 1650.930000  2.045000 1651.260000 2.465000 ;
      RECT 1651.350000  0.655000 1653.140000 0.905000 ;
      RECT 1651.440000  1.835000 1651.690000 2.635000 ;
      RECT 1651.910000  1.665000 1652.160000 2.465000 ;
      RECT 1652.380000  1.835000 1652.630000 2.635000 ;
      RECT 1652.810000  1.665000 1653.140000 2.465000 ;
      RECT 1652.905000  0.905000 1653.140000 1.445000 ;
      RECT 1653.325000  0.085000 1653.615000 0.810000 ;
      RECT 1653.325000  1.470000 1653.615000 2.635000 ;
      RECT 1653.785000  0.350000 1654.045000 1.440000 ;
      RECT 1653.785000  1.440000 1654.065000 2.465000 ;
      RECT 1654.215000  0.085000 1654.515000 0.525000 ;
      RECT 1654.215000  0.695000 1654.905000 0.865000 ;
      RECT 1654.215000  0.865000 1654.455000 1.330000 ;
      RECT 1654.235000  1.330000 1654.455000 1.875000 ;
      RECT 1654.235000  1.875000 1655.020000 2.045000 ;
      RECT 1654.235000  2.215000 1654.620000 2.635000 ;
      RECT 1654.685000  0.255000 1656.355000 0.425000 ;
      RECT 1654.685000  0.425000 1654.905000 0.695000 ;
      RECT 1654.685000  1.535000 1656.370000 1.705000 ;
      RECT 1654.800000  2.045000 1655.020000 2.235000 ;
      RECT 1654.800000  2.235000 1656.370000 2.405000 ;
      RECT 1655.075000  0.595000 1655.245000 1.535000 ;
      RECT 1655.360000  1.895000 1658.060000 2.065000 ;
      RECT 1655.415000  1.075000 1656.030000 1.325000 ;
      RECT 1655.545000  0.625000 1656.865000 0.795000 ;
      RECT 1655.545000  0.795000 1655.925000 0.905000 ;
      RECT 1655.870000  0.425000 1656.355000 0.455000 ;
      RECT 1656.200000  0.995000 1656.525000 1.325000 ;
      RECT 1656.200000  1.325000 1656.370000 1.535000 ;
      RECT 1656.575000  0.285000 1657.205000 0.455000 ;
      RECT 1656.590000  1.525000 1656.975000 1.695000 ;
      RECT 1656.695000  0.795000 1656.865000 1.375000 ;
      RECT 1656.695000  1.375000 1656.975000 1.525000 ;
      RECT 1657.035000  0.455000 1657.205000 1.035000 ;
      RECT 1657.035000  1.035000 1657.315000 1.205000 ;
      RECT 1657.125000  2.235000 1657.455000 2.635000 ;
      RECT 1657.145000  1.205000 1657.315000 1.895000 ;
      RECT 1657.375000  0.085000 1657.545000 0.865000 ;
      RECT 1657.545000  1.445000 1658.065000 1.715000 ;
      RECT 1657.775000  0.415000 1658.065000 1.445000 ;
      RECT 1657.890000  2.065000 1658.060000 2.275000 ;
      RECT 1657.890000  2.275000 1661.185000 2.445000 ;
      RECT 1658.245000  0.265000 1658.655000 0.485000 ;
      RECT 1658.245000  0.485000 1658.455000 0.595000 ;
      RECT 1658.245000  0.595000 1658.415000 2.105000 ;
      RECT 1658.585000  0.720000 1659.045000 0.825000 ;
      RECT 1658.585000  0.825000 1658.845000 0.890000 ;
      RECT 1658.585000  0.890000 1658.755000 2.275000 ;
      RECT 1658.625000  0.655000 1659.045000 0.720000 ;
      RECT 1658.875000  0.320000 1659.045000 0.655000 ;
      RECT 1658.985000  1.445000 1659.815000 1.615000 ;
      RECT 1658.985000  1.615000 1659.400000 2.045000 ;
      RECT 1659.000000  0.995000 1659.425000 1.270000 ;
      RECT 1659.215000  0.630000 1659.425000 0.995000 ;
      RECT 1659.645000  0.255000 1660.840000 0.425000 ;
      RECT 1659.645000  0.425000 1659.815000 1.445000 ;
      RECT 1659.985000  0.595000 1660.155000 1.935000 ;
      RECT 1659.985000  1.935000 1662.810000 2.105000 ;
      RECT 1660.325000  0.425000 1660.840000 0.465000 ;
      RECT 1660.325000  0.995000 1660.545000 1.445000 ;
      RECT 1660.325000  1.445000 1660.955000 1.615000 ;
      RECT 1660.715000  0.730000 1660.920000 0.945000 ;
      RECT 1660.715000  0.945000 1661.025000 1.275000 ;
      RECT 1661.175000  1.495000 1662.360000 1.705000 ;
      RECT 1661.195000  1.075000 1661.915000 1.325000 ;
      RECT 1661.215000  0.295000 1661.505000 0.735000 ;
      RECT 1661.215000  0.735000 1662.360000 0.750000 ;
      RECT 1661.255000  0.750000 1662.360000 0.905000 ;
      RECT 1661.615000  2.275000 1662.295000 2.635000 ;
      RECT 1661.750000  0.085000 1662.210000 0.565000 ;
      RECT 1662.190000  0.905000 1662.360000 0.995000 ;
      RECT 1662.190000  0.995000 1662.470000 1.325000 ;
      RECT 1662.190000  1.325000 1662.360000 1.495000 ;
      RECT 1662.275000  1.875000 1662.810000 1.935000 ;
      RECT 1662.510000  0.255000 1662.810000 0.585000 ;
      RECT 1662.515000  2.105000 1662.810000 2.465000 ;
      RECT 1662.640000  0.585000 1662.810000 1.875000 ;
      RECT 1662.985000  0.085000 1663.275000 0.810000 ;
      RECT 1662.985000  1.470000 1663.275000 2.635000 ;
      RECT 1663.445000  0.085000 1663.735000 0.735000 ;
      RECT 1663.445000  1.490000 1663.735000 2.635000 ;
      RECT 1663.905000  0.350000 1664.225000 2.465000 ;
      RECT 1664.395000  0.085000 1664.685000 0.525000 ;
      RECT 1664.405000  0.695000 1665.075000 0.865000 ;
      RECT 1664.405000  0.865000 1664.625000 1.875000 ;
      RECT 1664.405000  1.875000 1665.190000 2.045000 ;
      RECT 1664.405000  2.215000 1664.790000 2.635000 ;
      RECT 1664.855000  0.255000 1666.525000 0.425000 ;
      RECT 1664.855000  0.425000 1665.075000 0.695000 ;
      RECT 1664.855000  1.535000 1666.540000 1.705000 ;
      RECT 1664.970000  2.045000 1665.190000 2.235000 ;
      RECT 1664.970000  2.235000 1666.540000 2.405000 ;
      RECT 1665.245000  0.595000 1665.415000 1.535000 ;
      RECT 1665.530000  1.895000 1668.230000 2.065000 ;
      RECT 1665.585000  1.075000 1666.200000 1.325000 ;
      RECT 1665.715000  0.625000 1667.035000 0.795000 ;
      RECT 1665.715000  0.795000 1666.095000 0.905000 ;
      RECT 1666.040000  0.425000 1666.525000 0.455000 ;
      RECT 1666.370000  0.995000 1666.695000 1.325000 ;
      RECT 1666.370000  1.325000 1666.540000 1.535000 ;
      RECT 1666.745000  0.285000 1667.375000 0.455000 ;
      RECT 1666.760000  1.525000 1667.145000 1.695000 ;
      RECT 1666.865000  0.795000 1667.035000 1.375000 ;
      RECT 1666.865000  1.375000 1667.145000 1.525000 ;
      RECT 1667.205000  0.455000 1667.375000 1.035000 ;
      RECT 1667.205000  1.035000 1667.485000 1.205000 ;
      RECT 1667.295000  2.235000 1667.625000 2.635000 ;
      RECT 1667.315000  1.205000 1667.485000 1.895000 ;
      RECT 1667.545000  0.085000 1667.715000 0.865000 ;
      RECT 1667.715000  1.445000 1668.235000 1.715000 ;
      RECT 1667.945000  0.415000 1668.235000 1.445000 ;
      RECT 1668.060000  2.065000 1668.230000 2.275000 ;
      RECT 1668.060000  2.275000 1671.355000 2.445000 ;
      RECT 1668.415000  0.265000 1668.825000 0.485000 ;
      RECT 1668.415000  0.485000 1668.625000 0.595000 ;
      RECT 1668.415000  0.595000 1668.585000 2.105000 ;
      RECT 1668.755000  0.720000 1669.215000 0.825000 ;
      RECT 1668.755000  0.825000 1669.015000 0.890000 ;
      RECT 1668.755000  0.890000 1668.925000 2.275000 ;
      RECT 1668.795000  0.655000 1669.215000 0.720000 ;
      RECT 1669.045000  0.320000 1669.215000 0.655000 ;
      RECT 1669.155000  1.445000 1669.985000 1.615000 ;
      RECT 1669.155000  1.615000 1669.570000 2.045000 ;
      RECT 1669.170000  0.995000 1669.595000 1.270000 ;
      RECT 1669.385000  0.630000 1669.595000 0.995000 ;
      RECT 1669.815000  0.255000 1671.010000 0.425000 ;
      RECT 1669.815000  0.425000 1669.985000 1.445000 ;
      RECT 1670.155000  0.595000 1670.325000 1.935000 ;
      RECT 1670.155000  1.935000 1672.845000 2.105000 ;
      RECT 1670.495000  0.425000 1671.010000 0.465000 ;
      RECT 1670.495000  0.995000 1670.715000 1.445000 ;
      RECT 1670.495000  1.445000 1671.125000 1.615000 ;
      RECT 1670.885000  0.730000 1671.090000 0.945000 ;
      RECT 1670.885000  0.945000 1671.195000 1.275000 ;
      RECT 1671.345000  1.495000 1672.395000 1.705000 ;
      RECT 1671.385000  0.295000 1671.675000 0.735000 ;
      RECT 1671.385000  0.735000 1672.395000 0.750000 ;
      RECT 1671.415000  1.075000 1672.055000 1.325000 ;
      RECT 1671.425000  0.750000 1672.395000 0.905000 ;
      RECT 1671.815000  2.275000 1672.150000 2.635000 ;
      RECT 1671.895000  0.085000 1672.065000 0.565000 ;
      RECT 1672.225000  0.905000 1672.395000 0.995000 ;
      RECT 1672.225000  0.995000 1672.505000 1.325000 ;
      RECT 1672.225000  1.325000 1672.395000 1.495000 ;
      RECT 1672.310000  1.875000 1672.845000 1.935000 ;
      RECT 1672.545000  0.255000 1672.845000 0.585000 ;
      RECT 1672.550000  2.105000 1672.845000 2.465000 ;
      RECT 1672.675000  0.585000 1672.845000 1.875000 ;
      RECT 1673.105000  0.085000 1673.395000 0.810000 ;
      RECT 1673.105000  1.470000 1673.395000 2.635000 ;
      RECT 1673.765000  0.085000 1673.935000 0.735000 ;
      RECT 1673.765000  1.490000 1673.935000 2.635000 ;
      RECT 1674.105000  0.375000 1674.405000 0.995000 ;
      RECT 1674.105000  0.995000 1675.340000 1.325000 ;
      RECT 1674.105000  1.325000 1674.485000 2.425000 ;
      RECT 1674.705000  0.085000 1674.875000 0.735000 ;
      RECT 1674.705000  1.495000 1674.875000 2.635000 ;
      RECT 1675.045000  0.350000 1675.355000 0.925000 ;
      RECT 1675.045000  0.925000 1675.340000 0.995000 ;
      RECT 1675.045000  1.325000 1675.340000 1.440000 ;
      RECT 1675.045000  1.440000 1675.375000 2.465000 ;
      RECT 1675.510000  0.995000 1675.765000 1.325000 ;
      RECT 1675.525000  0.085000 1675.825000 0.525000 ;
      RECT 1675.540000  0.695000 1676.215000 0.865000 ;
      RECT 1675.540000  0.865000 1675.765000 0.995000 ;
      RECT 1675.545000  1.325000 1675.765000 1.875000 ;
      RECT 1675.545000  1.875000 1676.330000 2.045000 ;
      RECT 1675.545000  2.215000 1675.930000 2.635000 ;
      RECT 1675.995000  0.255000 1677.665000 0.425000 ;
      RECT 1675.995000  0.425000 1676.215000 0.695000 ;
      RECT 1675.995000  1.535000 1677.680000 1.705000 ;
      RECT 1676.110000  2.045000 1676.330000 2.235000 ;
      RECT 1676.110000  2.235000 1677.680000 2.405000 ;
      RECT 1676.385000  0.595000 1676.555000 1.535000 ;
      RECT 1676.670000  1.895000 1679.370000 2.065000 ;
      RECT 1676.725000  1.075000 1677.340000 1.325000 ;
      RECT 1676.855000  0.625000 1678.175000 0.795000 ;
      RECT 1676.855000  0.795000 1677.235000 0.905000 ;
      RECT 1677.180000  0.425000 1677.665000 0.455000 ;
      RECT 1677.510000  0.995000 1677.835000 1.325000 ;
      RECT 1677.510000  1.325000 1677.680000 1.535000 ;
      RECT 1677.885000  0.285000 1678.515000 0.455000 ;
      RECT 1677.900000  1.525000 1678.285000 1.695000 ;
      RECT 1678.005000  0.795000 1678.175000 1.375000 ;
      RECT 1678.005000  1.375000 1678.285000 1.525000 ;
      RECT 1678.345000  0.455000 1678.515000 1.035000 ;
      RECT 1678.345000  1.035000 1678.625000 1.205000 ;
      RECT 1678.435000  2.235000 1678.765000 2.635000 ;
      RECT 1678.455000  1.205000 1678.625000 1.895000 ;
      RECT 1678.685000  0.085000 1678.855000 0.865000 ;
      RECT 1678.855000  1.445000 1679.375000 1.715000 ;
      RECT 1679.085000  0.415000 1679.375000 1.445000 ;
      RECT 1679.200000  2.065000 1679.370000 2.275000 ;
      RECT 1679.200000  2.275000 1682.495000 2.445000 ;
      RECT 1679.555000  0.265000 1680.000000 0.485000 ;
      RECT 1679.555000  0.485000 1679.725000 2.105000 ;
      RECT 1679.895000  0.655000 1680.355000 0.825000 ;
      RECT 1679.895000  0.825000 1680.065000 2.275000 ;
      RECT 1680.185000  0.320000 1680.355000 0.655000 ;
      RECT 1680.295000  1.445000 1681.125000 1.615000 ;
      RECT 1680.295000  1.615000 1680.710000 2.045000 ;
      RECT 1680.310000  0.995000 1680.735000 1.270000 ;
      RECT 1680.525000  0.630000 1680.735000 0.995000 ;
      RECT 1680.955000  0.255000 1682.150000 0.425000 ;
      RECT 1680.955000  0.425000 1681.125000 1.445000 ;
      RECT 1681.295000  0.595000 1681.465000 1.935000 ;
      RECT 1681.295000  1.935000 1683.805000 2.105000 ;
      RECT 1681.635000  0.425000 1682.150000 0.465000 ;
      RECT 1681.635000  0.995000 1681.855000 1.445000 ;
      RECT 1681.635000  1.445000 1682.265000 1.615000 ;
      RECT 1682.025000  0.730000 1682.230000 0.945000 ;
      RECT 1682.025000  0.945000 1682.335000 1.275000 ;
      RECT 1682.485000  1.495000 1683.355000 1.705000 ;
      RECT 1682.525000  0.295000 1682.815000 0.735000 ;
      RECT 1682.525000  0.735000 1683.355000 0.750000 ;
      RECT 1682.555000  1.075000 1683.015000 1.325000 ;
      RECT 1682.565000  0.750000 1683.355000 0.905000 ;
      RECT 1682.905000  2.275000 1683.290000 2.635000 ;
      RECT 1683.035000  0.085000 1683.205000 0.565000 ;
      RECT 1683.185000  0.905000 1683.355000 0.995000 ;
      RECT 1683.185000  0.995000 1683.465000 1.325000 ;
      RECT 1683.185000  1.325000 1683.355000 1.495000 ;
      RECT 1683.270000  1.875000 1683.805000 1.935000 ;
      RECT 1683.505000  0.255000 1683.805000 0.585000 ;
      RECT 1683.510000  2.105000 1683.805000 2.465000 ;
      RECT 1683.635000  0.585000 1683.805000 1.875000 ;
      RECT 1684.145000  0.085000 1684.435000 0.810000 ;
      RECT 1684.145000  1.470000 1684.435000 2.635000 ;
      RECT 1684.605000  0.655000 1687.265000 0.825000 ;
      RECT 1684.605000  0.825000 1684.775000 1.785000 ;
      RECT 1684.605000  1.785000 1684.985000 2.465000 ;
      RECT 1684.655000  0.085000 1684.985000 0.475000 ;
      RECT 1684.945000  0.995000 1685.295000 1.445000 ;
      RECT 1684.945000  1.445000 1686.410000 1.615000 ;
      RECT 1685.205000  0.335000 1685.375000 0.655000 ;
      RECT 1685.475000  1.075000 1686.020000 1.275000 ;
      RECT 1685.555000  0.085000 1685.935000 0.475000 ;
      RECT 1685.685000  1.785000 1685.855000 2.635000 ;
      RECT 1686.025000  1.785000 1687.375000 1.955000 ;
      RECT 1686.025000  1.955000 1686.405000 2.465000 ;
      RECT 1686.240000  1.075000 1686.675000 1.245000 ;
      RECT 1686.240000  1.245000 1686.410000 1.445000 ;
      RECT 1686.400000  0.315000 1687.605000 0.485000 ;
      RECT 1686.635000  2.125000 1686.805000 2.635000 ;
      RECT 1686.975000  1.955000 1687.375000 2.465000 ;
      RECT 1687.035000  0.825000 1687.265000 1.325000 ;
      RECT 1687.435000  0.485000 1687.605000 1.365000 ;
      RECT 1687.435000  1.365000 1688.065000 1.535000 ;
      RECT 1687.745000  1.535000 1688.065000 2.465000 ;
      RECT 1687.775000  0.085000 1688.065000 0.920000 ;
      RECT 1688.285000  0.085000 1688.575000 0.810000 ;
      RECT 1688.285000  1.470000 1688.575000 2.635000 ;
      RECT 1688.780000  0.725000 1690.510000 0.905000 ;
      RECT 1688.780000  0.905000 1688.950000 1.785000 ;
      RECT 1688.780000  1.785000 1691.080000 1.955000 ;
      RECT 1688.780000  2.135000 1689.060000 2.465000 ;
      RECT 1688.805000  2.125000 1688.975000 2.135000 ;
      RECT 1688.850000  0.085000 1689.020000 0.555000 ;
      RECT 1689.190000  0.255000 1689.570000 0.725000 ;
      RECT 1689.205000  1.075000 1689.585000 1.275000 ;
      RECT 1689.280000  2.135000 1689.530000 2.635000 ;
      RECT 1689.415000  1.275000 1689.585000 1.445000 ;
      RECT 1689.415000  1.445000 1690.740000 1.615000 ;
      RECT 1689.750000  2.135000 1690.000000 2.295000 ;
      RECT 1689.750000  2.295000 1690.940000 2.465000 ;
      RECT 1689.790000  0.085000 1689.960000 0.555000 ;
      RECT 1689.805000  1.075000 1690.350000 1.275000 ;
      RECT 1689.825000  2.125000 1689.995000 2.135000 ;
      RECT 1690.130000  0.255000 1690.510000 0.725000 ;
      RECT 1690.220000  1.955000 1690.470000 2.125000 ;
      RECT 1690.520000  1.075000 1692.190000 1.275000 ;
      RECT 1690.520000  1.275000 1690.740000 1.445000 ;
      RECT 1690.690000  2.135000 1690.940000 2.295000 ;
      RECT 1690.730000  0.085000 1690.900000 0.555000 ;
      RECT 1690.910000  1.445000 1693.845000 1.615000 ;
      RECT 1690.910000  1.615000 1691.080000 1.785000 ;
      RECT 1691.145000  2.125000 1691.460000 2.465000 ;
      RECT 1691.170000  0.255000 1691.500000 0.725000 ;
      RECT 1691.170000  0.725000 1692.360000 0.905000 ;
      RECT 1691.250000  1.785000 1693.915000 1.955000 ;
      RECT 1691.250000  1.955000 1691.460000 2.125000 ;
      RECT 1691.680000  2.135000 1691.930000 2.635000 ;
      RECT 1691.720000  0.085000 1691.890000 0.555000 ;
      RECT 1692.060000  0.255000 1693.440000 0.475000 ;
      RECT 1692.060000  0.475000 1692.360000 0.725000 ;
      RECT 1692.150000  1.955000 1692.400000 2.465000 ;
      RECT 1692.380000  1.075000 1693.150000 1.275000 ;
      RECT 1692.620000  2.135000 1692.925000 2.635000 ;
      RECT 1692.635000  0.645000 1692.965000 0.725000 ;
      RECT 1692.635000  0.725000 1695.010000 0.905000 ;
      RECT 1693.145000  1.955000 1693.915000 2.295000 ;
      RECT 1693.145000  2.295000 1694.855000 2.465000 ;
      RECT 1693.675000  1.075000 1694.385000 1.245000 ;
      RECT 1693.675000  1.245000 1693.845000 1.445000 ;
      RECT 1693.705000  0.085000 1693.875000 0.555000 ;
      RECT 1694.045000  0.645000 1694.425000 0.725000 ;
      RECT 1694.135000  1.415000 1695.010000 1.625000 ;
      RECT 1694.135000  1.625000 1694.385000 2.125000 ;
      RECT 1694.605000  1.795000 1694.855000 2.295000 ;
      RECT 1694.645000  0.085000 1694.815000 0.555000 ;
      RECT 1694.645000  0.905000 1695.010000 1.415000 ;
      RECT 1695.185000  0.085000 1695.475000 0.810000 ;
      RECT 1695.185000  1.470000 1695.475000 2.635000 ;
      RECT 1695.645000  0.085000 1695.920000 0.565000 ;
      RECT 1695.645000  0.735000 1699.290000 0.905000 ;
      RECT 1695.645000  0.905000 1695.815000 1.445000 ;
      RECT 1695.645000  1.445000 1698.230000 1.615000 ;
      RECT 1695.645000  1.785000 1697.840000 2.005000 ;
      RECT 1695.645000  2.005000 1695.960000 2.465000 ;
      RECT 1695.985000  1.075000 1698.660000 1.275000 ;
      RECT 1696.090000  0.255000 1696.470000 0.725000 ;
      RECT 1696.090000  0.725000 1699.290000 0.735000 ;
      RECT 1696.180000  2.175000 1696.430000 2.635000 ;
      RECT 1696.650000  2.005000 1696.900000 2.465000 ;
      RECT 1696.690000  0.085000 1696.860000 0.555000 ;
      RECT 1697.030000  0.255000 1697.410000 0.725000 ;
      RECT 1697.120000  2.175000 1697.370000 2.635000 ;
      RECT 1697.590000  2.005000 1697.840000 2.295000 ;
      RECT 1697.590000  2.295000 1699.720000 2.465000 ;
      RECT 1697.630000  0.085000 1697.800000 0.555000 ;
      RECT 1697.970000  0.255000 1698.350000 0.725000 ;
      RECT 1698.060000  1.615000 1698.230000 1.785000 ;
      RECT 1698.060000  1.785000 1699.250000 1.955000 ;
      RECT 1698.060000  1.955000 1698.310000 2.125000 ;
      RECT 1698.440000  1.275000 1698.660000 1.445000 ;
      RECT 1698.440000  1.445000 1702.375000 1.615000 ;
      RECT 1698.530000  2.125000 1698.780000 2.295000 ;
      RECT 1698.570000  0.085000 1698.740000 0.555000 ;
      RECT 1698.830000  1.075000 1701.060000 1.105000 ;
      RECT 1698.830000  1.105000 1701.900000 1.275000 ;
      RECT 1698.910000  0.255000 1699.290000 0.725000 ;
      RECT 1699.000000  1.955000 1699.250000 2.125000 ;
      RECT 1699.470000  1.795000 1699.720000 2.295000 ;
      RECT 1699.510000  0.085000 1699.780000 0.895000 ;
      RECT 1699.950000  0.255000 1702.160000 0.475000 ;
      RECT 1699.990000  1.785000 1704.000000 2.005000 ;
      RECT 1699.990000  2.005000 1700.240000 2.465000 ;
      RECT 1700.125000  0.645000 1701.690000 0.905000 ;
      RECT 1700.460000  2.175000 1700.710000 2.635000 ;
      RECT 1700.930000  2.005000 1701.180000 2.465000 ;
      RECT 1701.210000  0.905000 1701.690000 0.935000 ;
      RECT 1701.400000  2.175000 1701.650000 2.635000 ;
      RECT 1701.870000  2.005000 1702.120000 2.465000 ;
      RECT 1701.910000  0.475000 1702.160000 0.725000 ;
      RECT 1701.910000  0.725000 1704.040000 0.905000 ;
      RECT 1702.155000  1.075000 1703.680000 1.275000 ;
      RECT 1702.155000  1.275000 1702.375000 1.445000 ;
      RECT 1702.340000  2.175000 1702.590000 2.635000 ;
      RECT 1702.380000  0.085000 1702.550000 0.555000 ;
      RECT 1702.720000  0.255000 1703.100000 0.725000 ;
      RECT 1702.810000  1.455000 1703.060000 1.785000 ;
      RECT 1702.810000  2.005000 1703.060000 2.465000 ;
      RECT 1703.280000  2.175000 1703.530000 2.635000 ;
      RECT 1703.320000  0.085000 1703.490000 0.555000 ;
      RECT 1703.570000  1.445000 1704.070000 1.615000 ;
      RECT 1703.660000  0.255000 1704.040000 0.725000 ;
      RECT 1703.750000  2.005000 1704.000000 2.295000 ;
      RECT 1703.750000  2.295000 1705.940000 2.465000 ;
      RECT 1703.900000  1.075000 1705.690000 1.275000 ;
      RECT 1703.900000  1.275000 1704.070000 1.445000 ;
      RECT 1704.210000  0.725000 1705.040000 0.735000 ;
      RECT 1704.210000  0.735000 1706.515000 0.905000 ;
      RECT 1704.240000  1.445000 1706.515000 1.625000 ;
      RECT 1704.240000  1.625000 1705.470000 1.665000 ;
      RECT 1704.240000  1.665000 1704.530000 2.125000 ;
      RECT 1704.320000  0.085000 1704.490000 0.555000 ;
      RECT 1704.660000  0.255000 1705.040000 0.725000 ;
      RECT 1704.750000  1.835000 1705.000000 2.295000 ;
      RECT 1705.220000  1.665000 1705.470000 2.125000 ;
      RECT 1705.260000  0.085000 1705.430000 0.555000 ;
      RECT 1705.600000  0.255000 1705.980000 0.735000 ;
      RECT 1705.690000  1.795000 1705.940000 2.295000 ;
      RECT 1706.110000  1.625000 1706.515000 2.465000 ;
      RECT 1706.195000  0.905000 1706.515000 1.445000 ;
      RECT 1706.200000  0.085000 1706.370000 0.555000 ;
      RECT 1706.685000  0.085000 1706.975000 0.810000 ;
      RECT 1706.685000  1.470000 1706.975000 2.635000 ;
      RECT 1707.145000  0.350000 1707.650000 0.925000 ;
      RECT 1707.145000  0.925000 1707.460000 1.440000 ;
      RECT 1707.145000  1.440000 1707.670000 2.465000 ;
      RECT 1707.860000  0.695000 1708.510000 0.865000 ;
      RECT 1707.860000  0.865000 1708.060000 1.875000 ;
      RECT 1707.860000  1.875000 1708.630000 2.045000 ;
      RECT 1707.870000  0.085000 1708.120000 0.525000 ;
      RECT 1707.890000  2.215000 1708.225000 2.635000 ;
      RECT 1708.290000  0.255000 1709.950000 0.425000 ;
      RECT 1708.290000  0.425000 1708.510000 0.695000 ;
      RECT 1708.295000  1.535000 1710.045000 1.705000 ;
      RECT 1708.410000  2.045000 1708.630000 2.235000 ;
      RECT 1708.410000  2.235000 1710.105000 2.405000 ;
      RECT 1708.680000  0.595000 1708.850000 1.535000 ;
      RECT 1709.020000  0.995000 1709.705000 1.325000 ;
      RECT 1709.030000  1.895000 1710.435000 2.065000 ;
      RECT 1709.130000  0.655000 1710.340000 0.825000 ;
      RECT 1709.550000  0.425000 1709.950000 0.455000 ;
      RECT 1709.875000  0.995000 1710.200000 1.325000 ;
      RECT 1709.875000  1.325000 1710.045000 1.535000 ;
      RECT 1710.120000  0.255000 1711.020000 0.425000 ;
      RECT 1710.120000  0.425000 1710.340000 0.655000 ;
      RECT 1710.265000  1.525000 1710.795000 1.695000 ;
      RECT 1710.265000  1.695000 1710.435000 1.895000 ;
      RECT 1710.370000  2.235000 1710.775000 2.405000 ;
      RECT 1710.510000  0.595000 1710.680000 1.375000 ;
      RECT 1710.510000  1.375000 1710.795000 1.525000 ;
      RECT 1710.605000  1.895000 1711.880000 2.065000 ;
      RECT 1710.605000  2.065000 1710.775000 2.235000 ;
      RECT 1710.850000  0.425000 1711.020000 1.035000 ;
      RECT 1710.850000  1.035000 1711.135000 1.205000 ;
      RECT 1710.945000  2.235000 1711.275000 2.635000 ;
      RECT 1710.965000  1.205000 1711.135000 1.895000 ;
      RECT 1711.190000  0.085000 1711.360000 0.865000 ;
      RECT 1711.365000  1.445000 1711.880000 1.715000 ;
      RECT 1711.590000  0.415000 1711.880000 1.445000 ;
      RECT 1711.710000  2.065000 1711.880000 2.275000 ;
      RECT 1711.710000  2.275000 1715.005000 2.445000 ;
      RECT 1712.055000  0.265000 1712.470000 0.485000 ;
      RECT 1712.055000  0.485000 1712.275000 0.595000 ;
      RECT 1712.055000  0.595000 1712.225000 2.105000 ;
      RECT 1712.395000  0.720000 1712.860000 0.825000 ;
      RECT 1712.395000  0.825000 1712.665000 0.890000 ;
      RECT 1712.395000  0.890000 1712.565000 2.275000 ;
      RECT 1712.445000  0.655000 1712.860000 0.720000 ;
      RECT 1712.690000  0.320000 1712.860000 0.655000 ;
      RECT 1712.805000  1.445000 1713.635000 1.615000 ;
      RECT 1712.805000  1.615000 1713.220000 2.045000 ;
      RECT 1712.820000  0.995000 1713.245000 1.270000 ;
      RECT 1713.030000  0.630000 1713.245000 0.995000 ;
      RECT 1713.465000  0.255000 1714.660000 0.425000 ;
      RECT 1713.465000  0.425000 1713.635000 1.445000 ;
      RECT 1713.805000  0.595000 1713.975000 1.935000 ;
      RECT 1713.805000  1.935000 1716.625000 2.105000 ;
      RECT 1714.145000  0.425000 1714.660000 0.465000 ;
      RECT 1714.145000  0.995000 1714.365000 1.445000 ;
      RECT 1714.145000  1.445000 1714.775000 1.725000 ;
      RECT 1714.535000  0.730000 1714.740000 0.945000 ;
      RECT 1714.535000  0.945000 1714.845000 1.275000 ;
      RECT 1714.995000  1.495000 1716.175000 1.705000 ;
      RECT 1715.035000  0.295000 1715.325000 0.735000 ;
      RECT 1715.035000  0.735000 1716.175000 0.750000 ;
      RECT 1715.065000  1.075000 1715.755000 1.325000 ;
      RECT 1715.075000  0.750000 1716.175000 0.905000 ;
      RECT 1715.415000  2.275000 1716.110000 2.635000 ;
      RECT 1715.545000  0.085000 1715.995000 0.565000 ;
      RECT 1716.005000  0.905000 1716.175000 0.995000 ;
      RECT 1716.005000  0.995000 1716.285000 1.325000 ;
      RECT 1716.005000  1.325000 1716.175000 1.495000 ;
      RECT 1716.090000  1.875000 1716.625000 1.935000 ;
      RECT 1716.325000  0.255000 1716.625000 0.585000 ;
      RECT 1716.330000  2.105000 1716.625000 2.465000 ;
      RECT 1716.455000  0.585000 1716.625000 1.875000 ;
      RECT 1716.805000  0.085000 1717.095000 0.810000 ;
      RECT 1716.805000  1.470000 1717.095000 2.635000 ;
      RECT 1717.285000  0.085000 1717.615000 0.465000 ;
      RECT 1717.285000  2.215000 1717.615000 2.635000 ;
      RECT 1717.510000  0.660000 1718.110000 0.925000 ;
      RECT 1717.510000  0.925000 1717.875000 1.440000 ;
      RECT 1717.510000  1.440000 1718.085000 2.045000 ;
      RECT 1717.835000  2.045000 1718.085000 2.465000 ;
      RECT 1717.860000  0.350000 1718.110000 0.660000 ;
      RECT 1718.275000  0.995000 1718.475000 1.325000 ;
      RECT 1718.285000  0.085000 1718.535000 0.525000 ;
      RECT 1718.305000  0.695000 1718.925000 0.865000 ;
      RECT 1718.305000  0.865000 1718.475000 0.995000 ;
      RECT 1718.305000  1.325000 1718.475000 1.875000 ;
      RECT 1718.305000  1.875000 1719.045000 2.045000 ;
      RECT 1718.305000  2.215000 1718.640000 2.635000 ;
      RECT 1718.705000  0.255000 1720.370000 0.425000 ;
      RECT 1718.705000  0.425000 1718.925000 0.695000 ;
      RECT 1718.710000  1.535000 1720.460000 1.705000 ;
      RECT 1718.825000  2.045000 1719.045000 2.235000 ;
      RECT 1718.825000  2.235000 1720.520000 2.405000 ;
      RECT 1719.095000  0.595000 1719.265000 1.535000 ;
      RECT 1719.435000  0.995000 1720.120000 1.325000 ;
      RECT 1719.445000  1.895000 1720.850000 2.065000 ;
      RECT 1719.545000  0.655000 1720.755000 0.825000 ;
      RECT 1719.965000  0.425000 1720.370000 0.455000 ;
      RECT 1720.290000  0.995000 1720.615000 1.325000 ;
      RECT 1720.290000  1.325000 1720.460000 1.535000 ;
      RECT 1720.540000  0.255000 1721.435000 0.425000 ;
      RECT 1720.540000  0.425000 1720.755000 0.655000 ;
      RECT 1720.680000  1.525000 1721.210000 1.695000 ;
      RECT 1720.680000  1.695000 1720.850000 1.895000 ;
      RECT 1720.785000  2.235000 1721.190000 2.405000 ;
      RECT 1720.925000  0.595000 1721.095000 1.375000 ;
      RECT 1720.925000  1.375000 1721.210000 1.525000 ;
      RECT 1721.020000  1.895000 1722.295000 2.065000 ;
      RECT 1721.020000  2.065000 1721.190000 2.235000 ;
      RECT 1721.265000  0.425000 1721.435000 1.035000 ;
      RECT 1721.265000  1.035000 1721.550000 1.205000 ;
      RECT 1721.360000  2.235000 1721.690000 2.635000 ;
      RECT 1721.380000  1.205000 1721.550000 1.895000 ;
      RECT 1721.605000  0.085000 1721.775000 0.865000 ;
      RECT 1721.780000  1.445000 1722.295000 1.715000 ;
      RECT 1722.005000  0.415000 1722.295000 1.445000 ;
      RECT 1722.125000  2.065000 1722.295000 2.275000 ;
      RECT 1722.125000  2.275000 1725.420000 2.445000 ;
      RECT 1722.470000  0.265000 1722.885000 0.485000 ;
      RECT 1722.470000  0.485000 1722.690000 0.595000 ;
      RECT 1722.470000  0.595000 1722.640000 2.105000 ;
      RECT 1722.810000  0.720000 1723.275000 0.825000 ;
      RECT 1722.810000  0.825000 1723.080000 0.890000 ;
      RECT 1722.810000  0.890000 1722.980000 2.275000 ;
      RECT 1722.860000  0.655000 1723.275000 0.720000 ;
      RECT 1723.105000  0.320000 1723.275000 0.655000 ;
      RECT 1723.220000  1.445000 1724.050000 1.615000 ;
      RECT 1723.220000  1.615000 1723.635000 2.045000 ;
      RECT 1723.235000  0.995000 1723.660000 1.270000 ;
      RECT 1723.445000  0.630000 1723.660000 0.995000 ;
      RECT 1723.880000  0.255000 1725.075000 0.425000 ;
      RECT 1723.880000  0.425000 1724.050000 1.445000 ;
      RECT 1724.220000  0.595000 1724.390000 1.935000 ;
      RECT 1724.220000  1.935000 1726.730000 2.105000 ;
      RECT 1724.560000  0.425000 1725.075000 0.465000 ;
      RECT 1724.560000  0.995000 1724.780000 1.445000 ;
      RECT 1724.560000  1.445000 1725.190000 1.665000 ;
      RECT 1724.950000  0.730000 1725.155000 0.945000 ;
      RECT 1724.950000  0.945000 1725.270000 1.275000 ;
      RECT 1725.410000  1.495000 1726.280000 1.705000 ;
      RECT 1725.450000  0.295000 1725.740000 0.735000 ;
      RECT 1725.450000  0.735000 1726.280000 0.750000 ;
      RECT 1725.480000  1.075000 1725.940000 1.325000 ;
      RECT 1725.490000  0.750000 1726.280000 0.905000 ;
      RECT 1725.830000  2.275000 1726.215000 2.635000 ;
      RECT 1725.960000  0.085000 1726.130000 0.565000 ;
      RECT 1726.110000  0.905000 1726.280000 0.995000 ;
      RECT 1726.110000  0.995000 1726.390000 1.325000 ;
      RECT 1726.110000  1.325000 1726.280000 1.495000 ;
      RECT 1726.195000  1.875000 1726.730000 1.935000 ;
      RECT 1726.430000  0.255000 1726.730000 0.585000 ;
      RECT 1726.435000  2.105000 1726.730000 2.465000 ;
      RECT 1726.560000  0.585000 1726.730000 1.875000 ;
      RECT 1726.925000  0.085000 1727.215000 0.810000 ;
      RECT 1726.925000  1.470000 1727.215000 2.635000 ;
      RECT 1727.475000  0.085000 1727.645000 0.545000 ;
      RECT 1727.575000  2.135000 1727.745000 2.635000 ;
      RECT 1727.945000  0.350000 1728.115000 0.660000 ;
      RECT 1727.945000  0.660000 1729.055000 0.925000 ;
      RECT 1728.045000  1.440000 1728.870000 1.455000 ;
      RECT 1728.045000  1.455000 1729.155000 2.045000 ;
      RECT 1728.045000  2.045000 1728.215000 2.465000 ;
      RECT 1728.285000  0.085000 1728.665000 0.465000 ;
      RECT 1728.435000  2.215000 1728.765000 2.635000 ;
      RECT 1728.505000  0.925000 1728.870000 1.440000 ;
      RECT 1728.885000  0.350000 1729.055000 0.660000 ;
      RECT 1728.985000  2.045000 1729.155000 2.465000 ;
      RECT 1729.320000  0.965000 1729.545000 1.325000 ;
      RECT 1729.355000  0.085000 1729.525000 0.525000 ;
      RECT 1729.375000  0.695000 1729.865000 0.865000 ;
      RECT 1729.375000  0.865000 1729.545000 0.965000 ;
      RECT 1729.375000  1.325000 1729.545000 1.875000 ;
      RECT 1729.375000  1.875000 1730.095000 2.045000 ;
      RECT 1729.375000  2.215000 1729.705000 2.635000 ;
      RECT 1729.695000  0.255000 1731.360000 0.425000 ;
      RECT 1729.695000  0.425000 1729.865000 0.695000 ;
      RECT 1729.870000  1.535000 1731.455000 1.705000 ;
      RECT 1729.875000  2.045000 1730.095000 2.235000 ;
      RECT 1729.875000  2.235000 1731.515000 2.405000 ;
      RECT 1730.090000  0.595000 1730.260000 1.535000 ;
      RECT 1730.430000  0.995000 1731.115000 1.325000 ;
      RECT 1730.440000  1.895000 1731.845000 2.065000 ;
      RECT 1730.540000  0.655000 1731.750000 0.825000 ;
      RECT 1730.960000  0.425000 1731.360000 0.455000 ;
      RECT 1731.285000  0.995000 1731.705000 1.325000 ;
      RECT 1731.285000  1.325000 1731.455000 1.535000 ;
      RECT 1731.530000  0.255000 1732.430000 0.425000 ;
      RECT 1731.530000  0.425000 1731.750000 0.655000 ;
      RECT 1731.675000  1.525000 1732.205000 1.695000 ;
      RECT 1731.675000  1.695000 1731.845000 1.895000 ;
      RECT 1731.780000  2.235000 1732.185000 2.405000 ;
      RECT 1731.920000  0.595000 1732.090000 1.375000 ;
      RECT 1731.920000  1.375000 1732.205000 1.525000 ;
      RECT 1732.015000  1.895000 1733.290000 2.065000 ;
      RECT 1732.015000  2.065000 1732.185000 2.235000 ;
      RECT 1732.260000  0.425000 1732.430000 1.035000 ;
      RECT 1732.260000  1.035000 1732.515000 1.040000 ;
      RECT 1732.260000  1.040000 1732.530000 1.045000 ;
      RECT 1732.260000  1.045000 1732.540000 1.050000 ;
      RECT 1732.260000  1.050000 1732.545000 1.205000 ;
      RECT 1732.355000  2.235000 1732.685000 2.635000 ;
      RECT 1732.375000  1.205000 1732.545000 1.895000 ;
      RECT 1732.600000  0.085000 1732.770000 0.885000 ;
      RECT 1732.775000  1.445000 1733.290000 1.715000 ;
      RECT 1733.000000  0.415000 1733.290000 1.445000 ;
      RECT 1733.120000  2.065000 1733.290000 2.275000 ;
      RECT 1733.120000  2.275000 1736.415000 2.445000 ;
      RECT 1733.465000  0.265000 1733.880000 0.485000 ;
      RECT 1733.465000  0.485000 1733.685000 0.595000 ;
      RECT 1733.465000  0.595000 1733.635000 2.105000 ;
      RECT 1733.825000  0.720000 1734.270000 0.825000 ;
      RECT 1733.825000  0.825000 1734.075000 0.890000 ;
      RECT 1733.825000  0.890000 1733.995000 2.275000 ;
      RECT 1733.855000  0.655000 1734.270000 0.720000 ;
      RECT 1734.100000  0.320000 1734.270000 0.655000 ;
      RECT 1734.215000  1.445000 1735.045000 1.615000 ;
      RECT 1734.215000  1.615000 1734.630000 2.045000 ;
      RECT 1734.230000  0.995000 1734.655000 1.270000 ;
      RECT 1734.440000  0.630000 1734.655000 0.995000 ;
      RECT 1734.875000  0.255000 1736.070000 0.425000 ;
      RECT 1734.875000  0.425000 1735.045000 1.445000 ;
      RECT 1735.215000  0.595000 1735.385000 1.935000 ;
      RECT 1735.215000  1.935000 1737.725000 2.105000 ;
      RECT 1735.555000  0.425000 1736.070000 0.465000 ;
      RECT 1735.555000  0.995000 1735.775000 1.445000 ;
      RECT 1735.555000  1.445000 1735.940000 1.615000 ;
      RECT 1735.945000  0.730000 1736.150000 0.945000 ;
      RECT 1735.945000  0.945000 1736.255000 1.275000 ;
      RECT 1736.405000  1.495000 1737.275000 1.705000 ;
      RECT 1736.445000  0.295000 1736.735000 0.735000 ;
      RECT 1736.445000  0.735000 1737.275000 0.750000 ;
      RECT 1736.475000  1.075000 1736.935000 1.325000 ;
      RECT 1736.485000  0.750000 1737.275000 0.905000 ;
      RECT 1736.915000  2.275000 1737.245000 2.635000 ;
      RECT 1736.995000  0.085000 1737.165000 0.565000 ;
      RECT 1737.105000  0.905000 1737.275000 0.995000 ;
      RECT 1737.105000  0.995000 1737.335000 1.325000 ;
      RECT 1737.105000  1.325000 1737.275000 1.495000 ;
      RECT 1737.190000  1.875000 1737.725000 1.935000 ;
      RECT 1737.465000  0.255000 1737.725000 0.585000 ;
      RECT 1737.465000  2.105000 1737.725000 2.465000 ;
      RECT 1737.555000  0.585000 1737.725000 1.875000 ;
      RECT 1737.965000  0.085000 1738.255000 0.810000 ;
      RECT 1737.965000  1.470000 1738.255000 2.635000 ;
      RECT 1738.430000  1.795000 1739.255000 1.965000 ;
      RECT 1738.430000  1.965000 1738.685000 2.465000 ;
      RECT 1738.435000  0.345000 1738.685000 0.635000 ;
      RECT 1738.435000  0.635000 1739.225000 0.805000 ;
      RECT 1738.480000  0.975000 1738.830000 1.625000 ;
      RECT 1738.855000  0.085000 1739.235000 0.465000 ;
      RECT 1738.870000  2.135000 1739.250000 2.635000 ;
      RECT 1739.050000  0.805000 1739.225000 0.995000 ;
      RECT 1739.050000  0.995000 1739.365000 1.325000 ;
      RECT 1739.050000  1.325000 1739.255000 1.795000 ;
      RECT 1739.455000  0.345000 1739.705000 0.675000 ;
      RECT 1739.475000  1.730000 1739.705000 2.465000 ;
      RECT 1739.535000  0.675000 1739.705000 1.730000 ;
      RECT 1739.925000  1.070000 1740.330000 1.335000 ;
      RECT 1739.925000  1.335000 1740.560000 1.745000 ;
      RECT 1740.035000  0.395000 1740.205000 0.730000 ;
      RECT 1740.035000  0.730000 1740.775000 0.900000 ;
      RECT 1740.375000  0.085000 1740.755000 0.560000 ;
      RECT 1740.450000  1.915000 1741.070000 2.085000 ;
      RECT 1740.450000  2.085000 1740.720000 2.400000 ;
      RECT 1740.605000  0.900000 1740.775000 0.995000 ;
      RECT 1740.605000  0.995000 1741.785000 1.165000 ;
      RECT 1740.815000  1.165000 1741.785000 1.185000 ;
      RECT 1740.815000  1.185000 1741.070000 1.915000 ;
      RECT 1740.940000  2.255000 1741.270000 2.635000 ;
      RECT 1740.995000  0.085000 1741.375000 0.825000 ;
      RECT 1741.460000  1.355000 1741.995000 2.465000 ;
      RECT 1741.615000  0.255000 1742.775000 0.425000 ;
      RECT 1741.615000  0.425000 1741.785000 0.995000 ;
      RECT 1742.005000  0.675000 1742.385000 1.075000 ;
      RECT 1742.210000  1.075000 1742.385000 1.935000 ;
      RECT 1742.210000  1.935000 1743.990000 2.105000 ;
      RECT 1742.210000  2.105000 1742.380000 2.465000 ;
      RECT 1742.605000  0.425000 1742.775000 1.685000 ;
      RECT 1742.950000  0.710000 1743.295000 1.700000 ;
      RECT 1743.195000  2.275000 1743.545000 2.635000 ;
      RECT 1743.345000  0.085000 1743.690000 0.540000 ;
      RECT 1743.480000  0.715000 1744.060000 0.895000 ;
      RECT 1743.480000  0.895000 1743.650000 1.935000 ;
      RECT 1743.820000  1.065000 1743.990000 1.395000 ;
      RECT 1743.820000  2.105000 1743.990000 2.185000 ;
      RECT 1743.820000  2.185000 1744.190000 2.435000 ;
      RECT 1743.890000  0.335000 1744.230000 0.505000 ;
      RECT 1743.890000  0.505000 1744.060000 0.715000 ;
      RECT 1744.160000  1.575000 1744.460000 1.955000 ;
      RECT 1744.240000  0.705000 1744.990000 1.035000 ;
      RECT 1744.240000  1.035000 1744.460000 1.575000 ;
      RECT 1744.435000  2.135000 1744.800000 2.465000 ;
      RECT 1744.450000  0.305000 1745.350000 0.475000 ;
      RECT 1744.630000  1.215000 1746.490000 1.385000 ;
      RECT 1744.630000  1.385000 1744.800000 2.135000 ;
      RECT 1745.020000  1.935000 1746.280000 2.105000 ;
      RECT 1745.020000  2.105000 1745.190000 2.375000 ;
      RECT 1745.180000  0.475000 1745.350000 1.215000 ;
      RECT 1745.300000  1.595000 1746.880000 1.765000 ;
      RECT 1745.475000  2.355000 1745.805000 2.635000 ;
      RECT 1745.570000  0.765000 1746.150000 1.045000 ;
      RECT 1746.030000  0.085000 1746.360000 0.545000 ;
      RECT 1746.110000  2.105000 1746.280000 2.375000 ;
      RECT 1746.320000  1.005000 1746.490000 1.215000 ;
      RECT 1746.490000  2.175000 1746.910000 2.635000 ;
      RECT 1746.570000  0.275000 1746.950000 0.445000 ;
      RECT 1746.570000  0.445000 1746.880000 0.835000 ;
      RECT 1746.570000  1.765000 1746.880000 1.835000 ;
      RECT 1746.570000  1.835000 1747.325000 2.005000 ;
      RECT 1746.710000  0.835000 1746.880000 1.595000 ;
      RECT 1747.050000  0.705000 1747.310000 1.495000 ;
      RECT 1747.050000  1.495000 1747.785000 1.660000 ;
      RECT 1747.050000  1.660000 1748.185000 1.665000 ;
      RECT 1747.120000  0.255000 1748.230000 0.535000 ;
      RECT 1747.155000  2.005000 1747.325000 2.465000 ;
      RECT 1747.525000  1.665000 1748.185000 1.955000 ;
      RECT 1747.535000  2.125000 1748.555000 2.465000 ;
      RECT 1747.575000  0.920000 1747.745000 1.325000 ;
      RECT 1748.010000  0.535000 1748.230000 1.315000 ;
      RECT 1748.010000  1.315000 1748.625000 1.485000 ;
      RECT 1748.380000  1.485000 1748.625000 1.575000 ;
      RECT 1748.380000  1.575000 1749.710000 1.745000 ;
      RECT 1748.380000  1.745000 1748.555000 2.125000 ;
      RECT 1748.450000  0.085000 1748.670000 0.525000 ;
      RECT 1748.490000  0.695000 1749.070000 0.865000 ;
      RECT 1748.490000  0.865000 1748.710000 1.145000 ;
      RECT 1748.755000  2.195000 1749.005000 2.635000 ;
      RECT 1748.900000  0.295000 1750.075000 0.465000 ;
      RECT 1748.900000  0.465000 1749.070000 0.695000 ;
      RECT 1748.940000  1.065000 1749.710000 1.275000 ;
      RECT 1749.250000  1.915000 1750.070000 2.085000 ;
      RECT 1749.250000  2.085000 1749.420000 2.375000 ;
      RECT 1749.405000  0.635000 1749.710000 1.065000 ;
      RECT 1749.595000  2.255000 1749.975000 2.635000 ;
      RECT 1749.900000  0.465000 1750.075000 0.995000 ;
      RECT 1749.900000  0.995000 1750.545000 1.325000 ;
      RECT 1749.900000  1.325000 1750.070000 1.915000 ;
      RECT 1750.245000  0.085000 1750.415000 0.545000 ;
      RECT 1750.245000  1.495000 1750.495000 2.635000 ;
      RECT 1750.765000  0.265000 1751.095000 0.995000 ;
      RECT 1750.765000  0.995000 1752.035000 1.325000 ;
      RECT 1750.765000  1.325000 1751.095000 2.325000 ;
      RECT 1751.315000  0.085000 1751.485000 0.545000 ;
      RECT 1751.315000  1.495000 1751.565000 2.635000 ;
      RECT 1751.785000  0.265000 1752.035000 0.995000 ;
      RECT 1751.785000  1.325000 1752.035000 2.325000 ;
      RECT 1752.255000  0.085000 1752.425000 0.545000 ;
      RECT 1752.255000  1.495000 1752.505000 2.635000 ;
      RECT 1752.685000  0.085000 1752.975000 0.810000 ;
      RECT 1752.685000  1.470000 1752.975000 2.635000 ;
      RECT 1753.160000  1.075000 1753.650000 1.325000 ;
      RECT 1753.160000  1.325000 1753.425000 1.685000 ;
      RECT 1753.185000  0.355000 1753.515000 0.715000 ;
      RECT 1753.185000  0.715000 1754.755000 0.905000 ;
      RECT 1753.185000  1.965000 1753.465000 2.635000 ;
      RECT 1753.685000  1.575000 1754.755000 1.745000 ;
      RECT 1753.685000  1.745000 1753.985000 2.295000 ;
      RECT 1753.915000  1.075000 1754.335000 1.325000 ;
      RECT 1754.235000  0.085000 1754.485000 0.545000 ;
      RECT 1754.235000  1.915000 1754.565000 2.635000 ;
      RECT 1754.585000  0.905000 1754.755000 1.575000 ;
      RECT 1754.655000  0.255000 1755.265000 0.545000 ;
      RECT 1754.805000  1.915000 1755.265000 2.465000 ;
      RECT 1755.015000  0.545000 1755.265000 1.915000 ;
      RECT 1755.445000  0.085000 1755.735000 0.810000 ;
      RECT 1755.445000  1.470000 1755.735000 2.635000 ;
      RECT 1755.910000  0.085000 1756.245000 0.590000 ;
      RECT 1755.965000  0.765000 1756.265000 1.615000 ;
      RECT 1755.995000  1.785000 1756.715000 2.015000 ;
      RECT 1755.995000  2.015000 1756.165000 2.445000 ;
      RECT 1756.335000  2.185000 1756.715000 2.635000 ;
      RECT 1756.465000  0.280000 1756.705000 0.805000 ;
      RECT 1756.465000  0.805000 1757.000000 1.135000 ;
      RECT 1756.465000  1.135000 1756.715000 1.785000 ;
      RECT 1756.885000  1.305000 1758.295000 1.325000 ;
      RECT 1756.885000  1.325000 1757.705000 1.475000 ;
      RECT 1756.885000  1.475000 1757.155000 2.420000 ;
      RECT 1756.985000  0.270000 1757.155000 0.415000 ;
      RECT 1756.985000  0.415000 1757.410000 0.610000 ;
      RECT 1757.170000  0.610000 1757.410000 0.945000 ;
      RECT 1757.170000  0.945000 1758.295000 1.305000 ;
      RECT 1757.325000  1.645000 1757.655000 1.955000 ;
      RECT 1757.385000  2.165000 1758.145000 2.635000 ;
      RECT 1757.890000  0.085000 1758.220000 0.580000 ;
      RECT 1758.325000  1.580000 1758.900000 2.365000 ;
      RECT 1758.440000  0.255000 1758.900000 0.775000 ;
      RECT 1758.725000  0.775000 1758.900000 1.580000 ;
      RECT 1759.125000  0.085000 1759.415000 0.810000 ;
      RECT 1759.125000  1.470000 1759.415000 2.635000 ;
      RECT 1759.590000  1.075000 1759.925000 1.325000 ;
      RECT 1759.590000  1.495000 1759.845000 2.635000 ;
      RECT 1759.610000  0.265000 1759.920000 0.735000 ;
      RECT 1759.610000  0.735000 1760.395000 0.905000 ;
      RECT 1760.040000  2.085000 1761.395000 2.415000 ;
      RECT 1760.140000  0.085000 1760.875000 0.565000 ;
      RECT 1760.145000  0.905000 1760.395000 0.995000 ;
      RECT 1760.145000  0.995000 1760.885000 1.325000 ;
      RECT 1760.145000  1.325000 1760.315000 1.885000 ;
      RECT 1760.540000  1.495000 1762.005000 1.665000 ;
      RECT 1760.540000  1.665000 1760.960000 1.915000 ;
      RECT 1761.155000  0.305000 1761.325000 0.655000 ;
      RECT 1761.155000  0.655000 1762.005000 0.825000 ;
      RECT 1761.495000  0.085000 1761.925000 0.485000 ;
      RECT 1761.625000  1.835000 1761.905000 2.635000 ;
      RECT 1761.835000  0.825000 1762.005000 1.495000 ;
      RECT 1762.175000  0.415000 1762.580000 0.760000 ;
      RECT 1762.175000  1.495000 1762.580000 2.465000 ;
      RECT 1762.410000  0.760000 1762.580000 1.495000 ;
      RECT 1762.805000  0.085000 1763.095000 0.810000 ;
      RECT 1762.805000  1.470000 1763.095000 2.635000 ;
      RECT 1763.265000  0.765000 1763.620000 1.325000 ;
      RECT 1763.330000  1.495000 1764.885000 1.665000 ;
      RECT 1763.330000  1.665000 1763.720000 1.840000 ;
      RECT 1763.370000  0.085000 1763.610000 0.595000 ;
      RECT 1763.790000  0.265000 1764.120000 0.595000 ;
      RECT 1763.790000  0.595000 1764.010000 1.495000 ;
      RECT 1764.180000  0.765000 1764.495000 1.325000 ;
      RECT 1764.365000  1.835000 1764.695000 2.635000 ;
      RECT 1764.400000  0.085000 1764.615000 0.595000 ;
      RECT 1764.715000  0.995000 1764.885000 1.495000 ;
      RECT 1764.845000  0.255000 1765.395000 0.825000 ;
      RECT 1764.975000  1.845000 1765.395000 2.465000 ;
      RECT 1765.080000  0.825000 1765.395000 1.845000 ;
      RECT 1765.565000  0.085000 1765.855000 0.810000 ;
      RECT 1765.565000  1.470000 1765.855000 2.635000 ;
      RECT 1766.040000  0.725000 1766.265000 1.325000 ;
      RECT 1766.270000  0.370000 1766.615000 0.545000 ;
      RECT 1766.355000  1.510000 1767.795000 1.680000 ;
      RECT 1766.355000  1.680000 1766.615000 1.905000 ;
      RECT 1766.435000  0.545000 1766.615000 1.510000 ;
      RECT 1766.845000  0.085000 1767.055000 0.895000 ;
      RECT 1766.865000  1.855000 1767.195000 2.635000 ;
      RECT 1766.950000  1.065000 1767.365000 1.325000 ;
      RECT 1767.225000  0.255000 1767.575000 0.645000 ;
      RECT 1767.225000  0.645000 1768.145000 0.815000 ;
      RECT 1767.575000  0.985000 1767.795000 1.510000 ;
      RECT 1767.695000  1.850000 1768.145000 2.465000 ;
      RECT 1767.745000  0.085000 1768.075000 0.475000 ;
      RECT 1767.965000  0.815000 1768.145000 1.850000 ;
      RECT 1768.325000  0.085000 1768.615000 0.810000 ;
      RECT 1768.325000  1.470000 1768.615000 2.635000 ;
      RECT 1768.785000  0.085000 1769.065000 0.895000 ;
      RECT 1768.785000  1.445000 1770.045000 1.655000 ;
      RECT 1768.785000  1.655000 1769.105000 2.465000 ;
      RECT 1769.180000  1.065000 1769.670000 1.275000 ;
      RECT 1769.235000  0.255000 1769.615000 0.725000 ;
      RECT 1769.235000  0.725000 1770.555000 0.895000 ;
      RECT 1769.325000  1.825000 1769.575000 2.635000 ;
      RECT 1769.795000  1.655000 1770.045000 2.295000 ;
      RECT 1769.795000  2.295000 1771.025000 2.465000 ;
      RECT 1769.835000  0.085000 1770.005000 0.555000 ;
      RECT 1770.175000  0.255000 1770.555000 0.725000 ;
      RECT 1770.225000  0.895000 1770.515000 2.125000 ;
      RECT 1770.735000  1.445000 1770.990000 1.890000 ;
      RECT 1770.735000  1.890000 1771.025000 2.295000 ;
      RECT 1770.775000  0.085000 1770.945000 0.895000 ;
      RECT 1770.775000  1.075000 1771.330000 1.245000 ;
      RECT 1771.115000  0.725000 1771.465000 0.895000 ;
      RECT 1771.115000  0.895000 1771.330000 1.075000 ;
      RECT 1771.160000  1.245000 1771.330000 1.445000 ;
      RECT 1771.160000  1.445000 1771.465000 1.615000 ;
      RECT 1771.295000  0.445000 1771.465000 0.725000 ;
      RECT 1771.295000  1.615000 1771.465000 2.460000 ;
      RECT 1771.500000  1.065000 1772.255000 1.275000 ;
      RECT 1771.725000  0.085000 1771.980000 0.845000 ;
      RECT 1771.725000  2.145000 1771.975000 2.635000 ;
      RECT 1772.040000  1.275000 1772.255000 1.965000 ;
      RECT 1772.465000  0.085000 1772.755000 0.810000 ;
      RECT 1772.465000  1.470000 1772.755000 2.635000 ;
      RECT 1772.925000  0.085000 1773.205000 0.905000 ;
      RECT 1772.925000  1.455000 1775.165000 1.665000 ;
      RECT 1772.925000  1.665000 1773.205000 2.465000 ;
      RECT 1773.200000  1.075000 1774.790000 1.275000 ;
      RECT 1773.375000  0.255000 1773.755000 0.725000 ;
      RECT 1773.375000  0.725000 1776.575000 0.905000 ;
      RECT 1773.375000  1.835000 1773.755000 2.635000 ;
      RECT 1773.975000  0.085000 1774.145000 0.555000 ;
      RECT 1773.975000  1.665000 1774.145000 2.465000 ;
      RECT 1774.315000  0.255000 1774.695000 0.725000 ;
      RECT 1774.315000  1.835000 1774.615000 2.635000 ;
      RECT 1774.785000  1.665000 1775.165000 2.295000 ;
      RECT 1774.785000  2.295000 1777.095000 2.465000 ;
      RECT 1774.915000  0.085000 1775.085000 0.555000 ;
      RECT 1775.255000  0.255000 1775.635000 0.725000 ;
      RECT 1775.385000  0.905000 1775.715000 1.445000 ;
      RECT 1775.385000  1.445000 1776.495000 1.745000 ;
      RECT 1775.385000  1.745000 1775.555000 2.125000 ;
      RECT 1775.725000  1.935000 1776.105000 2.295000 ;
      RECT 1775.855000  0.085000 1776.025000 0.555000 ;
      RECT 1775.935000  1.075000 1777.515000 1.275000 ;
      RECT 1776.195000  0.255000 1776.575000 0.725000 ;
      RECT 1776.325000  1.745000 1776.495000 2.125000 ;
      RECT 1776.665000  1.575000 1777.095000 2.295000 ;
      RECT 1776.795000  0.085000 1777.085000 0.905000 ;
      RECT 1777.265000  0.255000 1777.595000 0.815000 ;
      RECT 1777.265000  0.815000 1777.515000 1.075000 ;
      RECT 1777.265000  1.275000 1777.515000 1.575000 ;
      RECT 1777.265000  1.575000 1777.595000 2.465000 ;
      RECT 1777.685000  1.075000 1778.265000 1.320000 ;
      RECT 1777.815000  0.085000 1778.105000 0.905000 ;
      RECT 1777.815000  1.495000 1778.220000 2.635000 ;
      RECT 1778.445000  0.085000 1778.735000 0.810000 ;
      RECT 1778.445000  1.470000 1778.735000 2.635000 ;
      RECT 1778.905000  0.255000 1779.135000 1.065000 ;
      RECT 1778.905000  1.065000 1779.325000 1.285000 ;
      RECT 1778.945000  1.455000 1779.165000 2.635000 ;
      RECT 1779.305000  0.085000 1779.525000 0.895000 ;
      RECT 1779.335000  1.455000 1779.765000 2.465000 ;
      RECT 1779.545000  1.065000 1780.055000 1.075000 ;
      RECT 1779.545000  1.075000 1784.340000 1.285000 ;
      RECT 1779.545000  1.285000 1779.765000 1.455000 ;
      RECT 1779.695000  0.255000 1780.055000 1.065000 ;
      RECT 1779.985000  1.455000 1780.280000 2.635000 ;
      RECT 1780.265000  0.085000 1780.775000 0.905000 ;
      RECT 1780.495000  1.455000 1784.575000 1.665000 ;
      RECT 1780.495000  1.665000 1780.815000 2.465000 ;
      RECT 1780.945000  0.255000 1781.325000 0.725000 ;
      RECT 1780.945000  0.725000 1788.385000 0.905000 ;
      RECT 1781.035000  1.835000 1781.285000 2.635000 ;
      RECT 1781.505000  1.665000 1781.755000 2.465000 ;
      RECT 1781.545000  0.085000 1781.715000 0.555000 ;
      RECT 1781.885000  0.255000 1782.265000 0.725000 ;
      RECT 1781.975000  1.835000 1782.225000 2.635000 ;
      RECT 1782.445000  1.665000 1782.695000 2.465000 ;
      RECT 1782.485000  0.085000 1782.655000 0.555000 ;
      RECT 1782.825000  0.255000 1783.205000 0.725000 ;
      RECT 1782.915000  1.835000 1783.165000 2.635000 ;
      RECT 1783.385000  1.665000 1783.635000 2.465000 ;
      RECT 1783.425000  0.085000 1783.595000 0.555000 ;
      RECT 1783.765000  0.255000 1784.145000 0.725000 ;
      RECT 1783.855000  1.835000 1784.105000 2.635000 ;
      RECT 1784.325000  1.665000 1784.575000 2.295000 ;
      RECT 1784.325000  2.295000 1788.335000 2.465000 ;
      RECT 1784.365000  0.085000 1784.535000 0.555000 ;
      RECT 1784.610000  1.075000 1787.700000 1.275000 ;
      RECT 1784.705000  0.255000 1785.085000 0.725000 ;
      RECT 1784.795000  1.445000 1788.385000 1.615000 ;
      RECT 1784.795000  1.615000 1785.045000 2.125000 ;
      RECT 1785.265000  1.785000 1785.515000 2.295000 ;
      RECT 1785.305000  0.085000 1785.475000 0.555000 ;
      RECT 1785.645000  0.255000 1786.025000 0.725000 ;
      RECT 1785.735000  1.615000 1785.985000 2.125000 ;
      RECT 1786.205000  1.785000 1786.455000 2.295000 ;
      RECT 1786.245000  0.085000 1786.415000 0.555000 ;
      RECT 1786.585000  0.255000 1786.965000 0.725000 ;
      RECT 1786.675000  1.615000 1786.925000 2.125000 ;
      RECT 1787.145000  1.785000 1787.395000 2.295000 ;
      RECT 1787.185000  0.085000 1787.355000 0.555000 ;
      RECT 1787.525000  0.255000 1787.905000 0.725000 ;
      RECT 1787.615000  1.615000 1787.865000 2.125000 ;
      RECT 1787.870000  0.905000 1788.385000 1.445000 ;
      RECT 1788.085000  1.785000 1788.335000 2.295000 ;
      RECT 1788.125000  0.085000 1788.395000 0.555000 ;
      RECT 1788.565000  0.085000 1788.855000 0.810000 ;
      RECT 1788.565000  1.470000 1788.855000 2.635000 ;
      RECT 1789.025000  0.255000 1789.255000 0.995000 ;
      RECT 1789.025000  0.995000 1789.605000 1.325000 ;
      RECT 1789.240000  1.495000 1789.455000 2.635000 ;
      RECT 1789.425000  0.085000 1789.805000 0.825000 ;
      RECT 1789.625000  1.495000 1790.055000 2.465000 ;
      RECT 1789.825000  1.065000 1791.325000 1.075000 ;
      RECT 1789.825000  1.075000 1799.420000 1.285000 ;
      RECT 1789.825000  1.285000 1790.055000 1.495000 ;
      RECT 1790.025000  0.255000 1790.285000 1.065000 ;
      RECT 1790.275000  1.455000 1790.495000 2.635000 ;
      RECT 1790.505000  0.085000 1790.805000 0.895000 ;
      RECT 1790.665000  1.285000 1791.095000 2.465000 ;
      RECT 1791.025000  0.255000 1791.325000 1.065000 ;
      RECT 1791.315000  1.455000 1791.610000 2.635000 ;
      RECT 1791.545000  0.085000 1792.095000 0.905000 ;
      RECT 1791.815000  1.455000 1799.655000 1.665000 ;
      RECT 1791.815000  1.665000 1792.135000 2.465000 ;
      RECT 1792.265000  0.255000 1792.645000 0.725000 ;
      RECT 1792.265000  0.725000 1807.245000 0.905000 ;
      RECT 1792.355000  1.835000 1792.605000 2.635000 ;
      RECT 1792.825000  1.665000 1793.075000 2.465000 ;
      RECT 1792.865000  0.085000 1793.035000 0.555000 ;
      RECT 1793.205000  0.255000 1793.585000 0.725000 ;
      RECT 1793.295000  1.835000 1793.545000 2.635000 ;
      RECT 1793.765000  1.665000 1794.015000 2.465000 ;
      RECT 1793.805000  0.085000 1793.975000 0.555000 ;
      RECT 1794.145000  0.255000 1794.525000 0.725000 ;
      RECT 1794.235000  1.835000 1794.485000 2.635000 ;
      RECT 1794.705000  1.665000 1794.955000 2.465000 ;
      RECT 1794.745000  0.085000 1794.915000 0.555000 ;
      RECT 1795.085000  0.255000 1795.465000 0.725000 ;
      RECT 1795.175000  1.835000 1795.425000 2.635000 ;
      RECT 1795.645000  1.665000 1795.895000 2.465000 ;
      RECT 1795.685000  0.085000 1795.855000 0.555000 ;
      RECT 1796.025000  0.255000 1796.405000 0.725000 ;
      RECT 1796.115000  1.835000 1796.365000 2.635000 ;
      RECT 1796.585000  1.665000 1796.835000 2.465000 ;
      RECT 1796.625000  0.085000 1796.795000 0.555000 ;
      RECT 1796.965000  0.255000 1797.345000 0.725000 ;
      RECT 1797.055000  1.835000 1797.305000 2.635000 ;
      RECT 1797.525000  1.665000 1797.775000 2.465000 ;
      RECT 1797.565000  0.085000 1797.735000 0.555000 ;
      RECT 1797.905000  0.255000 1798.285000 0.725000 ;
      RECT 1797.995000  1.835000 1798.245000 2.635000 ;
      RECT 1798.465000  1.665000 1798.715000 2.465000 ;
      RECT 1798.505000  0.085000 1798.675000 0.555000 ;
      RECT 1798.845000  0.255000 1799.225000 0.725000 ;
      RECT 1798.935000  1.835000 1799.185000 2.635000 ;
      RECT 1799.405000  1.665000 1799.655000 2.295000 ;
      RECT 1799.405000  2.295000 1807.175000 2.465000 ;
      RECT 1799.445000  0.085000 1799.615000 0.555000 ;
      RECT 1799.590000  1.075000 1806.540000 1.285000 ;
      RECT 1799.785000  0.255000 1800.165000 0.725000 ;
      RECT 1799.875000  1.455000 1807.245000 1.625000 ;
      RECT 1799.875000  1.625000 1800.125000 2.125000 ;
      RECT 1800.345000  1.795000 1800.595000 2.295000 ;
      RECT 1800.385000  0.085000 1800.555000 0.555000 ;
      RECT 1800.725000  0.255000 1801.105000 0.725000 ;
      RECT 1800.815000  1.625000 1801.065000 2.125000 ;
      RECT 1801.285000  1.795000 1801.535000 2.295000 ;
      RECT 1801.325000  0.085000 1801.495000 0.555000 ;
      RECT 1801.665000  0.255000 1802.045000 0.725000 ;
      RECT 1801.755000  1.625000 1802.005000 2.125000 ;
      RECT 1802.225000  1.795000 1802.475000 2.295000 ;
      RECT 1802.265000  0.085000 1802.435000 0.555000 ;
      RECT 1802.605000  0.255000 1802.985000 0.725000 ;
      RECT 1802.695000  1.625000 1802.945000 2.125000 ;
      RECT 1803.165000  1.795000 1803.415000 2.295000 ;
      RECT 1803.205000  0.085000 1803.375000 0.555000 ;
      RECT 1803.545000  0.255000 1803.925000 0.725000 ;
      RECT 1803.635000  1.625000 1803.885000 2.125000 ;
      RECT 1804.105000  1.795000 1804.355000 2.295000 ;
      RECT 1804.145000  0.085000 1804.315000 0.555000 ;
      RECT 1804.485000  0.255000 1804.865000 0.725000 ;
      RECT 1804.575000  1.625000 1804.825000 2.125000 ;
      RECT 1805.045000  1.795000 1805.295000 2.295000 ;
      RECT 1805.085000  0.085000 1805.255000 0.555000 ;
      RECT 1805.425000  0.255000 1805.805000 0.725000 ;
      RECT 1805.515000  1.625000 1805.765000 2.125000 ;
      RECT 1805.985000  1.795000 1806.235000 2.295000 ;
      RECT 1806.025000  0.085000 1806.195000 0.555000 ;
      RECT 1806.365000  0.255000 1806.745000 0.725000 ;
      RECT 1806.455000  1.625000 1806.705000 2.125000 ;
      RECT 1806.710000  0.905000 1807.245000 1.455000 ;
      RECT 1806.925000  1.795000 1807.175000 2.295000 ;
      RECT 1806.965000  0.085000 1807.235000 0.555000 ;
      RECT 1807.425000  0.085000 1807.715000 0.810000 ;
      RECT 1807.425000  1.470000 1807.715000 2.635000 ;
      RECT 1807.885000  0.085000 1809.095000 0.835000 ;
      RECT 1807.885000  0.835000 1808.405000 1.375000 ;
      RECT 1807.885000  1.545000 1809.095000 2.635000 ;
      RECT 1808.575000  1.005000 1809.095000 1.545000 ;
      RECT 1809.265000  0.085000 1809.555000 0.810000 ;
      RECT 1809.265000  1.470000 1809.555000 2.635000 ;
      RECT 1809.725000  0.085000 1811.395000 0.855000 ;
      RECT 1809.725000  0.855000 1810.475000 1.375000 ;
      RECT 1809.725000  1.545000 1811.395000 2.635000 ;
      RECT 1810.645000  1.025000 1811.395000 1.545000 ;
      RECT 1811.565000  0.085000 1811.855000 0.810000 ;
      RECT 1811.565000  1.470000 1811.855000 2.635000 ;
      RECT 1812.025000  0.085000 1814.615000 0.855000 ;
      RECT 1812.025000  0.855000 1813.235000 1.375000 ;
      RECT 1812.025000  1.545000 1814.615000 2.635000 ;
      RECT 1813.405000  1.025000 1814.615000 1.545000 ;
      RECT 1814.785000  0.085000 1815.075000 0.810000 ;
      RECT 1814.785000  1.470000 1815.075000 2.635000 ;
      RECT 1815.245000  0.085000 1818.755000 0.855000 ;
      RECT 1815.245000  0.855000 1816.895000 1.375000 ;
      RECT 1815.245000  1.545000 1818.755000 2.635000 ;
      RECT 1817.065000  1.025000 1818.755000 1.545000 ;
      RECT 1818.925000  0.085000 1819.215000 0.810000 ;
      RECT 1818.925000  1.470000 1819.215000 2.635000 ;
      RECT 1819.385000  0.085000 1824.730000 0.855000 ;
      RECT 1819.385000  0.855000 1821.965000 1.375000 ;
      RECT 1819.385000  1.545000 1824.730000 2.635000 ;
      RECT 1822.135000  1.025000 1824.730000 1.545000 ;
      RECT 1824.905000  0.085000 1825.195000 0.810000 ;
      RECT 1824.905000  1.470000 1825.195000 2.635000 ;
      RECT 1832.265000  0.085000 1832.555000 0.810000 ;
      RECT 1832.265000  1.470000 1832.555000 2.635000 ;
      RECT 1832.725000  0.085000 1833.015000 0.810000 ;
      RECT 1832.725000  1.470000 1833.015000 2.635000 ;
      RECT 1833.195000  1.495000 1833.525000 2.635000 ;
      RECT 1833.230000  0.085000 1833.490000 0.885000 ;
      RECT 1833.435000  1.055000 1833.830000 1.325000 ;
      RECT 1833.660000  0.395000 1833.935000 0.625000 ;
      RECT 1833.660000  0.625000 1833.830000 1.055000 ;
      RECT 1834.000000  0.835000 1834.390000 1.005000 ;
      RECT 1834.000000  1.005000 1834.170000 1.755000 ;
      RECT 1834.000000  1.755000 1834.395000 1.805000 ;
      RECT 1834.000000  1.805000 1834.520000 1.985000 ;
      RECT 1834.145000  0.330000 1834.390000 0.835000 ;
      RECT 1834.190000  1.985000 1834.520000 2.465000 ;
      RECT 1834.340000  1.175000 1834.730000 1.465000 ;
      RECT 1834.340000  1.465000 1835.040000 1.505000 ;
      RECT 1834.560000  0.585000 1835.000000 0.755000 ;
      RECT 1834.560000  0.755000 1834.730000 1.175000 ;
      RECT 1834.560000  1.505000 1835.040000 1.635000 ;
      RECT 1834.710000  1.635000 1835.040000 2.465000 ;
      RECT 1834.750000  0.330000 1835.000000 0.585000 ;
      RECT 1834.905000  0.945000 1835.255000 1.295000 ;
      RECT 1835.235000  0.085000 1835.565000 0.660000 ;
      RECT 1835.265000  1.465000 1835.565000 2.635000 ;
      RECT 1835.545000  0.945000 1835.895000 1.295000 ;
      RECT 1835.760000  1.465000 1836.460000 1.505000 ;
      RECT 1835.760000  1.505000 1836.240000 1.635000 ;
      RECT 1835.760000  1.635000 1836.090000 2.465000 ;
      RECT 1835.800000  0.330000 1836.050000 0.585000 ;
      RECT 1835.800000  0.585000 1836.240000 0.755000 ;
      RECT 1836.070000  0.755000 1836.240000 1.175000 ;
      RECT 1836.070000  1.175000 1836.460000 1.465000 ;
      RECT 1836.280000  1.805000 1836.800000 1.985000 ;
      RECT 1836.280000  1.985000 1836.610000 2.465000 ;
      RECT 1836.405000  1.755000 1836.800000 1.805000 ;
      RECT 1836.410000  0.330000 1836.655000 0.835000 ;
      RECT 1836.410000  0.835000 1836.800000 1.005000 ;
      RECT 1836.630000  1.005000 1836.800000 1.755000 ;
      RECT 1836.865000  0.395000 1837.140000 0.625000 ;
      RECT 1836.970000  0.625000 1837.140000 1.055000 ;
      RECT 1836.970000  1.055000 1837.365000 1.325000 ;
      RECT 1837.275000  1.495000 1837.665000 2.635000 ;
      RECT 1837.310000  0.085000 1837.630000 0.885000 ;
      RECT 1837.575000  1.055000 1837.970000 1.325000 ;
      RECT 1837.800000  0.395000 1838.075000 0.625000 ;
      RECT 1837.800000  0.625000 1837.970000 1.055000 ;
      RECT 1838.140000  0.835000 1838.530000 1.005000 ;
      RECT 1838.140000  1.005000 1838.310000 1.755000 ;
      RECT 1838.140000  1.755000 1838.535000 1.805000 ;
      RECT 1838.140000  1.805000 1838.660000 1.985000 ;
      RECT 1838.285000  0.330000 1838.530000 0.835000 ;
      RECT 1838.330000  1.985000 1838.660000 2.465000 ;
      RECT 1838.480000  1.175000 1838.870000 1.465000 ;
      RECT 1838.480000  1.465000 1839.180000 1.505000 ;
      RECT 1838.700000  0.585000 1839.140000 0.755000 ;
      RECT 1838.700000  0.755000 1838.870000 1.175000 ;
      RECT 1838.700000  1.505000 1839.180000 1.635000 ;
      RECT 1838.850000  1.635000 1839.180000 2.465000 ;
      RECT 1838.890000  0.330000 1839.140000 0.585000 ;
      RECT 1839.045000  0.945000 1839.395000 1.295000 ;
      RECT 1839.375000  0.085000 1839.705000 0.660000 ;
      RECT 1839.375000  1.465000 1839.675000 2.635000 ;
      RECT 1839.685000  0.945000 1840.035000 1.295000 ;
      RECT 1839.900000  1.465000 1840.600000 1.505000 ;
      RECT 1839.900000  1.505000 1840.380000 1.635000 ;
      RECT 1839.900000  1.635000 1840.230000 2.465000 ;
      RECT 1839.940000  0.330000 1840.190000 0.585000 ;
      RECT 1839.940000  0.585000 1840.380000 0.755000 ;
      RECT 1840.210000  0.755000 1840.380000 1.175000 ;
      RECT 1840.210000  1.175000 1840.600000 1.465000 ;
      RECT 1840.420000  1.805000 1840.940000 1.985000 ;
      RECT 1840.420000  1.985000 1840.750000 2.465000 ;
      RECT 1840.545000  1.755000 1840.940000 1.805000 ;
      RECT 1840.550000  0.330000 1840.795000 0.835000 ;
      RECT 1840.550000  0.835000 1840.940000 1.005000 ;
      RECT 1840.770000  1.005000 1840.940000 1.755000 ;
      RECT 1841.005000  0.395000 1841.280000 0.625000 ;
      RECT 1841.110000  0.625000 1841.280000 1.055000 ;
      RECT 1841.110000  1.055000 1841.505000 1.325000 ;
      RECT 1841.415000  1.495000 1841.745000 2.635000 ;
      RECT 1841.450000  0.085000 1841.710000 0.885000 ;
      RECT 1841.925000  0.085000 1842.215000 0.810000 ;
      RECT 1841.925000  1.470000 1842.215000 2.635000 ;
      RECT 1842.395000  1.055000 1843.215000 1.325000 ;
      RECT 1842.395000  1.495000 1843.585000 1.665000 ;
      RECT 1842.395000  1.665000 1842.695000 2.210000 ;
      RECT 1842.395000  2.210000 1842.725000 2.465000 ;
      RECT 1842.445000  0.255000 1842.775000 0.715000 ;
      RECT 1842.445000  0.715000 1843.635000 0.885000 ;
      RECT 1842.865000  1.835000 1843.195000 2.105000 ;
      RECT 1842.895000  2.105000 1843.195000 2.635000 ;
      RECT 1842.945000  0.085000 1843.160000 0.545000 ;
      RECT 1843.330000  0.255000 1844.475000 0.425000 ;
      RECT 1843.330000  0.425000 1843.635000 0.715000 ;
      RECT 1843.330000  0.885000 1843.635000 0.925000 ;
      RECT 1843.415000  1.665000 1843.585000 2.295000 ;
      RECT 1843.415000  2.295000 1844.580000 2.465000 ;
      RECT 1843.765000  1.755000 1844.195000 2.125000 ;
      RECT 1843.805000  0.595000 1844.135000 0.885000 ;
      RECT 1843.885000  0.885000 1844.055000 1.755000 ;
      RECT 1844.305000  0.425000 1844.475000 0.770000 ;
      RECT 1844.400000  1.205000 1844.815000 1.305000 ;
      RECT 1844.400000  1.305000 1844.920000 1.465000 ;
      RECT 1844.400000  1.465000 1845.180000 1.475000 ;
      RECT 1844.410000  1.645000 1844.580000 2.295000 ;
      RECT 1844.645000  0.585000 1845.225000 0.755000 ;
      RECT 1844.645000  0.755000 1844.815000 1.205000 ;
      RECT 1844.750000  1.475000 1845.180000 1.635000 ;
      RECT 1844.850000  1.635000 1845.180000 2.465000 ;
      RECT 1844.975000  0.330000 1845.225000 0.585000 ;
      RECT 1845.090000  1.025000 1845.425000 1.295000 ;
      RECT 1845.355000  1.465000 1845.685000 2.635000 ;
      RECT 1845.395000  0.085000 1845.645000 0.660000 ;
      RECT 1845.615000  1.025000 1845.950000 1.295000 ;
      RECT 1845.815000  0.330000 1846.065000 0.585000 ;
      RECT 1845.815000  0.585000 1846.395000 0.755000 ;
      RECT 1845.860000  1.465000 1846.640000 1.475000 ;
      RECT 1845.860000  1.475000 1846.290000 1.635000 ;
      RECT 1845.860000  1.635000 1846.190000 2.465000 ;
      RECT 1846.120000  1.305000 1846.640000 1.465000 ;
      RECT 1846.225000  0.755000 1846.395000 1.205000 ;
      RECT 1846.225000  1.205000 1846.640000 1.305000 ;
      RECT 1846.460000  1.645000 1846.630000 2.295000 ;
      RECT 1846.460000  2.295000 1847.625000 2.465000 ;
      RECT 1846.565000  0.255000 1847.710000 0.425000 ;
      RECT 1846.565000  0.425000 1846.735000 0.770000 ;
      RECT 1846.845000  1.755000 1847.275000 2.125000 ;
      RECT 1846.905000  0.595000 1847.235000 0.885000 ;
      RECT 1846.985000  0.885000 1847.155000 1.755000 ;
      RECT 1847.405000  0.425000 1847.710000 0.715000 ;
      RECT 1847.405000  0.715000 1848.595000 0.885000 ;
      RECT 1847.405000  0.885000 1847.710000 0.925000 ;
      RECT 1847.455000  1.495000 1848.645000 1.665000 ;
      RECT 1847.455000  1.665000 1847.625000 2.295000 ;
      RECT 1847.825000  1.055000 1848.645000 1.325000 ;
      RECT 1847.845000  1.835000 1848.175000 2.105000 ;
      RECT 1847.845000  2.105000 1848.145000 2.635000 ;
      RECT 1847.880000  0.085000 1848.095000 0.545000 ;
      RECT 1848.265000  0.255000 1848.595000 0.715000 ;
      RECT 1848.315000  2.210000 1848.645000 2.465000 ;
      RECT 1848.345000  1.665000 1848.645000 2.210000 ;
      RECT 1848.835000  1.055000 1849.655000 1.325000 ;
      RECT 1848.835000  1.495000 1850.025000 1.665000 ;
      RECT 1848.835000  1.665000 1849.135000 2.210000 ;
      RECT 1848.835000  2.210000 1849.165000 2.465000 ;
      RECT 1848.885000  0.255000 1849.215000 0.715000 ;
      RECT 1848.885000  0.715000 1850.075000 0.885000 ;
      RECT 1849.305000  1.835000 1849.635000 2.105000 ;
      RECT 1849.335000  2.105000 1849.635000 2.635000 ;
      RECT 1849.385000  0.085000 1849.600000 0.545000 ;
      RECT 1849.770000  0.255000 1850.915000 0.425000 ;
      RECT 1849.770000  0.425000 1850.075000 0.715000 ;
      RECT 1849.770000  0.885000 1850.075000 0.925000 ;
      RECT 1849.855000  1.665000 1850.025000 2.295000 ;
      RECT 1849.855000  2.295000 1851.020000 2.465000 ;
      RECT 1850.205000  1.755000 1850.635000 2.125000 ;
      RECT 1850.245000  0.595000 1850.575000 0.885000 ;
      RECT 1850.325000  0.885000 1850.495000 1.755000 ;
      RECT 1850.745000  0.425000 1850.915000 0.770000 ;
      RECT 1850.840000  1.205000 1851.255000 1.305000 ;
      RECT 1850.840000  1.305000 1851.360000 1.465000 ;
      RECT 1850.840000  1.465000 1851.620000 1.475000 ;
      RECT 1850.850000  1.645000 1851.020000 2.295000 ;
      RECT 1851.085000  0.585000 1851.665000 0.755000 ;
      RECT 1851.085000  0.755000 1851.255000 1.205000 ;
      RECT 1851.190000  1.475000 1851.620000 1.635000 ;
      RECT 1851.290000  1.635000 1851.620000 2.465000 ;
      RECT 1851.415000  0.330000 1851.665000 0.585000 ;
      RECT 1851.530000  1.025000 1851.865000 1.295000 ;
      RECT 1851.795000  1.465000 1852.125000 2.635000 ;
      RECT 1851.835000  0.085000 1852.085000 0.660000 ;
      RECT 1852.055000  1.025000 1852.390000 1.295000 ;
      RECT 1852.255000  0.330000 1852.505000 0.585000 ;
      RECT 1852.255000  0.585000 1852.835000 0.755000 ;
      RECT 1852.300000  1.465000 1853.080000 1.475000 ;
      RECT 1852.300000  1.475000 1852.730000 1.635000 ;
      RECT 1852.300000  1.635000 1852.630000 2.465000 ;
      RECT 1852.560000  1.305000 1853.080000 1.465000 ;
      RECT 1852.665000  0.755000 1852.835000 1.205000 ;
      RECT 1852.665000  1.205000 1853.080000 1.305000 ;
      RECT 1852.900000  1.645000 1853.070000 2.295000 ;
      RECT 1852.900000  2.295000 1854.065000 2.465000 ;
      RECT 1853.005000  0.255000 1854.150000 0.425000 ;
      RECT 1853.005000  0.425000 1853.175000 0.770000 ;
      RECT 1853.285000  1.755000 1853.715000 2.125000 ;
      RECT 1853.345000  0.595000 1853.675000 0.885000 ;
      RECT 1853.425000  0.885000 1853.595000 1.755000 ;
      RECT 1853.845000  0.425000 1854.150000 0.715000 ;
      RECT 1853.845000  0.715000 1855.035000 0.885000 ;
      RECT 1853.845000  0.885000 1854.150000 0.925000 ;
      RECT 1853.895000  1.495000 1855.085000 1.665000 ;
      RECT 1853.895000  1.665000 1854.065000 2.295000 ;
      RECT 1854.265000  1.055000 1855.085000 1.325000 ;
      RECT 1854.285000  1.835000 1854.615000 2.105000 ;
      RECT 1854.285000  2.105000 1854.585000 2.635000 ;
      RECT 1854.320000  0.085000 1854.535000 0.545000 ;
      RECT 1854.705000  0.255000 1855.035000 0.715000 ;
      RECT 1854.755000  2.210000 1855.085000 2.465000 ;
      RECT 1854.785000  1.665000 1855.085000 2.210000 ;
      RECT 1855.265000  0.085000 1855.555000 0.810000 ;
      RECT 1855.265000  1.470000 1855.555000 2.635000 ;
      RECT 1855.765000  1.495000 1856.035000 2.635000 ;
      RECT 1855.785000  0.085000 1856.035000 0.885000 ;
      RECT 1856.035000  1.055000 1857.425000 1.325000 ;
      RECT 1856.205000  0.255000 1856.535000 0.715000 ;
      RECT 1856.205000  0.715000 1858.335000 0.885000 ;
      RECT 1856.205000  1.495000 1858.435000 1.665000 ;
      RECT 1856.205000  1.665000 1856.535000 2.465000 ;
      RECT 1856.705000  0.085000 1856.975000 0.545000 ;
      RECT 1856.705000  1.835000 1856.975000 2.635000 ;
      RECT 1857.145000  0.255000 1857.475000 0.715000 ;
      RECT 1857.145000  1.665000 1857.475000 2.465000 ;
      RECT 1857.645000  0.085000 1857.895000 0.545000 ;
      RECT 1857.645000  1.835000 1857.915000 2.635000 ;
      RECT 1858.065000  0.255000 1860.095000 0.425000 ;
      RECT 1858.065000  0.425000 1858.335000 0.715000 ;
      RECT 1858.135000  1.665000 1858.435000 2.295000 ;
      RECT 1858.135000  2.295000 1860.345000 2.465000 ;
      RECT 1858.505000  0.595000 1858.835000 0.885000 ;
      RECT 1858.605000  0.885000 1858.835000 1.065000 ;
      RECT 1858.605000  1.065000 1859.875000 1.365000 ;
      RECT 1858.605000  1.365000 1858.935000 2.125000 ;
      RECT 1859.005000  0.425000 1859.175000 0.770000 ;
      RECT 1859.105000  1.535000 1859.375000 2.295000 ;
      RECT 1859.345000  0.595000 1859.675000 1.065000 ;
      RECT 1859.545000  1.365000 1859.875000 2.125000 ;
      RECT 1859.845000  0.425000 1860.095000 0.770000 ;
      RECT 1860.045000  1.065000 1861.230000 1.395000 ;
      RECT 1860.045000  1.565000 1860.345000 2.295000 ;
      RECT 1860.590000  1.605000 1860.865000 2.635000 ;
      RECT 1860.600000  0.085000 1860.890000 0.610000 ;
      RECT 1861.060000  0.280000 1861.310000 0.825000 ;
      RECT 1861.060000  0.825000 1861.230000 1.065000 ;
      RECT 1861.060000  1.395000 1861.230000 1.605000 ;
      RECT 1861.060000  1.605000 1861.390000 2.465000 ;
      RECT 1861.400000  0.995000 1861.995000 1.325000 ;
      RECT 1861.520000  0.085000 1861.810000 0.610000 ;
      RECT 1861.560000  1.605000 1861.860000 2.635000 ;
      RECT 1862.165000  0.995000 1862.760000 1.325000 ;
      RECT 1862.300000  1.605000 1862.600000 2.635000 ;
      RECT 1862.350000  0.085000 1862.640000 0.610000 ;
      RECT 1862.770000  1.605000 1863.100000 2.465000 ;
      RECT 1862.850000  0.280000 1863.100000 0.825000 ;
      RECT 1862.930000  0.825000 1863.100000 1.065000 ;
      RECT 1862.930000  1.065000 1864.115000 1.395000 ;
      RECT 1862.930000  1.395000 1863.100000 1.605000 ;
      RECT 1863.270000  0.085000 1863.560000 0.610000 ;
      RECT 1863.295000  1.605000 1863.570000 2.635000 ;
      RECT 1863.815000  1.565000 1864.115000 2.295000 ;
      RECT 1863.815000  2.295000 1866.025000 2.465000 ;
      RECT 1864.065000  0.255000 1866.095000 0.425000 ;
      RECT 1864.065000  0.425000 1864.315000 0.770000 ;
      RECT 1864.285000  1.065000 1865.555000 1.365000 ;
      RECT 1864.285000  1.365000 1864.615000 2.125000 ;
      RECT 1864.485000  0.595000 1864.815000 1.065000 ;
      RECT 1864.785000  1.535000 1865.055000 2.295000 ;
      RECT 1864.985000  0.425000 1865.155000 0.770000 ;
      RECT 1865.225000  1.365000 1865.555000 2.125000 ;
      RECT 1865.325000  0.595000 1865.655000 0.885000 ;
      RECT 1865.325000  0.885000 1865.555000 1.065000 ;
      RECT 1865.725000  1.495000 1867.955000 1.665000 ;
      RECT 1865.725000  1.665000 1866.025000 2.295000 ;
      RECT 1865.825000  0.425000 1866.095000 0.715000 ;
      RECT 1865.825000  0.715000 1867.955000 0.885000 ;
      RECT 1866.245000  1.835000 1866.515000 2.635000 ;
      RECT 1866.265000  0.085000 1866.515000 0.545000 ;
      RECT 1866.685000  0.255000 1867.015000 0.715000 ;
      RECT 1866.685000  1.665000 1867.015000 2.465000 ;
      RECT 1866.735000  1.055000 1868.125000 1.325000 ;
      RECT 1867.185000  0.085000 1867.455000 0.545000 ;
      RECT 1867.185000  1.835000 1867.455000 2.635000 ;
      RECT 1867.625000  0.255000 1867.955000 0.715000 ;
      RECT 1867.625000  1.665000 1867.955000 2.465000 ;
      RECT 1868.125000  0.085000 1868.375000 0.885000 ;
      RECT 1868.125000  1.495000 1868.395000 2.635000 ;
      RECT 1868.645000  1.495000 1868.915000 2.635000 ;
      RECT 1868.665000  0.085000 1868.915000 0.885000 ;
      RECT 1868.915000  1.055000 1870.305000 1.325000 ;
      RECT 1869.085000  0.255000 1869.415000 0.715000 ;
      RECT 1869.085000  0.715000 1871.215000 0.885000 ;
      RECT 1869.085000  1.495000 1871.315000 1.665000 ;
      RECT 1869.085000  1.665000 1869.415000 2.465000 ;
      RECT 1869.585000  0.085000 1869.855000 0.545000 ;
      RECT 1869.585000  1.835000 1869.855000 2.635000 ;
      RECT 1870.025000  0.255000 1870.355000 0.715000 ;
      RECT 1870.025000  1.665000 1870.355000 2.465000 ;
      RECT 1870.525000  0.085000 1870.775000 0.545000 ;
      RECT 1870.525000  1.835000 1870.795000 2.635000 ;
      RECT 1870.945000  0.255000 1872.975000 0.425000 ;
      RECT 1870.945000  0.425000 1871.215000 0.715000 ;
      RECT 1871.015000  1.665000 1871.315000 2.295000 ;
      RECT 1871.015000  2.295000 1873.225000 2.465000 ;
      RECT 1871.385000  0.595000 1871.715000 0.885000 ;
      RECT 1871.485000  0.885000 1871.715000 1.065000 ;
      RECT 1871.485000  1.065000 1872.755000 1.365000 ;
      RECT 1871.485000  1.365000 1871.815000 2.125000 ;
      RECT 1871.885000  0.425000 1872.055000 0.770000 ;
      RECT 1871.985000  1.535000 1872.255000 2.295000 ;
      RECT 1872.225000  0.595000 1872.555000 1.065000 ;
      RECT 1872.425000  1.365000 1872.755000 2.125000 ;
      RECT 1872.725000  0.425000 1872.975000 0.770000 ;
      RECT 1872.925000  1.065000 1874.110000 1.395000 ;
      RECT 1872.925000  1.565000 1873.225000 2.295000 ;
      RECT 1873.470000  1.605000 1873.745000 2.635000 ;
      RECT 1873.480000  0.085000 1873.770000 0.610000 ;
      RECT 1873.940000  0.280000 1874.190000 0.825000 ;
      RECT 1873.940000  0.825000 1874.110000 1.065000 ;
      RECT 1873.940000  1.395000 1874.110000 1.605000 ;
      RECT 1873.940000  1.605000 1874.270000 2.465000 ;
      RECT 1874.280000  0.995000 1874.875000 1.325000 ;
      RECT 1874.400000  0.085000 1874.690000 0.610000 ;
      RECT 1874.440000  1.605000 1874.740000 2.635000 ;
      RECT 1875.045000  0.995000 1875.640000 1.325000 ;
      RECT 1875.180000  1.605000 1875.480000 2.635000 ;
      RECT 1875.230000  0.085000 1875.520000 0.610000 ;
      RECT 1875.650000  1.605000 1875.980000 2.465000 ;
      RECT 1875.730000  0.280000 1875.980000 0.825000 ;
      RECT 1875.810000  0.825000 1875.980000 1.065000 ;
      RECT 1875.810000  1.065000 1876.995000 1.395000 ;
      RECT 1875.810000  1.395000 1875.980000 1.605000 ;
      RECT 1876.150000  0.085000 1876.440000 0.610000 ;
      RECT 1876.175000  1.605000 1876.450000 2.635000 ;
      RECT 1876.695000  1.565000 1876.995000 2.295000 ;
      RECT 1876.695000  2.295000 1878.905000 2.465000 ;
      RECT 1876.945000  0.255000 1878.975000 0.425000 ;
      RECT 1876.945000  0.425000 1877.195000 0.770000 ;
      RECT 1877.165000  1.065000 1878.435000 1.365000 ;
      RECT 1877.165000  1.365000 1877.495000 2.125000 ;
      RECT 1877.365000  0.595000 1877.695000 1.065000 ;
      RECT 1877.665000  1.535000 1877.935000 2.295000 ;
      RECT 1877.865000  0.425000 1878.035000 0.770000 ;
      RECT 1878.105000  1.365000 1878.435000 2.125000 ;
      RECT 1878.205000  0.595000 1878.535000 0.885000 ;
      RECT 1878.205000  0.885000 1878.435000 1.065000 ;
      RECT 1878.605000  1.495000 1880.835000 1.665000 ;
      RECT 1878.605000  1.665000 1878.905000 2.295000 ;
      RECT 1878.705000  0.425000 1878.975000 0.715000 ;
      RECT 1878.705000  0.715000 1880.835000 0.885000 ;
      RECT 1879.125000  1.835000 1879.395000 2.635000 ;
      RECT 1879.145000  0.085000 1879.395000 0.545000 ;
      RECT 1879.565000  0.255000 1879.895000 0.715000 ;
      RECT 1879.565000  1.665000 1879.895000 2.465000 ;
      RECT 1879.615000  1.055000 1881.005000 1.325000 ;
      RECT 1880.065000  0.085000 1880.335000 0.545000 ;
      RECT 1880.065000  1.835000 1880.335000 2.635000 ;
      RECT 1880.505000  0.255000 1880.835000 0.715000 ;
      RECT 1880.505000  1.665000 1880.835000 2.465000 ;
      RECT 1881.005000  0.085000 1881.255000 0.885000 ;
      RECT 1881.005000  1.495000 1881.275000 2.635000 ;
      RECT 1881.485000  0.085000 1881.775000 0.810000 ;
      RECT 1881.485000  1.470000 1881.775000 2.635000 ;
      RECT 1881.955000  1.495000 1882.285000 2.635000 ;
      RECT 1881.990000  0.085000 1882.250000 0.885000 ;
      RECT 1882.195000  1.055000 1882.590000 1.325000 ;
      RECT 1882.420000  0.395000 1882.695000 0.625000 ;
      RECT 1882.420000  0.625000 1882.590000 1.055000 ;
      RECT 1882.760000  0.835000 1883.150000 1.005000 ;
      RECT 1882.760000  1.005000 1882.930000 1.755000 ;
      RECT 1882.760000  1.755000 1883.155000 1.805000 ;
      RECT 1882.760000  1.805000 1883.280000 1.985000 ;
      RECT 1882.905000  0.330000 1883.150000 0.835000 ;
      RECT 1882.950000  1.985000 1883.280000 2.465000 ;
      RECT 1883.100000  1.175000 1883.490000 1.465000 ;
      RECT 1883.100000  1.465000 1883.800000 1.505000 ;
      RECT 1883.320000  0.585000 1883.760000 0.755000 ;
      RECT 1883.320000  0.755000 1883.490000 1.175000 ;
      RECT 1883.320000  1.505000 1883.800000 1.635000 ;
      RECT 1883.470000  1.635000 1883.800000 2.465000 ;
      RECT 1883.510000  0.330000 1883.760000 0.585000 ;
      RECT 1883.665000  0.945000 1884.065000 1.295000 ;
      RECT 1883.995000  0.085000 1884.325000 0.660000 ;
      RECT 1883.995000  1.465000 1884.325000 2.635000 ;
      RECT 1884.255000  0.945000 1884.655000 1.295000 ;
      RECT 1884.520000  1.465000 1885.220000 1.505000 ;
      RECT 1884.520000  1.505000 1885.000000 1.635000 ;
      RECT 1884.520000  1.635000 1884.850000 2.465000 ;
      RECT 1884.560000  0.330000 1884.810000 0.585000 ;
      RECT 1884.560000  0.585000 1885.000000 0.755000 ;
      RECT 1884.830000  0.755000 1885.000000 1.175000 ;
      RECT 1884.830000  1.175000 1885.220000 1.465000 ;
      RECT 1885.040000  1.805000 1885.560000 1.985000 ;
      RECT 1885.040000  1.985000 1885.370000 2.465000 ;
      RECT 1885.165000  1.755000 1885.560000 1.805000 ;
      RECT 1885.170000  0.330000 1885.415000 0.835000 ;
      RECT 1885.170000  0.835000 1885.560000 1.005000 ;
      RECT 1885.390000  1.005000 1885.560000 1.755000 ;
      RECT 1885.625000  0.395000 1885.900000 0.625000 ;
      RECT 1885.730000  0.625000 1885.900000 1.055000 ;
      RECT 1885.730000  1.055000 1886.125000 1.325000 ;
      RECT 1886.035000  1.495000 1886.425000 2.635000 ;
      RECT 1886.070000  0.085000 1886.390000 0.885000 ;
      RECT 1886.335000  1.055000 1886.730000 1.325000 ;
      RECT 1886.560000  0.395000 1886.835000 0.625000 ;
      RECT 1886.560000  0.625000 1886.730000 1.055000 ;
      RECT 1886.900000  0.835000 1887.290000 1.005000 ;
      RECT 1886.900000  1.005000 1887.070000 1.755000 ;
      RECT 1886.900000  1.755000 1887.295000 1.805000 ;
      RECT 1886.900000  1.805000 1887.420000 1.985000 ;
      RECT 1887.045000  0.330000 1887.290000 0.835000 ;
      RECT 1887.090000  1.985000 1887.420000 2.465000 ;
      RECT 1887.240000  1.175000 1887.630000 1.465000 ;
      RECT 1887.240000  1.465000 1887.940000 1.505000 ;
      RECT 1887.460000  0.585000 1887.900000 0.755000 ;
      RECT 1887.460000  0.755000 1887.630000 1.175000 ;
      RECT 1887.460000  1.505000 1887.940000 1.635000 ;
      RECT 1887.610000  1.635000 1887.940000 2.465000 ;
      RECT 1887.650000  0.330000 1887.900000 0.585000 ;
      RECT 1887.805000  0.945000 1888.205000 1.295000 ;
      RECT 1888.135000  0.085000 1888.465000 0.660000 ;
      RECT 1888.135000  1.465000 1888.465000 2.635000 ;
      RECT 1888.395000  0.945000 1888.795000 1.295000 ;
      RECT 1888.660000  1.465000 1889.360000 1.505000 ;
      RECT 1888.660000  1.505000 1889.140000 1.635000 ;
      RECT 1888.660000  1.635000 1888.990000 2.465000 ;
      RECT 1888.700000  0.330000 1888.950000 0.585000 ;
      RECT 1888.700000  0.585000 1889.140000 0.755000 ;
      RECT 1888.970000  0.755000 1889.140000 1.175000 ;
      RECT 1888.970000  1.175000 1889.360000 1.465000 ;
      RECT 1889.180000  1.805000 1889.700000 1.985000 ;
      RECT 1889.180000  1.985000 1889.510000 2.465000 ;
      RECT 1889.305000  1.755000 1889.700000 1.805000 ;
      RECT 1889.310000  0.330000 1889.555000 0.835000 ;
      RECT 1889.310000  0.835000 1889.700000 1.005000 ;
      RECT 1889.530000  1.005000 1889.700000 1.755000 ;
      RECT 1889.765000  0.395000 1890.040000 0.625000 ;
      RECT 1889.870000  0.625000 1890.040000 1.055000 ;
      RECT 1889.870000  1.055000 1890.265000 1.325000 ;
      RECT 1890.175000  1.495000 1890.565000 2.635000 ;
      RECT 1890.210000  0.085000 1890.530000 0.885000 ;
      RECT 1890.475000  1.055000 1890.870000 1.325000 ;
      RECT 1890.700000  0.395000 1890.975000 0.625000 ;
      RECT 1890.700000  0.625000 1890.870000 1.055000 ;
      RECT 1891.040000  0.835000 1891.430000 1.005000 ;
      RECT 1891.040000  1.005000 1891.210000 1.755000 ;
      RECT 1891.040000  1.755000 1891.435000 1.805000 ;
      RECT 1891.040000  1.805000 1891.560000 1.985000 ;
      RECT 1891.185000  0.330000 1891.430000 0.835000 ;
      RECT 1891.230000  1.985000 1891.560000 2.465000 ;
      RECT 1891.380000  1.175000 1891.770000 1.465000 ;
      RECT 1891.380000  1.465000 1892.080000 1.505000 ;
      RECT 1891.600000  0.585000 1892.040000 0.755000 ;
      RECT 1891.600000  0.755000 1891.770000 1.175000 ;
      RECT 1891.600000  1.505000 1892.080000 1.635000 ;
      RECT 1891.750000  1.635000 1892.080000 2.465000 ;
      RECT 1891.790000  0.330000 1892.040000 0.585000 ;
      RECT 1891.945000  0.945000 1892.345000 1.295000 ;
      RECT 1892.275000  0.085000 1892.605000 0.660000 ;
      RECT 1892.275000  1.465000 1892.605000 2.635000 ;
      RECT 1892.535000  0.945000 1892.935000 1.295000 ;
      RECT 1892.800000  1.465000 1893.500000 1.505000 ;
      RECT 1892.800000  1.505000 1893.280000 1.635000 ;
      RECT 1892.800000  1.635000 1893.130000 2.465000 ;
      RECT 1892.840000  0.330000 1893.090000 0.585000 ;
      RECT 1892.840000  0.585000 1893.280000 0.755000 ;
      RECT 1893.110000  0.755000 1893.280000 1.175000 ;
      RECT 1893.110000  1.175000 1893.500000 1.465000 ;
      RECT 1893.320000  1.805000 1893.840000 1.985000 ;
      RECT 1893.320000  1.985000 1893.650000 2.465000 ;
      RECT 1893.445000  1.755000 1893.840000 1.805000 ;
      RECT 1893.450000  0.330000 1893.695000 0.835000 ;
      RECT 1893.450000  0.835000 1893.840000 1.005000 ;
      RECT 1893.670000  1.005000 1893.840000 1.755000 ;
      RECT 1893.905000  0.395000 1894.180000 0.625000 ;
      RECT 1894.010000  0.625000 1894.180000 1.055000 ;
      RECT 1894.010000  1.055000 1894.405000 1.325000 ;
      RECT 1894.315000  1.495000 1894.705000 2.635000 ;
      RECT 1894.350000  0.085000 1894.670000 0.885000 ;
      RECT 1894.615000  1.055000 1895.010000 1.325000 ;
      RECT 1894.840000  0.395000 1895.115000 0.625000 ;
      RECT 1894.840000  0.625000 1895.010000 1.055000 ;
      RECT 1895.180000  0.835000 1895.570000 1.005000 ;
      RECT 1895.180000  1.005000 1895.350000 1.755000 ;
      RECT 1895.180000  1.755000 1895.575000 1.805000 ;
      RECT 1895.180000  1.805000 1895.700000 1.985000 ;
      RECT 1895.325000  0.330000 1895.570000 0.835000 ;
      RECT 1895.370000  1.985000 1895.700000 2.465000 ;
      RECT 1895.520000  1.175000 1895.910000 1.465000 ;
      RECT 1895.520000  1.465000 1896.220000 1.505000 ;
      RECT 1895.740000  0.585000 1896.180000 0.755000 ;
      RECT 1895.740000  0.755000 1895.910000 1.175000 ;
      RECT 1895.740000  1.505000 1896.220000 1.635000 ;
      RECT 1895.890000  1.635000 1896.220000 2.465000 ;
      RECT 1895.930000  0.330000 1896.180000 0.585000 ;
      RECT 1896.085000  0.945000 1896.485000 1.295000 ;
      RECT 1896.415000  0.085000 1896.745000 0.660000 ;
      RECT 1896.415000  1.465000 1896.745000 2.635000 ;
      RECT 1896.675000  0.945000 1897.075000 1.295000 ;
      RECT 1896.940000  1.465000 1897.640000 1.505000 ;
      RECT 1896.940000  1.505000 1897.420000 1.635000 ;
      RECT 1896.940000  1.635000 1897.270000 2.465000 ;
      RECT 1896.980000  0.330000 1897.230000 0.585000 ;
      RECT 1896.980000  0.585000 1897.420000 0.755000 ;
      RECT 1897.250000  0.755000 1897.420000 1.175000 ;
      RECT 1897.250000  1.175000 1897.640000 1.465000 ;
      RECT 1897.460000  1.805000 1897.980000 1.985000 ;
      RECT 1897.460000  1.985000 1897.790000 2.465000 ;
      RECT 1897.585000  1.755000 1897.980000 1.805000 ;
      RECT 1897.590000  0.330000 1897.835000 0.835000 ;
      RECT 1897.590000  0.835000 1897.980000 1.005000 ;
      RECT 1897.810000  1.005000 1897.980000 1.755000 ;
      RECT 1898.045000  0.395000 1898.320000 0.625000 ;
      RECT 1898.150000  0.625000 1898.320000 1.055000 ;
      RECT 1898.150000  1.055000 1898.545000 1.325000 ;
      RECT 1898.455000  1.495000 1898.785000 2.635000 ;
      RECT 1898.490000  0.085000 1898.750000 0.885000 ;
      RECT 1898.965000  0.085000 1899.255000 0.810000 ;
      RECT 1898.965000  1.470000 1899.255000 2.635000 ;
      RECT 1899.435000  1.055000 1900.255000 1.325000 ;
      RECT 1899.435000  1.495000 1900.625000 1.665000 ;
      RECT 1899.435000  1.665000 1899.735000 2.210000 ;
      RECT 1899.435000  2.210000 1899.765000 2.465000 ;
      RECT 1899.485000  0.255000 1899.815000 0.715000 ;
      RECT 1899.485000  0.715000 1900.675000 0.885000 ;
      RECT 1899.905000  1.835000 1900.235000 2.105000 ;
      RECT 1899.935000  2.105000 1900.235000 2.635000 ;
      RECT 1899.985000  0.085000 1900.200000 0.545000 ;
      RECT 1900.370000  0.255000 1901.515000 0.425000 ;
      RECT 1900.370000  0.425000 1900.675000 0.715000 ;
      RECT 1900.370000  0.885000 1900.675000 0.925000 ;
      RECT 1900.455000  1.665000 1900.625000 2.295000 ;
      RECT 1900.455000  2.295000 1901.620000 2.465000 ;
      RECT 1900.805000  1.755000 1901.235000 2.125000 ;
      RECT 1900.845000  0.595000 1901.175000 0.885000 ;
      RECT 1900.925000  0.885000 1901.095000 1.755000 ;
      RECT 1901.345000  0.425000 1901.515000 0.770000 ;
      RECT 1901.440000  1.205000 1901.855000 1.305000 ;
      RECT 1901.440000  1.305000 1901.960000 1.465000 ;
      RECT 1901.440000  1.465000 1902.220000 1.475000 ;
      RECT 1901.450000  1.645000 1901.620000 2.295000 ;
      RECT 1901.685000  0.585000 1902.265000 0.755000 ;
      RECT 1901.685000  0.755000 1901.855000 1.205000 ;
      RECT 1901.790000  1.475000 1902.220000 1.635000 ;
      RECT 1901.890000  1.635000 1902.220000 2.465000 ;
      RECT 1902.015000  0.330000 1902.265000 0.585000 ;
      RECT 1902.130000  1.025000 1902.465000 1.295000 ;
      RECT 1902.395000  1.465000 1902.725000 2.635000 ;
      RECT 1902.435000  0.085000 1902.685000 0.660000 ;
      RECT 1902.655000  1.025000 1902.990000 1.295000 ;
      RECT 1902.855000  0.330000 1903.105000 0.585000 ;
      RECT 1902.855000  0.585000 1903.435000 0.755000 ;
      RECT 1902.900000  1.465000 1903.680000 1.475000 ;
      RECT 1902.900000  1.475000 1903.330000 1.635000 ;
      RECT 1902.900000  1.635000 1903.230000 2.465000 ;
      RECT 1903.160000  1.305000 1903.680000 1.465000 ;
      RECT 1903.265000  0.755000 1903.435000 1.205000 ;
      RECT 1903.265000  1.205000 1903.680000 1.305000 ;
      RECT 1903.500000  1.645000 1903.670000 2.295000 ;
      RECT 1903.500000  2.295000 1904.665000 2.465000 ;
      RECT 1903.605000  0.255000 1904.750000 0.425000 ;
      RECT 1903.605000  0.425000 1903.775000 0.770000 ;
      RECT 1903.885000  1.755000 1904.315000 2.125000 ;
      RECT 1903.945000  0.595000 1904.275000 0.885000 ;
      RECT 1904.025000  0.885000 1904.195000 1.755000 ;
      RECT 1904.445000  0.425000 1904.750000 0.715000 ;
      RECT 1904.445000  0.715000 1905.635000 0.885000 ;
      RECT 1904.445000  0.885000 1904.750000 0.925000 ;
      RECT 1904.495000  1.495000 1905.685000 1.665000 ;
      RECT 1904.495000  1.665000 1904.665000 2.295000 ;
      RECT 1904.865000  1.055000 1905.685000 1.325000 ;
      RECT 1904.885000  1.835000 1905.215000 2.105000 ;
      RECT 1904.885000  2.105000 1905.185000 2.635000 ;
      RECT 1904.920000  0.085000 1905.135000 0.545000 ;
      RECT 1905.305000  0.255000 1905.635000 0.715000 ;
      RECT 1905.355000  2.210000 1905.685000 2.465000 ;
      RECT 1905.385000  1.665000 1905.685000 2.210000 ;
      RECT 1905.875000  1.055000 1906.695000 1.325000 ;
      RECT 1905.875000  1.495000 1907.065000 1.665000 ;
      RECT 1905.875000  1.665000 1906.175000 2.210000 ;
      RECT 1905.875000  2.210000 1906.205000 2.465000 ;
      RECT 1905.925000  0.255000 1906.255000 0.715000 ;
      RECT 1905.925000  0.715000 1907.115000 0.885000 ;
      RECT 1906.345000  1.835000 1906.675000 2.105000 ;
      RECT 1906.375000  2.105000 1906.675000 2.635000 ;
      RECT 1906.425000  0.085000 1906.640000 0.545000 ;
      RECT 1906.810000  0.255000 1907.955000 0.425000 ;
      RECT 1906.810000  0.425000 1907.115000 0.715000 ;
      RECT 1906.810000  0.885000 1907.115000 0.925000 ;
      RECT 1906.895000  1.665000 1907.065000 2.295000 ;
      RECT 1906.895000  2.295000 1908.060000 2.465000 ;
      RECT 1907.245000  1.755000 1907.675000 2.125000 ;
      RECT 1907.285000  0.595000 1907.615000 0.885000 ;
      RECT 1907.365000  0.885000 1907.535000 1.755000 ;
      RECT 1907.785000  0.425000 1907.955000 0.770000 ;
      RECT 1907.880000  1.205000 1908.295000 1.305000 ;
      RECT 1907.880000  1.305000 1908.400000 1.465000 ;
      RECT 1907.880000  1.465000 1908.660000 1.475000 ;
      RECT 1907.890000  1.645000 1908.060000 2.295000 ;
      RECT 1908.125000  0.585000 1908.705000 0.755000 ;
      RECT 1908.125000  0.755000 1908.295000 1.205000 ;
      RECT 1908.230000  1.475000 1908.660000 1.635000 ;
      RECT 1908.330000  1.635000 1908.660000 2.465000 ;
      RECT 1908.455000  0.330000 1908.705000 0.585000 ;
      RECT 1908.570000  1.025000 1908.905000 1.295000 ;
      RECT 1908.835000  1.465000 1909.165000 2.635000 ;
      RECT 1908.875000  0.085000 1909.125000 0.660000 ;
      RECT 1909.095000  1.025000 1909.430000 1.295000 ;
      RECT 1909.295000  0.330000 1909.545000 0.585000 ;
      RECT 1909.295000  0.585000 1909.875000 0.755000 ;
      RECT 1909.340000  1.465000 1910.120000 1.475000 ;
      RECT 1909.340000  1.475000 1909.770000 1.635000 ;
      RECT 1909.340000  1.635000 1909.670000 2.465000 ;
      RECT 1909.600000  1.305000 1910.120000 1.465000 ;
      RECT 1909.705000  0.755000 1909.875000 1.205000 ;
      RECT 1909.705000  1.205000 1910.120000 1.305000 ;
      RECT 1909.940000  1.645000 1910.110000 2.295000 ;
      RECT 1909.940000  2.295000 1911.105000 2.465000 ;
      RECT 1910.045000  0.255000 1911.190000 0.425000 ;
      RECT 1910.045000  0.425000 1910.215000 0.770000 ;
      RECT 1910.325000  1.755000 1910.755000 2.125000 ;
      RECT 1910.385000  0.595000 1910.715000 0.885000 ;
      RECT 1910.465000  0.885000 1910.635000 1.755000 ;
      RECT 1910.885000  0.425000 1911.190000 0.715000 ;
      RECT 1910.885000  0.715000 1912.075000 0.885000 ;
      RECT 1910.885000  0.885000 1911.190000 0.925000 ;
      RECT 1910.935000  1.495000 1912.125000 1.665000 ;
      RECT 1910.935000  1.665000 1911.105000 2.295000 ;
      RECT 1911.305000  1.055000 1912.125000 1.325000 ;
      RECT 1911.325000  1.835000 1911.655000 2.105000 ;
      RECT 1911.325000  2.105000 1911.625000 2.635000 ;
      RECT 1911.360000  0.085000 1911.575000 0.545000 ;
      RECT 1911.745000  0.255000 1912.075000 0.715000 ;
      RECT 1911.795000  2.210000 1912.125000 2.465000 ;
      RECT 1911.825000  1.665000 1912.125000 2.210000 ;
      RECT 1912.315000  1.055000 1913.135000 1.325000 ;
      RECT 1912.315000  1.495000 1913.505000 1.665000 ;
      RECT 1912.315000  1.665000 1912.615000 2.210000 ;
      RECT 1912.315000  2.210000 1912.645000 2.465000 ;
      RECT 1912.365000  0.255000 1912.695000 0.715000 ;
      RECT 1912.365000  0.715000 1913.555000 0.885000 ;
      RECT 1912.785000  1.835000 1913.115000 2.105000 ;
      RECT 1912.815000  2.105000 1913.115000 2.635000 ;
      RECT 1912.865000  0.085000 1913.080000 0.545000 ;
      RECT 1913.250000  0.255000 1914.395000 0.425000 ;
      RECT 1913.250000  0.425000 1913.555000 0.715000 ;
      RECT 1913.250000  0.885000 1913.555000 0.925000 ;
      RECT 1913.335000  1.665000 1913.505000 2.295000 ;
      RECT 1913.335000  2.295000 1914.500000 2.465000 ;
      RECT 1913.685000  1.755000 1914.115000 2.125000 ;
      RECT 1913.725000  0.595000 1914.055000 0.885000 ;
      RECT 1913.805000  0.885000 1913.975000 1.755000 ;
      RECT 1914.225000  0.425000 1914.395000 0.770000 ;
      RECT 1914.320000  1.205000 1914.735000 1.305000 ;
      RECT 1914.320000  1.305000 1914.840000 1.465000 ;
      RECT 1914.320000  1.465000 1915.100000 1.475000 ;
      RECT 1914.330000  1.645000 1914.500000 2.295000 ;
      RECT 1914.565000  0.585000 1915.145000 0.755000 ;
      RECT 1914.565000  0.755000 1914.735000 1.205000 ;
      RECT 1914.670000  1.475000 1915.100000 1.635000 ;
      RECT 1914.770000  1.635000 1915.100000 2.465000 ;
      RECT 1914.895000  0.330000 1915.145000 0.585000 ;
      RECT 1915.010000  1.025000 1915.345000 1.295000 ;
      RECT 1915.275000  1.465000 1915.605000 2.635000 ;
      RECT 1915.315000  0.085000 1915.565000 0.660000 ;
      RECT 1915.535000  1.025000 1915.870000 1.295000 ;
      RECT 1915.735000  0.330000 1915.985000 0.585000 ;
      RECT 1915.735000  0.585000 1916.315000 0.755000 ;
      RECT 1915.780000  1.465000 1916.560000 1.475000 ;
      RECT 1915.780000  1.475000 1916.210000 1.635000 ;
      RECT 1915.780000  1.635000 1916.110000 2.465000 ;
      RECT 1916.040000  1.305000 1916.560000 1.465000 ;
      RECT 1916.145000  0.755000 1916.315000 1.205000 ;
      RECT 1916.145000  1.205000 1916.560000 1.305000 ;
      RECT 1916.380000  1.645000 1916.550000 2.295000 ;
      RECT 1916.380000  2.295000 1917.545000 2.465000 ;
      RECT 1916.485000  0.255000 1917.630000 0.425000 ;
      RECT 1916.485000  0.425000 1916.655000 0.770000 ;
      RECT 1916.765000  1.755000 1917.195000 2.125000 ;
      RECT 1916.825000  0.595000 1917.155000 0.885000 ;
      RECT 1916.905000  0.885000 1917.075000 1.755000 ;
      RECT 1917.325000  0.425000 1917.630000 0.715000 ;
      RECT 1917.325000  0.715000 1918.515000 0.885000 ;
      RECT 1917.325000  0.885000 1917.630000 0.925000 ;
      RECT 1917.375000  1.495000 1918.565000 1.665000 ;
      RECT 1917.375000  1.665000 1917.545000 2.295000 ;
      RECT 1917.745000  1.055000 1918.565000 1.325000 ;
      RECT 1917.765000  1.835000 1918.095000 2.105000 ;
      RECT 1917.765000  2.105000 1918.065000 2.635000 ;
      RECT 1917.800000  0.085000 1918.015000 0.545000 ;
      RECT 1918.185000  0.255000 1918.515000 0.715000 ;
      RECT 1918.235000  2.210000 1918.565000 2.465000 ;
      RECT 1918.265000  1.665000 1918.565000 2.210000 ;
      RECT 1918.755000  1.055000 1919.575000 1.325000 ;
      RECT 1918.755000  1.495000 1919.945000 1.665000 ;
      RECT 1918.755000  1.665000 1919.055000 2.210000 ;
      RECT 1918.755000  2.210000 1919.085000 2.465000 ;
      RECT 1918.805000  0.255000 1919.135000 0.715000 ;
      RECT 1918.805000  0.715000 1919.995000 0.885000 ;
      RECT 1919.225000  1.835000 1919.555000 2.105000 ;
      RECT 1919.255000  2.105000 1919.555000 2.635000 ;
      RECT 1919.305000  0.085000 1919.520000 0.545000 ;
      RECT 1919.690000  0.255000 1920.835000 0.425000 ;
      RECT 1919.690000  0.425000 1919.995000 0.715000 ;
      RECT 1919.690000  0.885000 1919.995000 0.925000 ;
      RECT 1919.775000  1.665000 1919.945000 2.295000 ;
      RECT 1919.775000  2.295000 1920.940000 2.465000 ;
      RECT 1920.125000  1.755000 1920.555000 2.125000 ;
      RECT 1920.165000  0.595000 1920.495000 0.885000 ;
      RECT 1920.245000  0.885000 1920.415000 1.755000 ;
      RECT 1920.665000  0.425000 1920.835000 0.770000 ;
      RECT 1920.760000  1.205000 1921.175000 1.305000 ;
      RECT 1920.760000  1.305000 1921.280000 1.465000 ;
      RECT 1920.760000  1.465000 1921.540000 1.475000 ;
      RECT 1920.770000  1.645000 1920.940000 2.295000 ;
      RECT 1921.005000  0.585000 1921.585000 0.755000 ;
      RECT 1921.005000  0.755000 1921.175000 1.205000 ;
      RECT 1921.110000  1.475000 1921.540000 1.635000 ;
      RECT 1921.210000  1.635000 1921.540000 2.465000 ;
      RECT 1921.335000  0.330000 1921.585000 0.585000 ;
      RECT 1921.450000  1.025000 1921.785000 1.295000 ;
      RECT 1921.715000  1.465000 1922.045000 2.635000 ;
      RECT 1921.755000  0.085000 1922.005000 0.660000 ;
      RECT 1921.975000  1.025000 1922.310000 1.295000 ;
      RECT 1922.175000  0.330000 1922.425000 0.585000 ;
      RECT 1922.175000  0.585000 1922.755000 0.755000 ;
      RECT 1922.220000  1.465000 1923.000000 1.475000 ;
      RECT 1922.220000  1.475000 1922.650000 1.635000 ;
      RECT 1922.220000  1.635000 1922.550000 2.465000 ;
      RECT 1922.480000  1.305000 1923.000000 1.465000 ;
      RECT 1922.585000  0.755000 1922.755000 1.205000 ;
      RECT 1922.585000  1.205000 1923.000000 1.305000 ;
      RECT 1922.820000  1.645000 1922.990000 2.295000 ;
      RECT 1922.820000  2.295000 1923.985000 2.465000 ;
      RECT 1922.925000  0.255000 1924.070000 0.425000 ;
      RECT 1922.925000  0.425000 1923.095000 0.770000 ;
      RECT 1923.205000  1.755000 1923.635000 2.125000 ;
      RECT 1923.265000  0.595000 1923.595000 0.885000 ;
      RECT 1923.345000  0.885000 1923.515000 1.755000 ;
      RECT 1923.765000  0.425000 1924.070000 0.715000 ;
      RECT 1923.765000  0.715000 1924.955000 0.885000 ;
      RECT 1923.765000  0.885000 1924.070000 0.925000 ;
      RECT 1923.815000  1.495000 1925.005000 1.665000 ;
      RECT 1923.815000  1.665000 1923.985000 2.295000 ;
      RECT 1924.185000  1.055000 1925.005000 1.325000 ;
      RECT 1924.205000  1.835000 1924.535000 2.105000 ;
      RECT 1924.205000  2.105000 1924.505000 2.635000 ;
      RECT 1924.240000  0.085000 1924.455000 0.545000 ;
      RECT 1924.625000  0.255000 1924.955000 0.715000 ;
      RECT 1924.675000  2.210000 1925.005000 2.465000 ;
      RECT 1924.705000  1.665000 1925.005000 2.210000 ;
      RECT 1925.185000  0.085000 1925.475000 0.810000 ;
      RECT 1925.185000  1.470000 1925.475000 2.635000 ;
      RECT 1925.650000  0.255000 1925.905000 1.495000 ;
      RECT 1925.650000  1.495000 1925.985000 2.465000 ;
      RECT 1926.075000  0.085000 1926.455000 0.485000 ;
      RECT 1926.075000  0.655000 1927.170000 0.825000 ;
      RECT 1926.075000  0.825000 1926.245000 1.325000 ;
      RECT 1926.205000  1.495000 1926.375000 2.635000 ;
      RECT 1926.555000  0.995000 1926.830000 1.325000 ;
      RECT 1926.630000  1.325000 1926.830000 2.295000 ;
      RECT 1926.630000  2.295000 1928.975000 2.465000 ;
      RECT 1926.995000  0.255000 1927.515000 0.620000 ;
      RECT 1926.995000  0.620000 1927.170000 0.655000 ;
      RECT 1927.000000  0.825000 1927.170000 1.955000 ;
      RECT 1927.000000  1.955000 1928.445000 2.125000 ;
      RECT 1927.340000  0.810000 1927.510000 1.615000 ;
      RECT 1927.340000  1.615000 1928.635000 1.785000 ;
      RECT 1927.850000  0.255000 1928.175000 1.415000 ;
      RECT 1928.345000  0.255000 1928.635000 1.615000 ;
      RECT 1928.805000  1.440000 1929.555000 1.630000 ;
      RECT 1928.805000  1.630000 1928.975000 2.295000 ;
      RECT 1928.810000  0.085000 1929.325000 0.525000 ;
      RECT 1928.885000  0.695000 1929.945000 0.865000 ;
      RECT 1928.885000  0.865000 1929.055000 1.185000 ;
      RECT 1929.145000  1.835000 1929.375000 2.635000 ;
      RECT 1929.365000  1.055000 1929.555000 1.440000 ;
      RECT 1929.545000  1.835000 1929.945000 2.465000 ;
      RECT 1929.595000  0.255000 1929.840000 0.695000 ;
      RECT 1929.775000  0.865000 1929.945000 1.835000 ;
      RECT 1930.245000  0.085000 1930.535000 0.810000 ;
      RECT 1930.245000  1.470000 1930.535000 2.635000 ;
      RECT 1930.755000  0.085000 1931.005000 0.655000 ;
      RECT 1930.755000  1.495000 1931.000000 2.635000 ;
      RECT 1931.175000  0.255000 1931.425000 1.495000 ;
      RECT 1931.175000  1.495000 1931.515000 2.465000 ;
      RECT 1931.595000  0.085000 1931.975000 0.485000 ;
      RECT 1931.595000  0.655000 1932.690000 0.825000 ;
      RECT 1931.595000  0.825000 1931.765000 1.325000 ;
      RECT 1931.695000  1.495000 1931.945000 2.635000 ;
      RECT 1932.075000  0.995000 1932.350000 1.325000 ;
      RECT 1932.150000  1.325000 1932.350000 2.295000 ;
      RECT 1932.150000  2.295000 1934.495000 2.465000 ;
      RECT 1932.515000  0.255000 1933.200000 0.620000 ;
      RECT 1932.515000  0.620000 1932.690000 0.655000 ;
      RECT 1932.520000  0.825000 1932.690000 1.955000 ;
      RECT 1932.520000  1.955000 1933.965000 2.125000 ;
      RECT 1932.860000  0.810000 1933.030000 1.615000 ;
      RECT 1932.860000  1.615000 1934.155000 1.785000 ;
      RECT 1933.370000  0.255000 1933.695000 1.415000 ;
      RECT 1933.865000  0.255000 1934.155000 1.615000 ;
      RECT 1934.325000  1.440000 1935.075000 1.630000 ;
      RECT 1934.325000  1.630000 1934.495000 2.295000 ;
      RECT 1934.330000  0.085000 1934.845000 0.525000 ;
      RECT 1934.405000  0.695000 1935.465000 0.865000 ;
      RECT 1934.405000  0.865000 1934.575000 1.185000 ;
      RECT 1934.665000  1.835000 1934.895000 2.635000 ;
      RECT 1934.885000  1.055000 1935.075000 1.440000 ;
      RECT 1935.065000  1.835000 1935.465000 2.465000 ;
      RECT 1935.115000  0.255000 1935.360000 0.695000 ;
      RECT 1935.295000  0.865000 1935.465000 1.835000 ;
      RECT 1935.765000  0.085000 1936.055000 0.810000 ;
      RECT 1935.765000  1.470000 1936.055000 2.635000 ;
      RECT 1936.275000  1.495000 1936.535000 2.635000 ;
      RECT 1936.315000  0.085000 1936.560000 0.655000 ;
      RECT 1936.705000  1.495000 1937.035000 2.465000 ;
      RECT 1936.730000  0.255000 1936.990000 1.065000 ;
      RECT 1936.730000  1.065000 1937.885000 1.325000 ;
      RECT 1936.730000  1.325000 1936.990000 1.495000 ;
      RECT 1937.195000  0.085000 1937.445000 0.655000 ;
      RECT 1937.205000  1.495000 1937.445000 2.635000 ;
      RECT 1937.615000  0.255000 1937.885000 1.065000 ;
      RECT 1937.615000  1.325000 1937.885000 1.495000 ;
      RECT 1937.615000  1.495000 1937.975000 2.465000 ;
      RECT 1938.055000  0.085000 1938.415000 0.485000 ;
      RECT 1938.055000  0.655000 1939.130000 0.825000 ;
      RECT 1938.055000  0.825000 1938.225000 1.325000 ;
      RECT 1938.145000  1.495000 1938.420000 2.635000 ;
      RECT 1938.515000  0.995000 1938.790000 1.325000 ;
      RECT 1938.590000  1.325000 1938.790000 2.295000 ;
      RECT 1938.590000  2.295000 1940.935000 2.465000 ;
      RECT 1938.955000  0.255000 1939.640000 0.620000 ;
      RECT 1938.955000  0.620000 1939.130000 0.655000 ;
      RECT 1938.960000  0.825000 1939.130000 1.955000 ;
      RECT 1938.960000  1.955000 1940.405000 2.125000 ;
      RECT 1939.300000  0.810000 1939.470000 1.615000 ;
      RECT 1939.300000  1.615000 1940.595000 1.785000 ;
      RECT 1939.810000  0.255000 1940.135000 1.415000 ;
      RECT 1940.305000  0.255000 1940.595000 1.615000 ;
      RECT 1940.765000  1.440000 1941.515000 1.630000 ;
      RECT 1940.765000  1.630000 1940.935000 2.295000 ;
      RECT 1940.770000  0.085000 1941.285000 0.525000 ;
      RECT 1940.845000  0.695000 1941.905000 0.865000 ;
      RECT 1940.845000  0.865000 1941.015000 1.185000 ;
      RECT 1941.105000  1.835000 1941.335000 2.635000 ;
      RECT 1941.325000  1.055000 1941.515000 1.440000 ;
      RECT 1941.505000  1.835000 1941.905000 2.465000 ;
      RECT 1941.555000  0.255000 1941.800000 0.695000 ;
      RECT 1941.735000  0.865000 1941.905000 1.835000 ;
      RECT 1942.120000  5.355000 2064.020000 5.525000 ;
      RECT 1942.205000  0.085000 1942.495000 0.810000 ;
      RECT 1942.205000  1.470000 1942.495000 2.635000 ;
      RECT 1942.205000  2.805000 1942.495000 3.970000 ;
      RECT 1942.205000  4.630000 1942.495000 5.355000 ;
      RECT 1942.665000  0.995000 1943.260000 1.325000 ;
      RECT 1942.665000  4.115000 1943.260000 4.445000 ;
      RECT 1942.800000  1.605000 1943.100000 2.635000 ;
      RECT 1942.800000  2.805000 1943.100000 3.835000 ;
      RECT 1942.850000  0.085000 1943.140000 0.610000 ;
      RECT 1942.850000  4.830000 1943.140000 5.355000 ;
      RECT 1943.270000  1.605000 1943.600000 2.465000 ;
      RECT 1943.270000  2.975000 1943.600000 3.835000 ;
      RECT 1943.350000  0.280000 1943.600000 0.825000 ;
      RECT 1943.350000  4.615000 1943.600000 5.160000 ;
      RECT 1943.430000  0.825000 1943.600000 1.065000 ;
      RECT 1943.430000  1.065000 1944.615000 1.395000 ;
      RECT 1943.430000  1.395000 1943.600000 1.605000 ;
      RECT 1943.430000  3.835000 1943.600000 4.045000 ;
      RECT 1943.430000  4.045000 1944.615000 4.375000 ;
      RECT 1943.430000  4.375000 1943.600000 4.615000 ;
      RECT 1943.770000  0.085000 1944.060000 0.610000 ;
      RECT 1943.770000  4.830000 1944.060000 5.355000 ;
      RECT 1943.795000  1.605000 1944.070000 2.635000 ;
      RECT 1943.795000  2.805000 1944.070000 3.835000 ;
      RECT 1944.315000  1.565000 1944.615000 2.465000 ;
      RECT 1944.315000  2.975000 1944.615000 3.875000 ;
      RECT 1944.565000  0.255000 1946.595000 0.425000 ;
      RECT 1944.565000  0.425000 1944.815000 0.770000 ;
      RECT 1944.565000  4.670000 1944.815000 5.015000 ;
      RECT 1944.565000  5.015000 1946.595000 5.185000 ;
      RECT 1944.785000  1.065000 1946.055000 1.365000 ;
      RECT 1944.785000  1.365000 1945.115000 4.075000 ;
      RECT 1944.785000  4.075000 1946.055000 4.375000 ;
      RECT 1944.985000  0.595000 1945.315000 1.065000 ;
      RECT 1944.985000  4.375000 1945.315000 4.845000 ;
      RECT 1945.285000  1.535000 1945.555000 2.465000 ;
      RECT 1945.285000  2.975000 1945.555000 3.905000 ;
      RECT 1945.485000  0.425000 1945.655000 0.770000 ;
      RECT 1945.485000  4.670000 1945.655000 5.015000 ;
      RECT 1945.725000  1.365000 1946.055000 4.075000 ;
      RECT 1945.825000  0.595000 1946.155000 0.885000 ;
      RECT 1945.825000  0.885000 1946.055000 1.065000 ;
      RECT 1945.825000  4.375000 1946.055000 4.555000 ;
      RECT 1945.825000  4.555000 1946.155000 4.845000 ;
      RECT 1946.225000  1.495000 1948.455000 1.665000 ;
      RECT 1946.225000  1.665000 1946.525000 2.465000 ;
      RECT 1946.225000  2.635000 1951.355000 2.805000 ;
      RECT 1946.225000  2.975000 1946.525000 3.775000 ;
      RECT 1946.225000  3.775000 1948.455000 3.945000 ;
      RECT 1946.325000  0.425000 1946.595000 0.715000 ;
      RECT 1946.325000  0.715000 1948.455000 0.885000 ;
      RECT 1946.325000  4.555000 1948.455000 4.725000 ;
      RECT 1946.325000  4.725000 1946.595000 5.015000 ;
      RECT 1946.745000  1.835000 1947.015000 2.635000 ;
      RECT 1946.745000  2.805000 1947.015000 3.605000 ;
      RECT 1946.765000  0.085000 1947.015000 0.545000 ;
      RECT 1946.765000  4.895000 1947.015000 5.355000 ;
      RECT 1947.185000  0.255000 1947.515000 0.715000 ;
      RECT 1947.185000  1.665000 1947.515000 2.465000 ;
      RECT 1947.185000  2.975000 1947.515000 3.775000 ;
      RECT 1947.185000  4.725000 1947.515000 5.185000 ;
      RECT 1947.235000  1.055000 1948.625000 1.325000 ;
      RECT 1947.235000  4.115000 1948.625000 4.385000 ;
      RECT 1947.685000  0.085000 1947.955000 0.545000 ;
      RECT 1947.685000  1.835000 1947.955000 2.635000 ;
      RECT 1947.685000  2.805000 1947.955000 3.605000 ;
      RECT 1947.685000  4.895000 1947.955000 5.355000 ;
      RECT 1948.125000  0.255000 1948.455000 0.715000 ;
      RECT 1948.125000  1.665000 1948.455000 2.465000 ;
      RECT 1948.125000  2.975000 1948.455000 3.775000 ;
      RECT 1948.125000  4.725000 1948.455000 5.185000 ;
      RECT 1948.625000  0.085000 1948.955000 0.885000 ;
      RECT 1948.625000  1.495000 1948.955000 2.635000 ;
      RECT 1948.625000  2.805000 1948.955000 3.945000 ;
      RECT 1948.625000  4.555000 1948.955000 5.355000 ;
      RECT 1948.955000  1.055000 1950.345000 1.325000 ;
      RECT 1948.955000  4.115000 1950.345000 4.385000 ;
      RECT 1949.125000  0.255000 1949.455000 0.715000 ;
      RECT 1949.125000  0.715000 1951.255000 0.885000 ;
      RECT 1949.125000  1.495000 1951.355000 1.665000 ;
      RECT 1949.125000  1.665000 1949.455000 2.465000 ;
      RECT 1949.125000  2.975000 1949.455000 3.775000 ;
      RECT 1949.125000  3.775000 1951.355000 3.945000 ;
      RECT 1949.125000  4.555000 1951.255000 4.725000 ;
      RECT 1949.125000  4.725000 1949.455000 5.185000 ;
      RECT 1949.625000  0.085000 1949.895000 0.545000 ;
      RECT 1949.625000  1.835000 1949.895000 2.635000 ;
      RECT 1949.625000  2.805000 1949.895000 3.605000 ;
      RECT 1949.625000  4.895000 1949.895000 5.355000 ;
      RECT 1950.065000  0.255000 1950.395000 0.715000 ;
      RECT 1950.065000  1.665000 1950.395000 2.465000 ;
      RECT 1950.065000  2.975000 1950.395000 3.775000 ;
      RECT 1950.065000  4.725000 1950.395000 5.185000 ;
      RECT 1950.565000  0.085000 1950.815000 0.545000 ;
      RECT 1950.565000  1.835000 1950.835000 2.635000 ;
      RECT 1950.565000  2.805000 1950.835000 3.605000 ;
      RECT 1950.565000  4.895000 1950.815000 5.355000 ;
      RECT 1950.985000  0.255000 1953.015000 0.425000 ;
      RECT 1950.985000  0.425000 1951.255000 0.715000 ;
      RECT 1950.985000  4.725000 1951.255000 5.015000 ;
      RECT 1950.985000  5.015000 1953.015000 5.185000 ;
      RECT 1951.055000  1.665000 1951.355000 2.465000 ;
      RECT 1951.055000  2.975000 1951.355000 3.775000 ;
      RECT 1951.425000  0.595000 1951.755000 0.885000 ;
      RECT 1951.425000  4.555000 1951.755000 4.845000 ;
      RECT 1951.525000  0.885000 1951.755000 1.065000 ;
      RECT 1951.525000  1.065000 1952.795000 1.365000 ;
      RECT 1951.525000  1.365000 1951.855000 4.075000 ;
      RECT 1951.525000  4.075000 1952.795000 4.375000 ;
      RECT 1951.525000  4.375000 1951.755000 4.555000 ;
      RECT 1951.925000  0.425000 1952.095000 0.770000 ;
      RECT 1951.925000  4.670000 1952.095000 5.015000 ;
      RECT 1952.025000  1.535000 1952.295000 2.465000 ;
      RECT 1952.025000  2.975000 1952.295000 3.905000 ;
      RECT 1952.265000  0.595000 1952.595000 1.065000 ;
      RECT 1952.265000  4.375000 1952.595000 4.845000 ;
      RECT 1952.465000  1.365000 1952.795000 4.075000 ;
      RECT 1952.765000  0.425000 1953.015000 0.770000 ;
      RECT 1952.765000  4.670000 1953.015000 5.015000 ;
      RECT 1952.965000  1.065000 1954.150000 1.395000 ;
      RECT 1952.965000  1.565000 1953.265000 2.465000 ;
      RECT 1952.965000  2.635000 1957.035000 2.805000 ;
      RECT 1952.965000  2.975000 1953.265000 3.875000 ;
      RECT 1952.965000  4.045000 1954.150000 4.375000 ;
      RECT 1953.510000  1.605000 1953.785000 2.635000 ;
      RECT 1953.510000  2.805000 1953.785000 3.835000 ;
      RECT 1953.520000  0.085000 1953.810000 0.610000 ;
      RECT 1953.520000  4.830000 1953.810000 5.355000 ;
      RECT 1953.980000  0.280000 1954.230000 0.825000 ;
      RECT 1953.980000  0.825000 1954.150000 1.065000 ;
      RECT 1953.980000  1.395000 1954.150000 1.605000 ;
      RECT 1953.980000  1.605000 1954.310000 2.465000 ;
      RECT 1953.980000  2.975000 1954.310000 3.835000 ;
      RECT 1953.980000  3.835000 1954.150000 4.045000 ;
      RECT 1953.980000  4.375000 1954.150000 4.615000 ;
      RECT 1953.980000  4.615000 1954.230000 5.160000 ;
      RECT 1954.320000  0.995000 1954.915000 1.325000 ;
      RECT 1954.320000  4.115000 1954.915000 4.445000 ;
      RECT 1954.440000  0.085000 1954.730000 0.610000 ;
      RECT 1954.440000  4.830000 1954.730000 5.355000 ;
      RECT 1954.480000  1.605000 1954.780000 2.635000 ;
      RECT 1954.480000  2.805000 1954.780000 3.835000 ;
      RECT 1955.085000  0.995000 1955.680000 1.325000 ;
      RECT 1955.085000  4.115000 1955.680000 4.445000 ;
      RECT 1955.220000  1.605000 1955.520000 2.635000 ;
      RECT 1955.220000  2.805000 1955.520000 3.835000 ;
      RECT 1955.270000  0.085000 1955.560000 0.610000 ;
      RECT 1955.270000  4.830000 1955.560000 5.355000 ;
      RECT 1955.690000  1.605000 1956.020000 2.465000 ;
      RECT 1955.690000  2.975000 1956.020000 3.835000 ;
      RECT 1955.770000  0.280000 1956.020000 0.825000 ;
      RECT 1955.770000  4.615000 1956.020000 5.160000 ;
      RECT 1955.850000  0.825000 1956.020000 1.065000 ;
      RECT 1955.850000  1.065000 1957.035000 1.395000 ;
      RECT 1955.850000  1.395000 1956.020000 1.605000 ;
      RECT 1955.850000  3.835000 1956.020000 4.045000 ;
      RECT 1955.850000  4.045000 1957.035000 4.375000 ;
      RECT 1955.850000  4.375000 1956.020000 4.615000 ;
      RECT 1956.190000  0.085000 1956.480000 0.610000 ;
      RECT 1956.190000  4.830000 1956.480000 5.355000 ;
      RECT 1956.215000  1.605000 1956.490000 2.635000 ;
      RECT 1956.215000  2.805000 1956.490000 3.835000 ;
      RECT 1956.735000  1.565000 1957.035000 2.465000 ;
      RECT 1956.735000  2.975000 1957.035000 3.875000 ;
      RECT 1956.985000  0.255000 1959.015000 0.425000 ;
      RECT 1956.985000  0.425000 1957.235000 0.770000 ;
      RECT 1956.985000  4.670000 1957.235000 5.015000 ;
      RECT 1956.985000  5.015000 1959.015000 5.185000 ;
      RECT 1957.205000  1.065000 1958.475000 1.365000 ;
      RECT 1957.205000  1.365000 1957.535000 4.075000 ;
      RECT 1957.205000  4.075000 1958.475000 4.375000 ;
      RECT 1957.405000  0.595000 1957.735000 1.065000 ;
      RECT 1957.405000  4.375000 1957.735000 4.845000 ;
      RECT 1957.705000  1.535000 1957.975000 2.465000 ;
      RECT 1957.705000  2.975000 1957.975000 3.905000 ;
      RECT 1957.905000  0.425000 1958.075000 0.770000 ;
      RECT 1957.905000  4.670000 1958.075000 5.015000 ;
      RECT 1958.145000  1.365000 1958.475000 4.075000 ;
      RECT 1958.245000  0.595000 1958.575000 0.885000 ;
      RECT 1958.245000  0.885000 1958.475000 1.065000 ;
      RECT 1958.245000  4.375000 1958.475000 4.555000 ;
      RECT 1958.245000  4.555000 1958.575000 4.845000 ;
      RECT 1958.645000  1.495000 1960.875000 1.665000 ;
      RECT 1958.645000  1.665000 1958.945000 2.465000 ;
      RECT 1958.645000  2.635000 1963.775000 2.805000 ;
      RECT 1958.645000  2.975000 1958.945000 3.775000 ;
      RECT 1958.645000  3.775000 1960.875000 3.945000 ;
      RECT 1958.745000  0.425000 1959.015000 0.715000 ;
      RECT 1958.745000  0.715000 1960.875000 0.885000 ;
      RECT 1958.745000  4.555000 1960.875000 4.725000 ;
      RECT 1958.745000  4.725000 1959.015000 5.015000 ;
      RECT 1959.165000  1.835000 1959.435000 2.635000 ;
      RECT 1959.165000  2.805000 1959.435000 3.605000 ;
      RECT 1959.185000  0.085000 1959.435000 0.545000 ;
      RECT 1959.185000  4.895000 1959.435000 5.355000 ;
      RECT 1959.605000  0.255000 1959.935000 0.715000 ;
      RECT 1959.605000  1.665000 1959.935000 2.465000 ;
      RECT 1959.605000  2.975000 1959.935000 3.775000 ;
      RECT 1959.605000  4.725000 1959.935000 5.185000 ;
      RECT 1959.655000  1.055000 1961.045000 1.325000 ;
      RECT 1959.655000  4.115000 1961.045000 4.385000 ;
      RECT 1960.105000  0.085000 1960.375000 0.545000 ;
      RECT 1960.105000  1.835000 1960.375000 2.635000 ;
      RECT 1960.105000  2.805000 1960.375000 3.605000 ;
      RECT 1960.105000  4.895000 1960.375000 5.355000 ;
      RECT 1960.545000  0.255000 1960.875000 0.715000 ;
      RECT 1960.545000  1.665000 1960.875000 2.465000 ;
      RECT 1960.545000  2.975000 1960.875000 3.775000 ;
      RECT 1960.545000  4.725000 1960.875000 5.185000 ;
      RECT 1961.045000  0.085000 1961.375000 0.885000 ;
      RECT 1961.045000  1.495000 1961.375000 2.635000 ;
      RECT 1961.045000  2.805000 1961.375000 3.945000 ;
      RECT 1961.045000  4.555000 1961.375000 5.355000 ;
      RECT 1961.375000  1.055000 1962.765000 1.325000 ;
      RECT 1961.375000  4.115000 1962.765000 4.385000 ;
      RECT 1961.545000  0.255000 1961.875000 0.715000 ;
      RECT 1961.545000  0.715000 1963.675000 0.885000 ;
      RECT 1961.545000  1.495000 1963.775000 1.665000 ;
      RECT 1961.545000  1.665000 1961.875000 2.465000 ;
      RECT 1961.545000  2.975000 1961.875000 3.775000 ;
      RECT 1961.545000  3.775000 1963.775000 3.945000 ;
      RECT 1961.545000  4.555000 1963.675000 4.725000 ;
      RECT 1961.545000  4.725000 1961.875000 5.185000 ;
      RECT 1962.045000  0.085000 1962.315000 0.545000 ;
      RECT 1962.045000  1.835000 1962.315000 2.635000 ;
      RECT 1962.045000  2.805000 1962.315000 3.605000 ;
      RECT 1962.045000  4.895000 1962.315000 5.355000 ;
      RECT 1962.485000  0.255000 1962.815000 0.715000 ;
      RECT 1962.485000  1.665000 1962.815000 2.465000 ;
      RECT 1962.485000  2.975000 1962.815000 3.775000 ;
      RECT 1962.485000  4.725000 1962.815000 5.185000 ;
      RECT 1962.985000  0.085000 1963.235000 0.545000 ;
      RECT 1962.985000  1.835000 1963.255000 2.635000 ;
      RECT 1962.985000  2.805000 1963.255000 3.605000 ;
      RECT 1962.985000  4.895000 1963.235000 5.355000 ;
      RECT 1963.405000  0.255000 1965.435000 0.425000 ;
      RECT 1963.405000  0.425000 1963.675000 0.715000 ;
      RECT 1963.405000  4.725000 1963.675000 5.015000 ;
      RECT 1963.405000  5.015000 1965.435000 5.185000 ;
      RECT 1963.475000  1.665000 1963.775000 2.465000 ;
      RECT 1963.475000  2.975000 1963.775000 3.775000 ;
      RECT 1963.845000  0.595000 1964.175000 0.885000 ;
      RECT 1963.845000  4.555000 1964.175000 4.845000 ;
      RECT 1963.945000  0.885000 1964.175000 1.065000 ;
      RECT 1963.945000  1.065000 1965.215000 1.365000 ;
      RECT 1963.945000  1.365000 1964.275000 4.075000 ;
      RECT 1963.945000  4.075000 1965.215000 4.375000 ;
      RECT 1963.945000  4.375000 1964.175000 4.555000 ;
      RECT 1964.345000  0.425000 1964.515000 0.770000 ;
      RECT 1964.345000  4.670000 1964.515000 5.015000 ;
      RECT 1964.445000  1.535000 1964.715000 2.465000 ;
      RECT 1964.445000  2.975000 1964.715000 3.905000 ;
      RECT 1964.685000  0.595000 1965.015000 1.065000 ;
      RECT 1964.685000  4.375000 1965.015000 4.845000 ;
      RECT 1964.885000  1.365000 1965.215000 4.075000 ;
      RECT 1965.185000  0.425000 1965.435000 0.770000 ;
      RECT 1965.185000  4.670000 1965.435000 5.015000 ;
      RECT 1965.385000  1.065000 1966.570000 1.395000 ;
      RECT 1965.385000  1.565000 1965.685000 2.465000 ;
      RECT 1965.385000  2.635000 1968.800000 2.805000 ;
      RECT 1965.385000  2.975000 1965.685000 3.875000 ;
      RECT 1965.385000  4.045000 1966.570000 4.375000 ;
      RECT 1965.930000  1.605000 1966.205000 2.635000 ;
      RECT 1965.930000  2.805000 1966.205000 3.835000 ;
      RECT 1965.940000  0.085000 1966.230000 0.610000 ;
      RECT 1965.940000  4.830000 1966.230000 5.355000 ;
      RECT 1966.400000  0.280000 1966.650000 0.825000 ;
      RECT 1966.400000  0.825000 1966.570000 1.065000 ;
      RECT 1966.400000  1.395000 1966.570000 1.605000 ;
      RECT 1966.400000  1.605000 1966.730000 2.465000 ;
      RECT 1966.400000  2.975000 1966.730000 3.835000 ;
      RECT 1966.400000  3.835000 1966.570000 4.045000 ;
      RECT 1966.400000  4.375000 1966.570000 4.615000 ;
      RECT 1966.400000  4.615000 1966.650000 5.160000 ;
      RECT 1966.740000  0.995000 1967.335000 1.325000 ;
      RECT 1966.740000  4.115000 1967.335000 4.445000 ;
      RECT 1966.860000  0.085000 1967.150000 0.610000 ;
      RECT 1966.860000  4.830000 1967.150000 5.355000 ;
      RECT 1966.900000  1.605000 1967.200000 2.635000 ;
      RECT 1966.900000  2.805000 1967.200000 3.835000 ;
      RECT 1967.505000  0.085000 1967.795000 0.810000 ;
      RECT 1967.505000  1.470000 1967.795000 2.635000 ;
      RECT 1967.505000  2.805000 1967.795000 3.970000 ;
      RECT 1967.505000  4.630000 1967.795000 5.355000 ;
      RECT 1967.975000  1.495000 1968.305000 2.635000 ;
      RECT 1967.975000  2.805000 1968.305000 3.945000 ;
      RECT 1968.010000  0.085000 1968.270000 0.885000 ;
      RECT 1968.010000  4.555000 1968.270000 5.355000 ;
      RECT 1968.215000  1.055000 1968.610000 1.325000 ;
      RECT 1968.215000  4.115000 1968.610000 4.385000 ;
      RECT 1968.440000  0.395000 1968.715000 0.625000 ;
      RECT 1968.440000  0.625000 1968.610000 1.055000 ;
      RECT 1968.440000  4.385000 1968.610000 4.815000 ;
      RECT 1968.440000  4.815000 1968.715000 5.045000 ;
      RECT 1968.780000  0.835000 1969.170000 1.005000 ;
      RECT 1968.780000  1.005000 1968.950000 1.755000 ;
      RECT 1968.780000  1.755000 1969.175000 1.805000 ;
      RECT 1968.780000  1.805000 1969.300000 1.985000 ;
      RECT 1968.780000  3.455000 1969.300000 3.635000 ;
      RECT 1968.780000  3.635000 1969.175000 3.685000 ;
      RECT 1968.780000  3.685000 1968.950000 4.435000 ;
      RECT 1968.780000  4.435000 1969.170000 4.605000 ;
      RECT 1968.925000  0.330000 1969.170000 0.835000 ;
      RECT 1968.925000  4.605000 1969.170000 5.110000 ;
      RECT 1968.970000  1.985000 1969.300000 2.465000 ;
      RECT 1968.970000  2.465000 1969.175000 2.975000 ;
      RECT 1968.970000  2.975000 1969.300000 3.455000 ;
      RECT 1969.120000  1.175000 1969.510000 1.465000 ;
      RECT 1969.120000  1.465000 1969.820000 1.505000 ;
      RECT 1969.120000  3.935000 1969.820000 3.975000 ;
      RECT 1969.120000  3.975000 1969.510000 4.265000 ;
      RECT 1969.340000  0.585000 1969.780000 0.755000 ;
      RECT 1969.340000  0.755000 1969.510000 1.175000 ;
      RECT 1969.340000  1.505000 1969.820000 1.635000 ;
      RECT 1969.340000  3.805000 1969.820000 3.935000 ;
      RECT 1969.340000  4.265000 1969.510000 4.685000 ;
      RECT 1969.340000  4.685000 1969.780000 4.855000 ;
      RECT 1969.345000  2.635000 1971.015000 2.805000 ;
      RECT 1969.490000  1.635000 1969.820000 2.465000 ;
      RECT 1969.490000  2.975000 1969.820000 3.805000 ;
      RECT 1969.530000  0.330000 1969.780000 0.585000 ;
      RECT 1969.530000  4.855000 1969.780000 5.110000 ;
      RECT 1969.685000  0.945000 1970.085000 1.295000 ;
      RECT 1969.685000  4.145000 1970.085000 4.495000 ;
      RECT 1970.015000  0.085000 1970.345000 0.660000 ;
      RECT 1970.015000  1.465000 1970.345000 2.635000 ;
      RECT 1970.015000  2.805000 1970.345000 3.975000 ;
      RECT 1970.015000  4.780000 1970.345000 5.355000 ;
      RECT 1970.275000  0.945000 1970.675000 1.295000 ;
      RECT 1970.275000  4.145000 1970.675000 4.495000 ;
      RECT 1970.540000  1.465000 1971.240000 1.505000 ;
      RECT 1970.540000  1.505000 1971.020000 1.635000 ;
      RECT 1970.540000  1.635000 1970.870000 2.465000 ;
      RECT 1970.540000  2.975000 1970.870000 3.805000 ;
      RECT 1970.540000  3.805000 1971.020000 3.935000 ;
      RECT 1970.540000  3.935000 1971.240000 3.975000 ;
      RECT 1970.580000  0.330000 1970.830000 0.585000 ;
      RECT 1970.580000  0.585000 1971.020000 0.755000 ;
      RECT 1970.580000  4.685000 1971.020000 4.855000 ;
      RECT 1970.580000  4.855000 1970.830000 5.110000 ;
      RECT 1970.850000  0.755000 1971.020000 1.175000 ;
      RECT 1970.850000  1.175000 1971.240000 1.465000 ;
      RECT 1970.850000  3.975000 1971.240000 4.265000 ;
      RECT 1970.850000  4.265000 1971.020000 4.685000 ;
      RECT 1971.060000  1.805000 1971.580000 1.985000 ;
      RECT 1971.060000  1.985000 1971.390000 2.465000 ;
      RECT 1971.060000  2.975000 1971.390000 3.455000 ;
      RECT 1971.060000  3.455000 1971.580000 3.635000 ;
      RECT 1971.185000  1.755000 1971.580000 1.805000 ;
      RECT 1971.185000  2.465000 1971.390000 2.975000 ;
      RECT 1971.185000  3.635000 1971.580000 3.685000 ;
      RECT 1971.190000  0.330000 1971.435000 0.835000 ;
      RECT 1971.190000  0.835000 1971.580000 1.005000 ;
      RECT 1971.190000  4.435000 1971.580000 4.605000 ;
      RECT 1971.190000  4.605000 1971.435000 5.110000 ;
      RECT 1971.410000  1.005000 1971.580000 1.755000 ;
      RECT 1971.410000  3.685000 1971.580000 4.435000 ;
      RECT 1971.560000  2.635000 1972.940000 2.805000 ;
      RECT 1971.645000  0.395000 1971.920000 0.625000 ;
      RECT 1971.645000  4.815000 1971.920000 5.045000 ;
      RECT 1971.750000  0.625000 1971.920000 1.055000 ;
      RECT 1971.750000  1.055000 1972.145000 1.325000 ;
      RECT 1971.750000  4.115000 1972.145000 4.385000 ;
      RECT 1971.750000  4.385000 1971.920000 4.815000 ;
      RECT 1972.055000  1.495000 1972.445000 2.635000 ;
      RECT 1972.055000  2.805000 1972.445000 3.945000 ;
      RECT 1972.090000  0.085000 1972.410000 0.885000 ;
      RECT 1972.090000  4.555000 1972.410000 5.355000 ;
      RECT 1972.355000  1.055000 1972.750000 1.325000 ;
      RECT 1972.355000  4.115000 1972.750000 4.385000 ;
      RECT 1972.580000  0.395000 1972.855000 0.625000 ;
      RECT 1972.580000  0.625000 1972.750000 1.055000 ;
      RECT 1972.580000  4.385000 1972.750000 4.815000 ;
      RECT 1972.580000  4.815000 1972.855000 5.045000 ;
      RECT 1972.920000  0.835000 1973.310000 1.005000 ;
      RECT 1972.920000  1.005000 1973.090000 1.755000 ;
      RECT 1972.920000  1.755000 1973.315000 1.805000 ;
      RECT 1972.920000  1.805000 1973.440000 1.985000 ;
      RECT 1972.920000  3.455000 1973.440000 3.635000 ;
      RECT 1972.920000  3.635000 1973.315000 3.685000 ;
      RECT 1972.920000  3.685000 1973.090000 4.435000 ;
      RECT 1972.920000  4.435000 1973.310000 4.605000 ;
      RECT 1973.065000  0.330000 1973.310000 0.835000 ;
      RECT 1973.065000  4.605000 1973.310000 5.110000 ;
      RECT 1973.110000  1.985000 1973.440000 2.465000 ;
      RECT 1973.110000  2.465000 1973.315000 2.975000 ;
      RECT 1973.110000  2.975000 1973.440000 3.455000 ;
      RECT 1973.260000  1.175000 1973.650000 1.465000 ;
      RECT 1973.260000  1.465000 1973.960000 1.505000 ;
      RECT 1973.260000  3.935000 1973.960000 3.975000 ;
      RECT 1973.260000  3.975000 1973.650000 4.265000 ;
      RECT 1973.480000  0.585000 1973.920000 0.755000 ;
      RECT 1973.480000  0.755000 1973.650000 1.175000 ;
      RECT 1973.480000  1.505000 1973.960000 1.635000 ;
      RECT 1973.480000  3.805000 1973.960000 3.935000 ;
      RECT 1973.480000  4.265000 1973.650000 4.685000 ;
      RECT 1973.480000  4.685000 1973.920000 4.855000 ;
      RECT 1973.485000  2.635000 1975.155000 2.805000 ;
      RECT 1973.630000  1.635000 1973.960000 2.465000 ;
      RECT 1973.630000  2.975000 1973.960000 3.805000 ;
      RECT 1973.670000  0.330000 1973.920000 0.585000 ;
      RECT 1973.670000  4.855000 1973.920000 5.110000 ;
      RECT 1973.825000  0.945000 1974.225000 1.295000 ;
      RECT 1973.825000  4.145000 1974.225000 4.495000 ;
      RECT 1974.155000  0.085000 1974.485000 0.660000 ;
      RECT 1974.155000  1.465000 1974.485000 2.635000 ;
      RECT 1974.155000  2.805000 1974.485000 3.975000 ;
      RECT 1974.155000  4.780000 1974.485000 5.355000 ;
      RECT 1974.415000  0.945000 1974.815000 1.295000 ;
      RECT 1974.415000  4.145000 1974.815000 4.495000 ;
      RECT 1974.680000  1.465000 1975.380000 1.505000 ;
      RECT 1974.680000  1.505000 1975.160000 1.635000 ;
      RECT 1974.680000  1.635000 1975.010000 2.465000 ;
      RECT 1974.680000  2.975000 1975.010000 3.805000 ;
      RECT 1974.680000  3.805000 1975.160000 3.935000 ;
      RECT 1974.680000  3.935000 1975.380000 3.975000 ;
      RECT 1974.720000  0.330000 1974.970000 0.585000 ;
      RECT 1974.720000  0.585000 1975.160000 0.755000 ;
      RECT 1974.720000  4.685000 1975.160000 4.855000 ;
      RECT 1974.720000  4.855000 1974.970000 5.110000 ;
      RECT 1974.990000  0.755000 1975.160000 1.175000 ;
      RECT 1974.990000  1.175000 1975.380000 1.465000 ;
      RECT 1974.990000  3.975000 1975.380000 4.265000 ;
      RECT 1974.990000  4.265000 1975.160000 4.685000 ;
      RECT 1975.200000  1.805000 1975.720000 1.985000 ;
      RECT 1975.200000  1.985000 1975.530000 2.465000 ;
      RECT 1975.200000  2.975000 1975.530000 3.455000 ;
      RECT 1975.200000  3.455000 1975.720000 3.635000 ;
      RECT 1975.325000  1.755000 1975.720000 1.805000 ;
      RECT 1975.325000  2.465000 1975.530000 2.975000 ;
      RECT 1975.325000  3.635000 1975.720000 3.685000 ;
      RECT 1975.330000  0.330000 1975.575000 0.835000 ;
      RECT 1975.330000  0.835000 1975.720000 1.005000 ;
      RECT 1975.330000  4.435000 1975.720000 4.605000 ;
      RECT 1975.330000  4.605000 1975.575000 5.110000 ;
      RECT 1975.550000  1.005000 1975.720000 1.755000 ;
      RECT 1975.550000  3.685000 1975.720000 4.435000 ;
      RECT 1975.700000  2.635000 1977.080000 2.805000 ;
      RECT 1975.785000  0.395000 1976.060000 0.625000 ;
      RECT 1975.785000  4.815000 1976.060000 5.045000 ;
      RECT 1975.890000  0.625000 1976.060000 1.055000 ;
      RECT 1975.890000  1.055000 1976.285000 1.325000 ;
      RECT 1975.890000  4.115000 1976.285000 4.385000 ;
      RECT 1975.890000  4.385000 1976.060000 4.815000 ;
      RECT 1976.195000  1.495000 1976.585000 2.635000 ;
      RECT 1976.195000  2.805000 1976.585000 3.945000 ;
      RECT 1976.230000  0.085000 1976.550000 0.885000 ;
      RECT 1976.230000  4.555000 1976.550000 5.355000 ;
      RECT 1976.495000  1.055000 1976.890000 1.325000 ;
      RECT 1976.495000  4.115000 1976.890000 4.385000 ;
      RECT 1976.720000  0.395000 1976.995000 0.625000 ;
      RECT 1976.720000  0.625000 1976.890000 1.055000 ;
      RECT 1976.720000  4.385000 1976.890000 4.815000 ;
      RECT 1976.720000  4.815000 1976.995000 5.045000 ;
      RECT 1977.060000  0.835000 1977.450000 1.005000 ;
      RECT 1977.060000  1.005000 1977.230000 1.755000 ;
      RECT 1977.060000  1.755000 1977.455000 1.805000 ;
      RECT 1977.060000  1.805000 1977.580000 1.985000 ;
      RECT 1977.060000  3.455000 1977.580000 3.635000 ;
      RECT 1977.060000  3.635000 1977.455000 3.685000 ;
      RECT 1977.060000  3.685000 1977.230000 4.435000 ;
      RECT 1977.060000  4.435000 1977.450000 4.605000 ;
      RECT 1977.205000  0.330000 1977.450000 0.835000 ;
      RECT 1977.205000  4.605000 1977.450000 5.110000 ;
      RECT 1977.250000  1.985000 1977.580000 2.465000 ;
      RECT 1977.250000  2.465000 1977.455000 2.975000 ;
      RECT 1977.250000  2.975000 1977.580000 3.455000 ;
      RECT 1977.400000  1.175000 1977.790000 1.465000 ;
      RECT 1977.400000  1.465000 1978.100000 1.505000 ;
      RECT 1977.400000  3.935000 1978.100000 3.975000 ;
      RECT 1977.400000  3.975000 1977.790000 4.265000 ;
      RECT 1977.620000  0.585000 1978.060000 0.755000 ;
      RECT 1977.620000  0.755000 1977.790000 1.175000 ;
      RECT 1977.620000  1.505000 1978.100000 1.635000 ;
      RECT 1977.620000  3.805000 1978.100000 3.935000 ;
      RECT 1977.620000  4.265000 1977.790000 4.685000 ;
      RECT 1977.620000  4.685000 1978.060000 4.855000 ;
      RECT 1977.625000  2.635000 1979.295000 2.805000 ;
      RECT 1977.770000  1.635000 1978.100000 2.465000 ;
      RECT 1977.770000  2.975000 1978.100000 3.805000 ;
      RECT 1977.810000  0.330000 1978.060000 0.585000 ;
      RECT 1977.810000  4.855000 1978.060000 5.110000 ;
      RECT 1977.965000  0.945000 1978.365000 1.295000 ;
      RECT 1977.965000  4.145000 1978.365000 4.495000 ;
      RECT 1978.295000  0.085000 1978.625000 0.660000 ;
      RECT 1978.295000  1.465000 1978.625000 2.635000 ;
      RECT 1978.295000  2.805000 1978.625000 3.975000 ;
      RECT 1978.295000  4.780000 1978.625000 5.355000 ;
      RECT 1978.555000  0.945000 1978.955000 1.295000 ;
      RECT 1978.555000  4.145000 1978.955000 4.495000 ;
      RECT 1978.820000  1.465000 1979.520000 1.505000 ;
      RECT 1978.820000  1.505000 1979.300000 1.635000 ;
      RECT 1978.820000  1.635000 1979.150000 2.465000 ;
      RECT 1978.820000  2.975000 1979.150000 3.805000 ;
      RECT 1978.820000  3.805000 1979.300000 3.935000 ;
      RECT 1978.820000  3.935000 1979.520000 3.975000 ;
      RECT 1978.860000  0.330000 1979.110000 0.585000 ;
      RECT 1978.860000  0.585000 1979.300000 0.755000 ;
      RECT 1978.860000  4.685000 1979.300000 4.855000 ;
      RECT 1978.860000  4.855000 1979.110000 5.110000 ;
      RECT 1979.130000  0.755000 1979.300000 1.175000 ;
      RECT 1979.130000  1.175000 1979.520000 1.465000 ;
      RECT 1979.130000  3.975000 1979.520000 4.265000 ;
      RECT 1979.130000  4.265000 1979.300000 4.685000 ;
      RECT 1979.340000  1.805000 1979.860000 1.985000 ;
      RECT 1979.340000  1.985000 1979.670000 2.465000 ;
      RECT 1979.340000  2.975000 1979.670000 3.455000 ;
      RECT 1979.340000  3.455000 1979.860000 3.635000 ;
      RECT 1979.465000  1.755000 1979.860000 1.805000 ;
      RECT 1979.465000  2.465000 1979.670000 2.975000 ;
      RECT 1979.465000  3.635000 1979.860000 3.685000 ;
      RECT 1979.470000  0.330000 1979.715000 0.835000 ;
      RECT 1979.470000  0.835000 1979.860000 1.005000 ;
      RECT 1979.470000  4.435000 1979.860000 4.605000 ;
      RECT 1979.470000  4.605000 1979.715000 5.110000 ;
      RECT 1979.690000  1.005000 1979.860000 1.755000 ;
      RECT 1979.690000  3.685000 1979.860000 4.435000 ;
      RECT 1979.840000  2.635000 1981.220000 2.805000 ;
      RECT 1979.925000  0.395000 1980.200000 0.625000 ;
      RECT 1979.925000  4.815000 1980.200000 5.045000 ;
      RECT 1980.030000  0.625000 1980.200000 1.055000 ;
      RECT 1980.030000  1.055000 1980.425000 1.325000 ;
      RECT 1980.030000  4.115000 1980.425000 4.385000 ;
      RECT 1980.030000  4.385000 1980.200000 4.815000 ;
      RECT 1980.335000  1.495000 1980.725000 2.635000 ;
      RECT 1980.335000  2.805000 1980.725000 3.945000 ;
      RECT 1980.370000  0.085000 1980.690000 0.885000 ;
      RECT 1980.370000  4.555000 1980.690000 5.355000 ;
      RECT 1980.635000  1.055000 1981.030000 1.325000 ;
      RECT 1980.635000  4.115000 1981.030000 4.385000 ;
      RECT 1980.860000  0.395000 1981.135000 0.625000 ;
      RECT 1980.860000  0.625000 1981.030000 1.055000 ;
      RECT 1980.860000  4.385000 1981.030000 4.815000 ;
      RECT 1980.860000  4.815000 1981.135000 5.045000 ;
      RECT 1981.200000  0.835000 1981.590000 1.005000 ;
      RECT 1981.200000  1.005000 1981.370000 1.755000 ;
      RECT 1981.200000  1.755000 1981.595000 1.805000 ;
      RECT 1981.200000  1.805000 1981.720000 1.985000 ;
      RECT 1981.200000  3.455000 1981.720000 3.635000 ;
      RECT 1981.200000  3.635000 1981.595000 3.685000 ;
      RECT 1981.200000  3.685000 1981.370000 4.435000 ;
      RECT 1981.200000  4.435000 1981.590000 4.605000 ;
      RECT 1981.345000  0.330000 1981.590000 0.835000 ;
      RECT 1981.345000  4.605000 1981.590000 5.110000 ;
      RECT 1981.390000  1.985000 1981.720000 2.465000 ;
      RECT 1981.390000  2.465000 1981.595000 2.975000 ;
      RECT 1981.390000  2.975000 1981.720000 3.455000 ;
      RECT 1981.540000  1.175000 1981.930000 1.465000 ;
      RECT 1981.540000  1.465000 1982.240000 1.505000 ;
      RECT 1981.540000  3.935000 1982.240000 3.975000 ;
      RECT 1981.540000  3.975000 1981.930000 4.265000 ;
      RECT 1981.760000  0.585000 1982.200000 0.755000 ;
      RECT 1981.760000  0.755000 1981.930000 1.175000 ;
      RECT 1981.760000  1.505000 1982.240000 1.635000 ;
      RECT 1981.760000  3.805000 1982.240000 3.935000 ;
      RECT 1981.760000  4.265000 1981.930000 4.685000 ;
      RECT 1981.760000  4.685000 1982.200000 4.855000 ;
      RECT 1981.765000  2.635000 1983.435000 2.805000 ;
      RECT 1981.910000  1.635000 1982.240000 2.465000 ;
      RECT 1981.910000  2.975000 1982.240000 3.805000 ;
      RECT 1981.950000  0.330000 1982.200000 0.585000 ;
      RECT 1981.950000  4.855000 1982.200000 5.110000 ;
      RECT 1982.105000  0.945000 1982.505000 1.295000 ;
      RECT 1982.105000  4.145000 1982.505000 4.495000 ;
      RECT 1982.435000  0.085000 1982.765000 0.660000 ;
      RECT 1982.435000  1.465000 1982.765000 2.635000 ;
      RECT 1982.435000  2.805000 1982.765000 3.975000 ;
      RECT 1982.435000  4.780000 1982.765000 5.355000 ;
      RECT 1982.695000  0.945000 1983.095000 1.295000 ;
      RECT 1982.695000  4.145000 1983.095000 4.495000 ;
      RECT 1982.960000  1.465000 1983.660000 1.505000 ;
      RECT 1982.960000  1.505000 1983.440000 1.635000 ;
      RECT 1982.960000  1.635000 1983.290000 2.465000 ;
      RECT 1982.960000  2.975000 1983.290000 3.805000 ;
      RECT 1982.960000  3.805000 1983.440000 3.935000 ;
      RECT 1982.960000  3.935000 1983.660000 3.975000 ;
      RECT 1983.000000  0.330000 1983.250000 0.585000 ;
      RECT 1983.000000  0.585000 1983.440000 0.755000 ;
      RECT 1983.000000  4.685000 1983.440000 4.855000 ;
      RECT 1983.000000  4.855000 1983.250000 5.110000 ;
      RECT 1983.270000  0.755000 1983.440000 1.175000 ;
      RECT 1983.270000  1.175000 1983.660000 1.465000 ;
      RECT 1983.270000  3.975000 1983.660000 4.265000 ;
      RECT 1983.270000  4.265000 1983.440000 4.685000 ;
      RECT 1983.480000  1.805000 1984.000000 1.985000 ;
      RECT 1983.480000  1.985000 1983.810000 2.465000 ;
      RECT 1983.480000  2.975000 1983.810000 3.455000 ;
      RECT 1983.480000  3.455000 1984.000000 3.635000 ;
      RECT 1983.605000  1.755000 1984.000000 1.805000 ;
      RECT 1983.605000  2.465000 1983.810000 2.975000 ;
      RECT 1983.605000  3.635000 1984.000000 3.685000 ;
      RECT 1983.610000  0.330000 1983.855000 0.835000 ;
      RECT 1983.610000  0.835000 1984.000000 1.005000 ;
      RECT 1983.610000  4.435000 1984.000000 4.605000 ;
      RECT 1983.610000  4.605000 1983.855000 5.110000 ;
      RECT 1983.830000  1.005000 1984.000000 1.755000 ;
      RECT 1983.830000  3.685000 1984.000000 4.435000 ;
      RECT 1983.980000  2.635000 1986.775000 2.805000 ;
      RECT 1984.065000  0.395000 1984.340000 0.625000 ;
      RECT 1984.065000  4.815000 1984.340000 5.045000 ;
      RECT 1984.170000  0.625000 1984.340000 1.055000 ;
      RECT 1984.170000  1.055000 1984.565000 1.325000 ;
      RECT 1984.170000  4.115000 1984.565000 4.385000 ;
      RECT 1984.170000  4.385000 1984.340000 4.815000 ;
      RECT 1984.475000  1.495000 1984.805000 2.635000 ;
      RECT 1984.475000  2.805000 1984.805000 3.945000 ;
      RECT 1984.510000  0.085000 1984.770000 0.885000 ;
      RECT 1984.510000  4.555000 1984.770000 5.355000 ;
      RECT 1984.985000  0.085000 1985.275000 0.810000 ;
      RECT 1984.985000  1.470000 1985.275000 2.635000 ;
      RECT 1984.985000  2.805000 1985.275000 3.970000 ;
      RECT 1984.985000  4.630000 1985.275000 5.355000 ;
      RECT 1985.455000  1.055000 1986.275000 1.325000 ;
      RECT 1985.455000  1.495000 1986.645000 1.665000 ;
      RECT 1985.455000  1.665000 1985.755000 2.210000 ;
      RECT 1985.455000  2.210000 1985.785000 2.465000 ;
      RECT 1985.455000  2.975000 1985.785000 3.230000 ;
      RECT 1985.455000  3.230000 1985.755000 3.775000 ;
      RECT 1985.455000  3.775000 1986.645000 3.945000 ;
      RECT 1985.455000  4.115000 1986.275000 4.385000 ;
      RECT 1985.505000  0.255000 1985.835000 0.715000 ;
      RECT 1985.505000  0.715000 1986.695000 0.885000 ;
      RECT 1985.505000  4.555000 1986.695000 4.725000 ;
      RECT 1985.505000  4.725000 1985.835000 5.185000 ;
      RECT 1985.925000  1.835000 1986.255000 2.105000 ;
      RECT 1985.925000  3.335000 1986.255000 3.605000 ;
      RECT 1985.955000  2.105000 1986.255000 2.635000 ;
      RECT 1985.955000  2.805000 1986.255000 3.335000 ;
      RECT 1986.005000  0.085000 1986.220000 0.545000 ;
      RECT 1986.005000  4.895000 1986.220000 5.355000 ;
      RECT 1986.390000  0.255000 1987.535000 0.425000 ;
      RECT 1986.390000  0.425000 1986.695000 0.715000 ;
      RECT 1986.390000  0.885000 1986.695000 0.925000 ;
      RECT 1986.390000  4.515000 1986.695000 4.555000 ;
      RECT 1986.390000  4.725000 1986.695000 5.015000 ;
      RECT 1986.390000  5.015000 1987.535000 5.185000 ;
      RECT 1986.475000  1.665000 1986.645000 2.295000 ;
      RECT 1986.475000  2.295000 1986.775000 2.465000 ;
      RECT 1986.475000  2.975000 1986.775000 3.145000 ;
      RECT 1986.475000  3.145000 1986.645000 3.775000 ;
      RECT 1986.825000  1.755000 1987.255000 2.125000 ;
      RECT 1986.825000  3.315000 1987.255000 3.685000 ;
      RECT 1986.865000  0.595000 1987.195000 0.885000 ;
      RECT 1986.865000  4.555000 1987.195000 4.845000 ;
      RECT 1986.945000  0.885000 1987.115000 1.755000 ;
      RECT 1986.945000  2.125000 1987.115000 3.315000 ;
      RECT 1986.945000  3.685000 1987.115000 4.555000 ;
      RECT 1987.285000  2.295000 1987.640000 2.465000 ;
      RECT 1987.285000  2.635000 1989.875000 2.805000 ;
      RECT 1987.285000  2.975000 1987.640000 3.145000 ;
      RECT 1987.365000  0.425000 1987.535000 0.770000 ;
      RECT 1987.365000  4.670000 1987.535000 5.015000 ;
      RECT 1987.460000  1.205000 1987.875000 1.305000 ;
      RECT 1987.460000  1.305000 1987.980000 1.465000 ;
      RECT 1987.460000  1.465000 1988.240000 1.475000 ;
      RECT 1987.460000  3.965000 1988.240000 3.975000 ;
      RECT 1987.460000  3.975000 1987.980000 4.135000 ;
      RECT 1987.460000  4.135000 1987.875000 4.235000 ;
      RECT 1987.470000  1.645000 1987.640000 2.295000 ;
      RECT 1987.470000  3.145000 1987.640000 3.795000 ;
      RECT 1987.705000  0.585000 1988.285000 0.755000 ;
      RECT 1987.705000  0.755000 1987.875000 1.205000 ;
      RECT 1987.705000  4.235000 1987.875000 4.685000 ;
      RECT 1987.705000  4.685000 1988.285000 4.855000 ;
      RECT 1987.810000  1.475000 1988.240000 1.635000 ;
      RECT 1987.810000  3.805000 1988.240000 3.965000 ;
      RECT 1987.910000  1.635000 1988.240000 2.465000 ;
      RECT 1987.910000  2.975000 1988.240000 3.805000 ;
      RECT 1988.035000  0.330000 1988.285000 0.585000 ;
      RECT 1988.035000  4.855000 1988.285000 5.110000 ;
      RECT 1988.150000  1.025000 1988.485000 1.295000 ;
      RECT 1988.150000  4.145000 1988.485000 4.415000 ;
      RECT 1988.415000  1.465000 1988.745000 2.635000 ;
      RECT 1988.415000  2.805000 1988.745000 3.975000 ;
      RECT 1988.455000  0.085000 1988.705000 0.660000 ;
      RECT 1988.455000  4.780000 1988.705000 5.355000 ;
      RECT 1988.675000  1.025000 1989.010000 1.295000 ;
      RECT 1988.675000  4.145000 1989.010000 4.415000 ;
      RECT 1988.875000  0.330000 1989.125000 0.585000 ;
      RECT 1988.875000  0.585000 1989.455000 0.755000 ;
      RECT 1988.875000  4.685000 1989.455000 4.855000 ;
      RECT 1988.875000  4.855000 1989.125000 5.110000 ;
      RECT 1988.920000  1.465000 1989.700000 1.475000 ;
      RECT 1988.920000  1.475000 1989.350000 1.635000 ;
      RECT 1988.920000  1.635000 1989.250000 2.465000 ;
      RECT 1988.920000  2.975000 1989.250000 3.805000 ;
      RECT 1988.920000  3.805000 1989.350000 3.965000 ;
      RECT 1988.920000  3.965000 1989.700000 3.975000 ;
      RECT 1989.180000  1.305000 1989.700000 1.465000 ;
      RECT 1989.180000  3.975000 1989.700000 4.135000 ;
      RECT 1989.285000  0.755000 1989.455000 1.205000 ;
      RECT 1989.285000  1.205000 1989.700000 1.305000 ;
      RECT 1989.285000  4.135000 1989.700000 4.235000 ;
      RECT 1989.285000  4.235000 1989.455000 4.685000 ;
      RECT 1989.520000  1.645000 1989.690000 2.295000 ;
      RECT 1989.520000  2.295000 1989.875000 2.465000 ;
      RECT 1989.520000  2.975000 1989.875000 3.145000 ;
      RECT 1989.520000  3.145000 1989.690000 3.795000 ;
      RECT 1989.625000  0.255000 1990.770000 0.425000 ;
      RECT 1989.625000  0.425000 1989.795000 0.770000 ;
      RECT 1989.625000  4.670000 1989.795000 5.015000 ;
      RECT 1989.625000  5.015000 1990.770000 5.185000 ;
      RECT 1989.905000  1.755000 1990.335000 2.125000 ;
      RECT 1989.905000  3.315000 1990.335000 3.685000 ;
      RECT 1989.965000  0.595000 1990.295000 0.885000 ;
      RECT 1989.965000  4.555000 1990.295000 4.845000 ;
      RECT 1990.045000  0.885000 1990.215000 1.755000 ;
      RECT 1990.045000  2.125000 1990.215000 3.315000 ;
      RECT 1990.045000  3.685000 1990.215000 4.555000 ;
      RECT 1990.385000  2.295000 1990.685000 2.465000 ;
      RECT 1990.385000  2.635000 1993.215000 2.805000 ;
      RECT 1990.385000  2.975000 1990.685000 3.145000 ;
      RECT 1990.465000  0.425000 1990.770000 0.715000 ;
      RECT 1990.465000  0.715000 1991.655000 0.885000 ;
      RECT 1990.465000  0.885000 1990.770000 0.925000 ;
      RECT 1990.465000  4.515000 1990.770000 4.555000 ;
      RECT 1990.465000  4.555000 1991.655000 4.725000 ;
      RECT 1990.465000  4.725000 1990.770000 5.015000 ;
      RECT 1990.515000  1.495000 1991.705000 1.665000 ;
      RECT 1990.515000  1.665000 1990.685000 2.295000 ;
      RECT 1990.515000  3.145000 1990.685000 3.775000 ;
      RECT 1990.515000  3.775000 1991.705000 3.945000 ;
      RECT 1990.885000  1.055000 1991.705000 1.325000 ;
      RECT 1990.885000  4.115000 1991.705000 4.385000 ;
      RECT 1990.905000  1.835000 1991.235000 2.105000 ;
      RECT 1990.905000  2.105000 1991.205000 2.635000 ;
      RECT 1990.905000  2.805000 1991.205000 3.335000 ;
      RECT 1990.905000  3.335000 1991.235000 3.605000 ;
      RECT 1990.940000  0.085000 1991.155000 0.545000 ;
      RECT 1990.940000  4.895000 1991.155000 5.355000 ;
      RECT 1991.325000  0.255000 1991.655000 0.715000 ;
      RECT 1991.325000  4.725000 1991.655000 5.185000 ;
      RECT 1991.375000  2.210000 1991.705000 2.465000 ;
      RECT 1991.375000  2.975000 1991.705000 3.230000 ;
      RECT 1991.405000  1.665000 1991.705000 2.210000 ;
      RECT 1991.405000  3.230000 1991.705000 3.775000 ;
      RECT 1991.895000  1.055000 1992.715000 1.325000 ;
      RECT 1991.895000  1.495000 1993.085000 1.665000 ;
      RECT 1991.895000  1.665000 1992.195000 2.210000 ;
      RECT 1991.895000  2.210000 1992.225000 2.465000 ;
      RECT 1991.895000  2.975000 1992.225000 3.230000 ;
      RECT 1991.895000  3.230000 1992.195000 3.775000 ;
      RECT 1991.895000  3.775000 1993.085000 3.945000 ;
      RECT 1991.895000  4.115000 1992.715000 4.385000 ;
      RECT 1991.945000  0.255000 1992.275000 0.715000 ;
      RECT 1991.945000  0.715000 1993.135000 0.885000 ;
      RECT 1991.945000  4.555000 1993.135000 4.725000 ;
      RECT 1991.945000  4.725000 1992.275000 5.185000 ;
      RECT 1992.365000  1.835000 1992.695000 2.105000 ;
      RECT 1992.365000  3.335000 1992.695000 3.605000 ;
      RECT 1992.395000  2.105000 1992.695000 2.635000 ;
      RECT 1992.395000  2.805000 1992.695000 3.335000 ;
      RECT 1992.445000  0.085000 1992.660000 0.545000 ;
      RECT 1992.445000  4.895000 1992.660000 5.355000 ;
      RECT 1992.830000  0.255000 1993.975000 0.425000 ;
      RECT 1992.830000  0.425000 1993.135000 0.715000 ;
      RECT 1992.830000  0.885000 1993.135000 0.925000 ;
      RECT 1992.830000  4.515000 1993.135000 4.555000 ;
      RECT 1992.830000  4.725000 1993.135000 5.015000 ;
      RECT 1992.830000  5.015000 1993.975000 5.185000 ;
      RECT 1992.915000  1.665000 1993.085000 2.295000 ;
      RECT 1992.915000  2.295000 1993.215000 2.465000 ;
      RECT 1992.915000  2.975000 1993.215000 3.145000 ;
      RECT 1992.915000  3.145000 1993.085000 3.775000 ;
      RECT 1993.265000  1.755000 1993.695000 2.125000 ;
      RECT 1993.265000  3.315000 1993.695000 3.685000 ;
      RECT 1993.305000  0.595000 1993.635000 0.885000 ;
      RECT 1993.305000  4.555000 1993.635000 4.845000 ;
      RECT 1993.385000  0.885000 1993.555000 1.755000 ;
      RECT 1993.385000  2.125000 1993.555000 3.315000 ;
      RECT 1993.385000  3.685000 1993.555000 4.555000 ;
      RECT 1993.725000  2.295000 1994.080000 2.465000 ;
      RECT 1993.725000  2.635000 1996.315000 2.805000 ;
      RECT 1993.725000  2.975000 1994.080000 3.145000 ;
      RECT 1993.805000  0.425000 1993.975000 0.770000 ;
      RECT 1993.805000  4.670000 1993.975000 5.015000 ;
      RECT 1993.900000  1.205000 1994.315000 1.305000 ;
      RECT 1993.900000  1.305000 1994.420000 1.465000 ;
      RECT 1993.900000  1.465000 1994.680000 1.475000 ;
      RECT 1993.900000  3.965000 1994.680000 3.975000 ;
      RECT 1993.900000  3.975000 1994.420000 4.135000 ;
      RECT 1993.900000  4.135000 1994.315000 4.235000 ;
      RECT 1993.910000  1.645000 1994.080000 2.295000 ;
      RECT 1993.910000  3.145000 1994.080000 3.795000 ;
      RECT 1994.145000  0.585000 1994.725000 0.755000 ;
      RECT 1994.145000  0.755000 1994.315000 1.205000 ;
      RECT 1994.145000  4.235000 1994.315000 4.685000 ;
      RECT 1994.145000  4.685000 1994.725000 4.855000 ;
      RECT 1994.250000  1.475000 1994.680000 1.635000 ;
      RECT 1994.250000  3.805000 1994.680000 3.965000 ;
      RECT 1994.350000  1.635000 1994.680000 2.465000 ;
      RECT 1994.350000  2.975000 1994.680000 3.805000 ;
      RECT 1994.475000  0.330000 1994.725000 0.585000 ;
      RECT 1994.475000  4.855000 1994.725000 5.110000 ;
      RECT 1994.590000  1.025000 1994.925000 1.295000 ;
      RECT 1994.590000  4.145000 1994.925000 4.415000 ;
      RECT 1994.855000  1.465000 1995.185000 2.635000 ;
      RECT 1994.855000  2.805000 1995.185000 3.975000 ;
      RECT 1994.895000  0.085000 1995.145000 0.660000 ;
      RECT 1994.895000  4.780000 1995.145000 5.355000 ;
      RECT 1995.115000  1.025000 1995.450000 1.295000 ;
      RECT 1995.115000  4.145000 1995.450000 4.415000 ;
      RECT 1995.315000  0.330000 1995.565000 0.585000 ;
      RECT 1995.315000  0.585000 1995.895000 0.755000 ;
      RECT 1995.315000  4.685000 1995.895000 4.855000 ;
      RECT 1995.315000  4.855000 1995.565000 5.110000 ;
      RECT 1995.360000  1.465000 1996.140000 1.475000 ;
      RECT 1995.360000  1.475000 1995.790000 1.635000 ;
      RECT 1995.360000  1.635000 1995.690000 2.465000 ;
      RECT 1995.360000  2.975000 1995.690000 3.805000 ;
      RECT 1995.360000  3.805000 1995.790000 3.965000 ;
      RECT 1995.360000  3.965000 1996.140000 3.975000 ;
      RECT 1995.620000  1.305000 1996.140000 1.465000 ;
      RECT 1995.620000  3.975000 1996.140000 4.135000 ;
      RECT 1995.725000  0.755000 1995.895000 1.205000 ;
      RECT 1995.725000  1.205000 1996.140000 1.305000 ;
      RECT 1995.725000  4.135000 1996.140000 4.235000 ;
      RECT 1995.725000  4.235000 1995.895000 4.685000 ;
      RECT 1995.960000  1.645000 1996.130000 2.295000 ;
      RECT 1995.960000  2.295000 1996.315000 2.465000 ;
      RECT 1995.960000  2.975000 1996.315000 3.145000 ;
      RECT 1995.960000  3.145000 1996.130000 3.795000 ;
      RECT 1996.065000  0.255000 1997.210000 0.425000 ;
      RECT 1996.065000  0.425000 1996.235000 0.770000 ;
      RECT 1996.065000  4.670000 1996.235000 5.015000 ;
      RECT 1996.065000  5.015000 1997.210000 5.185000 ;
      RECT 1996.345000  1.755000 1996.775000 2.125000 ;
      RECT 1996.345000  3.315000 1996.775000 3.685000 ;
      RECT 1996.405000  0.595000 1996.735000 0.885000 ;
      RECT 1996.405000  4.555000 1996.735000 4.845000 ;
      RECT 1996.485000  0.885000 1996.655000 1.755000 ;
      RECT 1996.485000  2.125000 1996.655000 3.315000 ;
      RECT 1996.485000  3.685000 1996.655000 4.555000 ;
      RECT 1996.825000  2.295000 1997.125000 2.465000 ;
      RECT 1996.825000  2.635000 1999.655000 2.805000 ;
      RECT 1996.825000  2.975000 1997.125000 3.145000 ;
      RECT 1996.905000  0.425000 1997.210000 0.715000 ;
      RECT 1996.905000  0.715000 1998.095000 0.885000 ;
      RECT 1996.905000  0.885000 1997.210000 0.925000 ;
      RECT 1996.905000  4.515000 1997.210000 4.555000 ;
      RECT 1996.905000  4.555000 1998.095000 4.725000 ;
      RECT 1996.905000  4.725000 1997.210000 5.015000 ;
      RECT 1996.955000  1.495000 1998.145000 1.665000 ;
      RECT 1996.955000  1.665000 1997.125000 2.295000 ;
      RECT 1996.955000  3.145000 1997.125000 3.775000 ;
      RECT 1996.955000  3.775000 1998.145000 3.945000 ;
      RECT 1997.325000  1.055000 1998.145000 1.325000 ;
      RECT 1997.325000  4.115000 1998.145000 4.385000 ;
      RECT 1997.345000  1.835000 1997.675000 2.105000 ;
      RECT 1997.345000  2.105000 1997.645000 2.635000 ;
      RECT 1997.345000  2.805000 1997.645000 3.335000 ;
      RECT 1997.345000  3.335000 1997.675000 3.605000 ;
      RECT 1997.380000  0.085000 1997.595000 0.545000 ;
      RECT 1997.380000  4.895000 1997.595000 5.355000 ;
      RECT 1997.765000  0.255000 1998.095000 0.715000 ;
      RECT 1997.765000  4.725000 1998.095000 5.185000 ;
      RECT 1997.815000  2.210000 1998.145000 2.465000 ;
      RECT 1997.815000  2.975000 1998.145000 3.230000 ;
      RECT 1997.845000  1.665000 1998.145000 2.210000 ;
      RECT 1997.845000  3.230000 1998.145000 3.775000 ;
      RECT 1998.335000  1.055000 1999.155000 1.325000 ;
      RECT 1998.335000  1.495000 1999.525000 1.665000 ;
      RECT 1998.335000  1.665000 1998.635000 2.210000 ;
      RECT 1998.335000  2.210000 1998.665000 2.465000 ;
      RECT 1998.335000  2.975000 1998.665000 3.230000 ;
      RECT 1998.335000  3.230000 1998.635000 3.775000 ;
      RECT 1998.335000  3.775000 1999.525000 3.945000 ;
      RECT 1998.335000  4.115000 1999.155000 4.385000 ;
      RECT 1998.385000  0.255000 1998.715000 0.715000 ;
      RECT 1998.385000  0.715000 1999.575000 0.885000 ;
      RECT 1998.385000  4.555000 1999.575000 4.725000 ;
      RECT 1998.385000  4.725000 1998.715000 5.185000 ;
      RECT 1998.805000  1.835000 1999.135000 2.105000 ;
      RECT 1998.805000  3.335000 1999.135000 3.605000 ;
      RECT 1998.835000  2.105000 1999.135000 2.635000 ;
      RECT 1998.835000  2.805000 1999.135000 3.335000 ;
      RECT 1998.885000  0.085000 1999.100000 0.545000 ;
      RECT 1998.885000  4.895000 1999.100000 5.355000 ;
      RECT 1999.270000  0.255000 2000.415000 0.425000 ;
      RECT 1999.270000  0.425000 1999.575000 0.715000 ;
      RECT 1999.270000  0.885000 1999.575000 0.925000 ;
      RECT 1999.270000  4.515000 1999.575000 4.555000 ;
      RECT 1999.270000  4.725000 1999.575000 5.015000 ;
      RECT 1999.270000  5.015000 2000.415000 5.185000 ;
      RECT 1999.355000  1.665000 1999.525000 2.295000 ;
      RECT 1999.355000  2.295000 1999.655000 2.465000 ;
      RECT 1999.355000  2.975000 1999.655000 3.145000 ;
      RECT 1999.355000  3.145000 1999.525000 3.775000 ;
      RECT 1999.705000  1.755000 2000.135000 2.125000 ;
      RECT 1999.705000  3.315000 2000.135000 3.685000 ;
      RECT 1999.745000  0.595000 2000.075000 0.885000 ;
      RECT 1999.745000  4.555000 2000.075000 4.845000 ;
      RECT 1999.825000  0.885000 1999.995000 1.755000 ;
      RECT 1999.825000  2.125000 1999.995000 3.315000 ;
      RECT 1999.825000  3.685000 1999.995000 4.555000 ;
      RECT 2000.165000  2.295000 2000.520000 2.465000 ;
      RECT 2000.165000  2.635000 2002.755000 2.805000 ;
      RECT 2000.165000  2.975000 2000.520000 3.145000 ;
      RECT 2000.245000  0.425000 2000.415000 0.770000 ;
      RECT 2000.245000  4.670000 2000.415000 5.015000 ;
      RECT 2000.340000  1.205000 2000.755000 1.305000 ;
      RECT 2000.340000  1.305000 2000.860000 1.465000 ;
      RECT 2000.340000  1.465000 2001.120000 1.475000 ;
      RECT 2000.340000  3.965000 2001.120000 3.975000 ;
      RECT 2000.340000  3.975000 2000.860000 4.135000 ;
      RECT 2000.340000  4.135000 2000.755000 4.235000 ;
      RECT 2000.350000  1.645000 2000.520000 2.295000 ;
      RECT 2000.350000  3.145000 2000.520000 3.795000 ;
      RECT 2000.585000  0.585000 2001.165000 0.755000 ;
      RECT 2000.585000  0.755000 2000.755000 1.205000 ;
      RECT 2000.585000  4.235000 2000.755000 4.685000 ;
      RECT 2000.585000  4.685000 2001.165000 4.855000 ;
      RECT 2000.690000  1.475000 2001.120000 1.635000 ;
      RECT 2000.690000  3.805000 2001.120000 3.965000 ;
      RECT 2000.790000  1.635000 2001.120000 2.465000 ;
      RECT 2000.790000  2.975000 2001.120000 3.805000 ;
      RECT 2000.915000  0.330000 2001.165000 0.585000 ;
      RECT 2000.915000  4.855000 2001.165000 5.110000 ;
      RECT 2001.030000  1.025000 2001.365000 1.295000 ;
      RECT 2001.030000  4.145000 2001.365000 4.415000 ;
      RECT 2001.295000  1.465000 2001.625000 2.635000 ;
      RECT 2001.295000  2.805000 2001.625000 3.975000 ;
      RECT 2001.335000  0.085000 2001.585000 0.660000 ;
      RECT 2001.335000  4.780000 2001.585000 5.355000 ;
      RECT 2001.555000  1.025000 2001.890000 1.295000 ;
      RECT 2001.555000  4.145000 2001.890000 4.415000 ;
      RECT 2001.755000  0.330000 2002.005000 0.585000 ;
      RECT 2001.755000  0.585000 2002.335000 0.755000 ;
      RECT 2001.755000  4.685000 2002.335000 4.855000 ;
      RECT 2001.755000  4.855000 2002.005000 5.110000 ;
      RECT 2001.800000  1.465000 2002.580000 1.475000 ;
      RECT 2001.800000  1.475000 2002.230000 1.635000 ;
      RECT 2001.800000  1.635000 2002.130000 2.465000 ;
      RECT 2001.800000  2.975000 2002.130000 3.805000 ;
      RECT 2001.800000  3.805000 2002.230000 3.965000 ;
      RECT 2001.800000  3.965000 2002.580000 3.975000 ;
      RECT 2002.060000  1.305000 2002.580000 1.465000 ;
      RECT 2002.060000  3.975000 2002.580000 4.135000 ;
      RECT 2002.165000  0.755000 2002.335000 1.205000 ;
      RECT 2002.165000  1.205000 2002.580000 1.305000 ;
      RECT 2002.165000  4.135000 2002.580000 4.235000 ;
      RECT 2002.165000  4.235000 2002.335000 4.685000 ;
      RECT 2002.400000  1.645000 2002.570000 2.295000 ;
      RECT 2002.400000  2.295000 2002.755000 2.465000 ;
      RECT 2002.400000  2.975000 2002.755000 3.145000 ;
      RECT 2002.400000  3.145000 2002.570000 3.795000 ;
      RECT 2002.505000  0.255000 2003.650000 0.425000 ;
      RECT 2002.505000  0.425000 2002.675000 0.770000 ;
      RECT 2002.505000  4.670000 2002.675000 5.015000 ;
      RECT 2002.505000  5.015000 2003.650000 5.185000 ;
      RECT 2002.785000  1.755000 2003.215000 2.125000 ;
      RECT 2002.785000  3.315000 2003.215000 3.685000 ;
      RECT 2002.845000  0.595000 2003.175000 0.885000 ;
      RECT 2002.845000  4.555000 2003.175000 4.845000 ;
      RECT 2002.925000  0.885000 2003.095000 1.755000 ;
      RECT 2002.925000  2.125000 2003.095000 3.315000 ;
      RECT 2002.925000  3.685000 2003.095000 4.555000 ;
      RECT 2003.265000  2.295000 2003.565000 2.465000 ;
      RECT 2003.265000  2.635000 2006.095000 2.805000 ;
      RECT 2003.265000  2.975000 2003.565000 3.145000 ;
      RECT 2003.345000  0.425000 2003.650000 0.715000 ;
      RECT 2003.345000  0.715000 2004.535000 0.885000 ;
      RECT 2003.345000  0.885000 2003.650000 0.925000 ;
      RECT 2003.345000  4.515000 2003.650000 4.555000 ;
      RECT 2003.345000  4.555000 2004.535000 4.725000 ;
      RECT 2003.345000  4.725000 2003.650000 5.015000 ;
      RECT 2003.395000  1.495000 2004.585000 1.665000 ;
      RECT 2003.395000  1.665000 2003.565000 2.295000 ;
      RECT 2003.395000  3.145000 2003.565000 3.775000 ;
      RECT 2003.395000  3.775000 2004.585000 3.945000 ;
      RECT 2003.765000  1.055000 2004.585000 1.325000 ;
      RECT 2003.765000  4.115000 2004.585000 4.385000 ;
      RECT 2003.785000  1.835000 2004.115000 2.105000 ;
      RECT 2003.785000  2.105000 2004.085000 2.635000 ;
      RECT 2003.785000  2.805000 2004.085000 3.335000 ;
      RECT 2003.785000  3.335000 2004.115000 3.605000 ;
      RECT 2003.820000  0.085000 2004.035000 0.545000 ;
      RECT 2003.820000  4.895000 2004.035000 5.355000 ;
      RECT 2004.205000  0.255000 2004.535000 0.715000 ;
      RECT 2004.205000  4.725000 2004.535000 5.185000 ;
      RECT 2004.255000  2.210000 2004.585000 2.465000 ;
      RECT 2004.255000  2.975000 2004.585000 3.230000 ;
      RECT 2004.285000  1.665000 2004.585000 2.210000 ;
      RECT 2004.285000  3.230000 2004.585000 3.775000 ;
      RECT 2004.775000  1.055000 2005.595000 1.325000 ;
      RECT 2004.775000  1.495000 2005.965000 1.665000 ;
      RECT 2004.775000  1.665000 2005.075000 2.210000 ;
      RECT 2004.775000  2.210000 2005.105000 2.465000 ;
      RECT 2004.775000  2.975000 2005.105000 3.230000 ;
      RECT 2004.775000  3.230000 2005.075000 3.775000 ;
      RECT 2004.775000  3.775000 2005.965000 3.945000 ;
      RECT 2004.775000  4.115000 2005.595000 4.385000 ;
      RECT 2004.825000  0.255000 2005.155000 0.715000 ;
      RECT 2004.825000  0.715000 2006.015000 0.885000 ;
      RECT 2004.825000  4.555000 2006.015000 4.725000 ;
      RECT 2004.825000  4.725000 2005.155000 5.185000 ;
      RECT 2005.245000  1.835000 2005.575000 2.105000 ;
      RECT 2005.245000  3.335000 2005.575000 3.605000 ;
      RECT 2005.275000  2.105000 2005.575000 2.635000 ;
      RECT 2005.275000  2.805000 2005.575000 3.335000 ;
      RECT 2005.325000  0.085000 2005.540000 0.545000 ;
      RECT 2005.325000  4.895000 2005.540000 5.355000 ;
      RECT 2005.710000  0.255000 2006.855000 0.425000 ;
      RECT 2005.710000  0.425000 2006.015000 0.715000 ;
      RECT 2005.710000  0.885000 2006.015000 0.925000 ;
      RECT 2005.710000  4.515000 2006.015000 4.555000 ;
      RECT 2005.710000  4.725000 2006.015000 5.015000 ;
      RECT 2005.710000  5.015000 2006.855000 5.185000 ;
      RECT 2005.795000  1.665000 2005.965000 2.295000 ;
      RECT 2005.795000  2.295000 2006.095000 2.465000 ;
      RECT 2005.795000  2.975000 2006.095000 3.145000 ;
      RECT 2005.795000  3.145000 2005.965000 3.775000 ;
      RECT 2006.145000  1.755000 2006.575000 2.125000 ;
      RECT 2006.145000  3.315000 2006.575000 3.685000 ;
      RECT 2006.185000  0.595000 2006.515000 0.885000 ;
      RECT 2006.185000  4.555000 2006.515000 4.845000 ;
      RECT 2006.265000  0.885000 2006.435000 1.755000 ;
      RECT 2006.265000  2.125000 2006.435000 3.315000 ;
      RECT 2006.265000  3.685000 2006.435000 4.555000 ;
      RECT 2006.605000  2.295000 2006.960000 2.465000 ;
      RECT 2006.605000  2.635000 2009.195000 2.805000 ;
      RECT 2006.605000  2.975000 2006.960000 3.145000 ;
      RECT 2006.685000  0.425000 2006.855000 0.770000 ;
      RECT 2006.685000  4.670000 2006.855000 5.015000 ;
      RECT 2006.780000  1.205000 2007.195000 1.305000 ;
      RECT 2006.780000  1.305000 2007.300000 1.465000 ;
      RECT 2006.780000  1.465000 2007.560000 1.475000 ;
      RECT 2006.780000  3.965000 2007.560000 3.975000 ;
      RECT 2006.780000  3.975000 2007.300000 4.135000 ;
      RECT 2006.780000  4.135000 2007.195000 4.235000 ;
      RECT 2006.790000  1.645000 2006.960000 2.295000 ;
      RECT 2006.790000  3.145000 2006.960000 3.795000 ;
      RECT 2007.025000  0.585000 2007.605000 0.755000 ;
      RECT 2007.025000  0.755000 2007.195000 1.205000 ;
      RECT 2007.025000  4.235000 2007.195000 4.685000 ;
      RECT 2007.025000  4.685000 2007.605000 4.855000 ;
      RECT 2007.130000  1.475000 2007.560000 1.635000 ;
      RECT 2007.130000  3.805000 2007.560000 3.965000 ;
      RECT 2007.230000  1.635000 2007.560000 2.465000 ;
      RECT 2007.230000  2.975000 2007.560000 3.805000 ;
      RECT 2007.355000  0.330000 2007.605000 0.585000 ;
      RECT 2007.355000  4.855000 2007.605000 5.110000 ;
      RECT 2007.470000  1.025000 2007.805000 1.295000 ;
      RECT 2007.470000  4.145000 2007.805000 4.415000 ;
      RECT 2007.735000  1.465000 2008.065000 2.635000 ;
      RECT 2007.735000  2.805000 2008.065000 3.975000 ;
      RECT 2007.775000  0.085000 2008.025000 0.660000 ;
      RECT 2007.775000  4.780000 2008.025000 5.355000 ;
      RECT 2007.995000  1.025000 2008.330000 1.295000 ;
      RECT 2007.995000  4.145000 2008.330000 4.415000 ;
      RECT 2008.195000  0.330000 2008.445000 0.585000 ;
      RECT 2008.195000  0.585000 2008.775000 0.755000 ;
      RECT 2008.195000  4.685000 2008.775000 4.855000 ;
      RECT 2008.195000  4.855000 2008.445000 5.110000 ;
      RECT 2008.240000  1.465000 2009.020000 1.475000 ;
      RECT 2008.240000  1.475000 2008.670000 1.635000 ;
      RECT 2008.240000  1.635000 2008.570000 2.465000 ;
      RECT 2008.240000  2.975000 2008.570000 3.805000 ;
      RECT 2008.240000  3.805000 2008.670000 3.965000 ;
      RECT 2008.240000  3.965000 2009.020000 3.975000 ;
      RECT 2008.500000  1.305000 2009.020000 1.465000 ;
      RECT 2008.500000  3.975000 2009.020000 4.135000 ;
      RECT 2008.605000  0.755000 2008.775000 1.205000 ;
      RECT 2008.605000  1.205000 2009.020000 1.305000 ;
      RECT 2008.605000  4.135000 2009.020000 4.235000 ;
      RECT 2008.605000  4.235000 2008.775000 4.685000 ;
      RECT 2008.840000  1.645000 2009.010000 2.295000 ;
      RECT 2008.840000  2.295000 2009.195000 2.465000 ;
      RECT 2008.840000  2.975000 2009.195000 3.145000 ;
      RECT 2008.840000  3.145000 2009.010000 3.795000 ;
      RECT 2008.945000  0.255000 2010.090000 0.425000 ;
      RECT 2008.945000  0.425000 2009.115000 0.770000 ;
      RECT 2008.945000  4.670000 2009.115000 5.015000 ;
      RECT 2008.945000  5.015000 2010.090000 5.185000 ;
      RECT 2009.225000  1.755000 2009.655000 2.125000 ;
      RECT 2009.225000  3.315000 2009.655000 3.685000 ;
      RECT 2009.285000  0.595000 2009.615000 0.885000 ;
      RECT 2009.285000  4.555000 2009.615000 4.845000 ;
      RECT 2009.365000  0.885000 2009.535000 1.755000 ;
      RECT 2009.365000  2.125000 2009.535000 3.315000 ;
      RECT 2009.365000  3.685000 2009.535000 4.555000 ;
      RECT 2009.705000  2.295000 2010.005000 2.465000 ;
      RECT 2009.705000  2.635000 2014.375000 2.805000 ;
      RECT 2009.705000  2.975000 2010.005000 3.145000 ;
      RECT 2009.785000  0.425000 2010.090000 0.715000 ;
      RECT 2009.785000  0.715000 2010.975000 0.885000 ;
      RECT 2009.785000  0.885000 2010.090000 0.925000 ;
      RECT 2009.785000  4.515000 2010.090000 4.555000 ;
      RECT 2009.785000  4.555000 2010.975000 4.725000 ;
      RECT 2009.785000  4.725000 2010.090000 5.015000 ;
      RECT 2009.835000  1.495000 2011.025000 1.665000 ;
      RECT 2009.835000  1.665000 2010.005000 2.295000 ;
      RECT 2009.835000  3.145000 2010.005000 3.775000 ;
      RECT 2009.835000  3.775000 2011.025000 3.945000 ;
      RECT 2010.205000  1.055000 2011.025000 1.325000 ;
      RECT 2010.205000  4.115000 2011.025000 4.385000 ;
      RECT 2010.225000  1.835000 2010.555000 2.105000 ;
      RECT 2010.225000  2.105000 2010.525000 2.635000 ;
      RECT 2010.225000  2.805000 2010.525000 3.335000 ;
      RECT 2010.225000  3.335000 2010.555000 3.605000 ;
      RECT 2010.260000  0.085000 2010.475000 0.545000 ;
      RECT 2010.260000  4.895000 2010.475000 5.355000 ;
      RECT 2010.645000  0.255000 2010.975000 0.715000 ;
      RECT 2010.645000  4.725000 2010.975000 5.185000 ;
      RECT 2010.695000  2.210000 2011.025000 2.465000 ;
      RECT 2010.695000  2.975000 2011.025000 3.230000 ;
      RECT 2010.725000  1.665000 2011.025000 2.210000 ;
      RECT 2010.725000  3.230000 2011.025000 3.775000 ;
      RECT 2011.205000  0.085000 2011.495000 0.810000 ;
      RECT 2011.205000  1.470000 2011.495000 2.635000 ;
      RECT 2011.205000  2.805000 2011.495000 3.970000 ;
      RECT 2011.205000  4.630000 2011.495000 5.355000 ;
      RECT 2011.705000  1.495000 2011.975000 2.635000 ;
      RECT 2011.705000  2.805000 2011.975000 3.945000 ;
      RECT 2011.725000  0.085000 2011.975000 0.885000 ;
      RECT 2011.725000  4.555000 2011.975000 5.355000 ;
      RECT 2011.975000  1.055000 2013.365000 1.325000 ;
      RECT 2011.975000  4.115000 2013.365000 4.385000 ;
      RECT 2012.145000  0.255000 2012.475000 0.715000 ;
      RECT 2012.145000  0.715000 2014.275000 0.885000 ;
      RECT 2012.145000  1.495000 2014.375000 1.665000 ;
      RECT 2012.145000  1.665000 2012.475000 2.465000 ;
      RECT 2012.145000  2.975000 2012.475000 3.775000 ;
      RECT 2012.145000  3.775000 2014.375000 3.945000 ;
      RECT 2012.145000  4.555000 2014.275000 4.725000 ;
      RECT 2012.145000  4.725000 2012.475000 5.185000 ;
      RECT 2012.645000  0.085000 2012.915000 0.545000 ;
      RECT 2012.645000  1.835000 2012.915000 2.635000 ;
      RECT 2012.645000  2.805000 2012.915000 3.605000 ;
      RECT 2012.645000  4.895000 2012.915000 5.355000 ;
      RECT 2013.085000  0.255000 2013.415000 0.715000 ;
      RECT 2013.085000  1.665000 2013.415000 2.465000 ;
      RECT 2013.085000  2.975000 2013.415000 3.775000 ;
      RECT 2013.085000  4.725000 2013.415000 5.185000 ;
      RECT 2013.585000  0.085000 2013.835000 0.545000 ;
      RECT 2013.585000  1.835000 2013.855000 2.635000 ;
      RECT 2013.585000  2.805000 2013.855000 3.605000 ;
      RECT 2013.585000  4.895000 2013.835000 5.355000 ;
      RECT 2014.005000  0.255000 2016.035000 0.425000 ;
      RECT 2014.005000  0.425000 2014.275000 0.715000 ;
      RECT 2014.005000  4.725000 2014.275000 5.015000 ;
      RECT 2014.005000  5.015000 2016.035000 5.185000 ;
      RECT 2014.075000  1.665000 2014.375000 2.465000 ;
      RECT 2014.075000  2.975000 2014.375000 3.775000 ;
      RECT 2014.445000  0.595000 2014.775000 0.885000 ;
      RECT 2014.445000  4.555000 2014.775000 4.845000 ;
      RECT 2014.545000  0.885000 2014.775000 1.065000 ;
      RECT 2014.545000  1.065000 2015.815000 1.365000 ;
      RECT 2014.545000  1.365000 2014.875000 4.075000 ;
      RECT 2014.545000  4.075000 2015.815000 4.375000 ;
      RECT 2014.545000  4.375000 2014.775000 4.555000 ;
      RECT 2014.945000  0.425000 2015.115000 0.770000 ;
      RECT 2014.945000  4.670000 2015.115000 5.015000 ;
      RECT 2015.045000  1.535000 2015.315000 2.465000 ;
      RECT 2015.045000  2.975000 2015.315000 3.905000 ;
      RECT 2015.285000  0.595000 2015.615000 1.065000 ;
      RECT 2015.285000  4.375000 2015.615000 4.845000 ;
      RECT 2015.485000  1.365000 2015.815000 4.075000 ;
      RECT 2015.785000  0.425000 2016.035000 0.770000 ;
      RECT 2015.785000  4.670000 2016.035000 5.015000 ;
      RECT 2015.985000  1.065000 2017.170000 1.395000 ;
      RECT 2015.985000  1.565000 2016.285000 2.465000 ;
      RECT 2015.985000  2.635000 2020.055000 2.805000 ;
      RECT 2015.985000  2.975000 2016.285000 3.875000 ;
      RECT 2015.985000  4.045000 2017.170000 4.375000 ;
      RECT 2016.530000  1.605000 2016.805000 2.635000 ;
      RECT 2016.530000  2.805000 2016.805000 3.835000 ;
      RECT 2016.540000  0.085000 2016.830000 0.610000 ;
      RECT 2016.540000  4.830000 2016.830000 5.355000 ;
      RECT 2017.000000  0.280000 2017.250000 0.825000 ;
      RECT 2017.000000  0.825000 2017.170000 1.065000 ;
      RECT 2017.000000  1.395000 2017.170000 1.605000 ;
      RECT 2017.000000  1.605000 2017.330000 2.465000 ;
      RECT 2017.000000  2.975000 2017.330000 3.835000 ;
      RECT 2017.000000  3.835000 2017.170000 4.045000 ;
      RECT 2017.000000  4.375000 2017.170000 4.615000 ;
      RECT 2017.000000  4.615000 2017.250000 5.160000 ;
      RECT 2017.340000  0.995000 2017.935000 1.325000 ;
      RECT 2017.340000  4.115000 2017.935000 4.445000 ;
      RECT 2017.460000  0.085000 2017.750000 0.610000 ;
      RECT 2017.460000  4.830000 2017.750000 5.355000 ;
      RECT 2017.500000  1.605000 2017.800000 2.635000 ;
      RECT 2017.500000  2.805000 2017.800000 3.835000 ;
      RECT 2018.105000  0.995000 2018.700000 1.325000 ;
      RECT 2018.105000  4.115000 2018.700000 4.445000 ;
      RECT 2018.240000  1.605000 2018.540000 2.635000 ;
      RECT 2018.240000  2.805000 2018.540000 3.835000 ;
      RECT 2018.290000  0.085000 2018.580000 0.610000 ;
      RECT 2018.290000  4.830000 2018.580000 5.355000 ;
      RECT 2018.710000  1.605000 2019.040000 2.465000 ;
      RECT 2018.710000  2.975000 2019.040000 3.835000 ;
      RECT 2018.790000  0.280000 2019.040000 0.825000 ;
      RECT 2018.790000  4.615000 2019.040000 5.160000 ;
      RECT 2018.870000  0.825000 2019.040000 1.065000 ;
      RECT 2018.870000  1.065000 2020.055000 1.395000 ;
      RECT 2018.870000  1.395000 2019.040000 1.605000 ;
      RECT 2018.870000  3.835000 2019.040000 4.045000 ;
      RECT 2018.870000  4.045000 2020.055000 4.375000 ;
      RECT 2018.870000  4.375000 2019.040000 4.615000 ;
      RECT 2019.210000  0.085000 2019.500000 0.610000 ;
      RECT 2019.210000  4.830000 2019.500000 5.355000 ;
      RECT 2019.235000  1.605000 2019.510000 2.635000 ;
      RECT 2019.235000  2.805000 2019.510000 3.835000 ;
      RECT 2019.755000  1.565000 2020.055000 2.465000 ;
      RECT 2019.755000  2.975000 2020.055000 3.875000 ;
      RECT 2020.005000  0.255000 2022.035000 0.425000 ;
      RECT 2020.005000  0.425000 2020.255000 0.770000 ;
      RECT 2020.005000  4.670000 2020.255000 5.015000 ;
      RECT 2020.005000  5.015000 2022.035000 5.185000 ;
      RECT 2020.225000  1.065000 2021.495000 1.365000 ;
      RECT 2020.225000  1.365000 2020.555000 4.075000 ;
      RECT 2020.225000  4.075000 2021.495000 4.375000 ;
      RECT 2020.425000  0.595000 2020.755000 1.065000 ;
      RECT 2020.425000  4.375000 2020.755000 4.845000 ;
      RECT 2020.725000  1.535000 2020.995000 2.465000 ;
      RECT 2020.725000  2.975000 2020.995000 3.905000 ;
      RECT 2020.925000  0.425000 2021.095000 0.770000 ;
      RECT 2020.925000  4.670000 2021.095000 5.015000 ;
      RECT 2021.165000  1.365000 2021.495000 4.075000 ;
      RECT 2021.265000  0.595000 2021.595000 0.885000 ;
      RECT 2021.265000  0.885000 2021.495000 1.065000 ;
      RECT 2021.265000  4.375000 2021.495000 4.555000 ;
      RECT 2021.265000  4.555000 2021.595000 4.845000 ;
      RECT 2021.665000  1.495000 2023.895000 1.665000 ;
      RECT 2021.665000  1.665000 2021.965000 2.465000 ;
      RECT 2021.665000  2.635000 2027.255000 2.805000 ;
      RECT 2021.665000  2.975000 2021.965000 3.775000 ;
      RECT 2021.665000  3.775000 2023.895000 3.945000 ;
      RECT 2021.765000  0.425000 2022.035000 0.715000 ;
      RECT 2021.765000  0.715000 2023.895000 0.885000 ;
      RECT 2021.765000  4.555000 2023.895000 4.725000 ;
      RECT 2021.765000  4.725000 2022.035000 5.015000 ;
      RECT 2022.185000  1.835000 2022.455000 2.635000 ;
      RECT 2022.185000  2.805000 2022.455000 3.605000 ;
      RECT 2022.205000  0.085000 2022.455000 0.545000 ;
      RECT 2022.205000  4.895000 2022.455000 5.355000 ;
      RECT 2022.625000  0.255000 2022.955000 0.715000 ;
      RECT 2022.625000  1.665000 2022.955000 2.465000 ;
      RECT 2022.625000  2.975000 2022.955000 3.775000 ;
      RECT 2022.625000  4.725000 2022.955000 5.185000 ;
      RECT 2022.675000  1.055000 2024.065000 1.325000 ;
      RECT 2022.675000  4.115000 2024.065000 4.385000 ;
      RECT 2023.125000  0.085000 2023.395000 0.545000 ;
      RECT 2023.125000  1.835000 2023.395000 2.635000 ;
      RECT 2023.125000  2.805000 2023.395000 3.605000 ;
      RECT 2023.125000  4.895000 2023.395000 5.355000 ;
      RECT 2023.565000  0.255000 2023.895000 0.715000 ;
      RECT 2023.565000  1.665000 2023.895000 2.465000 ;
      RECT 2023.565000  2.975000 2023.895000 3.775000 ;
      RECT 2023.565000  4.725000 2023.895000 5.185000 ;
      RECT 2024.065000  0.085000 2024.315000 0.885000 ;
      RECT 2024.065000  1.495000 2024.335000 2.635000 ;
      RECT 2024.065000  2.805000 2024.335000 3.945000 ;
      RECT 2024.065000  4.555000 2024.315000 5.355000 ;
      RECT 2024.585000  1.495000 2024.855000 2.635000 ;
      RECT 2024.585000  2.805000 2024.855000 3.945000 ;
      RECT 2024.605000  0.085000 2024.855000 0.885000 ;
      RECT 2024.605000  4.555000 2024.855000 5.355000 ;
      RECT 2024.855000  1.055000 2026.245000 1.325000 ;
      RECT 2024.855000  4.115000 2026.245000 4.385000 ;
      RECT 2025.025000  0.255000 2025.355000 0.715000 ;
      RECT 2025.025000  0.715000 2027.155000 0.885000 ;
      RECT 2025.025000  1.495000 2027.255000 1.665000 ;
      RECT 2025.025000  1.665000 2025.355000 2.465000 ;
      RECT 2025.025000  2.975000 2025.355000 3.775000 ;
      RECT 2025.025000  3.775000 2027.255000 3.945000 ;
      RECT 2025.025000  4.555000 2027.155000 4.725000 ;
      RECT 2025.025000  4.725000 2025.355000 5.185000 ;
      RECT 2025.525000  0.085000 2025.795000 0.545000 ;
      RECT 2025.525000  1.835000 2025.795000 2.635000 ;
      RECT 2025.525000  2.805000 2025.795000 3.605000 ;
      RECT 2025.525000  4.895000 2025.795000 5.355000 ;
      RECT 2025.965000  0.255000 2026.295000 0.715000 ;
      RECT 2025.965000  1.665000 2026.295000 2.465000 ;
      RECT 2025.965000  2.975000 2026.295000 3.775000 ;
      RECT 2025.965000  4.725000 2026.295000 5.185000 ;
      RECT 2026.465000  0.085000 2026.715000 0.545000 ;
      RECT 2026.465000  1.835000 2026.735000 2.635000 ;
      RECT 2026.465000  2.805000 2026.735000 3.605000 ;
      RECT 2026.465000  4.895000 2026.715000 5.355000 ;
      RECT 2026.885000  0.255000 2028.915000 0.425000 ;
      RECT 2026.885000  0.425000 2027.155000 0.715000 ;
      RECT 2026.885000  4.725000 2027.155000 5.015000 ;
      RECT 2026.885000  5.015000 2028.915000 5.185000 ;
      RECT 2026.955000  1.665000 2027.255000 2.465000 ;
      RECT 2026.955000  2.975000 2027.255000 3.775000 ;
      RECT 2027.325000  0.595000 2027.655000 0.885000 ;
      RECT 2027.325000  4.555000 2027.655000 4.845000 ;
      RECT 2027.425000  0.885000 2027.655000 1.065000 ;
      RECT 2027.425000  1.065000 2028.695000 1.365000 ;
      RECT 2027.425000  1.365000 2027.755000 4.075000 ;
      RECT 2027.425000  4.075000 2028.695000 4.375000 ;
      RECT 2027.425000  4.375000 2027.655000 4.555000 ;
      RECT 2027.825000  0.425000 2027.995000 0.770000 ;
      RECT 2027.825000  4.670000 2027.995000 5.015000 ;
      RECT 2027.925000  1.535000 2028.195000 2.465000 ;
      RECT 2027.925000  2.975000 2028.195000 3.905000 ;
      RECT 2028.165000  0.595000 2028.495000 1.065000 ;
      RECT 2028.165000  4.375000 2028.495000 4.845000 ;
      RECT 2028.365000  1.365000 2028.695000 4.075000 ;
      RECT 2028.665000  0.425000 2028.915000 0.770000 ;
      RECT 2028.665000  4.670000 2028.915000 5.015000 ;
      RECT 2028.865000  1.065000 2030.050000 1.395000 ;
      RECT 2028.865000  1.565000 2029.165000 2.465000 ;
      RECT 2028.865000  2.635000 2032.935000 2.805000 ;
      RECT 2028.865000  2.975000 2029.165000 3.875000 ;
      RECT 2028.865000  4.045000 2030.050000 4.375000 ;
      RECT 2029.410000  1.605000 2029.685000 2.635000 ;
      RECT 2029.410000  2.805000 2029.685000 3.835000 ;
      RECT 2029.420000  0.085000 2029.710000 0.610000 ;
      RECT 2029.420000  4.830000 2029.710000 5.355000 ;
      RECT 2029.880000  0.280000 2030.130000 0.825000 ;
      RECT 2029.880000  0.825000 2030.050000 1.065000 ;
      RECT 2029.880000  1.395000 2030.050000 1.605000 ;
      RECT 2029.880000  1.605000 2030.210000 2.465000 ;
      RECT 2029.880000  2.975000 2030.210000 3.835000 ;
      RECT 2029.880000  3.835000 2030.050000 4.045000 ;
      RECT 2029.880000  4.375000 2030.050000 4.615000 ;
      RECT 2029.880000  4.615000 2030.130000 5.160000 ;
      RECT 2030.220000  0.995000 2030.815000 1.325000 ;
      RECT 2030.220000  4.115000 2030.815000 4.445000 ;
      RECT 2030.340000  0.085000 2030.630000 0.610000 ;
      RECT 2030.340000  4.830000 2030.630000 5.355000 ;
      RECT 2030.380000  1.605000 2030.680000 2.635000 ;
      RECT 2030.380000  2.805000 2030.680000 3.835000 ;
      RECT 2030.985000  0.995000 2031.580000 1.325000 ;
      RECT 2030.985000  4.115000 2031.580000 4.445000 ;
      RECT 2031.120000  1.605000 2031.420000 2.635000 ;
      RECT 2031.120000  2.805000 2031.420000 3.835000 ;
      RECT 2031.170000  0.085000 2031.460000 0.610000 ;
      RECT 2031.170000  4.830000 2031.460000 5.355000 ;
      RECT 2031.590000  1.605000 2031.920000 2.465000 ;
      RECT 2031.590000  2.975000 2031.920000 3.835000 ;
      RECT 2031.670000  0.280000 2031.920000 0.825000 ;
      RECT 2031.670000  4.615000 2031.920000 5.160000 ;
      RECT 2031.750000  0.825000 2031.920000 1.065000 ;
      RECT 2031.750000  1.065000 2032.935000 1.395000 ;
      RECT 2031.750000  1.395000 2031.920000 1.605000 ;
      RECT 2031.750000  3.835000 2031.920000 4.045000 ;
      RECT 2031.750000  4.045000 2032.935000 4.375000 ;
      RECT 2031.750000  4.375000 2031.920000 4.615000 ;
      RECT 2032.090000  0.085000 2032.380000 0.610000 ;
      RECT 2032.090000  4.830000 2032.380000 5.355000 ;
      RECT 2032.115000  1.605000 2032.390000 2.635000 ;
      RECT 2032.115000  2.805000 2032.390000 3.835000 ;
      RECT 2032.635000  1.565000 2032.935000 2.465000 ;
      RECT 2032.635000  2.975000 2032.935000 3.875000 ;
      RECT 2032.885000  0.255000 2034.915000 0.425000 ;
      RECT 2032.885000  0.425000 2033.135000 0.770000 ;
      RECT 2032.885000  4.670000 2033.135000 5.015000 ;
      RECT 2032.885000  5.015000 2034.915000 5.185000 ;
      RECT 2033.105000  1.065000 2034.375000 1.365000 ;
      RECT 2033.105000  1.365000 2033.435000 4.075000 ;
      RECT 2033.105000  4.075000 2034.375000 4.375000 ;
      RECT 2033.305000  0.595000 2033.635000 1.065000 ;
      RECT 2033.305000  4.375000 2033.635000 4.845000 ;
      RECT 2033.605000  1.535000 2033.875000 2.465000 ;
      RECT 2033.605000  2.975000 2033.875000 3.905000 ;
      RECT 2033.805000  0.425000 2033.975000 0.770000 ;
      RECT 2033.805000  4.670000 2033.975000 5.015000 ;
      RECT 2034.045000  1.365000 2034.375000 4.075000 ;
      RECT 2034.145000  0.595000 2034.475000 0.885000 ;
      RECT 2034.145000  0.885000 2034.375000 1.065000 ;
      RECT 2034.145000  4.375000 2034.375000 4.555000 ;
      RECT 2034.145000  4.555000 2034.475000 4.845000 ;
      RECT 2034.545000  1.495000 2036.775000 1.665000 ;
      RECT 2034.545000  1.665000 2034.845000 2.465000 ;
      RECT 2034.545000  2.635000 2040.595000 2.805000 ;
      RECT 2034.545000  2.975000 2034.845000 3.775000 ;
      RECT 2034.545000  3.775000 2036.775000 3.945000 ;
      RECT 2034.645000  0.425000 2034.915000 0.715000 ;
      RECT 2034.645000  0.715000 2036.775000 0.885000 ;
      RECT 2034.645000  4.555000 2036.775000 4.725000 ;
      RECT 2034.645000  4.725000 2034.915000 5.015000 ;
      RECT 2035.065000  1.835000 2035.335000 2.635000 ;
      RECT 2035.065000  2.805000 2035.335000 3.605000 ;
      RECT 2035.085000  0.085000 2035.335000 0.545000 ;
      RECT 2035.085000  4.895000 2035.335000 5.355000 ;
      RECT 2035.505000  0.255000 2035.835000 0.715000 ;
      RECT 2035.505000  1.665000 2035.835000 2.465000 ;
      RECT 2035.505000  2.975000 2035.835000 3.775000 ;
      RECT 2035.505000  4.725000 2035.835000 5.185000 ;
      RECT 2035.555000  1.055000 2036.945000 1.325000 ;
      RECT 2035.555000  4.115000 2036.945000 4.385000 ;
      RECT 2036.005000  0.085000 2036.275000 0.545000 ;
      RECT 2036.005000  1.835000 2036.275000 2.635000 ;
      RECT 2036.005000  2.805000 2036.275000 3.605000 ;
      RECT 2036.005000  4.895000 2036.275000 5.355000 ;
      RECT 2036.445000  0.255000 2036.775000 0.715000 ;
      RECT 2036.445000  1.665000 2036.775000 2.465000 ;
      RECT 2036.445000  2.975000 2036.775000 3.775000 ;
      RECT 2036.445000  4.725000 2036.775000 5.185000 ;
      RECT 2036.945000  0.085000 2037.195000 0.885000 ;
      RECT 2036.945000  1.495000 2037.215000 2.635000 ;
      RECT 2036.945000  2.805000 2037.215000 3.945000 ;
      RECT 2036.945000  4.555000 2037.195000 5.355000 ;
      RECT 2037.425000  0.085000 2037.715000 0.810000 ;
      RECT 2037.425000  1.470000 2037.715000 2.635000 ;
      RECT 2037.425000  2.805000 2037.715000 3.970000 ;
      RECT 2037.425000  4.630000 2037.715000 5.355000 ;
      RECT 2037.925000  1.495000 2038.195000 2.635000 ;
      RECT 2037.925000  2.805000 2038.195000 3.945000 ;
      RECT 2037.945000  0.085000 2038.195000 0.885000 ;
      RECT 2037.945000  4.555000 2038.195000 5.355000 ;
      RECT 2038.195000  1.055000 2039.585000 1.325000 ;
      RECT 2038.195000  4.115000 2039.585000 4.385000 ;
      RECT 2038.365000  0.255000 2038.695000 0.715000 ;
      RECT 2038.365000  0.715000 2040.495000 0.885000 ;
      RECT 2038.365000  1.495000 2040.595000 1.665000 ;
      RECT 2038.365000  1.665000 2038.695000 2.465000 ;
      RECT 2038.365000  2.975000 2038.695000 3.775000 ;
      RECT 2038.365000  3.775000 2040.595000 3.945000 ;
      RECT 2038.365000  4.555000 2040.495000 4.725000 ;
      RECT 2038.365000  4.725000 2038.695000 5.185000 ;
      RECT 2038.865000  0.085000 2039.135000 0.545000 ;
      RECT 2038.865000  1.835000 2039.135000 2.635000 ;
      RECT 2038.865000  2.805000 2039.135000 3.605000 ;
      RECT 2038.865000  4.895000 2039.135000 5.355000 ;
      RECT 2039.305000  0.255000 2039.635000 0.715000 ;
      RECT 2039.305000  1.665000 2039.635000 2.465000 ;
      RECT 2039.305000  2.975000 2039.635000 3.775000 ;
      RECT 2039.305000  4.725000 2039.635000 5.185000 ;
      RECT 2039.805000  0.085000 2040.055000 0.545000 ;
      RECT 2039.805000  1.835000 2040.075000 2.635000 ;
      RECT 2039.805000  2.805000 2040.075000 3.605000 ;
      RECT 2039.805000  4.895000 2040.055000 5.355000 ;
      RECT 2040.225000  0.255000 2042.255000 0.425000 ;
      RECT 2040.225000  0.425000 2040.495000 0.715000 ;
      RECT 2040.225000  4.725000 2040.495000 5.015000 ;
      RECT 2040.225000  5.015000 2042.255000 5.185000 ;
      RECT 2040.295000  1.665000 2040.595000 2.465000 ;
      RECT 2040.295000  2.975000 2040.595000 3.775000 ;
      RECT 2040.665000  0.595000 2040.995000 0.885000 ;
      RECT 2040.665000  4.555000 2040.995000 4.845000 ;
      RECT 2040.765000  0.885000 2040.995000 1.065000 ;
      RECT 2040.765000  1.065000 2042.035000 1.365000 ;
      RECT 2040.765000  1.365000 2041.095000 4.075000 ;
      RECT 2040.765000  4.075000 2042.035000 4.375000 ;
      RECT 2040.765000  4.375000 2040.995000 4.555000 ;
      RECT 2041.165000  0.425000 2041.335000 0.770000 ;
      RECT 2041.165000  4.670000 2041.335000 5.015000 ;
      RECT 2041.265000  1.535000 2041.535000 2.465000 ;
      RECT 2041.265000  2.975000 2041.535000 3.905000 ;
      RECT 2041.505000  0.595000 2041.835000 1.065000 ;
      RECT 2041.505000  4.375000 2041.835000 4.845000 ;
      RECT 2041.705000  1.365000 2042.035000 4.075000 ;
      RECT 2042.005000  0.425000 2042.255000 0.770000 ;
      RECT 2042.005000  4.670000 2042.255000 5.015000 ;
      RECT 2042.205000  1.065000 2043.390000 1.395000 ;
      RECT 2042.205000  1.565000 2042.505000 2.465000 ;
      RECT 2042.205000  2.635000 2046.275000 2.805000 ;
      RECT 2042.205000  2.975000 2042.505000 3.875000 ;
      RECT 2042.205000  4.045000 2043.390000 4.375000 ;
      RECT 2042.750000  1.605000 2043.025000 2.635000 ;
      RECT 2042.750000  2.805000 2043.025000 3.835000 ;
      RECT 2042.760000  0.085000 2043.050000 0.610000 ;
      RECT 2042.760000  4.830000 2043.050000 5.355000 ;
      RECT 2043.220000  0.280000 2043.470000 0.825000 ;
      RECT 2043.220000  0.825000 2043.390000 1.065000 ;
      RECT 2043.220000  1.395000 2043.390000 1.605000 ;
      RECT 2043.220000  1.605000 2043.550000 2.465000 ;
      RECT 2043.220000  2.975000 2043.550000 3.835000 ;
      RECT 2043.220000  3.835000 2043.390000 4.045000 ;
      RECT 2043.220000  4.375000 2043.390000 4.615000 ;
      RECT 2043.220000  4.615000 2043.470000 5.160000 ;
      RECT 2043.560000  0.995000 2044.155000 1.325000 ;
      RECT 2043.560000  4.115000 2044.155000 4.445000 ;
      RECT 2043.680000  0.085000 2043.970000 0.610000 ;
      RECT 2043.680000  4.830000 2043.970000 5.355000 ;
      RECT 2043.720000  1.605000 2044.020000 2.635000 ;
      RECT 2043.720000  2.805000 2044.020000 3.835000 ;
      RECT 2044.325000  0.995000 2044.920000 1.325000 ;
      RECT 2044.325000  4.115000 2044.920000 4.445000 ;
      RECT 2044.460000  1.605000 2044.760000 2.635000 ;
      RECT 2044.460000  2.805000 2044.760000 3.835000 ;
      RECT 2044.510000  0.085000 2044.800000 0.610000 ;
      RECT 2044.510000  4.830000 2044.800000 5.355000 ;
      RECT 2044.930000  1.605000 2045.260000 2.465000 ;
      RECT 2044.930000  2.975000 2045.260000 3.835000 ;
      RECT 2045.010000  0.280000 2045.260000 0.825000 ;
      RECT 2045.010000  4.615000 2045.260000 5.160000 ;
      RECT 2045.090000  0.825000 2045.260000 1.065000 ;
      RECT 2045.090000  1.065000 2046.275000 1.395000 ;
      RECT 2045.090000  1.395000 2045.260000 1.605000 ;
      RECT 2045.090000  3.835000 2045.260000 4.045000 ;
      RECT 2045.090000  4.045000 2046.275000 4.375000 ;
      RECT 2045.090000  4.375000 2045.260000 4.615000 ;
      RECT 2045.430000  0.085000 2045.720000 0.610000 ;
      RECT 2045.430000  4.830000 2045.720000 5.355000 ;
      RECT 2045.455000  1.605000 2045.730000 2.635000 ;
      RECT 2045.455000  2.805000 2045.730000 3.835000 ;
      RECT 2045.975000  1.565000 2046.275000 2.465000 ;
      RECT 2045.975000  2.975000 2046.275000 3.875000 ;
      RECT 2046.225000  0.255000 2048.255000 0.425000 ;
      RECT 2046.225000  0.425000 2046.475000 0.770000 ;
      RECT 2046.225000  4.670000 2046.475000 5.015000 ;
      RECT 2046.225000  5.015000 2048.255000 5.185000 ;
      RECT 2046.445000  1.065000 2047.715000 1.365000 ;
      RECT 2046.445000  1.365000 2046.775000 4.075000 ;
      RECT 2046.445000  4.075000 2047.715000 4.375000 ;
      RECT 2046.645000  0.595000 2046.975000 1.065000 ;
      RECT 2046.645000  4.375000 2046.975000 4.845000 ;
      RECT 2046.945000  1.535000 2047.215000 2.465000 ;
      RECT 2046.945000  2.975000 2047.215000 3.905000 ;
      RECT 2047.145000  0.425000 2047.315000 0.770000 ;
      RECT 2047.145000  4.670000 2047.315000 5.015000 ;
      RECT 2047.385000  1.365000 2047.715000 4.075000 ;
      RECT 2047.485000  0.595000 2047.815000 0.885000 ;
      RECT 2047.485000  0.885000 2047.715000 1.065000 ;
      RECT 2047.485000  4.375000 2047.715000 4.555000 ;
      RECT 2047.485000  4.555000 2047.815000 4.845000 ;
      RECT 2047.885000  1.495000 2050.115000 1.665000 ;
      RECT 2047.885000  1.665000 2048.185000 2.465000 ;
      RECT 2047.885000  2.635000 2053.475000 2.805000 ;
      RECT 2047.885000  2.975000 2048.185000 3.775000 ;
      RECT 2047.885000  3.775000 2050.115000 3.945000 ;
      RECT 2047.985000  0.425000 2048.255000 0.715000 ;
      RECT 2047.985000  0.715000 2050.115000 0.885000 ;
      RECT 2047.985000  4.555000 2050.115000 4.725000 ;
      RECT 2047.985000  4.725000 2048.255000 5.015000 ;
      RECT 2048.405000  1.835000 2048.675000 2.635000 ;
      RECT 2048.405000  2.805000 2048.675000 3.605000 ;
      RECT 2048.425000  0.085000 2048.675000 0.545000 ;
      RECT 2048.425000  4.895000 2048.675000 5.355000 ;
      RECT 2048.845000  0.255000 2049.175000 0.715000 ;
      RECT 2048.845000  1.665000 2049.175000 2.465000 ;
      RECT 2048.845000  2.975000 2049.175000 3.775000 ;
      RECT 2048.845000  4.725000 2049.175000 5.185000 ;
      RECT 2048.895000  1.055000 2050.285000 1.325000 ;
      RECT 2048.895000  4.115000 2050.285000 4.385000 ;
      RECT 2049.345000  0.085000 2049.615000 0.545000 ;
      RECT 2049.345000  1.835000 2049.615000 2.635000 ;
      RECT 2049.345000  2.805000 2049.615000 3.605000 ;
      RECT 2049.345000  4.895000 2049.615000 5.355000 ;
      RECT 2049.785000  0.255000 2050.115000 0.715000 ;
      RECT 2049.785000  1.665000 2050.115000 2.465000 ;
      RECT 2049.785000  2.975000 2050.115000 3.775000 ;
      RECT 2049.785000  4.725000 2050.115000 5.185000 ;
      RECT 2050.285000  0.085000 2050.535000 0.885000 ;
      RECT 2050.285000  1.495000 2050.555000 2.635000 ;
      RECT 2050.285000  2.805000 2050.555000 3.945000 ;
      RECT 2050.285000  4.555000 2050.535000 5.355000 ;
      RECT 2050.805000  1.495000 2051.075000 2.635000 ;
      RECT 2050.805000  2.805000 2051.075000 3.945000 ;
      RECT 2050.825000  0.085000 2051.075000 0.885000 ;
      RECT 2050.825000  4.555000 2051.075000 5.355000 ;
      RECT 2051.075000  1.055000 2052.465000 1.325000 ;
      RECT 2051.075000  4.115000 2052.465000 4.385000 ;
      RECT 2051.245000  0.255000 2051.575000 0.715000 ;
      RECT 2051.245000  0.715000 2053.375000 0.885000 ;
      RECT 2051.245000  1.495000 2053.475000 1.665000 ;
      RECT 2051.245000  1.665000 2051.575000 2.465000 ;
      RECT 2051.245000  2.975000 2051.575000 3.775000 ;
      RECT 2051.245000  3.775000 2053.475000 3.945000 ;
      RECT 2051.245000  4.555000 2053.375000 4.725000 ;
      RECT 2051.245000  4.725000 2051.575000 5.185000 ;
      RECT 2051.745000  0.085000 2052.015000 0.545000 ;
      RECT 2051.745000  1.835000 2052.015000 2.635000 ;
      RECT 2051.745000  2.805000 2052.015000 3.605000 ;
      RECT 2051.745000  4.895000 2052.015000 5.355000 ;
      RECT 2052.185000  0.255000 2052.515000 0.715000 ;
      RECT 2052.185000  1.665000 2052.515000 2.465000 ;
      RECT 2052.185000  2.975000 2052.515000 3.775000 ;
      RECT 2052.185000  4.725000 2052.515000 5.185000 ;
      RECT 2052.685000  0.085000 2052.935000 0.545000 ;
      RECT 2052.685000  1.835000 2052.955000 2.635000 ;
      RECT 2052.685000  2.805000 2052.955000 3.605000 ;
      RECT 2052.685000  4.895000 2052.935000 5.355000 ;
      RECT 2053.105000  0.255000 2055.135000 0.425000 ;
      RECT 2053.105000  0.425000 2053.375000 0.715000 ;
      RECT 2053.105000  4.725000 2053.375000 5.015000 ;
      RECT 2053.105000  5.015000 2055.135000 5.185000 ;
      RECT 2053.175000  1.665000 2053.475000 2.465000 ;
      RECT 2053.175000  2.975000 2053.475000 3.775000 ;
      RECT 2053.545000  0.595000 2053.875000 0.885000 ;
      RECT 2053.545000  4.555000 2053.875000 4.845000 ;
      RECT 2053.645000  0.885000 2053.875000 1.065000 ;
      RECT 2053.645000  1.065000 2054.915000 1.365000 ;
      RECT 2053.645000  1.365000 2053.975000 4.075000 ;
      RECT 2053.645000  4.075000 2054.915000 4.375000 ;
      RECT 2053.645000  4.375000 2053.875000 4.555000 ;
      RECT 2054.045000  0.425000 2054.215000 0.770000 ;
      RECT 2054.045000  4.670000 2054.215000 5.015000 ;
      RECT 2054.145000  1.535000 2054.415000 2.465000 ;
      RECT 2054.145000  2.975000 2054.415000 3.905000 ;
      RECT 2054.385000  0.595000 2054.715000 1.065000 ;
      RECT 2054.385000  4.375000 2054.715000 4.845000 ;
      RECT 2054.585000  1.365000 2054.915000 4.075000 ;
      RECT 2054.885000  0.425000 2055.135000 0.770000 ;
      RECT 2054.885000  4.670000 2055.135000 5.015000 ;
      RECT 2055.085000  1.065000 2056.270000 1.395000 ;
      RECT 2055.085000  1.565000 2055.385000 2.465000 ;
      RECT 2055.085000  2.635000 2059.155000 2.805000 ;
      RECT 2055.085000  2.975000 2055.385000 3.875000 ;
      RECT 2055.085000  4.045000 2056.270000 4.375000 ;
      RECT 2055.630000  1.605000 2055.905000 2.635000 ;
      RECT 2055.630000  2.805000 2055.905000 3.835000 ;
      RECT 2055.640000  0.085000 2055.930000 0.610000 ;
      RECT 2055.640000  4.830000 2055.930000 5.355000 ;
      RECT 2056.100000  0.280000 2056.350000 0.825000 ;
      RECT 2056.100000  0.825000 2056.270000 1.065000 ;
      RECT 2056.100000  1.395000 2056.270000 1.605000 ;
      RECT 2056.100000  1.605000 2056.430000 2.465000 ;
      RECT 2056.100000  2.975000 2056.430000 3.835000 ;
      RECT 2056.100000  3.835000 2056.270000 4.045000 ;
      RECT 2056.100000  4.375000 2056.270000 4.615000 ;
      RECT 2056.100000  4.615000 2056.350000 5.160000 ;
      RECT 2056.440000  0.995000 2057.035000 1.325000 ;
      RECT 2056.440000  4.115000 2057.035000 4.445000 ;
      RECT 2056.560000  0.085000 2056.850000 0.610000 ;
      RECT 2056.560000  4.830000 2056.850000 5.355000 ;
      RECT 2056.600000  1.605000 2056.900000 2.635000 ;
      RECT 2056.600000  2.805000 2056.900000 3.835000 ;
      RECT 2057.205000  0.995000 2057.800000 1.325000 ;
      RECT 2057.205000  4.115000 2057.800000 4.445000 ;
      RECT 2057.340000  1.605000 2057.640000 2.635000 ;
      RECT 2057.340000  2.805000 2057.640000 3.835000 ;
      RECT 2057.390000  0.085000 2057.680000 0.610000 ;
      RECT 2057.390000  4.830000 2057.680000 5.355000 ;
      RECT 2057.810000  1.605000 2058.140000 2.465000 ;
      RECT 2057.810000  2.975000 2058.140000 3.835000 ;
      RECT 2057.890000  0.280000 2058.140000 0.825000 ;
      RECT 2057.890000  4.615000 2058.140000 5.160000 ;
      RECT 2057.970000  0.825000 2058.140000 1.065000 ;
      RECT 2057.970000  1.065000 2059.155000 1.395000 ;
      RECT 2057.970000  1.395000 2058.140000 1.605000 ;
      RECT 2057.970000  3.835000 2058.140000 4.045000 ;
      RECT 2057.970000  4.045000 2059.155000 4.375000 ;
      RECT 2057.970000  4.375000 2058.140000 4.615000 ;
      RECT 2058.310000  0.085000 2058.600000 0.610000 ;
      RECT 2058.310000  4.830000 2058.600000 5.355000 ;
      RECT 2058.335000  1.605000 2058.610000 2.635000 ;
      RECT 2058.335000  2.805000 2058.610000 3.835000 ;
      RECT 2058.855000  1.565000 2059.155000 2.465000 ;
      RECT 2058.855000  2.975000 2059.155000 3.875000 ;
      RECT 2059.105000  0.255000 2061.135000 0.425000 ;
      RECT 2059.105000  0.425000 2059.355000 0.770000 ;
      RECT 2059.105000  4.670000 2059.355000 5.015000 ;
      RECT 2059.105000  5.015000 2061.135000 5.185000 ;
      RECT 2059.325000  1.065000 2060.595000 1.365000 ;
      RECT 2059.325000  1.365000 2059.655000 4.075000 ;
      RECT 2059.325000  4.075000 2060.595000 4.375000 ;
      RECT 2059.525000  0.595000 2059.855000 1.065000 ;
      RECT 2059.525000  4.375000 2059.855000 4.845000 ;
      RECT 2059.825000  1.535000 2060.095000 2.465000 ;
      RECT 2059.825000  2.975000 2060.095000 3.905000 ;
      RECT 2060.025000  0.425000 2060.195000 0.770000 ;
      RECT 2060.025000  4.670000 2060.195000 5.015000 ;
      RECT 2060.265000  1.365000 2060.595000 4.075000 ;
      RECT 2060.365000  0.595000 2060.695000 0.885000 ;
      RECT 2060.365000  0.885000 2060.595000 1.065000 ;
      RECT 2060.365000  4.375000 2060.595000 4.555000 ;
      RECT 2060.365000  4.555000 2060.695000 4.845000 ;
      RECT 2060.765000  1.495000 2062.995000 1.665000 ;
      RECT 2060.765000  1.665000 2061.065000 2.465000 ;
      RECT 2060.765000  2.635000 2064.020000 2.805000 ;
      RECT 2060.765000  2.975000 2061.065000 3.775000 ;
      RECT 2060.765000  3.775000 2062.995000 3.945000 ;
      RECT 2060.865000  0.425000 2061.135000 0.715000 ;
      RECT 2060.865000  0.715000 2062.995000 0.885000 ;
      RECT 2060.865000  4.555000 2062.995000 4.725000 ;
      RECT 2060.865000  4.725000 2061.135000 5.015000 ;
      RECT 2061.285000  1.835000 2061.555000 2.635000 ;
      RECT 2061.285000  2.805000 2061.555000 3.605000 ;
      RECT 2061.305000  0.085000 2061.555000 0.545000 ;
      RECT 2061.305000  4.895000 2061.555000 5.355000 ;
      RECT 2061.725000  0.255000 2062.055000 0.715000 ;
      RECT 2061.725000  1.665000 2062.055000 2.465000 ;
      RECT 2061.725000  2.975000 2062.055000 3.775000 ;
      RECT 2061.725000  4.725000 2062.055000 5.185000 ;
      RECT 2061.775000  1.055000 2063.165000 1.325000 ;
      RECT 2061.775000  4.115000 2063.165000 4.385000 ;
      RECT 2062.225000  0.085000 2062.495000 0.545000 ;
      RECT 2062.225000  1.835000 2062.495000 2.635000 ;
      RECT 2062.225000  2.805000 2062.495000 3.605000 ;
      RECT 2062.225000  4.895000 2062.495000 5.355000 ;
      RECT 2062.665000  0.255000 2062.995000 0.715000 ;
      RECT 2062.665000  1.665000 2062.995000 2.465000 ;
      RECT 2062.665000  2.975000 2062.995000 3.775000 ;
      RECT 2062.665000  4.725000 2062.995000 5.185000 ;
      RECT 2063.165000  0.085000 2063.415000 0.885000 ;
      RECT 2063.165000  1.495000 2063.435000 2.635000 ;
      RECT 2063.165000  2.805000 2063.435000 3.945000 ;
      RECT 2063.165000  4.555000 2063.415000 5.355000 ;
      RECT 2063.645000  0.085000 2063.935000 0.810000 ;
      RECT 2063.645000  1.470000 2063.935000 2.635000 ;
      RECT 2063.645000  2.805000 2063.935000 3.970000 ;
      RECT 2063.645000  4.630000 2063.935000 5.355000 ;
    LAYER mcon ;
      RECT    0.145000 -0.085000    0.315000 0.085000 ;
      RECT    0.145000  2.635000    0.315000 2.805000 ;
      RECT    0.145000  5.355000    0.315000 5.525000 ;
      RECT    0.605000 -0.085000    0.775000 0.085000 ;
      RECT    0.605000  2.635000    0.775000 2.805000 ;
      RECT    0.605000  5.355000    0.775000 5.525000 ;
      RECT    1.065000 -0.085000    1.235000 0.085000 ;
      RECT    1.065000  2.635000    1.235000 2.805000 ;
      RECT    1.065000  5.355000    1.235000 5.525000 ;
      RECT    1.525000 -0.085000    1.695000 0.085000 ;
      RECT    1.525000  2.635000    1.695000 2.805000 ;
      RECT    1.525000  5.355000    1.695000 5.525000 ;
      RECT    1.985000 -0.085000    2.155000 0.085000 ;
      RECT    1.985000  2.635000    2.155000 2.805000 ;
      RECT    1.985000  5.355000    2.155000 5.525000 ;
      RECT    2.445000 -0.085000    2.615000 0.085000 ;
      RECT    2.445000  2.635000    2.615000 2.805000 ;
      RECT    2.445000  5.355000    2.615000 5.525000 ;
      RECT    2.905000 -0.085000    3.075000 0.085000 ;
      RECT    2.905000  2.635000    3.075000 2.805000 ;
      RECT    2.905000  5.355000    3.075000 5.525000 ;
      RECT    3.365000 -0.085000    3.535000 0.085000 ;
      RECT    3.365000  2.635000    3.535000 2.805000 ;
      RECT    3.365000  5.355000    3.535000 5.525000 ;
      RECT    3.825000 -0.085000    3.995000 0.085000 ;
      RECT    3.825000  2.635000    3.995000 2.805000 ;
      RECT    3.825000  5.355000    3.995000 5.525000 ;
      RECT    4.285000 -0.085000    4.455000 0.085000 ;
      RECT    4.285000  2.635000    4.455000 2.805000 ;
      RECT    4.285000  5.355000    4.455000 5.525000 ;
      RECT    4.745000 -0.085000    4.915000 0.085000 ;
      RECT    4.745000  2.635000    4.915000 2.805000 ;
      RECT    4.745000  5.355000    4.915000 5.525000 ;
      RECT    5.205000 -0.085000    5.375000 0.085000 ;
      RECT    5.205000  2.635000    5.375000 2.805000 ;
      RECT    5.205000  5.355000    5.375000 5.525000 ;
      RECT    5.665000 -0.085000    5.835000 0.085000 ;
      RECT    5.665000  2.635000    5.835000 2.805000 ;
      RECT    5.665000  5.355000    5.835000 5.525000 ;
      RECT    6.125000 -0.085000    6.295000 0.085000 ;
      RECT    6.125000  2.635000    6.295000 2.805000 ;
      RECT    6.125000  5.355000    6.295000 5.525000 ;
      RECT    6.585000 -0.085000    6.755000 0.085000 ;
      RECT    6.585000  2.635000    6.755000 2.805000 ;
      RECT    6.585000  5.355000    6.755000 5.525000 ;
      RECT    7.045000 -0.085000    7.215000 0.085000 ;
      RECT    7.045000  2.635000    7.215000 2.805000 ;
      RECT    7.045000  5.355000    7.215000 5.525000 ;
      RECT    7.505000 -0.085000    7.675000 0.085000 ;
      RECT    7.505000  2.635000    7.675000 2.805000 ;
      RECT    7.505000  5.355000    7.675000 5.525000 ;
      RECT    7.965000 -0.085000    8.135000 0.085000 ;
      RECT    7.965000  2.635000    8.135000 2.805000 ;
      RECT    7.965000  5.355000    8.135000 5.525000 ;
      RECT    8.425000 -0.085000    8.595000 0.085000 ;
      RECT    8.425000  2.635000    8.595000 2.805000 ;
      RECT    8.425000  5.355000    8.595000 5.525000 ;
      RECT    8.885000 -0.085000    9.055000 0.085000 ;
      RECT    8.885000  2.635000    9.055000 2.805000 ;
      RECT    8.885000  5.355000    9.055000 5.525000 ;
      RECT    9.345000 -0.085000    9.515000 0.085000 ;
      RECT    9.345000  2.635000    9.515000 2.805000 ;
      RECT    9.345000  5.355000    9.515000 5.525000 ;
      RECT    9.805000 -0.085000    9.975000 0.085000 ;
      RECT    9.805000  2.635000    9.975000 2.805000 ;
      RECT    9.805000  5.355000    9.975000 5.525000 ;
      RECT   10.265000 -0.085000   10.435000 0.085000 ;
      RECT   10.265000  2.635000   10.435000 2.805000 ;
      RECT   10.265000  5.355000   10.435000 5.525000 ;
      RECT   10.725000 -0.085000   10.895000 0.085000 ;
      RECT   10.725000  2.635000   10.895000 2.805000 ;
      RECT   10.725000  5.355000   10.895000 5.525000 ;
      RECT   11.185000 -0.085000   11.355000 0.085000 ;
      RECT   11.185000  2.635000   11.355000 2.805000 ;
      RECT   11.185000  5.355000   11.355000 5.525000 ;
      RECT   11.645000 -0.085000   11.815000 0.085000 ;
      RECT   11.645000  2.635000   11.815000 2.805000 ;
      RECT   11.645000  5.355000   11.815000 5.525000 ;
      RECT   12.105000 -0.085000   12.275000 0.085000 ;
      RECT   12.105000  2.635000   12.275000 2.805000 ;
      RECT   12.105000  5.355000   12.275000 5.525000 ;
      RECT   12.565000 -0.085000   12.735000 0.085000 ;
      RECT   12.565000  2.635000   12.735000 2.805000 ;
      RECT   12.565000  5.355000   12.735000 5.525000 ;
      RECT   13.025000 -0.085000   13.195000 0.085000 ;
      RECT   13.025000  2.635000   13.195000 2.805000 ;
      RECT   13.025000  5.355000   13.195000 5.525000 ;
      RECT   13.485000 -0.085000   13.655000 0.085000 ;
      RECT   13.485000  2.635000   13.655000 2.805000 ;
      RECT   13.485000  5.355000   13.655000 5.525000 ;
      RECT   13.945000 -0.085000   14.115000 0.085000 ;
      RECT   13.945000  2.635000   14.115000 2.805000 ;
      RECT   13.945000  5.355000   14.115000 5.525000 ;
      RECT   14.405000 -0.085000   14.575000 0.085000 ;
      RECT   14.405000  2.635000   14.575000 2.805000 ;
      RECT   14.405000  5.355000   14.575000 5.525000 ;
      RECT   14.865000 -0.085000   15.035000 0.085000 ;
      RECT   14.865000  2.635000   15.035000 2.805000 ;
      RECT   14.865000  5.355000   15.035000 5.525000 ;
      RECT   15.325000 -0.085000   15.495000 0.085000 ;
      RECT   15.325000  2.635000   15.495000 2.805000 ;
      RECT   15.325000  5.355000   15.495000 5.525000 ;
      RECT   15.785000 -0.085000   15.955000 0.085000 ;
      RECT   15.785000  2.635000   15.955000 2.805000 ;
      RECT   15.785000  5.355000   15.955000 5.525000 ;
      RECT   16.245000 -0.085000   16.415000 0.085000 ;
      RECT   16.245000  2.635000   16.415000 2.805000 ;
      RECT   16.245000  5.355000   16.415000 5.525000 ;
      RECT   16.705000 -0.085000   16.875000 0.085000 ;
      RECT   16.705000  2.635000   16.875000 2.805000 ;
      RECT   16.705000  5.355000   16.875000 5.525000 ;
      RECT   17.165000 -0.085000   17.335000 0.085000 ;
      RECT   17.165000  2.635000   17.335000 2.805000 ;
      RECT   17.165000  5.355000   17.335000 5.525000 ;
      RECT   17.625000 -0.085000   17.795000 0.085000 ;
      RECT   17.625000  2.635000   17.795000 2.805000 ;
      RECT   17.625000  5.355000   17.795000 5.525000 ;
      RECT   18.085000 -0.085000   18.255000 0.085000 ;
      RECT   18.085000  2.635000   18.255000 2.805000 ;
      RECT   18.085000  5.355000   18.255000 5.525000 ;
      RECT   18.545000 -0.085000   18.715000 0.085000 ;
      RECT   18.545000  2.635000   18.715000 2.805000 ;
      RECT   18.545000  5.355000   18.715000 5.525000 ;
      RECT   19.005000 -0.085000   19.175000 0.085000 ;
      RECT   19.005000  2.635000   19.175000 2.805000 ;
      RECT   19.005000  5.355000   19.175000 5.525000 ;
      RECT   19.465000 -0.085000   19.635000 0.085000 ;
      RECT   19.465000  2.635000   19.635000 2.805000 ;
      RECT   19.465000  5.355000   19.635000 5.525000 ;
      RECT   19.925000 -0.085000   20.095000 0.085000 ;
      RECT   19.925000  2.635000   20.095000 2.805000 ;
      RECT   19.925000  5.355000   20.095000 5.525000 ;
      RECT   20.385000 -0.085000   20.555000 0.085000 ;
      RECT   20.385000  2.635000   20.555000 2.805000 ;
      RECT   20.385000  5.355000   20.555000 5.525000 ;
      RECT   20.845000 -0.085000   21.015000 0.085000 ;
      RECT   20.845000  2.635000   21.015000 2.805000 ;
      RECT   20.845000  5.355000   21.015000 5.525000 ;
      RECT   21.305000 -0.085000   21.475000 0.085000 ;
      RECT   21.305000  2.635000   21.475000 2.805000 ;
      RECT   21.305000  5.355000   21.475000 5.525000 ;
      RECT   21.765000 -0.085000   21.935000 0.085000 ;
      RECT   21.765000  2.635000   21.935000 2.805000 ;
      RECT   21.765000  5.355000   21.935000 5.525000 ;
      RECT   22.225000 -0.085000   22.395000 0.085000 ;
      RECT   22.225000  2.635000   22.395000 2.805000 ;
      RECT   22.225000  5.355000   22.395000 5.525000 ;
      RECT   22.685000 -0.085000   22.855000 0.085000 ;
      RECT   22.685000  2.635000   22.855000 2.805000 ;
      RECT   22.685000  5.355000   22.855000 5.525000 ;
      RECT   23.145000 -0.085000   23.315000 0.085000 ;
      RECT   23.145000  2.635000   23.315000 2.805000 ;
      RECT   23.145000  5.355000   23.315000 5.525000 ;
      RECT   23.605000 -0.085000   23.775000 0.085000 ;
      RECT   23.605000  2.635000   23.775000 2.805000 ;
      RECT   23.605000  5.355000   23.775000 5.525000 ;
      RECT   24.065000 -0.085000   24.235000 0.085000 ;
      RECT   24.065000  2.635000   24.235000 2.805000 ;
      RECT   24.065000  5.355000   24.235000 5.525000 ;
      RECT   24.525000 -0.085000   24.695000 0.085000 ;
      RECT   24.525000  2.635000   24.695000 2.805000 ;
      RECT   24.525000  5.355000   24.695000 5.525000 ;
      RECT   24.985000 -0.085000   25.155000 0.085000 ;
      RECT   24.985000  2.635000   25.155000 2.805000 ;
      RECT   24.985000  5.355000   25.155000 5.525000 ;
      RECT   25.445000 -0.085000   25.615000 0.085000 ;
      RECT   25.445000  2.635000   25.615000 2.805000 ;
      RECT   25.445000  5.355000   25.615000 5.525000 ;
      RECT   25.905000 -0.085000   26.075000 0.085000 ;
      RECT   25.905000  2.635000   26.075000 2.805000 ;
      RECT   25.905000  5.355000   26.075000 5.525000 ;
      RECT   26.365000 -0.085000   26.535000 0.085000 ;
      RECT   26.365000  2.635000   26.535000 2.805000 ;
      RECT   26.365000  5.355000   26.535000 5.525000 ;
      RECT   26.825000 -0.085000   26.995000 0.085000 ;
      RECT   26.825000  2.635000   26.995000 2.805000 ;
      RECT   26.825000  5.355000   26.995000 5.525000 ;
      RECT   27.285000 -0.085000   27.455000 0.085000 ;
      RECT   27.285000  2.635000   27.455000 2.805000 ;
      RECT   27.285000  5.355000   27.455000 5.525000 ;
      RECT   27.745000 -0.085000   27.915000 0.085000 ;
      RECT   27.745000  2.635000   27.915000 2.805000 ;
      RECT   27.745000  5.355000   27.915000 5.525000 ;
      RECT   28.205000 -0.085000   28.375000 0.085000 ;
      RECT   28.205000  2.635000   28.375000 2.805000 ;
      RECT   28.205000  5.355000   28.375000 5.525000 ;
      RECT   28.665000 -0.085000   28.835000 0.085000 ;
      RECT   28.665000  2.635000   28.835000 2.805000 ;
      RECT   28.665000  5.355000   28.835000 5.525000 ;
      RECT   29.125000 -0.085000   29.295000 0.085000 ;
      RECT   29.125000  2.635000   29.295000 2.805000 ;
      RECT   29.125000  5.355000   29.295000 5.525000 ;
      RECT   29.585000 -0.085000   29.755000 0.085000 ;
      RECT   29.585000  1.445000   29.755000 1.615000 ;
      RECT   29.585000  2.635000   29.755000 2.805000 ;
      RECT   29.585000  5.355000   29.755000 5.525000 ;
      RECT   30.045000 -0.085000   30.215000 0.085000 ;
      RECT   30.045000  2.635000   30.215000 2.805000 ;
      RECT   30.045000  5.355000   30.215000 5.525000 ;
      RECT   30.505000 -0.085000   30.675000 0.085000 ;
      RECT   30.505000  2.635000   30.675000 2.805000 ;
      RECT   30.505000  5.355000   30.675000 5.525000 ;
      RECT   30.965000 -0.085000   31.135000 0.085000 ;
      RECT   30.965000  2.635000   31.135000 2.805000 ;
      RECT   30.965000  5.355000   31.135000 5.525000 ;
      RECT   31.425000 -0.085000   31.595000 0.085000 ;
      RECT   31.425000  2.635000   31.595000 2.805000 ;
      RECT   31.425000  5.355000   31.595000 5.525000 ;
      RECT   31.885000 -0.085000   32.055000 0.085000 ;
      RECT   31.885000  2.635000   32.055000 2.805000 ;
      RECT   31.885000  5.355000   32.055000 5.525000 ;
      RECT   32.345000 -0.085000   32.515000 0.085000 ;
      RECT   32.345000  2.635000   32.515000 2.805000 ;
      RECT   32.345000  5.355000   32.515000 5.525000 ;
      RECT   32.640000  1.445000   32.810000 1.615000 ;
      RECT   32.805000 -0.085000   32.975000 0.085000 ;
      RECT   32.805000  2.635000   32.975000 2.805000 ;
      RECT   32.805000  5.355000   32.975000 5.525000 ;
      RECT   33.265000 -0.085000   33.435000 0.085000 ;
      RECT   33.265000  2.635000   33.435000 2.805000 ;
      RECT   33.265000  5.355000   33.435000 5.525000 ;
      RECT   33.725000 -0.085000   33.895000 0.085000 ;
      RECT   33.725000  2.635000   33.895000 2.805000 ;
      RECT   33.725000  5.355000   33.895000 5.525000 ;
      RECT   34.185000 -0.085000   34.355000 0.085000 ;
      RECT   34.185000  2.635000   34.355000 2.805000 ;
      RECT   34.185000  5.355000   34.355000 5.525000 ;
      RECT   34.645000 -0.085000   34.815000 0.085000 ;
      RECT   34.645000  2.635000   34.815000 2.805000 ;
      RECT   34.645000  5.355000   34.815000 5.525000 ;
      RECT   35.105000 -0.085000   35.275000 0.085000 ;
      RECT   35.105000  2.635000   35.275000 2.805000 ;
      RECT   35.105000  5.355000   35.275000 5.525000 ;
      RECT   35.565000 -0.085000   35.735000 0.085000 ;
      RECT   35.565000  2.635000   35.735000 2.805000 ;
      RECT   35.565000  5.355000   35.735000 5.525000 ;
      RECT   36.025000 -0.085000   36.195000 0.085000 ;
      RECT   36.025000  2.635000   36.195000 2.805000 ;
      RECT   36.025000  5.355000   36.195000 5.525000 ;
      RECT   36.485000 -0.085000   36.655000 0.085000 ;
      RECT   36.485000  2.635000   36.655000 2.805000 ;
      RECT   36.485000  5.355000   36.655000 5.525000 ;
      RECT   36.945000 -0.085000   37.115000 0.085000 ;
      RECT   36.945000  2.635000   37.115000 2.805000 ;
      RECT   36.945000  5.355000   37.115000 5.525000 ;
      RECT   37.405000 -0.085000   37.575000 0.085000 ;
      RECT   37.405000  2.635000   37.575000 2.805000 ;
      RECT   37.405000  5.355000   37.575000 5.525000 ;
      RECT   37.865000 -0.085000   38.035000 0.085000 ;
      RECT   37.865000  2.635000   38.035000 2.805000 ;
      RECT   37.865000  5.355000   38.035000 5.525000 ;
      RECT   38.325000 -0.085000   38.495000 0.085000 ;
      RECT   38.325000  2.635000   38.495000 2.805000 ;
      RECT   38.325000  5.355000   38.495000 5.525000 ;
      RECT   38.785000 -0.085000   38.955000 0.085000 ;
      RECT   38.785000  2.635000   38.955000 2.805000 ;
      RECT   38.785000  5.355000   38.955000 5.525000 ;
      RECT   39.245000 -0.085000   39.415000 0.085000 ;
      RECT   39.245000  2.635000   39.415000 2.805000 ;
      RECT   39.245000  5.355000   39.415000 5.525000 ;
      RECT   39.705000 -0.085000   39.875000 0.085000 ;
      RECT   39.705000  2.635000   39.875000 2.805000 ;
      RECT   39.705000  5.355000   39.875000 5.525000 ;
      RECT   40.165000 -0.085000   40.335000 0.085000 ;
      RECT   40.165000  2.635000   40.335000 2.805000 ;
      RECT   40.165000  5.355000   40.335000 5.525000 ;
      RECT   40.625000 -0.085000   40.795000 0.085000 ;
      RECT   40.625000  2.635000   40.795000 2.805000 ;
      RECT   40.625000  5.355000   40.795000 5.525000 ;
      RECT   41.085000 -0.085000   41.255000 0.085000 ;
      RECT   41.085000  2.635000   41.255000 2.805000 ;
      RECT   41.085000  5.355000   41.255000 5.525000 ;
      RECT   41.545000 -0.085000   41.715000 0.085000 ;
      RECT   41.545000  2.635000   41.715000 2.805000 ;
      RECT   41.545000  5.355000   41.715000 5.525000 ;
      RECT   42.005000 -0.085000   42.175000 0.085000 ;
      RECT   42.005000  2.635000   42.175000 2.805000 ;
      RECT   42.005000  5.355000   42.175000 5.525000 ;
      RECT   42.465000 -0.085000   42.635000 0.085000 ;
      RECT   42.465000  2.635000   42.635000 2.805000 ;
      RECT   42.465000  5.355000   42.635000 5.525000 ;
      RECT   42.925000 -0.085000   43.095000 0.085000 ;
      RECT   42.925000  2.635000   43.095000 2.805000 ;
      RECT   42.925000  5.355000   43.095000 5.525000 ;
      RECT   43.385000 -0.085000   43.555000 0.085000 ;
      RECT   43.385000  2.635000   43.555000 2.805000 ;
      RECT   43.385000  5.355000   43.555000 5.525000 ;
      RECT   43.845000 -0.085000   44.015000 0.085000 ;
      RECT   43.845000  2.635000   44.015000 2.805000 ;
      RECT   43.845000  5.355000   44.015000 5.525000 ;
      RECT   44.305000 -0.085000   44.475000 0.085000 ;
      RECT   44.305000  2.635000   44.475000 2.805000 ;
      RECT   44.305000  5.355000   44.475000 5.525000 ;
      RECT   44.765000 -0.085000   44.935000 0.085000 ;
      RECT   44.765000  2.635000   44.935000 2.805000 ;
      RECT   44.765000  5.355000   44.935000 5.525000 ;
      RECT   45.225000 -0.085000   45.395000 0.085000 ;
      RECT   45.225000  2.635000   45.395000 2.805000 ;
      RECT   45.225000  5.355000   45.395000 5.525000 ;
      RECT   45.685000 -0.085000   45.855000 0.085000 ;
      RECT   45.685000  2.635000   45.855000 2.805000 ;
      RECT   45.685000  5.355000   45.855000 5.525000 ;
      RECT   46.145000 -0.085000   46.315000 0.085000 ;
      RECT   46.145000  2.635000   46.315000 2.805000 ;
      RECT   46.145000  5.355000   46.315000 5.525000 ;
      RECT   46.605000 -0.085000   46.775000 0.085000 ;
      RECT   46.605000  2.635000   46.775000 2.805000 ;
      RECT   46.605000  5.355000   46.775000 5.525000 ;
      RECT   47.065000 -0.085000   47.235000 0.085000 ;
      RECT   47.065000  2.635000   47.235000 2.805000 ;
      RECT   47.065000  5.355000   47.235000 5.525000 ;
      RECT   47.525000 -0.085000   47.695000 0.085000 ;
      RECT   47.525000  2.635000   47.695000 2.805000 ;
      RECT   47.525000  5.355000   47.695000 5.525000 ;
      RECT   47.985000 -0.085000   48.155000 0.085000 ;
      RECT   47.985000  2.635000   48.155000 2.805000 ;
      RECT   47.985000  5.355000   48.155000 5.525000 ;
      RECT   48.445000 -0.085000   48.615000 0.085000 ;
      RECT   48.445000  2.635000   48.615000 2.805000 ;
      RECT   48.445000  5.355000   48.615000 5.525000 ;
      RECT   48.905000 -0.085000   49.075000 0.085000 ;
      RECT   48.905000  2.635000   49.075000 2.805000 ;
      RECT   48.905000  5.355000   49.075000 5.525000 ;
      RECT   49.365000 -0.085000   49.535000 0.085000 ;
      RECT   49.365000  2.635000   49.535000 2.805000 ;
      RECT   49.365000  5.355000   49.535000 5.525000 ;
      RECT   49.825000 -0.085000   49.995000 0.085000 ;
      RECT   49.825000  2.635000   49.995000 2.805000 ;
      RECT   49.825000  5.355000   49.995000 5.525000 ;
      RECT   50.285000 -0.085000   50.455000 0.085000 ;
      RECT   50.285000  2.635000   50.455000 2.805000 ;
      RECT   50.285000  5.355000   50.455000 5.525000 ;
      RECT   50.745000 -0.085000   50.915000 0.085000 ;
      RECT   50.745000  2.635000   50.915000 2.805000 ;
      RECT   50.745000  5.355000   50.915000 5.525000 ;
      RECT   51.205000 -0.085000   51.375000 0.085000 ;
      RECT   51.205000  2.635000   51.375000 2.805000 ;
      RECT   51.205000  5.355000   51.375000 5.525000 ;
      RECT   51.665000 -0.085000   51.835000 0.085000 ;
      RECT   51.665000  2.635000   51.835000 2.805000 ;
      RECT   51.665000  5.355000   51.835000 5.525000 ;
      RECT   52.125000 -0.085000   52.295000 0.085000 ;
      RECT   52.125000  2.635000   52.295000 2.805000 ;
      RECT   52.125000  5.355000   52.295000 5.525000 ;
      RECT   52.155000  4.845000   52.325000 5.015000 ;
      RECT   52.585000 -0.085000   52.755000 0.085000 ;
      RECT   52.585000  2.635000   52.755000 2.805000 ;
      RECT   52.585000  5.355000   52.755000 5.525000 ;
      RECT   52.625000  3.485000   52.795000 3.655000 ;
      RECT   53.045000 -0.085000   53.215000 0.085000 ;
      RECT   53.045000  2.635000   53.215000 2.805000 ;
      RECT   53.045000  5.355000   53.215000 5.525000 ;
      RECT   53.505000 -0.085000   53.675000 0.085000 ;
      RECT   53.505000  2.635000   53.675000 2.805000 ;
      RECT   53.505000  5.355000   53.675000 5.525000 ;
      RECT   53.565000  3.485000   53.735000 3.655000 ;
      RECT   53.965000 -0.085000   54.135000 0.085000 ;
      RECT   53.965000  2.635000   54.135000 2.805000 ;
      RECT   53.965000  5.355000   54.135000 5.525000 ;
      RECT   54.425000 -0.085000   54.595000 0.085000 ;
      RECT   54.425000  2.635000   54.595000 2.805000 ;
      RECT   54.425000  5.355000   54.595000 5.525000 ;
      RECT   54.885000 -0.085000   55.055000 0.085000 ;
      RECT   54.885000  2.635000   55.055000 2.805000 ;
      RECT   54.885000  5.355000   55.055000 5.525000 ;
      RECT   55.025000  3.145000   55.195000 3.315000 ;
      RECT   55.345000 -0.085000   55.515000 0.085000 ;
      RECT   55.345000  2.635000   55.515000 2.805000 ;
      RECT   55.345000  5.355000   55.515000 5.525000 ;
      RECT   55.805000 -0.085000   55.975000 0.085000 ;
      RECT   55.805000  2.635000   55.975000 2.805000 ;
      RECT   55.805000  5.355000   55.975000 5.525000 ;
      RECT   55.965000  3.145000   56.135000 3.315000 ;
      RECT   56.265000 -0.085000   56.435000 0.085000 ;
      RECT   56.265000  2.635000   56.435000 2.805000 ;
      RECT   56.265000  5.355000   56.435000 5.525000 ;
      RECT   56.725000 -0.085000   56.895000 0.085000 ;
      RECT   56.725000  2.635000   56.895000 2.805000 ;
      RECT   56.725000  5.355000   56.895000 5.525000 ;
      RECT   57.185000 -0.085000   57.355000 0.085000 ;
      RECT   57.185000  2.635000   57.355000 2.805000 ;
      RECT   57.185000  5.355000   57.355000 5.525000 ;
      RECT   57.645000 -0.085000   57.815000 0.085000 ;
      RECT   57.645000  2.635000   57.815000 2.805000 ;
      RECT   57.645000  5.355000   57.815000 5.525000 ;
      RECT   57.845000  3.485000   58.015000 3.655000 ;
      RECT   58.105000 -0.085000   58.275000 0.085000 ;
      RECT   58.105000  2.635000   58.275000 2.805000 ;
      RECT   58.105000  5.355000   58.275000 5.525000 ;
      RECT   58.565000 -0.085000   58.735000 0.085000 ;
      RECT   58.565000  2.635000   58.735000 2.805000 ;
      RECT   58.565000  5.355000   58.735000 5.525000 ;
      RECT   58.785000  3.485000   58.955000 3.655000 ;
      RECT   59.025000 -0.085000   59.195000 0.085000 ;
      RECT   59.025000  2.635000   59.195000 2.805000 ;
      RECT   59.025000  5.355000   59.195000 5.525000 ;
      RECT   59.485000 -0.085000   59.655000 0.085000 ;
      RECT   59.485000  2.635000   59.655000 2.805000 ;
      RECT   59.485000  5.355000   59.655000 5.525000 ;
      RECT   59.945000 -0.085000   60.115000 0.085000 ;
      RECT   59.945000  2.635000   60.115000 2.805000 ;
      RECT   59.945000  5.355000   60.115000 5.525000 ;
      RECT   60.245000  3.485000   60.415000 3.655000 ;
      RECT   60.405000 -0.085000   60.575000 0.085000 ;
      RECT   60.405000  2.635000   60.575000 2.805000 ;
      RECT   60.405000  5.355000   60.575000 5.525000 ;
      RECT   60.865000 -0.085000   61.035000 0.085000 ;
      RECT   60.865000  2.635000   61.035000 2.805000 ;
      RECT   60.865000  5.355000   61.035000 5.525000 ;
      RECT   61.185000  3.485000   61.355000 3.655000 ;
      RECT   61.325000 -0.085000   61.495000 0.085000 ;
      RECT   61.325000  2.635000   61.495000 2.805000 ;
      RECT   61.325000  5.355000   61.495000 5.525000 ;
      RECT   61.655000  4.845000   61.825000 5.015000 ;
      RECT   61.785000 -0.085000   61.955000 0.085000 ;
      RECT   61.785000  2.635000   61.955000 2.805000 ;
      RECT   61.785000  5.355000   61.955000 5.525000 ;
      RECT   62.245000 -0.085000   62.415000 0.085000 ;
      RECT   62.245000  2.635000   62.415000 2.805000 ;
      RECT   62.245000  5.355000   62.415000 5.525000 ;
      RECT   62.705000 -0.085000   62.875000 0.085000 ;
      RECT   62.705000  2.635000   62.875000 2.805000 ;
      RECT   62.705000  5.355000   62.875000 5.525000 ;
      RECT   63.165000 -0.085000   63.335000 0.085000 ;
      RECT   63.165000  2.635000   63.335000 2.805000 ;
      RECT   63.165000  5.355000   63.335000 5.525000 ;
      RECT   63.625000 -0.085000   63.795000 0.085000 ;
      RECT   63.625000  2.635000   63.795000 2.805000 ;
      RECT   63.625000  5.355000   63.795000 5.525000 ;
      RECT   64.085000 -0.085000   64.255000 0.085000 ;
      RECT   64.085000  2.635000   64.255000 2.805000 ;
      RECT   64.085000  5.355000   64.255000 5.525000 ;
      RECT   64.545000 -0.085000   64.715000 0.085000 ;
      RECT   64.545000  2.635000   64.715000 2.805000 ;
      RECT   64.545000  5.355000   64.715000 5.525000 ;
      RECT   65.005000 -0.085000   65.175000 0.085000 ;
      RECT   65.005000  2.635000   65.175000 2.805000 ;
      RECT   65.005000  5.355000   65.175000 5.525000 ;
      RECT   65.465000 -0.085000   65.635000 0.085000 ;
      RECT   65.465000  2.635000   65.635000 2.805000 ;
      RECT   65.465000  5.355000   65.635000 5.525000 ;
      RECT   65.925000 -0.085000   66.095000 0.085000 ;
      RECT   65.925000  2.635000   66.095000 2.805000 ;
      RECT   65.925000  5.355000   66.095000 5.525000 ;
      RECT   66.385000 -0.085000   66.555000 0.085000 ;
      RECT   66.385000  2.635000   66.555000 2.805000 ;
      RECT   66.385000  5.355000   66.555000 5.525000 ;
      RECT   66.845000 -0.085000   67.015000 0.085000 ;
      RECT   66.845000  2.635000   67.015000 2.805000 ;
      RECT   66.845000  5.355000   67.015000 5.525000 ;
      RECT   67.305000 -0.085000   67.475000 0.085000 ;
      RECT   67.305000  2.635000   67.475000 2.805000 ;
      RECT   67.305000  5.355000   67.475000 5.525000 ;
      RECT   67.765000 -0.085000   67.935000 0.085000 ;
      RECT   67.765000  2.635000   67.935000 2.805000 ;
      RECT   67.765000  5.355000   67.935000 5.525000 ;
      RECT   68.225000 -0.085000   68.395000 0.085000 ;
      RECT   68.225000  2.635000   68.395000 2.805000 ;
      RECT   68.225000  5.355000   68.395000 5.525000 ;
      RECT   68.685000 -0.085000   68.855000 0.085000 ;
      RECT   68.685000  2.635000   68.855000 2.805000 ;
      RECT   68.685000  5.355000   68.855000 5.525000 ;
      RECT   69.145000 -0.085000   69.315000 0.085000 ;
      RECT   69.145000  2.635000   69.315000 2.805000 ;
      RECT   69.145000  5.355000   69.315000 5.525000 ;
      RECT   69.175000  4.845000   69.345000 5.015000 ;
      RECT   69.605000 -0.085000   69.775000 0.085000 ;
      RECT   69.605000  2.635000   69.775000 2.805000 ;
      RECT   69.605000  5.355000   69.775000 5.525000 ;
      RECT   69.645000  3.485000   69.815000 3.655000 ;
      RECT   70.065000 -0.085000   70.235000 0.085000 ;
      RECT   70.065000  2.635000   70.235000 2.805000 ;
      RECT   70.065000  5.355000   70.235000 5.525000 ;
      RECT   70.525000 -0.085000   70.695000 0.085000 ;
      RECT   70.525000  2.635000   70.695000 2.805000 ;
      RECT   70.525000  5.355000   70.695000 5.525000 ;
      RECT   70.585000  3.485000   70.755000 3.655000 ;
      RECT   70.985000 -0.085000   71.155000 0.085000 ;
      RECT   70.985000  2.635000   71.155000 2.805000 ;
      RECT   70.985000  5.355000   71.155000 5.525000 ;
      RECT   71.445000 -0.085000   71.615000 0.085000 ;
      RECT   71.445000  2.635000   71.615000 2.805000 ;
      RECT   71.445000  5.355000   71.615000 5.525000 ;
      RECT   71.905000 -0.085000   72.075000 0.085000 ;
      RECT   71.905000  2.635000   72.075000 2.805000 ;
      RECT   71.905000  5.355000   72.075000 5.525000 ;
      RECT   72.045000  3.145000   72.215000 3.315000 ;
      RECT   72.365000 -0.085000   72.535000 0.085000 ;
      RECT   72.365000  2.635000   72.535000 2.805000 ;
      RECT   72.365000  5.355000   72.535000 5.525000 ;
      RECT   72.825000 -0.085000   72.995000 0.085000 ;
      RECT   72.825000  2.635000   72.995000 2.805000 ;
      RECT   72.825000  5.355000   72.995000 5.525000 ;
      RECT   72.985000  3.145000   73.155000 3.315000 ;
      RECT   73.285000 -0.085000   73.455000 0.085000 ;
      RECT   73.285000  2.635000   73.455000 2.805000 ;
      RECT   73.285000  5.355000   73.455000 5.525000 ;
      RECT   73.745000 -0.085000   73.915000 0.085000 ;
      RECT   73.745000  2.635000   73.915000 2.805000 ;
      RECT   73.745000  5.355000   73.915000 5.525000 ;
      RECT   74.205000 -0.085000   74.375000 0.085000 ;
      RECT   74.205000  2.635000   74.375000 2.805000 ;
      RECT   74.205000  5.355000   74.375000 5.525000 ;
      RECT   74.665000 -0.085000   74.835000 0.085000 ;
      RECT   74.665000  2.635000   74.835000 2.805000 ;
      RECT   74.665000  5.355000   74.835000 5.525000 ;
      RECT   74.865000  3.485000   75.035000 3.655000 ;
      RECT   75.125000 -0.085000   75.295000 0.085000 ;
      RECT   75.125000  2.635000   75.295000 2.805000 ;
      RECT   75.125000  5.355000   75.295000 5.525000 ;
      RECT   75.585000 -0.085000   75.755000 0.085000 ;
      RECT   75.585000  2.635000   75.755000 2.805000 ;
      RECT   75.585000  5.355000   75.755000 5.525000 ;
      RECT   75.805000  3.485000   75.975000 3.655000 ;
      RECT   76.045000 -0.085000   76.215000 0.085000 ;
      RECT   76.045000  2.635000   76.215000 2.805000 ;
      RECT   76.045000  5.355000   76.215000 5.525000 ;
      RECT   76.505000 -0.085000   76.675000 0.085000 ;
      RECT   76.505000  2.635000   76.675000 2.805000 ;
      RECT   76.505000  5.355000   76.675000 5.525000 ;
      RECT   76.965000 -0.085000   77.135000 0.085000 ;
      RECT   76.965000  2.635000   77.135000 2.805000 ;
      RECT   76.965000  5.355000   77.135000 5.525000 ;
      RECT   77.265000  3.485000   77.435000 3.655000 ;
      RECT   77.425000 -0.085000   77.595000 0.085000 ;
      RECT   77.425000  2.635000   77.595000 2.805000 ;
      RECT   77.425000  5.355000   77.595000 5.525000 ;
      RECT   77.885000 -0.085000   78.055000 0.085000 ;
      RECT   77.885000  2.635000   78.055000 2.805000 ;
      RECT   77.885000  5.355000   78.055000 5.525000 ;
      RECT   78.205000  3.485000   78.375000 3.655000 ;
      RECT   78.345000 -0.085000   78.515000 0.085000 ;
      RECT   78.345000  2.635000   78.515000 2.805000 ;
      RECT   78.345000  5.355000   78.515000 5.525000 ;
      RECT   78.675000  4.845000   78.845000 5.015000 ;
      RECT   78.805000 -0.085000   78.975000 0.085000 ;
      RECT   78.805000  2.635000   78.975000 2.805000 ;
      RECT   78.805000  5.355000   78.975000 5.525000 ;
      RECT   79.265000 -0.085000   79.435000 0.085000 ;
      RECT   79.265000  2.635000   79.435000 2.805000 ;
      RECT   79.265000  5.355000   79.435000 5.525000 ;
      RECT   79.725000 -0.085000   79.895000 0.085000 ;
      RECT   79.725000  2.635000   79.895000 2.805000 ;
      RECT   79.725000  5.355000   79.895000 5.525000 ;
      RECT   80.185000 -0.085000   80.355000 0.085000 ;
      RECT   80.185000  2.635000   80.355000 2.805000 ;
      RECT   80.185000  5.355000   80.355000 5.525000 ;
      RECT   80.645000 -0.085000   80.815000 0.085000 ;
      RECT   80.645000  2.635000   80.815000 2.805000 ;
      RECT   80.645000  5.355000   80.815000 5.525000 ;
      RECT   81.105000 -0.085000   81.275000 0.085000 ;
      RECT   81.105000  2.635000   81.275000 2.805000 ;
      RECT   81.105000  5.355000   81.275000 5.525000 ;
      RECT   81.565000 -0.085000   81.735000 0.085000 ;
      RECT   81.565000  2.635000   81.735000 2.805000 ;
      RECT   81.565000  5.355000   81.735000 5.525000 ;
      RECT   82.025000 -0.085000   82.195000 0.085000 ;
      RECT   82.025000  2.635000   82.195000 2.805000 ;
      RECT   82.025000  5.355000   82.195000 5.525000 ;
      RECT   82.485000 -0.085000   82.655000 0.085000 ;
      RECT   82.485000  2.635000   82.655000 2.805000 ;
      RECT   82.485000  5.355000   82.655000 5.525000 ;
      RECT   82.945000 -0.085000   83.115000 0.085000 ;
      RECT   82.945000  2.635000   83.115000 2.805000 ;
      RECT   82.945000  5.355000   83.115000 5.525000 ;
      RECT   83.405000 -0.085000   83.575000 0.085000 ;
      RECT   83.405000  2.635000   83.575000 2.805000 ;
      RECT   83.405000  5.355000   83.575000 5.525000 ;
      RECT   83.865000 -0.085000   84.035000 0.085000 ;
      RECT   83.865000  2.635000   84.035000 2.805000 ;
      RECT   83.865000  5.355000   84.035000 5.525000 ;
      RECT   84.325000 -0.085000   84.495000 0.085000 ;
      RECT   84.325000  2.635000   84.495000 2.805000 ;
      RECT   84.325000  5.355000   84.495000 5.525000 ;
      RECT   84.785000 -0.085000   84.955000 0.085000 ;
      RECT   84.785000  2.635000   84.955000 2.805000 ;
      RECT   84.785000  5.355000   84.955000 5.525000 ;
      RECT   85.245000 -0.085000   85.415000 0.085000 ;
      RECT   85.245000  2.635000   85.415000 2.805000 ;
      RECT   85.245000  5.355000   85.415000 5.525000 ;
      RECT   85.705000 -0.085000   85.875000 0.085000 ;
      RECT   85.705000  2.635000   85.875000 2.805000 ;
      RECT   85.705000  5.355000   85.875000 5.525000 ;
      RECT   86.165000 -0.085000   86.335000 0.085000 ;
      RECT   86.165000  2.635000   86.335000 2.805000 ;
      RECT   86.165000  5.355000   86.335000 5.525000 ;
      RECT   86.625000 -0.085000   86.795000 0.085000 ;
      RECT   86.625000  2.635000   86.795000 2.805000 ;
      RECT   86.625000  5.355000   86.795000 5.525000 ;
      RECT   87.085000 -0.085000   87.255000 0.085000 ;
      RECT   87.085000  2.635000   87.255000 2.805000 ;
      RECT   87.085000  5.355000   87.255000 5.525000 ;
      RECT   87.545000 -0.085000   87.715000 0.085000 ;
      RECT   87.545000  2.635000   87.715000 2.805000 ;
      RECT   87.545000  5.355000   87.715000 5.525000 ;
      RECT   88.005000 -0.085000   88.175000 0.085000 ;
      RECT   88.005000  2.635000   88.175000 2.805000 ;
      RECT   88.005000  5.355000   88.175000 5.525000 ;
      RECT   88.465000 -0.085000   88.635000 0.085000 ;
      RECT   88.465000  2.635000   88.635000 2.805000 ;
      RECT   88.465000  5.355000   88.635000 5.525000 ;
      RECT   88.925000 -0.085000   89.095000 0.085000 ;
      RECT   88.925000  2.635000   89.095000 2.805000 ;
      RECT   88.925000  5.355000   89.095000 5.525000 ;
      RECT   89.385000 -0.085000   89.555000 0.085000 ;
      RECT   89.385000  2.635000   89.555000 2.805000 ;
      RECT   89.385000  5.355000   89.555000 5.525000 ;
      RECT   89.845000 -0.085000   90.015000 0.085000 ;
      RECT   89.845000  2.635000   90.015000 2.805000 ;
      RECT   89.845000  5.355000   90.015000 5.525000 ;
      RECT   90.305000 -0.085000   90.475000 0.085000 ;
      RECT   90.305000  2.635000   90.475000 2.805000 ;
      RECT   90.305000  5.355000   90.475000 5.525000 ;
      RECT   90.765000 -0.085000   90.935000 0.085000 ;
      RECT   90.765000  2.635000   90.935000 2.805000 ;
      RECT   90.765000  5.355000   90.935000 5.525000 ;
      RECT   91.225000 -0.085000   91.395000 0.085000 ;
      RECT   91.225000  2.635000   91.395000 2.805000 ;
      RECT   91.225000  5.355000   91.395000 5.525000 ;
      RECT   91.685000 -0.085000   91.855000 0.085000 ;
      RECT   91.685000  2.635000   91.855000 2.805000 ;
      RECT   91.685000  5.355000   91.855000 5.525000 ;
      RECT   92.145000 -0.085000   92.315000 0.085000 ;
      RECT   92.145000  2.635000   92.315000 2.805000 ;
      RECT   92.145000  5.355000   92.315000 5.525000 ;
      RECT   92.605000 -0.085000   92.775000 0.085000 ;
      RECT   92.605000  2.635000   92.775000 2.805000 ;
      RECT   92.605000  5.355000   92.775000 5.525000 ;
      RECT   93.065000 -0.085000   93.235000 0.085000 ;
      RECT   93.065000  2.635000   93.235000 2.805000 ;
      RECT   93.065000  5.355000   93.235000 5.525000 ;
      RECT   93.525000 -0.085000   93.695000 0.085000 ;
      RECT   93.525000  2.635000   93.695000 2.805000 ;
      RECT   93.525000  5.355000   93.695000 5.525000 ;
      RECT   93.985000 -0.085000   94.155000 0.085000 ;
      RECT   93.985000  2.635000   94.155000 2.805000 ;
      RECT   93.985000  5.355000   94.155000 5.525000 ;
      RECT   94.445000 -0.085000   94.615000 0.085000 ;
      RECT   94.445000  2.635000   94.615000 2.805000 ;
      RECT   94.445000  5.355000   94.615000 5.525000 ;
      RECT   94.905000 -0.085000   95.075000 0.085000 ;
      RECT   94.905000  2.635000   95.075000 2.805000 ;
      RECT   94.905000  5.355000   95.075000 5.525000 ;
      RECT   95.365000 -0.085000   95.535000 0.085000 ;
      RECT   95.365000  2.635000   95.535000 2.805000 ;
      RECT   95.365000  5.355000   95.535000 5.525000 ;
      RECT   95.825000 -0.085000   95.995000 0.085000 ;
      RECT   95.825000  2.635000   95.995000 2.805000 ;
      RECT   95.825000  5.355000   95.995000 5.525000 ;
      RECT   96.285000 -0.085000   96.455000 0.085000 ;
      RECT   96.285000  2.635000   96.455000 2.805000 ;
      RECT   96.285000  5.355000   96.455000 5.525000 ;
      RECT   96.745000 -0.085000   96.915000 0.085000 ;
      RECT   96.745000  2.635000   96.915000 2.805000 ;
      RECT   96.745000  5.355000   96.915000 5.525000 ;
      RECT   97.205000 -0.085000   97.375000 0.085000 ;
      RECT   97.205000  2.635000   97.375000 2.805000 ;
      RECT   97.205000  5.355000   97.375000 5.525000 ;
      RECT   97.665000 -0.085000   97.835000 0.085000 ;
      RECT   97.665000  2.635000   97.835000 2.805000 ;
      RECT   97.665000  5.355000   97.835000 5.525000 ;
      RECT   98.125000 -0.085000   98.295000 0.085000 ;
      RECT   98.125000  2.635000   98.295000 2.805000 ;
      RECT   98.125000  5.355000   98.295000 5.525000 ;
      RECT   98.585000 -0.085000   98.755000 0.085000 ;
      RECT   98.585000  2.635000   98.755000 2.805000 ;
      RECT   98.585000  5.355000   98.755000 5.525000 ;
      RECT   99.045000 -0.085000   99.215000 0.085000 ;
      RECT   99.045000  2.635000   99.215000 2.805000 ;
      RECT   99.045000  5.355000   99.215000 5.525000 ;
      RECT   99.505000 -0.085000   99.675000 0.085000 ;
      RECT   99.505000  2.635000   99.675000 2.805000 ;
      RECT   99.505000  5.355000   99.675000 5.525000 ;
      RECT   99.965000 -0.085000  100.135000 0.085000 ;
      RECT   99.965000  2.635000  100.135000 2.805000 ;
      RECT   99.965000  5.355000  100.135000 5.525000 ;
      RECT  100.425000 -0.085000  100.595000 0.085000 ;
      RECT  100.425000  2.635000  100.595000 2.805000 ;
      RECT  100.425000  5.355000  100.595000 5.525000 ;
      RECT  100.885000 -0.085000  101.055000 0.085000 ;
      RECT  100.885000  2.635000  101.055000 2.805000 ;
      RECT  100.885000  5.355000  101.055000 5.525000 ;
      RECT  101.345000 -0.085000  101.515000 0.085000 ;
      RECT  101.345000  2.635000  101.515000 2.805000 ;
      RECT  101.345000  5.355000  101.515000 5.525000 ;
      RECT  101.805000 -0.085000  101.975000 0.085000 ;
      RECT  101.805000  2.635000  101.975000 2.805000 ;
      RECT  101.805000  5.355000  101.975000 5.525000 ;
      RECT  102.265000 -0.085000  102.435000 0.085000 ;
      RECT  102.265000  2.635000  102.435000 2.805000 ;
      RECT  102.265000  5.355000  102.435000 5.525000 ;
      RECT  102.725000 -0.085000  102.895000 0.085000 ;
      RECT  102.725000  2.635000  102.895000 2.805000 ;
      RECT  102.725000  5.355000  102.895000 5.525000 ;
      RECT  103.185000 -0.085000  103.355000 0.085000 ;
      RECT  103.185000  2.635000  103.355000 2.805000 ;
      RECT  103.185000  5.355000  103.355000 5.525000 ;
      RECT  103.645000 -0.085000  103.815000 0.085000 ;
      RECT  103.645000  2.635000  103.815000 2.805000 ;
      RECT  103.645000  5.355000  103.815000 5.525000 ;
      RECT  104.105000 -0.085000  104.275000 0.085000 ;
      RECT  104.105000  2.635000  104.275000 2.805000 ;
      RECT  104.105000  5.355000  104.275000 5.525000 ;
      RECT  104.565000 -0.085000  104.735000 0.085000 ;
      RECT  104.565000  2.635000  104.735000 2.805000 ;
      RECT  104.565000  5.355000  104.735000 5.525000 ;
      RECT  105.025000 -0.085000  105.195000 0.085000 ;
      RECT  105.025000  2.635000  105.195000 2.805000 ;
      RECT  105.025000  5.355000  105.195000 5.525000 ;
      RECT  105.485000 -0.085000  105.655000 0.085000 ;
      RECT  105.485000  2.635000  105.655000 2.805000 ;
      RECT  105.485000  5.355000  105.655000 5.525000 ;
      RECT  105.945000 -0.085000  106.115000 0.085000 ;
      RECT  105.945000  2.635000  106.115000 2.805000 ;
      RECT  105.945000  5.355000  106.115000 5.525000 ;
      RECT  106.405000 -0.085000  106.575000 0.085000 ;
      RECT  106.405000  2.635000  106.575000 2.805000 ;
      RECT  106.405000  5.355000  106.575000 5.525000 ;
      RECT  106.865000 -0.085000  107.035000 0.085000 ;
      RECT  106.865000  2.635000  107.035000 2.805000 ;
      RECT  106.865000  5.355000  107.035000 5.525000 ;
      RECT  107.325000 -0.085000  107.495000 0.085000 ;
      RECT  107.325000  2.635000  107.495000 2.805000 ;
      RECT  107.325000  5.355000  107.495000 5.525000 ;
      RECT  107.785000 -0.085000  107.955000 0.085000 ;
      RECT  107.785000  2.635000  107.955000 2.805000 ;
      RECT  107.785000  5.355000  107.955000 5.525000 ;
      RECT  108.245000 -0.085000  108.415000 0.085000 ;
      RECT  108.245000  2.635000  108.415000 2.805000 ;
      RECT  108.245000  5.355000  108.415000 5.525000 ;
      RECT  108.705000 -0.085000  108.875000 0.085000 ;
      RECT  108.705000  2.635000  108.875000 2.805000 ;
      RECT  108.705000  5.355000  108.875000 5.525000 ;
      RECT  109.165000 -0.085000  109.335000 0.085000 ;
      RECT  109.165000  2.635000  109.335000 2.805000 ;
      RECT  109.165000  5.355000  109.335000 5.525000 ;
      RECT  109.625000 -0.085000  109.795000 0.085000 ;
      RECT  109.625000  2.635000  109.795000 2.805000 ;
      RECT  109.625000  5.355000  109.795000 5.525000 ;
      RECT  110.085000 -0.085000  110.255000 0.085000 ;
      RECT  110.085000  2.635000  110.255000 2.805000 ;
      RECT  110.085000  5.355000  110.255000 5.525000 ;
      RECT  110.545000 -0.085000  110.715000 0.085000 ;
      RECT  110.545000  2.635000  110.715000 2.805000 ;
      RECT  110.545000  5.355000  110.715000 5.525000 ;
      RECT  111.005000 -0.085000  111.175000 0.085000 ;
      RECT  111.005000  2.635000  111.175000 2.805000 ;
      RECT  111.005000  5.355000  111.175000 5.525000 ;
      RECT  111.465000 -0.085000  111.635000 0.085000 ;
      RECT  111.465000  2.635000  111.635000 2.805000 ;
      RECT  111.465000  5.355000  111.635000 5.525000 ;
      RECT  111.925000 -0.085000  112.095000 0.085000 ;
      RECT  111.925000  2.635000  112.095000 2.805000 ;
      RECT  111.925000  5.355000  112.095000 5.525000 ;
      RECT  112.385000 -0.085000  112.555000 0.085000 ;
      RECT  112.385000  2.635000  112.555000 2.805000 ;
      RECT  112.385000  5.355000  112.555000 5.525000 ;
      RECT  112.845000 -0.085000  113.015000 0.085000 ;
      RECT  112.845000  2.635000  113.015000 2.805000 ;
      RECT  112.845000  5.355000  113.015000 5.525000 ;
      RECT  113.305000 -0.085000  113.475000 0.085000 ;
      RECT  113.305000  2.635000  113.475000 2.805000 ;
      RECT  113.305000  5.355000  113.475000 5.525000 ;
      RECT  113.765000 -0.085000  113.935000 0.085000 ;
      RECT  113.765000  2.635000  113.935000 2.805000 ;
      RECT  113.765000  5.355000  113.935000 5.525000 ;
      RECT  114.225000 -0.085000  114.395000 0.085000 ;
      RECT  114.225000  2.635000  114.395000 2.805000 ;
      RECT  114.225000  5.355000  114.395000 5.525000 ;
      RECT  114.685000 -0.085000  114.855000 0.085000 ;
      RECT  114.685000  2.635000  114.855000 2.805000 ;
      RECT  114.685000  5.355000  114.855000 5.525000 ;
      RECT  115.145000 -0.085000  115.315000 0.085000 ;
      RECT  115.145000  2.635000  115.315000 2.805000 ;
      RECT  115.145000  5.355000  115.315000 5.525000 ;
      RECT  115.605000 -0.085000  115.775000 0.085000 ;
      RECT  115.605000  2.635000  115.775000 2.805000 ;
      RECT  115.605000  5.355000  115.775000 5.525000 ;
      RECT  116.065000 -0.085000  116.235000 0.085000 ;
      RECT  116.065000  2.635000  116.235000 2.805000 ;
      RECT  116.065000  5.355000  116.235000 5.525000 ;
      RECT  116.525000 -0.085000  116.695000 0.085000 ;
      RECT  116.525000  2.635000  116.695000 2.805000 ;
      RECT  116.525000  5.355000  116.695000 5.525000 ;
      RECT  116.985000 -0.085000  117.155000 0.085000 ;
      RECT  116.985000  2.635000  117.155000 2.805000 ;
      RECT  116.985000  5.355000  117.155000 5.525000 ;
      RECT  117.445000 -0.085000  117.615000 0.085000 ;
      RECT  117.445000  2.635000  117.615000 2.805000 ;
      RECT  117.445000  5.355000  117.615000 5.525000 ;
      RECT  117.905000 -0.085000  118.075000 0.085000 ;
      RECT  117.905000  2.635000  118.075000 2.805000 ;
      RECT  117.905000  5.355000  118.075000 5.525000 ;
      RECT  118.365000 -0.085000  118.535000 0.085000 ;
      RECT  118.365000  2.635000  118.535000 2.805000 ;
      RECT  118.365000  5.355000  118.535000 5.525000 ;
      RECT  118.825000 -0.085000  118.995000 0.085000 ;
      RECT  118.825000  2.635000  118.995000 2.805000 ;
      RECT  118.825000  5.355000  118.995000 5.525000 ;
      RECT  119.285000 -0.085000  119.455000 0.085000 ;
      RECT  119.285000  2.635000  119.455000 2.805000 ;
      RECT  119.285000  5.355000  119.455000 5.525000 ;
      RECT  119.745000 -0.085000  119.915000 0.085000 ;
      RECT  119.745000  2.635000  119.915000 2.805000 ;
      RECT  119.745000  5.355000  119.915000 5.525000 ;
      RECT  120.205000 -0.085000  120.375000 0.085000 ;
      RECT  120.205000  2.635000  120.375000 2.805000 ;
      RECT  120.205000  5.355000  120.375000 5.525000 ;
      RECT  120.665000 -0.085000  120.835000 0.085000 ;
      RECT  120.665000  2.635000  120.835000 2.805000 ;
      RECT  120.665000  5.355000  120.835000 5.525000 ;
      RECT  121.125000 -0.085000  121.295000 0.085000 ;
      RECT  121.125000  2.635000  121.295000 2.805000 ;
      RECT  121.125000  5.355000  121.295000 5.525000 ;
      RECT  121.585000 -0.085000  121.755000 0.085000 ;
      RECT  121.585000  2.635000  121.755000 2.805000 ;
      RECT  121.585000  5.355000  121.755000 5.525000 ;
      RECT  122.045000 -0.085000  122.215000 0.085000 ;
      RECT  122.045000  2.635000  122.215000 2.805000 ;
      RECT  122.045000  5.355000  122.215000 5.525000 ;
      RECT  122.505000 -0.085000  122.675000 0.085000 ;
      RECT  122.505000  2.635000  122.675000 2.805000 ;
      RECT  122.505000  5.355000  122.675000 5.525000 ;
      RECT  122.965000 -0.085000  123.135000 0.085000 ;
      RECT  122.965000  2.635000  123.135000 2.805000 ;
      RECT  122.965000  5.355000  123.135000 5.525000 ;
      RECT  123.425000 -0.085000  123.595000 0.085000 ;
      RECT  123.425000  2.635000  123.595000 2.805000 ;
      RECT  123.425000  5.355000  123.595000 5.525000 ;
      RECT  123.885000 -0.085000  124.055000 0.085000 ;
      RECT  123.885000  2.635000  124.055000 2.805000 ;
      RECT  123.885000  5.355000  124.055000 5.525000 ;
      RECT  124.345000 -0.085000  124.515000 0.085000 ;
      RECT  124.345000  2.635000  124.515000 2.805000 ;
      RECT  124.345000  5.355000  124.515000 5.525000 ;
      RECT  124.805000 -0.085000  124.975000 0.085000 ;
      RECT  124.805000  2.635000  124.975000 2.805000 ;
      RECT  124.805000  5.355000  124.975000 5.525000 ;
      RECT  125.265000 -0.085000  125.435000 0.085000 ;
      RECT  125.265000  2.635000  125.435000 2.805000 ;
      RECT  125.265000  5.355000  125.435000 5.525000 ;
      RECT  125.725000 -0.085000  125.895000 0.085000 ;
      RECT  125.725000  2.635000  125.895000 2.805000 ;
      RECT  125.725000  5.355000  125.895000 5.525000 ;
      RECT  126.185000 -0.085000  126.355000 0.085000 ;
      RECT  126.185000  2.635000  126.355000 2.805000 ;
      RECT  126.185000  5.355000  126.355000 5.525000 ;
      RECT  126.645000 -0.085000  126.815000 0.085000 ;
      RECT  126.645000  2.635000  126.815000 2.805000 ;
      RECT  126.645000  5.355000  126.815000 5.525000 ;
      RECT  127.105000 -0.085000  127.275000 0.085000 ;
      RECT  127.105000  2.635000  127.275000 2.805000 ;
      RECT  127.105000  5.355000  127.275000 5.525000 ;
      RECT  127.565000 -0.085000  127.735000 0.085000 ;
      RECT  127.565000  2.635000  127.735000 2.805000 ;
      RECT  127.565000  5.355000  127.735000 5.525000 ;
      RECT  128.025000 -0.085000  128.195000 0.085000 ;
      RECT  128.025000  2.635000  128.195000 2.805000 ;
      RECT  128.025000  5.355000  128.195000 5.525000 ;
      RECT  128.485000 -0.085000  128.655000 0.085000 ;
      RECT  128.485000  2.635000  128.655000 2.805000 ;
      RECT  128.485000  5.355000  128.655000 5.525000 ;
      RECT  128.945000 -0.085000  129.115000 0.085000 ;
      RECT  128.945000  2.635000  129.115000 2.805000 ;
      RECT  128.945000  5.355000  129.115000 5.525000 ;
      RECT  129.405000 -0.085000  129.575000 0.085000 ;
      RECT  129.405000  2.635000  129.575000 2.805000 ;
      RECT  129.405000  5.355000  129.575000 5.525000 ;
      RECT  129.865000 -0.085000  130.035000 0.085000 ;
      RECT  129.865000  2.635000  130.035000 2.805000 ;
      RECT  129.865000  5.355000  130.035000 5.525000 ;
      RECT  130.325000 -0.085000  130.495000 0.085000 ;
      RECT  130.325000  2.635000  130.495000 2.805000 ;
      RECT  130.325000  5.355000  130.495000 5.525000 ;
      RECT  130.785000 -0.085000  130.955000 0.085000 ;
      RECT  130.785000  2.635000  130.955000 2.805000 ;
      RECT  130.785000  5.355000  130.955000 5.525000 ;
      RECT  131.245000 -0.085000  131.415000 0.085000 ;
      RECT  131.245000  2.635000  131.415000 2.805000 ;
      RECT  131.245000  5.355000  131.415000 5.525000 ;
      RECT  131.705000 -0.085000  131.875000 0.085000 ;
      RECT  131.705000  2.635000  131.875000 2.805000 ;
      RECT  131.705000  5.355000  131.875000 5.525000 ;
      RECT  132.165000 -0.085000  132.335000 0.085000 ;
      RECT  132.165000  2.635000  132.335000 2.805000 ;
      RECT  132.165000  5.355000  132.335000 5.525000 ;
      RECT  132.625000 -0.085000  132.795000 0.085000 ;
      RECT  132.625000  2.635000  132.795000 2.805000 ;
      RECT  132.625000  5.355000  132.795000 5.525000 ;
      RECT  133.085000 -0.085000  133.255000 0.085000 ;
      RECT  133.085000  2.635000  133.255000 2.805000 ;
      RECT  133.085000  5.355000  133.255000 5.525000 ;
      RECT  133.545000 -0.085000  133.715000 0.085000 ;
      RECT  133.545000  2.635000  133.715000 2.805000 ;
      RECT  133.545000  5.355000  133.715000 5.525000 ;
      RECT  134.005000 -0.085000  134.175000 0.085000 ;
      RECT  134.005000  2.635000  134.175000 2.805000 ;
      RECT  134.005000  5.355000  134.175000 5.525000 ;
      RECT  134.465000 -0.085000  134.635000 0.085000 ;
      RECT  134.465000  2.635000  134.635000 2.805000 ;
      RECT  134.465000  5.355000  134.635000 5.525000 ;
      RECT  134.925000 -0.085000  135.095000 0.085000 ;
      RECT  134.925000  2.635000  135.095000 2.805000 ;
      RECT  134.925000  5.355000  135.095000 5.525000 ;
      RECT  135.385000 -0.085000  135.555000 0.085000 ;
      RECT  135.385000  2.635000  135.555000 2.805000 ;
      RECT  135.385000  5.355000  135.555000 5.525000 ;
      RECT  135.845000 -0.085000  136.015000 0.085000 ;
      RECT  135.845000  2.635000  136.015000 2.805000 ;
      RECT  135.845000  5.355000  136.015000 5.525000 ;
      RECT  136.305000 -0.085000  136.475000 0.085000 ;
      RECT  136.305000  2.635000  136.475000 2.805000 ;
      RECT  136.305000  5.355000  136.475000 5.525000 ;
      RECT  136.765000 -0.085000  136.935000 0.085000 ;
      RECT  136.765000  2.635000  136.935000 2.805000 ;
      RECT  136.765000  5.355000  136.935000 5.525000 ;
      RECT  137.225000 -0.085000  137.395000 0.085000 ;
      RECT  137.225000  2.635000  137.395000 2.805000 ;
      RECT  137.225000  5.355000  137.395000 5.525000 ;
      RECT  137.685000 -0.085000  137.855000 0.085000 ;
      RECT  137.685000  2.635000  137.855000 2.805000 ;
      RECT  137.685000  5.355000  137.855000 5.525000 ;
      RECT  138.145000 -0.085000  138.315000 0.085000 ;
      RECT  138.145000  2.635000  138.315000 2.805000 ;
      RECT  138.145000  5.355000  138.315000 5.525000 ;
      RECT  138.605000 -0.085000  138.775000 0.085000 ;
      RECT  138.605000  2.635000  138.775000 2.805000 ;
      RECT  138.605000  5.355000  138.775000 5.525000 ;
      RECT  139.065000 -0.085000  139.235000 0.085000 ;
      RECT  139.065000  2.635000  139.235000 2.805000 ;
      RECT  139.065000  5.355000  139.235000 5.525000 ;
      RECT  139.525000 -0.085000  139.695000 0.085000 ;
      RECT  139.525000  2.635000  139.695000 2.805000 ;
      RECT  139.525000  5.355000  139.695000 5.525000 ;
      RECT  139.985000 -0.085000  140.155000 0.085000 ;
      RECT  139.985000  2.635000  140.155000 2.805000 ;
      RECT  139.985000  5.355000  140.155000 5.525000 ;
      RECT  140.445000 -0.085000  140.615000 0.085000 ;
      RECT  140.445000  2.635000  140.615000 2.805000 ;
      RECT  140.445000  5.355000  140.615000 5.525000 ;
      RECT  140.905000 -0.085000  141.075000 0.085000 ;
      RECT  140.905000  2.635000  141.075000 2.805000 ;
      RECT  140.905000  5.355000  141.075000 5.525000 ;
      RECT  141.365000 -0.085000  141.535000 0.085000 ;
      RECT  141.365000  2.635000  141.535000 2.805000 ;
      RECT  141.365000  5.355000  141.535000 5.525000 ;
      RECT  141.825000 -0.085000  141.995000 0.085000 ;
      RECT  141.825000  2.635000  141.995000 2.805000 ;
      RECT  141.825000  5.355000  141.995000 5.525000 ;
      RECT  142.285000 -0.085000  142.455000 0.085000 ;
      RECT  142.285000  2.635000  142.455000 2.805000 ;
      RECT  142.285000  5.355000  142.455000 5.525000 ;
      RECT  142.745000 -0.085000  142.915000 0.085000 ;
      RECT  142.745000  2.635000  142.915000 2.805000 ;
      RECT  142.745000  5.355000  142.915000 5.525000 ;
      RECT  143.205000 -0.085000  143.375000 0.085000 ;
      RECT  143.205000  2.635000  143.375000 2.805000 ;
      RECT  143.205000  5.355000  143.375000 5.525000 ;
      RECT  143.665000 -0.085000  143.835000 0.085000 ;
      RECT  143.665000  2.635000  143.835000 2.805000 ;
      RECT  143.665000  5.355000  143.835000 5.525000 ;
      RECT  144.125000 -0.085000  144.295000 0.085000 ;
      RECT  144.125000  2.635000  144.295000 2.805000 ;
      RECT  144.125000  5.355000  144.295000 5.525000 ;
      RECT  144.585000 -0.085000  144.755000 0.085000 ;
      RECT  144.585000  2.635000  144.755000 2.805000 ;
      RECT  144.585000  5.355000  144.755000 5.525000 ;
      RECT  145.045000 -0.085000  145.215000 0.085000 ;
      RECT  145.045000  2.635000  145.215000 2.805000 ;
      RECT  145.045000  5.355000  145.215000 5.525000 ;
      RECT  145.505000 -0.085000  145.675000 0.085000 ;
      RECT  145.505000  2.635000  145.675000 2.805000 ;
      RECT  145.505000  5.355000  145.675000 5.525000 ;
      RECT  145.965000 -0.085000  146.135000 0.085000 ;
      RECT  145.965000  2.635000  146.135000 2.805000 ;
      RECT  145.965000  5.355000  146.135000 5.525000 ;
      RECT  146.425000 -0.085000  146.595000 0.085000 ;
      RECT  146.425000  2.635000  146.595000 2.805000 ;
      RECT  146.425000  5.355000  146.595000 5.525000 ;
      RECT  146.885000 -0.085000  147.055000 0.085000 ;
      RECT  146.885000  2.635000  147.055000 2.805000 ;
      RECT  146.885000  5.355000  147.055000 5.525000 ;
      RECT  147.345000 -0.085000  147.515000 0.085000 ;
      RECT  147.345000  2.635000  147.515000 2.805000 ;
      RECT  147.345000  5.355000  147.515000 5.525000 ;
      RECT  147.805000 -0.085000  147.975000 0.085000 ;
      RECT  147.805000  2.635000  147.975000 2.805000 ;
      RECT  147.805000  5.355000  147.975000 5.525000 ;
      RECT  148.265000 -0.085000  148.435000 0.085000 ;
      RECT  148.265000  2.635000  148.435000 2.805000 ;
      RECT  148.265000  5.355000  148.435000 5.525000 ;
      RECT  148.725000 -0.085000  148.895000 0.085000 ;
      RECT  148.725000  2.635000  148.895000 2.805000 ;
      RECT  148.725000  5.355000  148.895000 5.525000 ;
      RECT  149.185000 -0.085000  149.355000 0.085000 ;
      RECT  149.185000  2.635000  149.355000 2.805000 ;
      RECT  149.185000  5.355000  149.355000 5.525000 ;
      RECT  149.645000 -0.085000  149.815000 0.085000 ;
      RECT  149.645000  2.635000  149.815000 2.805000 ;
      RECT  149.645000  5.355000  149.815000 5.525000 ;
      RECT  150.105000 -0.085000  150.275000 0.085000 ;
      RECT  150.105000  2.635000  150.275000 2.805000 ;
      RECT  150.105000  5.355000  150.275000 5.525000 ;
      RECT  150.565000 -0.085000  150.735000 0.085000 ;
      RECT  150.565000  2.635000  150.735000 2.805000 ;
      RECT  150.565000  5.355000  150.735000 5.525000 ;
      RECT  151.025000 -0.085000  151.195000 0.085000 ;
      RECT  151.025000  2.635000  151.195000 2.805000 ;
      RECT  151.025000  5.355000  151.195000 5.525000 ;
      RECT  151.485000 -0.085000  151.655000 0.085000 ;
      RECT  151.485000  2.635000  151.655000 2.805000 ;
      RECT  151.485000  5.355000  151.655000 5.525000 ;
      RECT  151.945000 -0.085000  152.115000 0.085000 ;
      RECT  151.945000  2.635000  152.115000 2.805000 ;
      RECT  151.945000  5.355000  152.115000 5.525000 ;
      RECT  152.405000 -0.085000  152.575000 0.085000 ;
      RECT  152.405000  2.635000  152.575000 2.805000 ;
      RECT  152.405000  5.355000  152.575000 5.525000 ;
      RECT  152.865000 -0.085000  153.035000 0.085000 ;
      RECT  152.865000  2.635000  153.035000 2.805000 ;
      RECT  152.865000  5.355000  153.035000 5.525000 ;
      RECT  153.325000 -0.085000  153.495000 0.085000 ;
      RECT  153.325000  2.635000  153.495000 2.805000 ;
      RECT  153.325000  5.355000  153.495000 5.525000 ;
      RECT  153.785000 -0.085000  153.955000 0.085000 ;
      RECT  153.785000  2.635000  153.955000 2.805000 ;
      RECT  153.785000  5.355000  153.955000 5.525000 ;
      RECT  154.245000 -0.085000  154.415000 0.085000 ;
      RECT  154.245000  2.635000  154.415000 2.805000 ;
      RECT  154.245000  5.355000  154.415000 5.525000 ;
      RECT  154.705000 -0.085000  154.875000 0.085000 ;
      RECT  154.705000  2.635000  154.875000 2.805000 ;
      RECT  154.705000  5.355000  154.875000 5.525000 ;
      RECT  155.165000 -0.085000  155.335000 0.085000 ;
      RECT  155.165000  2.635000  155.335000 2.805000 ;
      RECT  155.165000  5.355000  155.335000 5.525000 ;
      RECT  155.625000 -0.085000  155.795000 0.085000 ;
      RECT  155.625000  2.635000  155.795000 2.805000 ;
      RECT  155.625000  5.355000  155.795000 5.525000 ;
      RECT  156.085000 -0.085000  156.255000 0.085000 ;
      RECT  156.085000  2.635000  156.255000 2.805000 ;
      RECT  156.085000  5.355000  156.255000 5.525000 ;
      RECT  156.545000 -0.085000  156.715000 0.085000 ;
      RECT  156.545000  2.635000  156.715000 2.805000 ;
      RECT  156.545000  5.355000  156.715000 5.525000 ;
      RECT  157.005000 -0.085000  157.175000 0.085000 ;
      RECT  157.005000  2.635000  157.175000 2.805000 ;
      RECT  157.005000  5.355000  157.175000 5.525000 ;
      RECT  157.280000  4.165000  157.450000 4.335000 ;
      RECT  157.465000 -0.085000  157.635000 0.085000 ;
      RECT  157.465000  2.635000  157.635000 2.805000 ;
      RECT  157.465000  5.355000  157.635000 5.525000 ;
      RECT  157.640000  4.165000  157.810000 4.335000 ;
      RECT  157.925000 -0.085000  158.095000 0.085000 ;
      RECT  157.925000  2.635000  158.095000 2.805000 ;
      RECT  157.925000  5.355000  158.095000 5.525000 ;
      RECT  158.385000 -0.085000  158.555000 0.085000 ;
      RECT  158.385000  2.635000  158.555000 2.805000 ;
      RECT  158.385000  5.355000  158.555000 5.525000 ;
      RECT  158.845000 -0.085000  159.015000 0.085000 ;
      RECT  158.845000  2.635000  159.015000 2.805000 ;
      RECT  158.845000  5.355000  159.015000 5.525000 ;
      RECT  159.305000 -0.085000  159.475000 0.085000 ;
      RECT  159.305000  2.635000  159.475000 2.805000 ;
      RECT  159.305000  5.355000  159.475000 5.525000 ;
      RECT  159.765000 -0.085000  159.935000 0.085000 ;
      RECT  159.765000  2.635000  159.935000 2.805000 ;
      RECT  159.765000  5.355000  159.935000 5.525000 ;
      RECT  160.225000 -0.085000  160.395000 0.085000 ;
      RECT  160.225000  2.635000  160.395000 2.805000 ;
      RECT  160.225000  5.355000  160.395000 5.525000 ;
      RECT  160.685000 -0.085000  160.855000 0.085000 ;
      RECT  160.685000  2.635000  160.855000 2.805000 ;
      RECT  160.685000  5.355000  160.855000 5.525000 ;
      RECT  161.145000 -0.085000  161.315000 0.085000 ;
      RECT  161.145000  2.635000  161.315000 2.805000 ;
      RECT  161.145000  5.355000  161.315000 5.525000 ;
      RECT  161.605000 -0.085000  161.775000 0.085000 ;
      RECT  161.605000  2.635000  161.775000 2.805000 ;
      RECT  161.605000  5.355000  161.775000 5.525000 ;
      RECT  162.065000 -0.085000  162.235000 0.085000 ;
      RECT  162.065000  2.635000  162.235000 2.805000 ;
      RECT  162.065000  5.355000  162.235000 5.525000 ;
      RECT  162.525000 -0.085000  162.695000 0.085000 ;
      RECT  162.525000  2.635000  162.695000 2.805000 ;
      RECT  162.525000  5.355000  162.695000 5.525000 ;
      RECT  162.985000 -0.085000  163.155000 0.085000 ;
      RECT  162.985000  2.635000  163.155000 2.805000 ;
      RECT  162.985000  5.355000  163.155000 5.525000 ;
      RECT  163.445000 -0.085000  163.615000 0.085000 ;
      RECT  163.445000  2.635000  163.615000 2.805000 ;
      RECT  163.445000  5.355000  163.615000 5.525000 ;
      RECT  163.905000 -0.085000  164.075000 0.085000 ;
      RECT  163.905000  2.635000  164.075000 2.805000 ;
      RECT  163.905000  5.355000  164.075000 5.525000 ;
      RECT  164.365000 -0.085000  164.535000 0.085000 ;
      RECT  164.365000  2.635000  164.535000 2.805000 ;
      RECT  164.365000  5.355000  164.535000 5.525000 ;
      RECT  164.825000 -0.085000  164.995000 0.085000 ;
      RECT  164.825000  2.635000  164.995000 2.805000 ;
      RECT  164.825000  5.355000  164.995000 5.525000 ;
      RECT  165.285000 -0.085000  165.455000 0.085000 ;
      RECT  165.285000  2.635000  165.455000 2.805000 ;
      RECT  165.285000  5.355000  165.455000 5.525000 ;
      RECT  165.745000 -0.085000  165.915000 0.085000 ;
      RECT  165.745000  2.635000  165.915000 2.805000 ;
      RECT  165.745000  5.355000  165.915000 5.525000 ;
      RECT  166.205000 -0.085000  166.375000 0.085000 ;
      RECT  166.205000  2.635000  166.375000 2.805000 ;
      RECT  166.205000  3.145000  166.375000 3.315000 ;
      RECT  166.205000  5.355000  166.375000 5.525000 ;
      RECT  166.665000 -0.085000  166.835000 0.085000 ;
      RECT  166.665000  2.635000  166.835000 2.805000 ;
      RECT  166.665000  3.485000  166.835000 3.655000 ;
      RECT  166.665000  5.355000  166.835000 5.525000 ;
      RECT  167.125000 -0.085000  167.295000 0.085000 ;
      RECT  167.125000  2.635000  167.295000 2.805000 ;
      RECT  167.125000  5.355000  167.295000 5.525000 ;
      RECT  167.585000 -0.085000  167.755000 0.085000 ;
      RECT  167.585000  2.635000  167.755000 2.805000 ;
      RECT  167.585000  5.355000  167.755000 5.525000 ;
      RECT  167.840000  1.445000  168.010000 1.615000 ;
      RECT  168.045000 -0.085000  168.215000 0.085000 ;
      RECT  168.045000  2.635000  168.215000 2.805000 ;
      RECT  168.045000  5.355000  168.215000 5.525000 ;
      RECT  168.505000 -0.085000  168.675000 0.085000 ;
      RECT  168.505000  2.635000  168.675000 2.805000 ;
      RECT  168.505000  5.355000  168.675000 5.525000 ;
      RECT  168.965000 -0.085000  169.135000 0.085000 ;
      RECT  168.965000  2.635000  169.135000 2.805000 ;
      RECT  168.965000  5.355000  169.135000 5.525000 ;
      RECT  169.425000 -0.085000  169.595000 0.085000 ;
      RECT  169.425000  2.635000  169.595000 2.805000 ;
      RECT  169.425000  5.355000  169.595000 5.525000 ;
      RECT  169.885000 -0.085000  170.055000 0.085000 ;
      RECT  169.885000  2.635000  170.055000 2.805000 ;
      RECT  169.885000  5.355000  170.055000 5.525000 ;
      RECT  170.345000 -0.085000  170.515000 0.085000 ;
      RECT  170.345000  2.635000  170.515000 2.805000 ;
      RECT  170.345000  5.355000  170.515000 5.525000 ;
      RECT  170.805000 -0.085000  170.975000 0.085000 ;
      RECT  170.805000  2.635000  170.975000 2.805000 ;
      RECT  170.805000  5.355000  170.975000 5.525000 ;
      RECT  170.870000  1.445000  171.040000 1.615000 ;
      RECT  171.265000 -0.085000  171.435000 0.085000 ;
      RECT  171.265000  2.635000  171.435000 2.805000 ;
      RECT  171.265000  5.355000  171.435000 5.525000 ;
      RECT  171.725000 -0.085000  171.895000 0.085000 ;
      RECT  171.725000  2.635000  171.895000 2.805000 ;
      RECT  171.725000  5.355000  171.895000 5.525000 ;
      RECT  172.185000 -0.085000  172.355000 0.085000 ;
      RECT  172.185000  2.635000  172.355000 2.805000 ;
      RECT  172.185000  5.355000  172.355000 5.525000 ;
      RECT  172.645000 -0.085000  172.815000 0.085000 ;
      RECT  172.645000  2.635000  172.815000 2.805000 ;
      RECT  172.645000  5.355000  172.815000 5.525000 ;
      RECT  173.105000 -0.085000  173.275000 0.085000 ;
      RECT  173.105000  2.635000  173.275000 2.805000 ;
      RECT  173.105000  5.355000  173.275000 5.525000 ;
      RECT  173.565000 -0.085000  173.735000 0.085000 ;
      RECT  173.565000  2.635000  173.735000 2.805000 ;
      RECT  173.565000  5.355000  173.735000 5.525000 ;
      RECT  174.025000 -0.085000  174.195000 0.085000 ;
      RECT  174.025000  2.635000  174.195000 2.805000 ;
      RECT  174.025000  5.355000  174.195000 5.525000 ;
      RECT  174.485000 -0.085000  174.655000 0.085000 ;
      RECT  174.485000  2.635000  174.655000 2.805000 ;
      RECT  174.485000  5.355000  174.655000 5.525000 ;
      RECT  174.945000 -0.085000  175.115000 0.085000 ;
      RECT  174.945000  2.635000  175.115000 2.805000 ;
      RECT  174.945000  5.355000  175.115000 5.525000 ;
      RECT  175.405000 -0.085000  175.575000 0.085000 ;
      RECT  175.405000  2.635000  175.575000 2.805000 ;
      RECT  175.405000  5.355000  175.575000 5.525000 ;
      RECT  175.865000 -0.085000  176.035000 0.085000 ;
      RECT  175.865000  2.635000  176.035000 2.805000 ;
      RECT  175.865000  5.355000  176.035000 5.525000 ;
      RECT  176.325000 -0.085000  176.495000 0.085000 ;
      RECT  176.325000  2.635000  176.495000 2.805000 ;
      RECT  176.325000  5.355000  176.495000 5.525000 ;
      RECT  176.785000 -0.085000  176.955000 0.085000 ;
      RECT  176.785000  2.635000  176.955000 2.805000 ;
      RECT  176.785000  5.355000  176.955000 5.525000 ;
      RECT  177.245000 -0.085000  177.415000 0.085000 ;
      RECT  177.245000  2.635000  177.415000 2.805000 ;
      RECT  177.245000  5.355000  177.415000 5.525000 ;
      RECT  177.705000 -0.085000  177.875000 0.085000 ;
      RECT  177.705000  2.635000  177.875000 2.805000 ;
      RECT  177.705000  5.355000  177.875000 5.525000 ;
      RECT  177.725000  4.165000  177.895000 4.335000 ;
      RECT  178.085000  4.165000  178.255000 4.335000 ;
      RECT  178.165000 -0.085000  178.335000 0.085000 ;
      RECT  178.165000  2.635000  178.335000 2.805000 ;
      RECT  178.165000  5.355000  178.335000 5.525000 ;
      RECT  178.625000 -0.085000  178.795000 0.085000 ;
      RECT  178.625000  2.635000  178.795000 2.805000 ;
      RECT  178.625000  5.355000  178.795000 5.525000 ;
      RECT  179.085000 -0.085000  179.255000 0.085000 ;
      RECT  179.085000  2.635000  179.255000 2.805000 ;
      RECT  179.085000  5.355000  179.255000 5.525000 ;
      RECT  179.545000 -0.085000  179.715000 0.085000 ;
      RECT  179.545000  2.635000  179.715000 2.805000 ;
      RECT  179.545000  5.355000  179.715000 5.525000 ;
      RECT  180.005000 -0.085000  180.175000 0.085000 ;
      RECT  180.005000  2.635000  180.175000 2.805000 ;
      RECT  180.005000  5.355000  180.175000 5.525000 ;
      RECT  180.465000 -0.085000  180.635000 0.085000 ;
      RECT  180.465000  2.635000  180.635000 2.805000 ;
      RECT  180.465000  5.355000  180.635000 5.525000 ;
      RECT  180.495000  3.485000  180.665000 3.655000 ;
      RECT  180.925000 -0.085000  181.095000 0.085000 ;
      RECT  180.925000  2.635000  181.095000 2.805000 ;
      RECT  180.925000  5.355000  181.095000 5.525000 ;
      RECT  180.955000  3.825000  181.125000 3.995000 ;
      RECT  181.385000 -0.085000  181.555000 0.085000 ;
      RECT  181.385000  2.635000  181.555000 2.805000 ;
      RECT  181.385000  5.355000  181.555000 5.525000 ;
      RECT  181.845000 -0.085000  182.015000 0.085000 ;
      RECT  181.845000  2.635000  182.015000 2.805000 ;
      RECT  181.845000  5.355000  182.015000 5.525000 ;
      RECT  182.305000 -0.085000  182.475000 0.085000 ;
      RECT  182.305000  2.635000  182.475000 2.805000 ;
      RECT  182.305000  5.355000  182.475000 5.525000 ;
      RECT  182.585000  3.825000  182.755000 3.995000 ;
      RECT  182.765000 -0.085000  182.935000 0.085000 ;
      RECT  182.765000  2.635000  182.935000 2.805000 ;
      RECT  182.765000  5.355000  182.935000 5.525000 ;
      RECT  183.140000  3.485000  183.310000 3.655000 ;
      RECT  183.225000 -0.085000  183.395000 0.085000 ;
      RECT  183.225000  2.635000  183.395000 2.805000 ;
      RECT  183.225000  5.355000  183.395000 5.525000 ;
      RECT  183.685000 -0.085000  183.855000 0.085000 ;
      RECT  183.685000  2.635000  183.855000 2.805000 ;
      RECT  183.685000  5.355000  183.855000 5.525000 ;
      RECT  184.145000 -0.085000  184.315000 0.085000 ;
      RECT  184.145000  2.635000  184.315000 2.805000 ;
      RECT  184.145000  5.355000  184.315000 5.525000 ;
      RECT  184.605000 -0.085000  184.775000 0.085000 ;
      RECT  184.605000  2.635000  184.775000 2.805000 ;
      RECT  184.605000  5.355000  184.775000 5.525000 ;
      RECT  185.065000 -0.085000  185.235000 0.085000 ;
      RECT  185.065000  2.635000  185.235000 2.805000 ;
      RECT  185.065000  5.355000  185.235000 5.525000 ;
      RECT  185.525000 -0.085000  185.695000 0.085000 ;
      RECT  185.525000  2.635000  185.695000 2.805000 ;
      RECT  185.525000  5.355000  185.695000 5.525000 ;
      RECT  185.985000 -0.085000  186.155000 0.085000 ;
      RECT  185.985000  2.635000  186.155000 2.805000 ;
      RECT  185.985000  5.355000  186.155000 5.525000 ;
      RECT  186.445000 -0.085000  186.615000 0.085000 ;
      RECT  186.445000  2.635000  186.615000 2.805000 ;
      RECT  186.445000  5.355000  186.615000 5.525000 ;
      RECT  186.905000 -0.085000  187.075000 0.085000 ;
      RECT  186.905000  2.635000  187.075000 2.805000 ;
      RECT  186.905000  5.355000  187.075000 5.525000 ;
      RECT  187.365000 -0.085000  187.535000 0.085000 ;
      RECT  187.365000  2.635000  187.535000 2.805000 ;
      RECT  187.365000  3.825000  187.535000 3.995000 ;
      RECT  187.365000  5.355000  187.535000 5.525000 ;
      RECT  187.825000 -0.085000  187.995000 0.085000 ;
      RECT  187.825000  2.635000  187.995000 2.805000 ;
      RECT  187.825000  5.355000  187.995000 5.525000 ;
      RECT  187.875000  3.485000  188.045000 3.655000 ;
      RECT  188.285000 -0.085000  188.455000 0.085000 ;
      RECT  188.285000  2.635000  188.455000 2.805000 ;
      RECT  188.285000  5.355000  188.455000 5.525000 ;
      RECT  188.745000 -0.085000  188.915000 0.085000 ;
      RECT  188.745000  2.635000  188.915000 2.805000 ;
      RECT  188.745000  5.355000  188.915000 5.525000 ;
      RECT  189.205000 -0.085000  189.375000 0.085000 ;
      RECT  189.205000  2.635000  189.375000 2.805000 ;
      RECT  189.205000  5.355000  189.375000 5.525000 ;
      RECT  189.485000  3.825000  189.655000 3.995000 ;
      RECT  189.665000 -0.085000  189.835000 0.085000 ;
      RECT  189.665000  2.635000  189.835000 2.805000 ;
      RECT  189.665000  5.355000  189.835000 5.525000 ;
      RECT  190.040000  3.485000  190.210000 3.655000 ;
      RECT  190.125000 -0.085000  190.295000 0.085000 ;
      RECT  190.125000  2.635000  190.295000 2.805000 ;
      RECT  190.125000  5.355000  190.295000 5.525000 ;
      RECT  190.585000 -0.085000  190.755000 0.085000 ;
      RECT  190.585000  2.635000  190.755000 2.805000 ;
      RECT  190.585000  5.355000  190.755000 5.525000 ;
      RECT  191.045000 -0.085000  191.215000 0.085000 ;
      RECT  191.045000  2.635000  191.215000 2.805000 ;
      RECT  191.045000  5.355000  191.215000 5.525000 ;
      RECT  191.505000 -0.085000  191.675000 0.085000 ;
      RECT  191.505000  2.635000  191.675000 2.805000 ;
      RECT  191.505000  5.355000  191.675000 5.525000 ;
      RECT  191.965000 -0.085000  192.135000 0.085000 ;
      RECT  191.965000  2.635000  192.135000 2.805000 ;
      RECT  191.965000  5.355000  192.135000 5.525000 ;
      RECT  192.425000 -0.085000  192.595000 0.085000 ;
      RECT  192.425000  2.635000  192.595000 2.805000 ;
      RECT  192.425000  5.355000  192.595000 5.525000 ;
      RECT  192.885000 -0.085000  193.055000 0.085000 ;
      RECT  192.885000  2.635000  193.055000 2.805000 ;
      RECT  192.885000  5.355000  193.055000 5.525000 ;
      RECT  193.345000 -0.085000  193.515000 0.085000 ;
      RECT  193.345000  2.635000  193.515000 2.805000 ;
      RECT  193.345000  5.355000  193.515000 5.525000 ;
      RECT  193.805000 -0.085000  193.975000 0.085000 ;
      RECT  193.805000  2.635000  193.975000 2.805000 ;
      RECT  193.805000  5.355000  193.975000 5.525000 ;
      RECT  194.265000 -0.085000  194.435000 0.085000 ;
      RECT  194.265000  2.635000  194.435000 2.805000 ;
      RECT  194.265000  5.355000  194.435000 5.525000 ;
      RECT  194.295000  3.485000  194.465000 3.655000 ;
      RECT  194.725000 -0.085000  194.895000 0.085000 ;
      RECT  194.725000  2.635000  194.895000 2.805000 ;
      RECT  194.725000  5.355000  194.895000 5.525000 ;
      RECT  194.755000  3.825000  194.925000 3.995000 ;
      RECT  195.185000 -0.085000  195.355000 0.085000 ;
      RECT  195.185000  2.635000  195.355000 2.805000 ;
      RECT  195.185000  5.355000  195.355000 5.525000 ;
      RECT  195.645000 -0.085000  195.815000 0.085000 ;
      RECT  195.645000  2.635000  195.815000 2.805000 ;
      RECT  195.645000  5.355000  195.815000 5.525000 ;
      RECT  196.105000 -0.085000  196.275000 0.085000 ;
      RECT  196.105000  2.635000  196.275000 2.805000 ;
      RECT  196.105000  5.355000  196.275000 5.525000 ;
      RECT  196.385000  3.825000  196.555000 3.995000 ;
      RECT  196.565000 -0.085000  196.735000 0.085000 ;
      RECT  196.565000  2.635000  196.735000 2.805000 ;
      RECT  196.565000  5.355000  196.735000 5.525000 ;
      RECT  196.940000  3.485000  197.110000 3.655000 ;
      RECT  197.025000 -0.085000  197.195000 0.085000 ;
      RECT  197.025000  2.635000  197.195000 2.805000 ;
      RECT  197.025000  5.355000  197.195000 5.525000 ;
      RECT  197.485000 -0.085000  197.655000 0.085000 ;
      RECT  197.485000  2.635000  197.655000 2.805000 ;
      RECT  197.485000  5.355000  197.655000 5.525000 ;
      RECT  197.945000 -0.085000  198.115000 0.085000 ;
      RECT  197.945000  2.635000  198.115000 2.805000 ;
      RECT  197.945000  5.355000  198.115000 5.525000 ;
      RECT  198.405000 -0.085000  198.575000 0.085000 ;
      RECT  198.405000  2.635000  198.575000 2.805000 ;
      RECT  198.405000  5.355000  198.575000 5.525000 ;
      RECT  198.865000 -0.085000  199.035000 0.085000 ;
      RECT  198.865000  2.635000  199.035000 2.805000 ;
      RECT  198.865000  5.355000  199.035000 5.525000 ;
      RECT  199.325000 -0.085000  199.495000 0.085000 ;
      RECT  199.325000  2.635000  199.495000 2.805000 ;
      RECT  199.325000  5.355000  199.495000 5.525000 ;
      RECT  199.785000 -0.085000  199.955000 0.085000 ;
      RECT  199.785000  2.635000  199.955000 2.805000 ;
      RECT  199.785000  5.355000  199.955000 5.525000 ;
      RECT  200.245000 -0.085000  200.415000 0.085000 ;
      RECT  200.245000  2.635000  200.415000 2.805000 ;
      RECT  200.245000  5.355000  200.415000 5.525000 ;
      RECT  200.705000 -0.085000  200.875000 0.085000 ;
      RECT  200.705000  2.635000  200.875000 2.805000 ;
      RECT  200.705000  5.355000  200.875000 5.525000 ;
      RECT  201.165000 -0.085000  201.335000 0.085000 ;
      RECT  201.165000  2.635000  201.335000 2.805000 ;
      RECT  201.165000  5.355000  201.335000 5.525000 ;
      RECT  201.625000 -0.085000  201.795000 0.085000 ;
      RECT  201.625000  2.635000  201.795000 2.805000 ;
      RECT  201.625000  3.825000  201.795000 3.995000 ;
      RECT  201.625000  5.355000  201.795000 5.525000 ;
      RECT  202.085000 -0.085000  202.255000 0.085000 ;
      RECT  202.085000  2.635000  202.255000 2.805000 ;
      RECT  202.085000  5.355000  202.255000 5.525000 ;
      RECT  202.135000  3.485000  202.305000 3.655000 ;
      RECT  202.545000 -0.085000  202.715000 0.085000 ;
      RECT  202.545000  2.635000  202.715000 2.805000 ;
      RECT  202.545000  5.355000  202.715000 5.525000 ;
      RECT  203.005000 -0.085000  203.175000 0.085000 ;
      RECT  203.005000  2.635000  203.175000 2.805000 ;
      RECT  203.005000  5.355000  203.175000 5.525000 ;
      RECT  203.465000 -0.085000  203.635000 0.085000 ;
      RECT  203.465000  2.635000  203.635000 2.805000 ;
      RECT  203.465000  5.355000  203.635000 5.525000 ;
      RECT  203.745000  3.825000  203.915000 3.995000 ;
      RECT  203.925000 -0.085000  204.095000 0.085000 ;
      RECT  203.925000  2.635000  204.095000 2.805000 ;
      RECT  203.925000  5.355000  204.095000 5.525000 ;
      RECT  204.300000  3.485000  204.470000 3.655000 ;
      RECT  204.385000 -0.085000  204.555000 0.085000 ;
      RECT  204.385000  2.635000  204.555000 2.805000 ;
      RECT  204.385000  5.355000  204.555000 5.525000 ;
      RECT  204.845000 -0.085000  205.015000 0.085000 ;
      RECT  204.845000  2.635000  205.015000 2.805000 ;
      RECT  204.845000  5.355000  205.015000 5.525000 ;
      RECT  205.305000 -0.085000  205.475000 0.085000 ;
      RECT  205.305000  2.635000  205.475000 2.805000 ;
      RECT  205.305000  5.355000  205.475000 5.525000 ;
      RECT  205.765000 -0.085000  205.935000 0.085000 ;
      RECT  205.765000  2.635000  205.935000 2.805000 ;
      RECT  205.765000  5.355000  205.935000 5.525000 ;
      RECT  206.225000 -0.085000  206.395000 0.085000 ;
      RECT  206.225000  2.635000  206.395000 2.805000 ;
      RECT  206.225000  5.355000  206.395000 5.525000 ;
      RECT  206.685000 -0.085000  206.855000 0.085000 ;
      RECT  206.685000  2.635000  206.855000 2.805000 ;
      RECT  206.685000  5.355000  206.855000 5.525000 ;
      RECT  207.145000 -0.085000  207.315000 0.085000 ;
      RECT  207.145000  2.635000  207.315000 2.805000 ;
      RECT  207.145000  5.355000  207.315000 5.525000 ;
      RECT  207.605000 -0.085000  207.775000 0.085000 ;
      RECT  207.605000  2.635000  207.775000 2.805000 ;
      RECT  207.605000  5.355000  207.775000 5.525000 ;
      RECT  208.065000 -0.085000  208.235000 0.085000 ;
      RECT  208.065000  2.635000  208.235000 2.805000 ;
      RECT  208.065000  5.355000  208.235000 5.525000 ;
      RECT  208.525000 -0.085000  208.695000 0.085000 ;
      RECT  208.525000  2.635000  208.695000 2.805000 ;
      RECT  208.525000  5.355000  208.695000 5.525000 ;
      RECT  208.985000 -0.085000  209.155000 0.085000 ;
      RECT  208.985000  2.635000  209.155000 2.805000 ;
      RECT  208.985000  5.355000  209.155000 5.525000 ;
      RECT  209.015000  3.485000  209.185000 3.655000 ;
      RECT  209.445000 -0.085000  209.615000 0.085000 ;
      RECT  209.445000  2.635000  209.615000 2.805000 ;
      RECT  209.445000  5.355000  209.615000 5.525000 ;
      RECT  209.475000  3.825000  209.645000 3.995000 ;
      RECT  209.905000 -0.085000  210.075000 0.085000 ;
      RECT  209.905000  2.635000  210.075000 2.805000 ;
      RECT  209.905000  5.355000  210.075000 5.525000 ;
      RECT  210.365000 -0.085000  210.535000 0.085000 ;
      RECT  210.365000  2.635000  210.535000 2.805000 ;
      RECT  210.365000  5.355000  210.535000 5.525000 ;
      RECT  210.825000 -0.085000  210.995000 0.085000 ;
      RECT  210.825000  2.635000  210.995000 2.805000 ;
      RECT  210.825000  5.355000  210.995000 5.525000 ;
      RECT  211.105000  3.825000  211.275000 3.995000 ;
      RECT  211.285000 -0.085000  211.455000 0.085000 ;
      RECT  211.285000  2.635000  211.455000 2.805000 ;
      RECT  211.285000  5.355000  211.455000 5.525000 ;
      RECT  211.660000  3.485000  211.830000 3.655000 ;
      RECT  211.745000 -0.085000  211.915000 0.085000 ;
      RECT  211.745000  2.635000  211.915000 2.805000 ;
      RECT  211.745000  5.355000  211.915000 5.525000 ;
      RECT  212.205000 -0.085000  212.375000 0.085000 ;
      RECT  212.205000  2.635000  212.375000 2.805000 ;
      RECT  212.205000  5.355000  212.375000 5.525000 ;
      RECT  212.665000 -0.085000  212.835000 0.085000 ;
      RECT  212.665000  2.635000  212.835000 2.805000 ;
      RECT  212.665000  5.355000  212.835000 5.525000 ;
      RECT  213.125000 -0.085000  213.295000 0.085000 ;
      RECT  213.125000  2.635000  213.295000 2.805000 ;
      RECT  213.125000  5.355000  213.295000 5.525000 ;
      RECT  213.585000 -0.085000  213.755000 0.085000 ;
      RECT  213.585000  2.635000  213.755000 2.805000 ;
      RECT  213.585000  5.355000  213.755000 5.525000 ;
      RECT  214.045000 -0.085000  214.215000 0.085000 ;
      RECT  214.045000  2.635000  214.215000 2.805000 ;
      RECT  214.045000  5.355000  214.215000 5.525000 ;
      RECT  214.505000 -0.085000  214.675000 0.085000 ;
      RECT  214.505000  2.635000  214.675000 2.805000 ;
      RECT  214.505000  5.355000  214.675000 5.525000 ;
      RECT  214.965000 -0.085000  215.135000 0.085000 ;
      RECT  214.965000  2.635000  215.135000 2.805000 ;
      RECT  214.965000  5.355000  215.135000 5.525000 ;
      RECT  215.425000 -0.085000  215.595000 0.085000 ;
      RECT  215.425000  2.635000  215.595000 2.805000 ;
      RECT  215.425000  5.355000  215.595000 5.525000 ;
      RECT  215.885000 -0.085000  216.055000 0.085000 ;
      RECT  215.885000  2.635000  216.055000 2.805000 ;
      RECT  215.885000  5.355000  216.055000 5.525000 ;
      RECT  216.345000 -0.085000  216.515000 0.085000 ;
      RECT  216.345000  2.635000  216.515000 2.805000 ;
      RECT  216.345000  5.355000  216.515000 5.525000 ;
      RECT  216.805000 -0.085000  216.975000 0.085000 ;
      RECT  216.805000  2.635000  216.975000 2.805000 ;
      RECT  216.805000  5.355000  216.975000 5.525000 ;
      RECT  217.265000 -0.085000  217.435000 0.085000 ;
      RECT  217.265000  2.635000  217.435000 2.805000 ;
      RECT  217.265000  3.825000  217.435000 3.995000 ;
      RECT  217.265000  5.355000  217.435000 5.525000 ;
      RECT  217.725000 -0.085000  217.895000 0.085000 ;
      RECT  217.725000  2.635000  217.895000 2.805000 ;
      RECT  217.725000  5.355000  217.895000 5.525000 ;
      RECT  217.775000  3.485000  217.945000 3.655000 ;
      RECT  218.185000 -0.085000  218.355000 0.085000 ;
      RECT  218.185000  2.635000  218.355000 2.805000 ;
      RECT  218.185000  5.355000  218.355000 5.525000 ;
      RECT  218.645000 -0.085000  218.815000 0.085000 ;
      RECT  218.645000  2.635000  218.815000 2.805000 ;
      RECT  218.645000  5.355000  218.815000 5.525000 ;
      RECT  219.105000 -0.085000  219.275000 0.085000 ;
      RECT  219.105000  2.635000  219.275000 2.805000 ;
      RECT  219.105000  5.355000  219.275000 5.525000 ;
      RECT  219.385000  3.825000  219.555000 3.995000 ;
      RECT  219.565000 -0.085000  219.735000 0.085000 ;
      RECT  219.565000  2.635000  219.735000 2.805000 ;
      RECT  219.565000  5.355000  219.735000 5.525000 ;
      RECT  219.940000  3.485000  220.110000 3.655000 ;
      RECT  220.025000 -0.085000  220.195000 0.085000 ;
      RECT  220.025000  2.635000  220.195000 2.805000 ;
      RECT  220.025000  5.355000  220.195000 5.525000 ;
      RECT  220.485000 -0.085000  220.655000 0.085000 ;
      RECT  220.485000  2.635000  220.655000 2.805000 ;
      RECT  220.485000  5.355000  220.655000 5.525000 ;
      RECT  220.945000 -0.085000  221.115000 0.085000 ;
      RECT  220.945000  2.635000  221.115000 2.805000 ;
      RECT  220.945000  5.355000  221.115000 5.525000 ;
      RECT  221.405000 -0.085000  221.575000 0.085000 ;
      RECT  221.405000  2.635000  221.575000 2.805000 ;
      RECT  221.405000  5.355000  221.575000 5.525000 ;
      RECT  221.865000 -0.085000  222.035000 0.085000 ;
      RECT  221.865000  2.635000  222.035000 2.805000 ;
      RECT  221.865000  5.355000  222.035000 5.525000 ;
      RECT  222.325000 -0.085000  222.495000 0.085000 ;
      RECT  222.325000  2.635000  222.495000 2.805000 ;
      RECT  222.325000  5.355000  222.495000 5.525000 ;
      RECT  222.785000 -0.085000  222.955000 0.085000 ;
      RECT  222.785000  2.635000  222.955000 2.805000 ;
      RECT  222.785000  5.355000  222.955000 5.525000 ;
      RECT  223.245000 -0.085000  223.415000 0.085000 ;
      RECT  223.245000  2.635000  223.415000 2.805000 ;
      RECT  223.245000  5.355000  223.415000 5.525000 ;
      RECT  223.705000 -0.085000  223.875000 0.085000 ;
      RECT  223.705000  2.635000  223.875000 2.805000 ;
      RECT  223.705000  5.355000  223.875000 5.525000 ;
      RECT  224.165000 -0.085000  224.335000 0.085000 ;
      RECT  224.165000  2.635000  224.335000 2.805000 ;
      RECT  224.165000  5.355000  224.335000 5.525000 ;
      RECT  224.625000 -0.085000  224.795000 0.085000 ;
      RECT  224.625000  2.635000  224.795000 2.805000 ;
      RECT  224.625000  5.355000  224.795000 5.525000 ;
      RECT  225.085000 -0.085000  225.255000 0.085000 ;
      RECT  225.085000  2.635000  225.255000 2.805000 ;
      RECT  225.085000  5.355000  225.255000 5.525000 ;
      RECT  225.545000 -0.085000  225.715000 0.085000 ;
      RECT  225.545000  2.635000  225.715000 2.805000 ;
      RECT  225.545000  5.355000  225.715000 5.525000 ;
      RECT  226.005000 -0.085000  226.175000 0.085000 ;
      RECT  226.005000  2.635000  226.175000 2.805000 ;
      RECT  226.005000  5.355000  226.175000 5.525000 ;
      RECT  226.465000 -0.085000  226.635000 0.085000 ;
      RECT  226.465000  2.635000  226.635000 2.805000 ;
      RECT  226.465000  5.355000  226.635000 5.525000 ;
      RECT  226.925000 -0.085000  227.095000 0.085000 ;
      RECT  226.925000  2.635000  227.095000 2.805000 ;
      RECT  226.925000  5.355000  227.095000 5.525000 ;
      RECT  227.385000 -0.085000  227.555000 0.085000 ;
      RECT  227.385000  2.635000  227.555000 2.805000 ;
      RECT  227.385000  5.355000  227.555000 5.525000 ;
      RECT  227.845000 -0.085000  228.015000 0.085000 ;
      RECT  227.845000  2.635000  228.015000 2.805000 ;
      RECT  227.845000  5.355000  228.015000 5.525000 ;
      RECT  228.305000 -0.085000  228.475000 0.085000 ;
      RECT  228.305000  2.635000  228.475000 2.805000 ;
      RECT  228.305000  5.355000  228.475000 5.525000 ;
      RECT  228.765000 -0.085000  228.935000 0.085000 ;
      RECT  228.765000  2.635000  228.935000 2.805000 ;
      RECT  228.765000  5.355000  228.935000 5.525000 ;
      RECT  229.225000 -0.085000  229.395000 0.085000 ;
      RECT  229.225000  2.635000  229.395000 2.805000 ;
      RECT  229.225000  5.355000  229.395000 5.525000 ;
      RECT  229.685000 -0.085000  229.855000 0.085000 ;
      RECT  229.685000  2.635000  229.855000 2.805000 ;
      RECT  229.685000  5.355000  229.855000 5.525000 ;
      RECT  230.145000 -0.085000  230.315000 0.085000 ;
      RECT  230.145000  2.635000  230.315000 2.805000 ;
      RECT  230.145000  5.355000  230.315000 5.525000 ;
      RECT  230.605000 -0.085000  230.775000 0.085000 ;
      RECT  230.605000  2.635000  230.775000 2.805000 ;
      RECT  230.605000  5.355000  230.775000 5.525000 ;
      RECT  231.065000 -0.085000  231.235000 0.085000 ;
      RECT  231.065000  2.635000  231.235000 2.805000 ;
      RECT  231.065000  5.355000  231.235000 5.525000 ;
      RECT  231.525000 -0.085000  231.695000 0.085000 ;
      RECT  231.525000  2.635000  231.695000 2.805000 ;
      RECT  231.525000  5.355000  231.695000 5.525000 ;
      RECT  231.985000 -0.085000  232.155000 0.085000 ;
      RECT  231.985000  2.635000  232.155000 2.805000 ;
      RECT  231.985000  5.355000  232.155000 5.525000 ;
      RECT  232.445000 -0.085000  232.615000 0.085000 ;
      RECT  232.445000  2.635000  232.615000 2.805000 ;
      RECT  232.445000  5.355000  232.615000 5.525000 ;
      RECT  232.905000 -0.085000  233.075000 0.085000 ;
      RECT  232.905000  2.635000  233.075000 2.805000 ;
      RECT  232.905000  5.355000  233.075000 5.525000 ;
      RECT  233.365000 -0.085000  233.535000 0.085000 ;
      RECT  233.365000  2.635000  233.535000 2.805000 ;
      RECT  233.365000  5.355000  233.535000 5.525000 ;
      RECT  233.825000 -0.085000  233.995000 0.085000 ;
      RECT  233.825000  2.635000  233.995000 2.805000 ;
      RECT  233.825000  5.355000  233.995000 5.525000 ;
      RECT  234.285000 -0.085000  234.455000 0.085000 ;
      RECT  234.285000  2.635000  234.455000 2.805000 ;
      RECT  234.285000  5.355000  234.455000 5.525000 ;
      RECT  234.745000 -0.085000  234.915000 0.085000 ;
      RECT  234.745000  2.635000  234.915000 2.805000 ;
      RECT  235.205000 -0.085000  235.375000 0.085000 ;
      RECT  235.205000  2.635000  235.375000 2.805000 ;
      RECT  235.665000 -0.085000  235.835000 0.085000 ;
      RECT  235.665000  2.635000  235.835000 2.805000 ;
      RECT  236.125000 -0.085000  236.295000 0.085000 ;
      RECT  236.125000  2.635000  236.295000 2.805000 ;
      RECT  236.585000 -0.085000  236.755000 0.085000 ;
      RECT  236.585000  2.635000  236.755000 2.805000 ;
      RECT  237.045000 -0.085000  237.215000 0.085000 ;
      RECT  237.045000  2.635000  237.215000 2.805000 ;
      RECT  237.505000 -0.085000  237.675000 0.085000 ;
      RECT  237.505000  2.635000  237.675000 2.805000 ;
      RECT  237.965000 -0.085000  238.135000 0.085000 ;
      RECT  237.965000  2.635000  238.135000 2.805000 ;
      RECT  238.425000 -0.085000  238.595000 0.085000 ;
      RECT  238.425000  2.635000  238.595000 2.805000 ;
      RECT  238.885000 -0.085000  239.055000 0.085000 ;
      RECT  238.885000  2.635000  239.055000 2.805000 ;
      RECT  239.345000 -0.085000  239.515000 0.085000 ;
      RECT  239.345000  2.635000  239.515000 2.805000 ;
      RECT  239.805000 -0.085000  239.975000 0.085000 ;
      RECT  239.805000  2.635000  239.975000 2.805000 ;
      RECT  240.265000 -0.085000  240.435000 0.085000 ;
      RECT  240.265000  2.635000  240.435000 2.805000 ;
      RECT  240.725000 -0.085000  240.895000 0.085000 ;
      RECT  240.725000  2.635000  240.895000 2.805000 ;
      RECT  241.185000 -0.085000  241.355000 0.085000 ;
      RECT  241.185000  2.635000  241.355000 2.805000 ;
      RECT  241.645000 -0.085000  241.815000 0.085000 ;
      RECT  241.645000  2.635000  241.815000 2.805000 ;
      RECT  242.105000 -0.085000  242.275000 0.085000 ;
      RECT  242.105000  2.635000  242.275000 2.805000 ;
      RECT  242.565000 -0.085000  242.735000 0.085000 ;
      RECT  242.565000  2.635000  242.735000 2.805000 ;
      RECT  243.025000 -0.085000  243.195000 0.085000 ;
      RECT  243.025000  2.635000  243.195000 2.805000 ;
      RECT  243.485000 -0.085000  243.655000 0.085000 ;
      RECT  243.485000  2.635000  243.655000 2.805000 ;
      RECT  243.945000 -0.085000  244.115000 0.085000 ;
      RECT  243.945000  2.635000  244.115000 2.805000 ;
      RECT  244.405000 -0.085000  244.575000 0.085000 ;
      RECT  244.405000  2.635000  244.575000 2.805000 ;
      RECT  244.865000 -0.085000  245.035000 0.085000 ;
      RECT  244.865000  2.635000  245.035000 2.805000 ;
      RECT  245.325000 -0.085000  245.495000 0.085000 ;
      RECT  245.325000  2.635000  245.495000 2.805000 ;
      RECT  245.785000 -0.085000  245.955000 0.085000 ;
      RECT  245.785000  2.635000  245.955000 2.805000 ;
      RECT  246.245000 -0.085000  246.415000 0.085000 ;
      RECT  246.245000  2.635000  246.415000 2.805000 ;
      RECT  246.705000 -0.085000  246.875000 0.085000 ;
      RECT  246.705000  2.635000  246.875000 2.805000 ;
      RECT  247.165000 -0.085000  247.335000 0.085000 ;
      RECT  247.165000  2.635000  247.335000 2.805000 ;
      RECT  247.625000 -0.085000  247.795000 0.085000 ;
      RECT  247.625000  2.635000  247.795000 2.805000 ;
      RECT  248.085000 -0.085000  248.255000 0.085000 ;
      RECT  248.085000  2.635000  248.255000 2.805000 ;
      RECT  248.545000 -0.085000  248.715000 0.085000 ;
      RECT  248.545000  2.635000  248.715000 2.805000 ;
      RECT  249.005000 -0.085000  249.175000 0.085000 ;
      RECT  249.005000  2.635000  249.175000 2.805000 ;
      RECT  249.465000 -0.085000  249.635000 0.085000 ;
      RECT  249.465000  2.635000  249.635000 2.805000 ;
      RECT  249.925000 -0.085000  250.095000 0.085000 ;
      RECT  249.925000  2.635000  250.095000 2.805000 ;
      RECT  250.385000 -0.085000  250.555000 0.085000 ;
      RECT  250.385000  2.635000  250.555000 2.805000 ;
      RECT  250.845000 -0.085000  251.015000 0.085000 ;
      RECT  250.845000  2.635000  251.015000 2.805000 ;
      RECT  251.305000 -0.085000  251.475000 0.085000 ;
      RECT  251.305000  2.635000  251.475000 2.805000 ;
      RECT  251.765000 -0.085000  251.935000 0.085000 ;
      RECT  251.765000  2.635000  251.935000 2.805000 ;
      RECT  252.225000 -0.085000  252.395000 0.085000 ;
      RECT  252.225000  2.635000  252.395000 2.805000 ;
      RECT  252.685000 -0.085000  252.855000 0.085000 ;
      RECT  252.685000  2.635000  252.855000 2.805000 ;
      RECT  253.145000 -0.085000  253.315000 0.085000 ;
      RECT  253.145000  2.635000  253.315000 2.805000 ;
      RECT  253.605000 -0.085000  253.775000 0.085000 ;
      RECT  253.605000  2.635000  253.775000 2.805000 ;
      RECT  254.065000 -0.085000  254.235000 0.085000 ;
      RECT  254.065000  2.635000  254.235000 2.805000 ;
      RECT  254.525000 -0.085000  254.695000 0.085000 ;
      RECT  254.525000  2.635000  254.695000 2.805000 ;
      RECT  254.985000 -0.085000  255.155000 0.085000 ;
      RECT  254.985000  2.635000  255.155000 2.805000 ;
      RECT  255.445000 -0.085000  255.615000 0.085000 ;
      RECT  255.445000  2.635000  255.615000 2.805000 ;
      RECT  255.905000 -0.085000  256.075000 0.085000 ;
      RECT  255.905000  2.635000  256.075000 2.805000 ;
      RECT  256.365000 -0.085000  256.535000 0.085000 ;
      RECT  256.365000  2.635000  256.535000 2.805000 ;
      RECT  256.825000 -0.085000  256.995000 0.085000 ;
      RECT  256.825000  2.635000  256.995000 2.805000 ;
      RECT  257.285000 -0.085000  257.455000 0.085000 ;
      RECT  257.285000  2.635000  257.455000 2.805000 ;
      RECT  257.745000 -0.085000  257.915000 0.085000 ;
      RECT  257.745000  2.635000  257.915000 2.805000 ;
      RECT  258.205000 -0.085000  258.375000 0.085000 ;
      RECT  258.205000  2.635000  258.375000 2.805000 ;
      RECT  258.665000 -0.085000  258.835000 0.085000 ;
      RECT  258.665000  2.635000  258.835000 2.805000 ;
      RECT  259.125000 -0.085000  259.295000 0.085000 ;
      RECT  259.125000  2.635000  259.295000 2.805000 ;
      RECT  259.585000 -0.085000  259.755000 0.085000 ;
      RECT  259.585000  2.635000  259.755000 2.805000 ;
      RECT  260.045000 -0.085000  260.215000 0.085000 ;
      RECT  260.045000  2.635000  260.215000 2.805000 ;
      RECT  260.505000 -0.085000  260.675000 0.085000 ;
      RECT  260.505000  2.635000  260.675000 2.805000 ;
      RECT  260.965000 -0.085000  261.135000 0.085000 ;
      RECT  260.965000  2.635000  261.135000 2.805000 ;
      RECT  261.425000 -0.085000  261.595000 0.085000 ;
      RECT  261.425000  2.635000  261.595000 2.805000 ;
      RECT  261.885000 -0.085000  262.055000 0.085000 ;
      RECT  261.885000  2.635000  262.055000 2.805000 ;
      RECT  262.345000 -0.085000  262.515000 0.085000 ;
      RECT  262.345000  2.635000  262.515000 2.805000 ;
      RECT  262.805000 -0.085000  262.975000 0.085000 ;
      RECT  262.805000  2.635000  262.975000 2.805000 ;
      RECT  263.265000 -0.085000  263.435000 0.085000 ;
      RECT  263.265000  2.635000  263.435000 2.805000 ;
      RECT  263.725000 -0.085000  263.895000 0.085000 ;
      RECT  263.725000  2.635000  263.895000 2.805000 ;
      RECT  264.185000 -0.085000  264.355000 0.085000 ;
      RECT  264.185000  2.635000  264.355000 2.805000 ;
      RECT  264.645000 -0.085000  264.815000 0.085000 ;
      RECT  264.645000  2.635000  264.815000 2.805000 ;
      RECT  265.105000 -0.085000  265.275000 0.085000 ;
      RECT  265.105000  2.635000  265.275000 2.805000 ;
      RECT  265.565000 -0.085000  265.735000 0.085000 ;
      RECT  265.565000  2.635000  265.735000 2.805000 ;
      RECT  266.025000 -0.085000  266.195000 0.085000 ;
      RECT  266.025000  2.635000  266.195000 2.805000 ;
      RECT  266.485000 -0.085000  266.655000 0.085000 ;
      RECT  266.485000  2.635000  266.655000 2.805000 ;
      RECT  266.945000 -0.085000  267.115000 0.085000 ;
      RECT  266.945000  2.635000  267.115000 2.805000 ;
      RECT  267.405000 -0.085000  267.575000 0.085000 ;
      RECT  267.405000  2.635000  267.575000 2.805000 ;
      RECT  267.865000 -0.085000  268.035000 0.085000 ;
      RECT  267.865000  2.635000  268.035000 2.805000 ;
      RECT  268.785000 -0.085000  268.955000 0.085000 ;
      RECT  268.785000  2.635000  268.955000 2.805000 ;
      RECT  269.245000 -0.085000  269.415000 0.085000 ;
      RECT  269.245000  2.635000  269.415000 2.805000 ;
      RECT  269.705000 -0.085000  269.875000 0.085000 ;
      RECT  269.705000  2.635000  269.875000 2.805000 ;
      RECT  270.165000 -0.085000  270.335000 0.085000 ;
      RECT  270.165000  2.635000  270.335000 2.805000 ;
      RECT  270.625000 -0.085000  270.795000 0.085000 ;
      RECT  270.625000  2.635000  270.795000 2.805000 ;
      RECT  271.085000 -0.085000  271.255000 0.085000 ;
      RECT  271.085000  2.635000  271.255000 2.805000 ;
      RECT  271.545000 -0.085000  271.715000 0.085000 ;
      RECT  271.545000  2.635000  271.715000 2.805000 ;
      RECT  272.005000 -0.085000  272.175000 0.085000 ;
      RECT  272.005000  2.635000  272.175000 2.805000 ;
      RECT  272.465000 -0.085000  272.635000 0.085000 ;
      RECT  272.465000  2.635000  272.635000 2.805000 ;
      RECT  272.925000 -0.085000  273.095000 0.085000 ;
      RECT  272.925000  2.635000  273.095000 2.805000 ;
      RECT  273.385000 -0.085000  273.555000 0.085000 ;
      RECT  273.385000  2.635000  273.555000 2.805000 ;
      RECT  273.845000 -0.085000  274.015000 0.085000 ;
      RECT  273.845000  2.635000  274.015000 2.805000 ;
      RECT  274.305000 -0.085000  274.475000 0.085000 ;
      RECT  274.305000  2.635000  274.475000 2.805000 ;
      RECT  274.765000 -0.085000  274.935000 0.085000 ;
      RECT  274.765000  2.635000  274.935000 2.805000 ;
      RECT  275.225000 -0.085000  275.395000 0.085000 ;
      RECT  275.225000  2.635000  275.395000 2.805000 ;
      RECT  275.685000 -0.085000  275.855000 0.085000 ;
      RECT  275.685000  2.635000  275.855000 2.805000 ;
      RECT  276.145000 -0.085000  276.315000 0.085000 ;
      RECT  276.145000  2.635000  276.315000 2.805000 ;
      RECT  276.605000 -0.085000  276.775000 0.085000 ;
      RECT  276.605000  2.635000  276.775000 2.805000 ;
      RECT  277.065000 -0.085000  277.235000 0.085000 ;
      RECT  277.065000  2.635000  277.235000 2.805000 ;
      RECT  277.525000 -0.085000  277.695000 0.085000 ;
      RECT  277.525000  2.635000  277.695000 2.805000 ;
      RECT  277.985000 -0.085000  278.155000 0.085000 ;
      RECT  277.985000  2.635000  278.155000 2.805000 ;
      RECT  278.445000 -0.085000  278.615000 0.085000 ;
      RECT  278.445000  2.635000  278.615000 2.805000 ;
      RECT  278.905000 -0.085000  279.075000 0.085000 ;
      RECT  278.905000  2.635000  279.075000 2.805000 ;
      RECT  279.365000 -0.085000  279.535000 0.085000 ;
      RECT  279.365000  2.635000  279.535000 2.805000 ;
      RECT  279.825000 -0.085000  279.995000 0.085000 ;
      RECT  279.825000  2.635000  279.995000 2.805000 ;
      RECT  280.285000 -0.085000  280.455000 0.085000 ;
      RECT  280.285000  2.635000  280.455000 2.805000 ;
      RECT  280.745000 -0.085000  280.915000 0.085000 ;
      RECT  280.745000  2.635000  280.915000 2.805000 ;
      RECT  281.205000 -0.085000  281.375000 0.085000 ;
      RECT  281.205000  2.635000  281.375000 2.805000 ;
      RECT  281.665000 -0.085000  281.835000 0.085000 ;
      RECT  281.665000  2.635000  281.835000 2.805000 ;
      RECT  282.125000 -0.085000  282.295000 0.085000 ;
      RECT  282.125000  2.635000  282.295000 2.805000 ;
      RECT  282.585000 -0.085000  282.755000 0.085000 ;
      RECT  282.585000  2.635000  282.755000 2.805000 ;
      RECT  283.045000 -0.085000  283.215000 0.085000 ;
      RECT  283.045000  2.635000  283.215000 2.805000 ;
      RECT  283.505000 -0.085000  283.675000 0.085000 ;
      RECT  283.505000  2.635000  283.675000 2.805000 ;
      RECT  283.965000 -0.085000  284.135000 0.085000 ;
      RECT  283.965000  2.635000  284.135000 2.805000 ;
      RECT  284.425000 -0.085000  284.595000 0.085000 ;
      RECT  284.425000  2.635000  284.595000 2.805000 ;
      RECT  284.885000 -0.085000  285.055000 0.085000 ;
      RECT  284.885000  2.635000  285.055000 2.805000 ;
      RECT  285.345000 -0.085000  285.515000 0.085000 ;
      RECT  285.345000  2.635000  285.515000 2.805000 ;
      RECT  285.805000 -0.085000  285.975000 0.085000 ;
      RECT  285.805000  2.635000  285.975000 2.805000 ;
      RECT  286.265000 -0.085000  286.435000 0.085000 ;
      RECT  286.265000  2.635000  286.435000 2.805000 ;
      RECT  286.725000 -0.085000  286.895000 0.085000 ;
      RECT  286.725000  2.635000  286.895000 2.805000 ;
      RECT  287.185000 -0.085000  287.355000 0.085000 ;
      RECT  287.185000  2.635000  287.355000 2.805000 ;
      RECT  287.645000 -0.085000  287.815000 0.085000 ;
      RECT  287.645000  2.635000  287.815000 2.805000 ;
      RECT  288.105000 -0.085000  288.275000 0.085000 ;
      RECT  288.105000  2.635000  288.275000 2.805000 ;
      RECT  288.565000 -0.085000  288.735000 0.085000 ;
      RECT  288.565000  2.635000  288.735000 2.805000 ;
      RECT  289.025000 -0.085000  289.195000 0.085000 ;
      RECT  289.025000  2.635000  289.195000 2.805000 ;
      RECT  289.485000 -0.085000  289.655000 0.085000 ;
      RECT  289.485000  2.635000  289.655000 2.805000 ;
      RECT  289.945000 -0.085000  290.115000 0.085000 ;
      RECT  289.945000  2.635000  290.115000 2.805000 ;
      RECT  290.405000 -0.085000  290.575000 0.085000 ;
      RECT  290.405000  2.635000  290.575000 2.805000 ;
      RECT  290.865000 -0.085000  291.035000 0.085000 ;
      RECT  290.865000  2.635000  291.035000 2.805000 ;
      RECT  291.325000 -0.085000  291.495000 0.085000 ;
      RECT  291.325000  2.635000  291.495000 2.805000 ;
      RECT  291.785000 -0.085000  291.955000 0.085000 ;
      RECT  291.785000  2.635000  291.955000 2.805000 ;
      RECT  292.245000 -0.085000  292.415000 0.085000 ;
      RECT  292.245000  2.635000  292.415000 2.805000 ;
      RECT  292.705000 -0.085000  292.875000 0.085000 ;
      RECT  292.705000  2.635000  292.875000 2.805000 ;
      RECT  293.165000 -0.085000  293.335000 0.085000 ;
      RECT  293.165000  2.635000  293.335000 2.805000 ;
      RECT  293.625000 -0.085000  293.795000 0.085000 ;
      RECT  293.625000  2.635000  293.795000 2.805000 ;
      RECT  294.085000 -0.085000  294.255000 0.085000 ;
      RECT  294.085000  2.635000  294.255000 2.805000 ;
      RECT  294.545000 -0.085000  294.715000 0.085000 ;
      RECT  294.545000  2.635000  294.715000 2.805000 ;
      RECT  295.005000 -0.085000  295.175000 0.085000 ;
      RECT  295.005000  2.635000  295.175000 2.805000 ;
      RECT  295.465000 -0.085000  295.635000 0.085000 ;
      RECT  295.465000  2.635000  295.635000 2.805000 ;
      RECT  295.925000 -0.085000  296.095000 0.085000 ;
      RECT  295.925000  2.635000  296.095000 2.805000 ;
      RECT  296.385000 -0.085000  296.555000 0.085000 ;
      RECT  296.385000  2.635000  296.555000 2.805000 ;
      RECT  296.845000 -0.085000  297.015000 0.085000 ;
      RECT  296.845000  2.635000  297.015000 2.805000 ;
      RECT  297.305000 -0.085000  297.475000 0.085000 ;
      RECT  297.305000  2.635000  297.475000 2.805000 ;
      RECT  297.765000 -0.085000  297.935000 0.085000 ;
      RECT  297.765000  2.635000  297.935000 2.805000 ;
      RECT  298.225000 -0.085000  298.395000 0.085000 ;
      RECT  298.225000  2.635000  298.395000 2.805000 ;
      RECT  298.685000 -0.085000  298.855000 0.085000 ;
      RECT  298.685000  2.635000  298.855000 2.805000 ;
      RECT  299.145000 -0.085000  299.315000 0.085000 ;
      RECT  299.145000  2.635000  299.315000 2.805000 ;
      RECT  299.605000 -0.085000  299.775000 0.085000 ;
      RECT  299.605000  2.635000  299.775000 2.805000 ;
      RECT  300.065000 -0.085000  300.235000 0.085000 ;
      RECT  300.065000  2.635000  300.235000 2.805000 ;
      RECT  300.525000 -0.085000  300.695000 0.085000 ;
      RECT  300.525000  2.635000  300.695000 2.805000 ;
      RECT  300.985000 -0.085000  301.155000 0.085000 ;
      RECT  300.985000  2.635000  301.155000 2.805000 ;
      RECT  301.445000 -0.085000  301.615000 0.085000 ;
      RECT  301.445000  2.635000  301.615000 2.805000 ;
      RECT  301.905000 -0.085000  302.075000 0.085000 ;
      RECT  301.905000  2.635000  302.075000 2.805000 ;
      RECT  302.365000 -0.085000  302.535000 0.085000 ;
      RECT  302.365000  2.635000  302.535000 2.805000 ;
      RECT  302.825000 -0.085000  302.995000 0.085000 ;
      RECT  302.825000  2.635000  302.995000 2.805000 ;
      RECT  303.285000 -0.085000  303.455000 0.085000 ;
      RECT  303.285000  2.635000  303.455000 2.805000 ;
      RECT  303.745000 -0.085000  303.915000 0.085000 ;
      RECT  303.745000  2.635000  303.915000 2.805000 ;
      RECT  304.205000 -0.085000  304.375000 0.085000 ;
      RECT  304.205000  2.635000  304.375000 2.805000 ;
      RECT  304.665000 -0.085000  304.835000 0.085000 ;
      RECT  304.665000  2.635000  304.835000 2.805000 ;
      RECT  305.125000 -0.085000  305.295000 0.085000 ;
      RECT  305.125000  2.635000  305.295000 2.805000 ;
      RECT  305.585000 -0.085000  305.755000 0.085000 ;
      RECT  305.585000  2.635000  305.755000 2.805000 ;
      RECT  306.045000 -0.085000  306.215000 0.085000 ;
      RECT  306.045000  2.635000  306.215000 2.805000 ;
      RECT  306.505000 -0.085000  306.675000 0.085000 ;
      RECT  306.505000  2.635000  306.675000 2.805000 ;
      RECT  306.965000 -0.085000  307.135000 0.085000 ;
      RECT  306.965000  2.635000  307.135000 2.805000 ;
      RECT  307.425000 -0.085000  307.595000 0.085000 ;
      RECT  307.425000  2.635000  307.595000 2.805000 ;
      RECT  307.885000 -0.085000  308.055000 0.085000 ;
      RECT  307.885000  2.635000  308.055000 2.805000 ;
      RECT  308.345000 -0.085000  308.515000 0.085000 ;
      RECT  308.345000  2.635000  308.515000 2.805000 ;
      RECT  308.805000 -0.085000  308.975000 0.085000 ;
      RECT  308.805000  2.635000  308.975000 2.805000 ;
      RECT  309.265000 -0.085000  309.435000 0.085000 ;
      RECT  309.265000  2.635000  309.435000 2.805000 ;
      RECT  309.725000 -0.085000  309.895000 0.085000 ;
      RECT  309.725000  2.635000  309.895000 2.805000 ;
      RECT  310.185000 -0.085000  310.355000 0.085000 ;
      RECT  310.185000  2.635000  310.355000 2.805000 ;
      RECT  310.645000 -0.085000  310.815000 0.085000 ;
      RECT  310.645000  2.635000  310.815000 2.805000 ;
      RECT  311.105000 -0.085000  311.275000 0.085000 ;
      RECT  311.105000  2.635000  311.275000 2.805000 ;
      RECT  311.565000 -0.085000  311.735000 0.085000 ;
      RECT  311.565000  2.635000  311.735000 2.805000 ;
      RECT  312.025000 -0.085000  312.195000 0.085000 ;
      RECT  312.025000  2.635000  312.195000 2.805000 ;
      RECT  312.485000 -0.085000  312.655000 0.085000 ;
      RECT  312.485000  2.635000  312.655000 2.805000 ;
      RECT  312.945000 -0.085000  313.115000 0.085000 ;
      RECT  312.945000  2.635000  313.115000 2.805000 ;
      RECT  313.405000 -0.085000  313.575000 0.085000 ;
      RECT  313.405000  2.635000  313.575000 2.805000 ;
      RECT  313.865000 -0.085000  314.035000 0.085000 ;
      RECT  313.865000  2.635000  314.035000 2.805000 ;
      RECT  314.325000 -0.085000  314.495000 0.085000 ;
      RECT  314.325000  2.635000  314.495000 2.805000 ;
      RECT  314.785000 -0.085000  314.955000 0.085000 ;
      RECT  314.785000  2.635000  314.955000 2.805000 ;
      RECT  315.245000 -0.085000  315.415000 0.085000 ;
      RECT  315.245000  2.635000  315.415000 2.805000 ;
      RECT  315.705000 -0.085000  315.875000 0.085000 ;
      RECT  315.705000  2.635000  315.875000 2.805000 ;
      RECT  316.165000 -0.085000  316.335000 0.085000 ;
      RECT  316.165000  2.635000  316.335000 2.805000 ;
      RECT  316.625000 -0.085000  316.795000 0.085000 ;
      RECT  316.625000  2.635000  316.795000 2.805000 ;
      RECT  317.085000 -0.085000  317.255000 0.085000 ;
      RECT  317.085000  2.635000  317.255000 2.805000 ;
      RECT  317.545000 -0.085000  317.715000 0.085000 ;
      RECT  317.545000  2.635000  317.715000 2.805000 ;
      RECT  318.005000 -0.085000  318.175000 0.085000 ;
      RECT  318.005000  2.635000  318.175000 2.805000 ;
      RECT  318.465000 -0.085000  318.635000 0.085000 ;
      RECT  318.465000  2.635000  318.635000 2.805000 ;
      RECT  318.925000 -0.085000  319.095000 0.085000 ;
      RECT  318.925000  2.635000  319.095000 2.805000 ;
      RECT  319.385000 -0.085000  319.555000 0.085000 ;
      RECT  319.385000  2.635000  319.555000 2.805000 ;
      RECT  319.845000 -0.085000  320.015000 0.085000 ;
      RECT  319.845000  2.635000  320.015000 2.805000 ;
      RECT  320.305000 -0.085000  320.475000 0.085000 ;
      RECT  320.305000  2.635000  320.475000 2.805000 ;
      RECT  320.765000 -0.085000  320.935000 0.085000 ;
      RECT  320.765000  2.635000  320.935000 2.805000 ;
      RECT  321.225000 -0.085000  321.395000 0.085000 ;
      RECT  321.225000  2.635000  321.395000 2.805000 ;
      RECT  321.685000 -0.085000  321.855000 0.085000 ;
      RECT  321.685000  2.635000  321.855000 2.805000 ;
      RECT  322.145000 -0.085000  322.315000 0.085000 ;
      RECT  322.145000  2.635000  322.315000 2.805000 ;
      RECT  322.605000 -0.085000  322.775000 0.085000 ;
      RECT  322.605000  2.635000  322.775000 2.805000 ;
      RECT  323.065000 -0.085000  323.235000 0.085000 ;
      RECT  323.065000  2.635000  323.235000 2.805000 ;
      RECT  323.525000 -0.085000  323.695000 0.085000 ;
      RECT  323.525000  2.635000  323.695000 2.805000 ;
      RECT  323.985000 -0.085000  324.155000 0.085000 ;
      RECT  323.985000  2.635000  324.155000 2.805000 ;
      RECT  324.445000 -0.085000  324.615000 0.085000 ;
      RECT  324.445000  2.635000  324.615000 2.805000 ;
      RECT  324.905000 -0.085000  325.075000 0.085000 ;
      RECT  324.905000  2.635000  325.075000 2.805000 ;
      RECT  325.365000 -0.085000  325.535000 0.085000 ;
      RECT  325.365000  2.635000  325.535000 2.805000 ;
      RECT  325.825000 -0.085000  325.995000 0.085000 ;
      RECT  325.825000  2.635000  325.995000 2.805000 ;
      RECT  326.285000 -0.085000  326.455000 0.085000 ;
      RECT  326.285000  2.635000  326.455000 2.805000 ;
      RECT  326.745000 -0.085000  326.915000 0.085000 ;
      RECT  326.745000  2.635000  326.915000 2.805000 ;
      RECT  327.205000 -0.085000  327.375000 0.085000 ;
      RECT  327.205000  2.635000  327.375000 2.805000 ;
      RECT  327.665000 -0.085000  327.835000 0.085000 ;
      RECT  327.665000  2.635000  327.835000 2.805000 ;
      RECT  328.125000 -0.085000  328.295000 0.085000 ;
      RECT  328.125000  2.635000  328.295000 2.805000 ;
      RECT  328.585000 -0.085000  328.755000 0.085000 ;
      RECT  328.585000  2.635000  328.755000 2.805000 ;
      RECT  329.045000 -0.085000  329.215000 0.085000 ;
      RECT  329.045000  2.635000  329.215000 2.805000 ;
      RECT  329.505000 -0.085000  329.675000 0.085000 ;
      RECT  329.505000  2.635000  329.675000 2.805000 ;
      RECT  329.965000 -0.085000  330.135000 0.085000 ;
      RECT  329.965000  2.635000  330.135000 2.805000 ;
      RECT  330.425000 -0.085000  330.595000 0.085000 ;
      RECT  330.425000  2.635000  330.595000 2.805000 ;
      RECT  330.885000 -0.085000  331.055000 0.085000 ;
      RECT  330.885000  2.635000  331.055000 2.805000 ;
      RECT  331.345000 -0.085000  331.515000 0.085000 ;
      RECT  331.345000  2.635000  331.515000 2.805000 ;
      RECT  331.805000 -0.085000  331.975000 0.085000 ;
      RECT  331.805000  2.635000  331.975000 2.805000 ;
      RECT  332.265000 -0.085000  332.435000 0.085000 ;
      RECT  332.265000  2.635000  332.435000 2.805000 ;
      RECT  332.725000 -0.085000  332.895000 0.085000 ;
      RECT  332.725000  2.635000  332.895000 2.805000 ;
      RECT  333.185000 -0.085000  333.355000 0.085000 ;
      RECT  333.185000  2.635000  333.355000 2.805000 ;
      RECT  333.645000 -0.085000  333.815000 0.085000 ;
      RECT  333.645000  2.635000  333.815000 2.805000 ;
      RECT  334.105000 -0.085000  334.275000 0.085000 ;
      RECT  334.105000  2.635000  334.275000 2.805000 ;
      RECT  334.565000 -0.085000  334.735000 0.085000 ;
      RECT  334.565000  2.635000  334.735000 2.805000 ;
      RECT  335.025000 -0.085000  335.195000 0.085000 ;
      RECT  335.025000  2.635000  335.195000 2.805000 ;
      RECT  335.485000 -0.085000  335.655000 0.085000 ;
      RECT  335.485000  2.635000  335.655000 2.805000 ;
      RECT  335.945000 -0.085000  336.115000 0.085000 ;
      RECT  335.945000  2.635000  336.115000 2.805000 ;
      RECT  336.405000 -0.085000  336.575000 0.085000 ;
      RECT  336.405000  2.635000  336.575000 2.805000 ;
      RECT  336.865000 -0.085000  337.035000 0.085000 ;
      RECT  336.865000  2.635000  337.035000 2.805000 ;
      RECT  337.325000 -0.085000  337.495000 0.085000 ;
      RECT  337.325000  2.635000  337.495000 2.805000 ;
      RECT  337.785000 -0.085000  337.955000 0.085000 ;
      RECT  337.785000  2.635000  337.955000 2.805000 ;
      RECT  338.245000 -0.085000  338.415000 0.085000 ;
      RECT  338.245000  2.635000  338.415000 2.805000 ;
      RECT  338.705000 -0.085000  338.875000 0.085000 ;
      RECT  338.705000  2.635000  338.875000 2.805000 ;
      RECT  339.165000 -0.085000  339.335000 0.085000 ;
      RECT  339.165000  2.635000  339.335000 2.805000 ;
      RECT  339.625000 -0.085000  339.795000 0.085000 ;
      RECT  339.625000  2.635000  339.795000 2.805000 ;
      RECT  340.085000 -0.085000  340.255000 0.085000 ;
      RECT  340.085000  2.635000  340.255000 2.805000 ;
      RECT  340.545000 -0.085000  340.715000 0.085000 ;
      RECT  340.545000  2.635000  340.715000 2.805000 ;
      RECT  341.005000 -0.085000  341.175000 0.085000 ;
      RECT  341.005000  2.635000  341.175000 2.805000 ;
      RECT  341.465000 -0.085000  341.635000 0.085000 ;
      RECT  341.465000  2.635000  341.635000 2.805000 ;
      RECT  341.925000 -0.085000  342.095000 0.085000 ;
      RECT  341.925000  2.635000  342.095000 2.805000 ;
      RECT  342.385000 -0.085000  342.555000 0.085000 ;
      RECT  342.385000  2.635000  342.555000 2.805000 ;
      RECT  342.845000 -0.085000  343.015000 0.085000 ;
      RECT  342.845000  2.635000  343.015000 2.805000 ;
      RECT  343.305000 -0.085000  343.475000 0.085000 ;
      RECT  343.305000  2.635000  343.475000 2.805000 ;
      RECT  343.765000 -0.085000  343.935000 0.085000 ;
      RECT  343.765000  2.635000  343.935000 2.805000 ;
      RECT  344.225000 -0.085000  344.395000 0.085000 ;
      RECT  344.225000  2.635000  344.395000 2.805000 ;
      RECT  344.685000 -0.085000  344.855000 0.085000 ;
      RECT  344.685000  2.635000  344.855000 2.805000 ;
      RECT  345.145000 -0.085000  345.315000 0.085000 ;
      RECT  345.145000  2.635000  345.315000 2.805000 ;
      RECT  345.605000 -0.085000  345.775000 0.085000 ;
      RECT  345.605000  2.635000  345.775000 2.805000 ;
      RECT  346.065000 -0.085000  346.235000 0.085000 ;
      RECT  346.065000  2.635000  346.235000 2.805000 ;
      RECT  346.525000 -0.085000  346.695000 0.085000 ;
      RECT  346.525000  2.635000  346.695000 2.805000 ;
      RECT  346.985000 -0.085000  347.155000 0.085000 ;
      RECT  346.985000  2.635000  347.155000 2.805000 ;
      RECT  347.445000 -0.085000  347.615000 0.085000 ;
      RECT  347.445000  2.635000  347.615000 2.805000 ;
      RECT  347.905000 -0.085000  348.075000 0.085000 ;
      RECT  347.905000  2.635000  348.075000 2.805000 ;
      RECT  348.365000 -0.085000  348.535000 0.085000 ;
      RECT  348.365000  2.635000  348.535000 2.805000 ;
      RECT  348.825000 -0.085000  348.995000 0.085000 ;
      RECT  348.825000  2.635000  348.995000 2.805000 ;
      RECT  349.285000 -0.085000  349.455000 0.085000 ;
      RECT  349.285000  2.635000  349.455000 2.805000 ;
      RECT  349.745000 -0.085000  349.915000 0.085000 ;
      RECT  349.745000  2.635000  349.915000 2.805000 ;
      RECT  350.205000 -0.085000  350.375000 0.085000 ;
      RECT  350.205000  2.635000  350.375000 2.805000 ;
      RECT  350.665000 -0.085000  350.835000 0.085000 ;
      RECT  350.665000  2.635000  350.835000 2.805000 ;
      RECT  351.125000 -0.085000  351.295000 0.085000 ;
      RECT  351.125000  2.635000  351.295000 2.805000 ;
      RECT  351.585000 -0.085000  351.755000 0.085000 ;
      RECT  351.585000  2.635000  351.755000 2.805000 ;
      RECT  352.045000 -0.085000  352.215000 0.085000 ;
      RECT  352.045000  2.635000  352.215000 2.805000 ;
      RECT  352.505000 -0.085000  352.675000 0.085000 ;
      RECT  352.505000  2.635000  352.675000 2.805000 ;
      RECT  352.965000 -0.085000  353.135000 0.085000 ;
      RECT  352.965000  2.635000  353.135000 2.805000 ;
      RECT  353.425000 -0.085000  353.595000 0.085000 ;
      RECT  353.425000  2.635000  353.595000 2.805000 ;
      RECT  353.885000 -0.085000  354.055000 0.085000 ;
      RECT  353.885000  2.635000  354.055000 2.805000 ;
      RECT  354.345000 -0.085000  354.515000 0.085000 ;
      RECT  354.345000  2.635000  354.515000 2.805000 ;
      RECT  354.805000 -0.085000  354.975000 0.085000 ;
      RECT  354.805000  2.635000  354.975000 2.805000 ;
      RECT  355.265000 -0.085000  355.435000 0.085000 ;
      RECT  355.265000  2.635000  355.435000 2.805000 ;
      RECT  355.725000 -0.085000  355.895000 0.085000 ;
      RECT  355.725000  2.635000  355.895000 2.805000 ;
      RECT  356.185000 -0.085000  356.355000 0.085000 ;
      RECT  356.185000  2.635000  356.355000 2.805000 ;
      RECT  356.645000 -0.085000  356.815000 0.085000 ;
      RECT  356.645000  2.635000  356.815000 2.805000 ;
      RECT  357.105000 -0.085000  357.275000 0.085000 ;
      RECT  357.105000  2.635000  357.275000 2.805000 ;
      RECT  357.565000 -0.085000  357.735000 0.085000 ;
      RECT  357.565000  2.635000  357.735000 2.805000 ;
      RECT  358.025000 -0.085000  358.195000 0.085000 ;
      RECT  358.025000  2.635000  358.195000 2.805000 ;
      RECT  358.485000 -0.085000  358.655000 0.085000 ;
      RECT  358.485000  2.635000  358.655000 2.805000 ;
      RECT  358.945000 -0.085000  359.115000 0.085000 ;
      RECT  358.945000  2.635000  359.115000 2.805000 ;
      RECT  359.405000 -0.085000  359.575000 0.085000 ;
      RECT  359.405000  2.635000  359.575000 2.805000 ;
      RECT  359.865000 -0.085000  360.035000 0.085000 ;
      RECT  359.865000  2.635000  360.035000 2.805000 ;
      RECT  360.325000 -0.085000  360.495000 0.085000 ;
      RECT  360.325000  2.635000  360.495000 2.805000 ;
      RECT  360.785000 -0.085000  360.955000 0.085000 ;
      RECT  360.785000  2.635000  360.955000 2.805000 ;
      RECT  361.245000 -0.085000  361.415000 0.085000 ;
      RECT  361.245000  2.635000  361.415000 2.805000 ;
      RECT  361.705000 -0.085000  361.875000 0.085000 ;
      RECT  361.705000  2.635000  361.875000 2.805000 ;
      RECT  362.165000 -0.085000  362.335000 0.085000 ;
      RECT  362.165000  2.635000  362.335000 2.805000 ;
      RECT  362.625000 -0.085000  362.795000 0.085000 ;
      RECT  362.625000  2.635000  362.795000 2.805000 ;
      RECT  363.085000 -0.085000  363.255000 0.085000 ;
      RECT  363.085000  2.635000  363.255000 2.805000 ;
      RECT  363.545000 -0.085000  363.715000 0.085000 ;
      RECT  363.545000  2.635000  363.715000 2.805000 ;
      RECT  364.005000 -0.085000  364.175000 0.085000 ;
      RECT  364.005000  2.635000  364.175000 2.805000 ;
      RECT  364.465000 -0.085000  364.635000 0.085000 ;
      RECT  364.465000  2.635000  364.635000 2.805000 ;
      RECT  364.925000 -0.085000  365.095000 0.085000 ;
      RECT  364.925000  2.635000  365.095000 2.805000 ;
      RECT  365.385000 -0.085000  365.555000 0.085000 ;
      RECT  365.385000  2.635000  365.555000 2.805000 ;
      RECT  365.845000 -0.085000  366.015000 0.085000 ;
      RECT  365.845000  2.635000  366.015000 2.805000 ;
      RECT  366.305000 -0.085000  366.475000 0.085000 ;
      RECT  366.305000  2.635000  366.475000 2.805000 ;
      RECT  366.765000 -0.085000  366.935000 0.085000 ;
      RECT  366.765000  2.635000  366.935000 2.805000 ;
      RECT  367.225000 -0.085000  367.395000 0.085000 ;
      RECT  367.225000  2.635000  367.395000 2.805000 ;
      RECT  367.685000 -0.085000  367.855000 0.085000 ;
      RECT  367.685000  2.635000  367.855000 2.805000 ;
      RECT  368.145000 -0.085000  368.315000 0.085000 ;
      RECT  368.145000  2.635000  368.315000 2.805000 ;
      RECT  368.605000 -0.085000  368.775000 0.085000 ;
      RECT  368.605000  2.635000  368.775000 2.805000 ;
      RECT  369.065000 -0.085000  369.235000 0.085000 ;
      RECT  369.065000  2.635000  369.235000 2.805000 ;
      RECT  369.525000 -0.085000  369.695000 0.085000 ;
      RECT  369.525000  2.635000  369.695000 2.805000 ;
      RECT  369.985000 -0.085000  370.155000 0.085000 ;
      RECT  369.985000  2.635000  370.155000 2.805000 ;
      RECT  370.445000 -0.085000  370.615000 0.085000 ;
      RECT  370.445000  2.635000  370.615000 2.805000 ;
      RECT  370.905000 -0.085000  371.075000 0.085000 ;
      RECT  370.905000  2.635000  371.075000 2.805000 ;
      RECT  371.365000 -0.085000  371.535000 0.085000 ;
      RECT  371.365000  2.635000  371.535000 2.805000 ;
      RECT  371.825000 -0.085000  371.995000 0.085000 ;
      RECT  371.825000  2.635000  371.995000 2.805000 ;
      RECT  372.285000 -0.085000  372.455000 0.085000 ;
      RECT  372.285000  2.635000  372.455000 2.805000 ;
      RECT  372.745000 -0.085000  372.915000 0.085000 ;
      RECT  372.745000  2.635000  372.915000 2.805000 ;
      RECT  373.205000 -0.085000  373.375000 0.085000 ;
      RECT  373.205000  2.635000  373.375000 2.805000 ;
      RECT  373.665000 -0.085000  373.835000 0.085000 ;
      RECT  373.665000  2.635000  373.835000 2.805000 ;
      RECT  374.125000 -0.085000  374.295000 0.085000 ;
      RECT  374.125000  2.635000  374.295000 2.805000 ;
      RECT  374.585000 -0.085000  374.755000 0.085000 ;
      RECT  374.585000  2.635000  374.755000 2.805000 ;
      RECT  375.045000 -0.085000  375.215000 0.085000 ;
      RECT  375.045000  2.635000  375.215000 2.805000 ;
      RECT  375.505000 -0.085000  375.675000 0.085000 ;
      RECT  375.505000  2.635000  375.675000 2.805000 ;
      RECT  375.965000 -0.085000  376.135000 0.085000 ;
      RECT  375.965000  2.635000  376.135000 2.805000 ;
      RECT  376.425000 -0.085000  376.595000 0.085000 ;
      RECT  376.425000  2.635000  376.595000 2.805000 ;
      RECT  376.885000 -0.085000  377.055000 0.085000 ;
      RECT  376.885000  2.635000  377.055000 2.805000 ;
      RECT  377.345000 -0.085000  377.515000 0.085000 ;
      RECT  377.345000  2.635000  377.515000 2.805000 ;
      RECT  377.805000 -0.085000  377.975000 0.085000 ;
      RECT  377.805000  2.635000  377.975000 2.805000 ;
      RECT  378.265000 -0.085000  378.435000 0.085000 ;
      RECT  378.265000  2.635000  378.435000 2.805000 ;
      RECT  378.725000 -0.085000  378.895000 0.085000 ;
      RECT  378.725000  2.635000  378.895000 2.805000 ;
      RECT  379.185000 -0.085000  379.355000 0.085000 ;
      RECT  379.185000  2.635000  379.355000 2.805000 ;
      RECT  379.645000 -0.085000  379.815000 0.085000 ;
      RECT  379.645000  2.635000  379.815000 2.805000 ;
      RECT  380.105000 -0.085000  380.275000 0.085000 ;
      RECT  380.105000  2.635000  380.275000 2.805000 ;
      RECT  380.565000 -0.085000  380.735000 0.085000 ;
      RECT  380.565000  2.635000  380.735000 2.805000 ;
      RECT  381.025000 -0.085000  381.195000 0.085000 ;
      RECT  381.025000  2.635000  381.195000 2.805000 ;
      RECT  381.485000 -0.085000  381.655000 0.085000 ;
      RECT  381.485000  2.635000  381.655000 2.805000 ;
      RECT  381.945000 -0.085000  382.115000 0.085000 ;
      RECT  381.945000  2.635000  382.115000 2.805000 ;
      RECT  382.405000 -0.085000  382.575000 0.085000 ;
      RECT  382.405000  2.635000  382.575000 2.805000 ;
      RECT  382.865000 -0.085000  383.035000 0.085000 ;
      RECT  382.865000  2.635000  383.035000 2.805000 ;
      RECT  383.325000 -0.085000  383.495000 0.085000 ;
      RECT  383.325000  2.635000  383.495000 2.805000 ;
      RECT  383.785000 -0.085000  383.955000 0.085000 ;
      RECT  383.785000  2.635000  383.955000 2.805000 ;
      RECT  384.245000 -0.085000  384.415000 0.085000 ;
      RECT  384.245000  2.635000  384.415000 2.805000 ;
      RECT  384.705000 -0.085000  384.875000 0.085000 ;
      RECT  384.705000  2.635000  384.875000 2.805000 ;
      RECT  385.165000 -0.085000  385.335000 0.085000 ;
      RECT  385.165000  2.635000  385.335000 2.805000 ;
      RECT  385.625000 -0.085000  385.795000 0.085000 ;
      RECT  385.625000  2.635000  385.795000 2.805000 ;
      RECT  386.085000 -0.085000  386.255000 0.085000 ;
      RECT  386.085000  2.635000  386.255000 2.805000 ;
      RECT  386.545000 -0.085000  386.715000 0.085000 ;
      RECT  386.545000  2.635000  386.715000 2.805000 ;
      RECT  387.005000 -0.085000  387.175000 0.085000 ;
      RECT  387.005000  2.635000  387.175000 2.805000 ;
      RECT  387.465000 -0.085000  387.635000 0.085000 ;
      RECT  387.465000  2.635000  387.635000 2.805000 ;
      RECT  387.925000 -0.085000  388.095000 0.085000 ;
      RECT  387.925000  2.635000  388.095000 2.805000 ;
      RECT  388.385000 -0.085000  388.555000 0.085000 ;
      RECT  388.385000  2.635000  388.555000 2.805000 ;
      RECT  388.845000 -0.085000  389.015000 0.085000 ;
      RECT  388.845000  2.635000  389.015000 2.805000 ;
      RECT  389.305000 -0.085000  389.475000 0.085000 ;
      RECT  389.305000  2.635000  389.475000 2.805000 ;
      RECT  389.765000 -0.085000  389.935000 0.085000 ;
      RECT  389.765000  2.635000  389.935000 2.805000 ;
      RECT  390.225000 -0.085000  390.395000 0.085000 ;
      RECT  390.225000  2.635000  390.395000 2.805000 ;
      RECT  390.685000 -0.085000  390.855000 0.085000 ;
      RECT  390.685000  2.635000  390.855000 2.805000 ;
      RECT  391.145000 -0.085000  391.315000 0.085000 ;
      RECT  391.145000  2.635000  391.315000 2.805000 ;
      RECT  391.605000 -0.085000  391.775000 0.085000 ;
      RECT  391.605000  2.635000  391.775000 2.805000 ;
      RECT  392.065000 -0.085000  392.235000 0.085000 ;
      RECT  392.065000  2.635000  392.235000 2.805000 ;
      RECT  392.525000 -0.085000  392.695000 0.085000 ;
      RECT  392.525000  2.635000  392.695000 2.805000 ;
      RECT  392.985000 -0.085000  393.155000 0.085000 ;
      RECT  392.985000  2.635000  393.155000 2.805000 ;
      RECT  393.445000 -0.085000  393.615000 0.085000 ;
      RECT  393.445000  2.635000  393.615000 2.805000 ;
      RECT  393.905000 -0.085000  394.075000 0.085000 ;
      RECT  393.905000  2.635000  394.075000 2.805000 ;
      RECT  394.365000 -0.085000  394.535000 0.085000 ;
      RECT  394.365000  2.635000  394.535000 2.805000 ;
      RECT  394.825000 -0.085000  394.995000 0.085000 ;
      RECT  394.825000  2.635000  394.995000 2.805000 ;
      RECT  395.285000 -0.085000  395.455000 0.085000 ;
      RECT  395.285000  2.635000  395.455000 2.805000 ;
      RECT  395.745000 -0.085000  395.915000 0.085000 ;
      RECT  395.745000  2.635000  395.915000 2.805000 ;
      RECT  396.205000 -0.085000  396.375000 0.085000 ;
      RECT  396.205000  2.635000  396.375000 2.805000 ;
      RECT  396.665000 -0.085000  396.835000 0.085000 ;
      RECT  396.665000  2.635000  396.835000 2.805000 ;
      RECT  397.125000 -0.085000  397.295000 0.085000 ;
      RECT  397.125000  2.635000  397.295000 2.805000 ;
      RECT  397.585000 -0.085000  397.755000 0.085000 ;
      RECT  397.585000  2.635000  397.755000 2.805000 ;
      RECT  398.045000 -0.085000  398.215000 0.085000 ;
      RECT  398.045000  2.635000  398.215000 2.805000 ;
      RECT  398.505000 -0.085000  398.675000 0.085000 ;
      RECT  398.505000  2.635000  398.675000 2.805000 ;
      RECT  398.965000 -0.085000  399.135000 0.085000 ;
      RECT  398.965000  2.635000  399.135000 2.805000 ;
      RECT  399.425000 -0.085000  399.595000 0.085000 ;
      RECT  399.425000  2.635000  399.595000 2.805000 ;
      RECT  399.885000 -0.085000  400.055000 0.085000 ;
      RECT  399.885000  2.635000  400.055000 2.805000 ;
      RECT  400.345000 -0.085000  400.515000 0.085000 ;
      RECT  400.345000  2.635000  400.515000 2.805000 ;
      RECT  400.805000 -0.085000  400.975000 0.085000 ;
      RECT  400.805000  2.635000  400.975000 2.805000 ;
      RECT  401.265000 -0.085000  401.435000 0.085000 ;
      RECT  401.265000  2.635000  401.435000 2.805000 ;
      RECT  401.725000 -0.085000  401.895000 0.085000 ;
      RECT  401.725000  2.635000  401.895000 2.805000 ;
      RECT  402.185000 -0.085000  402.355000 0.085000 ;
      RECT  402.185000  2.635000  402.355000 2.805000 ;
      RECT  402.645000 -0.085000  402.815000 0.085000 ;
      RECT  402.645000  2.635000  402.815000 2.805000 ;
      RECT  403.105000 -0.085000  403.275000 0.085000 ;
      RECT  403.105000  2.635000  403.275000 2.805000 ;
      RECT  403.565000 -0.085000  403.735000 0.085000 ;
      RECT  403.565000  2.635000  403.735000 2.805000 ;
      RECT  404.025000 -0.085000  404.195000 0.085000 ;
      RECT  404.025000  2.635000  404.195000 2.805000 ;
      RECT  404.485000 -0.085000  404.655000 0.085000 ;
      RECT  404.485000  2.635000  404.655000 2.805000 ;
      RECT  404.945000 -0.085000  405.115000 0.085000 ;
      RECT  404.945000  2.635000  405.115000 2.805000 ;
      RECT  405.405000 -0.085000  405.575000 0.085000 ;
      RECT  405.405000  2.635000  405.575000 2.805000 ;
      RECT  405.865000 -0.085000  406.035000 0.085000 ;
      RECT  405.865000  2.635000  406.035000 2.805000 ;
      RECT  406.325000 -0.085000  406.495000 0.085000 ;
      RECT  406.325000  2.635000  406.495000 2.805000 ;
      RECT  406.785000 -0.085000  406.955000 0.085000 ;
      RECT  406.785000  2.635000  406.955000 2.805000 ;
      RECT  407.245000 -0.085000  407.415000 0.085000 ;
      RECT  407.245000  2.635000  407.415000 2.805000 ;
      RECT  407.705000 -0.085000  407.875000 0.085000 ;
      RECT  407.705000  2.635000  407.875000 2.805000 ;
      RECT  408.165000 -0.085000  408.335000 0.085000 ;
      RECT  408.165000  2.635000  408.335000 2.805000 ;
      RECT  408.625000 -0.085000  408.795000 0.085000 ;
      RECT  408.625000  2.635000  408.795000 2.805000 ;
      RECT  409.085000 -0.085000  409.255000 0.085000 ;
      RECT  409.085000  2.635000  409.255000 2.805000 ;
      RECT  409.545000 -0.085000  409.715000 0.085000 ;
      RECT  409.545000  2.635000  409.715000 2.805000 ;
      RECT  410.005000 -0.085000  410.175000 0.085000 ;
      RECT  410.005000  2.635000  410.175000 2.805000 ;
      RECT  410.465000 -0.085000  410.635000 0.085000 ;
      RECT  410.465000  2.635000  410.635000 2.805000 ;
      RECT  410.925000 -0.085000  411.095000 0.085000 ;
      RECT  410.925000  2.635000  411.095000 2.805000 ;
      RECT  411.385000 -0.085000  411.555000 0.085000 ;
      RECT  411.385000  2.635000  411.555000 2.805000 ;
      RECT  411.845000 -0.085000  412.015000 0.085000 ;
      RECT  411.845000  2.635000  412.015000 2.805000 ;
      RECT  412.305000 -0.085000  412.475000 0.085000 ;
      RECT  412.305000  2.635000  412.475000 2.805000 ;
      RECT  412.765000 -0.085000  412.935000 0.085000 ;
      RECT  412.765000  2.635000  412.935000 2.805000 ;
      RECT  413.225000 -0.085000  413.395000 0.085000 ;
      RECT  413.225000  2.635000  413.395000 2.805000 ;
      RECT  413.685000 -0.085000  413.855000 0.085000 ;
      RECT  413.685000  2.635000  413.855000 2.805000 ;
      RECT  414.145000 -0.085000  414.315000 0.085000 ;
      RECT  414.145000  2.635000  414.315000 2.805000 ;
      RECT  414.605000 -0.085000  414.775000 0.085000 ;
      RECT  414.605000  2.635000  414.775000 2.805000 ;
      RECT  415.065000 -0.085000  415.235000 0.085000 ;
      RECT  415.065000  2.635000  415.235000 2.805000 ;
      RECT  415.525000 -0.085000  415.695000 0.085000 ;
      RECT  415.525000  2.635000  415.695000 2.805000 ;
      RECT  415.985000 -0.085000  416.155000 0.085000 ;
      RECT  415.985000  2.635000  416.155000 2.805000 ;
      RECT  416.445000 -0.085000  416.615000 0.085000 ;
      RECT  416.445000  2.635000  416.615000 2.805000 ;
      RECT  416.905000 -0.085000  417.075000 0.085000 ;
      RECT  416.905000  2.635000  417.075000 2.805000 ;
      RECT  417.365000 -0.085000  417.535000 0.085000 ;
      RECT  417.365000  2.635000  417.535000 2.805000 ;
      RECT  417.825000 -0.085000  417.995000 0.085000 ;
      RECT  417.825000  2.635000  417.995000 2.805000 ;
      RECT  418.285000 -0.085000  418.455000 0.085000 ;
      RECT  418.285000  2.635000  418.455000 2.805000 ;
      RECT  418.745000 -0.085000  418.915000 0.085000 ;
      RECT  418.745000  2.635000  418.915000 2.805000 ;
      RECT  419.205000 -0.085000  419.375000 0.085000 ;
      RECT  419.205000  2.635000  419.375000 2.805000 ;
      RECT  419.665000 -0.085000  419.835000 0.085000 ;
      RECT  419.665000  2.635000  419.835000 2.805000 ;
      RECT  420.125000 -0.085000  420.295000 0.085000 ;
      RECT  420.125000  2.635000  420.295000 2.805000 ;
      RECT  420.585000 -0.085000  420.755000 0.085000 ;
      RECT  420.585000  2.635000  420.755000 2.805000 ;
      RECT  421.045000 -0.085000  421.215000 0.085000 ;
      RECT  421.045000  2.635000  421.215000 2.805000 ;
      RECT  421.505000 -0.085000  421.675000 0.085000 ;
      RECT  421.505000  2.635000  421.675000 2.805000 ;
      RECT  421.965000 -0.085000  422.135000 0.085000 ;
      RECT  421.965000  2.635000  422.135000 2.805000 ;
      RECT  422.425000 -0.085000  422.595000 0.085000 ;
      RECT  422.425000  2.635000  422.595000 2.805000 ;
      RECT  422.885000 -0.085000  423.055000 0.085000 ;
      RECT  422.885000  2.635000  423.055000 2.805000 ;
      RECT  423.345000 -0.085000  423.515000 0.085000 ;
      RECT  423.345000  2.635000  423.515000 2.805000 ;
      RECT  423.805000 -0.085000  423.975000 0.085000 ;
      RECT  423.805000  2.635000  423.975000 2.805000 ;
      RECT  424.265000 -0.085000  424.435000 0.085000 ;
      RECT  424.265000  2.635000  424.435000 2.805000 ;
      RECT  424.725000 -0.085000  424.895000 0.085000 ;
      RECT  424.725000  2.635000  424.895000 2.805000 ;
      RECT  425.185000 -0.085000  425.355000 0.085000 ;
      RECT  425.185000  2.635000  425.355000 2.805000 ;
      RECT  425.645000 -0.085000  425.815000 0.085000 ;
      RECT  425.645000  2.635000  425.815000 2.805000 ;
      RECT  426.105000 -0.085000  426.275000 0.085000 ;
      RECT  426.105000  2.635000  426.275000 2.805000 ;
      RECT  426.565000 -0.085000  426.735000 0.085000 ;
      RECT  426.565000  2.635000  426.735000 2.805000 ;
      RECT  427.025000 -0.085000  427.195000 0.085000 ;
      RECT  427.025000  2.635000  427.195000 2.805000 ;
      RECT  427.485000 -0.085000  427.655000 0.085000 ;
      RECT  427.485000  2.635000  427.655000 2.805000 ;
      RECT  427.945000 -0.085000  428.115000 0.085000 ;
      RECT  427.945000  2.635000  428.115000 2.805000 ;
      RECT  428.405000 -0.085000  428.575000 0.085000 ;
      RECT  428.405000  2.635000  428.575000 2.805000 ;
      RECT  428.865000 -0.085000  429.035000 0.085000 ;
      RECT  428.865000  2.635000  429.035000 2.805000 ;
      RECT  429.325000 -0.085000  429.495000 0.085000 ;
      RECT  429.325000  2.635000  429.495000 2.805000 ;
      RECT  429.785000 -0.085000  429.955000 0.085000 ;
      RECT  429.785000  2.635000  429.955000 2.805000 ;
      RECT  430.245000 -0.085000  430.415000 0.085000 ;
      RECT  430.245000  2.635000  430.415000 2.805000 ;
      RECT  430.705000 -0.085000  430.875000 0.085000 ;
      RECT  430.705000  2.635000  430.875000 2.805000 ;
      RECT  431.165000 -0.085000  431.335000 0.085000 ;
      RECT  431.165000  2.635000  431.335000 2.805000 ;
      RECT  431.625000 -0.085000  431.795000 0.085000 ;
      RECT  431.625000  2.635000  431.795000 2.805000 ;
      RECT  432.085000 -0.085000  432.255000 0.085000 ;
      RECT  432.085000  2.635000  432.255000 2.805000 ;
      RECT  432.545000 -0.085000  432.715000 0.085000 ;
      RECT  432.545000  2.635000  432.715000 2.805000 ;
      RECT  433.005000 -0.085000  433.175000 0.085000 ;
      RECT  433.005000  2.635000  433.175000 2.805000 ;
      RECT  433.465000 -0.085000  433.635000 0.085000 ;
      RECT  433.465000  2.635000  433.635000 2.805000 ;
      RECT  433.925000 -0.085000  434.095000 0.085000 ;
      RECT  433.925000  2.635000  434.095000 2.805000 ;
      RECT  434.385000 -0.085000  434.555000 0.085000 ;
      RECT  434.385000  2.635000  434.555000 2.805000 ;
      RECT  434.845000 -0.085000  435.015000 0.085000 ;
      RECT  434.845000  2.635000  435.015000 2.805000 ;
      RECT  435.305000 -0.085000  435.475000 0.085000 ;
      RECT  435.305000  2.635000  435.475000 2.805000 ;
      RECT  435.765000 -0.085000  435.935000 0.085000 ;
      RECT  435.765000  2.635000  435.935000 2.805000 ;
      RECT  436.225000 -0.085000  436.395000 0.085000 ;
      RECT  436.225000  2.635000  436.395000 2.805000 ;
      RECT  436.685000 -0.085000  436.855000 0.085000 ;
      RECT  436.685000  2.635000  436.855000 2.805000 ;
      RECT  437.145000 -0.085000  437.315000 0.085000 ;
      RECT  437.145000  2.635000  437.315000 2.805000 ;
      RECT  437.605000 -0.085000  437.775000 0.085000 ;
      RECT  437.605000  2.635000  437.775000 2.805000 ;
      RECT  438.065000 -0.085000  438.235000 0.085000 ;
      RECT  438.065000  2.635000  438.235000 2.805000 ;
      RECT  438.525000 -0.085000  438.695000 0.085000 ;
      RECT  438.525000  2.635000  438.695000 2.805000 ;
      RECT  438.985000 -0.085000  439.155000 0.085000 ;
      RECT  438.985000  2.635000  439.155000 2.805000 ;
      RECT  439.445000 -0.085000  439.615000 0.085000 ;
      RECT  439.445000  2.635000  439.615000 2.805000 ;
      RECT  439.905000 -0.085000  440.075000 0.085000 ;
      RECT  439.905000  2.635000  440.075000 2.805000 ;
      RECT  440.365000 -0.085000  440.535000 0.085000 ;
      RECT  440.365000  2.635000  440.535000 2.805000 ;
      RECT  440.825000 -0.085000  440.995000 0.085000 ;
      RECT  440.825000  2.635000  440.995000 2.805000 ;
      RECT  441.285000 -0.085000  441.455000 0.085000 ;
      RECT  441.285000  2.635000  441.455000 2.805000 ;
      RECT  441.745000 -0.085000  441.915000 0.085000 ;
      RECT  441.745000  2.635000  441.915000 2.805000 ;
      RECT  442.205000 -0.085000  442.375000 0.085000 ;
      RECT  442.205000  2.635000  442.375000 2.805000 ;
      RECT  442.665000 -0.085000  442.835000 0.085000 ;
      RECT  442.665000  2.635000  442.835000 2.805000 ;
      RECT  443.125000 -0.085000  443.295000 0.085000 ;
      RECT  443.125000  2.635000  443.295000 2.805000 ;
      RECT  443.585000 -0.085000  443.755000 0.085000 ;
      RECT  443.585000  2.635000  443.755000 2.805000 ;
      RECT  444.045000 -0.085000  444.215000 0.085000 ;
      RECT  444.045000  2.635000  444.215000 2.805000 ;
      RECT  444.505000 -0.085000  444.675000 0.085000 ;
      RECT  444.505000  2.635000  444.675000 2.805000 ;
      RECT  444.965000 -0.085000  445.135000 0.085000 ;
      RECT  444.965000  2.635000  445.135000 2.805000 ;
      RECT  445.425000 -0.085000  445.595000 0.085000 ;
      RECT  445.425000  2.635000  445.595000 2.805000 ;
      RECT  445.885000 -0.085000  446.055000 0.085000 ;
      RECT  445.885000  2.635000  446.055000 2.805000 ;
      RECT  446.345000 -0.085000  446.515000 0.085000 ;
      RECT  446.345000  2.635000  446.515000 2.805000 ;
      RECT  446.805000 -0.085000  446.975000 0.085000 ;
      RECT  446.805000  2.635000  446.975000 2.805000 ;
      RECT  447.265000 -0.085000  447.435000 0.085000 ;
      RECT  447.265000  2.635000  447.435000 2.805000 ;
      RECT  447.725000 -0.085000  447.895000 0.085000 ;
      RECT  447.725000  2.635000  447.895000 2.805000 ;
      RECT  448.185000 -0.085000  448.355000 0.085000 ;
      RECT  448.185000  2.635000  448.355000 2.805000 ;
      RECT  448.645000 -0.085000  448.815000 0.085000 ;
      RECT  448.645000  2.635000  448.815000 2.805000 ;
      RECT  449.105000 -0.085000  449.275000 0.085000 ;
      RECT  449.105000  2.635000  449.275000 2.805000 ;
      RECT  449.565000 -0.085000  449.735000 0.085000 ;
      RECT  449.565000  2.635000  449.735000 2.805000 ;
      RECT  450.025000 -0.085000  450.195000 0.085000 ;
      RECT  450.025000  2.635000  450.195000 2.805000 ;
      RECT  450.485000 -0.085000  450.655000 0.085000 ;
      RECT  450.485000  2.635000  450.655000 2.805000 ;
      RECT  450.945000 -0.085000  451.115000 0.085000 ;
      RECT  450.945000  2.635000  451.115000 2.805000 ;
      RECT  451.405000 -0.085000  451.575000 0.085000 ;
      RECT  451.405000  2.635000  451.575000 2.805000 ;
      RECT  451.865000 -0.085000  452.035000 0.085000 ;
      RECT  451.865000  2.635000  452.035000 2.805000 ;
      RECT  452.325000 -0.085000  452.495000 0.085000 ;
      RECT  452.325000  2.635000  452.495000 2.805000 ;
      RECT  452.785000 -0.085000  452.955000 0.085000 ;
      RECT  452.785000  2.635000  452.955000 2.805000 ;
      RECT  453.245000 -0.085000  453.415000 0.085000 ;
      RECT  453.245000  2.635000  453.415000 2.805000 ;
      RECT  453.705000 -0.085000  453.875000 0.085000 ;
      RECT  453.705000  2.635000  453.875000 2.805000 ;
      RECT  454.165000 -0.085000  454.335000 0.085000 ;
      RECT  454.165000  2.635000  454.335000 2.805000 ;
      RECT  454.625000 -0.085000  454.795000 0.085000 ;
      RECT  454.625000  2.635000  454.795000 2.805000 ;
      RECT  455.085000 -0.085000  455.255000 0.085000 ;
      RECT  455.085000  2.635000  455.255000 2.805000 ;
      RECT  455.545000 -0.085000  455.715000 0.085000 ;
      RECT  455.545000  2.635000  455.715000 2.805000 ;
      RECT  456.005000 -0.085000  456.175000 0.085000 ;
      RECT  456.005000  2.635000  456.175000 2.805000 ;
      RECT  456.465000 -0.085000  456.635000 0.085000 ;
      RECT  456.465000  2.635000  456.635000 2.805000 ;
      RECT  456.925000 -0.085000  457.095000 0.085000 ;
      RECT  456.925000  2.635000  457.095000 2.805000 ;
      RECT  457.385000 -0.085000  457.555000 0.085000 ;
      RECT  457.385000  2.635000  457.555000 2.805000 ;
      RECT  457.845000 -0.085000  458.015000 0.085000 ;
      RECT  457.845000  2.635000  458.015000 2.805000 ;
      RECT  458.305000 -0.085000  458.475000 0.085000 ;
      RECT  458.305000  2.635000  458.475000 2.805000 ;
      RECT  458.765000 -0.085000  458.935000 0.085000 ;
      RECT  458.765000  2.635000  458.935000 2.805000 ;
      RECT  459.225000 -0.085000  459.395000 0.085000 ;
      RECT  459.225000  2.635000  459.395000 2.805000 ;
      RECT  459.685000 -0.085000  459.855000 0.085000 ;
      RECT  459.685000  2.635000  459.855000 2.805000 ;
      RECT  460.145000 -0.085000  460.315000 0.085000 ;
      RECT  460.145000  2.635000  460.315000 2.805000 ;
      RECT  460.605000 -0.085000  460.775000 0.085000 ;
      RECT  460.605000  2.635000  460.775000 2.805000 ;
      RECT  461.065000 -0.085000  461.235000 0.085000 ;
      RECT  461.065000  2.635000  461.235000 2.805000 ;
      RECT  461.525000 -0.085000  461.695000 0.085000 ;
      RECT  461.525000  2.635000  461.695000 2.805000 ;
      RECT  461.985000 -0.085000  462.155000 0.085000 ;
      RECT  461.985000  2.635000  462.155000 2.805000 ;
      RECT  462.445000 -0.085000  462.615000 0.085000 ;
      RECT  462.445000  2.635000  462.615000 2.805000 ;
      RECT  462.905000 -0.085000  463.075000 0.085000 ;
      RECT  462.905000  2.635000  463.075000 2.805000 ;
      RECT  463.365000 -0.085000  463.535000 0.085000 ;
      RECT  463.365000  2.635000  463.535000 2.805000 ;
      RECT  463.825000 -0.085000  463.995000 0.085000 ;
      RECT  463.825000  2.635000  463.995000 2.805000 ;
      RECT  464.285000 -0.085000  464.455000 0.085000 ;
      RECT  464.285000  2.635000  464.455000 2.805000 ;
      RECT  464.745000 -0.085000  464.915000 0.085000 ;
      RECT  464.745000  2.635000  464.915000 2.805000 ;
      RECT  465.205000 -0.085000  465.375000 0.085000 ;
      RECT  465.205000  2.635000  465.375000 2.805000 ;
      RECT  465.665000 -0.085000  465.835000 0.085000 ;
      RECT  465.665000  2.635000  465.835000 2.805000 ;
      RECT  466.125000 -0.085000  466.295000 0.085000 ;
      RECT  466.125000  2.635000  466.295000 2.805000 ;
      RECT  466.585000 -0.085000  466.755000 0.085000 ;
      RECT  466.585000  2.635000  466.755000 2.805000 ;
      RECT  467.045000 -0.085000  467.215000 0.085000 ;
      RECT  467.045000  2.635000  467.215000 2.805000 ;
      RECT  467.505000 -0.085000  467.675000 0.085000 ;
      RECT  467.505000  2.635000  467.675000 2.805000 ;
      RECT  467.965000 -0.085000  468.135000 0.085000 ;
      RECT  467.965000  2.635000  468.135000 2.805000 ;
      RECT  468.425000 -0.085000  468.595000 0.085000 ;
      RECT  468.425000  2.635000  468.595000 2.805000 ;
      RECT  468.885000 -0.085000  469.055000 0.085000 ;
      RECT  468.885000  2.635000  469.055000 2.805000 ;
      RECT  469.345000 -0.085000  469.515000 0.085000 ;
      RECT  469.345000  2.635000  469.515000 2.805000 ;
      RECT  469.805000 -0.085000  469.975000 0.085000 ;
      RECT  469.805000  2.635000  469.975000 2.805000 ;
      RECT  470.265000 -0.085000  470.435000 0.085000 ;
      RECT  470.265000  2.635000  470.435000 2.805000 ;
      RECT  470.725000 -0.085000  470.895000 0.085000 ;
      RECT  470.725000  2.635000  470.895000 2.805000 ;
      RECT  471.185000 -0.085000  471.355000 0.085000 ;
      RECT  471.185000  2.635000  471.355000 2.805000 ;
      RECT  471.645000 -0.085000  471.815000 0.085000 ;
      RECT  471.645000  2.635000  471.815000 2.805000 ;
      RECT  472.105000 -0.085000  472.275000 0.085000 ;
      RECT  472.105000  2.635000  472.275000 2.805000 ;
      RECT  472.565000 -0.085000  472.735000 0.085000 ;
      RECT  472.565000  2.635000  472.735000 2.805000 ;
      RECT  473.025000 -0.085000  473.195000 0.085000 ;
      RECT  473.025000  2.635000  473.195000 2.805000 ;
      RECT  473.485000 -0.085000  473.655000 0.085000 ;
      RECT  473.485000  2.635000  473.655000 2.805000 ;
      RECT  473.945000 -0.085000  474.115000 0.085000 ;
      RECT  473.945000  2.635000  474.115000 2.805000 ;
      RECT  474.405000 -0.085000  474.575000 0.085000 ;
      RECT  474.405000  2.635000  474.575000 2.805000 ;
      RECT  474.865000 -0.085000  475.035000 0.085000 ;
      RECT  474.865000  2.635000  475.035000 2.805000 ;
      RECT  475.325000 -0.085000  475.495000 0.085000 ;
      RECT  475.325000  2.635000  475.495000 2.805000 ;
      RECT  475.475000  1.105000  475.645000 1.275000 ;
      RECT  475.785000 -0.085000  475.955000 0.085000 ;
      RECT  475.785000  2.635000  475.955000 2.805000 ;
      RECT  475.985000  1.105000  476.155000 1.275000 ;
      RECT  476.245000 -0.085000  476.415000 0.085000 ;
      RECT  476.245000  2.635000  476.415000 2.805000 ;
      RECT  476.705000 -0.085000  476.875000 0.085000 ;
      RECT  476.705000  2.635000  476.875000 2.805000 ;
      RECT  477.165000 -0.085000  477.335000 0.085000 ;
      RECT  477.165000  2.635000  477.335000 2.805000 ;
      RECT  477.625000 -0.085000  477.795000 0.085000 ;
      RECT  477.625000  2.635000  477.795000 2.805000 ;
      RECT  478.085000 -0.085000  478.255000 0.085000 ;
      RECT  478.085000  2.635000  478.255000 2.805000 ;
      RECT  478.545000 -0.085000  478.715000 0.085000 ;
      RECT  478.545000  2.635000  478.715000 2.805000 ;
      RECT  479.005000 -0.085000  479.175000 0.085000 ;
      RECT  479.005000  2.635000  479.175000 2.805000 ;
      RECT  479.465000 -0.085000  479.635000 0.085000 ;
      RECT  479.465000  2.635000  479.635000 2.805000 ;
      RECT  479.925000 -0.085000  480.095000 0.085000 ;
      RECT  479.925000  2.635000  480.095000 2.805000 ;
      RECT  480.385000 -0.085000  480.555000 0.085000 ;
      RECT  480.385000  2.635000  480.555000 2.805000 ;
      RECT  480.845000 -0.085000  481.015000 0.085000 ;
      RECT  480.845000  2.635000  481.015000 2.805000 ;
      RECT  481.305000 -0.085000  481.475000 0.085000 ;
      RECT  481.305000  2.635000  481.475000 2.805000 ;
      RECT  481.765000 -0.085000  481.935000 0.085000 ;
      RECT  481.765000  2.635000  481.935000 2.805000 ;
      RECT  482.225000 -0.085000  482.395000 0.085000 ;
      RECT  482.225000  2.635000  482.395000 2.805000 ;
      RECT  482.685000 -0.085000  482.855000 0.085000 ;
      RECT  482.685000  2.635000  482.855000 2.805000 ;
      RECT  483.145000 -0.085000  483.315000 0.085000 ;
      RECT  483.145000  2.635000  483.315000 2.805000 ;
      RECT  483.605000 -0.085000  483.775000 0.085000 ;
      RECT  483.605000  2.635000  483.775000 2.805000 ;
      RECT  484.065000 -0.085000  484.235000 0.085000 ;
      RECT  484.065000  2.635000  484.235000 2.805000 ;
      RECT  484.195000  1.105000  484.365000 1.275000 ;
      RECT  484.525000 -0.085000  484.695000 0.085000 ;
      RECT  484.525000  2.635000  484.695000 2.805000 ;
      RECT  484.705000  1.105000  484.875000 1.275000 ;
      RECT  484.985000 -0.085000  485.155000 0.085000 ;
      RECT  484.985000  2.635000  485.155000 2.805000 ;
      RECT  485.445000 -0.085000  485.615000 0.085000 ;
      RECT  485.445000  2.635000  485.615000 2.805000 ;
      RECT  485.905000 -0.085000  486.075000 0.085000 ;
      RECT  485.905000  2.635000  486.075000 2.805000 ;
      RECT  486.365000 -0.085000  486.535000 0.085000 ;
      RECT  486.365000  2.635000  486.535000 2.805000 ;
      RECT  486.825000 -0.085000  486.995000 0.085000 ;
      RECT  486.825000  2.635000  486.995000 2.805000 ;
      RECT  487.285000 -0.085000  487.455000 0.085000 ;
      RECT  487.285000  2.635000  487.455000 2.805000 ;
      RECT  487.745000 -0.085000  487.915000 0.085000 ;
      RECT  487.745000  2.635000  487.915000 2.805000 ;
      RECT  488.205000 -0.085000  488.375000 0.085000 ;
      RECT  488.205000  2.635000  488.375000 2.805000 ;
      RECT  488.665000 -0.085000  488.835000 0.085000 ;
      RECT  488.665000  2.635000  488.835000 2.805000 ;
      RECT  489.125000 -0.085000  489.295000 0.085000 ;
      RECT  489.125000  2.635000  489.295000 2.805000 ;
      RECT  489.585000 -0.085000  489.755000 0.085000 ;
      RECT  489.585000  2.635000  489.755000 2.805000 ;
      RECT  490.045000 -0.085000  490.215000 0.085000 ;
      RECT  490.045000  2.635000  490.215000 2.805000 ;
      RECT  490.505000 -0.085000  490.675000 0.085000 ;
      RECT  490.505000  2.635000  490.675000 2.805000 ;
      RECT  490.965000 -0.085000  491.135000 0.085000 ;
      RECT  490.965000  2.635000  491.135000 2.805000 ;
      RECT  491.425000 -0.085000  491.595000 0.085000 ;
      RECT  491.425000  2.635000  491.595000 2.805000 ;
      RECT  491.885000 -0.085000  492.055000 0.085000 ;
      RECT  491.885000  2.635000  492.055000 2.805000 ;
      RECT  492.345000 -0.085000  492.515000 0.085000 ;
      RECT  492.345000  2.635000  492.515000 2.805000 ;
      RECT  492.805000 -0.085000  492.975000 0.085000 ;
      RECT  492.805000  2.635000  492.975000 2.805000 ;
      RECT  493.265000 -0.085000  493.435000 0.085000 ;
      RECT  493.265000  2.635000  493.435000 2.805000 ;
      RECT  493.725000 -0.085000  493.895000 0.085000 ;
      RECT  493.725000  2.635000  493.895000 2.805000 ;
      RECT  494.185000 -0.085000  494.355000 0.085000 ;
      RECT  494.185000  2.635000  494.355000 2.805000 ;
      RECT  494.645000 -0.085000  494.815000 0.085000 ;
      RECT  494.645000  2.635000  494.815000 2.805000 ;
      RECT  495.105000 -0.085000  495.275000 0.085000 ;
      RECT  495.105000  2.635000  495.275000 2.805000 ;
      RECT  495.565000 -0.085000  495.735000 0.085000 ;
      RECT  495.565000  2.635000  495.735000 2.805000 ;
      RECT  496.025000 -0.085000  496.195000 0.085000 ;
      RECT  496.025000  2.635000  496.195000 2.805000 ;
      RECT  496.485000 -0.085000  496.655000 0.085000 ;
      RECT  496.485000  2.635000  496.655000 2.805000 ;
      RECT  496.945000 -0.085000  497.115000 0.085000 ;
      RECT  496.945000  2.635000  497.115000 2.805000 ;
      RECT  497.405000 -0.085000  497.575000 0.085000 ;
      RECT  497.405000  2.635000  497.575000 2.805000 ;
      RECT  497.865000 -0.085000  498.035000 0.085000 ;
      RECT  497.865000  2.635000  498.035000 2.805000 ;
      RECT  498.325000 -0.085000  498.495000 0.085000 ;
      RECT  498.325000  2.635000  498.495000 2.805000 ;
      RECT  498.785000 -0.085000  498.955000 0.085000 ;
      RECT  498.785000  2.635000  498.955000 2.805000 ;
      RECT  499.245000 -0.085000  499.415000 0.085000 ;
      RECT  499.245000  2.635000  499.415000 2.805000 ;
      RECT  499.705000 -0.085000  499.875000 0.085000 ;
      RECT  499.705000  2.635000  499.875000 2.805000 ;
      RECT  500.165000 -0.085000  500.335000 0.085000 ;
      RECT  500.165000  2.635000  500.335000 2.805000 ;
      RECT  500.625000 -0.085000  500.795000 0.085000 ;
      RECT  500.625000  2.635000  500.795000 2.805000 ;
      RECT  501.085000 -0.085000  501.255000 0.085000 ;
      RECT  501.085000  2.635000  501.255000 2.805000 ;
      RECT  501.545000 -0.085000  501.715000 0.085000 ;
      RECT  501.545000  2.635000  501.715000 2.805000 ;
      RECT  502.005000 -0.085000  502.175000 0.085000 ;
      RECT  502.005000  2.635000  502.175000 2.805000 ;
      RECT  502.465000 -0.085000  502.635000 0.085000 ;
      RECT  502.465000  2.635000  502.635000 2.805000 ;
      RECT  502.925000 -0.085000  503.095000 0.085000 ;
      RECT  502.925000  2.635000  503.095000 2.805000 ;
      RECT  503.385000 -0.085000  503.555000 0.085000 ;
      RECT  503.385000  2.635000  503.555000 2.805000 ;
      RECT  503.845000 -0.085000  504.015000 0.085000 ;
      RECT  503.845000  2.635000  504.015000 2.805000 ;
      RECT  504.305000 -0.085000  504.475000 0.085000 ;
      RECT  504.305000  2.635000  504.475000 2.805000 ;
      RECT  504.765000 -0.085000  504.935000 0.085000 ;
      RECT  504.765000  2.635000  504.935000 2.805000 ;
      RECT  505.225000 -0.085000  505.395000 0.085000 ;
      RECT  505.225000  2.635000  505.395000 2.805000 ;
      RECT  505.685000 -0.085000  505.855000 0.085000 ;
      RECT  505.685000  2.635000  505.855000 2.805000 ;
      RECT  506.145000 -0.085000  506.315000 0.085000 ;
      RECT  506.145000  2.635000  506.315000 2.805000 ;
      RECT  506.605000 -0.085000  506.775000 0.085000 ;
      RECT  506.605000  2.635000  506.775000 2.805000 ;
      RECT  507.065000 -0.085000  507.235000 0.085000 ;
      RECT  507.065000  2.635000  507.235000 2.805000 ;
      RECT  507.525000 -0.085000  507.695000 0.085000 ;
      RECT  507.525000  2.635000  507.695000 2.805000 ;
      RECT  507.985000 -0.085000  508.155000 0.085000 ;
      RECT  507.985000  2.635000  508.155000 2.805000 ;
      RECT  508.445000 -0.085000  508.615000 0.085000 ;
      RECT  508.445000  2.635000  508.615000 2.805000 ;
      RECT  508.500000  1.105000  508.670000 1.275000 ;
      RECT  508.905000 -0.085000  509.075000 0.085000 ;
      RECT  508.905000  2.635000  509.075000 2.805000 ;
      RECT  508.955000  1.785000  509.125000 1.955000 ;
      RECT  509.365000 -0.085000  509.535000 0.085000 ;
      RECT  509.365000  2.635000  509.535000 2.805000 ;
      RECT  509.825000 -0.085000  509.995000 0.085000 ;
      RECT  509.825000  2.635000  509.995000 2.805000 ;
      RECT  510.285000 -0.085000  510.455000 0.085000 ;
      RECT  510.285000  2.635000  510.455000 2.805000 ;
      RECT  510.320000  1.105000  510.490000 1.275000 ;
      RECT  510.565000  1.785000  510.735000 1.955000 ;
      RECT  510.745000 -0.085000  510.915000 0.085000 ;
      RECT  510.745000  2.635000  510.915000 2.805000 ;
      RECT  511.205000 -0.085000  511.375000 0.085000 ;
      RECT  511.205000  2.635000  511.375000 2.805000 ;
      RECT  511.665000 -0.085000  511.835000 0.085000 ;
      RECT  511.665000  2.635000  511.835000 2.805000 ;
      RECT  511.945000  0.765000  512.115000 0.935000 ;
      RECT  512.125000 -0.085000  512.295000 0.085000 ;
      RECT  512.125000  2.635000  512.295000 2.805000 ;
      RECT  512.305000  0.765000  512.475000 0.935000 ;
      RECT  512.585000 -0.085000  512.755000 0.085000 ;
      RECT  512.585000  2.635000  512.755000 2.805000 ;
      RECT  513.045000 -0.085000  513.215000 0.085000 ;
      RECT  513.045000  2.635000  513.215000 2.805000 ;
      RECT  513.505000 -0.085000  513.675000 0.085000 ;
      RECT  513.505000  2.635000  513.675000 2.805000 ;
      RECT  513.860000  1.105000  514.030000 1.275000 ;
      RECT  513.965000 -0.085000  514.135000 0.085000 ;
      RECT  513.965000  2.635000  514.135000 2.805000 ;
      RECT  514.310000  1.785000  514.480000 1.955000 ;
      RECT  514.425000 -0.085000  514.595000 0.085000 ;
      RECT  514.425000  2.635000  514.595000 2.805000 ;
      RECT  514.885000 -0.085000  515.055000 0.085000 ;
      RECT  514.885000  2.635000  515.055000 2.805000 ;
      RECT  515.345000 -0.085000  515.515000 0.085000 ;
      RECT  515.345000  2.635000  515.515000 2.805000 ;
      RECT  515.475000  0.765000  515.645000 0.935000 ;
      RECT  515.805000 -0.085000  515.975000 0.085000 ;
      RECT  515.805000  2.635000  515.975000 2.805000 ;
      RECT  516.265000 -0.085000  516.435000 0.085000 ;
      RECT  516.265000  2.635000  516.435000 2.805000 ;
      RECT  516.725000 -0.085000  516.895000 0.085000 ;
      RECT  516.725000  2.635000  516.895000 2.805000 ;
      RECT  517.185000 -0.085000  517.355000 0.085000 ;
      RECT  517.185000  2.635000  517.355000 2.805000 ;
      RECT  517.645000 -0.085000  517.815000 0.085000 ;
      RECT  517.645000  2.635000  517.815000 2.805000 ;
      RECT  518.105000 -0.085000  518.275000 0.085000 ;
      RECT  518.105000  2.635000  518.275000 2.805000 ;
      RECT  518.565000 -0.085000  518.735000 0.085000 ;
      RECT  518.565000  2.635000  518.735000 2.805000 ;
      RECT  518.620000  1.105000  518.790000 1.275000 ;
      RECT  519.025000 -0.085000  519.195000 0.085000 ;
      RECT  519.025000  2.635000  519.195000 2.805000 ;
      RECT  519.075000  1.785000  519.245000 1.955000 ;
      RECT  519.485000 -0.085000  519.655000 0.085000 ;
      RECT  519.485000  2.635000  519.655000 2.805000 ;
      RECT  519.945000 -0.085000  520.115000 0.085000 ;
      RECT  519.945000  2.635000  520.115000 2.805000 ;
      RECT  520.405000 -0.085000  520.575000 0.085000 ;
      RECT  520.405000  2.635000  520.575000 2.805000 ;
      RECT  520.440000  1.105000  520.610000 1.275000 ;
      RECT  520.685000  1.785000  520.855000 1.955000 ;
      RECT  520.865000 -0.085000  521.035000 0.085000 ;
      RECT  520.865000  2.635000  521.035000 2.805000 ;
      RECT  521.325000 -0.085000  521.495000 0.085000 ;
      RECT  521.325000  2.635000  521.495000 2.805000 ;
      RECT  521.785000 -0.085000  521.955000 0.085000 ;
      RECT  521.785000  2.635000  521.955000 2.805000 ;
      RECT  522.065000  0.765000  522.235000 0.935000 ;
      RECT  522.245000 -0.085000  522.415000 0.085000 ;
      RECT  522.245000  2.635000  522.415000 2.805000 ;
      RECT  522.425000  0.765000  522.595000 0.935000 ;
      RECT  522.705000 -0.085000  522.875000 0.085000 ;
      RECT  522.705000  2.635000  522.875000 2.805000 ;
      RECT  523.165000 -0.085000  523.335000 0.085000 ;
      RECT  523.165000  2.635000  523.335000 2.805000 ;
      RECT  523.625000 -0.085000  523.795000 0.085000 ;
      RECT  523.625000  2.635000  523.795000 2.805000 ;
      RECT  523.980000  1.105000  524.150000 1.275000 ;
      RECT  524.085000 -0.085000  524.255000 0.085000 ;
      RECT  524.085000  2.635000  524.255000 2.805000 ;
      RECT  524.430000  1.785000  524.600000 1.955000 ;
      RECT  524.545000 -0.085000  524.715000 0.085000 ;
      RECT  524.545000  2.635000  524.715000 2.805000 ;
      RECT  525.005000 -0.085000  525.175000 0.085000 ;
      RECT  525.005000  2.635000  525.175000 2.805000 ;
      RECT  525.465000 -0.085000  525.635000 0.085000 ;
      RECT  525.465000  2.635000  525.635000 2.805000 ;
      RECT  525.595000  0.765000  525.765000 0.935000 ;
      RECT  525.925000 -0.085000  526.095000 0.085000 ;
      RECT  525.925000  2.635000  526.095000 2.805000 ;
      RECT  526.385000 -0.085000  526.555000 0.085000 ;
      RECT  526.385000  2.635000  526.555000 2.805000 ;
      RECT  526.845000 -0.085000  527.015000 0.085000 ;
      RECT  526.845000  2.635000  527.015000 2.805000 ;
      RECT  527.305000 -0.085000  527.475000 0.085000 ;
      RECT  527.305000  2.635000  527.475000 2.805000 ;
      RECT  527.765000 -0.085000  527.935000 0.085000 ;
      RECT  527.765000  2.635000  527.935000 2.805000 ;
      RECT  528.225000 -0.085000  528.395000 0.085000 ;
      RECT  528.225000  2.635000  528.395000 2.805000 ;
      RECT  528.685000 -0.085000  528.855000 0.085000 ;
      RECT  528.685000  2.635000  528.855000 2.805000 ;
      RECT  529.145000 -0.085000  529.315000 0.085000 ;
      RECT  529.145000  2.635000  529.315000 2.805000 ;
      RECT  529.200000  1.105000  529.370000 1.275000 ;
      RECT  529.605000 -0.085000  529.775000 0.085000 ;
      RECT  529.605000  2.635000  529.775000 2.805000 ;
      RECT  529.655000  1.785000  529.825000 1.955000 ;
      RECT  530.065000 -0.085000  530.235000 0.085000 ;
      RECT  530.065000  2.635000  530.235000 2.805000 ;
      RECT  530.525000 -0.085000  530.695000 0.085000 ;
      RECT  530.525000  2.635000  530.695000 2.805000 ;
      RECT  530.985000 -0.085000  531.155000 0.085000 ;
      RECT  530.985000  2.635000  531.155000 2.805000 ;
      RECT  531.135000  1.105000  531.305000 1.275000 ;
      RECT  531.445000 -0.085000  531.615000 0.085000 ;
      RECT  531.445000  2.635000  531.615000 2.805000 ;
      RECT  531.645000  1.785000  531.815000 1.955000 ;
      RECT  531.905000 -0.085000  532.075000 0.085000 ;
      RECT  531.905000  2.635000  532.075000 2.805000 ;
      RECT  532.365000 -0.085000  532.535000 0.085000 ;
      RECT  532.365000  2.635000  532.535000 2.805000 ;
      RECT  532.825000 -0.085000  532.995000 0.085000 ;
      RECT  532.825000  0.765000  532.995000 0.935000 ;
      RECT  532.825000  2.635000  532.995000 2.805000 ;
      RECT  533.185000  0.765000  533.355000 0.935000 ;
      RECT  533.285000 -0.085000  533.455000 0.085000 ;
      RECT  533.285000  2.635000  533.455000 2.805000 ;
      RECT  533.745000 -0.085000  533.915000 0.085000 ;
      RECT  533.745000  2.635000  533.915000 2.805000 ;
      RECT  534.205000 -0.085000  534.375000 0.085000 ;
      RECT  534.205000  2.635000  534.375000 2.805000 ;
      RECT  534.665000 -0.085000  534.835000 0.085000 ;
      RECT  534.665000  2.635000  534.835000 2.805000 ;
      RECT  535.065000  1.105000  535.235000 1.275000 ;
      RECT  535.065000  1.785000  535.235000 1.955000 ;
      RECT  535.125000 -0.085000  535.295000 0.085000 ;
      RECT  535.125000  2.635000  535.295000 2.805000 ;
      RECT  535.585000 -0.085000  535.755000 0.085000 ;
      RECT  535.585000  2.635000  535.755000 2.805000 ;
      RECT  536.045000 -0.085000  536.215000 0.085000 ;
      RECT  536.045000  2.635000  536.215000 2.805000 ;
      RECT  536.410000  1.080000  536.580000 1.250000 ;
      RECT  536.505000 -0.085000  536.675000 0.085000 ;
      RECT  536.505000  2.635000  536.675000 2.805000 ;
      RECT  536.705000  0.765000  536.875000 0.935000 ;
      RECT  536.965000 -0.085000  537.135000 0.085000 ;
      RECT  536.965000  2.635000  537.135000 2.805000 ;
      RECT  537.425000 -0.085000  537.595000 0.085000 ;
      RECT  537.425000  2.635000  537.595000 2.805000 ;
      RECT  537.885000 -0.085000  538.055000 0.085000 ;
      RECT  537.885000  2.635000  538.055000 2.805000 ;
      RECT  538.345000 -0.085000  538.515000 0.085000 ;
      RECT  538.345000  2.635000  538.515000 2.805000 ;
      RECT  538.805000 -0.085000  538.975000 0.085000 ;
      RECT  538.805000  2.635000  538.975000 2.805000 ;
      RECT  539.265000 -0.085000  539.435000 0.085000 ;
      RECT  539.265000  2.635000  539.435000 2.805000 ;
      RECT  539.725000 -0.085000  539.895000 0.085000 ;
      RECT  539.725000  2.635000  539.895000 2.805000 ;
      RECT  540.185000 -0.085000  540.355000 0.085000 ;
      RECT  540.185000  2.635000  540.355000 2.805000 ;
      RECT  540.645000 -0.085000  540.815000 0.085000 ;
      RECT  540.645000  2.635000  540.815000 2.805000 ;
      RECT  541.105000 -0.085000  541.275000 0.085000 ;
      RECT  541.105000  2.635000  541.275000 2.805000 ;
      RECT  541.165000  1.740000  541.335000 1.910000 ;
      RECT  541.565000 -0.085000  541.735000 0.085000 ;
      RECT  541.565000  2.635000  541.735000 2.805000 ;
      RECT  541.665000  0.720000  541.835000 0.890000 ;
      RECT  542.025000 -0.085000  542.195000 0.085000 ;
      RECT  542.025000  2.635000  542.195000 2.805000 ;
      RECT  542.485000 -0.085000  542.655000 0.085000 ;
      RECT  542.485000  2.635000  542.655000 2.805000 ;
      RECT  542.945000 -0.085000  543.115000 0.085000 ;
      RECT  542.945000  2.635000  543.115000 2.805000 ;
      RECT  543.145000  1.740000  543.315000 1.910000 ;
      RECT  543.405000 -0.085000  543.575000 0.085000 ;
      RECT  543.405000  2.635000  543.575000 2.805000 ;
      RECT  543.655000  0.720000  543.825000 0.890000 ;
      RECT  543.865000 -0.085000  544.035000 0.085000 ;
      RECT  543.865000  2.635000  544.035000 2.805000 ;
      RECT  544.325000 -0.085000  544.495000 0.085000 ;
      RECT  544.325000  2.635000  544.495000 2.805000 ;
      RECT  544.780000  0.765000  544.950000 0.935000 ;
      RECT  544.785000 -0.085000  544.955000 0.085000 ;
      RECT  544.785000  2.635000  544.955000 2.805000 ;
      RECT  545.245000 -0.085000  545.415000 0.085000 ;
      RECT  545.245000  2.635000  545.415000 2.805000 ;
      RECT  545.705000 -0.085000  545.875000 0.085000 ;
      RECT  545.705000  2.635000  545.875000 2.805000 ;
      RECT  546.165000 -0.085000  546.335000 0.085000 ;
      RECT  546.165000  2.635000  546.335000 2.805000 ;
      RECT  546.205000  1.740000  546.375000 1.910000 ;
      RECT  546.225000  1.110000  546.395000 1.280000 ;
      RECT  546.625000 -0.085000  546.795000 0.085000 ;
      RECT  546.625000  2.635000  546.795000 2.805000 ;
      RECT  547.085000 -0.085000  547.255000 0.085000 ;
      RECT  547.085000  2.635000  547.255000 2.805000 ;
      RECT  547.545000 -0.085000  547.715000 0.085000 ;
      RECT  547.545000  2.635000  547.715000 2.805000 ;
      RECT  548.005000 -0.085000  548.175000 0.085000 ;
      RECT  548.005000  0.765000  548.175000 0.935000 ;
      RECT  548.005000  2.635000  548.175000 2.805000 ;
      RECT  548.465000 -0.085000  548.635000 0.085000 ;
      RECT  548.465000  2.635000  548.635000 2.805000 ;
      RECT  548.925000 -0.085000  549.095000 0.085000 ;
      RECT  548.925000  2.635000  549.095000 2.805000 ;
      RECT  549.385000 -0.085000  549.555000 0.085000 ;
      RECT  549.385000  2.635000  549.555000 2.805000 ;
      RECT  549.845000 -0.085000  550.015000 0.085000 ;
      RECT  549.845000  2.635000  550.015000 2.805000 ;
      RECT  550.305000 -0.085000  550.475000 0.085000 ;
      RECT  550.305000  2.635000  550.475000 2.805000 ;
      RECT  550.765000 -0.085000  550.935000 0.085000 ;
      RECT  550.765000  2.635000  550.935000 2.805000 ;
      RECT  551.225000 -0.085000  551.395000 0.085000 ;
      RECT  551.225000  2.635000  551.395000 2.805000 ;
      RECT  551.685000 -0.085000  551.855000 0.085000 ;
      RECT  551.685000  2.635000  551.855000 2.805000 ;
      RECT  551.745000  1.740000  551.915000 1.910000 ;
      RECT  552.145000 -0.085000  552.315000 0.085000 ;
      RECT  552.145000  2.635000  552.315000 2.805000 ;
      RECT  552.245000  0.720000  552.415000 0.890000 ;
      RECT  552.605000 -0.085000  552.775000 0.085000 ;
      RECT  552.605000  2.635000  552.775000 2.805000 ;
      RECT  553.065000 -0.085000  553.235000 0.085000 ;
      RECT  553.065000  2.635000  553.235000 2.805000 ;
      RECT  553.525000 -0.085000  553.695000 0.085000 ;
      RECT  553.525000  2.635000  553.695000 2.805000 ;
      RECT  553.725000  1.740000  553.895000 1.910000 ;
      RECT  553.985000 -0.085000  554.155000 0.085000 ;
      RECT  553.985000  2.635000  554.155000 2.805000 ;
      RECT  554.235000  0.720000  554.405000 0.890000 ;
      RECT  554.445000 -0.085000  554.615000 0.085000 ;
      RECT  554.445000  2.635000  554.615000 2.805000 ;
      RECT  554.905000 -0.085000  555.075000 0.085000 ;
      RECT  554.905000  2.635000  555.075000 2.805000 ;
      RECT  555.360000  0.765000  555.530000 0.935000 ;
      RECT  555.365000 -0.085000  555.535000 0.085000 ;
      RECT  555.365000  2.635000  555.535000 2.805000 ;
      RECT  555.825000 -0.085000  555.995000 0.085000 ;
      RECT  555.825000  2.635000  555.995000 2.805000 ;
      RECT  556.285000 -0.085000  556.455000 0.085000 ;
      RECT  556.285000  2.635000  556.455000 2.805000 ;
      RECT  556.745000 -0.085000  556.915000 0.085000 ;
      RECT  556.745000  2.635000  556.915000 2.805000 ;
      RECT  556.785000  1.740000  556.955000 1.910000 ;
      RECT  556.805000  1.110000  556.975000 1.280000 ;
      RECT  557.205000 -0.085000  557.375000 0.085000 ;
      RECT  557.205000  2.635000  557.375000 2.805000 ;
      RECT  557.665000 -0.085000  557.835000 0.085000 ;
      RECT  557.665000  2.635000  557.835000 2.805000 ;
      RECT  558.125000 -0.085000  558.295000 0.085000 ;
      RECT  558.125000  2.635000  558.295000 2.805000 ;
      RECT  558.585000 -0.085000  558.755000 0.085000 ;
      RECT  558.585000  0.765000  558.755000 0.935000 ;
      RECT  558.585000  2.635000  558.755000 2.805000 ;
      RECT  559.045000 -0.085000  559.215000 0.085000 ;
      RECT  559.045000  2.635000  559.215000 2.805000 ;
      RECT  559.505000 -0.085000  559.675000 0.085000 ;
      RECT  559.505000  2.635000  559.675000 2.805000 ;
      RECT  559.965000 -0.085000  560.135000 0.085000 ;
      RECT  559.965000  2.635000  560.135000 2.805000 ;
      RECT  560.425000 -0.085000  560.595000 0.085000 ;
      RECT  560.425000  2.635000  560.595000 2.805000 ;
      RECT  560.885000 -0.085000  561.055000 0.085000 ;
      RECT  560.885000  2.635000  561.055000 2.805000 ;
      RECT  561.345000 -0.085000  561.515000 0.085000 ;
      RECT  561.345000  2.635000  561.515000 2.805000 ;
      RECT  561.805000 -0.085000  561.975000 0.085000 ;
      RECT  561.805000  2.635000  561.975000 2.805000 ;
      RECT  562.265000 -0.085000  562.435000 0.085000 ;
      RECT  562.265000  2.635000  562.435000 2.805000 ;
      RECT  562.725000 -0.085000  562.895000 0.085000 ;
      RECT  562.725000  2.635000  562.895000 2.805000 ;
      RECT  562.785000  1.740000  562.955000 1.910000 ;
      RECT  563.185000 -0.085000  563.355000 0.085000 ;
      RECT  563.185000  2.635000  563.355000 2.805000 ;
      RECT  563.285000  0.720000  563.455000 0.890000 ;
      RECT  563.645000 -0.085000  563.815000 0.085000 ;
      RECT  563.645000  2.635000  563.815000 2.805000 ;
      RECT  564.105000 -0.085000  564.275000 0.085000 ;
      RECT  564.105000  2.635000  564.275000 2.805000 ;
      RECT  564.565000 -0.085000  564.735000 0.085000 ;
      RECT  564.565000  2.635000  564.735000 2.805000 ;
      RECT  564.765000  1.740000  564.935000 1.910000 ;
      RECT  565.025000 -0.085000  565.195000 0.085000 ;
      RECT  565.025000  2.635000  565.195000 2.805000 ;
      RECT  565.275000  0.720000  565.445000 0.890000 ;
      RECT  565.485000 -0.085000  565.655000 0.085000 ;
      RECT  565.485000  2.635000  565.655000 2.805000 ;
      RECT  565.945000 -0.085000  566.115000 0.085000 ;
      RECT  565.945000  2.635000  566.115000 2.805000 ;
      RECT  566.400000  0.765000  566.570000 0.935000 ;
      RECT  566.405000 -0.085000  566.575000 0.085000 ;
      RECT  566.405000  2.635000  566.575000 2.805000 ;
      RECT  566.865000 -0.085000  567.035000 0.085000 ;
      RECT  566.865000  2.635000  567.035000 2.805000 ;
      RECT  567.325000 -0.085000  567.495000 0.085000 ;
      RECT  567.325000  2.635000  567.495000 2.805000 ;
      RECT  567.785000 -0.085000  567.955000 0.085000 ;
      RECT  567.785000  2.635000  567.955000 2.805000 ;
      RECT  567.825000  1.740000  567.995000 1.910000 ;
      RECT  567.845000  1.110000  568.015000 1.280000 ;
      RECT  568.245000 -0.085000  568.415000 0.085000 ;
      RECT  568.245000  2.635000  568.415000 2.805000 ;
      RECT  568.705000 -0.085000  568.875000 0.085000 ;
      RECT  568.705000  2.635000  568.875000 2.805000 ;
      RECT  569.165000 -0.085000  569.335000 0.085000 ;
      RECT  569.165000  2.635000  569.335000 2.805000 ;
      RECT  569.625000 -0.085000  569.795000 0.085000 ;
      RECT  569.625000  0.765000  569.795000 0.935000 ;
      RECT  569.625000  2.635000  569.795000 2.805000 ;
      RECT  570.085000 -0.085000  570.255000 0.085000 ;
      RECT  570.085000  2.635000  570.255000 2.805000 ;
      RECT  570.545000 -0.085000  570.715000 0.085000 ;
      RECT  570.545000  2.635000  570.715000 2.805000 ;
      RECT  571.005000 -0.085000  571.175000 0.085000 ;
      RECT  571.005000  2.635000  571.175000 2.805000 ;
      RECT  571.465000 -0.085000  571.635000 0.085000 ;
      RECT  571.465000  2.635000  571.635000 2.805000 ;
      RECT  571.925000 -0.085000  572.095000 0.085000 ;
      RECT  571.925000  2.635000  572.095000 2.805000 ;
      RECT  572.385000 -0.085000  572.555000 0.085000 ;
      RECT  572.385000  2.635000  572.555000 2.805000 ;
      RECT  572.845000 -0.085000  573.015000 0.085000 ;
      RECT  572.845000  2.635000  573.015000 2.805000 ;
      RECT  573.305000 -0.085000  573.475000 0.085000 ;
      RECT  573.305000  2.635000  573.475000 2.805000 ;
      RECT  573.765000 -0.085000  573.935000 0.085000 ;
      RECT  573.765000  2.635000  573.935000 2.805000 ;
      RECT  574.225000 -0.085000  574.395000 0.085000 ;
      RECT  574.225000  2.635000  574.395000 2.805000 ;
      RECT  574.685000 -0.085000  574.855000 0.085000 ;
      RECT  574.685000  2.635000  574.855000 2.805000 ;
      RECT  575.145000 -0.085000  575.315000 0.085000 ;
      RECT  575.145000  2.635000  575.315000 2.805000 ;
      RECT  575.200000  1.445000  575.370000 1.615000 ;
      RECT  575.605000 -0.085000  575.775000 0.085000 ;
      RECT  575.605000  2.635000  575.775000 2.805000 ;
      RECT  575.710000  1.785000  575.880000 1.955000 ;
      RECT  576.065000 -0.085000  576.235000 0.085000 ;
      RECT  576.065000  2.635000  576.235000 2.805000 ;
      RECT  576.525000 -0.085000  576.695000 0.085000 ;
      RECT  576.525000  2.635000  576.695000 2.805000 ;
      RECT  576.985000 -0.085000  577.155000 0.085000 ;
      RECT  576.985000  2.635000  577.155000 2.805000 ;
      RECT  577.210000  1.785000  577.380000 1.955000 ;
      RECT  577.445000 -0.085000  577.615000 0.085000 ;
      RECT  577.445000  2.635000  577.615000 2.805000 ;
      RECT  577.715000  1.445000  577.885000 1.615000 ;
      RECT  577.905000 -0.085000  578.075000 0.085000 ;
      RECT  577.905000  2.635000  578.075000 2.805000 ;
      RECT  578.365000 -0.085000  578.535000 0.085000 ;
      RECT  578.365000  2.635000  578.535000 2.805000 ;
      RECT  578.825000 -0.085000  578.995000 0.085000 ;
      RECT  578.825000  2.635000  578.995000 2.805000 ;
      RECT  579.285000 -0.085000  579.455000 0.085000 ;
      RECT  579.285000  2.635000  579.455000 2.805000 ;
      RECT  579.745000 -0.085000  579.915000 0.085000 ;
      RECT  579.745000  2.635000  579.915000 2.805000 ;
      RECT  580.205000 -0.085000  580.375000 0.085000 ;
      RECT  580.205000  2.635000  580.375000 2.805000 ;
      RECT  580.665000 -0.085000  580.835000 0.085000 ;
      RECT  580.665000  2.635000  580.835000 2.805000 ;
      RECT  581.125000 -0.085000  581.295000 0.085000 ;
      RECT  581.125000  2.635000  581.295000 2.805000 ;
      RECT  581.585000 -0.085000  581.755000 0.085000 ;
      RECT  581.585000  2.635000  581.755000 2.805000 ;
      RECT  581.640000  1.445000  581.810000 1.615000 ;
      RECT  582.045000 -0.085000  582.215000 0.085000 ;
      RECT  582.045000  2.635000  582.215000 2.805000 ;
      RECT  582.150000  1.785000  582.320000 1.955000 ;
      RECT  582.505000 -0.085000  582.675000 0.085000 ;
      RECT  582.505000  2.635000  582.675000 2.805000 ;
      RECT  582.965000 -0.085000  583.135000 0.085000 ;
      RECT  582.965000  2.635000  583.135000 2.805000 ;
      RECT  583.425000 -0.085000  583.595000 0.085000 ;
      RECT  583.425000  2.635000  583.595000 2.805000 ;
      RECT  583.650000  1.785000  583.820000 1.955000 ;
      RECT  583.885000 -0.085000  584.055000 0.085000 ;
      RECT  583.885000  2.635000  584.055000 2.805000 ;
      RECT  584.155000  1.445000  584.325000 1.615000 ;
      RECT  584.345000 -0.085000  584.515000 0.085000 ;
      RECT  584.345000  2.635000  584.515000 2.805000 ;
      RECT  584.805000 -0.085000  584.975000 0.085000 ;
      RECT  584.805000  2.635000  584.975000 2.805000 ;
      RECT  585.265000 -0.085000  585.435000 0.085000 ;
      RECT  585.265000  2.635000  585.435000 2.805000 ;
      RECT  585.725000 -0.085000  585.895000 0.085000 ;
      RECT  585.725000  2.635000  585.895000 2.805000 ;
      RECT  586.185000 -0.085000  586.355000 0.085000 ;
      RECT  586.185000  2.635000  586.355000 2.805000 ;
      RECT  586.645000 -0.085000  586.815000 0.085000 ;
      RECT  586.645000  2.635000  586.815000 2.805000 ;
      RECT  587.105000 -0.085000  587.275000 0.085000 ;
      RECT  587.105000  2.635000  587.275000 2.805000 ;
      RECT  587.565000 -0.085000  587.735000 0.085000 ;
      RECT  587.565000  2.635000  587.735000 2.805000 ;
      RECT  588.025000 -0.085000  588.195000 0.085000 ;
      RECT  588.025000  2.635000  588.195000 2.805000 ;
      RECT  588.485000 -0.085000  588.655000 0.085000 ;
      RECT  588.485000  2.635000  588.655000 2.805000 ;
      RECT  588.540000  1.400000  588.710000 1.570000 ;
      RECT  588.945000 -0.085000  589.115000 0.085000 ;
      RECT  588.945000  2.635000  589.115000 2.805000 ;
      RECT  588.995000  1.770000  589.165000 1.940000 ;
      RECT  589.405000 -0.085000  589.575000 0.085000 ;
      RECT  589.405000  2.635000  589.575000 2.805000 ;
      RECT  589.865000 -0.085000  590.035000 0.085000 ;
      RECT  589.865000  2.635000  590.035000 2.805000 ;
      RECT  590.325000 -0.085000  590.495000 0.085000 ;
      RECT  590.325000  2.635000  590.495000 2.805000 ;
      RECT  590.550000  1.770000  590.720000 1.940000 ;
      RECT  590.785000 -0.085000  590.955000 0.085000 ;
      RECT  590.785000  2.635000  590.955000 2.805000 ;
      RECT  591.055000  1.400000  591.225000 1.570000 ;
      RECT  591.245000 -0.085000  591.415000 0.085000 ;
      RECT  591.245000  2.635000  591.415000 2.805000 ;
      RECT  591.705000 -0.085000  591.875000 0.085000 ;
      RECT  591.705000  2.635000  591.875000 2.805000 ;
      RECT  592.165000 -0.085000  592.335000 0.085000 ;
      RECT  592.165000  2.635000  592.335000 2.805000 ;
      RECT  592.625000 -0.085000  592.795000 0.085000 ;
      RECT  592.625000  2.635000  592.795000 2.805000 ;
      RECT  593.085000 -0.085000  593.255000 0.085000 ;
      RECT  593.085000  2.635000  593.255000 2.805000 ;
      RECT  593.545000 -0.085000  593.715000 0.085000 ;
      RECT  593.545000  2.635000  593.715000 2.805000 ;
      RECT  594.005000 -0.085000  594.175000 0.085000 ;
      RECT  594.005000  2.635000  594.175000 2.805000 ;
      RECT  594.465000 -0.085000  594.635000 0.085000 ;
      RECT  594.465000  2.635000  594.635000 2.805000 ;
      RECT  594.925000 -0.085000  595.095000 0.085000 ;
      RECT  594.925000  2.635000  595.095000 2.805000 ;
      RECT  595.385000 -0.085000  595.555000 0.085000 ;
      RECT  595.385000  2.635000  595.555000 2.805000 ;
      RECT  595.845000 -0.085000  596.015000 0.085000 ;
      RECT  595.845000  2.635000  596.015000 2.805000 ;
      RECT  596.305000 -0.085000  596.475000 0.085000 ;
      RECT  596.305000  2.635000  596.475000 2.805000 ;
      RECT  596.765000 -0.085000  596.935000 0.085000 ;
      RECT  596.765000  2.635000  596.935000 2.805000 ;
      RECT  597.225000 -0.085000  597.395000 0.085000 ;
      RECT  597.225000  2.635000  597.395000 2.805000 ;
      RECT  597.685000 -0.085000  597.855000 0.085000 ;
      RECT  597.685000  2.635000  597.855000 2.805000 ;
      RECT  598.145000 -0.085000  598.315000 0.085000 ;
      RECT  598.145000  2.635000  598.315000 2.805000 ;
      RECT  598.605000 -0.085000  598.775000 0.085000 ;
      RECT  598.605000  2.635000  598.775000 2.805000 ;
      RECT  599.065000 -0.085000  599.235000 0.085000 ;
      RECT  599.065000  2.635000  599.235000 2.805000 ;
      RECT  599.525000 -0.085000  599.695000 0.085000 ;
      RECT  599.525000  2.635000  599.695000 2.805000 ;
      RECT  599.985000 -0.085000  600.155000 0.085000 ;
      RECT  599.985000  2.635000  600.155000 2.805000 ;
      RECT  600.445000 -0.085000  600.615000 0.085000 ;
      RECT  600.445000  2.635000  600.615000 2.805000 ;
      RECT  600.905000 -0.085000  601.075000 0.085000 ;
      RECT  600.905000  2.635000  601.075000 2.805000 ;
      RECT  601.365000 -0.085000  601.535000 0.085000 ;
      RECT  601.365000  2.635000  601.535000 2.805000 ;
      RECT  601.825000 -0.085000  601.995000 0.085000 ;
      RECT  601.825000  2.635000  601.995000 2.805000 ;
      RECT  602.285000 -0.085000  602.455000 0.085000 ;
      RECT  602.285000  2.635000  602.455000 2.805000 ;
      RECT  602.745000 -0.085000  602.915000 0.085000 ;
      RECT  602.745000  2.635000  602.915000 2.805000 ;
      RECT  603.205000 -0.085000  603.375000 0.085000 ;
      RECT  603.205000  2.635000  603.375000 2.805000 ;
      RECT  603.665000 -0.085000  603.835000 0.085000 ;
      RECT  603.665000  2.635000  603.835000 2.805000 ;
      RECT  604.125000 -0.085000  604.295000 0.085000 ;
      RECT  604.125000  2.635000  604.295000 2.805000 ;
      RECT  604.585000 -0.085000  604.755000 0.085000 ;
      RECT  604.585000  2.635000  604.755000 2.805000 ;
      RECT  605.045000 -0.085000  605.215000 0.085000 ;
      RECT  605.045000  2.635000  605.215000 2.805000 ;
      RECT  605.505000 -0.085000  605.675000 0.085000 ;
      RECT  605.505000  2.635000  605.675000 2.805000 ;
      RECT  605.965000 -0.085000  606.135000 0.085000 ;
      RECT  605.965000  2.635000  606.135000 2.805000 ;
      RECT  606.425000 -0.085000  606.595000 0.085000 ;
      RECT  606.425000  2.635000  606.595000 2.805000 ;
      RECT  606.885000 -0.085000  607.055000 0.085000 ;
      RECT  606.885000  2.635000  607.055000 2.805000 ;
      RECT  607.345000 -0.085000  607.515000 0.085000 ;
      RECT  607.345000  2.635000  607.515000 2.805000 ;
      RECT  607.805000 -0.085000  607.975000 0.085000 ;
      RECT  607.805000  2.635000  607.975000 2.805000 ;
      RECT  608.265000 -0.085000  608.435000 0.085000 ;
      RECT  608.265000  2.635000  608.435000 2.805000 ;
      RECT  608.725000 -0.085000  608.895000 0.085000 ;
      RECT  608.725000  2.635000  608.895000 2.805000 ;
      RECT  609.185000 -0.085000  609.355000 0.085000 ;
      RECT  609.185000  2.635000  609.355000 2.805000 ;
      RECT  609.645000 -0.085000  609.815000 0.085000 ;
      RECT  609.645000  2.635000  609.815000 2.805000 ;
      RECT  610.105000 -0.085000  610.275000 0.085000 ;
      RECT  610.105000  2.635000  610.275000 2.805000 ;
      RECT  610.565000 -0.085000  610.735000 0.085000 ;
      RECT  610.565000  2.635000  610.735000 2.805000 ;
      RECT  611.025000 -0.085000  611.195000 0.085000 ;
      RECT  611.025000  2.635000  611.195000 2.805000 ;
      RECT  611.485000 -0.085000  611.655000 0.085000 ;
      RECT  611.485000  2.635000  611.655000 2.805000 ;
      RECT  611.490000  1.060000  611.660000 1.230000 ;
      RECT  611.945000 -0.085000  612.115000 0.085000 ;
      RECT  611.945000  2.635000  612.115000 2.805000 ;
      RECT  612.405000 -0.085000  612.575000 0.085000 ;
      RECT  612.405000  2.635000  612.575000 2.805000 ;
      RECT  612.865000 -0.085000  613.035000 0.085000 ;
      RECT  612.865000  2.635000  613.035000 2.805000 ;
      RECT  613.325000 -0.085000  613.495000 0.085000 ;
      RECT  613.325000  2.635000  613.495000 2.805000 ;
      RECT  613.785000 -0.085000  613.955000 0.085000 ;
      RECT  613.785000  2.635000  613.955000 2.805000 ;
      RECT  614.245000 -0.085000  614.415000 0.085000 ;
      RECT  614.245000  2.635000  614.415000 2.805000 ;
      RECT  614.705000 -0.085000  614.875000 0.085000 ;
      RECT  614.705000  2.635000  614.875000 2.805000 ;
      RECT  615.020000  1.060000  615.190000 1.230000 ;
      RECT  615.165000 -0.085000  615.335000 0.085000 ;
      RECT  615.165000  2.635000  615.335000 2.805000 ;
      RECT  615.625000 -0.085000  615.795000 0.085000 ;
      RECT  615.625000  2.635000  615.795000 2.805000 ;
      RECT  616.085000 -0.085000  616.255000 0.085000 ;
      RECT  616.085000  2.635000  616.255000 2.805000 ;
      RECT  616.545000 -0.085000  616.715000 0.085000 ;
      RECT  616.545000  2.635000  616.715000 2.805000 ;
      RECT  616.550000  1.105000  616.720000 1.275000 ;
      RECT  617.005000 -0.085000  617.175000 0.085000 ;
      RECT  617.005000  2.635000  617.175000 2.805000 ;
      RECT  617.465000 -0.085000  617.635000 0.085000 ;
      RECT  617.465000  2.635000  617.635000 2.805000 ;
      RECT  617.925000 -0.085000  618.095000 0.085000 ;
      RECT  617.925000  2.635000  618.095000 2.805000 ;
      RECT  618.385000 -0.085000  618.555000 0.085000 ;
      RECT  618.385000  2.635000  618.555000 2.805000 ;
      RECT  618.845000 -0.085000  619.015000 0.085000 ;
      RECT  618.845000  2.635000  619.015000 2.805000 ;
      RECT  619.305000 -0.085000  619.475000 0.085000 ;
      RECT  619.305000  2.635000  619.475000 2.805000 ;
      RECT  619.765000 -0.085000  619.935000 0.085000 ;
      RECT  619.765000  2.635000  619.935000 2.805000 ;
      RECT  620.225000 -0.085000  620.395000 0.085000 ;
      RECT  620.225000  2.635000  620.395000 2.805000 ;
      RECT  620.685000 -0.085000  620.855000 0.085000 ;
      RECT  620.685000  2.635000  620.855000 2.805000 ;
      RECT  621.110000  1.105000  621.280000 1.275000 ;
      RECT  621.145000 -0.085000  621.315000 0.085000 ;
      RECT  621.145000  2.635000  621.315000 2.805000 ;
      RECT  621.605000 -0.085000  621.775000 0.085000 ;
      RECT  621.605000  2.635000  621.775000 2.805000 ;
      RECT  622.065000 -0.085000  622.235000 0.085000 ;
      RECT  622.065000  2.635000  622.235000 2.805000 ;
      RECT  622.525000 -0.085000  622.695000 0.085000 ;
      RECT  622.525000  2.635000  622.695000 2.805000 ;
      RECT  622.985000 -0.085000  623.155000 0.085000 ;
      RECT  622.985000  2.635000  623.155000 2.805000 ;
      RECT  623.445000 -0.085000  623.615000 0.085000 ;
      RECT  623.445000  2.635000  623.615000 2.805000 ;
      RECT  623.905000 -0.085000  624.075000 0.085000 ;
      RECT  623.905000  2.635000  624.075000 2.805000 ;
      RECT  623.955000  1.060000  624.125000 1.230000 ;
      RECT  624.365000 -0.085000  624.535000 0.085000 ;
      RECT  624.365000  2.635000  624.535000 2.805000 ;
      RECT  624.825000 -0.085000  624.995000 0.085000 ;
      RECT  624.825000  2.635000  624.995000 2.805000 ;
      RECT  625.285000 -0.085000  625.455000 0.085000 ;
      RECT  625.285000  2.635000  625.455000 2.805000 ;
      RECT  625.745000 -0.085000  625.915000 0.085000 ;
      RECT  625.745000  2.635000  625.915000 2.805000 ;
      RECT  626.205000 -0.085000  626.375000 0.085000 ;
      RECT  626.205000  2.635000  626.375000 2.805000 ;
      RECT  626.665000 -0.085000  626.835000 0.085000 ;
      RECT  626.665000  2.635000  626.835000 2.805000 ;
      RECT  627.125000 -0.085000  627.295000 0.085000 ;
      RECT  627.125000  2.635000  627.295000 2.805000 ;
      RECT  627.585000 -0.085000  627.755000 0.085000 ;
      RECT  627.585000  2.635000  627.755000 2.805000 ;
      RECT  628.045000 -0.085000  628.215000 0.085000 ;
      RECT  628.045000  2.635000  628.215000 2.805000 ;
      RECT  628.505000 -0.085000  628.675000 0.085000 ;
      RECT  628.505000  2.635000  628.675000 2.805000 ;
      RECT  628.965000 -0.085000  629.135000 0.085000 ;
      RECT  628.965000  2.635000  629.135000 2.805000 ;
      RECT  629.425000 -0.085000  629.595000 0.085000 ;
      RECT  629.425000  2.635000  629.595000 2.805000 ;
      RECT  629.885000 -0.085000  630.055000 0.085000 ;
      RECT  629.885000  2.635000  630.055000 2.805000 ;
      RECT  630.345000 -0.085000  630.515000 0.085000 ;
      RECT  630.345000  2.635000  630.515000 2.805000 ;
      RECT  630.805000 -0.085000  630.975000 0.085000 ;
      RECT  630.805000  2.635000  630.975000 2.805000 ;
      RECT  630.930000  1.060000  631.100000 1.230000 ;
      RECT  631.265000 -0.085000  631.435000 0.085000 ;
      RECT  631.265000  2.635000  631.435000 2.805000 ;
      RECT  631.725000 -0.085000  631.895000 0.085000 ;
      RECT  631.725000  2.635000  631.895000 2.805000 ;
      RECT  632.185000 -0.085000  632.355000 0.085000 ;
      RECT  632.185000  2.635000  632.355000 2.805000 ;
      RECT  632.645000 -0.085000  632.815000 0.085000 ;
      RECT  632.645000  2.635000  632.815000 2.805000 ;
      RECT  633.105000 -0.085000  633.275000 0.085000 ;
      RECT  633.105000  2.635000  633.275000 2.805000 ;
      RECT  633.565000 -0.085000  633.735000 0.085000 ;
      RECT  633.565000  2.635000  633.735000 2.805000 ;
      RECT  634.025000 -0.085000  634.195000 0.085000 ;
      RECT  634.025000  2.635000  634.195000 2.805000 ;
      RECT  634.485000 -0.085000  634.655000 0.085000 ;
      RECT  634.485000  2.635000  634.655000 2.805000 ;
      RECT  634.945000 -0.085000  635.115000 0.085000 ;
      RECT  634.945000  2.635000  635.115000 2.805000 ;
      RECT  635.405000 -0.085000  635.575000 0.085000 ;
      RECT  635.405000  2.635000  635.575000 2.805000 ;
      RECT  635.865000 -0.085000  636.035000 0.085000 ;
      RECT  635.865000  2.635000  636.035000 2.805000 ;
      RECT  636.325000 -0.085000  636.495000 0.085000 ;
      RECT  636.325000  2.635000  636.495000 2.805000 ;
      RECT  636.785000 -0.085000  636.955000 0.085000 ;
      RECT  636.785000  2.635000  636.955000 2.805000 ;
      RECT  637.245000 -0.085000  637.415000 0.085000 ;
      RECT  637.245000  2.635000  637.415000 2.805000 ;
      RECT  637.705000 -0.085000  637.875000 0.085000 ;
      RECT  637.705000  2.635000  637.875000 2.805000 ;
      RECT  638.165000 -0.085000  638.335000 0.085000 ;
      RECT  638.165000  2.635000  638.335000 2.805000 ;
      RECT  638.625000 -0.085000  638.795000 0.085000 ;
      RECT  638.625000  2.635000  638.795000 2.805000 ;
      RECT  639.085000 -0.085000  639.255000 0.085000 ;
      RECT  639.085000  2.635000  639.255000 2.805000 ;
      RECT  639.545000 -0.085000  639.715000 0.085000 ;
      RECT  639.545000  2.635000  639.715000 2.805000 ;
      RECT  640.005000 -0.085000  640.175000 0.085000 ;
      RECT  640.005000  2.635000  640.175000 2.805000 ;
      RECT  640.465000 -0.085000  640.635000 0.085000 ;
      RECT  640.465000  2.635000  640.635000 2.805000 ;
      RECT  640.925000 -0.085000  641.095000 0.085000 ;
      RECT  640.925000  2.635000  641.095000 2.805000 ;
      RECT  641.385000 -0.085000  641.555000 0.085000 ;
      RECT  641.385000  2.635000  641.555000 2.805000 ;
      RECT  641.845000 -0.085000  642.015000 0.085000 ;
      RECT  641.845000  2.635000  642.015000 2.805000 ;
      RECT  642.305000 -0.085000  642.475000 0.085000 ;
      RECT  642.305000  2.635000  642.475000 2.805000 ;
      RECT  642.765000 -0.085000  642.935000 0.085000 ;
      RECT  642.765000  2.635000  642.935000 2.805000 ;
      RECT  643.225000 -0.085000  643.395000 0.085000 ;
      RECT  643.225000  2.635000  643.395000 2.805000 ;
      RECT  643.685000 -0.085000  643.855000 0.085000 ;
      RECT  643.685000  2.635000  643.855000 2.805000 ;
      RECT  644.145000 -0.085000  644.315000 0.085000 ;
      RECT  644.145000  2.635000  644.315000 2.805000 ;
      RECT  644.605000 -0.085000  644.775000 0.085000 ;
      RECT  644.605000  2.635000  644.775000 2.805000 ;
      RECT  645.065000 -0.085000  645.235000 0.085000 ;
      RECT  645.065000  2.635000  645.235000 2.805000 ;
      RECT  645.525000 -0.085000  645.695000 0.085000 ;
      RECT  645.525000  2.635000  645.695000 2.805000 ;
      RECT  645.985000 -0.085000  646.155000 0.085000 ;
      RECT  645.985000  2.635000  646.155000 2.805000 ;
      RECT  646.445000 -0.085000  646.615000 0.085000 ;
      RECT  646.445000  2.635000  646.615000 2.805000 ;
      RECT  646.905000 -0.085000  647.075000 0.085000 ;
      RECT  646.905000  2.635000  647.075000 2.805000 ;
      RECT  647.365000 -0.085000  647.535000 0.085000 ;
      RECT  647.365000  2.635000  647.535000 2.805000 ;
      RECT  647.825000 -0.085000  647.995000 0.085000 ;
      RECT  647.825000  2.635000  647.995000 2.805000 ;
      RECT  648.285000 -0.085000  648.455000 0.085000 ;
      RECT  648.285000  2.635000  648.455000 2.805000 ;
      RECT  648.745000 -0.085000  648.915000 0.085000 ;
      RECT  648.745000  2.635000  648.915000 2.805000 ;
      RECT  649.205000 -0.085000  649.375000 0.085000 ;
      RECT  649.205000  2.635000  649.375000 2.805000 ;
      RECT  649.665000 -0.085000  649.835000 0.085000 ;
      RECT  649.665000  2.635000  649.835000 2.805000 ;
      RECT  650.125000 -0.085000  650.295000 0.085000 ;
      RECT  650.125000  2.635000  650.295000 2.805000 ;
      RECT  650.585000 -0.085000  650.755000 0.085000 ;
      RECT  650.585000  2.635000  650.755000 2.805000 ;
      RECT  651.045000 -0.085000  651.215000 0.085000 ;
      RECT  651.045000  2.635000  651.215000 2.805000 ;
      RECT  651.505000 -0.085000  651.675000 0.085000 ;
      RECT  651.505000  2.635000  651.675000 2.805000 ;
      RECT  651.965000 -0.085000  652.135000 0.085000 ;
      RECT  651.965000  2.635000  652.135000 2.805000 ;
      RECT  652.425000 -0.085000  652.595000 0.085000 ;
      RECT  652.425000  2.635000  652.595000 2.805000 ;
      RECT  652.885000 -0.085000  653.055000 0.085000 ;
      RECT  652.885000  2.635000  653.055000 2.805000 ;
      RECT  653.345000 -0.085000  653.515000 0.085000 ;
      RECT  653.345000  2.635000  653.515000 2.805000 ;
      RECT  653.805000 -0.085000  653.975000 0.085000 ;
      RECT  653.805000  2.635000  653.975000 2.805000 ;
      RECT  654.265000 -0.085000  654.435000 0.085000 ;
      RECT  654.265000  2.635000  654.435000 2.805000 ;
      RECT  654.725000 -0.085000  654.895000 0.085000 ;
      RECT  654.725000  2.635000  654.895000 2.805000 ;
      RECT  655.185000 -0.085000  655.355000 0.085000 ;
      RECT  655.185000  2.635000  655.355000 2.805000 ;
      RECT  655.645000 -0.085000  655.815000 0.085000 ;
      RECT  655.645000  2.635000  655.815000 2.805000 ;
      RECT  656.105000 -0.085000  656.275000 0.085000 ;
      RECT  656.105000  2.635000  656.275000 2.805000 ;
      RECT  656.565000 -0.085000  656.735000 0.085000 ;
      RECT  656.565000  2.635000  656.735000 2.805000 ;
      RECT  657.025000 -0.085000  657.195000 0.085000 ;
      RECT  657.025000  2.635000  657.195000 2.805000 ;
      RECT  657.485000 -0.085000  657.655000 0.085000 ;
      RECT  657.485000  2.635000  657.655000 2.805000 ;
      RECT  657.945000 -0.085000  658.115000 0.085000 ;
      RECT  657.945000  2.635000  658.115000 2.805000 ;
      RECT  658.405000 -0.085000  658.575000 0.085000 ;
      RECT  658.405000  2.635000  658.575000 2.805000 ;
      RECT  658.865000 -0.085000  659.035000 0.085000 ;
      RECT  658.865000  2.635000  659.035000 2.805000 ;
      RECT  659.325000 -0.085000  659.495000 0.085000 ;
      RECT  659.325000  2.635000  659.495000 2.805000 ;
      RECT  659.785000 -0.085000  659.955000 0.085000 ;
      RECT  659.785000  2.635000  659.955000 2.805000 ;
      RECT  660.245000 -0.085000  660.415000 0.085000 ;
      RECT  660.245000  2.635000  660.415000 2.805000 ;
      RECT  660.705000 -0.085000  660.875000 0.085000 ;
      RECT  660.705000  2.635000  660.875000 2.805000 ;
      RECT  661.165000 -0.085000  661.335000 0.085000 ;
      RECT  661.165000  2.635000  661.335000 2.805000 ;
      RECT  661.625000 -0.085000  661.795000 0.085000 ;
      RECT  661.625000  2.635000  661.795000 2.805000 ;
      RECT  662.085000 -0.085000  662.255000 0.085000 ;
      RECT  662.085000  2.635000  662.255000 2.805000 ;
      RECT  662.545000 -0.085000  662.715000 0.085000 ;
      RECT  662.545000  2.635000  662.715000 2.805000 ;
      RECT  663.005000 -0.085000  663.175000 0.085000 ;
      RECT  663.005000  2.635000  663.175000 2.805000 ;
      RECT  663.465000 -0.085000  663.635000 0.085000 ;
      RECT  663.465000  2.635000  663.635000 2.805000 ;
      RECT  663.925000 -0.085000  664.095000 0.085000 ;
      RECT  663.925000  2.635000  664.095000 2.805000 ;
      RECT  664.385000 -0.085000  664.555000 0.085000 ;
      RECT  664.385000  2.635000  664.555000 2.805000 ;
      RECT  664.845000 -0.085000  665.015000 0.085000 ;
      RECT  664.845000  2.635000  665.015000 2.805000 ;
      RECT  665.305000 -0.085000  665.475000 0.085000 ;
      RECT  665.305000  2.635000  665.475000 2.805000 ;
      RECT  665.765000 -0.085000  665.935000 0.085000 ;
      RECT  665.765000  2.635000  665.935000 2.805000 ;
      RECT  666.225000 -0.085000  666.395000 0.085000 ;
      RECT  666.225000  2.635000  666.395000 2.805000 ;
      RECT  666.685000 -0.085000  666.855000 0.085000 ;
      RECT  666.685000  2.635000  666.855000 2.805000 ;
      RECT  667.145000 -0.085000  667.315000 0.085000 ;
      RECT  667.145000  2.635000  667.315000 2.805000 ;
      RECT  667.605000 -0.085000  667.775000 0.085000 ;
      RECT  667.605000  2.635000  667.775000 2.805000 ;
      RECT  668.065000 -0.085000  668.235000 0.085000 ;
      RECT  668.065000  2.635000  668.235000 2.805000 ;
      RECT  668.525000 -0.085000  668.695000 0.085000 ;
      RECT  668.525000  2.635000  668.695000 2.805000 ;
      RECT  668.985000 -0.085000  669.155000 0.085000 ;
      RECT  668.985000  2.635000  669.155000 2.805000 ;
      RECT  669.445000 -0.085000  669.615000 0.085000 ;
      RECT  669.445000  2.635000  669.615000 2.805000 ;
      RECT  669.905000 -0.085000  670.075000 0.085000 ;
      RECT  669.905000  2.635000  670.075000 2.805000 ;
      RECT  670.365000 -0.085000  670.535000 0.085000 ;
      RECT  670.365000  2.635000  670.535000 2.805000 ;
      RECT  670.825000 -0.085000  670.995000 0.085000 ;
      RECT  670.825000  2.635000  670.995000 2.805000 ;
      RECT  671.285000 -0.085000  671.455000 0.085000 ;
      RECT  671.285000  2.635000  671.455000 2.805000 ;
      RECT  671.745000 -0.085000  671.915000 0.085000 ;
      RECT  671.745000  2.635000  671.915000 2.805000 ;
      RECT  672.205000 -0.085000  672.375000 0.085000 ;
      RECT  672.205000  2.635000  672.375000 2.805000 ;
      RECT  672.665000 -0.085000  672.835000 0.085000 ;
      RECT  672.665000  2.635000  672.835000 2.805000 ;
      RECT  673.125000 -0.085000  673.295000 0.085000 ;
      RECT  673.125000  2.635000  673.295000 2.805000 ;
      RECT  673.585000 -0.085000  673.755000 0.085000 ;
      RECT  673.585000  2.635000  673.755000 2.805000 ;
      RECT  674.045000 -0.085000  674.215000 0.085000 ;
      RECT  674.045000  2.635000  674.215000 2.805000 ;
      RECT  674.505000 -0.085000  674.675000 0.085000 ;
      RECT  674.505000  2.635000  674.675000 2.805000 ;
      RECT  674.965000 -0.085000  675.135000 0.085000 ;
      RECT  674.965000  2.635000  675.135000 2.805000 ;
      RECT  675.425000 -0.085000  675.595000 0.085000 ;
      RECT  675.425000  2.635000  675.595000 2.805000 ;
      RECT  675.885000 -0.085000  676.055000 0.085000 ;
      RECT  675.885000  2.635000  676.055000 2.805000 ;
      RECT  676.345000 -0.085000  676.515000 0.085000 ;
      RECT  676.345000  2.635000  676.515000 2.805000 ;
      RECT  676.805000 -0.085000  676.975000 0.085000 ;
      RECT  676.805000  2.635000  676.975000 2.805000 ;
      RECT  677.265000 -0.085000  677.435000 0.085000 ;
      RECT  677.265000  2.635000  677.435000 2.805000 ;
      RECT  677.725000 -0.085000  677.895000 0.085000 ;
      RECT  677.725000  2.635000  677.895000 2.805000 ;
      RECT  678.185000 -0.085000  678.355000 0.085000 ;
      RECT  678.185000  2.635000  678.355000 2.805000 ;
      RECT  678.645000 -0.085000  678.815000 0.085000 ;
      RECT  678.645000  2.635000  678.815000 2.805000 ;
      RECT  679.105000 -0.085000  679.275000 0.085000 ;
      RECT  679.105000  2.635000  679.275000 2.805000 ;
      RECT  679.565000 -0.085000  679.735000 0.085000 ;
      RECT  679.565000  2.635000  679.735000 2.805000 ;
      RECT  680.025000 -0.085000  680.195000 0.085000 ;
      RECT  680.025000  2.635000  680.195000 2.805000 ;
      RECT  680.485000 -0.085000  680.655000 0.085000 ;
      RECT  680.485000  2.635000  680.655000 2.805000 ;
      RECT  680.945000 -0.085000  681.115000 0.085000 ;
      RECT  680.945000  2.635000  681.115000 2.805000 ;
      RECT  681.405000 -0.085000  681.575000 0.085000 ;
      RECT  681.405000  2.635000  681.575000 2.805000 ;
      RECT  681.865000 -0.085000  682.035000 0.085000 ;
      RECT  681.865000  2.635000  682.035000 2.805000 ;
      RECT  682.325000 -0.085000  682.495000 0.085000 ;
      RECT  682.325000  2.635000  682.495000 2.805000 ;
      RECT  682.785000 -0.085000  682.955000 0.085000 ;
      RECT  682.785000  2.635000  682.955000 2.805000 ;
      RECT  683.245000 -0.085000  683.415000 0.085000 ;
      RECT  683.245000  2.635000  683.415000 2.805000 ;
      RECT  683.705000 -0.085000  683.875000 0.085000 ;
      RECT  683.705000  2.635000  683.875000 2.805000 ;
      RECT  684.165000 -0.085000  684.335000 0.085000 ;
      RECT  684.165000  2.635000  684.335000 2.805000 ;
      RECT  684.625000 -0.085000  684.795000 0.085000 ;
      RECT  684.625000  2.635000  684.795000 2.805000 ;
      RECT  685.085000 -0.085000  685.255000 0.085000 ;
      RECT  685.085000  2.635000  685.255000 2.805000 ;
      RECT  685.545000 -0.085000  685.715000 0.085000 ;
      RECT  685.545000  2.635000  685.715000 2.805000 ;
      RECT  686.005000 -0.085000  686.175000 0.085000 ;
      RECT  686.005000  2.635000  686.175000 2.805000 ;
      RECT  686.465000 -0.085000  686.635000 0.085000 ;
      RECT  686.465000  2.635000  686.635000 2.805000 ;
      RECT  686.925000 -0.085000  687.095000 0.085000 ;
      RECT  686.925000  2.635000  687.095000 2.805000 ;
      RECT  687.385000 -0.085000  687.555000 0.085000 ;
      RECT  687.385000  2.635000  687.555000 2.805000 ;
      RECT  687.845000 -0.085000  688.015000 0.085000 ;
      RECT  687.845000  2.635000  688.015000 2.805000 ;
      RECT  688.305000 -0.085000  688.475000 0.085000 ;
      RECT  688.305000  2.635000  688.475000 2.805000 ;
      RECT  688.765000 -0.085000  688.935000 0.085000 ;
      RECT  688.765000  2.635000  688.935000 2.805000 ;
      RECT  689.225000 -0.085000  689.395000 0.085000 ;
      RECT  689.225000  2.635000  689.395000 2.805000 ;
      RECT  689.685000 -0.085000  689.855000 0.085000 ;
      RECT  689.685000  2.635000  689.855000 2.805000 ;
      RECT  690.145000 -0.085000  690.315000 0.085000 ;
      RECT  690.145000  2.635000  690.315000 2.805000 ;
      RECT  690.605000 -0.085000  690.775000 0.085000 ;
      RECT  690.605000  2.635000  690.775000 2.805000 ;
      RECT  691.065000 -0.085000  691.235000 0.085000 ;
      RECT  691.065000  2.635000  691.235000 2.805000 ;
      RECT  691.525000 -0.085000  691.695000 0.085000 ;
      RECT  691.525000  2.635000  691.695000 2.805000 ;
      RECT  691.985000 -0.085000  692.155000 0.085000 ;
      RECT  691.985000  2.635000  692.155000 2.805000 ;
      RECT  692.445000 -0.085000  692.615000 0.085000 ;
      RECT  692.445000  2.635000  692.615000 2.805000 ;
      RECT  692.905000 -0.085000  693.075000 0.085000 ;
      RECT  692.905000  2.635000  693.075000 2.805000 ;
      RECT  693.365000 -0.085000  693.535000 0.085000 ;
      RECT  693.365000  2.635000  693.535000 2.805000 ;
      RECT  693.825000 -0.085000  693.995000 0.085000 ;
      RECT  693.825000  2.635000  693.995000 2.805000 ;
      RECT  694.285000 -0.085000  694.455000 0.085000 ;
      RECT  694.285000  2.635000  694.455000 2.805000 ;
      RECT  694.745000 -0.085000  694.915000 0.085000 ;
      RECT  694.745000  2.635000  694.915000 2.805000 ;
      RECT  695.205000 -0.085000  695.375000 0.085000 ;
      RECT  695.205000  2.635000  695.375000 2.805000 ;
      RECT  695.665000 -0.085000  695.835000 0.085000 ;
      RECT  695.665000  2.635000  695.835000 2.805000 ;
      RECT  696.125000 -0.085000  696.295000 0.085000 ;
      RECT  696.125000  2.635000  696.295000 2.805000 ;
      RECT  696.585000 -0.085000  696.755000 0.085000 ;
      RECT  696.585000  2.635000  696.755000 2.805000 ;
      RECT  697.045000 -0.085000  697.215000 0.085000 ;
      RECT  697.045000  2.635000  697.215000 2.805000 ;
      RECT  697.505000 -0.085000  697.675000 0.085000 ;
      RECT  697.505000  2.635000  697.675000 2.805000 ;
      RECT  697.965000 -0.085000  698.135000 0.085000 ;
      RECT  697.965000  2.635000  698.135000 2.805000 ;
      RECT  698.425000 -0.085000  698.595000 0.085000 ;
      RECT  698.425000  2.635000  698.595000 2.805000 ;
      RECT  698.885000 -0.085000  699.055000 0.085000 ;
      RECT  698.885000  2.635000  699.055000 2.805000 ;
      RECT  699.345000 -0.085000  699.515000 0.085000 ;
      RECT  699.345000  2.635000  699.515000 2.805000 ;
      RECT  699.805000 -0.085000  699.975000 0.085000 ;
      RECT  699.805000  2.635000  699.975000 2.805000 ;
      RECT  700.265000 -0.085000  700.435000 0.085000 ;
      RECT  700.265000  2.635000  700.435000 2.805000 ;
      RECT  700.725000 -0.085000  700.895000 0.085000 ;
      RECT  700.725000  2.635000  700.895000 2.805000 ;
      RECT  701.185000 -0.085000  701.355000 0.085000 ;
      RECT  701.185000  2.635000  701.355000 2.805000 ;
      RECT  701.645000 -0.085000  701.815000 0.085000 ;
      RECT  701.645000  2.635000  701.815000 2.805000 ;
      RECT  702.105000 -0.085000  702.275000 0.085000 ;
      RECT  702.105000  2.635000  702.275000 2.805000 ;
      RECT  702.565000 -0.085000  702.735000 0.085000 ;
      RECT  702.565000  2.635000  702.735000 2.805000 ;
      RECT  703.025000 -0.085000  703.195000 0.085000 ;
      RECT  703.025000  2.635000  703.195000 2.805000 ;
      RECT  703.485000 -0.085000  703.655000 0.085000 ;
      RECT  703.485000  2.635000  703.655000 2.805000 ;
      RECT  703.945000 -0.085000  704.115000 0.085000 ;
      RECT  703.945000  2.635000  704.115000 2.805000 ;
      RECT  704.405000 -0.085000  704.575000 0.085000 ;
      RECT  704.405000  2.635000  704.575000 2.805000 ;
      RECT  704.865000 -0.085000  705.035000 0.085000 ;
      RECT  704.865000  2.635000  705.035000 2.805000 ;
      RECT  705.325000 -0.085000  705.495000 0.085000 ;
      RECT  705.325000  2.635000  705.495000 2.805000 ;
      RECT  705.785000 -0.085000  705.955000 0.085000 ;
      RECT  705.785000  2.635000  705.955000 2.805000 ;
      RECT  706.245000 -0.085000  706.415000 0.085000 ;
      RECT  706.245000  2.635000  706.415000 2.805000 ;
      RECT  706.705000 -0.085000  706.875000 0.085000 ;
      RECT  706.705000  2.635000  706.875000 2.805000 ;
      RECT  707.165000 -0.085000  707.335000 0.085000 ;
      RECT  707.165000  2.635000  707.335000 2.805000 ;
      RECT  707.625000 -0.085000  707.795000 0.085000 ;
      RECT  707.625000  2.635000  707.795000 2.805000 ;
      RECT  708.085000 -0.085000  708.255000 0.085000 ;
      RECT  708.085000  2.635000  708.255000 2.805000 ;
      RECT  708.545000 -0.085000  708.715000 0.085000 ;
      RECT  708.545000  2.635000  708.715000 2.805000 ;
      RECT  709.005000 -0.085000  709.175000 0.085000 ;
      RECT  709.005000  2.635000  709.175000 2.805000 ;
      RECT  709.465000 -0.085000  709.635000 0.085000 ;
      RECT  709.465000  2.635000  709.635000 2.805000 ;
      RECT  709.925000 -0.085000  710.095000 0.085000 ;
      RECT  709.925000  2.635000  710.095000 2.805000 ;
      RECT  710.385000 -0.085000  710.555000 0.085000 ;
      RECT  710.385000  2.635000  710.555000 2.805000 ;
      RECT  710.845000 -0.085000  711.015000 0.085000 ;
      RECT  710.845000  2.635000  711.015000 2.805000 ;
      RECT  711.305000 -0.085000  711.475000 0.085000 ;
      RECT  711.305000  2.635000  711.475000 2.805000 ;
      RECT  711.765000 -0.085000  711.935000 0.085000 ;
      RECT  711.765000  2.635000  711.935000 2.805000 ;
      RECT  712.225000 -0.085000  712.395000 0.085000 ;
      RECT  712.225000  2.635000  712.395000 2.805000 ;
      RECT  712.685000 -0.085000  712.855000 0.085000 ;
      RECT  712.685000  2.635000  712.855000 2.805000 ;
      RECT  713.145000 -0.085000  713.315000 0.085000 ;
      RECT  713.145000  2.635000  713.315000 2.805000 ;
      RECT  713.605000 -0.085000  713.775000 0.085000 ;
      RECT  713.605000  2.635000  713.775000 2.805000 ;
      RECT  714.065000 -0.085000  714.235000 0.085000 ;
      RECT  714.065000  2.635000  714.235000 2.805000 ;
      RECT  714.525000 -0.085000  714.695000 0.085000 ;
      RECT  714.525000  2.635000  714.695000 2.805000 ;
      RECT  714.985000 -0.085000  715.155000 0.085000 ;
      RECT  714.985000  2.635000  715.155000 2.805000 ;
      RECT  715.445000 -0.085000  715.615000 0.085000 ;
      RECT  715.445000  2.635000  715.615000 2.805000 ;
      RECT  715.905000 -0.085000  716.075000 0.085000 ;
      RECT  715.905000  2.635000  716.075000 2.805000 ;
      RECT  716.365000 -0.085000  716.535000 0.085000 ;
      RECT  716.365000  2.635000  716.535000 2.805000 ;
      RECT  716.825000 -0.085000  716.995000 0.085000 ;
      RECT  716.825000  2.635000  716.995000 2.805000 ;
      RECT  717.285000 -0.085000  717.455000 0.085000 ;
      RECT  717.285000  2.635000  717.455000 2.805000 ;
      RECT  717.745000 -0.085000  717.915000 0.085000 ;
      RECT  717.745000  2.635000  717.915000 2.805000 ;
      RECT  718.205000 -0.085000  718.375000 0.085000 ;
      RECT  718.205000  2.635000  718.375000 2.805000 ;
      RECT  718.665000 -0.085000  718.835000 0.085000 ;
      RECT  718.665000  2.635000  718.835000 2.805000 ;
      RECT  719.125000 -0.085000  719.295000 0.085000 ;
      RECT  719.125000  2.635000  719.295000 2.805000 ;
      RECT  719.585000 -0.085000  719.755000 0.085000 ;
      RECT  719.585000  2.635000  719.755000 2.805000 ;
      RECT  720.045000 -0.085000  720.215000 0.085000 ;
      RECT  720.045000  2.635000  720.215000 2.805000 ;
      RECT  720.505000 -0.085000  720.675000 0.085000 ;
      RECT  720.505000  2.635000  720.675000 2.805000 ;
      RECT  720.965000 -0.085000  721.135000 0.085000 ;
      RECT  720.965000  2.635000  721.135000 2.805000 ;
      RECT  721.425000 -0.085000  721.595000 0.085000 ;
      RECT  721.425000  2.635000  721.595000 2.805000 ;
      RECT  721.885000 -0.085000  722.055000 0.085000 ;
      RECT  721.885000  2.635000  722.055000 2.805000 ;
      RECT  722.345000 -0.085000  722.515000 0.085000 ;
      RECT  722.345000  2.635000  722.515000 2.805000 ;
      RECT  722.805000 -0.085000  722.975000 0.085000 ;
      RECT  722.805000  2.635000  722.975000 2.805000 ;
      RECT  723.265000 -0.085000  723.435000 0.085000 ;
      RECT  723.265000  2.635000  723.435000 2.805000 ;
      RECT  723.725000 -0.085000  723.895000 0.085000 ;
      RECT  723.725000  2.635000  723.895000 2.805000 ;
      RECT  724.185000 -0.085000  724.355000 0.085000 ;
      RECT  724.185000  2.635000  724.355000 2.805000 ;
      RECT  724.645000 -0.085000  724.815000 0.085000 ;
      RECT  724.645000  2.635000  724.815000 2.805000 ;
      RECT  725.105000 -0.085000  725.275000 0.085000 ;
      RECT  725.105000  2.635000  725.275000 2.805000 ;
      RECT  725.565000 -0.085000  725.735000 0.085000 ;
      RECT  725.565000  2.635000  725.735000 2.805000 ;
      RECT  726.025000 -0.085000  726.195000 0.085000 ;
      RECT  726.025000  2.635000  726.195000 2.805000 ;
      RECT  726.485000 -0.085000  726.655000 0.085000 ;
      RECT  726.485000  2.635000  726.655000 2.805000 ;
      RECT  726.945000 -0.085000  727.115000 0.085000 ;
      RECT  726.945000  2.635000  727.115000 2.805000 ;
      RECT  727.405000 -0.085000  727.575000 0.085000 ;
      RECT  727.405000  2.635000  727.575000 2.805000 ;
      RECT  727.865000 -0.085000  728.035000 0.085000 ;
      RECT  727.865000  2.635000  728.035000 2.805000 ;
      RECT  728.325000 -0.085000  728.495000 0.085000 ;
      RECT  728.325000  2.635000  728.495000 2.805000 ;
      RECT  728.785000 -0.085000  728.955000 0.085000 ;
      RECT  728.785000  2.635000  728.955000 2.805000 ;
      RECT  729.245000 -0.085000  729.415000 0.085000 ;
      RECT  729.245000  2.635000  729.415000 2.805000 ;
      RECT  729.705000 -0.085000  729.875000 0.085000 ;
      RECT  729.705000  2.635000  729.875000 2.805000 ;
      RECT  730.165000 -0.085000  730.335000 0.085000 ;
      RECT  730.165000  2.635000  730.335000 2.805000 ;
      RECT  730.625000 -0.085000  730.795000 0.085000 ;
      RECT  730.625000  2.635000  730.795000 2.805000 ;
      RECT  731.085000 -0.085000  731.255000 0.085000 ;
      RECT  731.085000  2.635000  731.255000 2.805000 ;
      RECT  731.545000 -0.085000  731.715000 0.085000 ;
      RECT  731.545000  2.635000  731.715000 2.805000 ;
      RECT  732.005000 -0.085000  732.175000 0.085000 ;
      RECT  732.005000  2.635000  732.175000 2.805000 ;
      RECT  732.465000 -0.085000  732.635000 0.085000 ;
      RECT  732.465000  2.635000  732.635000 2.805000 ;
      RECT  732.925000 -0.085000  733.095000 0.085000 ;
      RECT  732.925000  2.635000  733.095000 2.805000 ;
      RECT  733.385000 -0.085000  733.555000 0.085000 ;
      RECT  733.385000  2.635000  733.555000 2.805000 ;
      RECT  733.845000 -0.085000  734.015000 0.085000 ;
      RECT  733.845000  2.635000  734.015000 2.805000 ;
      RECT  734.250000  1.105000  734.420000 1.275000 ;
      RECT  734.305000 -0.085000  734.475000 0.085000 ;
      RECT  734.305000  2.635000  734.475000 2.805000 ;
      RECT  734.730000  0.765000  734.900000 0.935000 ;
      RECT  734.765000 -0.085000  734.935000 0.085000 ;
      RECT  734.765000  2.635000  734.935000 2.805000 ;
      RECT  735.225000 -0.085000  735.395000 0.085000 ;
      RECT  735.225000  2.635000  735.395000 2.805000 ;
      RECT  735.685000 -0.085000  735.855000 0.085000 ;
      RECT  735.685000  2.635000  735.855000 2.805000 ;
      RECT  735.730000  1.445000  735.900000 1.615000 ;
      RECT  736.145000 -0.085000  736.315000 0.085000 ;
      RECT  736.145000  2.635000  736.315000 2.805000 ;
      RECT  736.605000 -0.085000  736.775000 0.085000 ;
      RECT  736.605000  2.635000  736.775000 2.805000 ;
      RECT  737.065000 -0.085000  737.235000 0.085000 ;
      RECT  737.065000  2.635000  737.235000 2.805000 ;
      RECT  737.525000 -0.085000  737.695000 0.085000 ;
      RECT  737.525000  2.635000  737.695000 2.805000 ;
      RECT  737.710000  0.765000  737.880000 0.935000 ;
      RECT  737.985000 -0.085000  738.155000 0.085000 ;
      RECT  737.985000  2.635000  738.155000 2.805000 ;
      RECT  738.445000 -0.085000  738.615000 0.085000 ;
      RECT  738.445000  1.105000  738.615000 1.275000 ;
      RECT  738.445000  2.635000  738.615000 2.805000 ;
      RECT  738.905000 -0.085000  739.075000 0.085000 ;
      RECT  738.905000  2.635000  739.075000 2.805000 ;
      RECT  739.365000 -0.085000  739.535000 0.085000 ;
      RECT  739.365000  1.445000  739.535000 1.615000 ;
      RECT  739.365000  2.635000  739.535000 2.805000 ;
      RECT  739.825000 -0.085000  739.995000 0.085000 ;
      RECT  739.825000  2.635000  739.995000 2.805000 ;
      RECT  740.285000 -0.085000  740.455000 0.085000 ;
      RECT  740.285000  2.635000  740.455000 2.805000 ;
      RECT  740.745000 -0.085000  740.915000 0.085000 ;
      RECT  740.745000  2.635000  740.915000 2.805000 ;
      RECT  741.205000 -0.085000  741.375000 0.085000 ;
      RECT  741.205000  2.635000  741.375000 2.805000 ;
      RECT  741.665000 -0.085000  741.835000 0.085000 ;
      RECT  741.665000  2.635000  741.835000 2.805000 ;
      RECT  742.125000 -0.085000  742.295000 0.085000 ;
      RECT  742.125000  2.635000  742.295000 2.805000 ;
      RECT  742.585000 -0.085000  742.755000 0.085000 ;
      RECT  742.585000  2.635000  742.755000 2.805000 ;
      RECT  743.045000 -0.085000  743.215000 0.085000 ;
      RECT  743.045000  2.635000  743.215000 2.805000 ;
      RECT  743.505000 -0.085000  743.675000 0.085000 ;
      RECT  743.505000  2.635000  743.675000 2.805000 ;
      RECT  743.965000 -0.085000  744.135000 0.085000 ;
      RECT  743.965000  2.635000  744.135000 2.805000 ;
      RECT  744.425000 -0.085000  744.595000 0.085000 ;
      RECT  744.425000  2.635000  744.595000 2.805000 ;
      RECT  744.885000 -0.085000  745.055000 0.085000 ;
      RECT  744.885000  2.635000  745.055000 2.805000 ;
      RECT  745.345000 -0.085000  745.515000 0.085000 ;
      RECT  745.345000  2.635000  745.515000 2.805000 ;
      RECT  745.805000 -0.085000  745.975000 0.085000 ;
      RECT  745.805000  2.635000  745.975000 2.805000 ;
      RECT  746.265000 -0.085000  746.435000 0.085000 ;
      RECT  746.265000  2.635000  746.435000 2.805000 ;
      RECT  746.370000  0.765000  746.540000 0.935000 ;
      RECT  746.725000 -0.085000  746.895000 0.085000 ;
      RECT  746.725000  2.635000  746.895000 2.805000 ;
      RECT  747.185000 -0.085000  747.355000 0.085000 ;
      RECT  747.185000  2.635000  747.355000 2.805000 ;
      RECT  747.645000 -0.085000  747.815000 0.085000 ;
      RECT  747.645000  2.635000  747.815000 2.805000 ;
      RECT  748.105000 -0.085000  748.275000 0.085000 ;
      RECT  748.105000  2.635000  748.275000 2.805000 ;
      RECT  748.565000 -0.085000  748.735000 0.085000 ;
      RECT  748.565000  2.635000  748.735000 2.805000 ;
      RECT  749.025000 -0.085000  749.195000 0.085000 ;
      RECT  749.025000  2.635000  749.195000 2.805000 ;
      RECT  749.400000  0.765000  749.570000 0.935000 ;
      RECT  749.485000 -0.085000  749.655000 0.085000 ;
      RECT  749.485000  2.635000  749.655000 2.805000 ;
      RECT  749.945000 -0.085000  750.115000 0.085000 ;
      RECT  749.945000  2.635000  750.115000 2.805000 ;
      RECT  750.405000 -0.085000  750.575000 0.085000 ;
      RECT  750.405000  2.635000  750.575000 2.805000 ;
      RECT  750.865000 -0.085000  751.035000 0.085000 ;
      RECT  750.865000  2.635000  751.035000 2.805000 ;
      RECT  751.325000 -0.085000  751.495000 0.085000 ;
      RECT  751.325000  2.635000  751.495000 2.805000 ;
      RECT  751.785000 -0.085000  751.955000 0.085000 ;
      RECT  751.785000  2.635000  751.955000 2.805000 ;
      RECT  752.245000 -0.085000  752.415000 0.085000 ;
      RECT  752.245000  2.635000  752.415000 2.805000 ;
      RECT  752.705000 -0.085000  752.875000 0.085000 ;
      RECT  752.705000  2.635000  752.875000 2.805000 ;
      RECT  752.860000  0.765000  753.030000 0.935000 ;
      RECT  753.165000 -0.085000  753.335000 0.085000 ;
      RECT  753.165000  2.635000  753.335000 2.805000 ;
      RECT  753.625000 -0.085000  753.795000 0.085000 ;
      RECT  753.625000  2.635000  753.795000 2.805000 ;
      RECT  754.085000 -0.085000  754.255000 0.085000 ;
      RECT  754.085000  2.635000  754.255000 2.805000 ;
      RECT  754.545000 -0.085000  754.715000 0.085000 ;
      RECT  754.545000  2.635000  754.715000 2.805000 ;
      RECT  755.005000 -0.085000  755.175000 0.085000 ;
      RECT  755.005000  2.635000  755.175000 2.805000 ;
      RECT  755.465000 -0.085000  755.635000 0.085000 ;
      RECT  755.465000  2.635000  755.635000 2.805000 ;
      RECT  755.925000 -0.085000  756.095000 0.085000 ;
      RECT  755.925000  2.635000  756.095000 2.805000 ;
      RECT  756.385000 -0.085000  756.555000 0.085000 ;
      RECT  756.385000  2.635000  756.555000 2.805000 ;
      RECT  756.845000 -0.085000  757.015000 0.085000 ;
      RECT  756.845000  2.635000  757.015000 2.805000 ;
      RECT  757.305000 -0.085000  757.475000 0.085000 ;
      RECT  757.305000  2.635000  757.475000 2.805000 ;
      RECT  757.765000 -0.085000  757.935000 0.085000 ;
      RECT  757.765000  2.635000  757.935000 2.805000 ;
      RECT  757.980000  0.765000  758.150000 0.935000 ;
      RECT  758.225000 -0.085000  758.395000 0.085000 ;
      RECT  758.225000  2.635000  758.395000 2.805000 ;
      RECT  758.685000 -0.085000  758.855000 0.085000 ;
      RECT  758.685000  2.635000  758.855000 2.805000 ;
      RECT  759.145000 -0.085000  759.315000 0.085000 ;
      RECT  759.145000  2.635000  759.315000 2.805000 ;
      RECT  759.605000 -0.085000  759.775000 0.085000 ;
      RECT  759.605000  2.635000  759.775000 2.805000 ;
      RECT  760.065000 -0.085000  760.235000 0.085000 ;
      RECT  760.065000  2.635000  760.235000 2.805000 ;
      RECT  760.525000 -0.085000  760.695000 0.085000 ;
      RECT  760.525000  2.635000  760.695000 2.805000 ;
      RECT  760.985000 -0.085000  761.155000 0.085000 ;
      RECT  760.985000  2.635000  761.155000 2.805000 ;
      RECT  761.445000 -0.085000  761.615000 0.085000 ;
      RECT  761.445000  2.635000  761.615000 2.805000 ;
      RECT  761.905000 -0.085000  762.075000 0.085000 ;
      RECT  761.905000  2.635000  762.075000 2.805000 ;
      RECT  762.365000 -0.085000  762.535000 0.085000 ;
      RECT  762.365000  2.635000  762.535000 2.805000 ;
      RECT  762.825000 -0.085000  762.995000 0.085000 ;
      RECT  762.825000  2.635000  762.995000 2.805000 ;
      RECT  763.285000 -0.085000  763.455000 0.085000 ;
      RECT  763.285000  2.635000  763.455000 2.805000 ;
      RECT  763.745000 -0.085000  763.915000 0.085000 ;
      RECT  763.745000  2.635000  763.915000 2.805000 ;
      RECT  764.205000 -0.085000  764.375000 0.085000 ;
      RECT  764.205000  2.635000  764.375000 2.805000 ;
      RECT  764.665000 -0.085000  764.835000 0.085000 ;
      RECT  764.665000  2.635000  764.835000 2.805000 ;
      RECT  765.125000 -0.085000  765.295000 0.085000 ;
      RECT  765.125000  2.635000  765.295000 2.805000 ;
      RECT  765.585000 -0.085000  765.755000 0.085000 ;
      RECT  765.585000  2.635000  765.755000 2.805000 ;
      RECT  766.045000 -0.085000  766.215000 0.085000 ;
      RECT  766.045000  2.635000  766.215000 2.805000 ;
      RECT  766.505000 -0.085000  766.675000 0.085000 ;
      RECT  766.505000  2.635000  766.675000 2.805000 ;
      RECT  766.965000 -0.085000  767.135000 0.085000 ;
      RECT  766.965000  2.635000  767.135000 2.805000 ;
      RECT  767.425000 -0.085000  767.595000 0.085000 ;
      RECT  767.425000  2.635000  767.595000 2.805000 ;
      RECT  767.885000 -0.085000  768.055000 0.085000 ;
      RECT  767.885000  2.635000  768.055000 2.805000 ;
      RECT  768.345000 -0.085000  768.515000 0.085000 ;
      RECT  768.345000  2.635000  768.515000 2.805000 ;
      RECT  768.805000 -0.085000  768.975000 0.085000 ;
      RECT  768.805000  2.635000  768.975000 2.805000 ;
      RECT  769.265000 -0.085000  769.435000 0.085000 ;
      RECT  769.265000  2.635000  769.435000 2.805000 ;
      RECT  769.725000 -0.085000  769.895000 0.085000 ;
      RECT  769.725000  2.635000  769.895000 2.805000 ;
      RECT  770.185000 -0.085000  770.355000 0.085000 ;
      RECT  770.185000  2.635000  770.355000 2.805000 ;
      RECT  770.645000 -0.085000  770.815000 0.085000 ;
      RECT  770.645000  2.635000  770.815000 2.805000 ;
      RECT  771.105000 -0.085000  771.275000 0.085000 ;
      RECT  771.105000  2.635000  771.275000 2.805000 ;
      RECT  771.565000 -0.085000  771.735000 0.085000 ;
      RECT  771.565000  2.635000  771.735000 2.805000 ;
      RECT  772.025000 -0.085000  772.195000 0.085000 ;
      RECT  772.025000  2.635000  772.195000 2.805000 ;
      RECT  772.485000 -0.085000  772.655000 0.085000 ;
      RECT  772.485000  2.635000  772.655000 2.805000 ;
      RECT  772.945000 -0.085000  773.115000 0.085000 ;
      RECT  772.945000  2.635000  773.115000 2.805000 ;
      RECT  773.405000 -0.085000  773.575000 0.085000 ;
      RECT  773.405000  2.635000  773.575000 2.805000 ;
      RECT  773.865000 -0.085000  774.035000 0.085000 ;
      RECT  773.865000  2.635000  774.035000 2.805000 ;
      RECT  774.325000 -0.085000  774.495000 0.085000 ;
      RECT  774.325000  2.635000  774.495000 2.805000 ;
      RECT  774.785000 -0.085000  774.955000 0.085000 ;
      RECT  774.785000  2.635000  774.955000 2.805000 ;
      RECT  775.245000 -0.085000  775.415000 0.085000 ;
      RECT  775.245000  2.635000  775.415000 2.805000 ;
      RECT  775.705000 -0.085000  775.875000 0.085000 ;
      RECT  775.705000  2.635000  775.875000 2.805000 ;
      RECT  776.165000 -0.085000  776.335000 0.085000 ;
      RECT  776.165000  2.635000  776.335000 2.805000 ;
      RECT  776.625000 -0.085000  776.795000 0.085000 ;
      RECT  776.625000  2.635000  776.795000 2.805000 ;
      RECT  777.085000 -0.085000  777.255000 0.085000 ;
      RECT  777.085000  2.635000  777.255000 2.805000 ;
      RECT  777.545000 -0.085000  777.715000 0.085000 ;
      RECT  777.545000  2.635000  777.715000 2.805000 ;
      RECT  778.005000 -0.085000  778.175000 0.085000 ;
      RECT  778.005000  2.635000  778.175000 2.805000 ;
      RECT  778.465000 -0.085000  778.635000 0.085000 ;
      RECT  778.465000  2.635000  778.635000 2.805000 ;
      RECT  778.925000 -0.085000  779.095000 0.085000 ;
      RECT  778.925000  2.635000  779.095000 2.805000 ;
      RECT  779.385000 -0.085000  779.555000 0.085000 ;
      RECT  779.385000  2.635000  779.555000 2.805000 ;
      RECT  779.845000 -0.085000  780.015000 0.085000 ;
      RECT  779.845000  2.635000  780.015000 2.805000 ;
      RECT  780.305000 -0.085000  780.475000 0.085000 ;
      RECT  780.305000  2.635000  780.475000 2.805000 ;
      RECT  780.765000 -0.085000  780.935000 0.085000 ;
      RECT  780.765000  2.635000  780.935000 2.805000 ;
      RECT  781.225000 -0.085000  781.395000 0.085000 ;
      RECT  781.225000  2.635000  781.395000 2.805000 ;
      RECT  781.685000 -0.085000  781.855000 0.085000 ;
      RECT  781.685000  2.635000  781.855000 2.805000 ;
      RECT  782.145000 -0.085000  782.315000 0.085000 ;
      RECT  782.145000  2.635000  782.315000 2.805000 ;
      RECT  782.605000 -0.085000  782.775000 0.085000 ;
      RECT  782.605000  2.635000  782.775000 2.805000 ;
      RECT  783.065000 -0.085000  783.235000 0.085000 ;
      RECT  783.065000  2.635000  783.235000 2.805000 ;
      RECT  783.525000 -0.085000  783.695000 0.085000 ;
      RECT  783.525000  2.635000  783.695000 2.805000 ;
      RECT  783.985000 -0.085000  784.155000 0.085000 ;
      RECT  783.985000  2.635000  784.155000 2.805000 ;
      RECT  784.445000 -0.085000  784.615000 0.085000 ;
      RECT  784.445000  2.635000  784.615000 2.805000 ;
      RECT  784.905000 -0.085000  785.075000 0.085000 ;
      RECT  784.905000  2.635000  785.075000 2.805000 ;
      RECT  785.365000 -0.085000  785.535000 0.085000 ;
      RECT  785.365000  2.635000  785.535000 2.805000 ;
      RECT  785.825000 -0.085000  785.995000 0.085000 ;
      RECT  785.825000  2.635000  785.995000 2.805000 ;
      RECT  786.285000 -0.085000  786.455000 0.085000 ;
      RECT  786.285000  2.635000  786.455000 2.805000 ;
      RECT  786.745000 -0.085000  786.915000 0.085000 ;
      RECT  786.745000  2.635000  786.915000 2.805000 ;
      RECT  787.205000 -0.085000  787.375000 0.085000 ;
      RECT  787.205000  2.635000  787.375000 2.805000 ;
      RECT  787.665000 -0.085000  787.835000 0.085000 ;
      RECT  787.665000  2.635000  787.835000 2.805000 ;
      RECT  788.125000 -0.085000  788.295000 0.085000 ;
      RECT  788.125000  2.635000  788.295000 2.805000 ;
      RECT  788.585000 -0.085000  788.755000 0.085000 ;
      RECT  788.585000  2.635000  788.755000 2.805000 ;
      RECT  789.045000 -0.085000  789.215000 0.085000 ;
      RECT  789.045000  2.635000  789.215000 2.805000 ;
      RECT  789.505000 -0.085000  789.675000 0.085000 ;
      RECT  789.505000  2.635000  789.675000 2.805000 ;
      RECT  789.965000 -0.085000  790.135000 0.085000 ;
      RECT  789.965000  2.635000  790.135000 2.805000 ;
      RECT  790.425000 -0.085000  790.595000 0.085000 ;
      RECT  790.425000  2.635000  790.595000 2.805000 ;
      RECT  790.885000 -0.085000  791.055000 0.085000 ;
      RECT  790.885000  2.635000  791.055000 2.805000 ;
      RECT  791.345000 -0.085000  791.515000 0.085000 ;
      RECT  791.345000  2.635000  791.515000 2.805000 ;
      RECT  791.805000 -0.085000  791.975000 0.085000 ;
      RECT  791.805000  2.635000  791.975000 2.805000 ;
      RECT  792.265000 -0.085000  792.435000 0.085000 ;
      RECT  792.265000  2.635000  792.435000 2.805000 ;
      RECT  792.725000 -0.085000  792.895000 0.085000 ;
      RECT  792.725000  2.635000  792.895000 2.805000 ;
      RECT  793.185000 -0.085000  793.355000 0.085000 ;
      RECT  793.185000  2.635000  793.355000 2.805000 ;
      RECT  793.645000 -0.085000  793.815000 0.085000 ;
      RECT  793.645000  2.635000  793.815000 2.805000 ;
      RECT  794.105000 -0.085000  794.275000 0.085000 ;
      RECT  794.105000  2.635000  794.275000 2.805000 ;
      RECT  794.565000 -0.085000  794.735000 0.085000 ;
      RECT  794.565000  2.635000  794.735000 2.805000 ;
      RECT  795.025000 -0.085000  795.195000 0.085000 ;
      RECT  795.025000  2.635000  795.195000 2.805000 ;
      RECT  795.485000 -0.085000  795.655000 0.085000 ;
      RECT  795.485000  2.635000  795.655000 2.805000 ;
      RECT  795.945000 -0.085000  796.115000 0.085000 ;
      RECT  795.945000  2.635000  796.115000 2.805000 ;
      RECT  796.405000 -0.085000  796.575000 0.085000 ;
      RECT  796.405000  2.635000  796.575000 2.805000 ;
      RECT  796.865000 -0.085000  797.035000 0.085000 ;
      RECT  796.865000  2.635000  797.035000 2.805000 ;
      RECT  797.325000 -0.085000  797.495000 0.085000 ;
      RECT  797.325000  2.635000  797.495000 2.805000 ;
      RECT  797.785000 -0.085000  797.955000 0.085000 ;
      RECT  797.785000  2.635000  797.955000 2.805000 ;
      RECT  798.245000 -0.085000  798.415000 0.085000 ;
      RECT  798.245000  2.635000  798.415000 2.805000 ;
      RECT  798.705000 -0.085000  798.875000 0.085000 ;
      RECT  798.705000  2.635000  798.875000 2.805000 ;
      RECT  799.165000 -0.085000  799.335000 0.085000 ;
      RECT  799.165000  2.635000  799.335000 2.805000 ;
      RECT  799.625000 -0.085000  799.795000 0.085000 ;
      RECT  799.625000  2.635000  799.795000 2.805000 ;
      RECT  800.085000 -0.085000  800.255000 0.085000 ;
      RECT  800.085000  2.635000  800.255000 2.805000 ;
      RECT  800.545000 -0.085000  800.715000 0.085000 ;
      RECT  800.545000  2.635000  800.715000 2.805000 ;
      RECT  801.005000 -0.085000  801.175000 0.085000 ;
      RECT  801.005000  2.635000  801.175000 2.805000 ;
      RECT  801.465000 -0.085000  801.635000 0.085000 ;
      RECT  801.465000  2.635000  801.635000 2.805000 ;
      RECT  801.925000 -0.085000  802.095000 0.085000 ;
      RECT  801.925000  2.635000  802.095000 2.805000 ;
      RECT  802.385000 -0.085000  802.555000 0.085000 ;
      RECT  802.385000  2.635000  802.555000 2.805000 ;
      RECT  802.845000 -0.085000  803.015000 0.085000 ;
      RECT  802.845000  2.635000  803.015000 2.805000 ;
      RECT  803.305000 -0.085000  803.475000 0.085000 ;
      RECT  803.305000  2.635000  803.475000 2.805000 ;
      RECT  803.765000 -0.085000  803.935000 0.085000 ;
      RECT  803.765000  2.635000  803.935000 2.805000 ;
      RECT  804.225000 -0.085000  804.395000 0.085000 ;
      RECT  804.225000  2.635000  804.395000 2.805000 ;
      RECT  804.685000 -0.085000  804.855000 0.085000 ;
      RECT  804.685000  2.635000  804.855000 2.805000 ;
      RECT  805.145000 -0.085000  805.315000 0.085000 ;
      RECT  805.145000  2.635000  805.315000 2.805000 ;
      RECT  805.605000 -0.085000  805.775000 0.085000 ;
      RECT  805.605000  2.635000  805.775000 2.805000 ;
      RECT  806.065000 -0.085000  806.235000 0.085000 ;
      RECT  806.065000  2.635000  806.235000 2.805000 ;
      RECT  806.525000 -0.085000  806.695000 0.085000 ;
      RECT  806.525000  2.635000  806.695000 2.805000 ;
      RECT  806.985000 -0.085000  807.155000 0.085000 ;
      RECT  806.985000  2.635000  807.155000 2.805000 ;
      RECT  807.445000 -0.085000  807.615000 0.085000 ;
      RECT  807.445000  2.635000  807.615000 2.805000 ;
      RECT  807.905000 -0.085000  808.075000 0.085000 ;
      RECT  807.905000  2.635000  808.075000 2.805000 ;
      RECT  808.365000 -0.085000  808.535000 0.085000 ;
      RECT  808.365000  2.635000  808.535000 2.805000 ;
      RECT  808.825000 -0.085000  808.995000 0.085000 ;
      RECT  808.825000  2.635000  808.995000 2.805000 ;
      RECT  809.285000 -0.085000  809.455000 0.085000 ;
      RECT  809.285000  2.635000  809.455000 2.805000 ;
      RECT  809.745000 -0.085000  809.915000 0.085000 ;
      RECT  809.745000  2.635000  809.915000 2.805000 ;
      RECT  810.205000 -0.085000  810.375000 0.085000 ;
      RECT  810.205000  2.635000  810.375000 2.805000 ;
      RECT  810.665000 -0.085000  810.835000 0.085000 ;
      RECT  810.665000  2.635000  810.835000 2.805000 ;
      RECT  811.125000 -0.085000  811.295000 0.085000 ;
      RECT  811.125000  2.635000  811.295000 2.805000 ;
      RECT  811.585000 -0.085000  811.755000 0.085000 ;
      RECT  811.585000  2.635000  811.755000 2.805000 ;
      RECT  812.045000 -0.085000  812.215000 0.085000 ;
      RECT  812.045000  2.635000  812.215000 2.805000 ;
      RECT  812.505000 -0.085000  812.675000 0.085000 ;
      RECT  812.505000  2.635000  812.675000 2.805000 ;
      RECT  812.965000 -0.085000  813.135000 0.085000 ;
      RECT  812.965000  2.635000  813.135000 2.805000 ;
      RECT  813.425000 -0.085000  813.595000 0.085000 ;
      RECT  813.425000  2.635000  813.595000 2.805000 ;
      RECT  813.885000 -0.085000  814.055000 0.085000 ;
      RECT  813.885000  2.635000  814.055000 2.805000 ;
      RECT  814.345000 -0.085000  814.515000 0.085000 ;
      RECT  814.345000  2.635000  814.515000 2.805000 ;
      RECT  814.805000 -0.085000  814.975000 0.085000 ;
      RECT  814.805000  2.635000  814.975000 2.805000 ;
      RECT  815.265000 -0.085000  815.435000 0.085000 ;
      RECT  815.265000  2.635000  815.435000 2.805000 ;
      RECT  815.725000 -0.085000  815.895000 0.085000 ;
      RECT  815.725000  2.635000  815.895000 2.805000 ;
      RECT  816.185000 -0.085000  816.355000 0.085000 ;
      RECT  816.185000  2.635000  816.355000 2.805000 ;
      RECT  816.645000 -0.085000  816.815000 0.085000 ;
      RECT  816.645000  2.635000  816.815000 2.805000 ;
      RECT  817.105000 -0.085000  817.275000 0.085000 ;
      RECT  817.105000  2.635000  817.275000 2.805000 ;
      RECT  817.565000 -0.085000  817.735000 0.085000 ;
      RECT  817.565000  2.635000  817.735000 2.805000 ;
      RECT  818.025000 -0.085000  818.195000 0.085000 ;
      RECT  818.025000  2.635000  818.195000 2.805000 ;
      RECT  818.485000 -0.085000  818.655000 0.085000 ;
      RECT  818.485000  2.635000  818.655000 2.805000 ;
      RECT  818.945000 -0.085000  819.115000 0.085000 ;
      RECT  818.945000  2.635000  819.115000 2.805000 ;
      RECT  819.405000 -0.085000  819.575000 0.085000 ;
      RECT  819.405000  2.635000  819.575000 2.805000 ;
      RECT  819.865000 -0.085000  820.035000 0.085000 ;
      RECT  819.865000  2.635000  820.035000 2.805000 ;
      RECT  820.325000 -0.085000  820.495000 0.085000 ;
      RECT  820.325000  2.635000  820.495000 2.805000 ;
      RECT  820.785000 -0.085000  820.955000 0.085000 ;
      RECT  820.785000  2.635000  820.955000 2.805000 ;
      RECT  821.245000 -0.085000  821.415000 0.085000 ;
      RECT  821.245000  2.635000  821.415000 2.805000 ;
      RECT  821.705000 -0.085000  821.875000 0.085000 ;
      RECT  821.705000  2.635000  821.875000 2.805000 ;
      RECT  822.165000 -0.085000  822.335000 0.085000 ;
      RECT  822.165000  2.635000  822.335000 2.805000 ;
      RECT  822.625000 -0.085000  822.795000 0.085000 ;
      RECT  822.625000  2.635000  822.795000 2.805000 ;
      RECT  823.085000 -0.085000  823.255000 0.085000 ;
      RECT  823.085000  2.635000  823.255000 2.805000 ;
      RECT  823.545000 -0.085000  823.715000 0.085000 ;
      RECT  823.545000  2.635000  823.715000 2.805000 ;
      RECT  824.005000 -0.085000  824.175000 0.085000 ;
      RECT  824.005000  2.635000  824.175000 2.805000 ;
      RECT  824.465000 -0.085000  824.635000 0.085000 ;
      RECT  824.465000  2.635000  824.635000 2.805000 ;
      RECT  824.925000 -0.085000  825.095000 0.085000 ;
      RECT  824.925000  2.635000  825.095000 2.805000 ;
      RECT  825.385000 -0.085000  825.555000 0.085000 ;
      RECT  825.385000  2.635000  825.555000 2.805000 ;
      RECT  825.845000 -0.085000  826.015000 0.085000 ;
      RECT  825.845000  2.635000  826.015000 2.805000 ;
      RECT  826.305000 -0.085000  826.475000 0.085000 ;
      RECT  826.305000  2.635000  826.475000 2.805000 ;
      RECT  826.765000 -0.085000  826.935000 0.085000 ;
      RECT  826.765000  2.635000  826.935000 2.805000 ;
      RECT  827.225000 -0.085000  827.395000 0.085000 ;
      RECT  827.225000  2.635000  827.395000 2.805000 ;
      RECT  827.685000 -0.085000  827.855000 0.085000 ;
      RECT  827.685000  2.635000  827.855000 2.805000 ;
      RECT  828.145000 -0.085000  828.315000 0.085000 ;
      RECT  828.145000  2.635000  828.315000 2.805000 ;
      RECT  828.605000 -0.085000  828.775000 0.085000 ;
      RECT  828.605000  2.635000  828.775000 2.805000 ;
      RECT  829.065000 -0.085000  829.235000 0.085000 ;
      RECT  829.065000  2.635000  829.235000 2.805000 ;
      RECT  829.525000 -0.085000  829.695000 0.085000 ;
      RECT  829.525000  2.635000  829.695000 2.805000 ;
      RECT  829.985000 -0.085000  830.155000 0.085000 ;
      RECT  829.985000  2.635000  830.155000 2.805000 ;
      RECT  830.445000 -0.085000  830.615000 0.085000 ;
      RECT  830.445000  2.635000  830.615000 2.805000 ;
      RECT  830.905000 -0.085000  831.075000 0.085000 ;
      RECT  830.905000  2.635000  831.075000 2.805000 ;
      RECT  831.365000 -0.085000  831.535000 0.085000 ;
      RECT  831.365000  2.635000  831.535000 2.805000 ;
      RECT  831.825000 -0.085000  831.995000 0.085000 ;
      RECT  831.825000  2.635000  831.995000 2.805000 ;
      RECT  832.285000 -0.085000  832.455000 0.085000 ;
      RECT  832.285000  2.635000  832.455000 2.805000 ;
      RECT  832.745000 -0.085000  832.915000 0.085000 ;
      RECT  832.745000  2.635000  832.915000 2.805000 ;
      RECT  833.205000 -0.085000  833.375000 0.085000 ;
      RECT  833.205000  2.635000  833.375000 2.805000 ;
      RECT  833.665000 -0.085000  833.835000 0.085000 ;
      RECT  833.665000  2.635000  833.835000 2.805000 ;
      RECT  834.125000 -0.085000  834.295000 0.085000 ;
      RECT  834.125000  2.635000  834.295000 2.805000 ;
      RECT  834.585000 -0.085000  834.755000 0.085000 ;
      RECT  834.585000  2.635000  834.755000 2.805000 ;
      RECT  835.045000 -0.085000  835.215000 0.085000 ;
      RECT  835.045000  2.635000  835.215000 2.805000 ;
      RECT  835.505000 -0.085000  835.675000 0.085000 ;
      RECT  835.505000  2.635000  835.675000 2.805000 ;
      RECT  835.965000 -0.085000  836.135000 0.085000 ;
      RECT  835.965000  2.635000  836.135000 2.805000 ;
      RECT  836.425000 -0.085000  836.595000 0.085000 ;
      RECT  836.425000  2.635000  836.595000 2.805000 ;
      RECT  836.885000 -0.085000  837.055000 0.085000 ;
      RECT  836.885000  2.635000  837.055000 2.805000 ;
      RECT  837.345000 -0.085000  837.515000 0.085000 ;
      RECT  837.345000  2.635000  837.515000 2.805000 ;
      RECT  837.805000 -0.085000  837.975000 0.085000 ;
      RECT  837.805000  2.635000  837.975000 2.805000 ;
      RECT  838.265000 -0.085000  838.435000 0.085000 ;
      RECT  838.265000  2.635000  838.435000 2.805000 ;
      RECT  838.725000 -0.085000  838.895000 0.085000 ;
      RECT  838.725000  2.635000  838.895000 2.805000 ;
      RECT  839.185000 -0.085000  839.355000 0.085000 ;
      RECT  839.185000  2.635000  839.355000 2.805000 ;
      RECT  839.645000 -0.085000  839.815000 0.085000 ;
      RECT  839.645000  2.635000  839.815000 2.805000 ;
      RECT  840.105000 -0.085000  840.275000 0.085000 ;
      RECT  840.105000  2.635000  840.275000 2.805000 ;
      RECT  840.565000 -0.085000  840.735000 0.085000 ;
      RECT  840.565000  2.635000  840.735000 2.805000 ;
      RECT  841.025000 -0.085000  841.195000 0.085000 ;
      RECT  841.025000  2.635000  841.195000 2.805000 ;
      RECT  841.485000 -0.085000  841.655000 0.085000 ;
      RECT  841.485000  2.635000  841.655000 2.805000 ;
      RECT  841.945000 -0.085000  842.115000 0.085000 ;
      RECT  841.945000  2.635000  842.115000 2.805000 ;
      RECT  842.405000 -0.085000  842.575000 0.085000 ;
      RECT  842.405000  2.635000  842.575000 2.805000 ;
      RECT  842.865000 -0.085000  843.035000 0.085000 ;
      RECT  842.865000  2.635000  843.035000 2.805000 ;
      RECT  843.325000 -0.085000  843.495000 0.085000 ;
      RECT  843.325000  2.635000  843.495000 2.805000 ;
      RECT  843.785000 -0.085000  843.955000 0.085000 ;
      RECT  843.785000  2.635000  843.955000 2.805000 ;
      RECT  844.245000 -0.085000  844.415000 0.085000 ;
      RECT  844.245000  2.635000  844.415000 2.805000 ;
      RECT  844.705000 -0.085000  844.875000 0.085000 ;
      RECT  844.705000  2.635000  844.875000 2.805000 ;
      RECT  845.165000 -0.085000  845.335000 0.085000 ;
      RECT  845.165000  2.635000  845.335000 2.805000 ;
      RECT  845.625000 -0.085000  845.795000 0.085000 ;
      RECT  845.625000  2.635000  845.795000 2.805000 ;
      RECT  846.085000 -0.085000  846.255000 0.085000 ;
      RECT  846.085000  2.635000  846.255000 2.805000 ;
      RECT  846.545000 -0.085000  846.715000 0.085000 ;
      RECT  846.545000  2.635000  846.715000 2.805000 ;
      RECT  847.005000 -0.085000  847.175000 0.085000 ;
      RECT  847.005000  2.635000  847.175000 2.805000 ;
      RECT  847.465000 -0.085000  847.635000 0.085000 ;
      RECT  847.465000  2.635000  847.635000 2.805000 ;
      RECT  847.925000 -0.085000  848.095000 0.085000 ;
      RECT  847.925000  2.635000  848.095000 2.805000 ;
      RECT  848.385000 -0.085000  848.555000 0.085000 ;
      RECT  848.385000  2.635000  848.555000 2.805000 ;
      RECT  848.845000 -0.085000  849.015000 0.085000 ;
      RECT  848.845000  2.635000  849.015000 2.805000 ;
      RECT  849.305000 -0.085000  849.475000 0.085000 ;
      RECT  849.305000  2.635000  849.475000 2.805000 ;
      RECT  849.765000 -0.085000  849.935000 0.085000 ;
      RECT  849.765000  2.635000  849.935000 2.805000 ;
      RECT  850.225000 -0.085000  850.395000 0.085000 ;
      RECT  850.225000  2.635000  850.395000 2.805000 ;
      RECT  850.685000 -0.085000  850.855000 0.085000 ;
      RECT  850.685000  2.635000  850.855000 2.805000 ;
      RECT  851.145000 -0.085000  851.315000 0.085000 ;
      RECT  851.145000  2.635000  851.315000 2.805000 ;
      RECT  851.605000 -0.085000  851.775000 0.085000 ;
      RECT  851.605000  2.635000  851.775000 2.805000 ;
      RECT  852.065000 -0.085000  852.235000 0.085000 ;
      RECT  852.065000  2.635000  852.235000 2.805000 ;
      RECT  852.525000 -0.085000  852.695000 0.085000 ;
      RECT  852.525000  2.635000  852.695000 2.805000 ;
      RECT  852.985000 -0.085000  853.155000 0.085000 ;
      RECT  852.985000  2.635000  853.155000 2.805000 ;
      RECT  853.445000 -0.085000  853.615000 0.085000 ;
      RECT  853.445000  2.635000  853.615000 2.805000 ;
      RECT  853.905000 -0.085000  854.075000 0.085000 ;
      RECT  853.905000  2.635000  854.075000 2.805000 ;
      RECT  854.365000 -0.085000  854.535000 0.085000 ;
      RECT  854.365000  2.635000  854.535000 2.805000 ;
      RECT  854.825000 -0.085000  854.995000 0.085000 ;
      RECT  854.825000  2.635000  854.995000 2.805000 ;
      RECT  855.285000 -0.085000  855.455000 0.085000 ;
      RECT  855.285000  2.635000  855.455000 2.805000 ;
      RECT  855.745000 -0.085000  855.915000 0.085000 ;
      RECT  855.745000  2.635000  855.915000 2.805000 ;
      RECT  856.205000 -0.085000  856.375000 0.085000 ;
      RECT  856.205000  2.635000  856.375000 2.805000 ;
      RECT  856.665000 -0.085000  856.835000 0.085000 ;
      RECT  856.665000  2.635000  856.835000 2.805000 ;
      RECT  857.125000 -0.085000  857.295000 0.085000 ;
      RECT  857.125000  2.635000  857.295000 2.805000 ;
      RECT  857.585000 -0.085000  857.755000 0.085000 ;
      RECT  857.585000  2.635000  857.755000 2.805000 ;
      RECT  858.045000 -0.085000  858.215000 0.085000 ;
      RECT  858.045000  2.635000  858.215000 2.805000 ;
      RECT  858.505000 -0.085000  858.675000 0.085000 ;
      RECT  858.505000  2.635000  858.675000 2.805000 ;
      RECT  858.965000 -0.085000  859.135000 0.085000 ;
      RECT  858.965000  2.635000  859.135000 2.805000 ;
      RECT  859.425000 -0.085000  859.595000 0.085000 ;
      RECT  859.425000  2.635000  859.595000 2.805000 ;
      RECT  859.885000 -0.085000  860.055000 0.085000 ;
      RECT  859.885000  2.635000  860.055000 2.805000 ;
      RECT  860.345000 -0.085000  860.515000 0.085000 ;
      RECT  860.345000  2.635000  860.515000 2.805000 ;
      RECT  860.805000 -0.085000  860.975000 0.085000 ;
      RECT  860.805000  2.635000  860.975000 2.805000 ;
      RECT  861.265000 -0.085000  861.435000 0.085000 ;
      RECT  861.265000  2.635000  861.435000 2.805000 ;
      RECT  861.725000 -0.085000  861.895000 0.085000 ;
      RECT  861.725000  2.635000  861.895000 2.805000 ;
      RECT  862.185000 -0.085000  862.355000 0.085000 ;
      RECT  862.185000  2.635000  862.355000 2.805000 ;
      RECT  862.645000 -0.085000  862.815000 0.085000 ;
      RECT  862.645000  2.635000  862.815000 2.805000 ;
      RECT  863.105000 -0.085000  863.275000 0.085000 ;
      RECT  863.105000  2.635000  863.275000 2.805000 ;
      RECT  863.565000 -0.085000  863.735000 0.085000 ;
      RECT  863.565000  2.635000  863.735000 2.805000 ;
      RECT  864.025000 -0.085000  864.195000 0.085000 ;
      RECT  864.025000  2.635000  864.195000 2.805000 ;
      RECT  864.485000 -0.085000  864.655000 0.085000 ;
      RECT  864.485000  2.635000  864.655000 2.805000 ;
      RECT  864.945000 -0.085000  865.115000 0.085000 ;
      RECT  864.945000  2.635000  865.115000 2.805000 ;
      RECT  865.405000 -0.085000  865.575000 0.085000 ;
      RECT  865.405000  2.635000  865.575000 2.805000 ;
      RECT  865.865000 -0.085000  866.035000 0.085000 ;
      RECT  865.865000  2.635000  866.035000 2.805000 ;
      RECT  866.325000 -0.085000  866.495000 0.085000 ;
      RECT  866.325000  2.635000  866.495000 2.805000 ;
      RECT  866.785000 -0.085000  866.955000 0.085000 ;
      RECT  866.785000  2.635000  866.955000 2.805000 ;
      RECT  867.245000 -0.085000  867.415000 0.085000 ;
      RECT  867.245000  2.635000  867.415000 2.805000 ;
      RECT  867.705000 -0.085000  867.875000 0.085000 ;
      RECT  867.705000  2.635000  867.875000 2.805000 ;
      RECT  867.800000  1.105000  867.970000 1.275000 ;
      RECT  868.165000 -0.085000  868.335000 0.085000 ;
      RECT  868.165000  2.635000  868.335000 2.805000 ;
      RECT  868.625000 -0.085000  868.795000 0.085000 ;
      RECT  868.625000  2.635000  868.795000 2.805000 ;
      RECT  869.085000 -0.085000  869.255000 0.085000 ;
      RECT  869.085000  2.635000  869.255000 2.805000 ;
      RECT  869.545000 -0.085000  869.715000 0.085000 ;
      RECT  869.545000  2.635000  869.715000 2.805000 ;
      RECT  869.795000  1.105000  869.965000 1.275000 ;
      RECT  870.005000 -0.085000  870.175000 0.085000 ;
      RECT  870.005000  2.635000  870.175000 2.805000 ;
      RECT  870.465000 -0.085000  870.635000 0.085000 ;
      RECT  870.465000  2.635000  870.635000 2.805000 ;
      RECT  870.925000 -0.085000  871.095000 0.085000 ;
      RECT  870.925000  2.635000  871.095000 2.805000 ;
      RECT  871.385000 -0.085000  871.555000 0.085000 ;
      RECT  871.385000  2.635000  871.555000 2.805000 ;
      RECT  871.845000 -0.085000  872.015000 0.085000 ;
      RECT  871.845000  2.635000  872.015000 2.805000 ;
      RECT  872.305000 -0.085000  872.475000 0.085000 ;
      RECT  872.305000  2.635000  872.475000 2.805000 ;
      RECT  872.765000 -0.085000  872.935000 0.085000 ;
      RECT  872.765000  2.635000  872.935000 2.805000 ;
      RECT  873.225000 -0.085000  873.395000 0.085000 ;
      RECT  873.225000  2.635000  873.395000 2.805000 ;
      RECT  873.685000 -0.085000  873.855000 0.085000 ;
      RECT  873.685000  2.635000  873.855000 2.805000 ;
      RECT  874.145000 -0.085000  874.315000 0.085000 ;
      RECT  874.145000  2.635000  874.315000 2.805000 ;
      RECT  874.605000 -0.085000  874.775000 0.085000 ;
      RECT  874.605000  2.635000  874.775000 2.805000 ;
      RECT  875.065000 -0.085000  875.235000 0.085000 ;
      RECT  875.065000  2.635000  875.235000 2.805000 ;
      RECT  875.335000  1.105000  875.505000 1.275000 ;
      RECT  875.525000 -0.085000  875.695000 0.085000 ;
      RECT  875.525000  2.635000  875.695000 2.805000 ;
      RECT  875.985000 -0.085000  876.155000 0.085000 ;
      RECT  875.985000  2.635000  876.155000 2.805000 ;
      RECT  876.445000 -0.085000  876.615000 0.085000 ;
      RECT  876.445000  2.635000  876.615000 2.805000 ;
      RECT  876.905000 -0.085000  877.075000 0.085000 ;
      RECT  876.905000  2.635000  877.075000 2.805000 ;
      RECT  877.365000 -0.085000  877.535000 0.085000 ;
      RECT  877.365000  2.635000  877.535000 2.805000 ;
      RECT  877.825000 -0.085000  877.995000 0.085000 ;
      RECT  877.825000  2.635000  877.995000 2.805000 ;
      RECT  877.870000  1.105000  878.040000 1.275000 ;
      RECT  878.285000 -0.085000  878.455000 0.085000 ;
      RECT  878.285000  2.635000  878.455000 2.805000 ;
      RECT  878.745000 -0.085000  878.915000 0.085000 ;
      RECT  878.745000  2.635000  878.915000 2.805000 ;
      RECT  879.205000 -0.085000  879.375000 0.085000 ;
      RECT  879.205000  2.635000  879.375000 2.805000 ;
      RECT  879.665000 -0.085000  879.835000 0.085000 ;
      RECT  879.665000  2.635000  879.835000 2.805000 ;
      RECT  880.125000 -0.085000  880.295000 0.085000 ;
      RECT  880.125000  2.635000  880.295000 2.805000 ;
      RECT  880.585000 -0.085000  880.755000 0.085000 ;
      RECT  880.585000  2.635000  880.755000 2.805000 ;
      RECT  881.045000 -0.085000  881.215000 0.085000 ;
      RECT  881.045000  2.635000  881.215000 2.805000 ;
      RECT  881.505000 -0.085000  881.675000 0.085000 ;
      RECT  881.505000  2.635000  881.675000 2.805000 ;
      RECT  881.965000 -0.085000  882.135000 0.085000 ;
      RECT  881.965000  2.635000  882.135000 2.805000 ;
      RECT  882.425000 -0.085000  882.595000 0.085000 ;
      RECT  882.425000  2.635000  882.595000 2.805000 ;
      RECT  882.885000 -0.085000  883.055000 0.085000 ;
      RECT  882.885000  2.635000  883.055000 2.805000 ;
      RECT  883.345000 -0.085000  883.515000 0.085000 ;
      RECT  883.345000  2.635000  883.515000 2.805000 ;
      RECT  883.805000 -0.085000  883.975000 0.085000 ;
      RECT  883.805000  2.635000  883.975000 2.805000 ;
      RECT  884.265000 -0.085000  884.435000 0.085000 ;
      RECT  884.265000  2.635000  884.435000 2.805000 ;
      RECT  884.725000 -0.085000  884.895000 0.085000 ;
      RECT  884.725000  2.635000  884.895000 2.805000 ;
      RECT  885.185000 -0.085000  885.355000 0.085000 ;
      RECT  885.185000  2.635000  885.355000 2.805000 ;
      RECT  885.645000 -0.085000  885.815000 0.085000 ;
      RECT  885.645000  2.635000  885.815000 2.805000 ;
      RECT  886.105000 -0.085000  886.275000 0.085000 ;
      RECT  886.105000  2.635000  886.275000 2.805000 ;
      RECT  886.565000 -0.085000  886.735000 0.085000 ;
      RECT  886.565000  2.635000  886.735000 2.805000 ;
      RECT  887.025000 -0.085000  887.195000 0.085000 ;
      RECT  887.025000  2.635000  887.195000 2.805000 ;
      RECT  887.485000 -0.085000  887.655000 0.085000 ;
      RECT  887.485000  2.635000  887.655000 2.805000 ;
      RECT  887.945000 -0.085000  888.115000 0.085000 ;
      RECT  887.945000  2.635000  888.115000 2.805000 ;
      RECT  888.405000 -0.085000  888.575000 0.085000 ;
      RECT  888.405000  2.635000  888.575000 2.805000 ;
      RECT  888.865000 -0.085000  889.035000 0.085000 ;
      RECT  888.865000  2.635000  889.035000 2.805000 ;
      RECT  889.325000 -0.085000  889.495000 0.085000 ;
      RECT  889.325000  2.635000  889.495000 2.805000 ;
      RECT  889.785000 -0.085000  889.955000 0.085000 ;
      RECT  889.785000  2.635000  889.955000 2.805000 ;
      RECT  890.245000 -0.085000  890.415000 0.085000 ;
      RECT  890.245000  2.635000  890.415000 2.805000 ;
      RECT  890.705000 -0.085000  890.875000 0.085000 ;
      RECT  890.705000  2.635000  890.875000 2.805000 ;
      RECT  891.165000 -0.085000  891.335000 0.085000 ;
      RECT  891.165000  2.635000  891.335000 2.805000 ;
      RECT  891.625000 -0.085000  891.795000 0.085000 ;
      RECT  891.625000  2.635000  891.795000 2.805000 ;
      RECT  892.085000 -0.085000  892.255000 0.085000 ;
      RECT  892.085000  2.635000  892.255000 2.805000 ;
      RECT  892.545000 -0.085000  892.715000 0.085000 ;
      RECT  892.545000  2.635000  892.715000 2.805000 ;
      RECT  893.005000 -0.085000  893.175000 0.085000 ;
      RECT  893.005000  2.635000  893.175000 2.805000 ;
      RECT  893.465000 -0.085000  893.635000 0.085000 ;
      RECT  893.465000  2.635000  893.635000 2.805000 ;
      RECT  893.925000 -0.085000  894.095000 0.085000 ;
      RECT  893.925000  2.635000  894.095000 2.805000 ;
      RECT  894.385000 -0.085000  894.555000 0.085000 ;
      RECT  894.385000  2.635000  894.555000 2.805000 ;
      RECT  894.845000 -0.085000  895.015000 0.085000 ;
      RECT  894.845000  2.635000  895.015000 2.805000 ;
      RECT  895.305000 -0.085000  895.475000 0.085000 ;
      RECT  895.305000  2.635000  895.475000 2.805000 ;
      RECT  895.765000 -0.085000  895.935000 0.085000 ;
      RECT  895.765000  2.635000  895.935000 2.805000 ;
      RECT  896.225000 -0.085000  896.395000 0.085000 ;
      RECT  896.225000  2.635000  896.395000 2.805000 ;
      RECT  896.685000 -0.085000  896.855000 0.085000 ;
      RECT  896.685000  2.635000  896.855000 2.805000 ;
      RECT  897.145000 -0.085000  897.315000 0.085000 ;
      RECT  897.145000  2.635000  897.315000 2.805000 ;
      RECT  897.605000 -0.085000  897.775000 0.085000 ;
      RECT  897.605000  2.635000  897.775000 2.805000 ;
      RECT  898.065000 -0.085000  898.235000 0.085000 ;
      RECT  898.065000  2.635000  898.235000 2.805000 ;
      RECT  898.525000 -0.085000  898.695000 0.085000 ;
      RECT  898.525000  2.635000  898.695000 2.805000 ;
      RECT  898.985000 -0.085000  899.155000 0.085000 ;
      RECT  898.985000  2.635000  899.155000 2.805000 ;
      RECT  899.445000 -0.085000  899.615000 0.085000 ;
      RECT  899.445000  2.635000  899.615000 2.805000 ;
      RECT  899.905000 -0.085000  900.075000 0.085000 ;
      RECT  899.905000  2.635000  900.075000 2.805000 ;
      RECT  900.365000 -0.085000  900.535000 0.085000 ;
      RECT  900.365000  2.635000  900.535000 2.805000 ;
      RECT  900.825000 -0.085000  900.995000 0.085000 ;
      RECT  900.825000  2.635000  900.995000 2.805000 ;
      RECT  901.285000 -0.085000  901.455000 0.085000 ;
      RECT  901.285000  2.635000  901.455000 2.805000 ;
      RECT  901.745000 -0.085000  901.915000 0.085000 ;
      RECT  901.745000  2.635000  901.915000 2.805000 ;
      RECT  902.205000 -0.085000  902.375000 0.085000 ;
      RECT  902.205000  2.635000  902.375000 2.805000 ;
      RECT  902.665000 -0.085000  902.835000 0.085000 ;
      RECT  902.665000  2.635000  902.835000 2.805000 ;
      RECT  903.125000 -0.085000  903.295000 0.085000 ;
      RECT  903.125000  2.635000  903.295000 2.805000 ;
      RECT  903.585000 -0.085000  903.755000 0.085000 ;
      RECT  903.585000  2.635000  903.755000 2.805000 ;
      RECT  904.045000 -0.085000  904.215000 0.085000 ;
      RECT  904.045000  2.635000  904.215000 2.805000 ;
      RECT  904.505000 -0.085000  904.675000 0.085000 ;
      RECT  904.505000  2.635000  904.675000 2.805000 ;
      RECT  904.965000 -0.085000  905.135000 0.085000 ;
      RECT  904.965000  2.635000  905.135000 2.805000 ;
      RECT  905.425000 -0.085000  905.595000 0.085000 ;
      RECT  905.425000  2.635000  905.595000 2.805000 ;
      RECT  905.885000 -0.085000  906.055000 0.085000 ;
      RECT  905.885000  2.635000  906.055000 2.805000 ;
      RECT  906.345000 -0.085000  906.515000 0.085000 ;
      RECT  906.345000  2.635000  906.515000 2.805000 ;
      RECT  906.805000 -0.085000  906.975000 0.085000 ;
      RECT  906.805000  2.635000  906.975000 2.805000 ;
      RECT  907.265000 -0.085000  907.435000 0.085000 ;
      RECT  907.265000  2.635000  907.435000 2.805000 ;
      RECT  907.725000 -0.085000  907.895000 0.085000 ;
      RECT  907.725000  2.635000  907.895000 2.805000 ;
      RECT  908.185000 -0.085000  908.355000 0.085000 ;
      RECT  908.185000  2.635000  908.355000 2.805000 ;
      RECT  908.645000 -0.085000  908.815000 0.085000 ;
      RECT  908.645000  2.635000  908.815000 2.805000 ;
      RECT  909.105000 -0.085000  909.275000 0.085000 ;
      RECT  909.105000  2.635000  909.275000 2.805000 ;
      RECT  909.565000 -0.085000  909.735000 0.085000 ;
      RECT  909.565000  2.635000  909.735000 2.805000 ;
      RECT  910.025000 -0.085000  910.195000 0.085000 ;
      RECT  910.025000  2.635000  910.195000 2.805000 ;
      RECT  910.485000 -0.085000  910.655000 0.085000 ;
      RECT  910.485000  2.635000  910.655000 2.805000 ;
      RECT  910.945000 -0.085000  911.115000 0.085000 ;
      RECT  910.945000  2.635000  911.115000 2.805000 ;
      RECT  911.405000 -0.085000  911.575000 0.085000 ;
      RECT  911.405000  2.635000  911.575000 2.805000 ;
      RECT  911.865000 -0.085000  912.035000 0.085000 ;
      RECT  911.865000  2.635000  912.035000 2.805000 ;
      RECT  912.325000 -0.085000  912.495000 0.085000 ;
      RECT  912.325000  2.635000  912.495000 2.805000 ;
      RECT  912.785000 -0.085000  912.955000 0.085000 ;
      RECT  912.785000  2.635000  912.955000 2.805000 ;
      RECT  913.245000 -0.085000  913.415000 0.085000 ;
      RECT  913.245000  2.635000  913.415000 2.805000 ;
      RECT  913.705000 -0.085000  913.875000 0.085000 ;
      RECT  913.705000  2.635000  913.875000 2.805000 ;
      RECT  914.165000 -0.085000  914.335000 0.085000 ;
      RECT  914.165000  2.635000  914.335000 2.805000 ;
      RECT  914.625000 -0.085000  914.795000 0.085000 ;
      RECT  914.625000  2.635000  914.795000 2.805000 ;
      RECT  915.085000 -0.085000  915.255000 0.085000 ;
      RECT  915.085000  2.635000  915.255000 2.805000 ;
      RECT  915.545000 -0.085000  915.715000 0.085000 ;
      RECT  915.545000  2.635000  915.715000 2.805000 ;
      RECT  916.005000 -0.085000  916.175000 0.085000 ;
      RECT  916.005000  2.635000  916.175000 2.805000 ;
      RECT  916.465000 -0.085000  916.635000 0.085000 ;
      RECT  916.465000  2.635000  916.635000 2.805000 ;
      RECT  916.925000 -0.085000  917.095000 0.085000 ;
      RECT  916.925000  2.635000  917.095000 2.805000 ;
      RECT  917.385000 -0.085000  917.555000 0.085000 ;
      RECT  917.385000  2.635000  917.555000 2.805000 ;
      RECT  917.845000 -0.085000  918.015000 0.085000 ;
      RECT  917.845000  2.635000  918.015000 2.805000 ;
      RECT  918.305000 -0.085000  918.475000 0.085000 ;
      RECT  918.305000  2.635000  918.475000 2.805000 ;
      RECT  918.765000 -0.085000  918.935000 0.085000 ;
      RECT  918.765000  2.635000  918.935000 2.805000 ;
      RECT  919.225000 -0.085000  919.395000 0.085000 ;
      RECT  919.225000  2.635000  919.395000 2.805000 ;
      RECT  919.685000 -0.085000  919.855000 0.085000 ;
      RECT  919.685000  2.635000  919.855000 2.805000 ;
      RECT  920.145000 -0.085000  920.315000 0.085000 ;
      RECT  920.145000  2.635000  920.315000 2.805000 ;
      RECT  920.605000 -0.085000  920.775000 0.085000 ;
      RECT  920.605000  2.635000  920.775000 2.805000 ;
      RECT  921.065000 -0.085000  921.235000 0.085000 ;
      RECT  921.065000  2.635000  921.235000 2.805000 ;
      RECT  921.525000 -0.085000  921.695000 0.085000 ;
      RECT  921.525000  2.635000  921.695000 2.805000 ;
      RECT  921.985000 -0.085000  922.155000 0.085000 ;
      RECT  921.985000  2.635000  922.155000 2.805000 ;
      RECT  922.445000 -0.085000  922.615000 0.085000 ;
      RECT  922.445000  2.635000  922.615000 2.805000 ;
      RECT  922.905000 -0.085000  923.075000 0.085000 ;
      RECT  922.905000  2.635000  923.075000 2.805000 ;
      RECT  923.365000 -0.085000  923.535000 0.085000 ;
      RECT  923.365000  2.635000  923.535000 2.805000 ;
      RECT  923.825000 -0.085000  923.995000 0.085000 ;
      RECT  923.825000  2.635000  923.995000 2.805000 ;
      RECT  924.285000 -0.085000  924.455000 0.085000 ;
      RECT  924.285000  2.635000  924.455000 2.805000 ;
      RECT  924.745000 -0.085000  924.915000 0.085000 ;
      RECT  924.745000  2.635000  924.915000 2.805000 ;
      RECT  925.205000 -0.085000  925.375000 0.085000 ;
      RECT  925.205000  2.635000  925.375000 2.805000 ;
      RECT  925.665000 -0.085000  925.835000 0.085000 ;
      RECT  925.665000  2.635000  925.835000 2.805000 ;
      RECT  926.125000 -0.085000  926.295000 0.085000 ;
      RECT  926.125000  2.635000  926.295000 2.805000 ;
      RECT  926.585000 -0.085000  926.755000 0.085000 ;
      RECT  926.585000  2.635000  926.755000 2.805000 ;
      RECT  926.835000  2.125000  927.005000 2.295000 ;
      RECT  927.045000 -0.085000  927.215000 0.085000 ;
      RECT  927.045000  2.635000  927.215000 2.805000 ;
      RECT  927.505000 -0.085000  927.675000 0.085000 ;
      RECT  927.505000  2.635000  927.675000 2.805000 ;
      RECT  927.965000 -0.085000  928.135000 0.085000 ;
      RECT  927.965000  2.635000  928.135000 2.805000 ;
      RECT  928.425000 -0.085000  928.595000 0.085000 ;
      RECT  928.425000  2.635000  928.595000 2.805000 ;
      RECT  928.885000 -0.085000  929.055000 0.085000 ;
      RECT  928.885000  2.635000  929.055000 2.805000 ;
      RECT  929.345000 -0.085000  929.515000 0.085000 ;
      RECT  929.345000  2.635000  929.515000 2.805000 ;
      RECT  929.805000 -0.085000  929.975000 0.085000 ;
      RECT  929.805000  2.635000  929.975000 2.805000 ;
      RECT  929.945000  2.125000  930.115000 2.295000 ;
      RECT  930.265000 -0.085000  930.435000 0.085000 ;
      RECT  930.265000  2.635000  930.435000 2.805000 ;
      RECT  930.725000 -0.085000  930.895000 0.085000 ;
      RECT  930.725000  2.635000  930.895000 2.805000 ;
      RECT  931.185000 -0.085000  931.355000 0.085000 ;
      RECT  931.185000  2.635000  931.355000 2.805000 ;
      RECT  931.645000 -0.085000  931.815000 0.085000 ;
      RECT  931.645000  2.635000  931.815000 2.805000 ;
      RECT  932.105000 -0.085000  932.275000 0.085000 ;
      RECT  932.105000  2.635000  932.275000 2.805000 ;
      RECT  932.565000 -0.085000  932.735000 0.085000 ;
      RECT  932.565000  2.635000  932.735000 2.805000 ;
      RECT  933.025000 -0.085000  933.195000 0.085000 ;
      RECT  933.025000  2.635000  933.195000 2.805000 ;
      RECT  933.485000 -0.085000  933.655000 0.085000 ;
      RECT  933.485000  2.635000  933.655000 2.805000 ;
      RECT  933.945000 -0.085000  934.115000 0.085000 ;
      RECT  933.945000  2.635000  934.115000 2.805000 ;
      RECT  934.405000 -0.085000  934.575000 0.085000 ;
      RECT  934.405000  2.635000  934.575000 2.805000 ;
      RECT  934.865000 -0.085000  935.035000 0.085000 ;
      RECT  934.865000  2.635000  935.035000 2.805000 ;
      RECT  935.325000 -0.085000  935.495000 0.085000 ;
      RECT  935.325000  2.635000  935.495000 2.805000 ;
      RECT  935.785000 -0.085000  935.955000 0.085000 ;
      RECT  935.785000  2.635000  935.955000 2.805000 ;
      RECT  936.245000 -0.085000  936.415000 0.085000 ;
      RECT  936.245000  2.635000  936.415000 2.805000 ;
      RECT  936.705000 -0.085000  936.875000 0.085000 ;
      RECT  936.705000  2.635000  936.875000 2.805000 ;
      RECT  937.165000 -0.085000  937.335000 0.085000 ;
      RECT  937.165000  2.635000  937.335000 2.805000 ;
      RECT  937.625000 -0.085000  937.795000 0.085000 ;
      RECT  937.625000  2.635000  937.795000 2.805000 ;
      RECT  938.085000 -0.085000  938.255000 0.085000 ;
      RECT  938.085000  2.635000  938.255000 2.805000 ;
      RECT  938.545000 -0.085000  938.715000 0.085000 ;
      RECT  938.545000  2.635000  938.715000 2.805000 ;
      RECT  939.005000 -0.085000  939.175000 0.085000 ;
      RECT  939.005000  2.635000  939.175000 2.805000 ;
      RECT  939.465000 -0.085000  939.635000 0.085000 ;
      RECT  939.465000  2.635000  939.635000 2.805000 ;
      RECT  939.925000 -0.085000  940.095000 0.085000 ;
      RECT  939.925000  2.635000  940.095000 2.805000 ;
      RECT  940.385000 -0.085000  940.555000 0.085000 ;
      RECT  940.385000  2.635000  940.555000 2.805000 ;
      RECT  940.845000 -0.085000  941.015000 0.085000 ;
      RECT  940.845000  2.635000  941.015000 2.805000 ;
      RECT  941.305000 -0.085000  941.475000 0.085000 ;
      RECT  941.305000  2.635000  941.475000 2.805000 ;
      RECT  941.765000 -0.085000  941.935000 0.085000 ;
      RECT  941.765000  2.635000  941.935000 2.805000 ;
      RECT  942.225000 -0.085000  942.395000 0.085000 ;
      RECT  942.225000  2.635000  942.395000 2.805000 ;
      RECT  942.685000 -0.085000  942.855000 0.085000 ;
      RECT  942.685000  2.635000  942.855000 2.805000 ;
      RECT  943.145000 -0.085000  943.315000 0.085000 ;
      RECT  943.145000  2.635000  943.315000 2.805000 ;
      RECT  943.605000 -0.085000  943.775000 0.085000 ;
      RECT  943.605000  2.635000  943.775000 2.805000 ;
      RECT  944.065000 -0.085000  944.235000 0.085000 ;
      RECT  944.065000  2.635000  944.235000 2.805000 ;
      RECT  944.525000 -0.085000  944.695000 0.085000 ;
      RECT  944.525000  2.635000  944.695000 2.805000 ;
      RECT  944.985000 -0.085000  945.155000 0.085000 ;
      RECT  944.985000  2.635000  945.155000 2.805000 ;
      RECT  945.445000 -0.085000  945.615000 0.085000 ;
      RECT  945.445000  2.635000  945.615000 2.805000 ;
      RECT  945.905000 -0.085000  946.075000 0.085000 ;
      RECT  945.905000  2.635000  946.075000 2.805000 ;
      RECT  946.365000 -0.085000  946.535000 0.085000 ;
      RECT  946.365000  2.635000  946.535000 2.805000 ;
      RECT  946.825000 -0.085000  946.995000 0.085000 ;
      RECT  946.825000  2.635000  946.995000 2.805000 ;
      RECT  947.285000 -0.085000  947.455000 0.085000 ;
      RECT  947.285000  2.635000  947.455000 2.805000 ;
      RECT  947.745000 -0.085000  947.915000 0.085000 ;
      RECT  947.745000  2.635000  947.915000 2.805000 ;
      RECT  948.205000 -0.085000  948.375000 0.085000 ;
      RECT  948.205000  2.635000  948.375000 2.805000 ;
      RECT  948.665000 -0.085000  948.835000 0.085000 ;
      RECT  948.665000  2.635000  948.835000 2.805000 ;
      RECT  949.125000 -0.085000  949.295000 0.085000 ;
      RECT  949.125000  2.635000  949.295000 2.805000 ;
      RECT  949.585000 -0.085000  949.755000 0.085000 ;
      RECT  949.585000  2.635000  949.755000 2.805000 ;
      RECT  950.045000 -0.085000  950.215000 0.085000 ;
      RECT  950.045000  2.635000  950.215000 2.805000 ;
      RECT  950.505000 -0.085000  950.675000 0.085000 ;
      RECT  950.505000  2.635000  950.675000 2.805000 ;
      RECT  950.965000 -0.085000  951.135000 0.085000 ;
      RECT  950.965000  2.635000  951.135000 2.805000 ;
      RECT  951.425000 -0.085000  951.595000 0.085000 ;
      RECT  951.425000  2.635000  951.595000 2.805000 ;
      RECT  951.885000 -0.085000  952.055000 0.085000 ;
      RECT  951.885000  2.635000  952.055000 2.805000 ;
      RECT  952.345000 -0.085000  952.515000 0.085000 ;
      RECT  952.345000  2.635000  952.515000 2.805000 ;
      RECT  952.805000 -0.085000  952.975000 0.085000 ;
      RECT  952.805000  2.635000  952.975000 2.805000 ;
      RECT  953.265000 -0.085000  953.435000 0.085000 ;
      RECT  953.265000  2.635000  953.435000 2.805000 ;
      RECT  953.725000 -0.085000  953.895000 0.085000 ;
      RECT  953.725000  2.635000  953.895000 2.805000 ;
      RECT  954.185000 -0.085000  954.355000 0.085000 ;
      RECT  954.185000  2.635000  954.355000 2.805000 ;
      RECT  954.645000 -0.085000  954.815000 0.085000 ;
      RECT  954.645000  2.635000  954.815000 2.805000 ;
      RECT  955.105000 -0.085000  955.275000 0.085000 ;
      RECT  955.105000  2.635000  955.275000 2.805000 ;
      RECT  955.565000 -0.085000  955.735000 0.085000 ;
      RECT  955.565000  2.635000  955.735000 2.805000 ;
      RECT  956.025000 -0.085000  956.195000 0.085000 ;
      RECT  956.025000  2.635000  956.195000 2.805000 ;
      RECT  956.485000 -0.085000  956.655000 0.085000 ;
      RECT  956.485000  2.635000  956.655000 2.805000 ;
      RECT  956.945000 -0.085000  957.115000 0.085000 ;
      RECT  956.945000  2.635000  957.115000 2.805000 ;
      RECT  957.405000 -0.085000  957.575000 0.085000 ;
      RECT  957.405000  2.635000  957.575000 2.805000 ;
      RECT  957.865000 -0.085000  958.035000 0.085000 ;
      RECT  957.865000  2.635000  958.035000 2.805000 ;
      RECT  958.325000 -0.085000  958.495000 0.085000 ;
      RECT  958.325000  2.635000  958.495000 2.805000 ;
      RECT  958.785000 -0.085000  958.955000 0.085000 ;
      RECT  958.785000  2.635000  958.955000 2.805000 ;
      RECT  959.245000 -0.085000  959.415000 0.085000 ;
      RECT  959.245000  2.635000  959.415000 2.805000 ;
      RECT  959.705000 -0.085000  959.875000 0.085000 ;
      RECT  959.705000  2.635000  959.875000 2.805000 ;
      RECT  960.165000 -0.085000  960.335000 0.085000 ;
      RECT  960.165000  2.635000  960.335000 2.805000 ;
      RECT  960.625000 -0.085000  960.795000 0.085000 ;
      RECT  960.625000  2.635000  960.795000 2.805000 ;
      RECT  961.085000 -0.085000  961.255000 0.085000 ;
      RECT  961.085000  2.635000  961.255000 2.805000 ;
      RECT  961.545000 -0.085000  961.715000 0.085000 ;
      RECT  961.545000  2.635000  961.715000 2.805000 ;
      RECT  962.005000 -0.085000  962.175000 0.085000 ;
      RECT  962.005000  2.635000  962.175000 2.805000 ;
      RECT  962.465000 -0.085000  962.635000 0.085000 ;
      RECT  962.465000  2.635000  962.635000 2.805000 ;
      RECT  962.925000 -0.085000  963.095000 0.085000 ;
      RECT  962.925000  2.635000  963.095000 2.805000 ;
      RECT  963.385000 -0.085000  963.555000 0.085000 ;
      RECT  963.385000  2.635000  963.555000 2.805000 ;
      RECT  963.845000 -0.085000  964.015000 0.085000 ;
      RECT  963.845000  2.635000  964.015000 2.805000 ;
      RECT  964.305000 -0.085000  964.475000 0.085000 ;
      RECT  964.305000  2.635000  964.475000 2.805000 ;
      RECT  964.765000 -0.085000  964.935000 0.085000 ;
      RECT  964.765000  2.635000  964.935000 2.805000 ;
      RECT  965.225000 -0.085000  965.395000 0.085000 ;
      RECT  965.225000  2.635000  965.395000 2.805000 ;
      RECT  965.685000 -0.085000  965.855000 0.085000 ;
      RECT  965.685000  2.635000  965.855000 2.805000 ;
      RECT  966.145000 -0.085000  966.315000 0.085000 ;
      RECT  966.145000  2.635000  966.315000 2.805000 ;
      RECT  966.605000 -0.085000  966.775000 0.085000 ;
      RECT  966.605000  2.635000  966.775000 2.805000 ;
      RECT  967.065000 -0.085000  967.235000 0.085000 ;
      RECT  967.065000  2.635000  967.235000 2.805000 ;
      RECT  967.525000 -0.085000  967.695000 0.085000 ;
      RECT  967.525000  2.635000  967.695000 2.805000 ;
      RECT  967.985000 -0.085000  968.155000 0.085000 ;
      RECT  967.985000  2.635000  968.155000 2.805000 ;
      RECT  968.445000 -0.085000  968.615000 0.085000 ;
      RECT  968.445000  2.635000  968.615000 2.805000 ;
      RECT  968.905000 -0.085000  969.075000 0.085000 ;
      RECT  968.905000  2.635000  969.075000 2.805000 ;
      RECT  969.365000 -0.085000  969.535000 0.085000 ;
      RECT  969.365000  2.635000  969.535000 2.805000 ;
      RECT  969.825000 -0.085000  969.995000 0.085000 ;
      RECT  969.825000  2.635000  969.995000 2.805000 ;
      RECT  970.285000 -0.085000  970.455000 0.085000 ;
      RECT  970.285000  2.635000  970.455000 2.805000 ;
      RECT  970.745000 -0.085000  970.915000 0.085000 ;
      RECT  970.745000  2.635000  970.915000 2.805000 ;
      RECT  971.205000 -0.085000  971.375000 0.085000 ;
      RECT  971.205000  2.635000  971.375000 2.805000 ;
      RECT  971.665000 -0.085000  971.835000 0.085000 ;
      RECT  971.665000  2.635000  971.835000 2.805000 ;
      RECT  972.125000 -0.085000  972.295000 0.085000 ;
      RECT  972.125000  2.635000  972.295000 2.805000 ;
      RECT  972.585000 -0.085000  972.755000 0.085000 ;
      RECT  972.585000  2.635000  972.755000 2.805000 ;
      RECT  973.045000 -0.085000  973.215000 0.085000 ;
      RECT  973.045000  2.635000  973.215000 2.805000 ;
      RECT  973.505000 -0.085000  973.675000 0.085000 ;
      RECT  973.505000  2.635000  973.675000 2.805000 ;
      RECT  973.965000 -0.085000  974.135000 0.085000 ;
      RECT  973.965000  2.635000  974.135000 2.805000 ;
      RECT  974.425000 -0.085000  974.595000 0.085000 ;
      RECT  974.425000  2.635000  974.595000 2.805000 ;
      RECT  974.885000 -0.085000  975.055000 0.085000 ;
      RECT  974.885000  2.635000  975.055000 2.805000 ;
      RECT  975.345000 -0.085000  975.515000 0.085000 ;
      RECT  975.345000  2.635000  975.515000 2.805000 ;
      RECT  975.805000 -0.085000  975.975000 0.085000 ;
      RECT  975.805000  2.635000  975.975000 2.805000 ;
      RECT  976.265000 -0.085000  976.435000 0.085000 ;
      RECT  976.265000  2.635000  976.435000 2.805000 ;
      RECT  976.725000 -0.085000  976.895000 0.085000 ;
      RECT  976.725000  2.635000  976.895000 2.805000 ;
      RECT  977.185000 -0.085000  977.355000 0.085000 ;
      RECT  977.185000  2.635000  977.355000 2.805000 ;
      RECT  977.645000 -0.085000  977.815000 0.085000 ;
      RECT  977.645000  2.635000  977.815000 2.805000 ;
      RECT  978.105000 -0.085000  978.275000 0.085000 ;
      RECT  978.105000  2.635000  978.275000 2.805000 ;
      RECT  978.565000 -0.085000  978.735000 0.085000 ;
      RECT  978.565000  2.635000  978.735000 2.805000 ;
      RECT  979.025000 -0.085000  979.195000 0.085000 ;
      RECT  979.025000  2.635000  979.195000 2.805000 ;
      RECT  979.485000 -0.085000  979.655000 0.085000 ;
      RECT  979.485000  2.635000  979.655000 2.805000 ;
      RECT  979.945000 -0.085000  980.115000 0.085000 ;
      RECT  979.945000  2.635000  980.115000 2.805000 ;
      RECT  980.405000 -0.085000  980.575000 0.085000 ;
      RECT  980.405000  2.635000  980.575000 2.805000 ;
      RECT  980.865000 -0.085000  981.035000 0.085000 ;
      RECT  980.865000  2.635000  981.035000 2.805000 ;
      RECT  981.325000 -0.085000  981.495000 0.085000 ;
      RECT  981.325000  2.635000  981.495000 2.805000 ;
      RECT  981.785000 -0.085000  981.955000 0.085000 ;
      RECT  981.785000  2.635000  981.955000 2.805000 ;
      RECT  982.245000 -0.085000  982.415000 0.085000 ;
      RECT  982.245000  2.635000  982.415000 2.805000 ;
      RECT  982.705000 -0.085000  982.875000 0.085000 ;
      RECT  982.705000  2.635000  982.875000 2.805000 ;
      RECT  983.165000 -0.085000  983.335000 0.085000 ;
      RECT  983.165000  2.635000  983.335000 2.805000 ;
      RECT  983.625000 -0.085000  983.795000 0.085000 ;
      RECT  983.625000  2.635000  983.795000 2.805000 ;
      RECT  984.085000 -0.085000  984.255000 0.085000 ;
      RECT  984.085000  2.635000  984.255000 2.805000 ;
      RECT  984.545000 -0.085000  984.715000 0.085000 ;
      RECT  984.545000  2.635000  984.715000 2.805000 ;
      RECT  985.005000 -0.085000  985.175000 0.085000 ;
      RECT  985.005000  2.635000  985.175000 2.805000 ;
      RECT  985.465000 -0.085000  985.635000 0.085000 ;
      RECT  985.465000  2.635000  985.635000 2.805000 ;
      RECT  985.925000 -0.085000  986.095000 0.085000 ;
      RECT  985.925000  2.635000  986.095000 2.805000 ;
      RECT  986.385000 -0.085000  986.555000 0.085000 ;
      RECT  986.385000  2.635000  986.555000 2.805000 ;
      RECT  986.845000 -0.085000  987.015000 0.085000 ;
      RECT  986.845000  2.635000  987.015000 2.805000 ;
      RECT  987.305000 -0.085000  987.475000 0.085000 ;
      RECT  987.305000  2.635000  987.475000 2.805000 ;
      RECT  987.765000 -0.085000  987.935000 0.085000 ;
      RECT  987.765000  2.635000  987.935000 2.805000 ;
      RECT  988.225000 -0.085000  988.395000 0.085000 ;
      RECT  988.225000  2.635000  988.395000 2.805000 ;
      RECT  988.685000 -0.085000  988.855000 0.085000 ;
      RECT  988.685000  2.635000  988.855000 2.805000 ;
      RECT  989.145000 -0.085000  989.315000 0.085000 ;
      RECT  989.145000  2.635000  989.315000 2.805000 ;
      RECT  989.605000 -0.085000  989.775000 0.085000 ;
      RECT  989.605000  2.635000  989.775000 2.805000 ;
      RECT  990.065000 -0.085000  990.235000 0.085000 ;
      RECT  990.065000  2.635000  990.235000 2.805000 ;
      RECT  990.525000 -0.085000  990.695000 0.085000 ;
      RECT  990.525000  2.635000  990.695000 2.805000 ;
      RECT  990.985000 -0.085000  991.155000 0.085000 ;
      RECT  990.985000  2.635000  991.155000 2.805000 ;
      RECT  991.445000 -0.085000  991.615000 0.085000 ;
      RECT  991.445000  2.635000  991.615000 2.805000 ;
      RECT  991.905000 -0.085000  992.075000 0.085000 ;
      RECT  991.905000  2.635000  992.075000 2.805000 ;
      RECT  992.365000 -0.085000  992.535000 0.085000 ;
      RECT  992.365000  2.635000  992.535000 2.805000 ;
      RECT  992.825000 -0.085000  992.995000 0.085000 ;
      RECT  992.825000  2.635000  992.995000 2.805000 ;
      RECT  993.285000 -0.085000  993.455000 0.085000 ;
      RECT  993.285000  2.635000  993.455000 2.805000 ;
      RECT  993.745000 -0.085000  993.915000 0.085000 ;
      RECT  993.745000  2.635000  993.915000 2.805000 ;
      RECT  994.205000 -0.085000  994.375000 0.085000 ;
      RECT  994.205000  2.635000  994.375000 2.805000 ;
      RECT  994.665000 -0.085000  994.835000 0.085000 ;
      RECT  994.665000  2.635000  994.835000 2.805000 ;
      RECT  995.125000 -0.085000  995.295000 0.085000 ;
      RECT  995.125000  2.635000  995.295000 2.805000 ;
      RECT  995.585000 -0.085000  995.755000 0.085000 ;
      RECT  995.585000  2.635000  995.755000 2.805000 ;
      RECT  996.045000 -0.085000  996.215000 0.085000 ;
      RECT  996.045000  2.635000  996.215000 2.805000 ;
      RECT  996.505000 -0.085000  996.675000 0.085000 ;
      RECT  996.505000  2.635000  996.675000 2.805000 ;
      RECT  996.965000 -0.085000  997.135000 0.085000 ;
      RECT  996.965000  2.635000  997.135000 2.805000 ;
      RECT  997.425000 -0.085000  997.595000 0.085000 ;
      RECT  997.425000  2.635000  997.595000 2.805000 ;
      RECT  997.885000 -0.085000  998.055000 0.085000 ;
      RECT  997.885000  2.635000  998.055000 2.805000 ;
      RECT  998.345000 -0.085000  998.515000 0.085000 ;
      RECT  998.345000  2.635000  998.515000 2.805000 ;
      RECT  998.805000 -0.085000  998.975000 0.085000 ;
      RECT  998.805000  2.635000  998.975000 2.805000 ;
      RECT  999.265000 -0.085000  999.435000 0.085000 ;
      RECT  999.265000  2.635000  999.435000 2.805000 ;
      RECT  999.725000 -0.085000  999.895000 0.085000 ;
      RECT  999.725000  2.635000  999.895000 2.805000 ;
      RECT 1000.185000 -0.085000 1000.355000 0.085000 ;
      RECT 1000.185000  2.635000 1000.355000 2.805000 ;
      RECT 1000.645000 -0.085000 1000.815000 0.085000 ;
      RECT 1000.645000  2.635000 1000.815000 2.805000 ;
      RECT 1001.105000 -0.085000 1001.275000 0.085000 ;
      RECT 1001.105000  2.635000 1001.275000 2.805000 ;
      RECT 1001.565000 -0.085000 1001.735000 0.085000 ;
      RECT 1001.565000  2.635000 1001.735000 2.805000 ;
      RECT 1002.025000 -0.085000 1002.195000 0.085000 ;
      RECT 1002.025000  2.635000 1002.195000 2.805000 ;
      RECT 1002.485000 -0.085000 1002.655000 0.085000 ;
      RECT 1002.485000  2.635000 1002.655000 2.805000 ;
      RECT 1002.945000 -0.085000 1003.115000 0.085000 ;
      RECT 1002.945000  2.635000 1003.115000 2.805000 ;
      RECT 1003.405000 -0.085000 1003.575000 0.085000 ;
      RECT 1003.405000  2.635000 1003.575000 2.805000 ;
      RECT 1003.865000 -0.085000 1004.035000 0.085000 ;
      RECT 1003.865000  2.635000 1004.035000 2.805000 ;
      RECT 1004.325000 -0.085000 1004.495000 0.085000 ;
      RECT 1004.325000  2.635000 1004.495000 2.805000 ;
      RECT 1004.785000 -0.085000 1004.955000 0.085000 ;
      RECT 1004.785000  2.635000 1004.955000 2.805000 ;
      RECT 1005.245000 -0.085000 1005.415000 0.085000 ;
      RECT 1005.245000  2.635000 1005.415000 2.805000 ;
      RECT 1005.705000 -0.085000 1005.875000 0.085000 ;
      RECT 1005.705000  2.635000 1005.875000 2.805000 ;
      RECT 1006.165000 -0.085000 1006.335000 0.085000 ;
      RECT 1006.165000  2.635000 1006.335000 2.805000 ;
      RECT 1006.625000 -0.085000 1006.795000 0.085000 ;
      RECT 1006.625000  2.635000 1006.795000 2.805000 ;
      RECT 1007.085000 -0.085000 1007.255000 0.085000 ;
      RECT 1007.085000  2.635000 1007.255000 2.805000 ;
      RECT 1007.545000 -0.085000 1007.715000 0.085000 ;
      RECT 1007.545000  2.635000 1007.715000 2.805000 ;
      RECT 1008.005000 -0.085000 1008.175000 0.085000 ;
      RECT 1008.005000  2.635000 1008.175000 2.805000 ;
      RECT 1008.465000 -0.085000 1008.635000 0.085000 ;
      RECT 1008.465000  2.635000 1008.635000 2.805000 ;
      RECT 1008.925000 -0.085000 1009.095000 0.085000 ;
      RECT 1008.925000  2.635000 1009.095000 2.805000 ;
      RECT 1009.385000 -0.085000 1009.555000 0.085000 ;
      RECT 1009.385000  2.635000 1009.555000 2.805000 ;
      RECT 1009.845000 -0.085000 1010.015000 0.085000 ;
      RECT 1009.845000  2.635000 1010.015000 2.805000 ;
      RECT 1010.305000 -0.085000 1010.475000 0.085000 ;
      RECT 1010.305000  2.635000 1010.475000 2.805000 ;
      RECT 1010.765000 -0.085000 1010.935000 0.085000 ;
      RECT 1010.765000  2.635000 1010.935000 2.805000 ;
      RECT 1011.225000 -0.085000 1011.395000 0.085000 ;
      RECT 1011.225000  2.635000 1011.395000 2.805000 ;
      RECT 1011.685000 -0.085000 1011.855000 0.085000 ;
      RECT 1011.685000  2.635000 1011.855000 2.805000 ;
      RECT 1012.145000 -0.085000 1012.315000 0.085000 ;
      RECT 1012.145000  2.635000 1012.315000 2.805000 ;
      RECT 1012.605000 -0.085000 1012.775000 0.085000 ;
      RECT 1012.605000  2.635000 1012.775000 2.805000 ;
      RECT 1013.065000 -0.085000 1013.235000 0.085000 ;
      RECT 1013.065000  2.635000 1013.235000 2.805000 ;
      RECT 1013.525000 -0.085000 1013.695000 0.085000 ;
      RECT 1013.525000  2.635000 1013.695000 2.805000 ;
      RECT 1013.985000 -0.085000 1014.155000 0.085000 ;
      RECT 1013.985000  2.635000 1014.155000 2.805000 ;
      RECT 1014.445000 -0.085000 1014.615000 0.085000 ;
      RECT 1014.445000  2.635000 1014.615000 2.805000 ;
      RECT 1014.905000 -0.085000 1015.075000 0.085000 ;
      RECT 1014.905000  2.635000 1015.075000 2.805000 ;
      RECT 1015.365000 -0.085000 1015.535000 0.085000 ;
      RECT 1015.365000  2.635000 1015.535000 2.805000 ;
      RECT 1015.825000 -0.085000 1015.995000 0.085000 ;
      RECT 1015.825000  2.635000 1015.995000 2.805000 ;
      RECT 1016.285000 -0.085000 1016.455000 0.085000 ;
      RECT 1016.285000  2.635000 1016.455000 2.805000 ;
      RECT 1016.745000 -0.085000 1016.915000 0.085000 ;
      RECT 1016.745000  2.635000 1016.915000 2.805000 ;
      RECT 1017.205000 -0.085000 1017.375000 0.085000 ;
      RECT 1017.205000  2.635000 1017.375000 2.805000 ;
      RECT 1017.665000 -0.085000 1017.835000 0.085000 ;
      RECT 1017.665000  2.635000 1017.835000 2.805000 ;
      RECT 1018.125000 -0.085000 1018.295000 0.085000 ;
      RECT 1018.125000  2.635000 1018.295000 2.805000 ;
      RECT 1018.585000 -0.085000 1018.755000 0.085000 ;
      RECT 1018.585000  2.635000 1018.755000 2.805000 ;
      RECT 1019.045000 -0.085000 1019.215000 0.085000 ;
      RECT 1019.045000  2.635000 1019.215000 2.805000 ;
      RECT 1019.505000 -0.085000 1019.675000 0.085000 ;
      RECT 1019.505000  2.635000 1019.675000 2.805000 ;
      RECT 1019.965000 -0.085000 1020.135000 0.085000 ;
      RECT 1019.965000  2.635000 1020.135000 2.805000 ;
      RECT 1020.425000 -0.085000 1020.595000 0.085000 ;
      RECT 1020.425000  2.635000 1020.595000 2.805000 ;
      RECT 1020.885000 -0.085000 1021.055000 0.085000 ;
      RECT 1020.885000  2.635000 1021.055000 2.805000 ;
      RECT 1021.345000 -0.085000 1021.515000 0.085000 ;
      RECT 1021.345000  2.635000 1021.515000 2.805000 ;
      RECT 1021.805000 -0.085000 1021.975000 0.085000 ;
      RECT 1021.805000  2.635000 1021.975000 2.805000 ;
      RECT 1022.265000 -0.085000 1022.435000 0.085000 ;
      RECT 1022.265000  2.635000 1022.435000 2.805000 ;
      RECT 1022.725000 -0.085000 1022.895000 0.085000 ;
      RECT 1022.725000  2.635000 1022.895000 2.805000 ;
      RECT 1023.185000 -0.085000 1023.355000 0.085000 ;
      RECT 1023.185000  2.635000 1023.355000 2.805000 ;
      RECT 1023.645000 -0.085000 1023.815000 0.085000 ;
      RECT 1023.645000  2.635000 1023.815000 2.805000 ;
      RECT 1024.105000 -0.085000 1024.275000 0.085000 ;
      RECT 1024.105000  2.635000 1024.275000 2.805000 ;
      RECT 1024.565000 -0.085000 1024.735000 0.085000 ;
      RECT 1024.565000  2.635000 1024.735000 2.805000 ;
      RECT 1025.025000 -0.085000 1025.195000 0.085000 ;
      RECT 1025.025000  2.635000 1025.195000 2.805000 ;
      RECT 1025.485000 -0.085000 1025.655000 0.085000 ;
      RECT 1025.485000  2.635000 1025.655000 2.805000 ;
      RECT 1025.945000 -0.085000 1026.115000 0.085000 ;
      RECT 1025.945000  2.635000 1026.115000 2.805000 ;
      RECT 1026.405000 -0.085000 1026.575000 0.085000 ;
      RECT 1026.405000  2.635000 1026.575000 2.805000 ;
      RECT 1026.865000 -0.085000 1027.035000 0.085000 ;
      RECT 1026.865000  2.635000 1027.035000 2.805000 ;
      RECT 1027.325000 -0.085000 1027.495000 0.085000 ;
      RECT 1027.325000  2.635000 1027.495000 2.805000 ;
      RECT 1027.785000 -0.085000 1027.955000 0.085000 ;
      RECT 1027.785000  2.635000 1027.955000 2.805000 ;
      RECT 1028.245000 -0.085000 1028.415000 0.085000 ;
      RECT 1028.245000  2.635000 1028.415000 2.805000 ;
      RECT 1028.705000 -0.085000 1028.875000 0.085000 ;
      RECT 1028.705000  2.635000 1028.875000 2.805000 ;
      RECT 1029.165000 -0.085000 1029.335000 0.085000 ;
      RECT 1029.165000  2.635000 1029.335000 2.805000 ;
      RECT 1029.625000 -0.085000 1029.795000 0.085000 ;
      RECT 1029.625000  2.635000 1029.795000 2.805000 ;
      RECT 1030.085000 -0.085000 1030.255000 0.085000 ;
      RECT 1030.085000  2.635000 1030.255000 2.805000 ;
      RECT 1030.545000 -0.085000 1030.715000 0.085000 ;
      RECT 1030.545000  2.635000 1030.715000 2.805000 ;
      RECT 1031.005000 -0.085000 1031.175000 0.085000 ;
      RECT 1031.005000  2.635000 1031.175000 2.805000 ;
      RECT 1031.465000 -0.085000 1031.635000 0.085000 ;
      RECT 1031.465000  2.635000 1031.635000 2.805000 ;
      RECT 1031.925000 -0.085000 1032.095000 0.085000 ;
      RECT 1031.925000  2.635000 1032.095000 2.805000 ;
      RECT 1032.385000 -0.085000 1032.555000 0.085000 ;
      RECT 1032.385000  2.635000 1032.555000 2.805000 ;
      RECT 1032.845000 -0.085000 1033.015000 0.085000 ;
      RECT 1032.845000  2.635000 1033.015000 2.805000 ;
      RECT 1033.305000 -0.085000 1033.475000 0.085000 ;
      RECT 1033.305000  2.635000 1033.475000 2.805000 ;
      RECT 1033.765000 -0.085000 1033.935000 0.085000 ;
      RECT 1033.765000  2.635000 1033.935000 2.805000 ;
      RECT 1034.225000 -0.085000 1034.395000 0.085000 ;
      RECT 1034.225000  2.635000 1034.395000 2.805000 ;
      RECT 1034.685000 -0.085000 1034.855000 0.085000 ;
      RECT 1034.685000  2.635000 1034.855000 2.805000 ;
      RECT 1034.790000  0.425000 1034.960000 0.595000 ;
      RECT 1035.145000 -0.085000 1035.315000 0.085000 ;
      RECT 1035.145000  2.635000 1035.315000 2.805000 ;
      RECT 1035.605000 -0.085000 1035.775000 0.085000 ;
      RECT 1035.605000  2.635000 1035.775000 2.805000 ;
      RECT 1036.065000 -0.085000 1036.235000 0.085000 ;
      RECT 1036.065000  2.635000 1036.235000 2.805000 ;
      RECT 1036.525000 -0.085000 1036.695000 0.085000 ;
      RECT 1036.525000  2.635000 1036.695000 2.805000 ;
      RECT 1036.985000 -0.085000 1037.155000 0.085000 ;
      RECT 1036.985000  2.635000 1037.155000 2.805000 ;
      RECT 1037.445000 -0.085000 1037.615000 0.085000 ;
      RECT 1037.445000  2.635000 1037.615000 2.805000 ;
      RECT 1037.905000 -0.085000 1038.075000 0.085000 ;
      RECT 1037.905000  2.635000 1038.075000 2.805000 ;
      RECT 1038.365000 -0.085000 1038.535000 0.085000 ;
      RECT 1038.365000  2.635000 1038.535000 2.805000 ;
      RECT 1038.825000 -0.085000 1038.995000 0.085000 ;
      RECT 1038.825000  2.635000 1038.995000 2.805000 ;
      RECT 1039.285000 -0.085000 1039.455000 0.085000 ;
      RECT 1039.285000  2.635000 1039.455000 2.805000 ;
      RECT 1039.745000 -0.085000 1039.915000 0.085000 ;
      RECT 1039.745000  2.635000 1039.915000 2.805000 ;
      RECT 1040.205000 -0.085000 1040.375000 0.085000 ;
      RECT 1040.205000  2.635000 1040.375000 2.805000 ;
      RECT 1040.665000 -0.085000 1040.835000 0.085000 ;
      RECT 1040.665000  2.635000 1040.835000 2.805000 ;
      RECT 1041.125000 -0.085000 1041.295000 0.085000 ;
      RECT 1041.125000  2.635000 1041.295000 2.805000 ;
      RECT 1041.585000 -0.085000 1041.755000 0.085000 ;
      RECT 1041.585000  2.635000 1041.755000 2.805000 ;
      RECT 1041.940000  0.425000 1042.110000 0.595000 ;
      RECT 1042.045000 -0.085000 1042.215000 0.085000 ;
      RECT 1042.045000  2.635000 1042.215000 2.805000 ;
      RECT 1042.505000 -0.085000 1042.675000 0.085000 ;
      RECT 1042.505000  2.635000 1042.675000 2.805000 ;
      RECT 1042.965000 -0.085000 1043.135000 0.085000 ;
      RECT 1042.965000  2.635000 1043.135000 2.805000 ;
      RECT 1043.425000 -0.085000 1043.595000 0.085000 ;
      RECT 1043.425000  2.635000 1043.595000 2.805000 ;
      RECT 1043.885000 -0.085000 1044.055000 0.085000 ;
      RECT 1043.885000  2.635000 1044.055000 2.805000 ;
      RECT 1044.345000 -0.085000 1044.515000 0.085000 ;
      RECT 1044.345000  2.635000 1044.515000 2.805000 ;
      RECT 1044.805000 -0.085000 1044.975000 0.085000 ;
      RECT 1044.805000  2.635000 1044.975000 2.805000 ;
      RECT 1045.265000 -0.085000 1045.435000 0.085000 ;
      RECT 1045.265000  2.635000 1045.435000 2.805000 ;
      RECT 1045.725000 -0.085000 1045.895000 0.085000 ;
      RECT 1045.725000  2.635000 1045.895000 2.805000 ;
      RECT 1046.185000 -0.085000 1046.355000 0.085000 ;
      RECT 1046.185000  2.635000 1046.355000 2.805000 ;
      RECT 1046.645000 -0.085000 1046.815000 0.085000 ;
      RECT 1046.645000  2.635000 1046.815000 2.805000 ;
      RECT 1047.105000 -0.085000 1047.275000 0.085000 ;
      RECT 1047.105000  2.635000 1047.275000 2.805000 ;
      RECT 1047.565000 -0.085000 1047.735000 0.085000 ;
      RECT 1047.565000  2.635000 1047.735000 2.805000 ;
      RECT 1048.025000 -0.085000 1048.195000 0.085000 ;
      RECT 1048.025000  2.635000 1048.195000 2.805000 ;
      RECT 1048.485000 -0.085000 1048.655000 0.085000 ;
      RECT 1048.485000  2.635000 1048.655000 2.805000 ;
      RECT 1048.945000 -0.085000 1049.115000 0.085000 ;
      RECT 1048.945000  2.635000 1049.115000 2.805000 ;
      RECT 1049.405000 -0.085000 1049.575000 0.085000 ;
      RECT 1049.405000  2.635000 1049.575000 2.805000 ;
      RECT 1049.865000 -0.085000 1050.035000 0.085000 ;
      RECT 1049.865000  2.635000 1050.035000 2.805000 ;
      RECT 1050.325000 -0.085000 1050.495000 0.085000 ;
      RECT 1050.325000  2.635000 1050.495000 2.805000 ;
      RECT 1050.785000 -0.085000 1050.955000 0.085000 ;
      RECT 1050.785000  2.635000 1050.955000 2.805000 ;
      RECT 1051.245000 -0.085000 1051.415000 0.085000 ;
      RECT 1051.245000  2.635000 1051.415000 2.805000 ;
      RECT 1051.705000 -0.085000 1051.875000 0.085000 ;
      RECT 1051.705000  2.635000 1051.875000 2.805000 ;
      RECT 1052.165000 -0.085000 1052.335000 0.085000 ;
      RECT 1052.165000  2.635000 1052.335000 2.805000 ;
      RECT 1052.625000 -0.085000 1052.795000 0.085000 ;
      RECT 1052.625000  2.635000 1052.795000 2.805000 ;
      RECT 1053.085000 -0.085000 1053.255000 0.085000 ;
      RECT 1053.085000  2.635000 1053.255000 2.805000 ;
      RECT 1053.545000 -0.085000 1053.715000 0.085000 ;
      RECT 1053.545000  2.635000 1053.715000 2.805000 ;
      RECT 1054.005000 -0.085000 1054.175000 0.085000 ;
      RECT 1054.005000  2.635000 1054.175000 2.805000 ;
      RECT 1054.465000 -0.085000 1054.635000 0.085000 ;
      RECT 1054.465000  2.635000 1054.635000 2.805000 ;
      RECT 1054.925000 -0.085000 1055.095000 0.085000 ;
      RECT 1054.925000  2.635000 1055.095000 2.805000 ;
      RECT 1055.385000 -0.085000 1055.555000 0.085000 ;
      RECT 1055.385000  2.635000 1055.555000 2.805000 ;
      RECT 1055.845000 -0.085000 1056.015000 0.085000 ;
      RECT 1055.845000  2.635000 1056.015000 2.805000 ;
      RECT 1056.305000 -0.085000 1056.475000 0.085000 ;
      RECT 1056.305000  2.635000 1056.475000 2.805000 ;
      RECT 1056.765000 -0.085000 1056.935000 0.085000 ;
      RECT 1056.765000  2.635000 1056.935000 2.805000 ;
      RECT 1057.225000 -0.085000 1057.395000 0.085000 ;
      RECT 1057.225000  2.635000 1057.395000 2.805000 ;
      RECT 1057.685000 -0.085000 1057.855000 0.085000 ;
      RECT 1057.685000  2.635000 1057.855000 2.805000 ;
      RECT 1058.145000 -0.085000 1058.315000 0.085000 ;
      RECT 1058.145000  2.635000 1058.315000 2.805000 ;
      RECT 1058.605000 -0.085000 1058.775000 0.085000 ;
      RECT 1058.605000  2.635000 1058.775000 2.805000 ;
      RECT 1059.065000 -0.085000 1059.235000 0.085000 ;
      RECT 1059.065000  2.635000 1059.235000 2.805000 ;
      RECT 1059.525000 -0.085000 1059.695000 0.085000 ;
      RECT 1059.525000  2.635000 1059.695000 2.805000 ;
      RECT 1059.985000 -0.085000 1060.155000 0.085000 ;
      RECT 1059.985000  2.635000 1060.155000 2.805000 ;
      RECT 1060.445000 -0.085000 1060.615000 0.085000 ;
      RECT 1060.445000  2.635000 1060.615000 2.805000 ;
      RECT 1060.905000 -0.085000 1061.075000 0.085000 ;
      RECT 1060.905000  2.635000 1061.075000 2.805000 ;
      RECT 1061.365000 -0.085000 1061.535000 0.085000 ;
      RECT 1061.365000  2.635000 1061.535000 2.805000 ;
      RECT 1061.825000 -0.085000 1061.995000 0.085000 ;
      RECT 1061.825000  2.635000 1061.995000 2.805000 ;
      RECT 1062.285000 -0.085000 1062.455000 0.085000 ;
      RECT 1062.285000  2.635000 1062.455000 2.805000 ;
      RECT 1062.745000 -0.085000 1062.915000 0.085000 ;
      RECT 1062.745000  2.635000 1062.915000 2.805000 ;
      RECT 1063.205000 -0.085000 1063.375000 0.085000 ;
      RECT 1063.205000  2.635000 1063.375000 2.805000 ;
      RECT 1063.665000 -0.085000 1063.835000 0.085000 ;
      RECT 1063.665000  2.635000 1063.835000 2.805000 ;
      RECT 1064.125000 -0.085000 1064.295000 0.085000 ;
      RECT 1064.125000  2.635000 1064.295000 2.805000 ;
      RECT 1064.585000 -0.085000 1064.755000 0.085000 ;
      RECT 1064.585000  2.635000 1064.755000 2.805000 ;
      RECT 1065.045000 -0.085000 1065.215000 0.085000 ;
      RECT 1065.045000  2.635000 1065.215000 2.805000 ;
      RECT 1065.505000 -0.085000 1065.675000 0.085000 ;
      RECT 1065.505000  2.635000 1065.675000 2.805000 ;
      RECT 1065.965000 -0.085000 1066.135000 0.085000 ;
      RECT 1065.965000  2.635000 1066.135000 2.805000 ;
      RECT 1066.425000 -0.085000 1066.595000 0.085000 ;
      RECT 1066.425000  2.635000 1066.595000 2.805000 ;
      RECT 1066.885000 -0.085000 1067.055000 0.085000 ;
      RECT 1066.885000  2.635000 1067.055000 2.805000 ;
      RECT 1067.345000 -0.085000 1067.515000 0.085000 ;
      RECT 1067.345000  2.635000 1067.515000 2.805000 ;
      RECT 1067.805000 -0.085000 1067.975000 0.085000 ;
      RECT 1067.805000  2.635000 1067.975000 2.805000 ;
      RECT 1068.265000 -0.085000 1068.435000 0.085000 ;
      RECT 1068.265000  2.635000 1068.435000 2.805000 ;
      RECT 1068.725000 -0.085000 1068.895000 0.085000 ;
      RECT 1068.725000  2.635000 1068.895000 2.805000 ;
      RECT 1069.185000 -0.085000 1069.355000 0.085000 ;
      RECT 1069.185000  2.635000 1069.355000 2.805000 ;
      RECT 1069.645000 -0.085000 1069.815000 0.085000 ;
      RECT 1069.645000  2.635000 1069.815000 2.805000 ;
      RECT 1070.105000 -0.085000 1070.275000 0.085000 ;
      RECT 1070.105000  2.635000 1070.275000 2.805000 ;
      RECT 1070.565000 -0.085000 1070.735000 0.085000 ;
      RECT 1070.565000  2.635000 1070.735000 2.805000 ;
      RECT 1071.025000 -0.085000 1071.195000 0.085000 ;
      RECT 1071.025000  2.635000 1071.195000 2.805000 ;
      RECT 1071.485000 -0.085000 1071.655000 0.085000 ;
      RECT 1071.485000  2.635000 1071.655000 2.805000 ;
      RECT 1071.945000 -0.085000 1072.115000 0.085000 ;
      RECT 1071.945000  2.635000 1072.115000 2.805000 ;
      RECT 1072.405000 -0.085000 1072.575000 0.085000 ;
      RECT 1072.405000  2.635000 1072.575000 2.805000 ;
      RECT 1072.865000 -0.085000 1073.035000 0.085000 ;
      RECT 1072.865000  2.635000 1073.035000 2.805000 ;
      RECT 1073.325000 -0.085000 1073.495000 0.085000 ;
      RECT 1073.325000  2.635000 1073.495000 2.805000 ;
      RECT 1073.785000 -0.085000 1073.955000 0.085000 ;
      RECT 1073.785000  2.635000 1073.955000 2.805000 ;
      RECT 1074.245000 -0.085000 1074.415000 0.085000 ;
      RECT 1074.245000  2.635000 1074.415000 2.805000 ;
      RECT 1074.705000 -0.085000 1074.875000 0.085000 ;
      RECT 1074.705000  2.635000 1074.875000 2.805000 ;
      RECT 1075.165000 -0.085000 1075.335000 0.085000 ;
      RECT 1075.165000  2.635000 1075.335000 2.805000 ;
      RECT 1075.625000 -0.085000 1075.795000 0.085000 ;
      RECT 1075.625000  2.635000 1075.795000 2.805000 ;
      RECT 1076.085000 -0.085000 1076.255000 0.085000 ;
      RECT 1076.085000  2.635000 1076.255000 2.805000 ;
      RECT 1076.545000 -0.085000 1076.715000 0.085000 ;
      RECT 1076.545000  2.635000 1076.715000 2.805000 ;
      RECT 1077.005000 -0.085000 1077.175000 0.085000 ;
      RECT 1077.005000  2.635000 1077.175000 2.805000 ;
      RECT 1077.465000 -0.085000 1077.635000 0.085000 ;
      RECT 1077.465000  2.635000 1077.635000 2.805000 ;
      RECT 1077.925000 -0.085000 1078.095000 0.085000 ;
      RECT 1077.925000  2.635000 1078.095000 2.805000 ;
      RECT 1078.385000 -0.085000 1078.555000 0.085000 ;
      RECT 1078.385000  2.635000 1078.555000 2.805000 ;
      RECT 1078.845000 -0.085000 1079.015000 0.085000 ;
      RECT 1078.845000  2.635000 1079.015000 2.805000 ;
      RECT 1079.305000 -0.085000 1079.475000 0.085000 ;
      RECT 1079.305000  2.635000 1079.475000 2.805000 ;
      RECT 1079.765000 -0.085000 1079.935000 0.085000 ;
      RECT 1079.765000  2.635000 1079.935000 2.805000 ;
      RECT 1080.225000 -0.085000 1080.395000 0.085000 ;
      RECT 1080.225000  2.635000 1080.395000 2.805000 ;
      RECT 1080.685000 -0.085000 1080.855000 0.085000 ;
      RECT 1080.685000  2.635000 1080.855000 2.805000 ;
      RECT 1081.145000 -0.085000 1081.315000 0.085000 ;
      RECT 1081.145000  2.635000 1081.315000 2.805000 ;
      RECT 1081.605000 -0.085000 1081.775000 0.085000 ;
      RECT 1081.605000  2.635000 1081.775000 2.805000 ;
      RECT 1082.065000 -0.085000 1082.235000 0.085000 ;
      RECT 1082.065000  2.635000 1082.235000 2.805000 ;
      RECT 1082.525000 -0.085000 1082.695000 0.085000 ;
      RECT 1082.525000  2.635000 1082.695000 2.805000 ;
      RECT 1082.985000 -0.085000 1083.155000 0.085000 ;
      RECT 1082.985000  2.635000 1083.155000 2.805000 ;
      RECT 1083.445000 -0.085000 1083.615000 0.085000 ;
      RECT 1083.445000  2.635000 1083.615000 2.805000 ;
      RECT 1083.905000 -0.085000 1084.075000 0.085000 ;
      RECT 1083.905000  2.635000 1084.075000 2.805000 ;
      RECT 1084.365000 -0.085000 1084.535000 0.085000 ;
      RECT 1084.365000  2.635000 1084.535000 2.805000 ;
      RECT 1084.825000 -0.085000 1084.995000 0.085000 ;
      RECT 1084.825000  2.635000 1084.995000 2.805000 ;
      RECT 1085.285000 -0.085000 1085.455000 0.085000 ;
      RECT 1085.285000  2.635000 1085.455000 2.805000 ;
      RECT 1085.745000 -0.085000 1085.915000 0.085000 ;
      RECT 1085.745000  2.635000 1085.915000 2.805000 ;
      RECT 1086.205000 -0.085000 1086.375000 0.085000 ;
      RECT 1086.205000  2.635000 1086.375000 2.805000 ;
      RECT 1086.665000 -0.085000 1086.835000 0.085000 ;
      RECT 1086.665000  2.635000 1086.835000 2.805000 ;
      RECT 1087.125000 -0.085000 1087.295000 0.085000 ;
      RECT 1087.125000  2.635000 1087.295000 2.805000 ;
      RECT 1087.585000 -0.085000 1087.755000 0.085000 ;
      RECT 1087.585000  2.635000 1087.755000 2.805000 ;
      RECT 1088.045000 -0.085000 1088.215000 0.085000 ;
      RECT 1088.045000  2.635000 1088.215000 2.805000 ;
      RECT 1088.505000 -0.085000 1088.675000 0.085000 ;
      RECT 1088.505000  2.635000 1088.675000 2.805000 ;
      RECT 1088.965000 -0.085000 1089.135000 0.085000 ;
      RECT 1088.965000  2.635000 1089.135000 2.805000 ;
      RECT 1089.425000 -0.085000 1089.595000 0.085000 ;
      RECT 1089.425000  2.635000 1089.595000 2.805000 ;
      RECT 1089.885000 -0.085000 1090.055000 0.085000 ;
      RECT 1089.885000  2.635000 1090.055000 2.805000 ;
      RECT 1090.345000 -0.085000 1090.515000 0.085000 ;
      RECT 1090.345000  2.635000 1090.515000 2.805000 ;
      RECT 1090.805000 -0.085000 1090.975000 0.085000 ;
      RECT 1090.805000  2.635000 1090.975000 2.805000 ;
      RECT 1091.265000 -0.085000 1091.435000 0.085000 ;
      RECT 1091.265000  2.635000 1091.435000 2.805000 ;
      RECT 1091.725000 -0.085000 1091.895000 0.085000 ;
      RECT 1091.725000  2.635000 1091.895000 2.805000 ;
      RECT 1092.185000 -0.085000 1092.355000 0.085000 ;
      RECT 1092.185000  2.635000 1092.355000 2.805000 ;
      RECT 1092.645000 -0.085000 1092.815000 0.085000 ;
      RECT 1092.645000  2.635000 1092.815000 2.805000 ;
      RECT 1093.105000 -0.085000 1093.275000 0.085000 ;
      RECT 1093.105000  2.635000 1093.275000 2.805000 ;
      RECT 1093.565000 -0.085000 1093.735000 0.085000 ;
      RECT 1093.565000  2.635000 1093.735000 2.805000 ;
      RECT 1094.025000 -0.085000 1094.195000 0.085000 ;
      RECT 1094.025000  2.635000 1094.195000 2.805000 ;
      RECT 1094.485000 -0.085000 1094.655000 0.085000 ;
      RECT 1094.485000  2.635000 1094.655000 2.805000 ;
      RECT 1094.945000 -0.085000 1095.115000 0.085000 ;
      RECT 1094.945000  2.635000 1095.115000 2.805000 ;
      RECT 1095.405000 -0.085000 1095.575000 0.085000 ;
      RECT 1095.405000  2.635000 1095.575000 2.805000 ;
      RECT 1095.865000 -0.085000 1096.035000 0.085000 ;
      RECT 1095.865000  2.635000 1096.035000 2.805000 ;
      RECT 1096.325000 -0.085000 1096.495000 0.085000 ;
      RECT 1096.325000  2.635000 1096.495000 2.805000 ;
      RECT 1096.785000 -0.085000 1096.955000 0.085000 ;
      RECT 1096.785000  2.635000 1096.955000 2.805000 ;
      RECT 1097.245000 -0.085000 1097.415000 0.085000 ;
      RECT 1097.245000  2.635000 1097.415000 2.805000 ;
      RECT 1097.705000 -0.085000 1097.875000 0.085000 ;
      RECT 1097.705000  2.635000 1097.875000 2.805000 ;
      RECT 1098.165000 -0.085000 1098.335000 0.085000 ;
      RECT 1098.165000  2.635000 1098.335000 2.805000 ;
      RECT 1098.625000 -0.085000 1098.795000 0.085000 ;
      RECT 1098.625000  2.635000 1098.795000 2.805000 ;
      RECT 1099.085000 -0.085000 1099.255000 0.085000 ;
      RECT 1099.085000  2.635000 1099.255000 2.805000 ;
      RECT 1099.545000 -0.085000 1099.715000 0.085000 ;
      RECT 1099.545000  2.635000 1099.715000 2.805000 ;
      RECT 1100.005000 -0.085000 1100.175000 0.085000 ;
      RECT 1100.005000  2.635000 1100.175000 2.805000 ;
      RECT 1100.465000 -0.085000 1100.635000 0.085000 ;
      RECT 1100.465000  2.635000 1100.635000 2.805000 ;
      RECT 1100.925000 -0.085000 1101.095000 0.085000 ;
      RECT 1100.925000  2.635000 1101.095000 2.805000 ;
      RECT 1101.385000 -0.085000 1101.555000 0.085000 ;
      RECT 1101.385000  2.635000 1101.555000 2.805000 ;
      RECT 1101.845000 -0.085000 1102.015000 0.085000 ;
      RECT 1101.845000  2.635000 1102.015000 2.805000 ;
      RECT 1102.305000 -0.085000 1102.475000 0.085000 ;
      RECT 1102.305000  2.635000 1102.475000 2.805000 ;
      RECT 1102.765000 -0.085000 1102.935000 0.085000 ;
      RECT 1102.765000  2.635000 1102.935000 2.805000 ;
      RECT 1103.225000 -0.085000 1103.395000 0.085000 ;
      RECT 1103.225000  2.635000 1103.395000 2.805000 ;
      RECT 1103.685000 -0.085000 1103.855000 0.085000 ;
      RECT 1103.685000  2.635000 1103.855000 2.805000 ;
      RECT 1104.145000 -0.085000 1104.315000 0.085000 ;
      RECT 1104.145000  2.635000 1104.315000 2.805000 ;
      RECT 1104.605000 -0.085000 1104.775000 0.085000 ;
      RECT 1104.605000  2.635000 1104.775000 2.805000 ;
      RECT 1105.065000 -0.085000 1105.235000 0.085000 ;
      RECT 1105.065000  2.635000 1105.235000 2.805000 ;
      RECT 1105.525000 -0.085000 1105.695000 0.085000 ;
      RECT 1105.525000  2.635000 1105.695000 2.805000 ;
      RECT 1105.985000 -0.085000 1106.155000 0.085000 ;
      RECT 1105.985000  2.635000 1106.155000 2.805000 ;
      RECT 1106.445000 -0.085000 1106.615000 0.085000 ;
      RECT 1106.445000  2.635000 1106.615000 2.805000 ;
      RECT 1106.905000 -0.085000 1107.075000 0.085000 ;
      RECT 1106.905000  2.635000 1107.075000 2.805000 ;
      RECT 1107.365000 -0.085000 1107.535000 0.085000 ;
      RECT 1107.365000  2.635000 1107.535000 2.805000 ;
      RECT 1107.825000 -0.085000 1107.995000 0.085000 ;
      RECT 1107.825000  2.635000 1107.995000 2.805000 ;
      RECT 1108.285000 -0.085000 1108.455000 0.085000 ;
      RECT 1108.285000  2.635000 1108.455000 2.805000 ;
      RECT 1108.745000 -0.085000 1108.915000 0.085000 ;
      RECT 1108.745000  2.635000 1108.915000 2.805000 ;
      RECT 1109.205000 -0.085000 1109.375000 0.085000 ;
      RECT 1109.205000  2.635000 1109.375000 2.805000 ;
      RECT 1109.665000 -0.085000 1109.835000 0.085000 ;
      RECT 1109.665000  2.635000 1109.835000 2.805000 ;
      RECT 1110.125000 -0.085000 1110.295000 0.085000 ;
      RECT 1110.125000  2.635000 1110.295000 2.805000 ;
      RECT 1110.585000 -0.085000 1110.755000 0.085000 ;
      RECT 1110.585000  2.635000 1110.755000 2.805000 ;
      RECT 1111.045000 -0.085000 1111.215000 0.085000 ;
      RECT 1111.045000  2.635000 1111.215000 2.805000 ;
      RECT 1111.505000 -0.085000 1111.675000 0.085000 ;
      RECT 1111.505000  2.635000 1111.675000 2.805000 ;
      RECT 1111.965000 -0.085000 1112.135000 0.085000 ;
      RECT 1111.965000  2.635000 1112.135000 2.805000 ;
      RECT 1112.425000 -0.085000 1112.595000 0.085000 ;
      RECT 1112.425000  2.635000 1112.595000 2.805000 ;
      RECT 1112.885000 -0.085000 1113.055000 0.085000 ;
      RECT 1112.885000  2.635000 1113.055000 2.805000 ;
      RECT 1113.345000 -0.085000 1113.515000 0.085000 ;
      RECT 1113.345000  2.635000 1113.515000 2.805000 ;
      RECT 1113.805000 -0.085000 1113.975000 0.085000 ;
      RECT 1113.805000  2.635000 1113.975000 2.805000 ;
      RECT 1114.265000 -0.085000 1114.435000 0.085000 ;
      RECT 1114.265000  2.635000 1114.435000 2.805000 ;
      RECT 1114.725000 -0.085000 1114.895000 0.085000 ;
      RECT 1114.725000  2.635000 1114.895000 2.805000 ;
      RECT 1115.185000 -0.085000 1115.355000 0.085000 ;
      RECT 1115.185000  2.635000 1115.355000 2.805000 ;
      RECT 1115.645000 -0.085000 1115.815000 0.085000 ;
      RECT 1115.645000  2.635000 1115.815000 2.805000 ;
      RECT 1116.105000 -0.085000 1116.275000 0.085000 ;
      RECT 1116.105000  2.635000 1116.275000 2.805000 ;
      RECT 1116.565000 -0.085000 1116.735000 0.085000 ;
      RECT 1116.565000  2.635000 1116.735000 2.805000 ;
      RECT 1117.025000 -0.085000 1117.195000 0.085000 ;
      RECT 1117.025000  2.635000 1117.195000 2.805000 ;
      RECT 1117.485000 -0.085000 1117.655000 0.085000 ;
      RECT 1117.485000  2.635000 1117.655000 2.805000 ;
      RECT 1117.945000 -0.085000 1118.115000 0.085000 ;
      RECT 1117.945000  2.635000 1118.115000 2.805000 ;
      RECT 1118.405000 -0.085000 1118.575000 0.085000 ;
      RECT 1118.405000  2.635000 1118.575000 2.805000 ;
      RECT 1118.865000 -0.085000 1119.035000 0.085000 ;
      RECT 1118.865000  2.635000 1119.035000 2.805000 ;
      RECT 1119.325000 -0.085000 1119.495000 0.085000 ;
      RECT 1119.325000  2.635000 1119.495000 2.805000 ;
      RECT 1119.785000 -0.085000 1119.955000 0.085000 ;
      RECT 1119.785000  2.635000 1119.955000 2.805000 ;
      RECT 1120.245000 -0.085000 1120.415000 0.085000 ;
      RECT 1120.245000  2.635000 1120.415000 2.805000 ;
      RECT 1120.705000 -0.085000 1120.875000 0.085000 ;
      RECT 1120.705000  2.635000 1120.875000 2.805000 ;
      RECT 1121.165000 -0.085000 1121.335000 0.085000 ;
      RECT 1121.165000  2.635000 1121.335000 2.805000 ;
      RECT 1121.625000 -0.085000 1121.795000 0.085000 ;
      RECT 1121.625000  2.635000 1121.795000 2.805000 ;
      RECT 1122.085000 -0.085000 1122.255000 0.085000 ;
      RECT 1122.085000  2.635000 1122.255000 2.805000 ;
      RECT 1122.545000 -0.085000 1122.715000 0.085000 ;
      RECT 1122.545000  2.635000 1122.715000 2.805000 ;
      RECT 1123.005000 -0.085000 1123.175000 0.085000 ;
      RECT 1123.005000  2.635000 1123.175000 2.805000 ;
      RECT 1123.465000 -0.085000 1123.635000 0.085000 ;
      RECT 1123.465000  2.635000 1123.635000 2.805000 ;
      RECT 1123.925000 -0.085000 1124.095000 0.085000 ;
      RECT 1123.925000  2.635000 1124.095000 2.805000 ;
      RECT 1124.385000 -0.085000 1124.555000 0.085000 ;
      RECT 1124.385000  2.635000 1124.555000 2.805000 ;
      RECT 1124.845000 -0.085000 1125.015000 0.085000 ;
      RECT 1124.845000  2.635000 1125.015000 2.805000 ;
      RECT 1125.305000 -0.085000 1125.475000 0.085000 ;
      RECT 1125.305000  2.635000 1125.475000 2.805000 ;
      RECT 1125.765000 -0.085000 1125.935000 0.085000 ;
      RECT 1125.765000  2.635000 1125.935000 2.805000 ;
      RECT 1126.225000 -0.085000 1126.395000 0.085000 ;
      RECT 1126.225000  2.635000 1126.395000 2.805000 ;
      RECT 1126.685000 -0.085000 1126.855000 0.085000 ;
      RECT 1126.685000  2.635000 1126.855000 2.805000 ;
      RECT 1127.145000 -0.085000 1127.315000 0.085000 ;
      RECT 1127.145000  2.635000 1127.315000 2.805000 ;
      RECT 1127.605000 -0.085000 1127.775000 0.085000 ;
      RECT 1127.605000  2.635000 1127.775000 2.805000 ;
      RECT 1128.065000 -0.085000 1128.235000 0.085000 ;
      RECT 1128.065000  2.635000 1128.235000 2.805000 ;
      RECT 1128.525000 -0.085000 1128.695000 0.085000 ;
      RECT 1128.525000  2.635000 1128.695000 2.805000 ;
      RECT 1128.985000 -0.085000 1129.155000 0.085000 ;
      RECT 1128.985000  2.635000 1129.155000 2.805000 ;
      RECT 1129.445000 -0.085000 1129.615000 0.085000 ;
      RECT 1129.445000  2.635000 1129.615000 2.805000 ;
      RECT 1129.905000 -0.085000 1130.075000 0.085000 ;
      RECT 1129.905000  2.635000 1130.075000 2.805000 ;
      RECT 1130.365000 -0.085000 1130.535000 0.085000 ;
      RECT 1130.365000  2.635000 1130.535000 2.805000 ;
      RECT 1130.825000 -0.085000 1130.995000 0.085000 ;
      RECT 1130.825000  2.635000 1130.995000 2.805000 ;
      RECT 1131.285000 -0.085000 1131.455000 0.085000 ;
      RECT 1131.285000  2.635000 1131.455000 2.805000 ;
      RECT 1131.745000 -0.085000 1131.915000 0.085000 ;
      RECT 1131.745000  2.635000 1131.915000 2.805000 ;
      RECT 1132.205000 -0.085000 1132.375000 0.085000 ;
      RECT 1132.205000  2.635000 1132.375000 2.805000 ;
      RECT 1132.665000 -0.085000 1132.835000 0.085000 ;
      RECT 1132.665000  2.635000 1132.835000 2.805000 ;
      RECT 1133.125000 -0.085000 1133.295000 0.085000 ;
      RECT 1133.125000  2.635000 1133.295000 2.805000 ;
      RECT 1133.585000 -0.085000 1133.755000 0.085000 ;
      RECT 1133.585000  2.635000 1133.755000 2.805000 ;
      RECT 1134.045000 -0.085000 1134.215000 0.085000 ;
      RECT 1134.045000  2.635000 1134.215000 2.805000 ;
      RECT 1134.505000 -0.085000 1134.675000 0.085000 ;
      RECT 1134.505000  2.635000 1134.675000 2.805000 ;
      RECT 1134.965000 -0.085000 1135.135000 0.085000 ;
      RECT 1134.965000  2.635000 1135.135000 2.805000 ;
      RECT 1135.425000 -0.085000 1135.595000 0.085000 ;
      RECT 1135.425000  2.635000 1135.595000 2.805000 ;
      RECT 1135.885000 -0.085000 1136.055000 0.085000 ;
      RECT 1135.885000  2.635000 1136.055000 2.805000 ;
      RECT 1136.345000 -0.085000 1136.515000 0.085000 ;
      RECT 1136.345000  2.635000 1136.515000 2.805000 ;
      RECT 1136.805000 -0.085000 1136.975000 0.085000 ;
      RECT 1136.805000  2.635000 1136.975000 2.805000 ;
      RECT 1137.265000 -0.085000 1137.435000 0.085000 ;
      RECT 1137.265000  2.635000 1137.435000 2.805000 ;
      RECT 1137.725000 -0.085000 1137.895000 0.085000 ;
      RECT 1137.725000  2.635000 1137.895000 2.805000 ;
      RECT 1138.185000 -0.085000 1138.355000 0.085000 ;
      RECT 1138.185000  2.635000 1138.355000 2.805000 ;
      RECT 1138.645000 -0.085000 1138.815000 0.085000 ;
      RECT 1138.645000  2.635000 1138.815000 2.805000 ;
      RECT 1139.105000 -0.085000 1139.275000 0.085000 ;
      RECT 1139.105000  2.635000 1139.275000 2.805000 ;
      RECT 1139.565000 -0.085000 1139.735000 0.085000 ;
      RECT 1139.565000  2.635000 1139.735000 2.805000 ;
      RECT 1140.025000 -0.085000 1140.195000 0.085000 ;
      RECT 1140.025000  2.635000 1140.195000 2.805000 ;
      RECT 1140.485000 -0.085000 1140.655000 0.085000 ;
      RECT 1140.485000  2.635000 1140.655000 2.805000 ;
      RECT 1140.945000 -0.085000 1141.115000 0.085000 ;
      RECT 1140.945000  2.635000 1141.115000 2.805000 ;
      RECT 1141.405000 -0.085000 1141.575000 0.085000 ;
      RECT 1141.405000  2.635000 1141.575000 2.805000 ;
      RECT 1141.865000 -0.085000 1142.035000 0.085000 ;
      RECT 1141.865000  2.635000 1142.035000 2.805000 ;
      RECT 1142.325000 -0.085000 1142.495000 0.085000 ;
      RECT 1142.325000  2.635000 1142.495000 2.805000 ;
      RECT 1142.785000 -0.085000 1142.955000 0.085000 ;
      RECT 1142.785000  2.635000 1142.955000 2.805000 ;
      RECT 1143.245000 -0.085000 1143.415000 0.085000 ;
      RECT 1143.245000  2.635000 1143.415000 2.805000 ;
      RECT 1143.705000 -0.085000 1143.875000 0.085000 ;
      RECT 1143.705000  2.635000 1143.875000 2.805000 ;
      RECT 1144.165000 -0.085000 1144.335000 0.085000 ;
      RECT 1144.165000  2.635000 1144.335000 2.805000 ;
      RECT 1144.625000 -0.085000 1144.795000 0.085000 ;
      RECT 1144.625000  2.635000 1144.795000 2.805000 ;
      RECT 1145.085000 -0.085000 1145.255000 0.085000 ;
      RECT 1145.085000  2.635000 1145.255000 2.805000 ;
      RECT 1145.545000 -0.085000 1145.715000 0.085000 ;
      RECT 1145.545000  2.635000 1145.715000 2.805000 ;
      RECT 1146.005000 -0.085000 1146.175000 0.085000 ;
      RECT 1146.005000  2.635000 1146.175000 2.805000 ;
      RECT 1146.465000 -0.085000 1146.635000 0.085000 ;
      RECT 1146.465000  2.635000 1146.635000 2.805000 ;
      RECT 1146.925000 -0.085000 1147.095000 0.085000 ;
      RECT 1146.925000  2.635000 1147.095000 2.805000 ;
      RECT 1147.385000 -0.085000 1147.555000 0.085000 ;
      RECT 1147.385000  2.635000 1147.555000 2.805000 ;
      RECT 1147.845000 -0.085000 1148.015000 0.085000 ;
      RECT 1147.845000  2.635000 1148.015000 2.805000 ;
      RECT 1148.305000 -0.085000 1148.475000 0.085000 ;
      RECT 1148.305000  2.635000 1148.475000 2.805000 ;
      RECT 1148.765000 -0.085000 1148.935000 0.085000 ;
      RECT 1148.765000  2.635000 1148.935000 2.805000 ;
      RECT 1149.225000 -0.085000 1149.395000 0.085000 ;
      RECT 1149.225000  2.635000 1149.395000 2.805000 ;
      RECT 1149.685000 -0.085000 1149.855000 0.085000 ;
      RECT 1149.685000  2.635000 1149.855000 2.805000 ;
      RECT 1150.145000 -0.085000 1150.315000 0.085000 ;
      RECT 1150.145000  2.635000 1150.315000 2.805000 ;
      RECT 1150.605000 -0.085000 1150.775000 0.085000 ;
      RECT 1150.605000  2.635000 1150.775000 2.805000 ;
      RECT 1151.065000 -0.085000 1151.235000 0.085000 ;
      RECT 1151.065000  2.635000 1151.235000 2.805000 ;
      RECT 1151.525000 -0.085000 1151.695000 0.085000 ;
      RECT 1151.525000  2.635000 1151.695000 2.805000 ;
      RECT 1151.985000 -0.085000 1152.155000 0.085000 ;
      RECT 1151.985000  2.635000 1152.155000 2.805000 ;
      RECT 1152.445000 -0.085000 1152.615000 0.085000 ;
      RECT 1152.445000  2.635000 1152.615000 2.805000 ;
      RECT 1152.905000 -0.085000 1153.075000 0.085000 ;
      RECT 1152.905000  2.635000 1153.075000 2.805000 ;
      RECT 1153.365000 -0.085000 1153.535000 0.085000 ;
      RECT 1153.365000  2.635000 1153.535000 2.805000 ;
      RECT 1153.825000 -0.085000 1153.995000 0.085000 ;
      RECT 1153.825000  2.635000 1153.995000 2.805000 ;
      RECT 1154.285000 -0.085000 1154.455000 0.085000 ;
      RECT 1154.285000  2.635000 1154.455000 2.805000 ;
      RECT 1154.745000 -0.085000 1154.915000 0.085000 ;
      RECT 1154.745000  2.635000 1154.915000 2.805000 ;
      RECT 1155.205000 -0.085000 1155.375000 0.085000 ;
      RECT 1155.205000  2.635000 1155.375000 2.805000 ;
      RECT 1155.665000 -0.085000 1155.835000 0.085000 ;
      RECT 1155.665000  2.635000 1155.835000 2.805000 ;
      RECT 1156.125000 -0.085000 1156.295000 0.085000 ;
      RECT 1156.125000  2.635000 1156.295000 2.805000 ;
      RECT 1156.585000 -0.085000 1156.755000 0.085000 ;
      RECT 1156.585000  2.635000 1156.755000 2.805000 ;
      RECT 1157.045000 -0.085000 1157.215000 0.085000 ;
      RECT 1157.045000  2.635000 1157.215000 2.805000 ;
      RECT 1157.505000 -0.085000 1157.675000 0.085000 ;
      RECT 1157.505000  2.635000 1157.675000 2.805000 ;
      RECT 1157.965000 -0.085000 1158.135000 0.085000 ;
      RECT 1157.965000  2.635000 1158.135000 2.805000 ;
      RECT 1158.425000 -0.085000 1158.595000 0.085000 ;
      RECT 1158.425000  2.635000 1158.595000 2.805000 ;
      RECT 1158.885000 -0.085000 1159.055000 0.085000 ;
      RECT 1158.885000  2.635000 1159.055000 2.805000 ;
      RECT 1159.345000 -0.085000 1159.515000 0.085000 ;
      RECT 1159.345000  2.635000 1159.515000 2.805000 ;
      RECT 1159.805000 -0.085000 1159.975000 0.085000 ;
      RECT 1159.805000  2.635000 1159.975000 2.805000 ;
      RECT 1160.265000 -0.085000 1160.435000 0.085000 ;
      RECT 1160.265000  2.635000 1160.435000 2.805000 ;
      RECT 1160.725000 -0.085000 1160.895000 0.085000 ;
      RECT 1160.725000  2.635000 1160.895000 2.805000 ;
      RECT 1161.185000 -0.085000 1161.355000 0.085000 ;
      RECT 1161.185000  2.635000 1161.355000 2.805000 ;
      RECT 1161.645000 -0.085000 1161.815000 0.085000 ;
      RECT 1161.645000  2.635000 1161.815000 2.805000 ;
      RECT 1162.105000 -0.085000 1162.275000 0.085000 ;
      RECT 1162.105000  2.635000 1162.275000 2.805000 ;
      RECT 1162.565000 -0.085000 1162.735000 0.085000 ;
      RECT 1162.565000  2.635000 1162.735000 2.805000 ;
      RECT 1163.025000 -0.085000 1163.195000 0.085000 ;
      RECT 1163.025000  2.635000 1163.195000 2.805000 ;
      RECT 1163.485000 -0.085000 1163.655000 0.085000 ;
      RECT 1163.485000  2.635000 1163.655000 2.805000 ;
      RECT 1163.945000 -0.085000 1164.115000 0.085000 ;
      RECT 1163.945000  2.635000 1164.115000 2.805000 ;
      RECT 1164.405000 -0.085000 1164.575000 0.085000 ;
      RECT 1164.405000  2.635000 1164.575000 2.805000 ;
      RECT 1164.865000 -0.085000 1165.035000 0.085000 ;
      RECT 1164.865000  2.635000 1165.035000 2.805000 ;
      RECT 1165.325000 -0.085000 1165.495000 0.085000 ;
      RECT 1165.325000  2.635000 1165.495000 2.805000 ;
      RECT 1165.785000 -0.085000 1165.955000 0.085000 ;
      RECT 1165.785000  2.635000 1165.955000 2.805000 ;
      RECT 1166.245000 -0.085000 1166.415000 0.085000 ;
      RECT 1166.245000  2.635000 1166.415000 2.805000 ;
      RECT 1166.705000 -0.085000 1166.875000 0.085000 ;
      RECT 1166.705000  2.635000 1166.875000 2.805000 ;
      RECT 1167.165000 -0.085000 1167.335000 0.085000 ;
      RECT 1167.165000  2.635000 1167.335000 2.805000 ;
      RECT 1167.625000 -0.085000 1167.795000 0.085000 ;
      RECT 1167.625000  2.635000 1167.795000 2.805000 ;
      RECT 1168.085000 -0.085000 1168.255000 0.085000 ;
      RECT 1168.085000  2.635000 1168.255000 2.805000 ;
      RECT 1168.545000 -0.085000 1168.715000 0.085000 ;
      RECT 1168.545000  2.635000 1168.715000 2.805000 ;
      RECT 1169.005000 -0.085000 1169.175000 0.085000 ;
      RECT 1169.005000  2.635000 1169.175000 2.805000 ;
      RECT 1169.465000 -0.085000 1169.635000 0.085000 ;
      RECT 1169.465000  2.635000 1169.635000 2.805000 ;
      RECT 1169.925000 -0.085000 1170.095000 0.085000 ;
      RECT 1169.925000  2.635000 1170.095000 2.805000 ;
      RECT 1170.385000 -0.085000 1170.555000 0.085000 ;
      RECT 1170.385000  2.635000 1170.555000 2.805000 ;
      RECT 1170.845000 -0.085000 1171.015000 0.085000 ;
      RECT 1170.845000  2.635000 1171.015000 2.805000 ;
      RECT 1171.305000 -0.085000 1171.475000 0.085000 ;
      RECT 1171.305000  2.635000 1171.475000 2.805000 ;
      RECT 1171.765000 -0.085000 1171.935000 0.085000 ;
      RECT 1171.765000  2.635000 1171.935000 2.805000 ;
      RECT 1172.225000 -0.085000 1172.395000 0.085000 ;
      RECT 1172.225000  2.635000 1172.395000 2.805000 ;
      RECT 1172.685000 -0.085000 1172.855000 0.085000 ;
      RECT 1172.685000  2.635000 1172.855000 2.805000 ;
      RECT 1173.145000 -0.085000 1173.315000 0.085000 ;
      RECT 1173.145000  2.635000 1173.315000 2.805000 ;
      RECT 1173.605000 -0.085000 1173.775000 0.085000 ;
      RECT 1173.605000  2.635000 1173.775000 2.805000 ;
      RECT 1174.065000 -0.085000 1174.235000 0.085000 ;
      RECT 1174.065000  2.635000 1174.235000 2.805000 ;
      RECT 1174.525000 -0.085000 1174.695000 0.085000 ;
      RECT 1174.525000  2.635000 1174.695000 2.805000 ;
      RECT 1174.985000 -0.085000 1175.155000 0.085000 ;
      RECT 1174.985000  2.635000 1175.155000 2.805000 ;
      RECT 1175.445000 -0.085000 1175.615000 0.085000 ;
      RECT 1175.445000  2.635000 1175.615000 2.805000 ;
      RECT 1175.905000 -0.085000 1176.075000 0.085000 ;
      RECT 1175.905000  2.635000 1176.075000 2.805000 ;
      RECT 1176.365000 -0.085000 1176.535000 0.085000 ;
      RECT 1176.365000  2.635000 1176.535000 2.805000 ;
      RECT 1176.825000 -0.085000 1176.995000 0.085000 ;
      RECT 1176.825000  2.635000 1176.995000 2.805000 ;
      RECT 1177.285000 -0.085000 1177.455000 0.085000 ;
      RECT 1177.285000  2.635000 1177.455000 2.805000 ;
      RECT 1177.745000 -0.085000 1177.915000 0.085000 ;
      RECT 1177.745000  2.635000 1177.915000 2.805000 ;
      RECT 1178.205000 -0.085000 1178.375000 0.085000 ;
      RECT 1178.205000  2.635000 1178.375000 2.805000 ;
      RECT 1178.665000 -0.085000 1178.835000 0.085000 ;
      RECT 1178.665000  2.635000 1178.835000 2.805000 ;
      RECT 1179.125000 -0.085000 1179.295000 0.085000 ;
      RECT 1179.125000  2.635000 1179.295000 2.805000 ;
      RECT 1179.585000 -0.085000 1179.755000 0.085000 ;
      RECT 1179.585000  2.635000 1179.755000 2.805000 ;
      RECT 1180.045000 -0.085000 1180.215000 0.085000 ;
      RECT 1180.045000  2.635000 1180.215000 2.805000 ;
      RECT 1180.505000 -0.085000 1180.675000 0.085000 ;
      RECT 1180.505000  2.635000 1180.675000 2.805000 ;
      RECT 1180.965000 -0.085000 1181.135000 0.085000 ;
      RECT 1180.965000  2.635000 1181.135000 2.805000 ;
      RECT 1181.425000 -0.085000 1181.595000 0.085000 ;
      RECT 1181.425000  2.635000 1181.595000 2.805000 ;
      RECT 1181.885000 -0.085000 1182.055000 0.085000 ;
      RECT 1181.885000  2.635000 1182.055000 2.805000 ;
      RECT 1182.345000 -0.085000 1182.515000 0.085000 ;
      RECT 1182.345000  2.635000 1182.515000 2.805000 ;
      RECT 1182.805000 -0.085000 1182.975000 0.085000 ;
      RECT 1182.805000  2.635000 1182.975000 2.805000 ;
      RECT 1183.265000 -0.085000 1183.435000 0.085000 ;
      RECT 1183.265000  2.635000 1183.435000 2.805000 ;
      RECT 1183.725000 -0.085000 1183.895000 0.085000 ;
      RECT 1183.725000  2.635000 1183.895000 2.805000 ;
      RECT 1184.185000 -0.085000 1184.355000 0.085000 ;
      RECT 1184.185000  2.635000 1184.355000 2.805000 ;
      RECT 1184.645000 -0.085000 1184.815000 0.085000 ;
      RECT 1184.645000  2.635000 1184.815000 2.805000 ;
      RECT 1185.105000 -0.085000 1185.275000 0.085000 ;
      RECT 1185.105000  2.635000 1185.275000 2.805000 ;
      RECT 1185.565000 -0.085000 1185.735000 0.085000 ;
      RECT 1185.565000  2.635000 1185.735000 2.805000 ;
      RECT 1186.025000 -0.085000 1186.195000 0.085000 ;
      RECT 1186.025000  2.635000 1186.195000 2.805000 ;
      RECT 1186.485000 -0.085000 1186.655000 0.085000 ;
      RECT 1186.485000  2.635000 1186.655000 2.805000 ;
      RECT 1186.945000 -0.085000 1187.115000 0.085000 ;
      RECT 1186.945000  2.635000 1187.115000 2.805000 ;
      RECT 1187.405000 -0.085000 1187.575000 0.085000 ;
      RECT 1187.405000  2.635000 1187.575000 2.805000 ;
      RECT 1187.865000 -0.085000 1188.035000 0.085000 ;
      RECT 1187.865000  2.635000 1188.035000 2.805000 ;
      RECT 1188.325000 -0.085000 1188.495000 0.085000 ;
      RECT 1188.325000  2.635000 1188.495000 2.805000 ;
      RECT 1188.575000  1.435000 1188.745000 1.605000 ;
      RECT 1188.785000 -0.085000 1188.955000 0.085000 ;
      RECT 1188.785000  2.635000 1188.955000 2.805000 ;
      RECT 1189.245000 -0.085000 1189.415000 0.085000 ;
      RECT 1189.245000  2.635000 1189.415000 2.805000 ;
      RECT 1189.705000 -0.085000 1189.875000 0.085000 ;
      RECT 1189.705000  2.635000 1189.875000 2.805000 ;
      RECT 1190.165000 -0.085000 1190.335000 0.085000 ;
      RECT 1190.165000  2.635000 1190.335000 2.805000 ;
      RECT 1190.625000 -0.085000 1190.795000 0.085000 ;
      RECT 1190.625000  2.635000 1190.795000 2.805000 ;
      RECT 1191.085000 -0.085000 1191.255000 0.085000 ;
      RECT 1191.085000  2.635000 1191.255000 2.805000 ;
      RECT 1191.545000 -0.085000 1191.715000 0.085000 ;
      RECT 1191.545000  2.635000 1191.715000 2.805000 ;
      RECT 1191.605000  1.445000 1191.775000 1.615000 ;
      RECT 1192.005000 -0.085000 1192.175000 0.085000 ;
      RECT 1192.005000  2.635000 1192.175000 2.805000 ;
      RECT 1192.465000 -0.085000 1192.635000 0.085000 ;
      RECT 1192.465000  2.635000 1192.635000 2.805000 ;
      RECT 1192.925000 -0.085000 1193.095000 0.085000 ;
      RECT 1192.925000  2.635000 1193.095000 2.805000 ;
      RECT 1193.385000 -0.085000 1193.555000 0.085000 ;
      RECT 1193.385000  2.635000 1193.555000 2.805000 ;
      RECT 1193.845000 -0.085000 1194.015000 0.085000 ;
      RECT 1193.845000  2.635000 1194.015000 2.805000 ;
      RECT 1194.305000 -0.085000 1194.475000 0.085000 ;
      RECT 1194.305000  2.635000 1194.475000 2.805000 ;
      RECT 1194.765000 -0.085000 1194.935000 0.085000 ;
      RECT 1194.765000  2.635000 1194.935000 2.805000 ;
      RECT 1195.225000 -0.085000 1195.395000 0.085000 ;
      RECT 1195.225000  2.635000 1195.395000 2.805000 ;
      RECT 1195.685000 -0.085000 1195.855000 0.085000 ;
      RECT 1195.685000  2.635000 1195.855000 2.805000 ;
      RECT 1196.145000 -0.085000 1196.315000 0.085000 ;
      RECT 1196.145000  2.635000 1196.315000 2.805000 ;
      RECT 1196.605000 -0.085000 1196.775000 0.085000 ;
      RECT 1196.605000  2.635000 1196.775000 2.805000 ;
      RECT 1197.065000 -0.085000 1197.235000 0.085000 ;
      RECT 1197.065000  2.635000 1197.235000 2.805000 ;
      RECT 1197.525000 -0.085000 1197.695000 0.085000 ;
      RECT 1197.525000  2.635000 1197.695000 2.805000 ;
      RECT 1197.985000 -0.085000 1198.155000 0.085000 ;
      RECT 1197.985000  2.635000 1198.155000 2.805000 ;
      RECT 1198.445000 -0.085000 1198.615000 0.085000 ;
      RECT 1198.445000  2.635000 1198.615000 2.805000 ;
      RECT 1198.905000 -0.085000 1199.075000 0.085000 ;
      RECT 1198.905000  2.635000 1199.075000 2.805000 ;
      RECT 1199.365000 -0.085000 1199.535000 0.085000 ;
      RECT 1199.365000  2.635000 1199.535000 2.805000 ;
      RECT 1199.825000 -0.085000 1199.995000 0.085000 ;
      RECT 1199.825000  2.635000 1199.995000 2.805000 ;
      RECT 1200.285000 -0.085000 1200.455000 0.085000 ;
      RECT 1200.285000  2.635000 1200.455000 2.805000 ;
      RECT 1200.745000 -0.085000 1200.915000 0.085000 ;
      RECT 1200.745000  2.635000 1200.915000 2.805000 ;
      RECT 1201.205000 -0.085000 1201.375000 0.085000 ;
      RECT 1201.205000  2.635000 1201.375000 2.805000 ;
      RECT 1201.665000 -0.085000 1201.835000 0.085000 ;
      RECT 1201.665000  2.635000 1201.835000 2.805000 ;
      RECT 1202.125000 -0.085000 1202.295000 0.085000 ;
      RECT 1202.125000  2.635000 1202.295000 2.805000 ;
      RECT 1202.585000 -0.085000 1202.755000 0.085000 ;
      RECT 1202.585000  2.635000 1202.755000 2.805000 ;
      RECT 1203.045000 -0.085000 1203.215000 0.085000 ;
      RECT 1203.045000  2.635000 1203.215000 2.805000 ;
      RECT 1203.505000 -0.085000 1203.675000 0.085000 ;
      RECT 1203.505000  2.635000 1203.675000 2.805000 ;
      RECT 1203.965000 -0.085000 1204.135000 0.085000 ;
      RECT 1203.965000  2.635000 1204.135000 2.805000 ;
      RECT 1204.425000 -0.085000 1204.595000 0.085000 ;
      RECT 1204.425000  2.635000 1204.595000 2.805000 ;
      RECT 1204.885000 -0.085000 1205.055000 0.085000 ;
      RECT 1204.885000  2.635000 1205.055000 2.805000 ;
      RECT 1205.345000 -0.085000 1205.515000 0.085000 ;
      RECT 1205.345000  2.635000 1205.515000 2.805000 ;
      RECT 1205.805000 -0.085000 1205.975000 0.085000 ;
      RECT 1205.805000  2.635000 1205.975000 2.805000 ;
      RECT 1206.265000 -0.085000 1206.435000 0.085000 ;
      RECT 1206.265000  2.635000 1206.435000 2.805000 ;
      RECT 1206.725000 -0.085000 1206.895000 0.085000 ;
      RECT 1206.725000  2.635000 1206.895000 2.805000 ;
      RECT 1207.185000 -0.085000 1207.355000 0.085000 ;
      RECT 1207.185000  2.635000 1207.355000 2.805000 ;
      RECT 1207.645000 -0.085000 1207.815000 0.085000 ;
      RECT 1207.645000  2.635000 1207.815000 2.805000 ;
      RECT 1208.105000 -0.085000 1208.275000 0.085000 ;
      RECT 1208.105000  2.635000 1208.275000 2.805000 ;
      RECT 1208.565000 -0.085000 1208.735000 0.085000 ;
      RECT 1208.565000  2.635000 1208.735000 2.805000 ;
      RECT 1209.025000 -0.085000 1209.195000 0.085000 ;
      RECT 1209.025000  2.635000 1209.195000 2.805000 ;
      RECT 1209.485000 -0.085000 1209.655000 0.085000 ;
      RECT 1209.485000  2.635000 1209.655000 2.805000 ;
      RECT 1209.945000 -0.085000 1210.115000 0.085000 ;
      RECT 1209.945000  2.635000 1210.115000 2.805000 ;
      RECT 1210.405000 -0.085000 1210.575000 0.085000 ;
      RECT 1210.405000  2.635000 1210.575000 2.805000 ;
      RECT 1210.865000 -0.085000 1211.035000 0.085000 ;
      RECT 1210.865000  2.635000 1211.035000 2.805000 ;
      RECT 1211.325000 -0.085000 1211.495000 0.085000 ;
      RECT 1211.325000  2.635000 1211.495000 2.805000 ;
      RECT 1211.785000 -0.085000 1211.955000 0.085000 ;
      RECT 1211.785000  2.635000 1211.955000 2.805000 ;
      RECT 1212.245000 -0.085000 1212.415000 0.085000 ;
      RECT 1212.245000  2.635000 1212.415000 2.805000 ;
      RECT 1212.705000 -0.085000 1212.875000 0.085000 ;
      RECT 1212.705000  2.635000 1212.875000 2.805000 ;
      RECT 1213.165000 -0.085000 1213.335000 0.085000 ;
      RECT 1213.165000  2.635000 1213.335000 2.805000 ;
      RECT 1213.625000 -0.085000 1213.795000 0.085000 ;
      RECT 1213.625000  2.635000 1213.795000 2.805000 ;
      RECT 1214.085000 -0.085000 1214.255000 0.085000 ;
      RECT 1214.085000  2.635000 1214.255000 2.805000 ;
      RECT 1214.545000 -0.085000 1214.715000 0.085000 ;
      RECT 1214.545000  2.635000 1214.715000 2.805000 ;
      RECT 1215.005000 -0.085000 1215.175000 0.085000 ;
      RECT 1215.005000  2.635000 1215.175000 2.805000 ;
      RECT 1215.465000 -0.085000 1215.635000 0.085000 ;
      RECT 1215.465000  2.635000 1215.635000 2.805000 ;
      RECT 1215.925000 -0.085000 1216.095000 0.085000 ;
      RECT 1215.925000  2.635000 1216.095000 2.805000 ;
      RECT 1216.385000 -0.085000 1216.555000 0.085000 ;
      RECT 1216.385000  2.635000 1216.555000 2.805000 ;
      RECT 1216.845000 -0.085000 1217.015000 0.085000 ;
      RECT 1216.845000  2.635000 1217.015000 2.805000 ;
      RECT 1217.305000 -0.085000 1217.475000 0.085000 ;
      RECT 1217.305000  2.635000 1217.475000 2.805000 ;
      RECT 1217.765000 -0.085000 1217.935000 0.085000 ;
      RECT 1217.765000  2.635000 1217.935000 2.805000 ;
      RECT 1218.225000 -0.085000 1218.395000 0.085000 ;
      RECT 1218.225000  2.635000 1218.395000 2.805000 ;
      RECT 1218.685000 -0.085000 1218.855000 0.085000 ;
      RECT 1218.685000  2.635000 1218.855000 2.805000 ;
      RECT 1219.145000 -0.085000 1219.315000 0.085000 ;
      RECT 1219.145000  2.635000 1219.315000 2.805000 ;
      RECT 1219.605000 -0.085000 1219.775000 0.085000 ;
      RECT 1219.605000  2.635000 1219.775000 2.805000 ;
      RECT 1220.065000 -0.085000 1220.235000 0.085000 ;
      RECT 1220.065000  2.635000 1220.235000 2.805000 ;
      RECT 1220.525000 -0.085000 1220.695000 0.085000 ;
      RECT 1220.525000  2.635000 1220.695000 2.805000 ;
      RECT 1220.985000 -0.085000 1221.155000 0.085000 ;
      RECT 1220.985000  2.635000 1221.155000 2.805000 ;
      RECT 1221.445000 -0.085000 1221.615000 0.085000 ;
      RECT 1221.445000  2.635000 1221.615000 2.805000 ;
      RECT 1221.905000 -0.085000 1222.075000 0.085000 ;
      RECT 1221.905000  2.635000 1222.075000 2.805000 ;
      RECT 1222.365000 -0.085000 1222.535000 0.085000 ;
      RECT 1222.365000  2.635000 1222.535000 2.805000 ;
      RECT 1222.825000 -0.085000 1222.995000 0.085000 ;
      RECT 1222.825000  2.635000 1222.995000 2.805000 ;
      RECT 1223.285000 -0.085000 1223.455000 0.085000 ;
      RECT 1223.285000  2.635000 1223.455000 2.805000 ;
      RECT 1223.745000 -0.085000 1223.915000 0.085000 ;
      RECT 1223.745000  2.635000 1223.915000 2.805000 ;
      RECT 1224.205000 -0.085000 1224.375000 0.085000 ;
      RECT 1224.205000  2.635000 1224.375000 2.805000 ;
      RECT 1224.665000 -0.085000 1224.835000 0.085000 ;
      RECT 1224.665000  2.635000 1224.835000 2.805000 ;
      RECT 1225.125000 -0.085000 1225.295000 0.085000 ;
      RECT 1225.125000  2.635000 1225.295000 2.805000 ;
      RECT 1225.585000 -0.085000 1225.755000 0.085000 ;
      RECT 1225.585000  2.635000 1225.755000 2.805000 ;
      RECT 1226.045000 -0.085000 1226.215000 0.085000 ;
      RECT 1226.045000  2.635000 1226.215000 2.805000 ;
      RECT 1226.505000 -0.085000 1226.675000 0.085000 ;
      RECT 1226.505000  2.635000 1226.675000 2.805000 ;
      RECT 1226.965000 -0.085000 1227.135000 0.085000 ;
      RECT 1226.965000  2.635000 1227.135000 2.805000 ;
      RECT 1227.425000 -0.085000 1227.595000 0.085000 ;
      RECT 1227.425000  2.635000 1227.595000 2.805000 ;
      RECT 1227.885000 -0.085000 1228.055000 0.085000 ;
      RECT 1227.885000  2.635000 1228.055000 2.805000 ;
      RECT 1228.345000 -0.085000 1228.515000 0.085000 ;
      RECT 1228.345000  2.635000 1228.515000 2.805000 ;
      RECT 1228.805000 -0.085000 1228.975000 0.085000 ;
      RECT 1228.805000  2.635000 1228.975000 2.805000 ;
      RECT 1229.265000 -0.085000 1229.435000 0.085000 ;
      RECT 1229.265000  2.635000 1229.435000 2.805000 ;
      RECT 1229.725000 -0.085000 1229.895000 0.085000 ;
      RECT 1229.725000  2.635000 1229.895000 2.805000 ;
      RECT 1230.185000 -0.085000 1230.355000 0.085000 ;
      RECT 1230.185000  2.635000 1230.355000 2.805000 ;
      RECT 1230.645000 -0.085000 1230.815000 0.085000 ;
      RECT 1230.645000  2.635000 1230.815000 2.805000 ;
      RECT 1231.105000 -0.085000 1231.275000 0.085000 ;
      RECT 1231.105000  2.635000 1231.275000 2.805000 ;
      RECT 1231.565000 -0.085000 1231.735000 0.085000 ;
      RECT 1231.565000  2.635000 1231.735000 2.805000 ;
      RECT 1232.025000 -0.085000 1232.195000 0.085000 ;
      RECT 1232.025000  2.635000 1232.195000 2.805000 ;
      RECT 1232.485000 -0.085000 1232.655000 0.085000 ;
      RECT 1232.485000  2.635000 1232.655000 2.805000 ;
      RECT 1232.945000 -0.085000 1233.115000 0.085000 ;
      RECT 1232.945000  2.635000 1233.115000 2.805000 ;
      RECT 1233.405000 -0.085000 1233.575000 0.085000 ;
      RECT 1233.405000  2.635000 1233.575000 2.805000 ;
      RECT 1233.865000 -0.085000 1234.035000 0.085000 ;
      RECT 1233.865000  2.635000 1234.035000 2.805000 ;
      RECT 1234.325000 -0.085000 1234.495000 0.085000 ;
      RECT 1234.325000  2.635000 1234.495000 2.805000 ;
      RECT 1234.785000 -0.085000 1234.955000 0.085000 ;
      RECT 1234.785000  2.635000 1234.955000 2.805000 ;
      RECT 1235.245000 -0.085000 1235.415000 0.085000 ;
      RECT 1235.245000  2.635000 1235.415000 2.805000 ;
      RECT 1235.705000 -0.085000 1235.875000 0.085000 ;
      RECT 1235.705000  2.635000 1235.875000 2.805000 ;
      RECT 1236.165000 -0.085000 1236.335000 0.085000 ;
      RECT 1236.165000  2.635000 1236.335000 2.805000 ;
      RECT 1236.625000 -0.085000 1236.795000 0.085000 ;
      RECT 1236.625000  2.635000 1236.795000 2.805000 ;
      RECT 1237.085000 -0.085000 1237.255000 0.085000 ;
      RECT 1237.085000  2.635000 1237.255000 2.805000 ;
      RECT 1237.545000 -0.085000 1237.715000 0.085000 ;
      RECT 1237.545000  2.635000 1237.715000 2.805000 ;
      RECT 1238.005000 -0.085000 1238.175000 0.085000 ;
      RECT 1238.005000  2.635000 1238.175000 2.805000 ;
      RECT 1238.465000 -0.085000 1238.635000 0.085000 ;
      RECT 1238.465000  2.635000 1238.635000 2.805000 ;
      RECT 1238.925000 -0.085000 1239.095000 0.085000 ;
      RECT 1238.925000  2.635000 1239.095000 2.805000 ;
      RECT 1239.385000 -0.085000 1239.555000 0.085000 ;
      RECT 1239.385000  2.635000 1239.555000 2.805000 ;
      RECT 1239.845000 -0.085000 1240.015000 0.085000 ;
      RECT 1239.845000  2.635000 1240.015000 2.805000 ;
      RECT 1240.305000 -0.085000 1240.475000 0.085000 ;
      RECT 1240.305000  2.635000 1240.475000 2.805000 ;
      RECT 1240.765000 -0.085000 1240.935000 0.085000 ;
      RECT 1240.765000  2.635000 1240.935000 2.805000 ;
      RECT 1241.225000 -0.085000 1241.395000 0.085000 ;
      RECT 1241.225000  2.635000 1241.395000 2.805000 ;
      RECT 1241.685000 -0.085000 1241.855000 0.085000 ;
      RECT 1241.685000  2.635000 1241.855000 2.805000 ;
      RECT 1242.145000 -0.085000 1242.315000 0.085000 ;
      RECT 1242.145000  2.635000 1242.315000 2.805000 ;
      RECT 1242.605000 -0.085000 1242.775000 0.085000 ;
      RECT 1242.605000  2.635000 1242.775000 2.805000 ;
      RECT 1243.065000 -0.085000 1243.235000 0.085000 ;
      RECT 1243.065000  2.635000 1243.235000 2.805000 ;
      RECT 1243.525000 -0.085000 1243.695000 0.085000 ;
      RECT 1243.525000  2.635000 1243.695000 2.805000 ;
      RECT 1243.985000 -0.085000 1244.155000 0.085000 ;
      RECT 1243.985000  2.635000 1244.155000 2.805000 ;
      RECT 1244.445000 -0.085000 1244.615000 0.085000 ;
      RECT 1244.445000  2.635000 1244.615000 2.805000 ;
      RECT 1244.905000 -0.085000 1245.075000 0.085000 ;
      RECT 1244.905000  2.635000 1245.075000 2.805000 ;
      RECT 1245.365000 -0.085000 1245.535000 0.085000 ;
      RECT 1245.365000  2.635000 1245.535000 2.805000 ;
      RECT 1245.825000 -0.085000 1245.995000 0.085000 ;
      RECT 1245.825000  2.635000 1245.995000 2.805000 ;
      RECT 1246.285000 -0.085000 1246.455000 0.085000 ;
      RECT 1246.285000  2.635000 1246.455000 2.805000 ;
      RECT 1246.745000 -0.085000 1246.915000 0.085000 ;
      RECT 1246.745000  2.635000 1246.915000 2.805000 ;
      RECT 1247.205000 -0.085000 1247.375000 0.085000 ;
      RECT 1247.205000  2.635000 1247.375000 2.805000 ;
      RECT 1247.665000 -0.085000 1247.835000 0.085000 ;
      RECT 1247.665000  2.635000 1247.835000 2.805000 ;
      RECT 1248.125000 -0.085000 1248.295000 0.085000 ;
      RECT 1248.125000  2.635000 1248.295000 2.805000 ;
      RECT 1248.585000 -0.085000 1248.755000 0.085000 ;
      RECT 1248.585000  2.635000 1248.755000 2.805000 ;
      RECT 1249.045000 -0.085000 1249.215000 0.085000 ;
      RECT 1249.045000  2.635000 1249.215000 2.805000 ;
      RECT 1249.505000 -0.085000 1249.675000 0.085000 ;
      RECT 1249.505000  2.635000 1249.675000 2.805000 ;
      RECT 1249.965000 -0.085000 1250.135000 0.085000 ;
      RECT 1249.965000  2.635000 1250.135000 2.805000 ;
      RECT 1250.425000 -0.085000 1250.595000 0.085000 ;
      RECT 1250.425000  2.635000 1250.595000 2.805000 ;
      RECT 1250.885000 -0.085000 1251.055000 0.085000 ;
      RECT 1250.885000  2.635000 1251.055000 2.805000 ;
      RECT 1251.345000 -0.085000 1251.515000 0.085000 ;
      RECT 1251.345000  2.635000 1251.515000 2.805000 ;
      RECT 1251.805000 -0.085000 1251.975000 0.085000 ;
      RECT 1251.805000  2.635000 1251.975000 2.805000 ;
      RECT 1252.265000 -0.085000 1252.435000 0.085000 ;
      RECT 1252.265000  2.635000 1252.435000 2.805000 ;
      RECT 1252.725000 -0.085000 1252.895000 0.085000 ;
      RECT 1252.725000  2.635000 1252.895000 2.805000 ;
      RECT 1253.185000 -0.085000 1253.355000 0.085000 ;
      RECT 1253.185000  2.635000 1253.355000 2.805000 ;
      RECT 1253.645000 -0.085000 1253.815000 0.085000 ;
      RECT 1253.645000  2.635000 1253.815000 2.805000 ;
      RECT 1254.105000 -0.085000 1254.275000 0.085000 ;
      RECT 1254.105000  2.635000 1254.275000 2.805000 ;
      RECT 1254.565000 -0.085000 1254.735000 0.085000 ;
      RECT 1254.565000  2.635000 1254.735000 2.805000 ;
      RECT 1255.025000 -0.085000 1255.195000 0.085000 ;
      RECT 1255.025000  2.635000 1255.195000 2.805000 ;
      RECT 1255.485000 -0.085000 1255.655000 0.085000 ;
      RECT 1255.485000  2.635000 1255.655000 2.805000 ;
      RECT 1255.945000 -0.085000 1256.115000 0.085000 ;
      RECT 1255.945000  2.635000 1256.115000 2.805000 ;
      RECT 1256.405000 -0.085000 1256.575000 0.085000 ;
      RECT 1256.405000  2.635000 1256.575000 2.805000 ;
      RECT 1256.865000 -0.085000 1257.035000 0.085000 ;
      RECT 1256.865000  2.635000 1257.035000 2.805000 ;
      RECT 1257.325000 -0.085000 1257.495000 0.085000 ;
      RECT 1257.325000  2.635000 1257.495000 2.805000 ;
      RECT 1257.785000 -0.085000 1257.955000 0.085000 ;
      RECT 1257.785000  2.635000 1257.955000 2.805000 ;
      RECT 1258.245000 -0.085000 1258.415000 0.085000 ;
      RECT 1258.245000  2.635000 1258.415000 2.805000 ;
      RECT 1258.705000 -0.085000 1258.875000 0.085000 ;
      RECT 1258.705000  2.635000 1258.875000 2.805000 ;
      RECT 1259.165000 -0.085000 1259.335000 0.085000 ;
      RECT 1259.165000  2.635000 1259.335000 2.805000 ;
      RECT 1259.625000 -0.085000 1259.795000 0.085000 ;
      RECT 1259.625000  2.635000 1259.795000 2.805000 ;
      RECT 1260.085000 -0.085000 1260.255000 0.085000 ;
      RECT 1260.085000  2.635000 1260.255000 2.805000 ;
      RECT 1260.545000 -0.085000 1260.715000 0.085000 ;
      RECT 1260.545000  2.635000 1260.715000 2.805000 ;
      RECT 1261.005000 -0.085000 1261.175000 0.085000 ;
      RECT 1261.005000  2.635000 1261.175000 2.805000 ;
      RECT 1261.465000 -0.085000 1261.635000 0.085000 ;
      RECT 1261.465000  2.635000 1261.635000 2.805000 ;
      RECT 1261.925000 -0.085000 1262.095000 0.085000 ;
      RECT 1261.925000  2.635000 1262.095000 2.805000 ;
      RECT 1262.385000 -0.085000 1262.555000 0.085000 ;
      RECT 1262.385000  2.635000 1262.555000 2.805000 ;
      RECT 1262.845000 -0.085000 1263.015000 0.085000 ;
      RECT 1262.845000  2.635000 1263.015000 2.805000 ;
      RECT 1263.305000 -0.085000 1263.475000 0.085000 ;
      RECT 1263.305000  2.635000 1263.475000 2.805000 ;
      RECT 1263.765000 -0.085000 1263.935000 0.085000 ;
      RECT 1263.765000  2.635000 1263.935000 2.805000 ;
      RECT 1264.225000 -0.085000 1264.395000 0.085000 ;
      RECT 1264.225000  2.635000 1264.395000 2.805000 ;
      RECT 1264.685000 -0.085000 1264.855000 0.085000 ;
      RECT 1264.685000  2.635000 1264.855000 2.805000 ;
      RECT 1265.145000 -0.085000 1265.315000 0.085000 ;
      RECT 1265.145000  2.635000 1265.315000 2.805000 ;
      RECT 1265.605000 -0.085000 1265.775000 0.085000 ;
      RECT 1265.605000  2.635000 1265.775000 2.805000 ;
      RECT 1266.065000 -0.085000 1266.235000 0.085000 ;
      RECT 1266.065000  2.635000 1266.235000 2.805000 ;
      RECT 1266.525000 -0.085000 1266.695000 0.085000 ;
      RECT 1266.525000  2.635000 1266.695000 2.805000 ;
      RECT 1266.985000 -0.085000 1267.155000 0.085000 ;
      RECT 1266.985000  2.635000 1267.155000 2.805000 ;
      RECT 1267.445000 -0.085000 1267.615000 0.085000 ;
      RECT 1267.445000  2.635000 1267.615000 2.805000 ;
      RECT 1267.905000 -0.085000 1268.075000 0.085000 ;
      RECT 1267.905000  2.635000 1268.075000 2.805000 ;
      RECT 1268.365000 -0.085000 1268.535000 0.085000 ;
      RECT 1268.365000  2.635000 1268.535000 2.805000 ;
      RECT 1268.825000 -0.085000 1268.995000 0.085000 ;
      RECT 1268.825000  2.635000 1268.995000 2.805000 ;
      RECT 1269.745000 -0.085000 1269.915000 0.085000 ;
      RECT 1269.745000  2.635000 1269.915000 2.805000 ;
      RECT 1270.205000 -0.085000 1270.375000 0.085000 ;
      RECT 1270.205000  2.635000 1270.375000 2.805000 ;
      RECT 1270.665000 -0.085000 1270.835000 0.085000 ;
      RECT 1270.665000  2.635000 1270.835000 2.805000 ;
      RECT 1271.125000 -0.085000 1271.295000 0.085000 ;
      RECT 1271.125000  2.635000 1271.295000 2.805000 ;
      RECT 1271.585000 -0.085000 1271.755000 0.085000 ;
      RECT 1271.585000  2.635000 1271.755000 2.805000 ;
      RECT 1272.045000 -0.085000 1272.215000 0.085000 ;
      RECT 1272.045000  2.635000 1272.215000 2.805000 ;
      RECT 1272.505000 -0.085000 1272.675000 0.085000 ;
      RECT 1272.505000  2.635000 1272.675000 2.805000 ;
      RECT 1272.965000 -0.085000 1273.135000 0.085000 ;
      RECT 1272.965000  2.635000 1273.135000 2.805000 ;
      RECT 1273.425000 -0.085000 1273.595000 0.085000 ;
      RECT 1273.425000  2.635000 1273.595000 2.805000 ;
      RECT 1273.885000 -0.085000 1274.055000 0.085000 ;
      RECT 1273.885000  2.635000 1274.055000 2.805000 ;
      RECT 1274.345000 -0.085000 1274.515000 0.085000 ;
      RECT 1274.345000  2.635000 1274.515000 2.805000 ;
      RECT 1274.805000 -0.085000 1274.975000 0.085000 ;
      RECT 1274.805000  2.635000 1274.975000 2.805000 ;
      RECT 1275.265000 -0.085000 1275.435000 0.085000 ;
      RECT 1275.265000  2.635000 1275.435000 2.805000 ;
      RECT 1275.725000 -0.085000 1275.895000 0.085000 ;
      RECT 1275.725000  2.635000 1275.895000 2.805000 ;
      RECT 1276.185000 -0.085000 1276.355000 0.085000 ;
      RECT 1276.185000  2.635000 1276.355000 2.805000 ;
      RECT 1276.645000 -0.085000 1276.815000 0.085000 ;
      RECT 1276.645000  2.635000 1276.815000 2.805000 ;
      RECT 1277.105000 -0.085000 1277.275000 0.085000 ;
      RECT 1277.105000  2.635000 1277.275000 2.805000 ;
      RECT 1277.565000 -0.085000 1277.735000 0.085000 ;
      RECT 1277.565000  2.635000 1277.735000 2.805000 ;
      RECT 1278.025000 -0.085000 1278.195000 0.085000 ;
      RECT 1278.025000  2.635000 1278.195000 2.805000 ;
      RECT 1278.485000 -0.085000 1278.655000 0.085000 ;
      RECT 1278.485000  2.635000 1278.655000 2.805000 ;
      RECT 1278.945000 -0.085000 1279.115000 0.085000 ;
      RECT 1278.945000  2.635000 1279.115000 2.805000 ;
      RECT 1279.405000 -0.085000 1279.575000 0.085000 ;
      RECT 1279.405000  2.635000 1279.575000 2.805000 ;
      RECT 1279.865000 -0.085000 1280.035000 0.085000 ;
      RECT 1279.865000  2.635000 1280.035000 2.805000 ;
      RECT 1280.325000 -0.085000 1280.495000 0.085000 ;
      RECT 1280.325000  2.635000 1280.495000 2.805000 ;
      RECT 1280.785000 -0.085000 1280.955000 0.085000 ;
      RECT 1280.785000  2.635000 1280.955000 2.805000 ;
      RECT 1281.245000 -0.085000 1281.415000 0.085000 ;
      RECT 1281.245000  2.635000 1281.415000 2.805000 ;
      RECT 1281.705000 -0.085000 1281.875000 0.085000 ;
      RECT 1281.705000  2.635000 1281.875000 2.805000 ;
      RECT 1282.165000 -0.085000 1282.335000 0.085000 ;
      RECT 1282.165000  2.635000 1282.335000 2.805000 ;
      RECT 1282.625000 -0.085000 1282.795000 0.085000 ;
      RECT 1282.625000  2.635000 1282.795000 2.805000 ;
      RECT 1283.085000 -0.085000 1283.255000 0.085000 ;
      RECT 1283.085000  2.635000 1283.255000 2.805000 ;
      RECT 1283.545000 -0.085000 1283.715000 0.085000 ;
      RECT 1283.545000  2.635000 1283.715000 2.805000 ;
      RECT 1284.005000 -0.085000 1284.175000 0.085000 ;
      RECT 1284.005000  2.635000 1284.175000 2.805000 ;
      RECT 1284.465000 -0.085000 1284.635000 0.085000 ;
      RECT 1284.465000  2.635000 1284.635000 2.805000 ;
      RECT 1284.925000 -0.085000 1285.095000 0.085000 ;
      RECT 1284.925000  2.635000 1285.095000 2.805000 ;
      RECT 1285.385000 -0.085000 1285.555000 0.085000 ;
      RECT 1285.385000  2.635000 1285.555000 2.805000 ;
      RECT 1285.845000 -0.085000 1286.015000 0.085000 ;
      RECT 1285.845000  2.635000 1286.015000 2.805000 ;
      RECT 1286.305000 -0.085000 1286.475000 0.085000 ;
      RECT 1286.305000  2.635000 1286.475000 2.805000 ;
      RECT 1286.765000 -0.085000 1286.935000 0.085000 ;
      RECT 1286.765000  2.635000 1286.935000 2.805000 ;
      RECT 1287.225000 -0.085000 1287.395000 0.085000 ;
      RECT 1287.225000  2.635000 1287.395000 2.805000 ;
      RECT 1287.685000 -0.085000 1287.855000 0.085000 ;
      RECT 1287.685000  2.635000 1287.855000 2.805000 ;
      RECT 1288.145000 -0.085000 1288.315000 0.085000 ;
      RECT 1288.145000  2.635000 1288.315000 2.805000 ;
      RECT 1288.605000 -0.085000 1288.775000 0.085000 ;
      RECT 1288.605000  2.635000 1288.775000 2.805000 ;
      RECT 1289.065000 -0.085000 1289.235000 0.085000 ;
      RECT 1289.065000  2.635000 1289.235000 2.805000 ;
      RECT 1289.525000 -0.085000 1289.695000 0.085000 ;
      RECT 1289.525000  2.635000 1289.695000 2.805000 ;
      RECT 1289.985000 -0.085000 1290.155000 0.085000 ;
      RECT 1289.985000  2.635000 1290.155000 2.805000 ;
      RECT 1290.445000 -0.085000 1290.615000 0.085000 ;
      RECT 1290.445000  2.635000 1290.615000 2.805000 ;
      RECT 1290.905000 -0.085000 1291.075000 0.085000 ;
      RECT 1290.905000  2.635000 1291.075000 2.805000 ;
      RECT 1291.365000 -0.085000 1291.535000 0.085000 ;
      RECT 1291.365000  2.635000 1291.535000 2.805000 ;
      RECT 1291.825000 -0.085000 1291.995000 0.085000 ;
      RECT 1291.825000  2.635000 1291.995000 2.805000 ;
      RECT 1292.285000 -0.085000 1292.455000 0.085000 ;
      RECT 1292.285000  2.635000 1292.455000 2.805000 ;
      RECT 1292.745000 -0.085000 1292.915000 0.085000 ;
      RECT 1292.745000  2.635000 1292.915000 2.805000 ;
      RECT 1293.205000 -0.085000 1293.375000 0.085000 ;
      RECT 1293.205000  2.635000 1293.375000 2.805000 ;
      RECT 1293.665000 -0.085000 1293.835000 0.085000 ;
      RECT 1293.665000  2.635000 1293.835000 2.805000 ;
      RECT 1294.125000 -0.085000 1294.295000 0.085000 ;
      RECT 1294.125000  2.635000 1294.295000 2.805000 ;
      RECT 1294.585000 -0.085000 1294.755000 0.085000 ;
      RECT 1294.585000  2.635000 1294.755000 2.805000 ;
      RECT 1295.045000 -0.085000 1295.215000 0.085000 ;
      RECT 1295.045000  2.635000 1295.215000 2.805000 ;
      RECT 1295.505000 -0.085000 1295.675000 0.085000 ;
      RECT 1295.505000  2.635000 1295.675000 2.805000 ;
      RECT 1295.965000 -0.085000 1296.135000 0.085000 ;
      RECT 1295.965000  2.635000 1296.135000 2.805000 ;
      RECT 1296.425000 -0.085000 1296.595000 0.085000 ;
      RECT 1296.425000  2.635000 1296.595000 2.805000 ;
      RECT 1296.885000 -0.085000 1297.055000 0.085000 ;
      RECT 1296.885000  2.635000 1297.055000 2.805000 ;
      RECT 1297.345000 -0.085000 1297.515000 0.085000 ;
      RECT 1297.345000  2.635000 1297.515000 2.805000 ;
      RECT 1297.805000 -0.085000 1297.975000 0.085000 ;
      RECT 1297.805000  2.635000 1297.975000 2.805000 ;
      RECT 1298.265000 -0.085000 1298.435000 0.085000 ;
      RECT 1298.265000  2.635000 1298.435000 2.805000 ;
      RECT 1298.725000 -0.085000 1298.895000 0.085000 ;
      RECT 1298.725000  2.635000 1298.895000 2.805000 ;
      RECT 1299.185000 -0.085000 1299.355000 0.085000 ;
      RECT 1299.185000  2.635000 1299.355000 2.805000 ;
      RECT 1299.645000 -0.085000 1299.815000 0.085000 ;
      RECT 1299.645000  2.635000 1299.815000 2.805000 ;
      RECT 1300.105000 -0.085000 1300.275000 0.085000 ;
      RECT 1300.105000  2.635000 1300.275000 2.805000 ;
      RECT 1300.565000 -0.085000 1300.735000 0.085000 ;
      RECT 1300.565000  2.635000 1300.735000 2.805000 ;
      RECT 1301.025000 -0.085000 1301.195000 0.085000 ;
      RECT 1301.025000  2.635000 1301.195000 2.805000 ;
      RECT 1301.485000 -0.085000 1301.655000 0.085000 ;
      RECT 1301.485000  2.635000 1301.655000 2.805000 ;
      RECT 1301.945000 -0.085000 1302.115000 0.085000 ;
      RECT 1301.945000  2.635000 1302.115000 2.805000 ;
      RECT 1302.405000 -0.085000 1302.575000 0.085000 ;
      RECT 1302.405000  2.635000 1302.575000 2.805000 ;
      RECT 1302.865000 -0.085000 1303.035000 0.085000 ;
      RECT 1302.865000  2.635000 1303.035000 2.805000 ;
      RECT 1303.325000 -0.085000 1303.495000 0.085000 ;
      RECT 1303.325000  2.635000 1303.495000 2.805000 ;
      RECT 1303.785000 -0.085000 1303.955000 0.085000 ;
      RECT 1303.785000  2.635000 1303.955000 2.805000 ;
      RECT 1304.245000 -0.085000 1304.415000 0.085000 ;
      RECT 1304.245000  2.635000 1304.415000 2.805000 ;
      RECT 1304.705000 -0.085000 1304.875000 0.085000 ;
      RECT 1304.705000  2.635000 1304.875000 2.805000 ;
      RECT 1305.165000 -0.085000 1305.335000 0.085000 ;
      RECT 1305.165000  2.635000 1305.335000 2.805000 ;
      RECT 1305.625000 -0.085000 1305.795000 0.085000 ;
      RECT 1305.625000  2.635000 1305.795000 2.805000 ;
      RECT 1306.085000 -0.085000 1306.255000 0.085000 ;
      RECT 1306.085000  2.635000 1306.255000 2.805000 ;
      RECT 1306.545000 -0.085000 1306.715000 0.085000 ;
      RECT 1306.545000  2.635000 1306.715000 2.805000 ;
      RECT 1307.005000 -0.085000 1307.175000 0.085000 ;
      RECT 1307.005000  2.635000 1307.175000 2.805000 ;
      RECT 1307.465000 -0.085000 1307.635000 0.085000 ;
      RECT 1307.465000  2.635000 1307.635000 2.805000 ;
      RECT 1307.925000 -0.085000 1308.095000 0.085000 ;
      RECT 1307.925000  2.635000 1308.095000 2.805000 ;
      RECT 1308.385000 -0.085000 1308.555000 0.085000 ;
      RECT 1308.385000  2.635000 1308.555000 2.805000 ;
      RECT 1308.845000 -0.085000 1309.015000 0.085000 ;
      RECT 1308.845000  2.635000 1309.015000 2.805000 ;
      RECT 1309.305000 -0.085000 1309.475000 0.085000 ;
      RECT 1309.305000  2.635000 1309.475000 2.805000 ;
      RECT 1309.765000 -0.085000 1309.935000 0.085000 ;
      RECT 1309.765000  2.635000 1309.935000 2.805000 ;
      RECT 1310.225000 -0.085000 1310.395000 0.085000 ;
      RECT 1310.225000  2.635000 1310.395000 2.805000 ;
      RECT 1310.685000 -0.085000 1310.855000 0.085000 ;
      RECT 1310.685000  2.635000 1310.855000 2.805000 ;
      RECT 1311.145000 -0.085000 1311.315000 0.085000 ;
      RECT 1311.145000  2.635000 1311.315000 2.805000 ;
      RECT 1311.605000 -0.085000 1311.775000 0.085000 ;
      RECT 1311.605000  2.635000 1311.775000 2.805000 ;
      RECT 1312.065000 -0.085000 1312.235000 0.085000 ;
      RECT 1312.065000  2.635000 1312.235000 2.805000 ;
      RECT 1312.525000 -0.085000 1312.695000 0.085000 ;
      RECT 1312.525000  2.635000 1312.695000 2.805000 ;
      RECT 1312.985000 -0.085000 1313.155000 0.085000 ;
      RECT 1312.985000  2.635000 1313.155000 2.805000 ;
      RECT 1313.445000 -0.085000 1313.615000 0.085000 ;
      RECT 1313.445000  2.635000 1313.615000 2.805000 ;
      RECT 1313.905000 -0.085000 1314.075000 0.085000 ;
      RECT 1313.905000  2.635000 1314.075000 2.805000 ;
      RECT 1314.365000 -0.085000 1314.535000 0.085000 ;
      RECT 1314.365000  2.635000 1314.535000 2.805000 ;
      RECT 1314.825000 -0.085000 1314.995000 0.085000 ;
      RECT 1314.825000  2.635000 1314.995000 2.805000 ;
      RECT 1315.285000 -0.085000 1315.455000 0.085000 ;
      RECT 1315.285000  2.635000 1315.455000 2.805000 ;
      RECT 1315.745000 -0.085000 1315.915000 0.085000 ;
      RECT 1315.745000  2.635000 1315.915000 2.805000 ;
      RECT 1316.205000 -0.085000 1316.375000 0.085000 ;
      RECT 1316.205000  2.635000 1316.375000 2.805000 ;
      RECT 1316.665000 -0.085000 1316.835000 0.085000 ;
      RECT 1316.665000  2.635000 1316.835000 2.805000 ;
      RECT 1317.125000 -0.085000 1317.295000 0.085000 ;
      RECT 1317.125000  2.635000 1317.295000 2.805000 ;
      RECT 1317.585000 -0.085000 1317.755000 0.085000 ;
      RECT 1317.585000  2.635000 1317.755000 2.805000 ;
      RECT 1318.045000 -0.085000 1318.215000 0.085000 ;
      RECT 1318.045000  2.635000 1318.215000 2.805000 ;
      RECT 1318.505000 -0.085000 1318.675000 0.085000 ;
      RECT 1318.505000  2.635000 1318.675000 2.805000 ;
      RECT 1318.965000 -0.085000 1319.135000 0.085000 ;
      RECT 1318.965000  2.635000 1319.135000 2.805000 ;
      RECT 1319.425000 -0.085000 1319.595000 0.085000 ;
      RECT 1319.425000  2.635000 1319.595000 2.805000 ;
      RECT 1319.885000 -0.085000 1320.055000 0.085000 ;
      RECT 1319.885000  2.635000 1320.055000 2.805000 ;
      RECT 1320.345000 -0.085000 1320.515000 0.085000 ;
      RECT 1320.345000  2.635000 1320.515000 2.805000 ;
      RECT 1320.805000 -0.085000 1320.975000 0.085000 ;
      RECT 1320.805000  2.635000 1320.975000 2.805000 ;
      RECT 1321.265000 -0.085000 1321.435000 0.085000 ;
      RECT 1321.265000  2.635000 1321.435000 2.805000 ;
      RECT 1321.725000 -0.085000 1321.895000 0.085000 ;
      RECT 1321.725000  2.635000 1321.895000 2.805000 ;
      RECT 1322.185000 -0.085000 1322.355000 0.085000 ;
      RECT 1322.185000  2.635000 1322.355000 2.805000 ;
      RECT 1322.645000 -0.085000 1322.815000 0.085000 ;
      RECT 1322.645000  2.635000 1322.815000 2.805000 ;
      RECT 1323.105000 -0.085000 1323.275000 0.085000 ;
      RECT 1323.105000  2.635000 1323.275000 2.805000 ;
      RECT 1323.565000 -0.085000 1323.735000 0.085000 ;
      RECT 1323.565000  2.635000 1323.735000 2.805000 ;
      RECT 1324.025000 -0.085000 1324.195000 0.085000 ;
      RECT 1324.025000  2.635000 1324.195000 2.805000 ;
      RECT 1324.485000 -0.085000 1324.655000 0.085000 ;
      RECT 1324.485000  2.635000 1324.655000 2.805000 ;
      RECT 1324.945000 -0.085000 1325.115000 0.085000 ;
      RECT 1324.945000  2.635000 1325.115000 2.805000 ;
      RECT 1325.405000 -0.085000 1325.575000 0.085000 ;
      RECT 1325.405000  2.635000 1325.575000 2.805000 ;
      RECT 1325.865000 -0.085000 1326.035000 0.085000 ;
      RECT 1325.865000  2.635000 1326.035000 2.805000 ;
      RECT 1326.325000 -0.085000 1326.495000 0.085000 ;
      RECT 1326.325000  2.635000 1326.495000 2.805000 ;
      RECT 1326.785000 -0.085000 1326.955000 0.085000 ;
      RECT 1326.785000  2.635000 1326.955000 2.805000 ;
      RECT 1327.245000 -0.085000 1327.415000 0.085000 ;
      RECT 1327.245000  2.635000 1327.415000 2.805000 ;
      RECT 1327.705000 -0.085000 1327.875000 0.085000 ;
      RECT 1327.705000  2.635000 1327.875000 2.805000 ;
      RECT 1328.165000 -0.085000 1328.335000 0.085000 ;
      RECT 1328.165000  2.635000 1328.335000 2.805000 ;
      RECT 1328.625000 -0.085000 1328.795000 0.085000 ;
      RECT 1328.625000  2.635000 1328.795000 2.805000 ;
      RECT 1329.085000 -0.085000 1329.255000 0.085000 ;
      RECT 1329.085000  2.635000 1329.255000 2.805000 ;
      RECT 1329.545000 -0.085000 1329.715000 0.085000 ;
      RECT 1329.545000  2.635000 1329.715000 2.805000 ;
      RECT 1330.005000 -0.085000 1330.175000 0.085000 ;
      RECT 1330.005000  2.635000 1330.175000 2.805000 ;
      RECT 1330.465000 -0.085000 1330.635000 0.085000 ;
      RECT 1330.465000  2.635000 1330.635000 2.805000 ;
      RECT 1330.925000 -0.085000 1331.095000 0.085000 ;
      RECT 1330.925000  2.635000 1331.095000 2.805000 ;
      RECT 1331.385000 -0.085000 1331.555000 0.085000 ;
      RECT 1331.385000  2.635000 1331.555000 2.805000 ;
      RECT 1331.845000 -0.085000 1332.015000 0.085000 ;
      RECT 1331.845000  2.635000 1332.015000 2.805000 ;
      RECT 1332.305000 -0.085000 1332.475000 0.085000 ;
      RECT 1332.305000  2.635000 1332.475000 2.805000 ;
      RECT 1332.765000 -0.085000 1332.935000 0.085000 ;
      RECT 1332.765000  2.635000 1332.935000 2.805000 ;
      RECT 1333.225000 -0.085000 1333.395000 0.085000 ;
      RECT 1333.225000  2.635000 1333.395000 2.805000 ;
      RECT 1333.685000 -0.085000 1333.855000 0.085000 ;
      RECT 1333.685000  2.635000 1333.855000 2.805000 ;
      RECT 1334.145000 -0.085000 1334.315000 0.085000 ;
      RECT 1334.145000  2.635000 1334.315000 2.805000 ;
      RECT 1334.605000 -0.085000 1334.775000 0.085000 ;
      RECT 1334.605000  2.635000 1334.775000 2.805000 ;
      RECT 1335.065000 -0.085000 1335.235000 0.085000 ;
      RECT 1335.065000  2.635000 1335.235000 2.805000 ;
      RECT 1335.525000 -0.085000 1335.695000 0.085000 ;
      RECT 1335.525000  2.635000 1335.695000 2.805000 ;
      RECT 1335.985000 -0.085000 1336.155000 0.085000 ;
      RECT 1335.985000  2.635000 1336.155000 2.805000 ;
      RECT 1336.445000 -0.085000 1336.615000 0.085000 ;
      RECT 1336.445000  2.635000 1336.615000 2.805000 ;
      RECT 1336.905000 -0.085000 1337.075000 0.085000 ;
      RECT 1336.905000  2.635000 1337.075000 2.805000 ;
      RECT 1337.365000 -0.085000 1337.535000 0.085000 ;
      RECT 1337.365000  2.635000 1337.535000 2.805000 ;
      RECT 1337.825000 -0.085000 1337.995000 0.085000 ;
      RECT 1337.825000  2.635000 1337.995000 2.805000 ;
      RECT 1338.285000 -0.085000 1338.455000 0.085000 ;
      RECT 1338.285000  2.635000 1338.455000 2.805000 ;
      RECT 1338.745000 -0.085000 1338.915000 0.085000 ;
      RECT 1338.745000  2.635000 1338.915000 2.805000 ;
      RECT 1339.205000 -0.085000 1339.375000 0.085000 ;
      RECT 1339.205000  2.635000 1339.375000 2.805000 ;
      RECT 1339.665000 -0.085000 1339.835000 0.085000 ;
      RECT 1339.665000  2.635000 1339.835000 2.805000 ;
      RECT 1340.125000 -0.085000 1340.295000 0.085000 ;
      RECT 1340.125000  2.635000 1340.295000 2.805000 ;
      RECT 1340.585000 -0.085000 1340.755000 0.085000 ;
      RECT 1340.585000  2.635000 1340.755000 2.805000 ;
      RECT 1341.045000 -0.085000 1341.215000 0.085000 ;
      RECT 1341.045000  2.635000 1341.215000 2.805000 ;
      RECT 1341.505000 -0.085000 1341.675000 0.085000 ;
      RECT 1341.505000  2.635000 1341.675000 2.805000 ;
      RECT 1341.965000 -0.085000 1342.135000 0.085000 ;
      RECT 1341.965000  2.635000 1342.135000 2.805000 ;
      RECT 1342.425000 -0.085000 1342.595000 0.085000 ;
      RECT 1342.425000  2.635000 1342.595000 2.805000 ;
      RECT 1342.885000 -0.085000 1343.055000 0.085000 ;
      RECT 1342.885000  2.635000 1343.055000 2.805000 ;
      RECT 1343.345000 -0.085000 1343.515000 0.085000 ;
      RECT 1343.345000  2.635000 1343.515000 2.805000 ;
      RECT 1343.805000 -0.085000 1343.975000 0.085000 ;
      RECT 1343.805000  2.635000 1343.975000 2.805000 ;
      RECT 1344.265000 -0.085000 1344.435000 0.085000 ;
      RECT 1344.265000  2.635000 1344.435000 2.805000 ;
      RECT 1344.725000 -0.085000 1344.895000 0.085000 ;
      RECT 1344.725000  2.635000 1344.895000 2.805000 ;
      RECT 1345.185000 -0.085000 1345.355000 0.085000 ;
      RECT 1345.185000  2.635000 1345.355000 2.805000 ;
      RECT 1345.645000 -0.085000 1345.815000 0.085000 ;
      RECT 1345.645000  2.635000 1345.815000 2.805000 ;
      RECT 1346.105000 -0.085000 1346.275000 0.085000 ;
      RECT 1346.105000  2.635000 1346.275000 2.805000 ;
      RECT 1346.565000 -0.085000 1346.735000 0.085000 ;
      RECT 1346.565000  2.635000 1346.735000 2.805000 ;
      RECT 1347.025000 -0.085000 1347.195000 0.085000 ;
      RECT 1347.025000  2.635000 1347.195000 2.805000 ;
      RECT 1347.485000 -0.085000 1347.655000 0.085000 ;
      RECT 1347.485000  2.635000 1347.655000 2.805000 ;
      RECT 1347.945000 -0.085000 1348.115000 0.085000 ;
      RECT 1347.945000  2.635000 1348.115000 2.805000 ;
      RECT 1348.405000 -0.085000 1348.575000 0.085000 ;
      RECT 1348.405000  2.635000 1348.575000 2.805000 ;
      RECT 1348.865000 -0.085000 1349.035000 0.085000 ;
      RECT 1348.865000  2.635000 1349.035000 2.805000 ;
      RECT 1349.325000 -0.085000 1349.495000 0.085000 ;
      RECT 1349.325000  2.635000 1349.495000 2.805000 ;
      RECT 1349.785000 -0.085000 1349.955000 0.085000 ;
      RECT 1349.785000  2.635000 1349.955000 2.805000 ;
      RECT 1350.245000 -0.085000 1350.415000 0.085000 ;
      RECT 1350.245000  2.635000 1350.415000 2.805000 ;
      RECT 1350.295000  1.785000 1350.465000 1.955000 ;
      RECT 1350.705000 -0.085000 1350.875000 0.085000 ;
      RECT 1350.705000  2.635000 1350.875000 2.805000 ;
      RECT 1350.790000  0.765000 1350.960000 0.935000 ;
      RECT 1351.165000 -0.085000 1351.335000 0.085000 ;
      RECT 1351.165000  2.635000 1351.335000 2.805000 ;
      RECT 1351.625000 -0.085000 1351.795000 0.085000 ;
      RECT 1351.625000  2.635000 1351.795000 2.805000 ;
      RECT 1352.085000 -0.085000 1352.255000 0.085000 ;
      RECT 1352.085000  2.635000 1352.255000 2.805000 ;
      RECT 1352.545000 -0.085000 1352.715000 0.085000 ;
      RECT 1352.545000  2.635000 1352.715000 2.805000 ;
      RECT 1352.745000  1.105000 1352.915000 1.275000 ;
      RECT 1353.005000 -0.085000 1353.175000 0.085000 ;
      RECT 1353.005000  2.635000 1353.175000 2.805000 ;
      RECT 1353.465000 -0.085000 1353.635000 0.085000 ;
      RECT 1353.465000  2.635000 1353.635000 2.805000 ;
      RECT 1353.925000 -0.085000 1354.095000 0.085000 ;
      RECT 1353.925000  2.635000 1354.095000 2.805000 ;
      RECT 1354.285000  1.105000 1354.455000 1.275000 ;
      RECT 1354.385000 -0.085000 1354.555000 0.085000 ;
      RECT 1354.385000  2.635000 1354.555000 2.805000 ;
      RECT 1354.785000  1.785000 1354.955000 1.955000 ;
      RECT 1354.845000 -0.085000 1355.015000 0.085000 ;
      RECT 1354.845000  2.635000 1355.015000 2.805000 ;
      RECT 1355.295000  0.765000 1355.465000 0.935000 ;
      RECT 1355.305000 -0.085000 1355.475000 0.085000 ;
      RECT 1355.305000  2.635000 1355.475000 2.805000 ;
      RECT 1355.765000 -0.085000 1355.935000 0.085000 ;
      RECT 1355.765000  2.635000 1355.935000 2.805000 ;
      RECT 1356.225000 -0.085000 1356.395000 0.085000 ;
      RECT 1356.225000  0.765000 1356.395000 0.935000 ;
      RECT 1356.225000  2.635000 1356.395000 2.805000 ;
      RECT 1356.685000 -0.085000 1356.855000 0.085000 ;
      RECT 1356.685000  2.635000 1356.855000 2.805000 ;
      RECT 1357.145000 -0.085000 1357.315000 0.085000 ;
      RECT 1357.145000  2.635000 1357.315000 2.805000 ;
      RECT 1357.605000 -0.085000 1357.775000 0.085000 ;
      RECT 1357.605000  2.635000 1357.775000 2.805000 ;
      RECT 1358.065000 -0.085000 1358.235000 0.085000 ;
      RECT 1358.065000  2.635000 1358.235000 2.805000 ;
      RECT 1358.355000  1.445000 1358.525000 1.615000 ;
      RECT 1358.525000 -0.085000 1358.695000 0.085000 ;
      RECT 1358.525000  2.635000 1358.695000 2.805000 ;
      RECT 1358.815000  1.105000 1358.985000 1.275000 ;
      RECT 1358.815000  1.785000 1358.985000 1.955000 ;
      RECT 1358.985000 -0.085000 1359.155000 0.085000 ;
      RECT 1358.985000  2.635000 1359.155000 2.805000 ;
      RECT 1359.445000 -0.085000 1359.615000 0.085000 ;
      RECT 1359.445000  2.635000 1359.615000 2.805000 ;
      RECT 1359.905000 -0.085000 1360.075000 0.085000 ;
      RECT 1359.905000  2.635000 1360.075000 2.805000 ;
      RECT 1360.355000  0.765000 1360.525000 0.935000 ;
      RECT 1360.365000 -0.085000 1360.535000 0.085000 ;
      RECT 1360.365000  2.635000 1360.535000 2.805000 ;
      RECT 1360.825000 -0.085000 1360.995000 0.085000 ;
      RECT 1360.825000  2.635000 1360.995000 2.805000 ;
      RECT 1361.285000 -0.085000 1361.455000 0.085000 ;
      RECT 1361.285000  2.635000 1361.455000 2.805000 ;
      RECT 1361.745000 -0.085000 1361.915000 0.085000 ;
      RECT 1361.745000  2.635000 1361.915000 2.805000 ;
      RECT 1361.805000  1.445000 1361.975000 1.615000 ;
      RECT 1362.205000 -0.085000 1362.375000 0.085000 ;
      RECT 1362.205000  2.635000 1362.375000 2.805000 ;
      RECT 1362.665000 -0.085000 1362.835000 0.085000 ;
      RECT 1362.665000  2.635000 1362.835000 2.805000 ;
      RECT 1363.125000 -0.085000 1363.295000 0.085000 ;
      RECT 1363.125000  2.635000 1363.295000 2.805000 ;
      RECT 1363.585000 -0.085000 1363.755000 0.085000 ;
      RECT 1363.585000  2.635000 1363.755000 2.805000 ;
      RECT 1364.045000 -0.085000 1364.215000 0.085000 ;
      RECT 1364.045000  2.635000 1364.215000 2.805000 ;
      RECT 1364.505000 -0.085000 1364.675000 0.085000 ;
      RECT 1364.505000  2.635000 1364.675000 2.805000 ;
      RECT 1364.965000 -0.085000 1365.135000 0.085000 ;
      RECT 1364.965000  2.635000 1365.135000 2.805000 ;
      RECT 1365.425000 -0.085000 1365.595000 0.085000 ;
      RECT 1365.425000  2.635000 1365.595000 2.805000 ;
      RECT 1365.885000 -0.085000 1366.055000 0.085000 ;
      RECT 1365.885000  2.635000 1366.055000 2.805000 ;
      RECT 1366.345000 -0.085000 1366.515000 0.085000 ;
      RECT 1366.345000  2.635000 1366.515000 2.805000 ;
      RECT 1366.595000  1.105000 1366.765000 1.275000 ;
      RECT 1366.805000 -0.085000 1366.975000 0.085000 ;
      RECT 1366.805000  2.635000 1366.975000 2.805000 ;
      RECT 1366.875000  1.785000 1367.045000 1.955000 ;
      RECT 1367.265000 -0.085000 1367.435000 0.085000 ;
      RECT 1367.265000  2.635000 1367.435000 2.805000 ;
      RECT 1367.725000 -0.085000 1367.895000 0.085000 ;
      RECT 1367.725000  2.635000 1367.895000 2.805000 ;
      RECT 1368.185000 -0.085000 1368.355000 0.085000 ;
      RECT 1368.185000  2.635000 1368.355000 2.805000 ;
      RECT 1368.645000 -0.085000 1368.815000 0.085000 ;
      RECT 1368.645000  2.635000 1368.815000 2.805000 ;
      RECT 1369.105000 -0.085000 1369.275000 0.085000 ;
      RECT 1369.105000  2.635000 1369.275000 2.805000 ;
      RECT 1369.565000 -0.085000 1369.735000 0.085000 ;
      RECT 1369.565000  2.635000 1369.735000 2.805000 ;
      RECT 1370.025000 -0.085000 1370.195000 0.085000 ;
      RECT 1370.025000  2.635000 1370.195000 2.805000 ;
      RECT 1370.485000 -0.085000 1370.655000 0.085000 ;
      RECT 1370.485000  2.635000 1370.655000 2.805000 ;
      RECT 1370.945000 -0.085000 1371.115000 0.085000 ;
      RECT 1370.945000  2.635000 1371.115000 2.805000 ;
      RECT 1371.220000  1.105000 1371.390000 1.275000 ;
      RECT 1371.405000 -0.085000 1371.575000 0.085000 ;
      RECT 1371.405000  2.635000 1371.575000 2.805000 ;
      RECT 1371.690000  1.785000 1371.860000 1.955000 ;
      RECT 1371.865000 -0.085000 1372.035000 0.085000 ;
      RECT 1371.865000  2.635000 1372.035000 2.805000 ;
      RECT 1372.325000 -0.085000 1372.495000 0.085000 ;
      RECT 1372.325000  2.635000 1372.495000 2.805000 ;
      RECT 1372.785000 -0.085000 1372.955000 0.085000 ;
      RECT 1372.785000  2.635000 1372.955000 2.805000 ;
      RECT 1372.995000  0.765000 1373.165000 0.935000 ;
      RECT 1373.245000 -0.085000 1373.415000 0.085000 ;
      RECT 1373.245000  2.635000 1373.415000 2.805000 ;
      RECT 1373.355000  0.765000 1373.525000 0.935000 ;
      RECT 1373.705000 -0.085000 1373.875000 0.085000 ;
      RECT 1373.705000  2.635000 1373.875000 2.805000 ;
      RECT 1374.165000 -0.085000 1374.335000 0.085000 ;
      RECT 1374.165000  2.635000 1374.335000 2.805000 ;
      RECT 1374.625000 -0.085000 1374.795000 0.085000 ;
      RECT 1374.625000  2.635000 1374.795000 2.805000 ;
      RECT 1374.975000  1.105000 1375.145000 1.275000 ;
      RECT 1375.085000 -0.085000 1375.255000 0.085000 ;
      RECT 1375.085000  2.635000 1375.255000 2.805000 ;
      RECT 1375.305000  1.785000 1375.475000 1.955000 ;
      RECT 1375.545000 -0.085000 1375.715000 0.085000 ;
      RECT 1375.545000  2.635000 1375.715000 2.805000 ;
      RECT 1376.005000 -0.085000 1376.175000 0.085000 ;
      RECT 1376.005000  2.635000 1376.175000 2.805000 ;
      RECT 1376.465000 -0.085000 1376.635000 0.085000 ;
      RECT 1376.465000  2.635000 1376.635000 2.805000 ;
      RECT 1376.915000  0.765000 1377.085000 0.935000 ;
      RECT 1376.925000 -0.085000 1377.095000 0.085000 ;
      RECT 1376.925000  2.635000 1377.095000 2.805000 ;
      RECT 1377.385000 -0.085000 1377.555000 0.085000 ;
      RECT 1377.385000  2.635000 1377.555000 2.805000 ;
      RECT 1377.845000 -0.085000 1378.015000 0.085000 ;
      RECT 1377.845000  2.635000 1378.015000 2.805000 ;
      RECT 1378.305000 -0.085000 1378.475000 0.085000 ;
      RECT 1378.305000  2.635000 1378.475000 2.805000 ;
      RECT 1378.765000 -0.085000 1378.935000 0.085000 ;
      RECT 1378.765000  2.635000 1378.935000 2.805000 ;
      RECT 1379.225000 -0.085000 1379.395000 0.085000 ;
      RECT 1379.225000  2.635000 1379.395000 2.805000 ;
      RECT 1379.685000 -0.085000 1379.855000 0.085000 ;
      RECT 1379.685000  2.635000 1379.855000 2.805000 ;
      RECT 1380.145000 -0.085000 1380.315000 0.085000 ;
      RECT 1380.145000  2.635000 1380.315000 2.805000 ;
      RECT 1380.605000 -0.085000 1380.775000 0.085000 ;
      RECT 1380.605000  2.635000 1380.775000 2.805000 ;
      RECT 1381.065000 -0.085000 1381.235000 0.085000 ;
      RECT 1381.065000  2.635000 1381.235000 2.805000 ;
      RECT 1381.315000  1.105000 1381.485000 1.275000 ;
      RECT 1381.525000 -0.085000 1381.695000 0.085000 ;
      RECT 1381.525000  2.635000 1381.695000 2.805000 ;
      RECT 1381.595000  1.785000 1381.765000 1.955000 ;
      RECT 1381.985000 -0.085000 1382.155000 0.085000 ;
      RECT 1381.985000  2.635000 1382.155000 2.805000 ;
      RECT 1382.445000 -0.085000 1382.615000 0.085000 ;
      RECT 1382.445000  2.635000 1382.615000 2.805000 ;
      RECT 1382.905000 -0.085000 1383.075000 0.085000 ;
      RECT 1382.905000  2.635000 1383.075000 2.805000 ;
      RECT 1383.365000 -0.085000 1383.535000 0.085000 ;
      RECT 1383.365000  2.635000 1383.535000 2.805000 ;
      RECT 1383.825000 -0.085000 1383.995000 0.085000 ;
      RECT 1383.825000  2.635000 1383.995000 2.805000 ;
      RECT 1384.285000 -0.085000 1384.455000 0.085000 ;
      RECT 1384.285000  2.635000 1384.455000 2.805000 ;
      RECT 1384.745000 -0.085000 1384.915000 0.085000 ;
      RECT 1384.745000  2.635000 1384.915000 2.805000 ;
      RECT 1385.205000 -0.085000 1385.375000 0.085000 ;
      RECT 1385.205000  2.635000 1385.375000 2.805000 ;
      RECT 1385.665000 -0.085000 1385.835000 0.085000 ;
      RECT 1385.665000  2.635000 1385.835000 2.805000 ;
      RECT 1385.940000  1.105000 1386.110000 1.275000 ;
      RECT 1386.125000 -0.085000 1386.295000 0.085000 ;
      RECT 1386.125000  2.635000 1386.295000 2.805000 ;
      RECT 1386.410000  1.785000 1386.580000 1.955000 ;
      RECT 1386.585000 -0.085000 1386.755000 0.085000 ;
      RECT 1386.585000  2.635000 1386.755000 2.805000 ;
      RECT 1387.045000 -0.085000 1387.215000 0.085000 ;
      RECT 1387.045000  2.635000 1387.215000 2.805000 ;
      RECT 1387.505000 -0.085000 1387.675000 0.085000 ;
      RECT 1387.505000  2.635000 1387.675000 2.805000 ;
      RECT 1387.715000  0.765000 1387.885000 0.935000 ;
      RECT 1387.965000 -0.085000 1388.135000 0.085000 ;
      RECT 1387.965000  2.635000 1388.135000 2.805000 ;
      RECT 1388.075000  0.765000 1388.245000 0.935000 ;
      RECT 1388.425000 -0.085000 1388.595000 0.085000 ;
      RECT 1388.425000  2.635000 1388.595000 2.805000 ;
      RECT 1388.885000 -0.085000 1389.055000 0.085000 ;
      RECT 1388.885000  2.635000 1389.055000 2.805000 ;
      RECT 1389.345000 -0.085000 1389.515000 0.085000 ;
      RECT 1389.345000  2.635000 1389.515000 2.805000 ;
      RECT 1389.695000  1.105000 1389.865000 1.275000 ;
      RECT 1389.805000 -0.085000 1389.975000 0.085000 ;
      RECT 1389.805000  2.635000 1389.975000 2.805000 ;
      RECT 1390.025000  1.785000 1390.195000 1.955000 ;
      RECT 1390.265000 -0.085000 1390.435000 0.085000 ;
      RECT 1390.265000  2.635000 1390.435000 2.805000 ;
      RECT 1390.725000 -0.085000 1390.895000 0.085000 ;
      RECT 1390.725000  2.635000 1390.895000 2.805000 ;
      RECT 1391.185000 -0.085000 1391.355000 0.085000 ;
      RECT 1391.185000  2.635000 1391.355000 2.805000 ;
      RECT 1391.635000  0.765000 1391.805000 0.935000 ;
      RECT 1391.645000 -0.085000 1391.815000 0.085000 ;
      RECT 1391.645000  2.635000 1391.815000 2.805000 ;
      RECT 1392.105000 -0.085000 1392.275000 0.085000 ;
      RECT 1392.105000  2.635000 1392.275000 2.805000 ;
      RECT 1392.565000 -0.085000 1392.735000 0.085000 ;
      RECT 1392.565000  2.635000 1392.735000 2.805000 ;
      RECT 1393.025000 -0.085000 1393.195000 0.085000 ;
      RECT 1393.025000  2.635000 1393.195000 2.805000 ;
      RECT 1393.485000 -0.085000 1393.655000 0.085000 ;
      RECT 1393.485000  2.635000 1393.655000 2.805000 ;
      RECT 1393.945000 -0.085000 1394.115000 0.085000 ;
      RECT 1393.945000  2.635000 1394.115000 2.805000 ;
      RECT 1394.405000 -0.085000 1394.575000 0.085000 ;
      RECT 1394.405000  2.635000 1394.575000 2.805000 ;
      RECT 1394.865000 -0.085000 1395.035000 0.085000 ;
      RECT 1394.865000  2.635000 1395.035000 2.805000 ;
      RECT 1395.325000 -0.085000 1395.495000 0.085000 ;
      RECT 1395.325000  2.635000 1395.495000 2.805000 ;
      RECT 1395.785000 -0.085000 1395.955000 0.085000 ;
      RECT 1395.785000  2.635000 1395.955000 2.805000 ;
      RECT 1396.245000 -0.085000 1396.415000 0.085000 ;
      RECT 1396.245000  2.635000 1396.415000 2.805000 ;
      RECT 1396.365000  1.785000 1396.535000 1.955000 ;
      RECT 1396.705000 -0.085000 1396.875000 0.085000 ;
      RECT 1396.705000  2.635000 1396.875000 2.805000 ;
      RECT 1396.835000  1.105000 1397.005000 1.275000 ;
      RECT 1397.165000 -0.085000 1397.335000 0.085000 ;
      RECT 1397.165000  2.635000 1397.335000 2.805000 ;
      RECT 1397.625000 -0.085000 1397.795000 0.085000 ;
      RECT 1397.625000  2.635000 1397.795000 2.805000 ;
      RECT 1398.085000 -0.085000 1398.255000 0.085000 ;
      RECT 1398.085000  2.635000 1398.255000 2.805000 ;
      RECT 1398.545000 -0.085000 1398.715000 0.085000 ;
      RECT 1398.545000  2.635000 1398.715000 2.805000 ;
      RECT 1399.005000 -0.085000 1399.175000 0.085000 ;
      RECT 1399.005000  2.635000 1399.175000 2.805000 ;
      RECT 1399.465000 -0.085000 1399.635000 0.085000 ;
      RECT 1399.465000  2.635000 1399.635000 2.805000 ;
      RECT 1399.925000 -0.085000 1400.095000 0.085000 ;
      RECT 1399.925000  2.635000 1400.095000 2.805000 ;
      RECT 1400.385000 -0.085000 1400.555000 0.085000 ;
      RECT 1400.385000  2.635000 1400.555000 2.805000 ;
      RECT 1400.845000 -0.085000 1401.015000 0.085000 ;
      RECT 1400.845000  2.635000 1401.015000 2.805000 ;
      RECT 1401.120000  1.105000 1401.290000 1.275000 ;
      RECT 1401.305000 -0.085000 1401.475000 0.085000 ;
      RECT 1401.305000  2.635000 1401.475000 2.805000 ;
      RECT 1401.590000  1.785000 1401.760000 1.955000 ;
      RECT 1401.765000 -0.085000 1401.935000 0.085000 ;
      RECT 1401.765000  2.635000 1401.935000 2.805000 ;
      RECT 1402.225000 -0.085000 1402.395000 0.085000 ;
      RECT 1402.225000  2.635000 1402.395000 2.805000 ;
      RECT 1402.685000 -0.085000 1402.855000 0.085000 ;
      RECT 1402.685000  2.635000 1402.855000 2.805000 ;
      RECT 1402.895000  0.765000 1403.065000 0.935000 ;
      RECT 1403.145000 -0.085000 1403.315000 0.085000 ;
      RECT 1403.145000  2.635000 1403.315000 2.805000 ;
      RECT 1403.255000  0.765000 1403.425000 0.935000 ;
      RECT 1403.605000 -0.085000 1403.775000 0.085000 ;
      RECT 1403.605000  2.635000 1403.775000 2.805000 ;
      RECT 1404.065000 -0.085000 1404.235000 0.085000 ;
      RECT 1404.065000  2.635000 1404.235000 2.805000 ;
      RECT 1404.525000 -0.085000 1404.695000 0.085000 ;
      RECT 1404.525000  2.635000 1404.695000 2.805000 ;
      RECT 1404.875000  1.105000 1405.045000 1.275000 ;
      RECT 1404.985000 -0.085000 1405.155000 0.085000 ;
      RECT 1404.985000  2.635000 1405.155000 2.805000 ;
      RECT 1405.205000  1.785000 1405.375000 1.955000 ;
      RECT 1405.445000 -0.085000 1405.615000 0.085000 ;
      RECT 1405.445000  2.635000 1405.615000 2.805000 ;
      RECT 1405.905000 -0.085000 1406.075000 0.085000 ;
      RECT 1405.905000  2.635000 1406.075000 2.805000 ;
      RECT 1406.365000 -0.085000 1406.535000 0.085000 ;
      RECT 1406.365000  2.635000 1406.535000 2.805000 ;
      RECT 1406.815000  0.765000 1406.985000 0.935000 ;
      RECT 1406.825000 -0.085000 1406.995000 0.085000 ;
      RECT 1406.825000  2.635000 1406.995000 2.805000 ;
      RECT 1407.285000 -0.085000 1407.455000 0.085000 ;
      RECT 1407.285000  2.635000 1407.455000 2.805000 ;
      RECT 1407.745000 -0.085000 1407.915000 0.085000 ;
      RECT 1407.745000  2.635000 1407.915000 2.805000 ;
      RECT 1408.205000 -0.085000 1408.375000 0.085000 ;
      RECT 1408.205000  2.635000 1408.375000 2.805000 ;
      RECT 1408.665000 -0.085000 1408.835000 0.085000 ;
      RECT 1408.665000  2.635000 1408.835000 2.805000 ;
      RECT 1409.125000 -0.085000 1409.295000 0.085000 ;
      RECT 1409.125000  2.635000 1409.295000 2.805000 ;
      RECT 1409.585000 -0.085000 1409.755000 0.085000 ;
      RECT 1409.585000  2.635000 1409.755000 2.805000 ;
      RECT 1409.835000  1.105000 1410.005000 1.275000 ;
      RECT 1410.045000 -0.085000 1410.215000 0.085000 ;
      RECT 1410.045000  2.635000 1410.215000 2.805000 ;
      RECT 1410.115000  1.785000 1410.285000 1.955000 ;
      RECT 1410.505000 -0.085000 1410.675000 0.085000 ;
      RECT 1410.505000  2.635000 1410.675000 2.805000 ;
      RECT 1410.965000 -0.085000 1411.135000 0.085000 ;
      RECT 1410.965000  2.635000 1411.135000 2.805000 ;
      RECT 1411.425000 -0.085000 1411.595000 0.085000 ;
      RECT 1411.425000  2.635000 1411.595000 2.805000 ;
      RECT 1411.885000 -0.085000 1412.055000 0.085000 ;
      RECT 1411.885000  2.635000 1412.055000 2.805000 ;
      RECT 1412.345000 -0.085000 1412.515000 0.085000 ;
      RECT 1412.345000  2.635000 1412.515000 2.805000 ;
      RECT 1412.805000 -0.085000 1412.975000 0.085000 ;
      RECT 1412.805000  2.635000 1412.975000 2.805000 ;
      RECT 1413.265000 -0.085000 1413.435000 0.085000 ;
      RECT 1413.265000  2.635000 1413.435000 2.805000 ;
      RECT 1413.725000 -0.085000 1413.895000 0.085000 ;
      RECT 1413.725000  2.635000 1413.895000 2.805000 ;
      RECT 1414.185000 -0.085000 1414.355000 0.085000 ;
      RECT 1414.185000  2.635000 1414.355000 2.805000 ;
      RECT 1414.460000  1.105000 1414.630000 1.275000 ;
      RECT 1414.645000 -0.085000 1414.815000 0.085000 ;
      RECT 1414.645000  2.635000 1414.815000 2.805000 ;
      RECT 1414.930000  1.785000 1415.100000 1.955000 ;
      RECT 1415.105000 -0.085000 1415.275000 0.085000 ;
      RECT 1415.105000  2.635000 1415.275000 2.805000 ;
      RECT 1415.565000 -0.085000 1415.735000 0.085000 ;
      RECT 1415.565000  2.635000 1415.735000 2.805000 ;
      RECT 1416.025000 -0.085000 1416.195000 0.085000 ;
      RECT 1416.025000  2.635000 1416.195000 2.805000 ;
      RECT 1416.235000  0.765000 1416.405000 0.935000 ;
      RECT 1416.485000 -0.085000 1416.655000 0.085000 ;
      RECT 1416.485000  2.635000 1416.655000 2.805000 ;
      RECT 1416.595000  0.765000 1416.765000 0.935000 ;
      RECT 1416.945000 -0.085000 1417.115000 0.085000 ;
      RECT 1416.945000  2.635000 1417.115000 2.805000 ;
      RECT 1417.405000 -0.085000 1417.575000 0.085000 ;
      RECT 1417.405000  2.635000 1417.575000 2.805000 ;
      RECT 1417.865000 -0.085000 1418.035000 0.085000 ;
      RECT 1417.865000  2.635000 1418.035000 2.805000 ;
      RECT 1418.215000  1.105000 1418.385000 1.275000 ;
      RECT 1418.325000 -0.085000 1418.495000 0.085000 ;
      RECT 1418.325000  2.635000 1418.495000 2.805000 ;
      RECT 1418.545000  1.785000 1418.715000 1.955000 ;
      RECT 1418.785000 -0.085000 1418.955000 0.085000 ;
      RECT 1418.785000  2.635000 1418.955000 2.805000 ;
      RECT 1419.245000 -0.085000 1419.415000 0.085000 ;
      RECT 1419.245000  2.635000 1419.415000 2.805000 ;
      RECT 1419.705000 -0.085000 1419.875000 0.085000 ;
      RECT 1419.705000  2.635000 1419.875000 2.805000 ;
      RECT 1420.155000  0.765000 1420.325000 0.935000 ;
      RECT 1420.165000 -0.085000 1420.335000 0.085000 ;
      RECT 1420.165000  2.635000 1420.335000 2.805000 ;
      RECT 1420.625000 -0.085000 1420.795000 0.085000 ;
      RECT 1420.625000  2.635000 1420.795000 2.805000 ;
      RECT 1421.085000 -0.085000 1421.255000 0.085000 ;
      RECT 1421.085000  2.635000 1421.255000 2.805000 ;
      RECT 1421.545000 -0.085000 1421.715000 0.085000 ;
      RECT 1421.545000  2.635000 1421.715000 2.805000 ;
      RECT 1422.005000 -0.085000 1422.175000 0.085000 ;
      RECT 1422.005000  2.635000 1422.175000 2.805000 ;
      RECT 1422.465000 -0.085000 1422.635000 0.085000 ;
      RECT 1422.465000  2.635000 1422.635000 2.805000 ;
      RECT 1422.925000 -0.085000 1423.095000 0.085000 ;
      RECT 1422.925000  2.635000 1423.095000 2.805000 ;
      RECT 1423.175000  1.105000 1423.345000 1.275000 ;
      RECT 1423.385000 -0.085000 1423.555000 0.085000 ;
      RECT 1423.385000  2.635000 1423.555000 2.805000 ;
      RECT 1423.455000  1.785000 1423.625000 1.955000 ;
      RECT 1423.845000 -0.085000 1424.015000 0.085000 ;
      RECT 1423.845000  2.635000 1424.015000 2.805000 ;
      RECT 1424.305000 -0.085000 1424.475000 0.085000 ;
      RECT 1424.305000  2.635000 1424.475000 2.805000 ;
      RECT 1424.765000 -0.085000 1424.935000 0.085000 ;
      RECT 1424.765000  2.635000 1424.935000 2.805000 ;
      RECT 1425.225000 -0.085000 1425.395000 0.085000 ;
      RECT 1425.225000  2.635000 1425.395000 2.805000 ;
      RECT 1425.685000 -0.085000 1425.855000 0.085000 ;
      RECT 1425.685000  2.635000 1425.855000 2.805000 ;
      RECT 1426.145000 -0.085000 1426.315000 0.085000 ;
      RECT 1426.145000  2.635000 1426.315000 2.805000 ;
      RECT 1426.605000 -0.085000 1426.775000 0.085000 ;
      RECT 1426.605000  2.635000 1426.775000 2.805000 ;
      RECT 1427.065000 -0.085000 1427.235000 0.085000 ;
      RECT 1427.065000  2.635000 1427.235000 2.805000 ;
      RECT 1427.525000 -0.085000 1427.695000 0.085000 ;
      RECT 1427.525000  2.635000 1427.695000 2.805000 ;
      RECT 1427.800000  1.105000 1427.970000 1.275000 ;
      RECT 1427.985000 -0.085000 1428.155000 0.085000 ;
      RECT 1427.985000  2.635000 1428.155000 2.805000 ;
      RECT 1428.270000  1.785000 1428.440000 1.955000 ;
      RECT 1428.445000 -0.085000 1428.615000 0.085000 ;
      RECT 1428.445000  2.635000 1428.615000 2.805000 ;
      RECT 1428.905000 -0.085000 1429.075000 0.085000 ;
      RECT 1428.905000  2.635000 1429.075000 2.805000 ;
      RECT 1429.365000 -0.085000 1429.535000 0.085000 ;
      RECT 1429.365000  2.635000 1429.535000 2.805000 ;
      RECT 1429.575000  0.765000 1429.745000 0.935000 ;
      RECT 1429.825000 -0.085000 1429.995000 0.085000 ;
      RECT 1429.825000  2.635000 1429.995000 2.805000 ;
      RECT 1429.935000  0.765000 1430.105000 0.935000 ;
      RECT 1430.285000 -0.085000 1430.455000 0.085000 ;
      RECT 1430.285000  2.635000 1430.455000 2.805000 ;
      RECT 1430.745000 -0.085000 1430.915000 0.085000 ;
      RECT 1430.745000  2.635000 1430.915000 2.805000 ;
      RECT 1431.205000 -0.085000 1431.375000 0.085000 ;
      RECT 1431.205000  2.635000 1431.375000 2.805000 ;
      RECT 1431.555000  1.105000 1431.725000 1.275000 ;
      RECT 1431.665000 -0.085000 1431.835000 0.085000 ;
      RECT 1431.665000  2.635000 1431.835000 2.805000 ;
      RECT 1431.885000  1.785000 1432.055000 1.955000 ;
      RECT 1432.125000 -0.085000 1432.295000 0.085000 ;
      RECT 1432.125000  2.635000 1432.295000 2.805000 ;
      RECT 1432.585000 -0.085000 1432.755000 0.085000 ;
      RECT 1432.585000  2.635000 1432.755000 2.805000 ;
      RECT 1433.045000 -0.085000 1433.215000 0.085000 ;
      RECT 1433.045000  2.635000 1433.215000 2.805000 ;
      RECT 1433.460000  0.765000 1433.630000 0.935000 ;
      RECT 1433.505000 -0.085000 1433.675000 0.085000 ;
      RECT 1433.505000  2.635000 1433.675000 2.805000 ;
      RECT 1433.965000 -0.085000 1434.135000 0.085000 ;
      RECT 1433.965000  2.635000 1434.135000 2.805000 ;
      RECT 1434.425000 -0.085000 1434.595000 0.085000 ;
      RECT 1434.425000  2.635000 1434.595000 2.805000 ;
      RECT 1434.885000 -0.085000 1435.055000 0.085000 ;
      RECT 1434.885000  2.635000 1435.055000 2.805000 ;
      RECT 1435.345000 -0.085000 1435.515000 0.085000 ;
      RECT 1435.345000  2.635000 1435.515000 2.805000 ;
      RECT 1435.805000 -0.085000 1435.975000 0.085000 ;
      RECT 1435.805000  2.635000 1435.975000 2.805000 ;
      RECT 1436.265000 -0.085000 1436.435000 0.085000 ;
      RECT 1436.265000  2.635000 1436.435000 2.805000 ;
      RECT 1436.725000 -0.085000 1436.895000 0.085000 ;
      RECT 1436.725000  2.635000 1436.895000 2.805000 ;
      RECT 1436.750000  1.105000 1436.920000 1.275000 ;
      RECT 1437.185000 -0.085000 1437.355000 0.085000 ;
      RECT 1437.185000  2.635000 1437.355000 2.805000 ;
      RECT 1437.645000 -0.085000 1437.815000 0.085000 ;
      RECT 1437.645000  2.635000 1437.815000 2.805000 ;
      RECT 1437.795000  1.445000 1437.965000 1.615000 ;
      RECT 1438.105000 -0.085000 1438.275000 0.085000 ;
      RECT 1438.105000  2.635000 1438.275000 2.805000 ;
      RECT 1438.565000 -0.085000 1438.735000 0.085000 ;
      RECT 1438.565000  2.635000 1438.735000 2.805000 ;
      RECT 1438.765000  1.105000 1438.935000 1.275000 ;
      RECT 1439.025000 -0.085000 1439.195000 0.085000 ;
      RECT 1439.025000  2.635000 1439.195000 2.805000 ;
      RECT 1439.485000 -0.085000 1439.655000 0.085000 ;
      RECT 1439.485000  2.635000 1439.655000 2.805000 ;
      RECT 1439.945000 -0.085000 1440.115000 0.085000 ;
      RECT 1439.945000  2.635000 1440.115000 2.805000 ;
      RECT 1440.245000  1.785000 1440.415000 1.955000 ;
      RECT 1440.405000 -0.085000 1440.575000 0.085000 ;
      RECT 1440.405000  2.635000 1440.575000 2.805000 ;
      RECT 1440.705000  1.105000 1440.875000 1.275000 ;
      RECT 1440.865000 -0.085000 1441.035000 0.085000 ;
      RECT 1440.865000  2.635000 1441.035000 2.805000 ;
      RECT 1441.130000  1.445000 1441.300000 1.615000 ;
      RECT 1441.325000 -0.085000 1441.495000 0.085000 ;
      RECT 1441.325000  2.635000 1441.495000 2.805000 ;
      RECT 1441.725000  1.785000 1441.895000 1.955000 ;
      RECT 1441.785000 -0.085000 1441.955000 0.085000 ;
      RECT 1441.785000  2.635000 1441.955000 2.805000 ;
      RECT 1442.245000 -0.085000 1442.415000 0.085000 ;
      RECT 1442.245000  2.635000 1442.415000 2.805000 ;
      RECT 1442.705000 -0.085000 1442.875000 0.085000 ;
      RECT 1442.705000  2.635000 1442.875000 2.805000 ;
      RECT 1443.165000 -0.085000 1443.335000 0.085000 ;
      RECT 1443.165000  2.635000 1443.335000 2.805000 ;
      RECT 1443.565000  1.445000 1443.735000 1.615000 ;
      RECT 1443.625000 -0.085000 1443.795000 0.085000 ;
      RECT 1443.625000  2.635000 1443.795000 2.805000 ;
      RECT 1444.085000 -0.085000 1444.255000 0.085000 ;
      RECT 1444.085000  2.635000 1444.255000 2.805000 ;
      RECT 1444.325000  1.785000 1444.495000 1.955000 ;
      RECT 1444.545000 -0.085000 1444.715000 0.085000 ;
      RECT 1444.545000  2.635000 1444.715000 2.805000 ;
      RECT 1445.005000 -0.085000 1445.175000 0.085000 ;
      RECT 1445.005000  2.635000 1445.175000 2.805000 ;
      RECT 1445.345000  1.105000 1445.515000 1.275000 ;
      RECT 1445.465000 -0.085000 1445.635000 0.085000 ;
      RECT 1445.465000  2.635000 1445.635000 2.805000 ;
      RECT 1445.855000  1.445000 1446.025000 1.615000 ;
      RECT 1445.925000 -0.085000 1446.095000 0.085000 ;
      RECT 1445.925000  2.635000 1446.095000 2.805000 ;
      RECT 1446.385000 -0.085000 1446.555000 0.085000 ;
      RECT 1446.385000  2.635000 1446.555000 2.805000 ;
      RECT 1446.845000 -0.085000 1447.015000 0.085000 ;
      RECT 1446.845000  2.635000 1447.015000 2.805000 ;
      RECT 1447.305000 -0.085000 1447.475000 0.085000 ;
      RECT 1447.305000  2.635000 1447.475000 2.805000 ;
      RECT 1447.765000 -0.085000 1447.935000 0.085000 ;
      RECT 1447.765000  2.635000 1447.935000 2.805000 ;
      RECT 1448.225000 -0.085000 1448.395000 0.085000 ;
      RECT 1448.225000  2.635000 1448.395000 2.805000 ;
      RECT 1448.685000 -0.085000 1448.855000 0.085000 ;
      RECT 1448.685000  2.635000 1448.855000 2.805000 ;
      RECT 1449.145000 -0.085000 1449.315000 0.085000 ;
      RECT 1449.145000  2.635000 1449.315000 2.805000 ;
      RECT 1449.605000 -0.085000 1449.775000 0.085000 ;
      RECT 1449.605000  2.635000 1449.775000 2.805000 ;
      RECT 1450.065000 -0.085000 1450.235000 0.085000 ;
      RECT 1450.065000  2.635000 1450.235000 2.805000 ;
      RECT 1450.525000 -0.085000 1450.695000 0.085000 ;
      RECT 1450.525000  2.635000 1450.695000 2.805000 ;
      RECT 1450.985000 -0.085000 1451.155000 0.085000 ;
      RECT 1450.985000  2.635000 1451.155000 2.805000 ;
      RECT 1451.445000 -0.085000 1451.615000 0.085000 ;
      RECT 1451.445000  2.635000 1451.615000 2.805000 ;
      RECT 1451.905000 -0.085000 1452.075000 0.085000 ;
      RECT 1451.905000  2.635000 1452.075000 2.805000 ;
      RECT 1451.930000  1.105000 1452.100000 1.275000 ;
      RECT 1452.365000 -0.085000 1452.535000 0.085000 ;
      RECT 1452.365000  2.635000 1452.535000 2.805000 ;
      RECT 1452.825000 -0.085000 1452.995000 0.085000 ;
      RECT 1452.825000  2.635000 1452.995000 2.805000 ;
      RECT 1452.975000  1.445000 1453.145000 1.615000 ;
      RECT 1453.285000 -0.085000 1453.455000 0.085000 ;
      RECT 1453.285000  2.635000 1453.455000 2.805000 ;
      RECT 1453.745000 -0.085000 1453.915000 0.085000 ;
      RECT 1453.745000  2.635000 1453.915000 2.805000 ;
      RECT 1453.945000  1.105000 1454.115000 1.275000 ;
      RECT 1454.205000 -0.085000 1454.375000 0.085000 ;
      RECT 1454.205000  2.635000 1454.375000 2.805000 ;
      RECT 1454.665000 -0.085000 1454.835000 0.085000 ;
      RECT 1454.665000  2.635000 1454.835000 2.805000 ;
      RECT 1455.125000 -0.085000 1455.295000 0.085000 ;
      RECT 1455.125000  2.635000 1455.295000 2.805000 ;
      RECT 1455.425000  1.785000 1455.595000 1.955000 ;
      RECT 1455.585000 -0.085000 1455.755000 0.085000 ;
      RECT 1455.585000  2.635000 1455.755000 2.805000 ;
      RECT 1455.885000  1.105000 1456.055000 1.275000 ;
      RECT 1456.045000 -0.085000 1456.215000 0.085000 ;
      RECT 1456.045000  2.635000 1456.215000 2.805000 ;
      RECT 1456.310000  1.445000 1456.480000 1.615000 ;
      RECT 1456.505000 -0.085000 1456.675000 0.085000 ;
      RECT 1456.505000  2.635000 1456.675000 2.805000 ;
      RECT 1456.905000  1.785000 1457.075000 1.955000 ;
      RECT 1456.965000 -0.085000 1457.135000 0.085000 ;
      RECT 1456.965000  2.635000 1457.135000 2.805000 ;
      RECT 1457.425000 -0.085000 1457.595000 0.085000 ;
      RECT 1457.425000  2.635000 1457.595000 2.805000 ;
      RECT 1457.885000 -0.085000 1458.055000 0.085000 ;
      RECT 1457.885000  2.635000 1458.055000 2.805000 ;
      RECT 1458.345000 -0.085000 1458.515000 0.085000 ;
      RECT 1458.345000  2.635000 1458.515000 2.805000 ;
      RECT 1458.745000  1.445000 1458.915000 1.615000 ;
      RECT 1458.805000 -0.085000 1458.975000 0.085000 ;
      RECT 1458.805000  2.635000 1458.975000 2.805000 ;
      RECT 1459.265000 -0.085000 1459.435000 0.085000 ;
      RECT 1459.265000  2.635000 1459.435000 2.805000 ;
      RECT 1459.505000  1.785000 1459.675000 1.955000 ;
      RECT 1459.725000 -0.085000 1459.895000 0.085000 ;
      RECT 1459.725000  2.635000 1459.895000 2.805000 ;
      RECT 1460.185000 -0.085000 1460.355000 0.085000 ;
      RECT 1460.185000  2.635000 1460.355000 2.805000 ;
      RECT 1460.525000  1.105000 1460.695000 1.275000 ;
      RECT 1460.645000 -0.085000 1460.815000 0.085000 ;
      RECT 1460.645000  2.635000 1460.815000 2.805000 ;
      RECT 1461.035000  1.445000 1461.205000 1.615000 ;
      RECT 1461.105000 -0.085000 1461.275000 0.085000 ;
      RECT 1461.105000  2.635000 1461.275000 2.805000 ;
      RECT 1461.565000 -0.085000 1461.735000 0.085000 ;
      RECT 1461.565000  2.635000 1461.735000 2.805000 ;
      RECT 1462.025000 -0.085000 1462.195000 0.085000 ;
      RECT 1462.025000  2.635000 1462.195000 2.805000 ;
      RECT 1462.485000 -0.085000 1462.655000 0.085000 ;
      RECT 1462.485000  2.635000 1462.655000 2.805000 ;
      RECT 1462.945000 -0.085000 1463.115000 0.085000 ;
      RECT 1462.945000  2.635000 1463.115000 2.805000 ;
      RECT 1463.405000 -0.085000 1463.575000 0.085000 ;
      RECT 1463.405000  2.635000 1463.575000 2.805000 ;
      RECT 1463.865000 -0.085000 1464.035000 0.085000 ;
      RECT 1463.865000  2.635000 1464.035000 2.805000 ;
      RECT 1464.325000 -0.085000 1464.495000 0.085000 ;
      RECT 1464.325000  2.635000 1464.495000 2.805000 ;
      RECT 1464.785000 -0.085000 1464.955000 0.085000 ;
      RECT 1464.785000  2.635000 1464.955000 2.805000 ;
      RECT 1465.245000 -0.085000 1465.415000 0.085000 ;
      RECT 1465.245000  2.635000 1465.415000 2.805000 ;
      RECT 1465.705000 -0.085000 1465.875000 0.085000 ;
      RECT 1465.705000  2.635000 1465.875000 2.805000 ;
      RECT 1466.165000 -0.085000 1466.335000 0.085000 ;
      RECT 1466.165000  2.635000 1466.335000 2.805000 ;
      RECT 1466.625000 -0.085000 1466.795000 0.085000 ;
      RECT 1466.625000  2.635000 1466.795000 2.805000 ;
      RECT 1467.085000 -0.085000 1467.255000 0.085000 ;
      RECT 1467.085000  2.635000 1467.255000 2.805000 ;
      RECT 1467.545000 -0.085000 1467.715000 0.085000 ;
      RECT 1467.545000  2.635000 1467.715000 2.805000 ;
      RECT 1468.005000 -0.085000 1468.175000 0.085000 ;
      RECT 1468.005000  2.635000 1468.175000 2.805000 ;
      RECT 1468.040000  1.105000 1468.210000 1.275000 ;
      RECT 1468.465000 -0.085000 1468.635000 0.085000 ;
      RECT 1468.465000  2.635000 1468.635000 2.805000 ;
      RECT 1468.925000 -0.085000 1469.095000 0.085000 ;
      RECT 1468.925000  2.635000 1469.095000 2.805000 ;
      RECT 1469.075000  1.445000 1469.245000 1.615000 ;
      RECT 1469.385000 -0.085000 1469.555000 0.085000 ;
      RECT 1469.385000  2.635000 1469.555000 2.805000 ;
      RECT 1469.845000 -0.085000 1470.015000 0.085000 ;
      RECT 1469.845000  2.635000 1470.015000 2.805000 ;
      RECT 1470.045000  1.105000 1470.215000 1.275000 ;
      RECT 1470.305000 -0.085000 1470.475000 0.085000 ;
      RECT 1470.305000  2.635000 1470.475000 2.805000 ;
      RECT 1470.765000 -0.085000 1470.935000 0.085000 ;
      RECT 1470.765000  2.635000 1470.935000 2.805000 ;
      RECT 1471.225000 -0.085000 1471.395000 0.085000 ;
      RECT 1471.225000  2.635000 1471.395000 2.805000 ;
      RECT 1471.525000  1.785000 1471.695000 1.955000 ;
      RECT 1471.685000 -0.085000 1471.855000 0.085000 ;
      RECT 1471.685000  2.635000 1471.855000 2.805000 ;
      RECT 1472.035000  1.100000 1472.205000 1.270000 ;
      RECT 1472.145000 -0.085000 1472.315000 0.085000 ;
      RECT 1472.145000  2.635000 1472.315000 2.805000 ;
      RECT 1472.410000  1.445000 1472.580000 1.615000 ;
      RECT 1472.605000 -0.085000 1472.775000 0.085000 ;
      RECT 1472.605000  2.635000 1472.775000 2.805000 ;
      RECT 1473.005000  1.785000 1473.175000 1.955000 ;
      RECT 1473.065000 -0.085000 1473.235000 0.085000 ;
      RECT 1473.065000  2.635000 1473.235000 2.805000 ;
      RECT 1473.525000 -0.085000 1473.695000 0.085000 ;
      RECT 1473.525000  2.635000 1473.695000 2.805000 ;
      RECT 1473.985000 -0.085000 1474.155000 0.085000 ;
      RECT 1473.985000  2.635000 1474.155000 2.805000 ;
      RECT 1474.445000 -0.085000 1474.615000 0.085000 ;
      RECT 1474.445000  2.635000 1474.615000 2.805000 ;
      RECT 1474.835000  1.445000 1475.005000 1.615000 ;
      RECT 1474.905000 -0.085000 1475.075000 0.085000 ;
      RECT 1474.905000  2.635000 1475.075000 2.805000 ;
      RECT 1475.365000 -0.085000 1475.535000 0.085000 ;
      RECT 1475.365000  2.635000 1475.535000 2.805000 ;
      RECT 1475.610000  1.785000 1475.780000 1.955000 ;
      RECT 1475.825000 -0.085000 1475.995000 0.085000 ;
      RECT 1475.825000  2.635000 1475.995000 2.805000 ;
      RECT 1476.285000 -0.085000 1476.455000 0.085000 ;
      RECT 1476.285000  2.635000 1476.455000 2.805000 ;
      RECT 1476.450000  1.105000 1476.620000 1.275000 ;
      RECT 1476.745000 -0.085000 1476.915000 0.085000 ;
      RECT 1476.745000  2.635000 1476.915000 2.805000 ;
      RECT 1477.025000  1.445000 1477.195000 1.615000 ;
      RECT 1477.205000 -0.085000 1477.375000 0.085000 ;
      RECT 1477.205000  2.635000 1477.375000 2.805000 ;
      RECT 1477.665000 -0.085000 1477.835000 0.085000 ;
      RECT 1477.665000  2.635000 1477.835000 2.805000 ;
      RECT 1478.125000 -0.085000 1478.295000 0.085000 ;
      RECT 1478.125000  2.635000 1478.295000 2.805000 ;
      RECT 1478.585000 -0.085000 1478.755000 0.085000 ;
      RECT 1478.585000  2.635000 1478.755000 2.805000 ;
      RECT 1479.045000 -0.085000 1479.215000 0.085000 ;
      RECT 1479.045000  2.635000 1479.215000 2.805000 ;
      RECT 1479.505000 -0.085000 1479.675000 0.085000 ;
      RECT 1479.505000  2.635000 1479.675000 2.805000 ;
      RECT 1479.965000 -0.085000 1480.135000 0.085000 ;
      RECT 1479.965000  2.635000 1480.135000 2.805000 ;
      RECT 1480.425000 -0.085000 1480.595000 0.085000 ;
      RECT 1480.425000  2.635000 1480.595000 2.805000 ;
      RECT 1480.885000 -0.085000 1481.055000 0.085000 ;
      RECT 1480.885000  2.635000 1481.055000 2.805000 ;
      RECT 1481.345000 -0.085000 1481.515000 0.085000 ;
      RECT 1481.345000  2.635000 1481.515000 2.805000 ;
      RECT 1481.805000 -0.085000 1481.975000 0.085000 ;
      RECT 1481.805000  2.635000 1481.975000 2.805000 ;
      RECT 1481.840000  1.105000 1482.010000 1.275000 ;
      RECT 1482.265000 -0.085000 1482.435000 0.085000 ;
      RECT 1482.265000  2.635000 1482.435000 2.805000 ;
      RECT 1482.725000 -0.085000 1482.895000 0.085000 ;
      RECT 1482.725000  2.635000 1482.895000 2.805000 ;
      RECT 1482.875000  1.445000 1483.045000 1.615000 ;
      RECT 1483.185000 -0.085000 1483.355000 0.085000 ;
      RECT 1483.185000  2.635000 1483.355000 2.805000 ;
      RECT 1483.645000 -0.085000 1483.815000 0.085000 ;
      RECT 1483.645000  2.635000 1483.815000 2.805000 ;
      RECT 1483.845000  1.105000 1484.015000 1.275000 ;
      RECT 1484.105000 -0.085000 1484.275000 0.085000 ;
      RECT 1484.105000  2.635000 1484.275000 2.805000 ;
      RECT 1484.565000 -0.085000 1484.735000 0.085000 ;
      RECT 1484.565000  2.635000 1484.735000 2.805000 ;
      RECT 1485.025000 -0.085000 1485.195000 0.085000 ;
      RECT 1485.025000  2.635000 1485.195000 2.805000 ;
      RECT 1485.325000  1.785000 1485.495000 1.955000 ;
      RECT 1485.485000 -0.085000 1485.655000 0.085000 ;
      RECT 1485.485000  2.635000 1485.655000 2.805000 ;
      RECT 1485.835000  1.100000 1486.005000 1.270000 ;
      RECT 1485.945000 -0.085000 1486.115000 0.085000 ;
      RECT 1485.945000  2.635000 1486.115000 2.805000 ;
      RECT 1486.210000  1.445000 1486.380000 1.615000 ;
      RECT 1486.405000 -0.085000 1486.575000 0.085000 ;
      RECT 1486.405000  2.635000 1486.575000 2.805000 ;
      RECT 1486.805000  1.785000 1486.975000 1.955000 ;
      RECT 1486.865000 -0.085000 1487.035000 0.085000 ;
      RECT 1486.865000  2.635000 1487.035000 2.805000 ;
      RECT 1487.325000 -0.085000 1487.495000 0.085000 ;
      RECT 1487.325000  2.635000 1487.495000 2.805000 ;
      RECT 1487.785000 -0.085000 1487.955000 0.085000 ;
      RECT 1487.785000  2.635000 1487.955000 2.805000 ;
      RECT 1488.245000 -0.085000 1488.415000 0.085000 ;
      RECT 1488.245000  2.635000 1488.415000 2.805000 ;
      RECT 1488.635000  1.445000 1488.805000 1.615000 ;
      RECT 1488.705000 -0.085000 1488.875000 0.085000 ;
      RECT 1488.705000  2.635000 1488.875000 2.805000 ;
      RECT 1489.165000 -0.085000 1489.335000 0.085000 ;
      RECT 1489.165000  2.635000 1489.335000 2.805000 ;
      RECT 1489.410000  1.785000 1489.580000 1.955000 ;
      RECT 1489.625000 -0.085000 1489.795000 0.085000 ;
      RECT 1489.625000  2.635000 1489.795000 2.805000 ;
      RECT 1490.085000 -0.085000 1490.255000 0.085000 ;
      RECT 1490.085000  2.635000 1490.255000 2.805000 ;
      RECT 1490.480000  1.105000 1490.650000 1.275000 ;
      RECT 1490.545000 -0.085000 1490.715000 0.085000 ;
      RECT 1490.545000  2.635000 1490.715000 2.805000 ;
      RECT 1490.990000  1.445000 1491.160000 1.615000 ;
      RECT 1491.005000 -0.085000 1491.175000 0.085000 ;
      RECT 1491.005000  2.635000 1491.175000 2.805000 ;
      RECT 1491.465000 -0.085000 1491.635000 0.085000 ;
      RECT 1491.465000  2.635000 1491.635000 2.805000 ;
      RECT 1491.925000 -0.085000 1492.095000 0.085000 ;
      RECT 1491.925000  2.635000 1492.095000 2.805000 ;
      RECT 1492.385000 -0.085000 1492.555000 0.085000 ;
      RECT 1492.385000  2.635000 1492.555000 2.805000 ;
      RECT 1492.845000 -0.085000 1493.015000 0.085000 ;
      RECT 1492.845000  2.635000 1493.015000 2.805000 ;
      RECT 1493.305000 -0.085000 1493.475000 0.085000 ;
      RECT 1493.305000  2.635000 1493.475000 2.805000 ;
      RECT 1493.765000 -0.085000 1493.935000 0.085000 ;
      RECT 1493.765000  2.635000 1493.935000 2.805000 ;
      RECT 1494.225000 -0.085000 1494.395000 0.085000 ;
      RECT 1494.225000  2.635000 1494.395000 2.805000 ;
      RECT 1494.685000 -0.085000 1494.855000 0.085000 ;
      RECT 1494.685000  2.635000 1494.855000 2.805000 ;
      RECT 1495.145000 -0.085000 1495.315000 0.085000 ;
      RECT 1495.145000  2.635000 1495.315000 2.805000 ;
      RECT 1495.605000 -0.085000 1495.775000 0.085000 ;
      RECT 1495.605000  2.635000 1495.775000 2.805000 ;
      RECT 1496.065000 -0.085000 1496.235000 0.085000 ;
      RECT 1496.065000  2.635000 1496.235000 2.805000 ;
      RECT 1496.525000 -0.085000 1496.695000 0.085000 ;
      RECT 1496.525000  2.635000 1496.695000 2.805000 ;
      RECT 1496.560000  1.105000 1496.730000 1.275000 ;
      RECT 1496.985000 -0.085000 1497.155000 0.085000 ;
      RECT 1496.985000  2.635000 1497.155000 2.805000 ;
      RECT 1497.445000 -0.085000 1497.615000 0.085000 ;
      RECT 1497.445000  2.635000 1497.615000 2.805000 ;
      RECT 1497.595000  1.445000 1497.765000 1.615000 ;
      RECT 1497.905000 -0.085000 1498.075000 0.085000 ;
      RECT 1497.905000  2.635000 1498.075000 2.805000 ;
      RECT 1498.365000 -0.085000 1498.535000 0.085000 ;
      RECT 1498.365000  2.635000 1498.535000 2.805000 ;
      RECT 1498.565000  1.105000 1498.735000 1.275000 ;
      RECT 1498.825000 -0.085000 1498.995000 0.085000 ;
      RECT 1498.825000  2.635000 1498.995000 2.805000 ;
      RECT 1499.285000 -0.085000 1499.455000 0.085000 ;
      RECT 1499.285000  2.635000 1499.455000 2.805000 ;
      RECT 1499.745000 -0.085000 1499.915000 0.085000 ;
      RECT 1499.745000  2.635000 1499.915000 2.805000 ;
      RECT 1500.045000  1.785000 1500.215000 1.955000 ;
      RECT 1500.205000 -0.085000 1500.375000 0.085000 ;
      RECT 1500.205000  2.635000 1500.375000 2.805000 ;
      RECT 1500.555000  1.100000 1500.725000 1.270000 ;
      RECT 1500.665000 -0.085000 1500.835000 0.085000 ;
      RECT 1500.665000  2.635000 1500.835000 2.805000 ;
      RECT 1500.930000  1.445000 1501.100000 1.615000 ;
      RECT 1501.125000 -0.085000 1501.295000 0.085000 ;
      RECT 1501.125000  2.635000 1501.295000 2.805000 ;
      RECT 1501.525000  1.785000 1501.695000 1.955000 ;
      RECT 1501.585000 -0.085000 1501.755000 0.085000 ;
      RECT 1501.585000  2.635000 1501.755000 2.805000 ;
      RECT 1502.045000 -0.085000 1502.215000 0.085000 ;
      RECT 1502.045000  2.635000 1502.215000 2.805000 ;
      RECT 1502.505000 -0.085000 1502.675000 0.085000 ;
      RECT 1502.505000  2.635000 1502.675000 2.805000 ;
      RECT 1502.965000 -0.085000 1503.135000 0.085000 ;
      RECT 1502.965000  2.635000 1503.135000 2.805000 ;
      RECT 1503.355000  1.445000 1503.525000 1.615000 ;
      RECT 1503.425000 -0.085000 1503.595000 0.085000 ;
      RECT 1503.425000  2.635000 1503.595000 2.805000 ;
      RECT 1503.885000 -0.085000 1504.055000 0.085000 ;
      RECT 1503.885000  2.635000 1504.055000 2.805000 ;
      RECT 1504.130000  1.785000 1504.300000 1.955000 ;
      RECT 1504.345000 -0.085000 1504.515000 0.085000 ;
      RECT 1504.345000  2.635000 1504.515000 2.805000 ;
      RECT 1504.805000 -0.085000 1504.975000 0.085000 ;
      RECT 1504.805000  2.635000 1504.975000 2.805000 ;
      RECT 1505.200000  1.105000 1505.370000 1.275000 ;
      RECT 1505.265000 -0.085000 1505.435000 0.085000 ;
      RECT 1505.265000  2.635000 1505.435000 2.805000 ;
      RECT 1505.710000  1.445000 1505.880000 1.615000 ;
      RECT 1505.725000 -0.085000 1505.895000 0.085000 ;
      RECT 1505.725000  2.635000 1505.895000 2.805000 ;
      RECT 1506.185000 -0.085000 1506.355000 0.085000 ;
      RECT 1506.185000  2.635000 1506.355000 2.805000 ;
      RECT 1506.645000 -0.085000 1506.815000 0.085000 ;
      RECT 1506.645000  2.635000 1506.815000 2.805000 ;
      RECT 1507.105000 -0.085000 1507.275000 0.085000 ;
      RECT 1507.105000  2.635000 1507.275000 2.805000 ;
      RECT 1507.565000 -0.085000 1507.735000 0.085000 ;
      RECT 1507.565000  2.635000 1507.735000 2.805000 ;
      RECT 1508.025000 -0.085000 1508.195000 0.085000 ;
      RECT 1508.025000  2.635000 1508.195000 2.805000 ;
      RECT 1508.485000 -0.085000 1508.655000 0.085000 ;
      RECT 1508.485000  2.635000 1508.655000 2.805000 ;
      RECT 1508.945000 -0.085000 1509.115000 0.085000 ;
      RECT 1508.945000  2.635000 1509.115000 2.805000 ;
      RECT 1509.405000 -0.085000 1509.575000 0.085000 ;
      RECT 1509.405000  2.635000 1509.575000 2.805000 ;
      RECT 1509.865000 -0.085000 1510.035000 0.085000 ;
      RECT 1509.865000  2.635000 1510.035000 2.805000 ;
      RECT 1510.325000 -0.085000 1510.495000 0.085000 ;
      RECT 1510.325000  2.635000 1510.495000 2.805000 ;
      RECT 1510.785000 -0.085000 1510.955000 0.085000 ;
      RECT 1510.785000  2.635000 1510.955000 2.805000 ;
      RECT 1511.245000 -0.085000 1511.415000 0.085000 ;
      RECT 1511.245000  2.635000 1511.415000 2.805000 ;
      RECT 1511.705000 -0.085000 1511.875000 0.085000 ;
      RECT 1511.705000  2.635000 1511.875000 2.805000 ;
      RECT 1512.165000 -0.085000 1512.335000 0.085000 ;
      RECT 1512.165000  2.635000 1512.335000 2.805000 ;
      RECT 1512.255000  1.785000 1512.425000 1.955000 ;
      RECT 1512.625000 -0.085000 1512.795000 0.085000 ;
      RECT 1512.625000  2.635000 1512.795000 2.805000 ;
      RECT 1512.675000  0.425000 1512.845000 0.595000 ;
      RECT 1513.085000 -0.085000 1513.255000 0.085000 ;
      RECT 1513.085000  2.635000 1513.255000 2.805000 ;
      RECT 1513.545000 -0.085000 1513.715000 0.085000 ;
      RECT 1513.545000  2.635000 1513.715000 2.805000 ;
      RECT 1514.005000 -0.085000 1514.175000 0.085000 ;
      RECT 1514.005000  2.635000 1514.175000 2.805000 ;
      RECT 1514.465000 -0.085000 1514.635000 0.085000 ;
      RECT 1514.465000  2.635000 1514.635000 2.805000 ;
      RECT 1514.925000 -0.085000 1515.095000 0.085000 ;
      RECT 1514.925000  2.635000 1515.095000 2.805000 ;
      RECT 1515.385000 -0.085000 1515.555000 0.085000 ;
      RECT 1515.385000  2.635000 1515.555000 2.805000 ;
      RECT 1515.845000 -0.085000 1516.015000 0.085000 ;
      RECT 1515.845000  2.635000 1516.015000 2.805000 ;
      RECT 1516.305000 -0.085000 1516.475000 0.085000 ;
      RECT 1516.305000  2.635000 1516.475000 2.805000 ;
      RECT 1516.765000 -0.085000 1516.935000 0.085000 ;
      RECT 1516.765000  0.765000 1516.935000 0.935000 ;
      RECT 1516.765000  2.635000 1516.935000 2.805000 ;
      RECT 1517.175000  1.785000 1517.345000 1.955000 ;
      RECT 1517.225000 -0.085000 1517.395000 0.085000 ;
      RECT 1517.225000  2.635000 1517.395000 2.805000 ;
      RECT 1517.685000 -0.085000 1517.855000 0.085000 ;
      RECT 1517.685000  2.635000 1517.855000 2.805000 ;
      RECT 1518.145000 -0.085000 1518.315000 0.085000 ;
      RECT 1518.145000  2.635000 1518.315000 2.805000 ;
      RECT 1518.605000 -0.085000 1518.775000 0.085000 ;
      RECT 1518.605000  2.635000 1518.775000 2.805000 ;
      RECT 1518.735000  1.785000 1518.905000 1.955000 ;
      RECT 1518.745000  0.765000 1518.915000 0.935000 ;
      RECT 1519.065000 -0.085000 1519.235000 0.085000 ;
      RECT 1519.065000  2.635000 1519.235000 2.805000 ;
      RECT 1519.525000 -0.085000 1519.695000 0.085000 ;
      RECT 1519.525000  2.635000 1519.695000 2.805000 ;
      RECT 1519.985000 -0.085000 1520.155000 0.085000 ;
      RECT 1519.985000  2.635000 1520.155000 2.805000 ;
      RECT 1520.445000 -0.085000 1520.615000 0.085000 ;
      RECT 1520.445000  2.635000 1520.615000 2.805000 ;
      RECT 1520.905000 -0.085000 1521.075000 0.085000 ;
      RECT 1520.905000  2.635000 1521.075000 2.805000 ;
      RECT 1521.365000 -0.085000 1521.535000 0.085000 ;
      RECT 1521.365000  2.635000 1521.535000 2.805000 ;
      RECT 1521.825000 -0.085000 1521.995000 0.085000 ;
      RECT 1521.825000  2.635000 1521.995000 2.805000 ;
      RECT 1522.285000 -0.085000 1522.455000 0.085000 ;
      RECT 1522.285000  2.635000 1522.455000 2.805000 ;
      RECT 1522.745000 -0.085000 1522.915000 0.085000 ;
      RECT 1522.745000  2.635000 1522.915000 2.805000 ;
      RECT 1523.205000 -0.085000 1523.375000 0.085000 ;
      RECT 1523.205000  2.635000 1523.375000 2.805000 ;
      RECT 1523.665000 -0.085000 1523.835000 0.085000 ;
      RECT 1523.665000  2.635000 1523.835000 2.805000 ;
      RECT 1524.125000 -0.085000 1524.295000 0.085000 ;
      RECT 1524.125000  2.635000 1524.295000 2.805000 ;
      RECT 1524.585000 -0.085000 1524.755000 0.085000 ;
      RECT 1524.585000  2.635000 1524.755000 2.805000 ;
      RECT 1524.675000  1.785000 1524.845000 1.955000 ;
      RECT 1525.045000 -0.085000 1525.215000 0.085000 ;
      RECT 1525.045000  2.635000 1525.215000 2.805000 ;
      RECT 1525.095000  0.425000 1525.265000 0.595000 ;
      RECT 1525.505000 -0.085000 1525.675000 0.085000 ;
      RECT 1525.505000  2.635000 1525.675000 2.805000 ;
      RECT 1525.965000 -0.085000 1526.135000 0.085000 ;
      RECT 1525.965000  2.635000 1526.135000 2.805000 ;
      RECT 1526.425000 -0.085000 1526.595000 0.085000 ;
      RECT 1526.425000  2.635000 1526.595000 2.805000 ;
      RECT 1526.885000 -0.085000 1527.055000 0.085000 ;
      RECT 1526.885000  2.635000 1527.055000 2.805000 ;
      RECT 1527.345000 -0.085000 1527.515000 0.085000 ;
      RECT 1527.345000  2.635000 1527.515000 2.805000 ;
      RECT 1527.805000 -0.085000 1527.975000 0.085000 ;
      RECT 1527.805000  2.635000 1527.975000 2.805000 ;
      RECT 1528.265000 -0.085000 1528.435000 0.085000 ;
      RECT 1528.265000  2.635000 1528.435000 2.805000 ;
      RECT 1528.725000 -0.085000 1528.895000 0.085000 ;
      RECT 1528.725000  2.635000 1528.895000 2.805000 ;
      RECT 1529.125000  0.765000 1529.295000 0.935000 ;
      RECT 1529.185000 -0.085000 1529.355000 0.085000 ;
      RECT 1529.185000  2.635000 1529.355000 2.805000 ;
      RECT 1529.595000  1.785000 1529.765000 1.955000 ;
      RECT 1529.645000 -0.085000 1529.815000 0.085000 ;
      RECT 1529.645000  2.635000 1529.815000 2.805000 ;
      RECT 1530.105000 -0.085000 1530.275000 0.085000 ;
      RECT 1530.105000  2.635000 1530.275000 2.805000 ;
      RECT 1530.565000 -0.085000 1530.735000 0.085000 ;
      RECT 1530.565000  2.635000 1530.735000 2.805000 ;
      RECT 1531.025000 -0.085000 1531.195000 0.085000 ;
      RECT 1531.025000  2.635000 1531.195000 2.805000 ;
      RECT 1531.155000  1.785000 1531.325000 1.955000 ;
      RECT 1531.165000  0.765000 1531.335000 0.935000 ;
      RECT 1531.485000 -0.085000 1531.655000 0.085000 ;
      RECT 1531.485000  2.635000 1531.655000 2.805000 ;
      RECT 1531.945000 -0.085000 1532.115000 0.085000 ;
      RECT 1531.945000  2.635000 1532.115000 2.805000 ;
      RECT 1532.405000 -0.085000 1532.575000 0.085000 ;
      RECT 1532.405000  2.635000 1532.575000 2.805000 ;
      RECT 1532.865000 -0.085000 1533.035000 0.085000 ;
      RECT 1532.865000  2.635000 1533.035000 2.805000 ;
      RECT 1533.325000 -0.085000 1533.495000 0.085000 ;
      RECT 1533.325000  2.635000 1533.495000 2.805000 ;
      RECT 1533.785000 -0.085000 1533.955000 0.085000 ;
      RECT 1533.785000  2.635000 1533.955000 2.805000 ;
      RECT 1534.245000 -0.085000 1534.415000 0.085000 ;
      RECT 1534.245000  2.635000 1534.415000 2.805000 ;
      RECT 1534.705000 -0.085000 1534.875000 0.085000 ;
      RECT 1534.705000  2.635000 1534.875000 2.805000 ;
      RECT 1535.165000 -0.085000 1535.335000 0.085000 ;
      RECT 1535.165000  2.635000 1535.335000 2.805000 ;
      RECT 1535.625000 -0.085000 1535.795000 0.085000 ;
      RECT 1535.625000  2.635000 1535.795000 2.805000 ;
      RECT 1536.085000 -0.085000 1536.255000 0.085000 ;
      RECT 1536.085000  2.635000 1536.255000 2.805000 ;
      RECT 1536.545000 -0.085000 1536.715000 0.085000 ;
      RECT 1536.545000  2.635000 1536.715000 2.805000 ;
      RECT 1537.005000 -0.085000 1537.175000 0.085000 ;
      RECT 1537.005000  2.635000 1537.175000 2.805000 ;
      RECT 1537.465000 -0.085000 1537.635000 0.085000 ;
      RECT 1537.465000  2.635000 1537.635000 2.805000 ;
      RECT 1537.925000 -0.085000 1538.095000 0.085000 ;
      RECT 1537.925000  2.635000 1538.095000 2.805000 ;
      RECT 1538.385000 -0.085000 1538.555000 0.085000 ;
      RECT 1538.385000  2.635000 1538.555000 2.805000 ;
      RECT 1538.445000  1.740000 1538.615000 1.910000 ;
      RECT 1538.845000 -0.085000 1539.015000 0.085000 ;
      RECT 1538.845000  2.635000 1539.015000 2.805000 ;
      RECT 1538.935000  0.720000 1539.105000 0.890000 ;
      RECT 1539.305000 -0.085000 1539.475000 0.085000 ;
      RECT 1539.305000  2.635000 1539.475000 2.805000 ;
      RECT 1539.765000 -0.085000 1539.935000 0.085000 ;
      RECT 1539.765000  2.635000 1539.935000 2.805000 ;
      RECT 1540.225000 -0.085000 1540.395000 0.085000 ;
      RECT 1540.225000  2.635000 1540.395000 2.805000 ;
      RECT 1540.685000 -0.085000 1540.855000 0.085000 ;
      RECT 1540.685000  2.635000 1540.855000 2.805000 ;
      RECT 1541.145000 -0.085000 1541.315000 0.085000 ;
      RECT 1541.145000  2.635000 1541.315000 2.805000 ;
      RECT 1541.605000 -0.085000 1541.775000 0.085000 ;
      RECT 1541.605000  2.635000 1541.775000 2.805000 ;
      RECT 1542.065000 -0.085000 1542.235000 0.085000 ;
      RECT 1542.065000  2.635000 1542.235000 2.805000 ;
      RECT 1542.525000 -0.085000 1542.695000 0.085000 ;
      RECT 1542.525000  2.635000 1542.695000 2.805000 ;
      RECT 1542.935000  0.720000 1543.105000 0.890000 ;
      RECT 1542.985000 -0.085000 1543.155000 0.085000 ;
      RECT 1542.985000  2.635000 1543.155000 2.805000 ;
      RECT 1543.445000 -0.085000 1543.615000 0.085000 ;
      RECT 1543.445000  1.740000 1543.615000 1.910000 ;
      RECT 1543.445000  2.635000 1543.615000 2.805000 ;
      RECT 1543.905000 -0.085000 1544.075000 0.085000 ;
      RECT 1543.905000  2.635000 1544.075000 2.805000 ;
      RECT 1544.365000 -0.085000 1544.535000 0.085000 ;
      RECT 1544.365000  2.635000 1544.535000 2.805000 ;
      RECT 1544.825000 -0.085000 1544.995000 0.085000 ;
      RECT 1544.825000  2.635000 1544.995000 2.805000 ;
      RECT 1545.020000  1.740000 1545.190000 1.910000 ;
      RECT 1545.090000  0.720000 1545.260000 0.890000 ;
      RECT 1545.285000 -0.085000 1545.455000 0.085000 ;
      RECT 1545.285000  2.635000 1545.455000 2.805000 ;
      RECT 1545.745000 -0.085000 1545.915000 0.085000 ;
      RECT 1545.745000  2.635000 1545.915000 2.805000 ;
      RECT 1546.205000 -0.085000 1546.375000 0.085000 ;
      RECT 1546.205000  2.635000 1546.375000 2.805000 ;
      RECT 1546.665000 -0.085000 1546.835000 0.085000 ;
      RECT 1546.665000  2.635000 1546.835000 2.805000 ;
      RECT 1547.125000 -0.085000 1547.295000 0.085000 ;
      RECT 1547.125000  2.635000 1547.295000 2.805000 ;
      RECT 1547.585000 -0.085000 1547.755000 0.085000 ;
      RECT 1547.585000  2.635000 1547.755000 2.805000 ;
      RECT 1548.045000 -0.085000 1548.215000 0.085000 ;
      RECT 1548.045000  2.635000 1548.215000 2.805000 ;
      RECT 1548.505000 -0.085000 1548.675000 0.085000 ;
      RECT 1548.505000  2.635000 1548.675000 2.805000 ;
      RECT 1548.965000 -0.085000 1549.135000 0.085000 ;
      RECT 1548.965000  2.635000 1549.135000 2.805000 ;
      RECT 1549.425000 -0.085000 1549.595000 0.085000 ;
      RECT 1549.425000  2.635000 1549.595000 2.805000 ;
      RECT 1549.485000  1.740000 1549.655000 1.910000 ;
      RECT 1549.885000 -0.085000 1550.055000 0.085000 ;
      RECT 1549.885000  2.635000 1550.055000 2.805000 ;
      RECT 1549.975000  0.720000 1550.145000 0.890000 ;
      RECT 1550.345000 -0.085000 1550.515000 0.085000 ;
      RECT 1550.345000  2.635000 1550.515000 2.805000 ;
      RECT 1550.805000 -0.085000 1550.975000 0.085000 ;
      RECT 1550.805000  2.635000 1550.975000 2.805000 ;
      RECT 1551.265000 -0.085000 1551.435000 0.085000 ;
      RECT 1551.265000  2.635000 1551.435000 2.805000 ;
      RECT 1551.725000 -0.085000 1551.895000 0.085000 ;
      RECT 1551.725000  2.635000 1551.895000 2.805000 ;
      RECT 1552.185000 -0.085000 1552.355000 0.085000 ;
      RECT 1552.185000  2.635000 1552.355000 2.805000 ;
      RECT 1552.645000 -0.085000 1552.815000 0.085000 ;
      RECT 1552.645000  2.635000 1552.815000 2.805000 ;
      RECT 1553.105000 -0.085000 1553.275000 0.085000 ;
      RECT 1553.105000  2.635000 1553.275000 2.805000 ;
      RECT 1553.565000 -0.085000 1553.735000 0.085000 ;
      RECT 1553.565000  2.635000 1553.735000 2.805000 ;
      RECT 1553.975000  0.720000 1554.145000 0.890000 ;
      RECT 1554.025000 -0.085000 1554.195000 0.085000 ;
      RECT 1554.025000  2.635000 1554.195000 2.805000 ;
      RECT 1554.485000 -0.085000 1554.655000 0.085000 ;
      RECT 1554.485000  1.740000 1554.655000 1.910000 ;
      RECT 1554.485000  2.635000 1554.655000 2.805000 ;
      RECT 1554.945000 -0.085000 1555.115000 0.085000 ;
      RECT 1554.945000  2.635000 1555.115000 2.805000 ;
      RECT 1555.405000 -0.085000 1555.575000 0.085000 ;
      RECT 1555.405000  2.635000 1555.575000 2.805000 ;
      RECT 1555.865000 -0.085000 1556.035000 0.085000 ;
      RECT 1555.865000  2.635000 1556.035000 2.805000 ;
      RECT 1556.045000  0.720000 1556.215000 0.890000 ;
      RECT 1556.045000  1.740000 1556.215000 1.910000 ;
      RECT 1556.325000 -0.085000 1556.495000 0.085000 ;
      RECT 1556.325000  2.635000 1556.495000 2.805000 ;
      RECT 1556.785000 -0.085000 1556.955000 0.085000 ;
      RECT 1556.785000  2.635000 1556.955000 2.805000 ;
      RECT 1557.245000 -0.085000 1557.415000 0.085000 ;
      RECT 1557.245000  2.635000 1557.415000 2.805000 ;
      RECT 1557.705000 -0.085000 1557.875000 0.085000 ;
      RECT 1557.705000  2.635000 1557.875000 2.805000 ;
      RECT 1558.165000 -0.085000 1558.335000 0.085000 ;
      RECT 1558.165000  2.635000 1558.335000 2.805000 ;
      RECT 1558.625000 -0.085000 1558.795000 0.085000 ;
      RECT 1558.625000  2.635000 1558.795000 2.805000 ;
      RECT 1559.085000 -0.085000 1559.255000 0.085000 ;
      RECT 1559.085000  2.635000 1559.255000 2.805000 ;
      RECT 1559.545000 -0.085000 1559.715000 0.085000 ;
      RECT 1559.545000  2.635000 1559.715000 2.805000 ;
      RECT 1560.005000 -0.085000 1560.175000 0.085000 ;
      RECT 1560.005000  2.635000 1560.175000 2.805000 ;
      RECT 1560.465000 -0.085000 1560.635000 0.085000 ;
      RECT 1560.465000  2.635000 1560.635000 2.805000 ;
      RECT 1560.925000 -0.085000 1561.095000 0.085000 ;
      RECT 1560.925000  2.635000 1561.095000 2.805000 ;
      RECT 1560.985000  1.740000 1561.155000 1.910000 ;
      RECT 1561.385000 -0.085000 1561.555000 0.085000 ;
      RECT 1561.385000  2.635000 1561.555000 2.805000 ;
      RECT 1561.475000  0.720000 1561.645000 0.890000 ;
      RECT 1561.845000 -0.085000 1562.015000 0.085000 ;
      RECT 1561.845000  2.635000 1562.015000 2.805000 ;
      RECT 1562.305000 -0.085000 1562.475000 0.085000 ;
      RECT 1562.305000  2.635000 1562.475000 2.805000 ;
      RECT 1562.765000 -0.085000 1562.935000 0.085000 ;
      RECT 1562.765000  2.635000 1562.935000 2.805000 ;
      RECT 1563.225000 -0.085000 1563.395000 0.085000 ;
      RECT 1563.225000  2.635000 1563.395000 2.805000 ;
      RECT 1563.685000 -0.085000 1563.855000 0.085000 ;
      RECT 1563.685000  2.635000 1563.855000 2.805000 ;
      RECT 1564.145000 -0.085000 1564.315000 0.085000 ;
      RECT 1564.145000  2.635000 1564.315000 2.805000 ;
      RECT 1564.605000 -0.085000 1564.775000 0.085000 ;
      RECT 1564.605000  2.635000 1564.775000 2.805000 ;
      RECT 1565.065000 -0.085000 1565.235000 0.085000 ;
      RECT 1565.065000  2.635000 1565.235000 2.805000 ;
      RECT 1565.475000  0.720000 1565.645000 0.890000 ;
      RECT 1565.525000 -0.085000 1565.695000 0.085000 ;
      RECT 1565.525000  2.635000 1565.695000 2.805000 ;
      RECT 1565.985000 -0.085000 1566.155000 0.085000 ;
      RECT 1565.985000  1.740000 1566.155000 1.910000 ;
      RECT 1565.985000  2.635000 1566.155000 2.805000 ;
      RECT 1566.445000 -0.085000 1566.615000 0.085000 ;
      RECT 1566.445000  2.635000 1566.615000 2.805000 ;
      RECT 1566.905000 -0.085000 1567.075000 0.085000 ;
      RECT 1566.905000  2.635000 1567.075000 2.805000 ;
      RECT 1567.365000 -0.085000 1567.535000 0.085000 ;
      RECT 1567.365000  2.635000 1567.535000 2.805000 ;
      RECT 1567.545000  0.720000 1567.715000 0.890000 ;
      RECT 1567.545000  1.740000 1567.715000 1.910000 ;
      RECT 1567.825000 -0.085000 1567.995000 0.085000 ;
      RECT 1567.825000  2.635000 1567.995000 2.805000 ;
      RECT 1568.285000 -0.085000 1568.455000 0.085000 ;
      RECT 1568.285000  2.635000 1568.455000 2.805000 ;
      RECT 1568.745000 -0.085000 1568.915000 0.085000 ;
      RECT 1568.745000  2.635000 1568.915000 2.805000 ;
      RECT 1569.205000 -0.085000 1569.375000 0.085000 ;
      RECT 1569.205000  2.635000 1569.375000 2.805000 ;
      RECT 1569.665000 -0.085000 1569.835000 0.085000 ;
      RECT 1569.665000  2.635000 1569.835000 2.805000 ;
      RECT 1570.125000 -0.085000 1570.295000 0.085000 ;
      RECT 1570.125000  2.635000 1570.295000 2.805000 ;
      RECT 1570.585000 -0.085000 1570.755000 0.085000 ;
      RECT 1570.585000  2.635000 1570.755000 2.805000 ;
      RECT 1571.045000 -0.085000 1571.215000 0.085000 ;
      RECT 1571.045000  2.635000 1571.215000 2.805000 ;
      RECT 1571.505000 -0.085000 1571.675000 0.085000 ;
      RECT 1571.505000  2.635000 1571.675000 2.805000 ;
      RECT 1571.965000 -0.085000 1572.135000 0.085000 ;
      RECT 1571.965000  2.635000 1572.135000 2.805000 ;
      RECT 1572.425000 -0.085000 1572.595000 0.085000 ;
      RECT 1572.425000  2.635000 1572.595000 2.805000 ;
      RECT 1572.885000 -0.085000 1573.055000 0.085000 ;
      RECT 1572.885000  2.635000 1573.055000 2.805000 ;
      RECT 1573.345000 -0.085000 1573.515000 0.085000 ;
      RECT 1573.345000  2.635000 1573.515000 2.805000 ;
      RECT 1573.805000 -0.085000 1573.975000 0.085000 ;
      RECT 1573.805000  2.635000 1573.975000 2.805000 ;
      RECT 1574.265000 -0.085000 1574.435000 0.085000 ;
      RECT 1574.265000  2.635000 1574.435000 2.805000 ;
      RECT 1574.365000  1.445000 1574.535000 1.615000 ;
      RECT 1574.725000 -0.085000 1574.895000 0.085000 ;
      RECT 1574.725000  2.635000 1574.895000 2.805000 ;
      RECT 1574.875000  0.765000 1575.045000 0.935000 ;
      RECT 1575.185000 -0.085000 1575.355000 0.085000 ;
      RECT 1575.185000  2.635000 1575.355000 2.805000 ;
      RECT 1575.645000 -0.085000 1575.815000 0.085000 ;
      RECT 1575.645000  2.635000 1575.815000 2.805000 ;
      RECT 1576.105000 -0.085000 1576.275000 0.085000 ;
      RECT 1576.105000  2.635000 1576.275000 2.805000 ;
      RECT 1576.540000  0.765000 1576.710000 0.935000 ;
      RECT 1576.565000 -0.085000 1576.735000 0.085000 ;
      RECT 1576.565000  2.635000 1576.735000 2.805000 ;
      RECT 1577.025000 -0.085000 1577.195000 0.085000 ;
      RECT 1577.025000  2.635000 1577.195000 2.805000 ;
      RECT 1577.105000  1.445000 1577.275000 1.615000 ;
      RECT 1577.485000 -0.085000 1577.655000 0.085000 ;
      RECT 1577.485000  2.635000 1577.655000 2.805000 ;
      RECT 1577.545000  1.105000 1577.715000 1.275000 ;
      RECT 1577.945000 -0.085000 1578.115000 0.085000 ;
      RECT 1577.945000  2.635000 1578.115000 2.805000 ;
      RECT 1578.405000 -0.085000 1578.575000 0.085000 ;
      RECT 1578.405000  2.635000 1578.575000 2.805000 ;
      RECT 1578.740000  1.105000 1578.910000 1.275000 ;
      RECT 1578.865000 -0.085000 1579.035000 0.085000 ;
      RECT 1578.865000  2.635000 1579.035000 2.805000 ;
      RECT 1579.325000 -0.085000 1579.495000 0.085000 ;
      RECT 1579.325000  2.635000 1579.495000 2.805000 ;
      RECT 1579.785000 -0.085000 1579.955000 0.085000 ;
      RECT 1579.785000  2.635000 1579.955000 2.805000 ;
      RECT 1580.245000 -0.085000 1580.415000 0.085000 ;
      RECT 1580.245000  2.635000 1580.415000 2.805000 ;
      RECT 1580.705000 -0.085000 1580.875000 0.085000 ;
      RECT 1580.705000  2.635000 1580.875000 2.805000 ;
      RECT 1581.165000 -0.085000 1581.335000 0.085000 ;
      RECT 1581.165000  2.635000 1581.335000 2.805000 ;
      RECT 1581.625000 -0.085000 1581.795000 0.085000 ;
      RECT 1581.625000  2.635000 1581.795000 2.805000 ;
      RECT 1582.085000 -0.085000 1582.255000 0.085000 ;
      RECT 1582.085000  2.635000 1582.255000 2.805000 ;
      RECT 1582.185000  1.445000 1582.355000 1.615000 ;
      RECT 1582.545000 -0.085000 1582.715000 0.085000 ;
      RECT 1582.545000  2.635000 1582.715000 2.805000 ;
      RECT 1582.695000  0.765000 1582.865000 0.935000 ;
      RECT 1583.005000 -0.085000 1583.175000 0.085000 ;
      RECT 1583.005000  2.635000 1583.175000 2.805000 ;
      RECT 1583.465000 -0.085000 1583.635000 0.085000 ;
      RECT 1583.465000  2.635000 1583.635000 2.805000 ;
      RECT 1583.925000 -0.085000 1584.095000 0.085000 ;
      RECT 1583.925000  2.635000 1584.095000 2.805000 ;
      RECT 1584.385000 -0.085000 1584.555000 0.085000 ;
      RECT 1584.385000  2.635000 1584.555000 2.805000 ;
      RECT 1584.550000  0.765000 1584.720000 0.935000 ;
      RECT 1584.845000 -0.085000 1585.015000 0.085000 ;
      RECT 1584.845000  2.635000 1585.015000 2.805000 ;
      RECT 1585.060000  1.445000 1585.230000 1.615000 ;
      RECT 1585.305000 -0.085000 1585.475000 0.085000 ;
      RECT 1585.305000  2.635000 1585.475000 2.805000 ;
      RECT 1585.570000  1.105000 1585.740000 1.275000 ;
      RECT 1585.765000 -0.085000 1585.935000 0.085000 ;
      RECT 1585.765000  2.635000 1585.935000 2.805000 ;
      RECT 1586.225000 -0.085000 1586.395000 0.085000 ;
      RECT 1586.225000  2.635000 1586.395000 2.805000 ;
      RECT 1586.560000  1.105000 1586.730000 1.275000 ;
      RECT 1586.685000 -0.085000 1586.855000 0.085000 ;
      RECT 1586.685000  2.635000 1586.855000 2.805000 ;
      RECT 1587.145000 -0.085000 1587.315000 0.085000 ;
      RECT 1587.145000  2.635000 1587.315000 2.805000 ;
      RECT 1587.605000 -0.085000 1587.775000 0.085000 ;
      RECT 1587.605000  2.635000 1587.775000 2.805000 ;
      RECT 1588.065000 -0.085000 1588.235000 0.085000 ;
      RECT 1588.065000  2.635000 1588.235000 2.805000 ;
      RECT 1588.525000 -0.085000 1588.695000 0.085000 ;
      RECT 1588.525000  2.635000 1588.695000 2.805000 ;
      RECT 1588.985000 -0.085000 1589.155000 0.085000 ;
      RECT 1588.985000  2.635000 1589.155000 2.805000 ;
      RECT 1589.445000 -0.085000 1589.615000 0.085000 ;
      RECT 1589.445000  2.635000 1589.615000 2.805000 ;
      RECT 1589.905000 -0.085000 1590.075000 0.085000 ;
      RECT 1589.905000  2.635000 1590.075000 2.805000 ;
      RECT 1590.365000 -0.085000 1590.535000 0.085000 ;
      RECT 1590.365000  2.635000 1590.535000 2.805000 ;
      RECT 1590.520000  1.445000 1590.690000 1.615000 ;
      RECT 1590.825000 -0.085000 1590.995000 0.085000 ;
      RECT 1590.825000  2.635000 1590.995000 2.805000 ;
      RECT 1591.030000  0.765000 1591.200000 0.935000 ;
      RECT 1591.285000 -0.085000 1591.455000 0.085000 ;
      RECT 1591.285000  2.635000 1591.455000 2.805000 ;
      RECT 1591.745000 -0.085000 1591.915000 0.085000 ;
      RECT 1591.745000  2.635000 1591.915000 2.805000 ;
      RECT 1592.205000 -0.085000 1592.375000 0.085000 ;
      RECT 1592.205000  2.635000 1592.375000 2.805000 ;
      RECT 1592.665000 -0.085000 1592.835000 0.085000 ;
      RECT 1592.665000  2.635000 1592.835000 2.805000 ;
      RECT 1592.990000  0.765000 1593.160000 0.935000 ;
      RECT 1593.125000 -0.085000 1593.295000 0.085000 ;
      RECT 1593.125000  2.635000 1593.295000 2.805000 ;
      RECT 1593.500000  1.445000 1593.670000 1.615000 ;
      RECT 1593.585000 -0.085000 1593.755000 0.085000 ;
      RECT 1593.585000  2.635000 1593.755000 2.805000 ;
      RECT 1593.955000  1.105000 1594.125000 1.275000 ;
      RECT 1594.045000 -0.085000 1594.215000 0.085000 ;
      RECT 1594.045000  2.635000 1594.215000 2.805000 ;
      RECT 1594.505000 -0.085000 1594.675000 0.085000 ;
      RECT 1594.505000  2.635000 1594.675000 2.805000 ;
      RECT 1594.965000 -0.085000 1595.135000 0.085000 ;
      RECT 1594.965000  2.635000 1595.135000 2.805000 ;
      RECT 1595.000000  1.105000 1595.170000 1.275000 ;
      RECT 1595.425000 -0.085000 1595.595000 0.085000 ;
      RECT 1595.425000  2.635000 1595.595000 2.805000 ;
      RECT 1595.885000 -0.085000 1596.055000 0.085000 ;
      RECT 1595.885000  2.635000 1596.055000 2.805000 ;
      RECT 1596.345000 -0.085000 1596.515000 0.085000 ;
      RECT 1596.345000  2.635000 1596.515000 2.805000 ;
      RECT 1596.805000 -0.085000 1596.975000 0.085000 ;
      RECT 1596.805000  2.635000 1596.975000 2.805000 ;
      RECT 1597.265000 -0.085000 1597.435000 0.085000 ;
      RECT 1597.265000  2.635000 1597.435000 2.805000 ;
      RECT 1597.725000 -0.085000 1597.895000 0.085000 ;
      RECT 1597.725000  2.635000 1597.895000 2.805000 ;
      RECT 1598.185000 -0.085000 1598.355000 0.085000 ;
      RECT 1598.185000  2.635000 1598.355000 2.805000 ;
      RECT 1598.645000 -0.085000 1598.815000 0.085000 ;
      RECT 1598.645000  2.635000 1598.815000 2.805000 ;
      RECT 1599.105000 -0.085000 1599.275000 0.085000 ;
      RECT 1599.105000  2.635000 1599.275000 2.805000 ;
      RECT 1599.185000  1.785000 1599.355000 1.955000 ;
      RECT 1599.565000 -0.085000 1599.735000 0.085000 ;
      RECT 1599.565000  2.635000 1599.735000 2.805000 ;
      RECT 1599.615000  1.445000 1599.785000 1.615000 ;
      RECT 1599.955000  0.425000 1600.125000 0.595000 ;
      RECT 1600.025000 -0.085000 1600.195000 0.085000 ;
      RECT 1600.025000  2.635000 1600.195000 2.805000 ;
      RECT 1600.485000 -0.085000 1600.655000 0.085000 ;
      RECT 1600.485000  2.635000 1600.655000 2.805000 ;
      RECT 1600.945000 -0.085000 1601.115000 0.085000 ;
      RECT 1600.945000  2.635000 1601.115000 2.805000 ;
      RECT 1601.405000 -0.085000 1601.575000 0.085000 ;
      RECT 1601.405000  2.635000 1601.575000 2.805000 ;
      RECT 1601.865000 -0.085000 1602.035000 0.085000 ;
      RECT 1601.865000  2.635000 1602.035000 2.805000 ;
      RECT 1602.325000 -0.085000 1602.495000 0.085000 ;
      RECT 1602.325000  2.635000 1602.495000 2.805000 ;
      RECT 1602.605000  0.765000 1602.775000 0.935000 ;
      RECT 1602.785000 -0.085000 1602.955000 0.085000 ;
      RECT 1602.785000  2.635000 1602.955000 2.805000 ;
      RECT 1603.035000  0.425000 1603.205000 0.595000 ;
      RECT 1603.245000 -0.085000 1603.415000 0.085000 ;
      RECT 1603.245000  2.635000 1603.415000 2.805000 ;
      RECT 1603.515000  0.425000 1603.685000 0.595000 ;
      RECT 1603.705000 -0.085000 1603.875000 0.085000 ;
      RECT 1603.705000  2.635000 1603.875000 2.805000 ;
      RECT 1604.165000 -0.085000 1604.335000 0.085000 ;
      RECT 1604.165000  2.635000 1604.335000 2.805000 ;
      RECT 1604.625000 -0.085000 1604.795000 0.085000 ;
      RECT 1604.625000  2.635000 1604.795000 2.805000 ;
      RECT 1605.085000 -0.085000 1605.255000 0.085000 ;
      RECT 1605.085000  2.635000 1605.255000 2.805000 ;
      RECT 1605.545000 -0.085000 1605.715000 0.085000 ;
      RECT 1605.545000  2.635000 1605.715000 2.805000 ;
      RECT 1605.815000  0.425000 1605.985000 0.595000 ;
      RECT 1606.005000 -0.085000 1606.175000 0.085000 ;
      RECT 1606.005000  2.635000 1606.175000 2.805000 ;
      RECT 1606.410000  1.445000 1606.580000 1.615000 ;
      RECT 1606.465000 -0.085000 1606.635000 0.085000 ;
      RECT 1606.465000  2.635000 1606.635000 2.805000 ;
      RECT 1606.845000  1.785000 1607.015000 1.955000 ;
      RECT 1606.925000 -0.085000 1607.095000 0.085000 ;
      RECT 1606.925000  2.635000 1607.095000 2.805000 ;
      RECT 1607.385000 -0.085000 1607.555000 0.085000 ;
      RECT 1607.385000  2.635000 1607.555000 2.805000 ;
      RECT 1607.845000 -0.085000 1608.015000 0.085000 ;
      RECT 1607.845000  2.635000 1608.015000 2.805000 ;
      RECT 1608.305000 -0.085000 1608.475000 0.085000 ;
      RECT 1608.305000  2.635000 1608.475000 2.805000 ;
      RECT 1608.765000 -0.085000 1608.935000 0.085000 ;
      RECT 1608.765000  2.635000 1608.935000 2.805000 ;
      RECT 1609.225000 -0.085000 1609.395000 0.085000 ;
      RECT 1609.225000  2.635000 1609.395000 2.805000 ;
      RECT 1609.660000  1.785000 1609.830000 1.955000 ;
      RECT 1609.685000 -0.085000 1609.855000 0.085000 ;
      RECT 1609.685000  2.635000 1609.855000 2.805000 ;
      RECT 1610.130000  1.445000 1610.300000 1.615000 ;
      RECT 1610.145000 -0.085000 1610.315000 0.085000 ;
      RECT 1610.145000  2.635000 1610.315000 2.805000 ;
      RECT 1610.605000 -0.085000 1610.775000 0.085000 ;
      RECT 1610.605000  2.635000 1610.775000 2.805000 ;
      RECT 1610.665000  1.105000 1610.835000 1.275000 ;
      RECT 1611.065000 -0.085000 1611.235000 0.085000 ;
      RECT 1611.065000  2.635000 1611.235000 2.805000 ;
      RECT 1611.525000 -0.085000 1611.695000 0.085000 ;
      RECT 1611.525000  2.635000 1611.695000 2.805000 ;
      RECT 1611.985000 -0.085000 1612.155000 0.085000 ;
      RECT 1611.985000  2.635000 1612.155000 2.805000 ;
      RECT 1612.200000  0.765000 1612.370000 0.935000 ;
      RECT 1612.445000 -0.085000 1612.615000 0.085000 ;
      RECT 1612.445000  2.635000 1612.615000 2.805000 ;
      RECT 1612.695000  1.105000 1612.865000 1.275000 ;
      RECT 1612.905000 -0.085000 1613.075000 0.085000 ;
      RECT 1612.905000  2.635000 1613.075000 2.805000 ;
      RECT 1613.365000 -0.085000 1613.535000 0.085000 ;
      RECT 1613.365000  2.635000 1613.535000 2.805000 ;
      RECT 1613.825000 -0.085000 1613.995000 0.085000 ;
      RECT 1613.825000  2.635000 1613.995000 2.805000 ;
      RECT 1614.285000 -0.085000 1614.455000 0.085000 ;
      RECT 1614.285000  2.635000 1614.455000 2.805000 ;
      RECT 1614.745000 -0.085000 1614.915000 0.085000 ;
      RECT 1614.745000  2.635000 1614.915000 2.805000 ;
      RECT 1614.825000  1.785000 1614.995000 1.955000 ;
      RECT 1615.205000 -0.085000 1615.375000 0.085000 ;
      RECT 1615.205000  2.635000 1615.375000 2.805000 ;
      RECT 1615.255000  1.445000 1615.425000 1.615000 ;
      RECT 1615.595000  0.425000 1615.765000 0.595000 ;
      RECT 1615.665000 -0.085000 1615.835000 0.085000 ;
      RECT 1615.665000  2.635000 1615.835000 2.805000 ;
      RECT 1616.125000 -0.085000 1616.295000 0.085000 ;
      RECT 1616.125000  2.635000 1616.295000 2.805000 ;
      RECT 1616.585000 -0.085000 1616.755000 0.085000 ;
      RECT 1616.585000  2.635000 1616.755000 2.805000 ;
      RECT 1617.045000 -0.085000 1617.215000 0.085000 ;
      RECT 1617.045000  2.635000 1617.215000 2.805000 ;
      RECT 1617.505000 -0.085000 1617.675000 0.085000 ;
      RECT 1617.505000  2.635000 1617.675000 2.805000 ;
      RECT 1617.965000 -0.085000 1618.135000 0.085000 ;
      RECT 1617.965000  2.635000 1618.135000 2.805000 ;
      RECT 1618.245000  0.765000 1618.415000 0.935000 ;
      RECT 1618.425000 -0.085000 1618.595000 0.085000 ;
      RECT 1618.425000  2.635000 1618.595000 2.805000 ;
      RECT 1618.675000  0.425000 1618.845000 0.595000 ;
      RECT 1618.885000 -0.085000 1619.055000 0.085000 ;
      RECT 1618.885000  2.635000 1619.055000 2.805000 ;
      RECT 1619.155000  0.425000 1619.325000 0.595000 ;
      RECT 1619.345000 -0.085000 1619.515000 0.085000 ;
      RECT 1619.345000  2.635000 1619.515000 2.805000 ;
      RECT 1619.805000 -0.085000 1619.975000 0.085000 ;
      RECT 1619.805000  2.635000 1619.975000 2.805000 ;
      RECT 1620.265000 -0.085000 1620.435000 0.085000 ;
      RECT 1620.265000  2.635000 1620.435000 2.805000 ;
      RECT 1620.725000 -0.085000 1620.895000 0.085000 ;
      RECT 1620.725000  2.635000 1620.895000 2.805000 ;
      RECT 1621.185000 -0.085000 1621.355000 0.085000 ;
      RECT 1621.185000  2.635000 1621.355000 2.805000 ;
      RECT 1621.455000  0.425000 1621.625000 0.595000 ;
      RECT 1621.645000 -0.085000 1621.815000 0.085000 ;
      RECT 1621.645000  2.635000 1621.815000 2.805000 ;
      RECT 1622.050000  1.445000 1622.220000 1.615000 ;
      RECT 1622.105000 -0.085000 1622.275000 0.085000 ;
      RECT 1622.105000  2.635000 1622.275000 2.805000 ;
      RECT 1622.485000  1.785000 1622.655000 1.955000 ;
      RECT 1622.565000 -0.085000 1622.735000 0.085000 ;
      RECT 1622.565000  2.635000 1622.735000 2.805000 ;
      RECT 1623.025000 -0.085000 1623.195000 0.085000 ;
      RECT 1623.025000  2.635000 1623.195000 2.805000 ;
      RECT 1623.485000 -0.085000 1623.655000 0.085000 ;
      RECT 1623.485000  2.635000 1623.655000 2.805000 ;
      RECT 1623.945000 -0.085000 1624.115000 0.085000 ;
      RECT 1623.945000  2.635000 1624.115000 2.805000 ;
      RECT 1624.405000 -0.085000 1624.575000 0.085000 ;
      RECT 1624.405000  2.635000 1624.575000 2.805000 ;
      RECT 1624.865000 -0.085000 1625.035000 0.085000 ;
      RECT 1624.865000  2.635000 1625.035000 2.805000 ;
      RECT 1625.300000  1.785000 1625.470000 1.955000 ;
      RECT 1625.325000 -0.085000 1625.495000 0.085000 ;
      RECT 1625.325000  2.635000 1625.495000 2.805000 ;
      RECT 1625.770000  1.445000 1625.940000 1.615000 ;
      RECT 1625.785000 -0.085000 1625.955000 0.085000 ;
      RECT 1625.785000  2.635000 1625.955000 2.805000 ;
      RECT 1626.245000 -0.085000 1626.415000 0.085000 ;
      RECT 1626.245000  2.635000 1626.415000 2.805000 ;
      RECT 1626.305000  1.785000 1626.475000 1.955000 ;
      RECT 1626.705000 -0.085000 1626.875000 0.085000 ;
      RECT 1626.705000  2.635000 1626.875000 2.805000 ;
      RECT 1627.165000 -0.085000 1627.335000 0.085000 ;
      RECT 1627.165000  2.635000 1627.335000 2.805000 ;
      RECT 1627.625000 -0.085000 1627.795000 0.085000 ;
      RECT 1627.625000  2.635000 1627.795000 2.805000 ;
      RECT 1628.085000 -0.085000 1628.255000 0.085000 ;
      RECT 1628.085000  2.635000 1628.255000 2.805000 ;
      RECT 1628.125000  1.785000 1628.295000 1.955000 ;
      RECT 1628.545000 -0.085000 1628.715000 0.085000 ;
      RECT 1628.545000  2.635000 1628.715000 2.805000 ;
      RECT 1628.585000  0.765000 1628.755000 0.935000 ;
      RECT 1629.005000 -0.085000 1629.175000 0.085000 ;
      RECT 1629.005000  2.635000 1629.175000 2.805000 ;
      RECT 1629.465000 -0.085000 1629.635000 0.085000 ;
      RECT 1629.465000  2.635000 1629.635000 2.805000 ;
      RECT 1629.925000 -0.085000 1630.095000 0.085000 ;
      RECT 1629.925000  2.635000 1630.095000 2.805000 ;
      RECT 1630.385000 -0.085000 1630.555000 0.085000 ;
      RECT 1630.385000  2.635000 1630.555000 2.805000 ;
      RECT 1630.845000 -0.085000 1631.015000 0.085000 ;
      RECT 1630.845000  2.635000 1631.015000 2.805000 ;
      RECT 1631.305000 -0.085000 1631.475000 0.085000 ;
      RECT 1631.305000  2.635000 1631.475000 2.805000 ;
      RECT 1631.765000 -0.085000 1631.935000 0.085000 ;
      RECT 1631.765000  2.635000 1631.935000 2.805000 ;
      RECT 1632.225000 -0.085000 1632.395000 0.085000 ;
      RECT 1632.225000  2.635000 1632.395000 2.805000 ;
      RECT 1632.685000 -0.085000 1632.855000 0.085000 ;
      RECT 1632.685000  2.635000 1632.855000 2.805000 ;
      RECT 1633.145000 -0.085000 1633.315000 0.085000 ;
      RECT 1633.145000  2.635000 1633.315000 2.805000 ;
      RECT 1633.605000 -0.085000 1633.775000 0.085000 ;
      RECT 1633.605000  2.635000 1633.775000 2.805000 ;
      RECT 1634.065000 -0.085000 1634.235000 0.085000 ;
      RECT 1634.065000  2.635000 1634.235000 2.805000 ;
      RECT 1634.525000 -0.085000 1634.695000 0.085000 ;
      RECT 1634.525000  2.635000 1634.695000 2.805000 ;
      RECT 1634.985000 -0.085000 1635.155000 0.085000 ;
      RECT 1634.985000  2.635000 1635.155000 2.805000 ;
      RECT 1635.445000 -0.085000 1635.615000 0.085000 ;
      RECT 1635.445000  2.635000 1635.615000 2.805000 ;
      RECT 1635.905000 -0.085000 1636.075000 0.085000 ;
      RECT 1635.905000  2.635000 1636.075000 2.805000 ;
      RECT 1636.365000 -0.085000 1636.535000 0.085000 ;
      RECT 1636.365000  2.635000 1636.535000 2.805000 ;
      RECT 1636.825000 -0.085000 1636.995000 0.085000 ;
      RECT 1636.825000  2.635000 1636.995000 2.805000 ;
      RECT 1637.285000 -0.085000 1637.455000 0.085000 ;
      RECT 1637.285000  2.635000 1637.455000 2.805000 ;
      RECT 1637.745000 -0.085000 1637.915000 0.085000 ;
      RECT 1637.745000  2.635000 1637.915000 2.805000 ;
      RECT 1637.965000  2.125000 1638.135000 2.295000 ;
      RECT 1638.205000 -0.085000 1638.375000 0.085000 ;
      RECT 1638.205000  2.635000 1638.375000 2.805000 ;
      RECT 1638.665000 -0.085000 1638.835000 0.085000 ;
      RECT 1638.665000  2.635000 1638.835000 2.805000 ;
      RECT 1638.985000  2.125000 1639.155000 2.295000 ;
      RECT 1639.125000 -0.085000 1639.295000 0.085000 ;
      RECT 1639.125000  2.635000 1639.295000 2.805000 ;
      RECT 1639.585000 -0.085000 1639.755000 0.085000 ;
      RECT 1639.585000  2.635000 1639.755000 2.805000 ;
      RECT 1640.045000 -0.085000 1640.215000 0.085000 ;
      RECT 1640.045000  2.635000 1640.215000 2.805000 ;
      RECT 1640.505000 -0.085000 1640.675000 0.085000 ;
      RECT 1640.505000  2.635000 1640.675000 2.805000 ;
      RECT 1640.965000 -0.085000 1641.135000 0.085000 ;
      RECT 1640.965000  2.635000 1641.135000 2.805000 ;
      RECT 1641.425000 -0.085000 1641.595000 0.085000 ;
      RECT 1641.425000  2.635000 1641.595000 2.805000 ;
      RECT 1641.885000 -0.085000 1642.055000 0.085000 ;
      RECT 1641.885000  2.635000 1642.055000 2.805000 ;
      RECT 1642.345000 -0.085000 1642.515000 0.085000 ;
      RECT 1642.345000  2.635000 1642.515000 2.805000 ;
      RECT 1642.805000 -0.085000 1642.975000 0.085000 ;
      RECT 1642.805000  2.635000 1642.975000 2.805000 ;
      RECT 1643.265000 -0.085000 1643.435000 0.085000 ;
      RECT 1643.265000  2.635000 1643.435000 2.805000 ;
      RECT 1643.365000  1.445000 1643.535000 1.615000 ;
      RECT 1643.725000 -0.085000 1643.895000 0.085000 ;
      RECT 1643.725000  2.635000 1643.895000 2.805000 ;
      RECT 1644.185000 -0.085000 1644.355000 0.085000 ;
      RECT 1644.185000  2.635000 1644.355000 2.805000 ;
      RECT 1644.645000 -0.085000 1644.815000 0.085000 ;
      RECT 1644.645000  2.635000 1644.815000 2.805000 ;
      RECT 1645.105000 -0.085000 1645.275000 0.085000 ;
      RECT 1645.105000  2.635000 1645.275000 2.805000 ;
      RECT 1645.565000 -0.085000 1645.735000 0.085000 ;
      RECT 1645.565000  2.635000 1645.735000 2.805000 ;
      RECT 1646.025000 -0.085000 1646.195000 0.085000 ;
      RECT 1646.025000  2.635000 1646.195000 2.805000 ;
      RECT 1646.485000 -0.085000 1646.655000 0.085000 ;
      RECT 1646.485000  2.635000 1646.655000 2.805000 ;
      RECT 1646.945000 -0.085000 1647.115000 0.085000 ;
      RECT 1646.945000  2.635000 1647.115000 2.805000 ;
      RECT 1647.405000 -0.085000 1647.575000 0.085000 ;
      RECT 1647.405000  2.635000 1647.575000 2.805000 ;
      RECT 1647.865000 -0.085000 1648.035000 0.085000 ;
      RECT 1647.865000  2.635000 1648.035000 2.805000 ;
      RECT 1648.325000 -0.085000 1648.495000 0.085000 ;
      RECT 1648.325000  2.635000 1648.495000 2.805000 ;
      RECT 1648.785000 -0.085000 1648.955000 0.085000 ;
      RECT 1648.785000  2.635000 1648.955000 2.805000 ;
      RECT 1648.925000  1.445000 1649.095000 1.615000 ;
      RECT 1649.245000 -0.085000 1649.415000 0.085000 ;
      RECT 1649.245000  2.635000 1649.415000 2.805000 ;
      RECT 1649.705000 -0.085000 1649.875000 0.085000 ;
      RECT 1649.705000  2.635000 1649.875000 2.805000 ;
      RECT 1650.165000 -0.085000 1650.335000 0.085000 ;
      RECT 1650.165000  2.635000 1650.335000 2.805000 ;
      RECT 1650.625000 -0.085000 1650.795000 0.085000 ;
      RECT 1650.625000  2.635000 1650.795000 2.805000 ;
      RECT 1651.085000 -0.085000 1651.255000 0.085000 ;
      RECT 1651.085000  2.635000 1651.255000 2.805000 ;
      RECT 1651.545000 -0.085000 1651.715000 0.085000 ;
      RECT 1651.545000  2.635000 1651.715000 2.805000 ;
      RECT 1652.005000 -0.085000 1652.175000 0.085000 ;
      RECT 1652.005000  2.635000 1652.175000 2.805000 ;
      RECT 1652.465000 -0.085000 1652.635000 0.085000 ;
      RECT 1652.465000  2.635000 1652.635000 2.805000 ;
      RECT 1652.925000 -0.085000 1653.095000 0.085000 ;
      RECT 1652.925000  2.635000 1653.095000 2.805000 ;
      RECT 1653.385000 -0.085000 1653.555000 0.085000 ;
      RECT 1653.385000  2.635000 1653.555000 2.805000 ;
      RECT 1653.845000 -0.085000 1654.015000 0.085000 ;
      RECT 1653.845000  2.635000 1654.015000 2.805000 ;
      RECT 1654.305000 -0.085000 1654.475000 0.085000 ;
      RECT 1654.305000  2.635000 1654.475000 2.805000 ;
      RECT 1654.765000 -0.085000 1654.935000 0.085000 ;
      RECT 1654.765000  2.635000 1654.935000 2.805000 ;
      RECT 1655.225000 -0.085000 1655.395000 0.085000 ;
      RECT 1655.225000  2.635000 1655.395000 2.805000 ;
      RECT 1655.685000 -0.085000 1655.855000 0.085000 ;
      RECT 1655.685000  2.635000 1655.855000 2.805000 ;
      RECT 1656.145000 -0.085000 1656.315000 0.085000 ;
      RECT 1656.145000  2.635000 1656.315000 2.805000 ;
      RECT 1656.605000 -0.085000 1656.775000 0.085000 ;
      RECT 1656.605000  2.635000 1656.775000 2.805000 ;
      RECT 1656.805000  1.445000 1656.975000 1.615000 ;
      RECT 1657.065000 -0.085000 1657.235000 0.085000 ;
      RECT 1657.065000  2.635000 1657.235000 2.805000 ;
      RECT 1657.525000 -0.085000 1657.695000 0.085000 ;
      RECT 1657.525000  2.635000 1657.695000 2.805000 ;
      RECT 1657.775000  0.765000 1657.945000 0.935000 ;
      RECT 1657.985000 -0.085000 1658.155000 0.085000 ;
      RECT 1657.985000  2.635000 1658.155000 2.805000 ;
      RECT 1658.285000  0.425000 1658.455000 0.595000 ;
      RECT 1658.445000 -0.085000 1658.615000 0.085000 ;
      RECT 1658.445000  2.635000 1658.615000 2.805000 ;
      RECT 1658.905000 -0.085000 1659.075000 0.085000 ;
      RECT 1658.905000  2.635000 1659.075000 2.805000 ;
      RECT 1659.255000  0.765000 1659.425000 0.935000 ;
      RECT 1659.255000  1.445000 1659.425000 1.615000 ;
      RECT 1659.365000 -0.085000 1659.535000 0.085000 ;
      RECT 1659.365000  2.635000 1659.535000 2.805000 ;
      RECT 1659.825000 -0.085000 1659.995000 0.085000 ;
      RECT 1659.825000  2.635000 1659.995000 2.805000 ;
      RECT 1660.285000 -0.085000 1660.455000 0.085000 ;
      RECT 1660.285000  2.635000 1660.455000 2.805000 ;
      RECT 1660.735000  0.765000 1660.905000 0.935000 ;
      RECT 1660.745000 -0.085000 1660.915000 0.085000 ;
      RECT 1660.745000  2.635000 1660.915000 2.805000 ;
      RECT 1661.205000 -0.085000 1661.375000 0.085000 ;
      RECT 1661.205000  2.635000 1661.375000 2.805000 ;
      RECT 1661.245000  0.425000 1661.415000 0.595000 ;
      RECT 1661.665000 -0.085000 1661.835000 0.085000 ;
      RECT 1661.665000  2.635000 1661.835000 2.805000 ;
      RECT 1662.125000 -0.085000 1662.295000 0.085000 ;
      RECT 1662.125000  2.635000 1662.295000 2.805000 ;
      RECT 1662.585000 -0.085000 1662.755000 0.085000 ;
      RECT 1662.585000  2.635000 1662.755000 2.805000 ;
      RECT 1663.045000 -0.085000 1663.215000 0.085000 ;
      RECT 1663.045000  2.635000 1663.215000 2.805000 ;
      RECT 1663.505000 -0.085000 1663.675000 0.085000 ;
      RECT 1663.505000  2.635000 1663.675000 2.805000 ;
      RECT 1663.965000 -0.085000 1664.135000 0.085000 ;
      RECT 1663.965000  2.635000 1664.135000 2.805000 ;
      RECT 1664.425000 -0.085000 1664.595000 0.085000 ;
      RECT 1664.425000  2.635000 1664.595000 2.805000 ;
      RECT 1664.885000 -0.085000 1665.055000 0.085000 ;
      RECT 1664.885000  2.635000 1665.055000 2.805000 ;
      RECT 1665.345000 -0.085000 1665.515000 0.085000 ;
      RECT 1665.345000  2.635000 1665.515000 2.805000 ;
      RECT 1665.805000 -0.085000 1665.975000 0.085000 ;
      RECT 1665.805000  2.635000 1665.975000 2.805000 ;
      RECT 1666.265000 -0.085000 1666.435000 0.085000 ;
      RECT 1666.265000  2.635000 1666.435000 2.805000 ;
      RECT 1666.725000 -0.085000 1666.895000 0.085000 ;
      RECT 1666.725000  2.635000 1666.895000 2.805000 ;
      RECT 1666.975000  1.445000 1667.145000 1.615000 ;
      RECT 1667.185000 -0.085000 1667.355000 0.085000 ;
      RECT 1667.185000  2.635000 1667.355000 2.805000 ;
      RECT 1667.645000 -0.085000 1667.815000 0.085000 ;
      RECT 1667.645000  2.635000 1667.815000 2.805000 ;
      RECT 1667.945000  0.765000 1668.115000 0.935000 ;
      RECT 1668.105000 -0.085000 1668.275000 0.085000 ;
      RECT 1668.105000  2.635000 1668.275000 2.805000 ;
      RECT 1668.455000  0.425000 1668.625000 0.595000 ;
      RECT 1668.565000 -0.085000 1668.735000 0.085000 ;
      RECT 1668.565000  2.635000 1668.735000 2.805000 ;
      RECT 1669.025000 -0.085000 1669.195000 0.085000 ;
      RECT 1669.025000  2.635000 1669.195000 2.805000 ;
      RECT 1669.425000  0.765000 1669.595000 0.935000 ;
      RECT 1669.425000  1.445000 1669.595000 1.615000 ;
      RECT 1669.485000 -0.085000 1669.655000 0.085000 ;
      RECT 1669.485000  2.635000 1669.655000 2.805000 ;
      RECT 1669.945000 -0.085000 1670.115000 0.085000 ;
      RECT 1669.945000  2.635000 1670.115000 2.805000 ;
      RECT 1670.405000 -0.085000 1670.575000 0.085000 ;
      RECT 1670.405000  2.635000 1670.575000 2.805000 ;
      RECT 1670.865000 -0.085000 1671.035000 0.085000 ;
      RECT 1670.865000  2.635000 1671.035000 2.805000 ;
      RECT 1670.905000  0.765000 1671.075000 0.935000 ;
      RECT 1671.325000 -0.085000 1671.495000 0.085000 ;
      RECT 1671.325000  2.635000 1671.495000 2.805000 ;
      RECT 1671.415000  0.425000 1671.585000 0.595000 ;
      RECT 1671.785000 -0.085000 1671.955000 0.085000 ;
      RECT 1671.785000  2.635000 1671.955000 2.805000 ;
      RECT 1672.245000 -0.085000 1672.415000 0.085000 ;
      RECT 1672.245000  2.635000 1672.415000 2.805000 ;
      RECT 1672.705000 -0.085000 1672.875000 0.085000 ;
      RECT 1672.705000  2.635000 1672.875000 2.805000 ;
      RECT 1673.165000 -0.085000 1673.335000 0.085000 ;
      RECT 1673.165000  2.635000 1673.335000 2.805000 ;
      RECT 1673.625000 -0.085000 1673.795000 0.085000 ;
      RECT 1673.625000  2.635000 1673.795000 2.805000 ;
      RECT 1674.085000 -0.085000 1674.255000 0.085000 ;
      RECT 1674.085000  2.635000 1674.255000 2.805000 ;
      RECT 1674.545000 -0.085000 1674.715000 0.085000 ;
      RECT 1674.545000  2.635000 1674.715000 2.805000 ;
      RECT 1675.005000 -0.085000 1675.175000 0.085000 ;
      RECT 1675.005000  2.635000 1675.175000 2.805000 ;
      RECT 1675.465000 -0.085000 1675.635000 0.085000 ;
      RECT 1675.465000  2.635000 1675.635000 2.805000 ;
      RECT 1675.925000 -0.085000 1676.095000 0.085000 ;
      RECT 1675.925000  2.635000 1676.095000 2.805000 ;
      RECT 1676.385000 -0.085000 1676.555000 0.085000 ;
      RECT 1676.385000  2.635000 1676.555000 2.805000 ;
      RECT 1676.845000 -0.085000 1677.015000 0.085000 ;
      RECT 1676.845000  2.635000 1677.015000 2.805000 ;
      RECT 1677.305000 -0.085000 1677.475000 0.085000 ;
      RECT 1677.305000  2.635000 1677.475000 2.805000 ;
      RECT 1677.765000 -0.085000 1677.935000 0.085000 ;
      RECT 1677.765000  2.635000 1677.935000 2.805000 ;
      RECT 1678.115000  1.445000 1678.285000 1.615000 ;
      RECT 1678.225000 -0.085000 1678.395000 0.085000 ;
      RECT 1678.225000  2.635000 1678.395000 2.805000 ;
      RECT 1678.685000 -0.085000 1678.855000 0.085000 ;
      RECT 1678.685000  2.635000 1678.855000 2.805000 ;
      RECT 1679.085000  0.765000 1679.255000 0.935000 ;
      RECT 1679.145000 -0.085000 1679.315000 0.085000 ;
      RECT 1679.145000  2.635000 1679.315000 2.805000 ;
      RECT 1679.555000  0.425000 1679.725000 0.595000 ;
      RECT 1679.605000 -0.085000 1679.775000 0.085000 ;
      RECT 1679.605000  2.635000 1679.775000 2.805000 ;
      RECT 1680.065000 -0.085000 1680.235000 0.085000 ;
      RECT 1680.065000  2.635000 1680.235000 2.805000 ;
      RECT 1680.525000 -0.085000 1680.695000 0.085000 ;
      RECT 1680.525000  2.635000 1680.695000 2.805000 ;
      RECT 1680.565000  0.765000 1680.735000 0.935000 ;
      RECT 1680.565000  1.445000 1680.735000 1.615000 ;
      RECT 1680.985000 -0.085000 1681.155000 0.085000 ;
      RECT 1680.985000  2.635000 1681.155000 2.805000 ;
      RECT 1681.445000 -0.085000 1681.615000 0.085000 ;
      RECT 1681.445000  2.635000 1681.615000 2.805000 ;
      RECT 1681.905000 -0.085000 1682.075000 0.085000 ;
      RECT 1681.905000  2.635000 1682.075000 2.805000 ;
      RECT 1682.045000  0.765000 1682.215000 0.935000 ;
      RECT 1682.365000 -0.085000 1682.535000 0.085000 ;
      RECT 1682.365000  2.635000 1682.535000 2.805000 ;
      RECT 1682.555000  0.425000 1682.725000 0.595000 ;
      RECT 1682.825000 -0.085000 1682.995000 0.085000 ;
      RECT 1682.825000  2.635000 1682.995000 2.805000 ;
      RECT 1683.285000 -0.085000 1683.455000 0.085000 ;
      RECT 1683.285000  2.635000 1683.455000 2.805000 ;
      RECT 1683.745000 -0.085000 1683.915000 0.085000 ;
      RECT 1683.745000  2.635000 1683.915000 2.805000 ;
      RECT 1684.205000 -0.085000 1684.375000 0.085000 ;
      RECT 1684.205000  2.635000 1684.375000 2.805000 ;
      RECT 1684.665000 -0.085000 1684.835000 0.085000 ;
      RECT 1684.665000  2.635000 1684.835000 2.805000 ;
      RECT 1685.125000 -0.085000 1685.295000 0.085000 ;
      RECT 1685.125000  2.635000 1685.295000 2.805000 ;
      RECT 1685.585000 -0.085000 1685.755000 0.085000 ;
      RECT 1685.585000  2.635000 1685.755000 2.805000 ;
      RECT 1686.045000 -0.085000 1686.215000 0.085000 ;
      RECT 1686.045000  2.635000 1686.215000 2.805000 ;
      RECT 1686.505000 -0.085000 1686.675000 0.085000 ;
      RECT 1686.505000  2.635000 1686.675000 2.805000 ;
      RECT 1686.965000 -0.085000 1687.135000 0.085000 ;
      RECT 1686.965000  2.635000 1687.135000 2.805000 ;
      RECT 1687.425000 -0.085000 1687.595000 0.085000 ;
      RECT 1687.425000  2.635000 1687.595000 2.805000 ;
      RECT 1687.885000 -0.085000 1688.055000 0.085000 ;
      RECT 1687.885000  2.635000 1688.055000 2.805000 ;
      RECT 1688.345000 -0.085000 1688.515000 0.085000 ;
      RECT 1688.345000  2.635000 1688.515000 2.805000 ;
      RECT 1688.805000 -0.085000 1688.975000 0.085000 ;
      RECT 1688.805000  2.635000 1688.975000 2.805000 ;
      RECT 1689.265000 -0.085000 1689.435000 0.085000 ;
      RECT 1689.265000  2.635000 1689.435000 2.805000 ;
      RECT 1689.725000 -0.085000 1689.895000 0.085000 ;
      RECT 1689.725000  2.635000 1689.895000 2.805000 ;
      RECT 1689.825000  1.105000 1689.995000 1.275000 ;
      RECT 1690.185000 -0.085000 1690.355000 0.085000 ;
      RECT 1690.185000  2.635000 1690.355000 2.805000 ;
      RECT 1690.645000 -0.085000 1690.815000 0.085000 ;
      RECT 1690.645000  2.635000 1690.815000 2.805000 ;
      RECT 1691.105000 -0.085000 1691.275000 0.085000 ;
      RECT 1691.105000  2.635000 1691.275000 2.805000 ;
      RECT 1691.565000 -0.085000 1691.735000 0.085000 ;
      RECT 1691.565000  2.635000 1691.735000 2.805000 ;
      RECT 1692.025000 -0.085000 1692.195000 0.085000 ;
      RECT 1692.025000  2.635000 1692.195000 2.805000 ;
      RECT 1692.485000 -0.085000 1692.655000 0.085000 ;
      RECT 1692.485000  1.105000 1692.655000 1.275000 ;
      RECT 1692.485000  2.635000 1692.655000 2.805000 ;
      RECT 1692.945000 -0.085000 1693.115000 0.085000 ;
      RECT 1692.945000  2.635000 1693.115000 2.805000 ;
      RECT 1693.405000 -0.085000 1693.575000 0.085000 ;
      RECT 1693.405000  2.635000 1693.575000 2.805000 ;
      RECT 1693.865000 -0.085000 1694.035000 0.085000 ;
      RECT 1693.865000  2.635000 1694.035000 2.805000 ;
      RECT 1694.325000 -0.085000 1694.495000 0.085000 ;
      RECT 1694.325000  2.635000 1694.495000 2.805000 ;
      RECT 1694.785000 -0.085000 1694.955000 0.085000 ;
      RECT 1694.785000  2.635000 1694.955000 2.805000 ;
      RECT 1695.245000 -0.085000 1695.415000 0.085000 ;
      RECT 1695.245000  2.635000 1695.415000 2.805000 ;
      RECT 1695.705000 -0.085000 1695.875000 0.085000 ;
      RECT 1695.705000  2.635000 1695.875000 2.805000 ;
      RECT 1696.165000 -0.085000 1696.335000 0.085000 ;
      RECT 1696.165000  2.635000 1696.335000 2.805000 ;
      RECT 1696.625000 -0.085000 1696.795000 0.085000 ;
      RECT 1696.625000  2.635000 1696.795000 2.805000 ;
      RECT 1697.085000 -0.085000 1697.255000 0.085000 ;
      RECT 1697.085000  2.635000 1697.255000 2.805000 ;
      RECT 1697.545000 -0.085000 1697.715000 0.085000 ;
      RECT 1697.545000  2.635000 1697.715000 2.805000 ;
      RECT 1697.745000  1.445000 1697.915000 1.615000 ;
      RECT 1698.005000 -0.085000 1698.175000 0.085000 ;
      RECT 1698.005000  2.635000 1698.175000 2.805000 ;
      RECT 1698.465000 -0.085000 1698.635000 0.085000 ;
      RECT 1698.465000  2.635000 1698.635000 2.805000 ;
      RECT 1698.925000 -0.085000 1699.095000 0.085000 ;
      RECT 1698.925000  2.635000 1699.095000 2.805000 ;
      RECT 1699.385000 -0.085000 1699.555000 0.085000 ;
      RECT 1699.385000  2.635000 1699.555000 2.805000 ;
      RECT 1699.845000 -0.085000 1700.015000 0.085000 ;
      RECT 1699.845000  2.635000 1700.015000 2.805000 ;
      RECT 1700.305000 -0.085000 1700.475000 0.085000 ;
      RECT 1700.305000  2.635000 1700.475000 2.805000 ;
      RECT 1700.765000 -0.085000 1700.935000 0.085000 ;
      RECT 1700.765000  2.635000 1700.935000 2.805000 ;
      RECT 1701.225000 -0.085000 1701.395000 0.085000 ;
      RECT 1701.225000  2.635000 1701.395000 2.805000 ;
      RECT 1701.265000  0.725000 1701.435000 0.895000 ;
      RECT 1701.685000 -0.085000 1701.855000 0.085000 ;
      RECT 1701.685000  2.635000 1701.855000 2.805000 ;
      RECT 1702.145000 -0.085000 1702.315000 0.085000 ;
      RECT 1702.145000  2.635000 1702.315000 2.805000 ;
      RECT 1702.605000 -0.085000 1702.775000 0.085000 ;
      RECT 1702.605000  2.635000 1702.775000 2.805000 ;
      RECT 1703.065000 -0.085000 1703.235000 0.085000 ;
      RECT 1703.065000  2.635000 1703.235000 2.805000 ;
      RECT 1703.525000 -0.085000 1703.695000 0.085000 ;
      RECT 1703.525000  2.635000 1703.695000 2.805000 ;
      RECT 1703.865000  1.445000 1704.035000 1.615000 ;
      RECT 1703.985000 -0.085000 1704.155000 0.085000 ;
      RECT 1703.985000  2.635000 1704.155000 2.805000 ;
      RECT 1704.325000  0.725000 1704.495000 0.895000 ;
      RECT 1704.445000 -0.085000 1704.615000 0.085000 ;
      RECT 1704.445000  2.635000 1704.615000 2.805000 ;
      RECT 1704.905000 -0.085000 1705.075000 0.085000 ;
      RECT 1704.905000  2.635000 1705.075000 2.805000 ;
      RECT 1705.365000 -0.085000 1705.535000 0.085000 ;
      RECT 1705.365000  2.635000 1705.535000 2.805000 ;
      RECT 1705.825000 -0.085000 1705.995000 0.085000 ;
      RECT 1705.825000  2.635000 1705.995000 2.805000 ;
      RECT 1706.285000 -0.085000 1706.455000 0.085000 ;
      RECT 1706.285000  2.635000 1706.455000 2.805000 ;
      RECT 1706.745000 -0.085000 1706.915000 0.085000 ;
      RECT 1706.745000  2.635000 1706.915000 2.805000 ;
      RECT 1707.205000 -0.085000 1707.375000 0.085000 ;
      RECT 1707.205000  2.635000 1707.375000 2.805000 ;
      RECT 1707.665000 -0.085000 1707.835000 0.085000 ;
      RECT 1707.665000  2.635000 1707.835000 2.805000 ;
      RECT 1708.125000 -0.085000 1708.295000 0.085000 ;
      RECT 1708.125000  2.635000 1708.295000 2.805000 ;
      RECT 1708.585000 -0.085000 1708.755000 0.085000 ;
      RECT 1708.585000  2.635000 1708.755000 2.805000 ;
      RECT 1709.045000 -0.085000 1709.215000 0.085000 ;
      RECT 1709.045000  2.635000 1709.215000 2.805000 ;
      RECT 1709.505000 -0.085000 1709.675000 0.085000 ;
      RECT 1709.505000  2.635000 1709.675000 2.805000 ;
      RECT 1709.965000 -0.085000 1710.135000 0.085000 ;
      RECT 1709.965000  2.635000 1710.135000 2.805000 ;
      RECT 1710.425000 -0.085000 1710.595000 0.085000 ;
      RECT 1710.425000  2.635000 1710.595000 2.805000 ;
      RECT 1710.625000  1.445000 1710.795000 1.615000 ;
      RECT 1710.885000 -0.085000 1711.055000 0.085000 ;
      RECT 1710.885000  2.635000 1711.055000 2.805000 ;
      RECT 1711.345000 -0.085000 1711.515000 0.085000 ;
      RECT 1711.345000  2.635000 1711.515000 2.805000 ;
      RECT 1711.595000  0.765000 1711.765000 0.935000 ;
      RECT 1711.805000 -0.085000 1711.975000 0.085000 ;
      RECT 1711.805000  2.635000 1711.975000 2.805000 ;
      RECT 1712.105000  0.425000 1712.275000 0.595000 ;
      RECT 1712.265000 -0.085000 1712.435000 0.085000 ;
      RECT 1712.265000  2.635000 1712.435000 2.805000 ;
      RECT 1712.725000 -0.085000 1712.895000 0.085000 ;
      RECT 1712.725000  2.635000 1712.895000 2.805000 ;
      RECT 1713.075000  0.765000 1713.245000 0.935000 ;
      RECT 1713.075000  1.445000 1713.245000 1.615000 ;
      RECT 1713.185000 -0.085000 1713.355000 0.085000 ;
      RECT 1713.185000  2.635000 1713.355000 2.805000 ;
      RECT 1713.645000 -0.085000 1713.815000 0.085000 ;
      RECT 1713.645000  2.635000 1713.815000 2.805000 ;
      RECT 1714.105000 -0.085000 1714.275000 0.085000 ;
      RECT 1714.105000  2.635000 1714.275000 2.805000 ;
      RECT 1714.555000  0.765000 1714.725000 0.935000 ;
      RECT 1714.565000 -0.085000 1714.735000 0.085000 ;
      RECT 1714.565000  2.635000 1714.735000 2.805000 ;
      RECT 1715.025000 -0.085000 1715.195000 0.085000 ;
      RECT 1715.025000  2.635000 1715.195000 2.805000 ;
      RECT 1715.065000  0.425000 1715.235000 0.595000 ;
      RECT 1715.485000 -0.085000 1715.655000 0.085000 ;
      RECT 1715.485000  2.635000 1715.655000 2.805000 ;
      RECT 1715.945000 -0.085000 1716.115000 0.085000 ;
      RECT 1715.945000  2.635000 1716.115000 2.805000 ;
      RECT 1716.405000 -0.085000 1716.575000 0.085000 ;
      RECT 1716.405000  2.635000 1716.575000 2.805000 ;
      RECT 1716.865000 -0.085000 1717.035000 0.085000 ;
      RECT 1716.865000  2.635000 1717.035000 2.805000 ;
      RECT 1717.325000 -0.085000 1717.495000 0.085000 ;
      RECT 1717.325000  2.635000 1717.495000 2.805000 ;
      RECT 1717.785000 -0.085000 1717.955000 0.085000 ;
      RECT 1717.785000  2.635000 1717.955000 2.805000 ;
      RECT 1718.245000 -0.085000 1718.415000 0.085000 ;
      RECT 1718.245000  2.635000 1718.415000 2.805000 ;
      RECT 1718.705000 -0.085000 1718.875000 0.085000 ;
      RECT 1718.705000  2.635000 1718.875000 2.805000 ;
      RECT 1719.165000 -0.085000 1719.335000 0.085000 ;
      RECT 1719.165000  2.635000 1719.335000 2.805000 ;
      RECT 1719.625000 -0.085000 1719.795000 0.085000 ;
      RECT 1719.625000  2.635000 1719.795000 2.805000 ;
      RECT 1720.085000 -0.085000 1720.255000 0.085000 ;
      RECT 1720.085000  2.635000 1720.255000 2.805000 ;
      RECT 1720.545000 -0.085000 1720.715000 0.085000 ;
      RECT 1720.545000  2.635000 1720.715000 2.805000 ;
      RECT 1721.005000 -0.085000 1721.175000 0.085000 ;
      RECT 1721.005000  2.635000 1721.175000 2.805000 ;
      RECT 1721.040000  1.445000 1721.210000 1.615000 ;
      RECT 1721.465000 -0.085000 1721.635000 0.085000 ;
      RECT 1721.465000  2.635000 1721.635000 2.805000 ;
      RECT 1721.925000 -0.085000 1722.095000 0.085000 ;
      RECT 1721.925000  2.635000 1722.095000 2.805000 ;
      RECT 1722.010000  0.765000 1722.180000 0.935000 ;
      RECT 1722.385000 -0.085000 1722.555000 0.085000 ;
      RECT 1722.385000  2.635000 1722.555000 2.805000 ;
      RECT 1722.520000  0.425000 1722.690000 0.595000 ;
      RECT 1722.845000 -0.085000 1723.015000 0.085000 ;
      RECT 1722.845000  2.635000 1723.015000 2.805000 ;
      RECT 1723.305000 -0.085000 1723.475000 0.085000 ;
      RECT 1723.305000  2.635000 1723.475000 2.805000 ;
      RECT 1723.490000  0.765000 1723.660000 0.935000 ;
      RECT 1723.490000  1.445000 1723.660000 1.615000 ;
      RECT 1723.765000 -0.085000 1723.935000 0.085000 ;
      RECT 1723.765000  2.635000 1723.935000 2.805000 ;
      RECT 1724.225000 -0.085000 1724.395000 0.085000 ;
      RECT 1724.225000  2.635000 1724.395000 2.805000 ;
      RECT 1724.685000 -0.085000 1724.855000 0.085000 ;
      RECT 1724.685000  2.635000 1724.855000 2.805000 ;
      RECT 1724.970000  0.765000 1725.140000 0.935000 ;
      RECT 1725.145000 -0.085000 1725.315000 0.085000 ;
      RECT 1725.145000  2.635000 1725.315000 2.805000 ;
      RECT 1725.480000  0.425000 1725.650000 0.595000 ;
      RECT 1725.605000 -0.085000 1725.775000 0.085000 ;
      RECT 1725.605000  2.635000 1725.775000 2.805000 ;
      RECT 1726.065000 -0.085000 1726.235000 0.085000 ;
      RECT 1726.065000  2.635000 1726.235000 2.805000 ;
      RECT 1726.525000 -0.085000 1726.695000 0.085000 ;
      RECT 1726.525000  2.635000 1726.695000 2.805000 ;
      RECT 1726.985000 -0.085000 1727.155000 0.085000 ;
      RECT 1726.985000  2.635000 1727.155000 2.805000 ;
      RECT 1727.445000 -0.085000 1727.615000 0.085000 ;
      RECT 1727.445000  2.635000 1727.615000 2.805000 ;
      RECT 1727.905000 -0.085000 1728.075000 0.085000 ;
      RECT 1727.905000  2.635000 1728.075000 2.805000 ;
      RECT 1728.365000 -0.085000 1728.535000 0.085000 ;
      RECT 1728.365000  2.635000 1728.535000 2.805000 ;
      RECT 1728.825000 -0.085000 1728.995000 0.085000 ;
      RECT 1728.825000  2.635000 1728.995000 2.805000 ;
      RECT 1729.285000 -0.085000 1729.455000 0.085000 ;
      RECT 1729.285000  2.635000 1729.455000 2.805000 ;
      RECT 1729.745000 -0.085000 1729.915000 0.085000 ;
      RECT 1729.745000  2.635000 1729.915000 2.805000 ;
      RECT 1730.205000 -0.085000 1730.375000 0.085000 ;
      RECT 1730.205000  2.635000 1730.375000 2.805000 ;
      RECT 1730.665000 -0.085000 1730.835000 0.085000 ;
      RECT 1730.665000  2.635000 1730.835000 2.805000 ;
      RECT 1731.125000 -0.085000 1731.295000 0.085000 ;
      RECT 1731.125000  2.635000 1731.295000 2.805000 ;
      RECT 1731.585000 -0.085000 1731.755000 0.085000 ;
      RECT 1731.585000  2.635000 1731.755000 2.805000 ;
      RECT 1732.035000  1.445000 1732.205000 1.615000 ;
      RECT 1732.045000 -0.085000 1732.215000 0.085000 ;
      RECT 1732.045000  2.635000 1732.215000 2.805000 ;
      RECT 1732.505000 -0.085000 1732.675000 0.085000 ;
      RECT 1732.505000  2.635000 1732.675000 2.805000 ;
      RECT 1732.965000 -0.085000 1733.135000 0.085000 ;
      RECT 1732.965000  2.635000 1733.135000 2.805000 ;
      RECT 1733.005000  0.765000 1733.175000 0.935000 ;
      RECT 1733.425000 -0.085000 1733.595000 0.085000 ;
      RECT 1733.425000  2.635000 1733.595000 2.805000 ;
      RECT 1733.515000  0.425000 1733.685000 0.595000 ;
      RECT 1733.885000 -0.085000 1734.055000 0.085000 ;
      RECT 1733.885000  2.635000 1734.055000 2.805000 ;
      RECT 1734.345000 -0.085000 1734.515000 0.085000 ;
      RECT 1734.345000  2.635000 1734.515000 2.805000 ;
      RECT 1734.485000  0.765000 1734.655000 0.935000 ;
      RECT 1734.485000  1.445000 1734.655000 1.615000 ;
      RECT 1734.805000 -0.085000 1734.975000 0.085000 ;
      RECT 1734.805000  2.635000 1734.975000 2.805000 ;
      RECT 1735.265000 -0.085000 1735.435000 0.085000 ;
      RECT 1735.265000  2.635000 1735.435000 2.805000 ;
      RECT 1735.725000 -0.085000 1735.895000 0.085000 ;
      RECT 1735.725000  2.635000 1735.895000 2.805000 ;
      RECT 1735.965000  0.765000 1736.135000 0.935000 ;
      RECT 1736.185000 -0.085000 1736.355000 0.085000 ;
      RECT 1736.185000  2.635000 1736.355000 2.805000 ;
      RECT 1736.475000  0.425000 1736.645000 0.595000 ;
      RECT 1736.645000 -0.085000 1736.815000 0.085000 ;
      RECT 1736.645000  2.635000 1736.815000 2.805000 ;
      RECT 1737.105000 -0.085000 1737.275000 0.085000 ;
      RECT 1737.105000  2.635000 1737.275000 2.805000 ;
      RECT 1737.565000 -0.085000 1737.735000 0.085000 ;
      RECT 1737.565000  2.635000 1737.735000 2.805000 ;
      RECT 1738.025000 -0.085000 1738.195000 0.085000 ;
      RECT 1738.025000  2.635000 1738.195000 2.805000 ;
      RECT 1738.485000 -0.085000 1738.655000 0.085000 ;
      RECT 1738.485000  2.635000 1738.655000 2.805000 ;
      RECT 1738.945000 -0.085000 1739.115000 0.085000 ;
      RECT 1738.945000  2.635000 1739.115000 2.805000 ;
      RECT 1739.195000  1.105000 1739.365000 1.275000 ;
      RECT 1739.405000 -0.085000 1739.575000 0.085000 ;
      RECT 1739.405000  2.635000 1739.575000 2.805000 ;
      RECT 1739.475000  1.785000 1739.645000 1.955000 ;
      RECT 1739.865000 -0.085000 1740.035000 0.085000 ;
      RECT 1739.865000  2.635000 1740.035000 2.805000 ;
      RECT 1740.325000 -0.085000 1740.495000 0.085000 ;
      RECT 1740.325000  2.635000 1740.495000 2.805000 ;
      RECT 1740.785000 -0.085000 1740.955000 0.085000 ;
      RECT 1740.785000  2.635000 1740.955000 2.805000 ;
      RECT 1741.245000 -0.085000 1741.415000 0.085000 ;
      RECT 1741.245000  2.635000 1741.415000 2.805000 ;
      RECT 1741.705000 -0.085000 1741.875000 0.085000 ;
      RECT 1741.705000  2.635000 1741.875000 2.805000 ;
      RECT 1742.165000 -0.085000 1742.335000 0.085000 ;
      RECT 1742.165000  2.635000 1742.335000 2.805000 ;
      RECT 1742.625000 -0.085000 1742.795000 0.085000 ;
      RECT 1742.625000  2.635000 1742.795000 2.805000 ;
      RECT 1743.085000 -0.085000 1743.255000 0.085000 ;
      RECT 1743.085000  2.635000 1743.255000 2.805000 ;
      RECT 1743.545000 -0.085000 1743.715000 0.085000 ;
      RECT 1743.545000  2.635000 1743.715000 2.805000 ;
      RECT 1743.820000  1.105000 1743.990000 1.275000 ;
      RECT 1744.005000 -0.085000 1744.175000 0.085000 ;
      RECT 1744.005000  2.635000 1744.175000 2.805000 ;
      RECT 1744.290000  1.785000 1744.460000 1.955000 ;
      RECT 1744.465000 -0.085000 1744.635000 0.085000 ;
      RECT 1744.465000  2.635000 1744.635000 2.805000 ;
      RECT 1744.925000 -0.085000 1745.095000 0.085000 ;
      RECT 1744.925000  2.635000 1745.095000 2.805000 ;
      RECT 1745.385000 -0.085000 1745.555000 0.085000 ;
      RECT 1745.385000  2.635000 1745.555000 2.805000 ;
      RECT 1745.595000  0.765000 1745.765000 0.935000 ;
      RECT 1745.845000 -0.085000 1746.015000 0.085000 ;
      RECT 1745.845000  2.635000 1746.015000 2.805000 ;
      RECT 1745.955000  0.765000 1746.125000 0.935000 ;
      RECT 1746.305000 -0.085000 1746.475000 0.085000 ;
      RECT 1746.305000  2.635000 1746.475000 2.805000 ;
      RECT 1746.765000 -0.085000 1746.935000 0.085000 ;
      RECT 1746.765000  2.635000 1746.935000 2.805000 ;
      RECT 1747.225000 -0.085000 1747.395000 0.085000 ;
      RECT 1747.225000  2.635000 1747.395000 2.805000 ;
      RECT 1747.575000  1.105000 1747.745000 1.275000 ;
      RECT 1747.685000 -0.085000 1747.855000 0.085000 ;
      RECT 1747.685000  2.635000 1747.855000 2.805000 ;
      RECT 1747.905000  1.785000 1748.075000 1.955000 ;
      RECT 1748.145000 -0.085000 1748.315000 0.085000 ;
      RECT 1748.145000  2.635000 1748.315000 2.805000 ;
      RECT 1748.605000 -0.085000 1748.775000 0.085000 ;
      RECT 1748.605000  2.635000 1748.775000 2.805000 ;
      RECT 1749.065000 -0.085000 1749.235000 0.085000 ;
      RECT 1749.065000  2.635000 1749.235000 2.805000 ;
      RECT 1749.175000  1.085000 1749.345000 1.255000 ;
      RECT 1749.515000  0.765000 1749.685000 0.935000 ;
      RECT 1749.525000 -0.085000 1749.695000 0.085000 ;
      RECT 1749.525000  2.635000 1749.695000 2.805000 ;
      RECT 1749.985000 -0.085000 1750.155000 0.085000 ;
      RECT 1749.985000  2.635000 1750.155000 2.805000 ;
      RECT 1750.445000 -0.085000 1750.615000 0.085000 ;
      RECT 1750.445000  2.635000 1750.615000 2.805000 ;
      RECT 1750.905000 -0.085000 1751.075000 0.085000 ;
      RECT 1750.905000  2.635000 1751.075000 2.805000 ;
      RECT 1751.365000 -0.085000 1751.535000 0.085000 ;
      RECT 1751.365000  2.635000 1751.535000 2.805000 ;
      RECT 1751.825000 -0.085000 1751.995000 0.085000 ;
      RECT 1751.825000  2.635000 1751.995000 2.805000 ;
      RECT 1752.285000 -0.085000 1752.455000 0.085000 ;
      RECT 1752.285000  2.635000 1752.455000 2.805000 ;
      RECT 1752.745000 -0.085000 1752.915000 0.085000 ;
      RECT 1752.745000  2.635000 1752.915000 2.805000 ;
      RECT 1753.205000 -0.085000 1753.375000 0.085000 ;
      RECT 1753.205000  2.635000 1753.375000 2.805000 ;
      RECT 1753.665000 -0.085000 1753.835000 0.085000 ;
      RECT 1753.665000  2.635000 1753.835000 2.805000 ;
      RECT 1754.125000 -0.085000 1754.295000 0.085000 ;
      RECT 1754.125000  2.635000 1754.295000 2.805000 ;
      RECT 1754.585000 -0.085000 1754.755000 0.085000 ;
      RECT 1754.585000  2.635000 1754.755000 2.805000 ;
      RECT 1755.045000 -0.085000 1755.215000 0.085000 ;
      RECT 1755.045000  2.635000 1755.215000 2.805000 ;
      RECT 1755.505000 -0.085000 1755.675000 0.085000 ;
      RECT 1755.505000  2.635000 1755.675000 2.805000 ;
      RECT 1755.965000 -0.085000 1756.135000 0.085000 ;
      RECT 1755.965000  2.635000 1756.135000 2.805000 ;
      RECT 1756.425000 -0.085000 1756.595000 0.085000 ;
      RECT 1756.425000  2.635000 1756.595000 2.805000 ;
      RECT 1756.885000 -0.085000 1757.055000 0.085000 ;
      RECT 1756.885000  2.635000 1757.055000 2.805000 ;
      RECT 1757.345000 -0.085000 1757.515000 0.085000 ;
      RECT 1757.345000  2.635000 1757.515000 2.805000 ;
      RECT 1757.805000 -0.085000 1757.975000 0.085000 ;
      RECT 1757.805000  2.635000 1757.975000 2.805000 ;
      RECT 1758.265000 -0.085000 1758.435000 0.085000 ;
      RECT 1758.265000  2.635000 1758.435000 2.805000 ;
      RECT 1758.725000 -0.085000 1758.895000 0.085000 ;
      RECT 1758.725000  2.635000 1758.895000 2.805000 ;
      RECT 1759.185000 -0.085000 1759.355000 0.085000 ;
      RECT 1759.185000  2.635000 1759.355000 2.805000 ;
      RECT 1759.645000 -0.085000 1759.815000 0.085000 ;
      RECT 1759.645000  2.635000 1759.815000 2.805000 ;
      RECT 1760.105000 -0.085000 1760.275000 0.085000 ;
      RECT 1760.105000  2.635000 1760.275000 2.805000 ;
      RECT 1760.565000 -0.085000 1760.735000 0.085000 ;
      RECT 1760.565000  2.635000 1760.735000 2.805000 ;
      RECT 1761.025000 -0.085000 1761.195000 0.085000 ;
      RECT 1761.025000  2.635000 1761.195000 2.805000 ;
      RECT 1761.485000 -0.085000 1761.655000 0.085000 ;
      RECT 1761.485000  2.635000 1761.655000 2.805000 ;
      RECT 1761.945000 -0.085000 1762.115000 0.085000 ;
      RECT 1761.945000  2.635000 1762.115000 2.805000 ;
      RECT 1762.405000 -0.085000 1762.575000 0.085000 ;
      RECT 1762.405000  2.635000 1762.575000 2.805000 ;
      RECT 1762.865000 -0.085000 1763.035000 0.085000 ;
      RECT 1762.865000  2.635000 1763.035000 2.805000 ;
      RECT 1763.325000 -0.085000 1763.495000 0.085000 ;
      RECT 1763.325000  2.635000 1763.495000 2.805000 ;
      RECT 1763.785000 -0.085000 1763.955000 0.085000 ;
      RECT 1763.785000  2.635000 1763.955000 2.805000 ;
      RECT 1764.245000 -0.085000 1764.415000 0.085000 ;
      RECT 1764.245000  2.635000 1764.415000 2.805000 ;
      RECT 1764.705000 -0.085000 1764.875000 0.085000 ;
      RECT 1764.705000  2.635000 1764.875000 2.805000 ;
      RECT 1765.165000 -0.085000 1765.335000 0.085000 ;
      RECT 1765.165000  2.635000 1765.335000 2.805000 ;
      RECT 1765.625000 -0.085000 1765.795000 0.085000 ;
      RECT 1765.625000  2.635000 1765.795000 2.805000 ;
      RECT 1766.085000 -0.085000 1766.255000 0.085000 ;
      RECT 1766.085000  2.635000 1766.255000 2.805000 ;
      RECT 1766.545000 -0.085000 1766.715000 0.085000 ;
      RECT 1766.545000  2.635000 1766.715000 2.805000 ;
      RECT 1767.005000 -0.085000 1767.175000 0.085000 ;
      RECT 1767.005000  2.635000 1767.175000 2.805000 ;
      RECT 1767.465000 -0.085000 1767.635000 0.085000 ;
      RECT 1767.465000  2.635000 1767.635000 2.805000 ;
      RECT 1767.925000 -0.085000 1768.095000 0.085000 ;
      RECT 1767.925000  2.635000 1768.095000 2.805000 ;
      RECT 1768.385000 -0.085000 1768.555000 0.085000 ;
      RECT 1768.385000  2.635000 1768.555000 2.805000 ;
      RECT 1768.845000 -0.085000 1769.015000 0.085000 ;
      RECT 1768.845000  2.635000 1769.015000 2.805000 ;
      RECT 1769.305000 -0.085000 1769.475000 0.085000 ;
      RECT 1769.305000  2.635000 1769.475000 2.805000 ;
      RECT 1769.765000 -0.085000 1769.935000 0.085000 ;
      RECT 1769.765000  2.635000 1769.935000 2.805000 ;
      RECT 1770.225000 -0.085000 1770.395000 0.085000 ;
      RECT 1770.225000  2.635000 1770.395000 2.805000 ;
      RECT 1770.685000 -0.085000 1770.855000 0.085000 ;
      RECT 1770.685000  2.635000 1770.855000 2.805000 ;
      RECT 1771.145000 -0.085000 1771.315000 0.085000 ;
      RECT 1771.145000  2.635000 1771.315000 2.805000 ;
      RECT 1771.605000 -0.085000 1771.775000 0.085000 ;
      RECT 1771.605000  2.635000 1771.775000 2.805000 ;
      RECT 1772.065000 -0.085000 1772.235000 0.085000 ;
      RECT 1772.065000  2.635000 1772.235000 2.805000 ;
      RECT 1772.525000 -0.085000 1772.695000 0.085000 ;
      RECT 1772.525000  2.635000 1772.695000 2.805000 ;
      RECT 1772.985000 -0.085000 1773.155000 0.085000 ;
      RECT 1772.985000  2.635000 1773.155000 2.805000 ;
      RECT 1773.445000 -0.085000 1773.615000 0.085000 ;
      RECT 1773.445000  2.635000 1773.615000 2.805000 ;
      RECT 1773.905000 -0.085000 1774.075000 0.085000 ;
      RECT 1773.905000  2.635000 1774.075000 2.805000 ;
      RECT 1774.365000 -0.085000 1774.535000 0.085000 ;
      RECT 1774.365000  2.635000 1774.535000 2.805000 ;
      RECT 1774.825000 -0.085000 1774.995000 0.085000 ;
      RECT 1774.825000  2.635000 1774.995000 2.805000 ;
      RECT 1775.285000 -0.085000 1775.455000 0.085000 ;
      RECT 1775.285000  2.635000 1775.455000 2.805000 ;
      RECT 1775.745000 -0.085000 1775.915000 0.085000 ;
      RECT 1775.745000  2.635000 1775.915000 2.805000 ;
      RECT 1776.205000 -0.085000 1776.375000 0.085000 ;
      RECT 1776.205000  2.635000 1776.375000 2.805000 ;
      RECT 1776.665000 -0.085000 1776.835000 0.085000 ;
      RECT 1776.665000  2.635000 1776.835000 2.805000 ;
      RECT 1777.125000 -0.085000 1777.295000 0.085000 ;
      RECT 1777.125000  2.635000 1777.295000 2.805000 ;
      RECT 1777.585000 -0.085000 1777.755000 0.085000 ;
      RECT 1777.585000  2.635000 1777.755000 2.805000 ;
      RECT 1778.045000 -0.085000 1778.215000 0.085000 ;
      RECT 1778.045000  2.635000 1778.215000 2.805000 ;
      RECT 1778.505000 -0.085000 1778.675000 0.085000 ;
      RECT 1778.505000  2.635000 1778.675000 2.805000 ;
      RECT 1778.965000 -0.085000 1779.135000 0.085000 ;
      RECT 1778.965000  2.635000 1779.135000 2.805000 ;
      RECT 1779.425000 -0.085000 1779.595000 0.085000 ;
      RECT 1779.425000  2.635000 1779.595000 2.805000 ;
      RECT 1779.885000 -0.085000 1780.055000 0.085000 ;
      RECT 1779.885000  2.635000 1780.055000 2.805000 ;
      RECT 1780.345000 -0.085000 1780.515000 0.085000 ;
      RECT 1780.345000  2.635000 1780.515000 2.805000 ;
      RECT 1780.805000 -0.085000 1780.975000 0.085000 ;
      RECT 1780.805000  2.635000 1780.975000 2.805000 ;
      RECT 1781.265000 -0.085000 1781.435000 0.085000 ;
      RECT 1781.265000  2.635000 1781.435000 2.805000 ;
      RECT 1781.725000 -0.085000 1781.895000 0.085000 ;
      RECT 1781.725000  2.635000 1781.895000 2.805000 ;
      RECT 1782.185000 -0.085000 1782.355000 0.085000 ;
      RECT 1782.185000  2.635000 1782.355000 2.805000 ;
      RECT 1782.645000 -0.085000 1782.815000 0.085000 ;
      RECT 1782.645000  2.635000 1782.815000 2.805000 ;
      RECT 1783.105000 -0.085000 1783.275000 0.085000 ;
      RECT 1783.105000  2.635000 1783.275000 2.805000 ;
      RECT 1783.565000 -0.085000 1783.735000 0.085000 ;
      RECT 1783.565000  2.635000 1783.735000 2.805000 ;
      RECT 1784.025000 -0.085000 1784.195000 0.085000 ;
      RECT 1784.025000  2.635000 1784.195000 2.805000 ;
      RECT 1784.485000 -0.085000 1784.655000 0.085000 ;
      RECT 1784.485000  2.635000 1784.655000 2.805000 ;
      RECT 1784.945000 -0.085000 1785.115000 0.085000 ;
      RECT 1784.945000  2.635000 1785.115000 2.805000 ;
      RECT 1785.405000 -0.085000 1785.575000 0.085000 ;
      RECT 1785.405000  2.635000 1785.575000 2.805000 ;
      RECT 1785.865000 -0.085000 1786.035000 0.085000 ;
      RECT 1785.865000  2.635000 1786.035000 2.805000 ;
      RECT 1786.325000 -0.085000 1786.495000 0.085000 ;
      RECT 1786.325000  2.635000 1786.495000 2.805000 ;
      RECT 1786.785000 -0.085000 1786.955000 0.085000 ;
      RECT 1786.785000  2.635000 1786.955000 2.805000 ;
      RECT 1787.245000 -0.085000 1787.415000 0.085000 ;
      RECT 1787.245000  2.635000 1787.415000 2.805000 ;
      RECT 1787.705000 -0.085000 1787.875000 0.085000 ;
      RECT 1787.705000  2.635000 1787.875000 2.805000 ;
      RECT 1788.165000 -0.085000 1788.335000 0.085000 ;
      RECT 1788.165000  2.635000 1788.335000 2.805000 ;
      RECT 1788.625000 -0.085000 1788.795000 0.085000 ;
      RECT 1788.625000  2.635000 1788.795000 2.805000 ;
      RECT 1789.085000 -0.085000 1789.255000 0.085000 ;
      RECT 1789.085000  2.635000 1789.255000 2.805000 ;
      RECT 1789.545000 -0.085000 1789.715000 0.085000 ;
      RECT 1789.545000  2.635000 1789.715000 2.805000 ;
      RECT 1790.005000 -0.085000 1790.175000 0.085000 ;
      RECT 1790.005000  2.635000 1790.175000 2.805000 ;
      RECT 1790.465000 -0.085000 1790.635000 0.085000 ;
      RECT 1790.465000  2.635000 1790.635000 2.805000 ;
      RECT 1790.925000 -0.085000 1791.095000 0.085000 ;
      RECT 1790.925000  2.635000 1791.095000 2.805000 ;
      RECT 1791.385000 -0.085000 1791.555000 0.085000 ;
      RECT 1791.385000  2.635000 1791.555000 2.805000 ;
      RECT 1791.845000 -0.085000 1792.015000 0.085000 ;
      RECT 1791.845000  2.635000 1792.015000 2.805000 ;
      RECT 1792.305000 -0.085000 1792.475000 0.085000 ;
      RECT 1792.305000  2.635000 1792.475000 2.805000 ;
      RECT 1792.765000 -0.085000 1792.935000 0.085000 ;
      RECT 1792.765000  2.635000 1792.935000 2.805000 ;
      RECT 1793.225000 -0.085000 1793.395000 0.085000 ;
      RECT 1793.225000  2.635000 1793.395000 2.805000 ;
      RECT 1793.685000 -0.085000 1793.855000 0.085000 ;
      RECT 1793.685000  2.635000 1793.855000 2.805000 ;
      RECT 1794.145000 -0.085000 1794.315000 0.085000 ;
      RECT 1794.145000  2.635000 1794.315000 2.805000 ;
      RECT 1794.605000 -0.085000 1794.775000 0.085000 ;
      RECT 1794.605000  2.635000 1794.775000 2.805000 ;
      RECT 1795.065000 -0.085000 1795.235000 0.085000 ;
      RECT 1795.065000  2.635000 1795.235000 2.805000 ;
      RECT 1795.525000 -0.085000 1795.695000 0.085000 ;
      RECT 1795.525000  2.635000 1795.695000 2.805000 ;
      RECT 1795.985000 -0.085000 1796.155000 0.085000 ;
      RECT 1795.985000  2.635000 1796.155000 2.805000 ;
      RECT 1796.445000 -0.085000 1796.615000 0.085000 ;
      RECT 1796.445000  2.635000 1796.615000 2.805000 ;
      RECT 1796.905000 -0.085000 1797.075000 0.085000 ;
      RECT 1796.905000  2.635000 1797.075000 2.805000 ;
      RECT 1797.365000 -0.085000 1797.535000 0.085000 ;
      RECT 1797.365000  2.635000 1797.535000 2.805000 ;
      RECT 1797.825000 -0.085000 1797.995000 0.085000 ;
      RECT 1797.825000  2.635000 1797.995000 2.805000 ;
      RECT 1798.285000 -0.085000 1798.455000 0.085000 ;
      RECT 1798.285000  2.635000 1798.455000 2.805000 ;
      RECT 1798.745000 -0.085000 1798.915000 0.085000 ;
      RECT 1798.745000  2.635000 1798.915000 2.805000 ;
      RECT 1799.205000 -0.085000 1799.375000 0.085000 ;
      RECT 1799.205000  2.635000 1799.375000 2.805000 ;
      RECT 1799.665000 -0.085000 1799.835000 0.085000 ;
      RECT 1799.665000  2.635000 1799.835000 2.805000 ;
      RECT 1800.125000 -0.085000 1800.295000 0.085000 ;
      RECT 1800.125000  2.635000 1800.295000 2.805000 ;
      RECT 1800.585000 -0.085000 1800.755000 0.085000 ;
      RECT 1800.585000  2.635000 1800.755000 2.805000 ;
      RECT 1801.045000 -0.085000 1801.215000 0.085000 ;
      RECT 1801.045000  2.635000 1801.215000 2.805000 ;
      RECT 1801.505000 -0.085000 1801.675000 0.085000 ;
      RECT 1801.505000  2.635000 1801.675000 2.805000 ;
      RECT 1801.965000 -0.085000 1802.135000 0.085000 ;
      RECT 1801.965000  2.635000 1802.135000 2.805000 ;
      RECT 1802.425000 -0.085000 1802.595000 0.085000 ;
      RECT 1802.425000  2.635000 1802.595000 2.805000 ;
      RECT 1802.885000 -0.085000 1803.055000 0.085000 ;
      RECT 1802.885000  2.635000 1803.055000 2.805000 ;
      RECT 1803.345000 -0.085000 1803.515000 0.085000 ;
      RECT 1803.345000  2.635000 1803.515000 2.805000 ;
      RECT 1803.805000 -0.085000 1803.975000 0.085000 ;
      RECT 1803.805000  2.635000 1803.975000 2.805000 ;
      RECT 1804.265000 -0.085000 1804.435000 0.085000 ;
      RECT 1804.265000  2.635000 1804.435000 2.805000 ;
      RECT 1804.725000 -0.085000 1804.895000 0.085000 ;
      RECT 1804.725000  2.635000 1804.895000 2.805000 ;
      RECT 1805.185000 -0.085000 1805.355000 0.085000 ;
      RECT 1805.185000  2.635000 1805.355000 2.805000 ;
      RECT 1805.645000 -0.085000 1805.815000 0.085000 ;
      RECT 1805.645000  2.635000 1805.815000 2.805000 ;
      RECT 1806.105000 -0.085000 1806.275000 0.085000 ;
      RECT 1806.105000  2.635000 1806.275000 2.805000 ;
      RECT 1806.565000 -0.085000 1806.735000 0.085000 ;
      RECT 1806.565000  2.635000 1806.735000 2.805000 ;
      RECT 1807.025000 -0.085000 1807.195000 0.085000 ;
      RECT 1807.025000  2.635000 1807.195000 2.805000 ;
      RECT 1807.485000 -0.085000 1807.655000 0.085000 ;
      RECT 1807.485000  2.635000 1807.655000 2.805000 ;
      RECT 1807.945000 -0.085000 1808.115000 0.085000 ;
      RECT 1807.945000  2.635000 1808.115000 2.805000 ;
      RECT 1808.405000 -0.085000 1808.575000 0.085000 ;
      RECT 1808.405000  2.635000 1808.575000 2.805000 ;
      RECT 1808.865000 -0.085000 1809.035000 0.085000 ;
      RECT 1808.865000  2.635000 1809.035000 2.805000 ;
      RECT 1809.325000 -0.085000 1809.495000 0.085000 ;
      RECT 1809.325000  2.635000 1809.495000 2.805000 ;
      RECT 1809.785000 -0.085000 1809.955000 0.085000 ;
      RECT 1809.785000  2.635000 1809.955000 2.805000 ;
      RECT 1810.245000 -0.085000 1810.415000 0.085000 ;
      RECT 1810.245000  2.635000 1810.415000 2.805000 ;
      RECT 1810.705000 -0.085000 1810.875000 0.085000 ;
      RECT 1810.705000  2.635000 1810.875000 2.805000 ;
      RECT 1811.165000 -0.085000 1811.335000 0.085000 ;
      RECT 1811.165000  2.635000 1811.335000 2.805000 ;
      RECT 1811.625000 -0.085000 1811.795000 0.085000 ;
      RECT 1811.625000  2.635000 1811.795000 2.805000 ;
      RECT 1812.085000 -0.085000 1812.255000 0.085000 ;
      RECT 1812.085000  2.635000 1812.255000 2.805000 ;
      RECT 1812.545000 -0.085000 1812.715000 0.085000 ;
      RECT 1812.545000  2.635000 1812.715000 2.805000 ;
      RECT 1813.005000 -0.085000 1813.175000 0.085000 ;
      RECT 1813.005000  2.635000 1813.175000 2.805000 ;
      RECT 1813.465000 -0.085000 1813.635000 0.085000 ;
      RECT 1813.465000  2.635000 1813.635000 2.805000 ;
      RECT 1813.925000 -0.085000 1814.095000 0.085000 ;
      RECT 1813.925000  2.635000 1814.095000 2.805000 ;
      RECT 1814.385000 -0.085000 1814.555000 0.085000 ;
      RECT 1814.385000  2.635000 1814.555000 2.805000 ;
      RECT 1814.845000 -0.085000 1815.015000 0.085000 ;
      RECT 1814.845000  2.635000 1815.015000 2.805000 ;
      RECT 1815.305000 -0.085000 1815.475000 0.085000 ;
      RECT 1815.305000  2.635000 1815.475000 2.805000 ;
      RECT 1815.765000 -0.085000 1815.935000 0.085000 ;
      RECT 1815.765000  2.635000 1815.935000 2.805000 ;
      RECT 1816.225000 -0.085000 1816.395000 0.085000 ;
      RECT 1816.225000  2.635000 1816.395000 2.805000 ;
      RECT 1816.685000 -0.085000 1816.855000 0.085000 ;
      RECT 1816.685000  2.635000 1816.855000 2.805000 ;
      RECT 1817.145000 -0.085000 1817.315000 0.085000 ;
      RECT 1817.145000  2.635000 1817.315000 2.805000 ;
      RECT 1817.605000 -0.085000 1817.775000 0.085000 ;
      RECT 1817.605000  2.635000 1817.775000 2.805000 ;
      RECT 1818.065000 -0.085000 1818.235000 0.085000 ;
      RECT 1818.065000  2.635000 1818.235000 2.805000 ;
      RECT 1818.525000 -0.085000 1818.695000 0.085000 ;
      RECT 1818.525000  2.635000 1818.695000 2.805000 ;
      RECT 1818.985000 -0.085000 1819.155000 0.085000 ;
      RECT 1818.985000  2.635000 1819.155000 2.805000 ;
      RECT 1819.445000 -0.085000 1819.615000 0.085000 ;
      RECT 1819.445000  2.635000 1819.615000 2.805000 ;
      RECT 1819.905000 -0.085000 1820.075000 0.085000 ;
      RECT 1819.905000  2.635000 1820.075000 2.805000 ;
      RECT 1820.365000 -0.085000 1820.535000 0.085000 ;
      RECT 1820.365000  2.635000 1820.535000 2.805000 ;
      RECT 1820.825000 -0.085000 1820.995000 0.085000 ;
      RECT 1820.825000  2.635000 1820.995000 2.805000 ;
      RECT 1821.285000 -0.085000 1821.455000 0.085000 ;
      RECT 1821.285000  2.635000 1821.455000 2.805000 ;
      RECT 1821.745000 -0.085000 1821.915000 0.085000 ;
      RECT 1821.745000  2.635000 1821.915000 2.805000 ;
      RECT 1822.205000 -0.085000 1822.375000 0.085000 ;
      RECT 1822.205000  2.635000 1822.375000 2.805000 ;
      RECT 1822.665000 -0.085000 1822.835000 0.085000 ;
      RECT 1822.665000  2.635000 1822.835000 2.805000 ;
      RECT 1823.125000 -0.085000 1823.295000 0.085000 ;
      RECT 1823.125000  2.635000 1823.295000 2.805000 ;
      RECT 1823.585000 -0.085000 1823.755000 0.085000 ;
      RECT 1823.585000  2.635000 1823.755000 2.805000 ;
      RECT 1824.045000 -0.085000 1824.215000 0.085000 ;
      RECT 1824.045000  2.635000 1824.215000 2.805000 ;
      RECT 1824.505000 -0.085000 1824.675000 0.085000 ;
      RECT 1824.505000  2.635000 1824.675000 2.805000 ;
      RECT 1824.965000 -0.085000 1825.135000 0.085000 ;
      RECT 1824.965000  2.635000 1825.135000 2.805000 ;
      RECT 1825.425000 -0.085000 1825.595000 0.085000 ;
      RECT 1825.425000  2.635000 1825.595000 2.805000 ;
      RECT 1825.885000 -0.085000 1826.055000 0.085000 ;
      RECT 1825.885000  2.635000 1826.055000 2.805000 ;
      RECT 1826.345000 -0.085000 1826.515000 0.085000 ;
      RECT 1826.345000  2.635000 1826.515000 2.805000 ;
      RECT 1826.805000 -0.085000 1826.975000 0.085000 ;
      RECT 1826.805000  2.635000 1826.975000 2.805000 ;
      RECT 1827.265000 -0.085000 1827.435000 0.085000 ;
      RECT 1827.265000  2.635000 1827.435000 2.805000 ;
      RECT 1827.725000 -0.085000 1827.895000 0.085000 ;
      RECT 1827.725000  2.635000 1827.895000 2.805000 ;
      RECT 1828.185000 -0.085000 1828.355000 0.085000 ;
      RECT 1828.185000  2.635000 1828.355000 2.805000 ;
      RECT 1828.645000 -0.085000 1828.815000 0.085000 ;
      RECT 1828.645000  2.635000 1828.815000 2.805000 ;
      RECT 1829.105000 -0.085000 1829.275000 0.085000 ;
      RECT 1829.105000  2.635000 1829.275000 2.805000 ;
      RECT 1829.565000 -0.085000 1829.735000 0.085000 ;
      RECT 1829.565000  2.635000 1829.735000 2.805000 ;
      RECT 1830.025000 -0.085000 1830.195000 0.085000 ;
      RECT 1830.025000  2.635000 1830.195000 2.805000 ;
      RECT 1830.485000 -0.085000 1830.655000 0.085000 ;
      RECT 1830.485000  2.635000 1830.655000 2.805000 ;
      RECT 1830.945000 -0.085000 1831.115000 0.085000 ;
      RECT 1830.945000  2.635000 1831.115000 2.805000 ;
      RECT 1831.405000 -0.085000 1831.575000 0.085000 ;
      RECT 1831.405000  2.635000 1831.575000 2.805000 ;
      RECT 1831.865000 -0.085000 1832.035000 0.085000 ;
      RECT 1831.865000  2.635000 1832.035000 2.805000 ;
      RECT 1832.325000 -0.085000 1832.495000 0.085000 ;
      RECT 1832.325000  2.635000 1832.495000 2.805000 ;
      RECT 1832.785000 -0.085000 1832.955000 0.085000 ;
      RECT 1832.785000  2.635000 1832.955000 2.805000 ;
      RECT 1833.245000 -0.085000 1833.415000 0.085000 ;
      RECT 1833.245000  2.635000 1833.415000 2.805000 ;
      RECT 1833.705000 -0.085000 1833.875000 0.085000 ;
      RECT 1833.705000  2.635000 1833.875000 2.805000 ;
      RECT 1834.165000 -0.085000 1834.335000 0.085000 ;
      RECT 1834.165000  1.785000 1834.335000 1.955000 ;
      RECT 1834.165000  2.635000 1834.335000 2.805000 ;
      RECT 1834.625000 -0.085000 1834.795000 0.085000 ;
      RECT 1834.625000  2.635000 1834.795000 2.805000 ;
      RECT 1835.085000 -0.085000 1835.255000 0.085000 ;
      RECT 1835.085000  2.635000 1835.255000 2.805000 ;
      RECT 1835.545000 -0.085000 1835.715000 0.085000 ;
      RECT 1835.545000  2.635000 1835.715000 2.805000 ;
      RECT 1836.005000 -0.085000 1836.175000 0.085000 ;
      RECT 1836.005000  2.635000 1836.175000 2.805000 ;
      RECT 1836.465000 -0.085000 1836.635000 0.085000 ;
      RECT 1836.465000  1.785000 1836.635000 1.955000 ;
      RECT 1836.465000  2.635000 1836.635000 2.805000 ;
      RECT 1836.925000 -0.085000 1837.095000 0.085000 ;
      RECT 1836.925000  2.635000 1837.095000 2.805000 ;
      RECT 1837.385000 -0.085000 1837.555000 0.085000 ;
      RECT 1837.385000  2.635000 1837.555000 2.805000 ;
      RECT 1837.845000 -0.085000 1838.015000 0.085000 ;
      RECT 1837.845000  2.635000 1838.015000 2.805000 ;
      RECT 1838.305000 -0.085000 1838.475000 0.085000 ;
      RECT 1838.305000  1.785000 1838.475000 1.955000 ;
      RECT 1838.305000  2.635000 1838.475000 2.805000 ;
      RECT 1838.765000 -0.085000 1838.935000 0.085000 ;
      RECT 1838.765000  2.635000 1838.935000 2.805000 ;
      RECT 1839.225000 -0.085000 1839.395000 0.085000 ;
      RECT 1839.225000  2.635000 1839.395000 2.805000 ;
      RECT 1839.685000 -0.085000 1839.855000 0.085000 ;
      RECT 1839.685000  2.635000 1839.855000 2.805000 ;
      RECT 1840.145000 -0.085000 1840.315000 0.085000 ;
      RECT 1840.145000  2.635000 1840.315000 2.805000 ;
      RECT 1840.605000 -0.085000 1840.775000 0.085000 ;
      RECT 1840.605000  1.785000 1840.775000 1.955000 ;
      RECT 1840.605000  2.635000 1840.775000 2.805000 ;
      RECT 1841.065000 -0.085000 1841.235000 0.085000 ;
      RECT 1841.065000  2.635000 1841.235000 2.805000 ;
      RECT 1841.525000 -0.085000 1841.695000 0.085000 ;
      RECT 1841.525000  2.635000 1841.695000 2.805000 ;
      RECT 1841.985000 -0.085000 1842.155000 0.085000 ;
      RECT 1841.985000  2.635000 1842.155000 2.805000 ;
      RECT 1842.445000 -0.085000 1842.615000 0.085000 ;
      RECT 1842.445000  2.635000 1842.615000 2.805000 ;
      RECT 1842.905000 -0.085000 1843.075000 0.085000 ;
      RECT 1842.905000  2.635000 1843.075000 2.805000 ;
      RECT 1843.365000 -0.085000 1843.535000 0.085000 ;
      RECT 1843.365000  2.635000 1843.535000 2.805000 ;
      RECT 1843.825000 -0.085000 1843.995000 0.085000 ;
      RECT 1843.825000  1.785000 1843.995000 1.955000 ;
      RECT 1843.825000  2.635000 1843.995000 2.805000 ;
      RECT 1844.285000 -0.085000 1844.455000 0.085000 ;
      RECT 1844.285000  2.635000 1844.455000 2.805000 ;
      RECT 1844.745000 -0.085000 1844.915000 0.085000 ;
      RECT 1844.745000  2.635000 1844.915000 2.805000 ;
      RECT 1845.205000 -0.085000 1845.375000 0.085000 ;
      RECT 1845.205000  2.635000 1845.375000 2.805000 ;
      RECT 1845.665000 -0.085000 1845.835000 0.085000 ;
      RECT 1845.665000  2.635000 1845.835000 2.805000 ;
      RECT 1846.125000 -0.085000 1846.295000 0.085000 ;
      RECT 1846.125000  2.635000 1846.295000 2.805000 ;
      RECT 1846.585000 -0.085000 1846.755000 0.085000 ;
      RECT 1846.585000  2.635000 1846.755000 2.805000 ;
      RECT 1847.045000 -0.085000 1847.215000 0.085000 ;
      RECT 1847.045000  1.785000 1847.215000 1.955000 ;
      RECT 1847.045000  2.635000 1847.215000 2.805000 ;
      RECT 1847.505000 -0.085000 1847.675000 0.085000 ;
      RECT 1847.505000  2.635000 1847.675000 2.805000 ;
      RECT 1847.965000 -0.085000 1848.135000 0.085000 ;
      RECT 1847.965000  2.635000 1848.135000 2.805000 ;
      RECT 1848.425000 -0.085000 1848.595000 0.085000 ;
      RECT 1848.425000  2.635000 1848.595000 2.805000 ;
      RECT 1848.885000 -0.085000 1849.055000 0.085000 ;
      RECT 1848.885000  2.635000 1849.055000 2.805000 ;
      RECT 1849.345000 -0.085000 1849.515000 0.085000 ;
      RECT 1849.345000  2.635000 1849.515000 2.805000 ;
      RECT 1849.805000 -0.085000 1849.975000 0.085000 ;
      RECT 1849.805000  2.635000 1849.975000 2.805000 ;
      RECT 1850.265000 -0.085000 1850.435000 0.085000 ;
      RECT 1850.265000  1.785000 1850.435000 1.955000 ;
      RECT 1850.265000  2.635000 1850.435000 2.805000 ;
      RECT 1850.725000 -0.085000 1850.895000 0.085000 ;
      RECT 1850.725000  2.635000 1850.895000 2.805000 ;
      RECT 1851.185000 -0.085000 1851.355000 0.085000 ;
      RECT 1851.185000  2.635000 1851.355000 2.805000 ;
      RECT 1851.645000 -0.085000 1851.815000 0.085000 ;
      RECT 1851.645000  2.635000 1851.815000 2.805000 ;
      RECT 1852.105000 -0.085000 1852.275000 0.085000 ;
      RECT 1852.105000  2.635000 1852.275000 2.805000 ;
      RECT 1852.565000 -0.085000 1852.735000 0.085000 ;
      RECT 1852.565000  2.635000 1852.735000 2.805000 ;
      RECT 1853.025000 -0.085000 1853.195000 0.085000 ;
      RECT 1853.025000  2.635000 1853.195000 2.805000 ;
      RECT 1853.485000 -0.085000 1853.655000 0.085000 ;
      RECT 1853.485000  1.785000 1853.655000 1.955000 ;
      RECT 1853.485000  2.635000 1853.655000 2.805000 ;
      RECT 1853.945000 -0.085000 1854.115000 0.085000 ;
      RECT 1853.945000  2.635000 1854.115000 2.805000 ;
      RECT 1854.405000 -0.085000 1854.575000 0.085000 ;
      RECT 1854.405000  2.635000 1854.575000 2.805000 ;
      RECT 1854.865000 -0.085000 1855.035000 0.085000 ;
      RECT 1854.865000  2.635000 1855.035000 2.805000 ;
      RECT 1855.325000 -0.085000 1855.495000 0.085000 ;
      RECT 1855.325000  2.635000 1855.495000 2.805000 ;
      RECT 1855.785000 -0.085000 1855.955000 0.085000 ;
      RECT 1855.785000  2.635000 1855.955000 2.805000 ;
      RECT 1856.245000 -0.085000 1856.415000 0.085000 ;
      RECT 1856.245000  2.635000 1856.415000 2.805000 ;
      RECT 1856.705000 -0.085000 1856.875000 0.085000 ;
      RECT 1856.705000  2.635000 1856.875000 2.805000 ;
      RECT 1857.165000 -0.085000 1857.335000 0.085000 ;
      RECT 1857.165000  2.635000 1857.335000 2.805000 ;
      RECT 1857.625000 -0.085000 1857.795000 0.085000 ;
      RECT 1857.625000  2.635000 1857.795000 2.805000 ;
      RECT 1858.085000 -0.085000 1858.255000 0.085000 ;
      RECT 1858.085000  2.635000 1858.255000 2.805000 ;
      RECT 1858.545000 -0.085000 1858.715000 0.085000 ;
      RECT 1858.545000  2.635000 1858.715000 2.805000 ;
      RECT 1858.685000  1.785000 1858.855000 1.955000 ;
      RECT 1859.005000 -0.085000 1859.175000 0.085000 ;
      RECT 1859.005000  2.635000 1859.175000 2.805000 ;
      RECT 1859.465000 -0.085000 1859.635000 0.085000 ;
      RECT 1859.465000  2.635000 1859.635000 2.805000 ;
      RECT 1859.625000  1.785000 1859.795000 1.955000 ;
      RECT 1859.925000 -0.085000 1860.095000 0.085000 ;
      RECT 1859.925000  2.635000 1860.095000 2.805000 ;
      RECT 1860.385000 -0.085000 1860.555000 0.085000 ;
      RECT 1860.385000  2.635000 1860.555000 2.805000 ;
      RECT 1860.845000 -0.085000 1861.015000 0.085000 ;
      RECT 1860.845000  2.635000 1861.015000 2.805000 ;
      RECT 1861.305000 -0.085000 1861.475000 0.085000 ;
      RECT 1861.305000  2.635000 1861.475000 2.805000 ;
      RECT 1861.765000 -0.085000 1861.935000 0.085000 ;
      RECT 1861.765000  2.635000 1861.935000 2.805000 ;
      RECT 1862.225000 -0.085000 1862.395000 0.085000 ;
      RECT 1862.225000  2.635000 1862.395000 2.805000 ;
      RECT 1862.685000 -0.085000 1862.855000 0.085000 ;
      RECT 1862.685000  2.635000 1862.855000 2.805000 ;
      RECT 1863.145000 -0.085000 1863.315000 0.085000 ;
      RECT 1863.145000  2.635000 1863.315000 2.805000 ;
      RECT 1863.605000 -0.085000 1863.775000 0.085000 ;
      RECT 1863.605000  2.635000 1863.775000 2.805000 ;
      RECT 1864.065000 -0.085000 1864.235000 0.085000 ;
      RECT 1864.065000  2.635000 1864.235000 2.805000 ;
      RECT 1864.365000  1.785000 1864.535000 1.955000 ;
      RECT 1864.525000 -0.085000 1864.695000 0.085000 ;
      RECT 1864.525000  2.635000 1864.695000 2.805000 ;
      RECT 1864.985000 -0.085000 1865.155000 0.085000 ;
      RECT 1864.985000  2.635000 1865.155000 2.805000 ;
      RECT 1865.305000  1.785000 1865.475000 1.955000 ;
      RECT 1865.445000 -0.085000 1865.615000 0.085000 ;
      RECT 1865.445000  2.635000 1865.615000 2.805000 ;
      RECT 1865.905000 -0.085000 1866.075000 0.085000 ;
      RECT 1865.905000  2.635000 1866.075000 2.805000 ;
      RECT 1866.365000 -0.085000 1866.535000 0.085000 ;
      RECT 1866.365000  2.635000 1866.535000 2.805000 ;
      RECT 1866.825000 -0.085000 1866.995000 0.085000 ;
      RECT 1866.825000  2.635000 1866.995000 2.805000 ;
      RECT 1867.285000 -0.085000 1867.455000 0.085000 ;
      RECT 1867.285000  2.635000 1867.455000 2.805000 ;
      RECT 1867.745000 -0.085000 1867.915000 0.085000 ;
      RECT 1867.745000  2.635000 1867.915000 2.805000 ;
      RECT 1868.205000 -0.085000 1868.375000 0.085000 ;
      RECT 1868.205000  2.635000 1868.375000 2.805000 ;
      RECT 1868.665000 -0.085000 1868.835000 0.085000 ;
      RECT 1868.665000  2.635000 1868.835000 2.805000 ;
      RECT 1869.125000 -0.085000 1869.295000 0.085000 ;
      RECT 1869.125000  2.635000 1869.295000 2.805000 ;
      RECT 1869.585000 -0.085000 1869.755000 0.085000 ;
      RECT 1869.585000  2.635000 1869.755000 2.805000 ;
      RECT 1870.045000 -0.085000 1870.215000 0.085000 ;
      RECT 1870.045000  2.635000 1870.215000 2.805000 ;
      RECT 1870.505000 -0.085000 1870.675000 0.085000 ;
      RECT 1870.505000  2.635000 1870.675000 2.805000 ;
      RECT 1870.965000 -0.085000 1871.135000 0.085000 ;
      RECT 1870.965000  2.635000 1871.135000 2.805000 ;
      RECT 1871.425000 -0.085000 1871.595000 0.085000 ;
      RECT 1871.425000  2.635000 1871.595000 2.805000 ;
      RECT 1871.565000  1.785000 1871.735000 1.955000 ;
      RECT 1871.885000 -0.085000 1872.055000 0.085000 ;
      RECT 1871.885000  2.635000 1872.055000 2.805000 ;
      RECT 1872.345000 -0.085000 1872.515000 0.085000 ;
      RECT 1872.345000  2.635000 1872.515000 2.805000 ;
      RECT 1872.505000  1.785000 1872.675000 1.955000 ;
      RECT 1872.805000 -0.085000 1872.975000 0.085000 ;
      RECT 1872.805000  2.635000 1872.975000 2.805000 ;
      RECT 1873.265000 -0.085000 1873.435000 0.085000 ;
      RECT 1873.265000  2.635000 1873.435000 2.805000 ;
      RECT 1873.725000 -0.085000 1873.895000 0.085000 ;
      RECT 1873.725000  2.635000 1873.895000 2.805000 ;
      RECT 1874.185000 -0.085000 1874.355000 0.085000 ;
      RECT 1874.185000  2.635000 1874.355000 2.805000 ;
      RECT 1874.645000 -0.085000 1874.815000 0.085000 ;
      RECT 1874.645000  2.635000 1874.815000 2.805000 ;
      RECT 1875.105000 -0.085000 1875.275000 0.085000 ;
      RECT 1875.105000  2.635000 1875.275000 2.805000 ;
      RECT 1875.565000 -0.085000 1875.735000 0.085000 ;
      RECT 1875.565000  2.635000 1875.735000 2.805000 ;
      RECT 1876.025000 -0.085000 1876.195000 0.085000 ;
      RECT 1876.025000  2.635000 1876.195000 2.805000 ;
      RECT 1876.485000 -0.085000 1876.655000 0.085000 ;
      RECT 1876.485000  2.635000 1876.655000 2.805000 ;
      RECT 1876.945000 -0.085000 1877.115000 0.085000 ;
      RECT 1876.945000  2.635000 1877.115000 2.805000 ;
      RECT 1877.245000  1.785000 1877.415000 1.955000 ;
      RECT 1877.405000 -0.085000 1877.575000 0.085000 ;
      RECT 1877.405000  2.635000 1877.575000 2.805000 ;
      RECT 1877.865000 -0.085000 1878.035000 0.085000 ;
      RECT 1877.865000  2.635000 1878.035000 2.805000 ;
      RECT 1878.185000  1.785000 1878.355000 1.955000 ;
      RECT 1878.325000 -0.085000 1878.495000 0.085000 ;
      RECT 1878.325000  2.635000 1878.495000 2.805000 ;
      RECT 1878.785000 -0.085000 1878.955000 0.085000 ;
      RECT 1878.785000  2.635000 1878.955000 2.805000 ;
      RECT 1879.245000 -0.085000 1879.415000 0.085000 ;
      RECT 1879.245000  2.635000 1879.415000 2.805000 ;
      RECT 1879.705000 -0.085000 1879.875000 0.085000 ;
      RECT 1879.705000  2.635000 1879.875000 2.805000 ;
      RECT 1880.165000 -0.085000 1880.335000 0.085000 ;
      RECT 1880.165000  2.635000 1880.335000 2.805000 ;
      RECT 1880.625000 -0.085000 1880.795000 0.085000 ;
      RECT 1880.625000  2.635000 1880.795000 2.805000 ;
      RECT 1881.085000 -0.085000 1881.255000 0.085000 ;
      RECT 1881.085000  2.635000 1881.255000 2.805000 ;
      RECT 1881.545000 -0.085000 1881.715000 0.085000 ;
      RECT 1881.545000  2.635000 1881.715000 2.805000 ;
      RECT 1882.005000 -0.085000 1882.175000 0.085000 ;
      RECT 1882.005000  2.635000 1882.175000 2.805000 ;
      RECT 1882.465000 -0.085000 1882.635000 0.085000 ;
      RECT 1882.465000  2.635000 1882.635000 2.805000 ;
      RECT 1882.925000 -0.085000 1883.095000 0.085000 ;
      RECT 1882.925000  1.785000 1883.095000 1.955000 ;
      RECT 1882.925000  2.635000 1883.095000 2.805000 ;
      RECT 1883.385000 -0.085000 1883.555000 0.085000 ;
      RECT 1883.385000  2.635000 1883.555000 2.805000 ;
      RECT 1883.845000 -0.085000 1884.015000 0.085000 ;
      RECT 1883.845000  2.635000 1884.015000 2.805000 ;
      RECT 1884.305000 -0.085000 1884.475000 0.085000 ;
      RECT 1884.305000  2.635000 1884.475000 2.805000 ;
      RECT 1884.765000 -0.085000 1884.935000 0.085000 ;
      RECT 1884.765000  2.635000 1884.935000 2.805000 ;
      RECT 1885.225000 -0.085000 1885.395000 0.085000 ;
      RECT 1885.225000  1.785000 1885.395000 1.955000 ;
      RECT 1885.225000  2.635000 1885.395000 2.805000 ;
      RECT 1885.685000 -0.085000 1885.855000 0.085000 ;
      RECT 1885.685000  2.635000 1885.855000 2.805000 ;
      RECT 1886.145000 -0.085000 1886.315000 0.085000 ;
      RECT 1886.145000  2.635000 1886.315000 2.805000 ;
      RECT 1886.605000 -0.085000 1886.775000 0.085000 ;
      RECT 1886.605000  2.635000 1886.775000 2.805000 ;
      RECT 1887.065000 -0.085000 1887.235000 0.085000 ;
      RECT 1887.065000  1.785000 1887.235000 1.955000 ;
      RECT 1887.065000  2.635000 1887.235000 2.805000 ;
      RECT 1887.525000 -0.085000 1887.695000 0.085000 ;
      RECT 1887.525000  2.635000 1887.695000 2.805000 ;
      RECT 1887.985000 -0.085000 1888.155000 0.085000 ;
      RECT 1887.985000  2.635000 1888.155000 2.805000 ;
      RECT 1888.445000 -0.085000 1888.615000 0.085000 ;
      RECT 1888.445000  2.635000 1888.615000 2.805000 ;
      RECT 1888.905000 -0.085000 1889.075000 0.085000 ;
      RECT 1888.905000  2.635000 1889.075000 2.805000 ;
      RECT 1889.365000 -0.085000 1889.535000 0.085000 ;
      RECT 1889.365000  1.785000 1889.535000 1.955000 ;
      RECT 1889.365000  2.635000 1889.535000 2.805000 ;
      RECT 1889.825000 -0.085000 1889.995000 0.085000 ;
      RECT 1889.825000  2.635000 1889.995000 2.805000 ;
      RECT 1890.285000 -0.085000 1890.455000 0.085000 ;
      RECT 1890.285000  2.635000 1890.455000 2.805000 ;
      RECT 1890.745000 -0.085000 1890.915000 0.085000 ;
      RECT 1890.745000  2.635000 1890.915000 2.805000 ;
      RECT 1891.205000 -0.085000 1891.375000 0.085000 ;
      RECT 1891.205000  1.785000 1891.375000 1.955000 ;
      RECT 1891.205000  2.635000 1891.375000 2.805000 ;
      RECT 1891.665000 -0.085000 1891.835000 0.085000 ;
      RECT 1891.665000  2.635000 1891.835000 2.805000 ;
      RECT 1892.125000 -0.085000 1892.295000 0.085000 ;
      RECT 1892.125000  2.635000 1892.295000 2.805000 ;
      RECT 1892.585000 -0.085000 1892.755000 0.085000 ;
      RECT 1892.585000  2.635000 1892.755000 2.805000 ;
      RECT 1893.045000 -0.085000 1893.215000 0.085000 ;
      RECT 1893.045000  2.635000 1893.215000 2.805000 ;
      RECT 1893.505000 -0.085000 1893.675000 0.085000 ;
      RECT 1893.505000  1.785000 1893.675000 1.955000 ;
      RECT 1893.505000  2.635000 1893.675000 2.805000 ;
      RECT 1893.965000 -0.085000 1894.135000 0.085000 ;
      RECT 1893.965000  2.635000 1894.135000 2.805000 ;
      RECT 1894.425000 -0.085000 1894.595000 0.085000 ;
      RECT 1894.425000  2.635000 1894.595000 2.805000 ;
      RECT 1894.885000 -0.085000 1895.055000 0.085000 ;
      RECT 1894.885000  2.635000 1895.055000 2.805000 ;
      RECT 1895.345000 -0.085000 1895.515000 0.085000 ;
      RECT 1895.345000  1.785000 1895.515000 1.955000 ;
      RECT 1895.345000  2.635000 1895.515000 2.805000 ;
      RECT 1895.805000 -0.085000 1895.975000 0.085000 ;
      RECT 1895.805000  2.635000 1895.975000 2.805000 ;
      RECT 1896.265000 -0.085000 1896.435000 0.085000 ;
      RECT 1896.265000  2.635000 1896.435000 2.805000 ;
      RECT 1896.725000 -0.085000 1896.895000 0.085000 ;
      RECT 1896.725000  2.635000 1896.895000 2.805000 ;
      RECT 1897.185000 -0.085000 1897.355000 0.085000 ;
      RECT 1897.185000  2.635000 1897.355000 2.805000 ;
      RECT 1897.645000 -0.085000 1897.815000 0.085000 ;
      RECT 1897.645000  1.785000 1897.815000 1.955000 ;
      RECT 1897.645000  2.635000 1897.815000 2.805000 ;
      RECT 1898.105000 -0.085000 1898.275000 0.085000 ;
      RECT 1898.105000  2.635000 1898.275000 2.805000 ;
      RECT 1898.565000 -0.085000 1898.735000 0.085000 ;
      RECT 1898.565000  2.635000 1898.735000 2.805000 ;
      RECT 1899.025000 -0.085000 1899.195000 0.085000 ;
      RECT 1899.025000  2.635000 1899.195000 2.805000 ;
      RECT 1899.485000 -0.085000 1899.655000 0.085000 ;
      RECT 1899.485000  2.635000 1899.655000 2.805000 ;
      RECT 1899.945000 -0.085000 1900.115000 0.085000 ;
      RECT 1899.945000  2.635000 1900.115000 2.805000 ;
      RECT 1900.405000 -0.085000 1900.575000 0.085000 ;
      RECT 1900.405000  2.635000 1900.575000 2.805000 ;
      RECT 1900.865000 -0.085000 1901.035000 0.085000 ;
      RECT 1900.865000  1.785000 1901.035000 1.955000 ;
      RECT 1900.865000  2.635000 1901.035000 2.805000 ;
      RECT 1901.325000 -0.085000 1901.495000 0.085000 ;
      RECT 1901.325000  2.635000 1901.495000 2.805000 ;
      RECT 1901.785000 -0.085000 1901.955000 0.085000 ;
      RECT 1901.785000  2.635000 1901.955000 2.805000 ;
      RECT 1902.245000 -0.085000 1902.415000 0.085000 ;
      RECT 1902.245000  2.635000 1902.415000 2.805000 ;
      RECT 1902.705000 -0.085000 1902.875000 0.085000 ;
      RECT 1902.705000  2.635000 1902.875000 2.805000 ;
      RECT 1903.165000 -0.085000 1903.335000 0.085000 ;
      RECT 1903.165000  2.635000 1903.335000 2.805000 ;
      RECT 1903.625000 -0.085000 1903.795000 0.085000 ;
      RECT 1903.625000  2.635000 1903.795000 2.805000 ;
      RECT 1904.085000 -0.085000 1904.255000 0.085000 ;
      RECT 1904.085000  1.785000 1904.255000 1.955000 ;
      RECT 1904.085000  2.635000 1904.255000 2.805000 ;
      RECT 1904.545000 -0.085000 1904.715000 0.085000 ;
      RECT 1904.545000  2.635000 1904.715000 2.805000 ;
      RECT 1905.005000 -0.085000 1905.175000 0.085000 ;
      RECT 1905.005000  2.635000 1905.175000 2.805000 ;
      RECT 1905.465000 -0.085000 1905.635000 0.085000 ;
      RECT 1905.465000  2.635000 1905.635000 2.805000 ;
      RECT 1905.925000 -0.085000 1906.095000 0.085000 ;
      RECT 1905.925000  2.635000 1906.095000 2.805000 ;
      RECT 1906.385000 -0.085000 1906.555000 0.085000 ;
      RECT 1906.385000  2.635000 1906.555000 2.805000 ;
      RECT 1906.845000 -0.085000 1907.015000 0.085000 ;
      RECT 1906.845000  2.635000 1907.015000 2.805000 ;
      RECT 1907.305000 -0.085000 1907.475000 0.085000 ;
      RECT 1907.305000  1.785000 1907.475000 1.955000 ;
      RECT 1907.305000  2.635000 1907.475000 2.805000 ;
      RECT 1907.765000 -0.085000 1907.935000 0.085000 ;
      RECT 1907.765000  2.635000 1907.935000 2.805000 ;
      RECT 1908.225000 -0.085000 1908.395000 0.085000 ;
      RECT 1908.225000  2.635000 1908.395000 2.805000 ;
      RECT 1908.685000 -0.085000 1908.855000 0.085000 ;
      RECT 1908.685000  2.635000 1908.855000 2.805000 ;
      RECT 1909.145000 -0.085000 1909.315000 0.085000 ;
      RECT 1909.145000  2.635000 1909.315000 2.805000 ;
      RECT 1909.605000 -0.085000 1909.775000 0.085000 ;
      RECT 1909.605000  2.635000 1909.775000 2.805000 ;
      RECT 1910.065000 -0.085000 1910.235000 0.085000 ;
      RECT 1910.065000  2.635000 1910.235000 2.805000 ;
      RECT 1910.525000 -0.085000 1910.695000 0.085000 ;
      RECT 1910.525000  1.785000 1910.695000 1.955000 ;
      RECT 1910.525000  2.635000 1910.695000 2.805000 ;
      RECT 1910.985000 -0.085000 1911.155000 0.085000 ;
      RECT 1910.985000  2.635000 1911.155000 2.805000 ;
      RECT 1911.445000 -0.085000 1911.615000 0.085000 ;
      RECT 1911.445000  2.635000 1911.615000 2.805000 ;
      RECT 1911.905000 -0.085000 1912.075000 0.085000 ;
      RECT 1911.905000  2.635000 1912.075000 2.805000 ;
      RECT 1912.365000 -0.085000 1912.535000 0.085000 ;
      RECT 1912.365000  2.635000 1912.535000 2.805000 ;
      RECT 1912.825000 -0.085000 1912.995000 0.085000 ;
      RECT 1912.825000  2.635000 1912.995000 2.805000 ;
      RECT 1913.285000 -0.085000 1913.455000 0.085000 ;
      RECT 1913.285000  2.635000 1913.455000 2.805000 ;
      RECT 1913.745000 -0.085000 1913.915000 0.085000 ;
      RECT 1913.745000  1.785000 1913.915000 1.955000 ;
      RECT 1913.745000  2.635000 1913.915000 2.805000 ;
      RECT 1914.205000 -0.085000 1914.375000 0.085000 ;
      RECT 1914.205000  2.635000 1914.375000 2.805000 ;
      RECT 1914.665000 -0.085000 1914.835000 0.085000 ;
      RECT 1914.665000  2.635000 1914.835000 2.805000 ;
      RECT 1915.125000 -0.085000 1915.295000 0.085000 ;
      RECT 1915.125000  2.635000 1915.295000 2.805000 ;
      RECT 1915.585000 -0.085000 1915.755000 0.085000 ;
      RECT 1915.585000  2.635000 1915.755000 2.805000 ;
      RECT 1916.045000 -0.085000 1916.215000 0.085000 ;
      RECT 1916.045000  2.635000 1916.215000 2.805000 ;
      RECT 1916.505000 -0.085000 1916.675000 0.085000 ;
      RECT 1916.505000  2.635000 1916.675000 2.805000 ;
      RECT 1916.965000 -0.085000 1917.135000 0.085000 ;
      RECT 1916.965000  1.785000 1917.135000 1.955000 ;
      RECT 1916.965000  2.635000 1917.135000 2.805000 ;
      RECT 1917.425000 -0.085000 1917.595000 0.085000 ;
      RECT 1917.425000  2.635000 1917.595000 2.805000 ;
      RECT 1917.885000 -0.085000 1918.055000 0.085000 ;
      RECT 1917.885000  2.635000 1918.055000 2.805000 ;
      RECT 1918.345000 -0.085000 1918.515000 0.085000 ;
      RECT 1918.345000  2.635000 1918.515000 2.805000 ;
      RECT 1918.805000 -0.085000 1918.975000 0.085000 ;
      RECT 1918.805000  2.635000 1918.975000 2.805000 ;
      RECT 1919.265000 -0.085000 1919.435000 0.085000 ;
      RECT 1919.265000  2.635000 1919.435000 2.805000 ;
      RECT 1919.725000 -0.085000 1919.895000 0.085000 ;
      RECT 1919.725000  2.635000 1919.895000 2.805000 ;
      RECT 1920.185000 -0.085000 1920.355000 0.085000 ;
      RECT 1920.185000  1.785000 1920.355000 1.955000 ;
      RECT 1920.185000  2.635000 1920.355000 2.805000 ;
      RECT 1920.645000 -0.085000 1920.815000 0.085000 ;
      RECT 1920.645000  2.635000 1920.815000 2.805000 ;
      RECT 1921.105000 -0.085000 1921.275000 0.085000 ;
      RECT 1921.105000  2.635000 1921.275000 2.805000 ;
      RECT 1921.565000 -0.085000 1921.735000 0.085000 ;
      RECT 1921.565000  2.635000 1921.735000 2.805000 ;
      RECT 1922.025000 -0.085000 1922.195000 0.085000 ;
      RECT 1922.025000  2.635000 1922.195000 2.805000 ;
      RECT 1922.485000 -0.085000 1922.655000 0.085000 ;
      RECT 1922.485000  2.635000 1922.655000 2.805000 ;
      RECT 1922.945000 -0.085000 1923.115000 0.085000 ;
      RECT 1922.945000  2.635000 1923.115000 2.805000 ;
      RECT 1923.405000 -0.085000 1923.575000 0.085000 ;
      RECT 1923.405000  1.785000 1923.575000 1.955000 ;
      RECT 1923.405000  2.635000 1923.575000 2.805000 ;
      RECT 1923.865000 -0.085000 1924.035000 0.085000 ;
      RECT 1923.865000  2.635000 1924.035000 2.805000 ;
      RECT 1924.325000 -0.085000 1924.495000 0.085000 ;
      RECT 1924.325000  2.635000 1924.495000 2.805000 ;
      RECT 1924.785000 -0.085000 1924.955000 0.085000 ;
      RECT 1924.785000  2.635000 1924.955000 2.805000 ;
      RECT 1925.245000 -0.085000 1925.415000 0.085000 ;
      RECT 1925.245000  2.635000 1925.415000 2.805000 ;
      RECT 1925.705000 -0.085000 1925.875000 0.085000 ;
      RECT 1925.705000  2.635000 1925.875000 2.805000 ;
      RECT 1926.165000 -0.085000 1926.335000 0.085000 ;
      RECT 1926.165000  2.635000 1926.335000 2.805000 ;
      RECT 1926.625000 -0.085000 1926.795000 0.085000 ;
      RECT 1926.625000  2.635000 1926.795000 2.805000 ;
      RECT 1927.085000 -0.085000 1927.255000 0.085000 ;
      RECT 1927.085000  2.635000 1927.255000 2.805000 ;
      RECT 1927.545000 -0.085000 1927.715000 0.085000 ;
      RECT 1927.545000  2.635000 1927.715000 2.805000 ;
      RECT 1928.005000 -0.085000 1928.175000 0.085000 ;
      RECT 1928.005000  2.635000 1928.175000 2.805000 ;
      RECT 1928.465000 -0.085000 1928.635000 0.085000 ;
      RECT 1928.465000  2.635000 1928.635000 2.805000 ;
      RECT 1928.925000 -0.085000 1929.095000 0.085000 ;
      RECT 1928.925000  2.635000 1929.095000 2.805000 ;
      RECT 1929.385000 -0.085000 1929.555000 0.085000 ;
      RECT 1929.385000  2.635000 1929.555000 2.805000 ;
      RECT 1929.845000 -0.085000 1930.015000 0.085000 ;
      RECT 1929.845000  2.635000 1930.015000 2.805000 ;
      RECT 1930.305000 -0.085000 1930.475000 0.085000 ;
      RECT 1930.305000  2.635000 1930.475000 2.805000 ;
      RECT 1930.765000 -0.085000 1930.935000 0.085000 ;
      RECT 1930.765000  2.635000 1930.935000 2.805000 ;
      RECT 1931.225000 -0.085000 1931.395000 0.085000 ;
      RECT 1931.225000  2.635000 1931.395000 2.805000 ;
      RECT 1931.685000 -0.085000 1931.855000 0.085000 ;
      RECT 1931.685000  2.635000 1931.855000 2.805000 ;
      RECT 1932.145000 -0.085000 1932.315000 0.085000 ;
      RECT 1932.145000  2.635000 1932.315000 2.805000 ;
      RECT 1932.605000 -0.085000 1932.775000 0.085000 ;
      RECT 1932.605000  2.635000 1932.775000 2.805000 ;
      RECT 1933.065000 -0.085000 1933.235000 0.085000 ;
      RECT 1933.065000  2.635000 1933.235000 2.805000 ;
      RECT 1933.525000 -0.085000 1933.695000 0.085000 ;
      RECT 1933.525000  2.635000 1933.695000 2.805000 ;
      RECT 1933.985000 -0.085000 1934.155000 0.085000 ;
      RECT 1933.985000  2.635000 1934.155000 2.805000 ;
      RECT 1934.445000 -0.085000 1934.615000 0.085000 ;
      RECT 1934.445000  2.635000 1934.615000 2.805000 ;
      RECT 1934.905000 -0.085000 1935.075000 0.085000 ;
      RECT 1934.905000  2.635000 1935.075000 2.805000 ;
      RECT 1935.365000 -0.085000 1935.535000 0.085000 ;
      RECT 1935.365000  2.635000 1935.535000 2.805000 ;
      RECT 1935.825000 -0.085000 1935.995000 0.085000 ;
      RECT 1935.825000  2.635000 1935.995000 2.805000 ;
      RECT 1936.285000 -0.085000 1936.455000 0.085000 ;
      RECT 1936.285000  2.635000 1936.455000 2.805000 ;
      RECT 1936.745000 -0.085000 1936.915000 0.085000 ;
      RECT 1936.745000  2.635000 1936.915000 2.805000 ;
      RECT 1937.205000 -0.085000 1937.375000 0.085000 ;
      RECT 1937.205000  2.635000 1937.375000 2.805000 ;
      RECT 1937.665000 -0.085000 1937.835000 0.085000 ;
      RECT 1937.665000  2.635000 1937.835000 2.805000 ;
      RECT 1938.125000 -0.085000 1938.295000 0.085000 ;
      RECT 1938.125000  2.635000 1938.295000 2.805000 ;
      RECT 1938.585000 -0.085000 1938.755000 0.085000 ;
      RECT 1938.585000  2.635000 1938.755000 2.805000 ;
      RECT 1939.045000 -0.085000 1939.215000 0.085000 ;
      RECT 1939.045000  2.635000 1939.215000 2.805000 ;
      RECT 1939.505000 -0.085000 1939.675000 0.085000 ;
      RECT 1939.505000  2.635000 1939.675000 2.805000 ;
      RECT 1939.965000 -0.085000 1940.135000 0.085000 ;
      RECT 1939.965000  2.635000 1940.135000 2.805000 ;
      RECT 1940.425000 -0.085000 1940.595000 0.085000 ;
      RECT 1940.425000  2.635000 1940.595000 2.805000 ;
      RECT 1940.885000 -0.085000 1941.055000 0.085000 ;
      RECT 1940.885000  2.635000 1941.055000 2.805000 ;
      RECT 1941.345000 -0.085000 1941.515000 0.085000 ;
      RECT 1941.345000  2.635000 1941.515000 2.805000 ;
      RECT 1941.805000 -0.085000 1941.975000 0.085000 ;
      RECT 1941.805000  2.635000 1941.975000 2.805000 ;
      RECT 1942.265000 -0.085000 1942.435000 0.085000 ;
      RECT 1942.265000  2.635000 1942.435000 2.805000 ;
      RECT 1942.265000  5.355000 1942.435000 5.525000 ;
      RECT 1942.725000 -0.085000 1942.895000 0.085000 ;
      RECT 1942.725000  2.635000 1942.895000 2.805000 ;
      RECT 1942.725000  5.355000 1942.895000 5.525000 ;
      RECT 1943.185000 -0.085000 1943.355000 0.085000 ;
      RECT 1943.185000  2.635000 1943.355000 2.805000 ;
      RECT 1943.185000  5.355000 1943.355000 5.525000 ;
      RECT 1943.645000 -0.085000 1943.815000 0.085000 ;
      RECT 1943.645000  2.635000 1943.815000 2.805000 ;
      RECT 1943.645000  5.355000 1943.815000 5.525000 ;
      RECT 1944.105000 -0.085000 1944.275000 0.085000 ;
      RECT 1944.105000  2.635000 1944.275000 2.805000 ;
      RECT 1944.105000  5.355000 1944.275000 5.525000 ;
      RECT 1944.385000  2.140000 1944.555000 2.310000 ;
      RECT 1944.385000  3.130000 1944.555000 3.300000 ;
      RECT 1944.565000 -0.085000 1944.735000 0.085000 ;
      RECT 1944.565000  5.355000 1944.735000 5.525000 ;
      RECT 1944.865000  1.785000 1945.035000 1.955000 ;
      RECT 1944.865000  3.485000 1945.035000 3.655000 ;
      RECT 1945.025000 -0.085000 1945.195000 0.085000 ;
      RECT 1945.025000  5.355000 1945.195000 5.525000 ;
      RECT 1945.335000  2.140000 1945.505000 2.310000 ;
      RECT 1945.335000  3.130000 1945.505000 3.300000 ;
      RECT 1945.485000 -0.085000 1945.655000 0.085000 ;
      RECT 1945.485000  5.355000 1945.655000 5.525000 ;
      RECT 1945.805000  1.785000 1945.975000 1.955000 ;
      RECT 1945.805000  3.485000 1945.975000 3.655000 ;
      RECT 1945.945000 -0.085000 1946.115000 0.085000 ;
      RECT 1945.945000  5.355000 1946.115000 5.525000 ;
      RECT 1946.285000  2.140000 1946.455000 2.310000 ;
      RECT 1946.285000  3.130000 1946.455000 3.300000 ;
      RECT 1946.405000 -0.085000 1946.575000 0.085000 ;
      RECT 1946.405000  2.635000 1946.575000 2.805000 ;
      RECT 1946.405000  5.355000 1946.575000 5.525000 ;
      RECT 1946.865000 -0.085000 1947.035000 0.085000 ;
      RECT 1946.865000  2.635000 1947.035000 2.805000 ;
      RECT 1946.865000  5.355000 1947.035000 5.525000 ;
      RECT 1947.265000  2.140000 1947.435000 2.310000 ;
      RECT 1947.265000  3.130000 1947.435000 3.300000 ;
      RECT 1947.325000 -0.085000 1947.495000 0.085000 ;
      RECT 1947.325000  2.635000 1947.495000 2.805000 ;
      RECT 1947.325000  5.355000 1947.495000 5.525000 ;
      RECT 1947.785000 -0.085000 1947.955000 0.085000 ;
      RECT 1947.785000  2.635000 1947.955000 2.805000 ;
      RECT 1947.785000  5.355000 1947.955000 5.525000 ;
      RECT 1948.205000  2.140000 1948.375000 2.310000 ;
      RECT 1948.205000  3.130000 1948.375000 3.300000 ;
      RECT 1948.245000 -0.085000 1948.415000 0.085000 ;
      RECT 1948.245000  2.635000 1948.415000 2.805000 ;
      RECT 1948.245000  5.355000 1948.415000 5.525000 ;
      RECT 1948.705000 -0.085000 1948.875000 0.085000 ;
      RECT 1948.705000  2.635000 1948.875000 2.805000 ;
      RECT 1948.705000  5.355000 1948.875000 5.525000 ;
      RECT 1949.165000 -0.085000 1949.335000 0.085000 ;
      RECT 1949.165000  2.635000 1949.335000 2.805000 ;
      RECT 1949.165000  5.355000 1949.335000 5.525000 ;
      RECT 1949.205000  2.140000 1949.375000 2.310000 ;
      RECT 1949.205000  3.130000 1949.375000 3.300000 ;
      RECT 1949.625000 -0.085000 1949.795000 0.085000 ;
      RECT 1949.625000  2.635000 1949.795000 2.805000 ;
      RECT 1949.625000  5.355000 1949.795000 5.525000 ;
      RECT 1950.085000 -0.085000 1950.255000 0.085000 ;
      RECT 1950.085000  2.635000 1950.255000 2.805000 ;
      RECT 1950.085000  5.355000 1950.255000 5.525000 ;
      RECT 1950.145000  2.140000 1950.315000 2.310000 ;
      RECT 1950.145000  3.130000 1950.315000 3.300000 ;
      RECT 1950.545000 -0.085000 1950.715000 0.085000 ;
      RECT 1950.545000  2.635000 1950.715000 2.805000 ;
      RECT 1950.545000  5.355000 1950.715000 5.525000 ;
      RECT 1951.005000 -0.085000 1951.175000 0.085000 ;
      RECT 1951.005000  2.635000 1951.175000 2.805000 ;
      RECT 1951.005000  5.355000 1951.175000 5.525000 ;
      RECT 1951.125000  2.140000 1951.295000 2.310000 ;
      RECT 1951.125000  3.130000 1951.295000 3.300000 ;
      RECT 1951.465000 -0.085000 1951.635000 0.085000 ;
      RECT 1951.465000  5.355000 1951.635000 5.525000 ;
      RECT 1951.605000  1.785000 1951.775000 1.955000 ;
      RECT 1951.605000  3.485000 1951.775000 3.655000 ;
      RECT 1951.925000 -0.085000 1952.095000 0.085000 ;
      RECT 1951.925000  5.355000 1952.095000 5.525000 ;
      RECT 1952.075000  2.140000 1952.245000 2.310000 ;
      RECT 1952.075000  3.130000 1952.245000 3.300000 ;
      RECT 1952.385000 -0.085000 1952.555000 0.085000 ;
      RECT 1952.385000  5.355000 1952.555000 5.525000 ;
      RECT 1952.545000  1.785000 1952.715000 1.955000 ;
      RECT 1952.545000  3.485000 1952.715000 3.655000 ;
      RECT 1952.845000 -0.085000 1953.015000 0.085000 ;
      RECT 1952.845000  5.355000 1953.015000 5.525000 ;
      RECT 1953.025000  2.140000 1953.195000 2.310000 ;
      RECT 1953.025000  3.130000 1953.195000 3.300000 ;
      RECT 1953.305000 -0.085000 1953.475000 0.085000 ;
      RECT 1953.305000  2.635000 1953.475000 2.805000 ;
      RECT 1953.305000  5.355000 1953.475000 5.525000 ;
      RECT 1953.765000 -0.085000 1953.935000 0.085000 ;
      RECT 1953.765000  2.635000 1953.935000 2.805000 ;
      RECT 1953.765000  5.355000 1953.935000 5.525000 ;
      RECT 1954.225000 -0.085000 1954.395000 0.085000 ;
      RECT 1954.225000  2.635000 1954.395000 2.805000 ;
      RECT 1954.225000  5.355000 1954.395000 5.525000 ;
      RECT 1954.685000 -0.085000 1954.855000 0.085000 ;
      RECT 1954.685000  2.635000 1954.855000 2.805000 ;
      RECT 1954.685000  5.355000 1954.855000 5.525000 ;
      RECT 1955.145000 -0.085000 1955.315000 0.085000 ;
      RECT 1955.145000  2.635000 1955.315000 2.805000 ;
      RECT 1955.145000  5.355000 1955.315000 5.525000 ;
      RECT 1955.605000 -0.085000 1955.775000 0.085000 ;
      RECT 1955.605000  2.635000 1955.775000 2.805000 ;
      RECT 1955.605000  5.355000 1955.775000 5.525000 ;
      RECT 1956.065000 -0.085000 1956.235000 0.085000 ;
      RECT 1956.065000  2.635000 1956.235000 2.805000 ;
      RECT 1956.065000  5.355000 1956.235000 5.525000 ;
      RECT 1956.525000 -0.085000 1956.695000 0.085000 ;
      RECT 1956.525000  2.635000 1956.695000 2.805000 ;
      RECT 1956.525000  5.355000 1956.695000 5.525000 ;
      RECT 1956.805000  2.140000 1956.975000 2.310000 ;
      RECT 1956.805000  3.130000 1956.975000 3.300000 ;
      RECT 1956.985000 -0.085000 1957.155000 0.085000 ;
      RECT 1956.985000  5.355000 1957.155000 5.525000 ;
      RECT 1957.285000  1.785000 1957.455000 1.955000 ;
      RECT 1957.285000  3.485000 1957.455000 3.655000 ;
      RECT 1957.445000 -0.085000 1957.615000 0.085000 ;
      RECT 1957.445000  5.355000 1957.615000 5.525000 ;
      RECT 1957.755000  2.140000 1957.925000 2.310000 ;
      RECT 1957.755000  3.130000 1957.925000 3.300000 ;
      RECT 1957.905000 -0.085000 1958.075000 0.085000 ;
      RECT 1957.905000  5.355000 1958.075000 5.525000 ;
      RECT 1958.225000  1.785000 1958.395000 1.955000 ;
      RECT 1958.225000  3.485000 1958.395000 3.655000 ;
      RECT 1958.365000 -0.085000 1958.535000 0.085000 ;
      RECT 1958.365000  5.355000 1958.535000 5.525000 ;
      RECT 1958.705000  2.140000 1958.875000 2.310000 ;
      RECT 1958.705000  3.130000 1958.875000 3.300000 ;
      RECT 1958.825000 -0.085000 1958.995000 0.085000 ;
      RECT 1958.825000  2.635000 1958.995000 2.805000 ;
      RECT 1958.825000  5.355000 1958.995000 5.525000 ;
      RECT 1959.285000 -0.085000 1959.455000 0.085000 ;
      RECT 1959.285000  2.635000 1959.455000 2.805000 ;
      RECT 1959.285000  5.355000 1959.455000 5.525000 ;
      RECT 1959.685000  2.140000 1959.855000 2.310000 ;
      RECT 1959.685000  3.130000 1959.855000 3.300000 ;
      RECT 1959.745000 -0.085000 1959.915000 0.085000 ;
      RECT 1959.745000  2.635000 1959.915000 2.805000 ;
      RECT 1959.745000  5.355000 1959.915000 5.525000 ;
      RECT 1960.205000 -0.085000 1960.375000 0.085000 ;
      RECT 1960.205000  2.635000 1960.375000 2.805000 ;
      RECT 1960.205000  5.355000 1960.375000 5.525000 ;
      RECT 1960.625000  2.140000 1960.795000 2.310000 ;
      RECT 1960.625000  3.130000 1960.795000 3.300000 ;
      RECT 1960.665000 -0.085000 1960.835000 0.085000 ;
      RECT 1960.665000  2.635000 1960.835000 2.805000 ;
      RECT 1960.665000  5.355000 1960.835000 5.525000 ;
      RECT 1961.125000 -0.085000 1961.295000 0.085000 ;
      RECT 1961.125000  2.635000 1961.295000 2.805000 ;
      RECT 1961.125000  5.355000 1961.295000 5.525000 ;
      RECT 1961.585000 -0.085000 1961.755000 0.085000 ;
      RECT 1961.585000  2.635000 1961.755000 2.805000 ;
      RECT 1961.585000  5.355000 1961.755000 5.525000 ;
      RECT 1961.625000  2.140000 1961.795000 2.310000 ;
      RECT 1961.625000  3.130000 1961.795000 3.300000 ;
      RECT 1962.045000 -0.085000 1962.215000 0.085000 ;
      RECT 1962.045000  2.635000 1962.215000 2.805000 ;
      RECT 1962.045000  5.355000 1962.215000 5.525000 ;
      RECT 1962.505000 -0.085000 1962.675000 0.085000 ;
      RECT 1962.505000  2.635000 1962.675000 2.805000 ;
      RECT 1962.505000  5.355000 1962.675000 5.525000 ;
      RECT 1962.565000  2.140000 1962.735000 2.310000 ;
      RECT 1962.565000  3.130000 1962.735000 3.300000 ;
      RECT 1962.965000 -0.085000 1963.135000 0.085000 ;
      RECT 1962.965000  2.635000 1963.135000 2.805000 ;
      RECT 1962.965000  5.355000 1963.135000 5.525000 ;
      RECT 1963.425000 -0.085000 1963.595000 0.085000 ;
      RECT 1963.425000  2.635000 1963.595000 2.805000 ;
      RECT 1963.425000  5.355000 1963.595000 5.525000 ;
      RECT 1963.545000  2.140000 1963.715000 2.310000 ;
      RECT 1963.545000  3.130000 1963.715000 3.300000 ;
      RECT 1963.885000 -0.085000 1964.055000 0.085000 ;
      RECT 1963.885000  5.355000 1964.055000 5.525000 ;
      RECT 1964.025000  1.785000 1964.195000 1.955000 ;
      RECT 1964.025000  3.485000 1964.195000 3.655000 ;
      RECT 1964.345000 -0.085000 1964.515000 0.085000 ;
      RECT 1964.345000  5.355000 1964.515000 5.525000 ;
      RECT 1964.495000  2.140000 1964.665000 2.310000 ;
      RECT 1964.495000  3.130000 1964.665000 3.300000 ;
      RECT 1964.805000 -0.085000 1964.975000 0.085000 ;
      RECT 1964.805000  5.355000 1964.975000 5.525000 ;
      RECT 1964.965000  1.785000 1965.135000 1.955000 ;
      RECT 1964.965000  3.485000 1965.135000 3.655000 ;
      RECT 1965.265000 -0.085000 1965.435000 0.085000 ;
      RECT 1965.265000  5.355000 1965.435000 5.525000 ;
      RECT 1965.445000  2.140000 1965.615000 2.310000 ;
      RECT 1965.445000  3.130000 1965.615000 3.300000 ;
      RECT 1965.725000 -0.085000 1965.895000 0.085000 ;
      RECT 1965.725000  2.635000 1965.895000 2.805000 ;
      RECT 1965.725000  5.355000 1965.895000 5.525000 ;
      RECT 1966.185000 -0.085000 1966.355000 0.085000 ;
      RECT 1966.185000  2.635000 1966.355000 2.805000 ;
      RECT 1966.185000  5.355000 1966.355000 5.525000 ;
      RECT 1966.645000 -0.085000 1966.815000 0.085000 ;
      RECT 1966.645000  2.635000 1966.815000 2.805000 ;
      RECT 1966.645000  5.355000 1966.815000 5.525000 ;
      RECT 1967.105000 -0.085000 1967.275000 0.085000 ;
      RECT 1967.105000  2.635000 1967.275000 2.805000 ;
      RECT 1967.105000  5.355000 1967.275000 5.525000 ;
      RECT 1967.565000 -0.085000 1967.735000 0.085000 ;
      RECT 1967.565000  2.635000 1967.735000 2.805000 ;
      RECT 1967.565000  5.355000 1967.735000 5.525000 ;
      RECT 1968.025000 -0.085000 1968.195000 0.085000 ;
      RECT 1968.025000  2.635000 1968.195000 2.805000 ;
      RECT 1968.025000  5.355000 1968.195000 5.525000 ;
      RECT 1968.485000 -0.085000 1968.655000 0.085000 ;
      RECT 1968.485000  2.635000 1968.655000 2.805000 ;
      RECT 1968.485000  5.355000 1968.655000 5.525000 ;
      RECT 1968.945000 -0.085000 1969.115000 0.085000 ;
      RECT 1968.945000  1.785000 1969.115000 1.955000 ;
      RECT 1968.945000  3.485000 1969.115000 3.655000 ;
      RECT 1968.945000  5.355000 1969.115000 5.525000 ;
      RECT 1969.405000 -0.085000 1969.575000 0.085000 ;
      RECT 1969.405000  2.635000 1969.575000 2.805000 ;
      RECT 1969.405000  5.355000 1969.575000 5.525000 ;
      RECT 1969.865000 -0.085000 1970.035000 0.085000 ;
      RECT 1969.865000  2.635000 1970.035000 2.805000 ;
      RECT 1969.865000  5.355000 1970.035000 5.525000 ;
      RECT 1970.325000 -0.085000 1970.495000 0.085000 ;
      RECT 1970.325000  2.635000 1970.495000 2.805000 ;
      RECT 1970.325000  5.355000 1970.495000 5.525000 ;
      RECT 1970.785000 -0.085000 1970.955000 0.085000 ;
      RECT 1970.785000  2.635000 1970.955000 2.805000 ;
      RECT 1970.785000  5.355000 1970.955000 5.525000 ;
      RECT 1971.245000 -0.085000 1971.415000 0.085000 ;
      RECT 1971.245000  1.785000 1971.415000 1.955000 ;
      RECT 1971.245000  3.485000 1971.415000 3.655000 ;
      RECT 1971.245000  5.355000 1971.415000 5.525000 ;
      RECT 1971.705000 -0.085000 1971.875000 0.085000 ;
      RECT 1971.705000  2.635000 1971.875000 2.805000 ;
      RECT 1971.705000  5.355000 1971.875000 5.525000 ;
      RECT 1972.165000 -0.085000 1972.335000 0.085000 ;
      RECT 1972.165000  2.635000 1972.335000 2.805000 ;
      RECT 1972.165000  5.355000 1972.335000 5.525000 ;
      RECT 1972.625000 -0.085000 1972.795000 0.085000 ;
      RECT 1972.625000  2.635000 1972.795000 2.805000 ;
      RECT 1972.625000  5.355000 1972.795000 5.525000 ;
      RECT 1973.085000 -0.085000 1973.255000 0.085000 ;
      RECT 1973.085000  1.785000 1973.255000 1.955000 ;
      RECT 1973.085000  3.485000 1973.255000 3.655000 ;
      RECT 1973.085000  5.355000 1973.255000 5.525000 ;
      RECT 1973.545000 -0.085000 1973.715000 0.085000 ;
      RECT 1973.545000  2.635000 1973.715000 2.805000 ;
      RECT 1973.545000  5.355000 1973.715000 5.525000 ;
      RECT 1974.005000 -0.085000 1974.175000 0.085000 ;
      RECT 1974.005000  2.635000 1974.175000 2.805000 ;
      RECT 1974.005000  5.355000 1974.175000 5.525000 ;
      RECT 1974.465000 -0.085000 1974.635000 0.085000 ;
      RECT 1974.465000  2.635000 1974.635000 2.805000 ;
      RECT 1974.465000  5.355000 1974.635000 5.525000 ;
      RECT 1974.925000 -0.085000 1975.095000 0.085000 ;
      RECT 1974.925000  2.635000 1975.095000 2.805000 ;
      RECT 1974.925000  5.355000 1975.095000 5.525000 ;
      RECT 1975.385000 -0.085000 1975.555000 0.085000 ;
      RECT 1975.385000  1.785000 1975.555000 1.955000 ;
      RECT 1975.385000  3.485000 1975.555000 3.655000 ;
      RECT 1975.385000  5.355000 1975.555000 5.525000 ;
      RECT 1975.845000 -0.085000 1976.015000 0.085000 ;
      RECT 1975.845000  2.635000 1976.015000 2.805000 ;
      RECT 1975.845000  5.355000 1976.015000 5.525000 ;
      RECT 1976.305000 -0.085000 1976.475000 0.085000 ;
      RECT 1976.305000  2.635000 1976.475000 2.805000 ;
      RECT 1976.305000  5.355000 1976.475000 5.525000 ;
      RECT 1976.765000 -0.085000 1976.935000 0.085000 ;
      RECT 1976.765000  2.635000 1976.935000 2.805000 ;
      RECT 1976.765000  5.355000 1976.935000 5.525000 ;
      RECT 1977.225000 -0.085000 1977.395000 0.085000 ;
      RECT 1977.225000  1.785000 1977.395000 1.955000 ;
      RECT 1977.225000  3.485000 1977.395000 3.655000 ;
      RECT 1977.225000  5.355000 1977.395000 5.525000 ;
      RECT 1977.685000 -0.085000 1977.855000 0.085000 ;
      RECT 1977.685000  2.635000 1977.855000 2.805000 ;
      RECT 1977.685000  5.355000 1977.855000 5.525000 ;
      RECT 1978.145000 -0.085000 1978.315000 0.085000 ;
      RECT 1978.145000  2.635000 1978.315000 2.805000 ;
      RECT 1978.145000  5.355000 1978.315000 5.525000 ;
      RECT 1978.605000 -0.085000 1978.775000 0.085000 ;
      RECT 1978.605000  2.635000 1978.775000 2.805000 ;
      RECT 1978.605000  5.355000 1978.775000 5.525000 ;
      RECT 1979.065000 -0.085000 1979.235000 0.085000 ;
      RECT 1979.065000  2.635000 1979.235000 2.805000 ;
      RECT 1979.065000  5.355000 1979.235000 5.525000 ;
      RECT 1979.525000 -0.085000 1979.695000 0.085000 ;
      RECT 1979.525000  1.785000 1979.695000 1.955000 ;
      RECT 1979.525000  3.485000 1979.695000 3.655000 ;
      RECT 1979.525000  5.355000 1979.695000 5.525000 ;
      RECT 1979.985000 -0.085000 1980.155000 0.085000 ;
      RECT 1979.985000  2.635000 1980.155000 2.805000 ;
      RECT 1979.985000  5.355000 1980.155000 5.525000 ;
      RECT 1980.445000 -0.085000 1980.615000 0.085000 ;
      RECT 1980.445000  2.635000 1980.615000 2.805000 ;
      RECT 1980.445000  5.355000 1980.615000 5.525000 ;
      RECT 1980.905000 -0.085000 1981.075000 0.085000 ;
      RECT 1980.905000  2.635000 1981.075000 2.805000 ;
      RECT 1980.905000  5.355000 1981.075000 5.525000 ;
      RECT 1981.365000 -0.085000 1981.535000 0.085000 ;
      RECT 1981.365000  1.785000 1981.535000 1.955000 ;
      RECT 1981.365000  3.485000 1981.535000 3.655000 ;
      RECT 1981.365000  5.355000 1981.535000 5.525000 ;
      RECT 1981.825000 -0.085000 1981.995000 0.085000 ;
      RECT 1981.825000  2.635000 1981.995000 2.805000 ;
      RECT 1981.825000  5.355000 1981.995000 5.525000 ;
      RECT 1982.285000 -0.085000 1982.455000 0.085000 ;
      RECT 1982.285000  2.635000 1982.455000 2.805000 ;
      RECT 1982.285000  5.355000 1982.455000 5.525000 ;
      RECT 1982.745000 -0.085000 1982.915000 0.085000 ;
      RECT 1982.745000  2.635000 1982.915000 2.805000 ;
      RECT 1982.745000  5.355000 1982.915000 5.525000 ;
      RECT 1983.205000 -0.085000 1983.375000 0.085000 ;
      RECT 1983.205000  2.635000 1983.375000 2.805000 ;
      RECT 1983.205000  5.355000 1983.375000 5.525000 ;
      RECT 1983.665000 -0.085000 1983.835000 0.085000 ;
      RECT 1983.665000  1.785000 1983.835000 1.955000 ;
      RECT 1983.665000  3.485000 1983.835000 3.655000 ;
      RECT 1983.665000  5.355000 1983.835000 5.525000 ;
      RECT 1984.125000 -0.085000 1984.295000 0.085000 ;
      RECT 1984.125000  2.635000 1984.295000 2.805000 ;
      RECT 1984.125000  5.355000 1984.295000 5.525000 ;
      RECT 1984.585000 -0.085000 1984.755000 0.085000 ;
      RECT 1984.585000  2.635000 1984.755000 2.805000 ;
      RECT 1984.585000  5.355000 1984.755000 5.525000 ;
      RECT 1985.045000 -0.085000 1985.215000 0.085000 ;
      RECT 1985.045000  2.635000 1985.215000 2.805000 ;
      RECT 1985.045000  5.355000 1985.215000 5.525000 ;
      RECT 1985.505000 -0.085000 1985.675000 0.085000 ;
      RECT 1985.505000  2.635000 1985.675000 2.805000 ;
      RECT 1985.505000  5.355000 1985.675000 5.525000 ;
      RECT 1985.535000  2.140000 1985.705000 2.310000 ;
      RECT 1985.535000  3.130000 1985.705000 3.300000 ;
      RECT 1985.965000 -0.085000 1986.135000 0.085000 ;
      RECT 1985.965000  2.635000 1986.135000 2.805000 ;
      RECT 1985.965000  5.355000 1986.135000 5.525000 ;
      RECT 1986.425000 -0.085000 1986.595000 0.085000 ;
      RECT 1986.425000  2.635000 1986.595000 2.805000 ;
      RECT 1986.425000  5.355000 1986.595000 5.525000 ;
      RECT 1986.475000  2.140000 1986.645000 2.310000 ;
      RECT 1986.475000  3.130000 1986.645000 3.300000 ;
      RECT 1986.885000 -0.085000 1987.055000 0.085000 ;
      RECT 1986.885000  1.785000 1987.055000 1.955000 ;
      RECT 1986.885000  3.485000 1987.055000 3.655000 ;
      RECT 1986.885000  5.355000 1987.055000 5.525000 ;
      RECT 1987.345000 -0.085000 1987.515000 0.085000 ;
      RECT 1987.345000  2.635000 1987.515000 2.805000 ;
      RECT 1987.345000  5.355000 1987.515000 5.525000 ;
      RECT 1987.470000  2.140000 1987.640000 2.310000 ;
      RECT 1987.470000  3.130000 1987.640000 3.300000 ;
      RECT 1987.805000 -0.085000 1987.975000 0.085000 ;
      RECT 1987.805000  2.635000 1987.975000 2.805000 ;
      RECT 1987.805000  5.355000 1987.975000 5.525000 ;
      RECT 1988.265000 -0.085000 1988.435000 0.085000 ;
      RECT 1988.265000  2.635000 1988.435000 2.805000 ;
      RECT 1988.265000  5.355000 1988.435000 5.525000 ;
      RECT 1988.725000 -0.085000 1988.895000 0.085000 ;
      RECT 1988.725000  2.635000 1988.895000 2.805000 ;
      RECT 1988.725000  5.355000 1988.895000 5.525000 ;
      RECT 1989.185000 -0.085000 1989.355000 0.085000 ;
      RECT 1989.185000  2.635000 1989.355000 2.805000 ;
      RECT 1989.185000  5.355000 1989.355000 5.525000 ;
      RECT 1989.520000  2.140000 1989.690000 2.310000 ;
      RECT 1989.520000  3.130000 1989.690000 3.300000 ;
      RECT 1989.645000 -0.085000 1989.815000 0.085000 ;
      RECT 1989.645000  2.635000 1989.815000 2.805000 ;
      RECT 1989.645000  5.355000 1989.815000 5.525000 ;
      RECT 1990.105000 -0.085000 1990.275000 0.085000 ;
      RECT 1990.105000  1.785000 1990.275000 1.955000 ;
      RECT 1990.105000  3.485000 1990.275000 3.655000 ;
      RECT 1990.105000  5.355000 1990.275000 5.525000 ;
      RECT 1990.515000  2.140000 1990.685000 2.310000 ;
      RECT 1990.515000  3.130000 1990.685000 3.300000 ;
      RECT 1990.565000 -0.085000 1990.735000 0.085000 ;
      RECT 1990.565000  2.635000 1990.735000 2.805000 ;
      RECT 1990.565000  5.355000 1990.735000 5.525000 ;
      RECT 1991.025000 -0.085000 1991.195000 0.085000 ;
      RECT 1991.025000  2.635000 1991.195000 2.805000 ;
      RECT 1991.025000  5.355000 1991.195000 5.525000 ;
      RECT 1991.455000  2.140000 1991.625000 2.310000 ;
      RECT 1991.455000  3.130000 1991.625000 3.300000 ;
      RECT 1991.485000 -0.085000 1991.655000 0.085000 ;
      RECT 1991.485000  2.635000 1991.655000 2.805000 ;
      RECT 1991.485000  5.355000 1991.655000 5.525000 ;
      RECT 1991.945000 -0.085000 1992.115000 0.085000 ;
      RECT 1991.945000  2.635000 1992.115000 2.805000 ;
      RECT 1991.945000  5.355000 1992.115000 5.525000 ;
      RECT 1991.975000  2.140000 1992.145000 2.310000 ;
      RECT 1991.975000  3.130000 1992.145000 3.300000 ;
      RECT 1992.405000 -0.085000 1992.575000 0.085000 ;
      RECT 1992.405000  2.635000 1992.575000 2.805000 ;
      RECT 1992.405000  5.355000 1992.575000 5.525000 ;
      RECT 1992.865000 -0.085000 1993.035000 0.085000 ;
      RECT 1992.865000  2.635000 1993.035000 2.805000 ;
      RECT 1992.865000  5.355000 1993.035000 5.525000 ;
      RECT 1992.915000  2.140000 1993.085000 2.310000 ;
      RECT 1992.915000  3.130000 1993.085000 3.300000 ;
      RECT 1993.325000 -0.085000 1993.495000 0.085000 ;
      RECT 1993.325000  1.785000 1993.495000 1.955000 ;
      RECT 1993.325000  3.485000 1993.495000 3.655000 ;
      RECT 1993.325000  5.355000 1993.495000 5.525000 ;
      RECT 1993.785000 -0.085000 1993.955000 0.085000 ;
      RECT 1993.785000  2.635000 1993.955000 2.805000 ;
      RECT 1993.785000  5.355000 1993.955000 5.525000 ;
      RECT 1993.910000  2.140000 1994.080000 2.310000 ;
      RECT 1993.910000  3.130000 1994.080000 3.300000 ;
      RECT 1994.245000 -0.085000 1994.415000 0.085000 ;
      RECT 1994.245000  2.635000 1994.415000 2.805000 ;
      RECT 1994.245000  5.355000 1994.415000 5.525000 ;
      RECT 1994.705000 -0.085000 1994.875000 0.085000 ;
      RECT 1994.705000  2.635000 1994.875000 2.805000 ;
      RECT 1994.705000  5.355000 1994.875000 5.525000 ;
      RECT 1995.165000 -0.085000 1995.335000 0.085000 ;
      RECT 1995.165000  2.635000 1995.335000 2.805000 ;
      RECT 1995.165000  5.355000 1995.335000 5.525000 ;
      RECT 1995.625000 -0.085000 1995.795000 0.085000 ;
      RECT 1995.625000  2.635000 1995.795000 2.805000 ;
      RECT 1995.625000  5.355000 1995.795000 5.525000 ;
      RECT 1995.960000  2.140000 1996.130000 2.310000 ;
      RECT 1995.960000  3.130000 1996.130000 3.300000 ;
      RECT 1996.085000 -0.085000 1996.255000 0.085000 ;
      RECT 1996.085000  2.635000 1996.255000 2.805000 ;
      RECT 1996.085000  5.355000 1996.255000 5.525000 ;
      RECT 1996.545000 -0.085000 1996.715000 0.085000 ;
      RECT 1996.545000  1.785000 1996.715000 1.955000 ;
      RECT 1996.545000  3.485000 1996.715000 3.655000 ;
      RECT 1996.545000  5.355000 1996.715000 5.525000 ;
      RECT 1996.955000  2.140000 1997.125000 2.310000 ;
      RECT 1996.955000  3.130000 1997.125000 3.300000 ;
      RECT 1997.005000 -0.085000 1997.175000 0.085000 ;
      RECT 1997.005000  2.635000 1997.175000 2.805000 ;
      RECT 1997.005000  5.355000 1997.175000 5.525000 ;
      RECT 1997.465000 -0.085000 1997.635000 0.085000 ;
      RECT 1997.465000  2.635000 1997.635000 2.805000 ;
      RECT 1997.465000  5.355000 1997.635000 5.525000 ;
      RECT 1997.895000  2.140000 1998.065000 2.310000 ;
      RECT 1997.895000  3.130000 1998.065000 3.300000 ;
      RECT 1997.925000 -0.085000 1998.095000 0.085000 ;
      RECT 1997.925000  2.635000 1998.095000 2.805000 ;
      RECT 1997.925000  5.355000 1998.095000 5.525000 ;
      RECT 1998.385000 -0.085000 1998.555000 0.085000 ;
      RECT 1998.385000  2.635000 1998.555000 2.805000 ;
      RECT 1998.385000  5.355000 1998.555000 5.525000 ;
      RECT 1998.415000  2.140000 1998.585000 2.310000 ;
      RECT 1998.415000  3.130000 1998.585000 3.300000 ;
      RECT 1998.845000 -0.085000 1999.015000 0.085000 ;
      RECT 1998.845000  2.635000 1999.015000 2.805000 ;
      RECT 1998.845000  5.355000 1999.015000 5.525000 ;
      RECT 1999.305000 -0.085000 1999.475000 0.085000 ;
      RECT 1999.305000  2.635000 1999.475000 2.805000 ;
      RECT 1999.305000  5.355000 1999.475000 5.525000 ;
      RECT 1999.355000  2.140000 1999.525000 2.310000 ;
      RECT 1999.355000  3.130000 1999.525000 3.300000 ;
      RECT 1999.765000 -0.085000 1999.935000 0.085000 ;
      RECT 1999.765000  1.785000 1999.935000 1.955000 ;
      RECT 1999.765000  3.485000 1999.935000 3.655000 ;
      RECT 1999.765000  5.355000 1999.935000 5.525000 ;
      RECT 2000.225000 -0.085000 2000.395000 0.085000 ;
      RECT 2000.225000  2.635000 2000.395000 2.805000 ;
      RECT 2000.225000  5.355000 2000.395000 5.525000 ;
      RECT 2000.350000  2.140000 2000.520000 2.310000 ;
      RECT 2000.350000  3.130000 2000.520000 3.300000 ;
      RECT 2000.685000 -0.085000 2000.855000 0.085000 ;
      RECT 2000.685000  2.635000 2000.855000 2.805000 ;
      RECT 2000.685000  5.355000 2000.855000 5.525000 ;
      RECT 2001.145000 -0.085000 2001.315000 0.085000 ;
      RECT 2001.145000  2.635000 2001.315000 2.805000 ;
      RECT 2001.145000  5.355000 2001.315000 5.525000 ;
      RECT 2001.605000 -0.085000 2001.775000 0.085000 ;
      RECT 2001.605000  2.635000 2001.775000 2.805000 ;
      RECT 2001.605000  5.355000 2001.775000 5.525000 ;
      RECT 2002.065000 -0.085000 2002.235000 0.085000 ;
      RECT 2002.065000  2.635000 2002.235000 2.805000 ;
      RECT 2002.065000  5.355000 2002.235000 5.525000 ;
      RECT 2002.400000  2.140000 2002.570000 2.310000 ;
      RECT 2002.400000  3.130000 2002.570000 3.300000 ;
      RECT 2002.525000 -0.085000 2002.695000 0.085000 ;
      RECT 2002.525000  2.635000 2002.695000 2.805000 ;
      RECT 2002.525000  5.355000 2002.695000 5.525000 ;
      RECT 2002.985000 -0.085000 2003.155000 0.085000 ;
      RECT 2002.985000  1.785000 2003.155000 1.955000 ;
      RECT 2002.985000  3.485000 2003.155000 3.655000 ;
      RECT 2002.985000  5.355000 2003.155000 5.525000 ;
      RECT 2003.395000  2.140000 2003.565000 2.310000 ;
      RECT 2003.395000  3.130000 2003.565000 3.300000 ;
      RECT 2003.445000 -0.085000 2003.615000 0.085000 ;
      RECT 2003.445000  2.635000 2003.615000 2.805000 ;
      RECT 2003.445000  5.355000 2003.615000 5.525000 ;
      RECT 2003.905000 -0.085000 2004.075000 0.085000 ;
      RECT 2003.905000  2.635000 2004.075000 2.805000 ;
      RECT 2003.905000  5.355000 2004.075000 5.525000 ;
      RECT 2004.335000  2.140000 2004.505000 2.310000 ;
      RECT 2004.335000  3.130000 2004.505000 3.300000 ;
      RECT 2004.365000 -0.085000 2004.535000 0.085000 ;
      RECT 2004.365000  2.635000 2004.535000 2.805000 ;
      RECT 2004.365000  5.355000 2004.535000 5.525000 ;
      RECT 2004.825000 -0.085000 2004.995000 0.085000 ;
      RECT 2004.825000  2.635000 2004.995000 2.805000 ;
      RECT 2004.825000  5.355000 2004.995000 5.525000 ;
      RECT 2004.855000  2.140000 2005.025000 2.310000 ;
      RECT 2004.855000  3.130000 2005.025000 3.300000 ;
      RECT 2005.285000 -0.085000 2005.455000 0.085000 ;
      RECT 2005.285000  2.635000 2005.455000 2.805000 ;
      RECT 2005.285000  5.355000 2005.455000 5.525000 ;
      RECT 2005.745000 -0.085000 2005.915000 0.085000 ;
      RECT 2005.745000  2.635000 2005.915000 2.805000 ;
      RECT 2005.745000  5.355000 2005.915000 5.525000 ;
      RECT 2005.795000  2.140000 2005.965000 2.310000 ;
      RECT 2005.795000  3.130000 2005.965000 3.300000 ;
      RECT 2006.205000 -0.085000 2006.375000 0.085000 ;
      RECT 2006.205000  1.785000 2006.375000 1.955000 ;
      RECT 2006.205000  3.485000 2006.375000 3.655000 ;
      RECT 2006.205000  5.355000 2006.375000 5.525000 ;
      RECT 2006.665000 -0.085000 2006.835000 0.085000 ;
      RECT 2006.665000  2.635000 2006.835000 2.805000 ;
      RECT 2006.665000  5.355000 2006.835000 5.525000 ;
      RECT 2006.790000  2.140000 2006.960000 2.310000 ;
      RECT 2006.790000  3.130000 2006.960000 3.300000 ;
      RECT 2007.125000 -0.085000 2007.295000 0.085000 ;
      RECT 2007.125000  2.635000 2007.295000 2.805000 ;
      RECT 2007.125000  5.355000 2007.295000 5.525000 ;
      RECT 2007.585000 -0.085000 2007.755000 0.085000 ;
      RECT 2007.585000  2.635000 2007.755000 2.805000 ;
      RECT 2007.585000  5.355000 2007.755000 5.525000 ;
      RECT 2008.045000 -0.085000 2008.215000 0.085000 ;
      RECT 2008.045000  2.635000 2008.215000 2.805000 ;
      RECT 2008.045000  5.355000 2008.215000 5.525000 ;
      RECT 2008.505000 -0.085000 2008.675000 0.085000 ;
      RECT 2008.505000  2.635000 2008.675000 2.805000 ;
      RECT 2008.505000  5.355000 2008.675000 5.525000 ;
      RECT 2008.840000  2.140000 2009.010000 2.310000 ;
      RECT 2008.840000  3.130000 2009.010000 3.300000 ;
      RECT 2008.965000 -0.085000 2009.135000 0.085000 ;
      RECT 2008.965000  2.635000 2009.135000 2.805000 ;
      RECT 2008.965000  5.355000 2009.135000 5.525000 ;
      RECT 2009.425000 -0.085000 2009.595000 0.085000 ;
      RECT 2009.425000  1.785000 2009.595000 1.955000 ;
      RECT 2009.425000  3.485000 2009.595000 3.655000 ;
      RECT 2009.425000  5.355000 2009.595000 5.525000 ;
      RECT 2009.835000  2.140000 2010.005000 2.310000 ;
      RECT 2009.835000  3.130000 2010.005000 3.300000 ;
      RECT 2009.885000 -0.085000 2010.055000 0.085000 ;
      RECT 2009.885000  2.635000 2010.055000 2.805000 ;
      RECT 2009.885000  5.355000 2010.055000 5.525000 ;
      RECT 2010.345000 -0.085000 2010.515000 0.085000 ;
      RECT 2010.345000  2.635000 2010.515000 2.805000 ;
      RECT 2010.345000  5.355000 2010.515000 5.525000 ;
      RECT 2010.775000  2.140000 2010.945000 2.310000 ;
      RECT 2010.775000  3.130000 2010.945000 3.300000 ;
      RECT 2010.805000 -0.085000 2010.975000 0.085000 ;
      RECT 2010.805000  2.635000 2010.975000 2.805000 ;
      RECT 2010.805000  5.355000 2010.975000 5.525000 ;
      RECT 2011.265000 -0.085000 2011.435000 0.085000 ;
      RECT 2011.265000  2.635000 2011.435000 2.805000 ;
      RECT 2011.265000  5.355000 2011.435000 5.525000 ;
      RECT 2011.725000 -0.085000 2011.895000 0.085000 ;
      RECT 2011.725000  2.635000 2011.895000 2.805000 ;
      RECT 2011.725000  5.355000 2011.895000 5.525000 ;
      RECT 2012.185000 -0.085000 2012.355000 0.085000 ;
      RECT 2012.185000  2.635000 2012.355000 2.805000 ;
      RECT 2012.185000  5.355000 2012.355000 5.525000 ;
      RECT 2012.225000  2.140000 2012.395000 2.310000 ;
      RECT 2012.225000  3.130000 2012.395000 3.300000 ;
      RECT 2012.645000 -0.085000 2012.815000 0.085000 ;
      RECT 2012.645000  2.635000 2012.815000 2.805000 ;
      RECT 2012.645000  5.355000 2012.815000 5.525000 ;
      RECT 2013.105000 -0.085000 2013.275000 0.085000 ;
      RECT 2013.105000  2.635000 2013.275000 2.805000 ;
      RECT 2013.105000  5.355000 2013.275000 5.525000 ;
      RECT 2013.165000  2.140000 2013.335000 2.310000 ;
      RECT 2013.165000  3.130000 2013.335000 3.300000 ;
      RECT 2013.565000 -0.085000 2013.735000 0.085000 ;
      RECT 2013.565000  2.635000 2013.735000 2.805000 ;
      RECT 2013.565000  5.355000 2013.735000 5.525000 ;
      RECT 2014.025000 -0.085000 2014.195000 0.085000 ;
      RECT 2014.025000  2.635000 2014.195000 2.805000 ;
      RECT 2014.025000  5.355000 2014.195000 5.525000 ;
      RECT 2014.145000  2.140000 2014.315000 2.310000 ;
      RECT 2014.145000  3.130000 2014.315000 3.300000 ;
      RECT 2014.485000 -0.085000 2014.655000 0.085000 ;
      RECT 2014.485000  5.355000 2014.655000 5.525000 ;
      RECT 2014.625000  1.785000 2014.795000 1.955000 ;
      RECT 2014.625000  3.485000 2014.795000 3.655000 ;
      RECT 2014.945000 -0.085000 2015.115000 0.085000 ;
      RECT 2014.945000  5.355000 2015.115000 5.525000 ;
      RECT 2015.095000  2.140000 2015.265000 2.310000 ;
      RECT 2015.095000  3.130000 2015.265000 3.300000 ;
      RECT 2015.405000 -0.085000 2015.575000 0.085000 ;
      RECT 2015.405000  5.355000 2015.575000 5.525000 ;
      RECT 2015.565000  1.785000 2015.735000 1.955000 ;
      RECT 2015.565000  3.485000 2015.735000 3.655000 ;
      RECT 2015.865000 -0.085000 2016.035000 0.085000 ;
      RECT 2015.865000  5.355000 2016.035000 5.525000 ;
      RECT 2016.045000  2.140000 2016.215000 2.310000 ;
      RECT 2016.045000  3.130000 2016.215000 3.300000 ;
      RECT 2016.325000 -0.085000 2016.495000 0.085000 ;
      RECT 2016.325000  2.635000 2016.495000 2.805000 ;
      RECT 2016.325000  5.355000 2016.495000 5.525000 ;
      RECT 2016.785000 -0.085000 2016.955000 0.085000 ;
      RECT 2016.785000  2.635000 2016.955000 2.805000 ;
      RECT 2016.785000  5.355000 2016.955000 5.525000 ;
      RECT 2017.245000 -0.085000 2017.415000 0.085000 ;
      RECT 2017.245000  2.635000 2017.415000 2.805000 ;
      RECT 2017.245000  5.355000 2017.415000 5.525000 ;
      RECT 2017.705000 -0.085000 2017.875000 0.085000 ;
      RECT 2017.705000  2.635000 2017.875000 2.805000 ;
      RECT 2017.705000  5.355000 2017.875000 5.525000 ;
      RECT 2018.165000 -0.085000 2018.335000 0.085000 ;
      RECT 2018.165000  2.635000 2018.335000 2.805000 ;
      RECT 2018.165000  5.355000 2018.335000 5.525000 ;
      RECT 2018.625000 -0.085000 2018.795000 0.085000 ;
      RECT 2018.625000  2.635000 2018.795000 2.805000 ;
      RECT 2018.625000  5.355000 2018.795000 5.525000 ;
      RECT 2019.085000 -0.085000 2019.255000 0.085000 ;
      RECT 2019.085000  2.635000 2019.255000 2.805000 ;
      RECT 2019.085000  5.355000 2019.255000 5.525000 ;
      RECT 2019.545000 -0.085000 2019.715000 0.085000 ;
      RECT 2019.545000  2.635000 2019.715000 2.805000 ;
      RECT 2019.545000  5.355000 2019.715000 5.525000 ;
      RECT 2019.825000  2.140000 2019.995000 2.310000 ;
      RECT 2019.825000  3.130000 2019.995000 3.300000 ;
      RECT 2020.005000 -0.085000 2020.175000 0.085000 ;
      RECT 2020.005000  5.355000 2020.175000 5.525000 ;
      RECT 2020.305000  1.785000 2020.475000 1.955000 ;
      RECT 2020.305000  3.485000 2020.475000 3.655000 ;
      RECT 2020.465000 -0.085000 2020.635000 0.085000 ;
      RECT 2020.465000  5.355000 2020.635000 5.525000 ;
      RECT 2020.775000  2.140000 2020.945000 2.310000 ;
      RECT 2020.775000  3.130000 2020.945000 3.300000 ;
      RECT 2020.925000 -0.085000 2021.095000 0.085000 ;
      RECT 2020.925000  5.355000 2021.095000 5.525000 ;
      RECT 2021.245000  1.785000 2021.415000 1.955000 ;
      RECT 2021.245000  3.485000 2021.415000 3.655000 ;
      RECT 2021.385000 -0.085000 2021.555000 0.085000 ;
      RECT 2021.385000  5.355000 2021.555000 5.525000 ;
      RECT 2021.725000  2.140000 2021.895000 2.310000 ;
      RECT 2021.725000  3.130000 2021.895000 3.300000 ;
      RECT 2021.845000 -0.085000 2022.015000 0.085000 ;
      RECT 2021.845000  2.635000 2022.015000 2.805000 ;
      RECT 2021.845000  5.355000 2022.015000 5.525000 ;
      RECT 2022.305000 -0.085000 2022.475000 0.085000 ;
      RECT 2022.305000  2.635000 2022.475000 2.805000 ;
      RECT 2022.305000  5.355000 2022.475000 5.525000 ;
      RECT 2022.705000  2.140000 2022.875000 2.310000 ;
      RECT 2022.705000  3.130000 2022.875000 3.300000 ;
      RECT 2022.765000 -0.085000 2022.935000 0.085000 ;
      RECT 2022.765000  2.635000 2022.935000 2.805000 ;
      RECT 2022.765000  5.355000 2022.935000 5.525000 ;
      RECT 2023.225000 -0.085000 2023.395000 0.085000 ;
      RECT 2023.225000  2.635000 2023.395000 2.805000 ;
      RECT 2023.225000  5.355000 2023.395000 5.525000 ;
      RECT 2023.645000  2.140000 2023.815000 2.310000 ;
      RECT 2023.645000  3.130000 2023.815000 3.300000 ;
      RECT 2023.685000 -0.085000 2023.855000 0.085000 ;
      RECT 2023.685000  2.635000 2023.855000 2.805000 ;
      RECT 2023.685000  5.355000 2023.855000 5.525000 ;
      RECT 2024.145000 -0.085000 2024.315000 0.085000 ;
      RECT 2024.145000  2.635000 2024.315000 2.805000 ;
      RECT 2024.145000  5.355000 2024.315000 5.525000 ;
      RECT 2024.605000 -0.085000 2024.775000 0.085000 ;
      RECT 2024.605000  2.635000 2024.775000 2.805000 ;
      RECT 2024.605000  5.355000 2024.775000 5.525000 ;
      RECT 2025.065000 -0.085000 2025.235000 0.085000 ;
      RECT 2025.065000  2.635000 2025.235000 2.805000 ;
      RECT 2025.065000  5.355000 2025.235000 5.525000 ;
      RECT 2025.105000  2.140000 2025.275000 2.310000 ;
      RECT 2025.105000  3.130000 2025.275000 3.300000 ;
      RECT 2025.525000 -0.085000 2025.695000 0.085000 ;
      RECT 2025.525000  2.635000 2025.695000 2.805000 ;
      RECT 2025.525000  5.355000 2025.695000 5.525000 ;
      RECT 2025.985000 -0.085000 2026.155000 0.085000 ;
      RECT 2025.985000  2.635000 2026.155000 2.805000 ;
      RECT 2025.985000  5.355000 2026.155000 5.525000 ;
      RECT 2026.045000  2.140000 2026.215000 2.310000 ;
      RECT 2026.045000  3.130000 2026.215000 3.300000 ;
      RECT 2026.445000 -0.085000 2026.615000 0.085000 ;
      RECT 2026.445000  2.635000 2026.615000 2.805000 ;
      RECT 2026.445000  5.355000 2026.615000 5.525000 ;
      RECT 2026.905000 -0.085000 2027.075000 0.085000 ;
      RECT 2026.905000  2.635000 2027.075000 2.805000 ;
      RECT 2026.905000  5.355000 2027.075000 5.525000 ;
      RECT 2027.025000  2.140000 2027.195000 2.310000 ;
      RECT 2027.025000  3.130000 2027.195000 3.300000 ;
      RECT 2027.365000 -0.085000 2027.535000 0.085000 ;
      RECT 2027.365000  5.355000 2027.535000 5.525000 ;
      RECT 2027.505000  1.785000 2027.675000 1.955000 ;
      RECT 2027.505000  3.485000 2027.675000 3.655000 ;
      RECT 2027.825000 -0.085000 2027.995000 0.085000 ;
      RECT 2027.825000  5.355000 2027.995000 5.525000 ;
      RECT 2027.975000  2.140000 2028.145000 2.310000 ;
      RECT 2027.975000  3.130000 2028.145000 3.300000 ;
      RECT 2028.285000 -0.085000 2028.455000 0.085000 ;
      RECT 2028.285000  5.355000 2028.455000 5.525000 ;
      RECT 2028.445000  1.785000 2028.615000 1.955000 ;
      RECT 2028.445000  3.485000 2028.615000 3.655000 ;
      RECT 2028.745000 -0.085000 2028.915000 0.085000 ;
      RECT 2028.745000  5.355000 2028.915000 5.525000 ;
      RECT 2028.925000  2.140000 2029.095000 2.310000 ;
      RECT 2028.925000  3.130000 2029.095000 3.300000 ;
      RECT 2029.205000 -0.085000 2029.375000 0.085000 ;
      RECT 2029.205000  2.635000 2029.375000 2.805000 ;
      RECT 2029.205000  5.355000 2029.375000 5.525000 ;
      RECT 2029.665000 -0.085000 2029.835000 0.085000 ;
      RECT 2029.665000  2.635000 2029.835000 2.805000 ;
      RECT 2029.665000  5.355000 2029.835000 5.525000 ;
      RECT 2030.125000 -0.085000 2030.295000 0.085000 ;
      RECT 2030.125000  2.635000 2030.295000 2.805000 ;
      RECT 2030.125000  5.355000 2030.295000 5.525000 ;
      RECT 2030.585000 -0.085000 2030.755000 0.085000 ;
      RECT 2030.585000  2.635000 2030.755000 2.805000 ;
      RECT 2030.585000  5.355000 2030.755000 5.525000 ;
      RECT 2031.045000 -0.085000 2031.215000 0.085000 ;
      RECT 2031.045000  2.635000 2031.215000 2.805000 ;
      RECT 2031.045000  5.355000 2031.215000 5.525000 ;
      RECT 2031.505000 -0.085000 2031.675000 0.085000 ;
      RECT 2031.505000  2.635000 2031.675000 2.805000 ;
      RECT 2031.505000  5.355000 2031.675000 5.525000 ;
      RECT 2031.965000 -0.085000 2032.135000 0.085000 ;
      RECT 2031.965000  2.635000 2032.135000 2.805000 ;
      RECT 2031.965000  5.355000 2032.135000 5.525000 ;
      RECT 2032.425000 -0.085000 2032.595000 0.085000 ;
      RECT 2032.425000  2.635000 2032.595000 2.805000 ;
      RECT 2032.425000  5.355000 2032.595000 5.525000 ;
      RECT 2032.705000  2.140000 2032.875000 2.310000 ;
      RECT 2032.705000  3.130000 2032.875000 3.300000 ;
      RECT 2032.885000 -0.085000 2033.055000 0.085000 ;
      RECT 2032.885000  5.355000 2033.055000 5.525000 ;
      RECT 2033.185000  1.785000 2033.355000 1.955000 ;
      RECT 2033.185000  3.485000 2033.355000 3.655000 ;
      RECT 2033.345000 -0.085000 2033.515000 0.085000 ;
      RECT 2033.345000  5.355000 2033.515000 5.525000 ;
      RECT 2033.655000  2.140000 2033.825000 2.310000 ;
      RECT 2033.655000  3.130000 2033.825000 3.300000 ;
      RECT 2033.805000 -0.085000 2033.975000 0.085000 ;
      RECT 2033.805000  5.355000 2033.975000 5.525000 ;
      RECT 2034.125000  1.785000 2034.295000 1.955000 ;
      RECT 2034.125000  3.485000 2034.295000 3.655000 ;
      RECT 2034.265000 -0.085000 2034.435000 0.085000 ;
      RECT 2034.265000  5.355000 2034.435000 5.525000 ;
      RECT 2034.605000  2.140000 2034.775000 2.310000 ;
      RECT 2034.605000  3.130000 2034.775000 3.300000 ;
      RECT 2034.725000 -0.085000 2034.895000 0.085000 ;
      RECT 2034.725000  2.635000 2034.895000 2.805000 ;
      RECT 2034.725000  5.355000 2034.895000 5.525000 ;
      RECT 2035.185000 -0.085000 2035.355000 0.085000 ;
      RECT 2035.185000  2.635000 2035.355000 2.805000 ;
      RECT 2035.185000  5.355000 2035.355000 5.525000 ;
      RECT 2035.585000  2.140000 2035.755000 2.310000 ;
      RECT 2035.585000  3.130000 2035.755000 3.300000 ;
      RECT 2035.645000 -0.085000 2035.815000 0.085000 ;
      RECT 2035.645000  2.635000 2035.815000 2.805000 ;
      RECT 2035.645000  5.355000 2035.815000 5.525000 ;
      RECT 2036.105000 -0.085000 2036.275000 0.085000 ;
      RECT 2036.105000  2.635000 2036.275000 2.805000 ;
      RECT 2036.105000  5.355000 2036.275000 5.525000 ;
      RECT 2036.525000  2.140000 2036.695000 2.310000 ;
      RECT 2036.525000  3.130000 2036.695000 3.300000 ;
      RECT 2036.565000 -0.085000 2036.735000 0.085000 ;
      RECT 2036.565000  2.635000 2036.735000 2.805000 ;
      RECT 2036.565000  5.355000 2036.735000 5.525000 ;
      RECT 2037.025000 -0.085000 2037.195000 0.085000 ;
      RECT 2037.025000  2.635000 2037.195000 2.805000 ;
      RECT 2037.025000  5.355000 2037.195000 5.525000 ;
      RECT 2037.485000 -0.085000 2037.655000 0.085000 ;
      RECT 2037.485000  2.635000 2037.655000 2.805000 ;
      RECT 2037.485000  5.355000 2037.655000 5.525000 ;
      RECT 2037.945000 -0.085000 2038.115000 0.085000 ;
      RECT 2037.945000  2.635000 2038.115000 2.805000 ;
      RECT 2037.945000  5.355000 2038.115000 5.525000 ;
      RECT 2038.405000 -0.085000 2038.575000 0.085000 ;
      RECT 2038.405000  2.635000 2038.575000 2.805000 ;
      RECT 2038.405000  5.355000 2038.575000 5.525000 ;
      RECT 2038.445000  2.140000 2038.615000 2.310000 ;
      RECT 2038.445000  3.130000 2038.615000 3.300000 ;
      RECT 2038.865000 -0.085000 2039.035000 0.085000 ;
      RECT 2038.865000  2.635000 2039.035000 2.805000 ;
      RECT 2038.865000  5.355000 2039.035000 5.525000 ;
      RECT 2039.325000 -0.085000 2039.495000 0.085000 ;
      RECT 2039.325000  2.635000 2039.495000 2.805000 ;
      RECT 2039.325000  5.355000 2039.495000 5.525000 ;
      RECT 2039.385000  2.140000 2039.555000 2.310000 ;
      RECT 2039.385000  3.130000 2039.555000 3.300000 ;
      RECT 2039.785000 -0.085000 2039.955000 0.085000 ;
      RECT 2039.785000  2.635000 2039.955000 2.805000 ;
      RECT 2039.785000  5.355000 2039.955000 5.525000 ;
      RECT 2040.245000 -0.085000 2040.415000 0.085000 ;
      RECT 2040.245000  2.635000 2040.415000 2.805000 ;
      RECT 2040.245000  5.355000 2040.415000 5.525000 ;
      RECT 2040.365000  2.140000 2040.535000 2.310000 ;
      RECT 2040.365000  3.130000 2040.535000 3.300000 ;
      RECT 2040.705000 -0.085000 2040.875000 0.085000 ;
      RECT 2040.705000  5.355000 2040.875000 5.525000 ;
      RECT 2040.845000  1.785000 2041.015000 1.955000 ;
      RECT 2040.845000  3.485000 2041.015000 3.655000 ;
      RECT 2041.165000 -0.085000 2041.335000 0.085000 ;
      RECT 2041.165000  5.355000 2041.335000 5.525000 ;
      RECT 2041.315000  2.140000 2041.485000 2.310000 ;
      RECT 2041.315000  3.130000 2041.485000 3.300000 ;
      RECT 2041.625000 -0.085000 2041.795000 0.085000 ;
      RECT 2041.625000  5.355000 2041.795000 5.525000 ;
      RECT 2041.785000  1.785000 2041.955000 1.955000 ;
      RECT 2041.785000  3.485000 2041.955000 3.655000 ;
      RECT 2042.085000 -0.085000 2042.255000 0.085000 ;
      RECT 2042.085000  5.355000 2042.255000 5.525000 ;
      RECT 2042.265000  2.140000 2042.435000 2.310000 ;
      RECT 2042.265000  3.130000 2042.435000 3.300000 ;
      RECT 2042.545000 -0.085000 2042.715000 0.085000 ;
      RECT 2042.545000  2.635000 2042.715000 2.805000 ;
      RECT 2042.545000  5.355000 2042.715000 5.525000 ;
      RECT 2043.005000 -0.085000 2043.175000 0.085000 ;
      RECT 2043.005000  2.635000 2043.175000 2.805000 ;
      RECT 2043.005000  5.355000 2043.175000 5.525000 ;
      RECT 2043.465000 -0.085000 2043.635000 0.085000 ;
      RECT 2043.465000  2.635000 2043.635000 2.805000 ;
      RECT 2043.465000  5.355000 2043.635000 5.525000 ;
      RECT 2043.925000 -0.085000 2044.095000 0.085000 ;
      RECT 2043.925000  2.635000 2044.095000 2.805000 ;
      RECT 2043.925000  5.355000 2044.095000 5.525000 ;
      RECT 2044.385000 -0.085000 2044.555000 0.085000 ;
      RECT 2044.385000  2.635000 2044.555000 2.805000 ;
      RECT 2044.385000  5.355000 2044.555000 5.525000 ;
      RECT 2044.845000 -0.085000 2045.015000 0.085000 ;
      RECT 2044.845000  2.635000 2045.015000 2.805000 ;
      RECT 2044.845000  5.355000 2045.015000 5.525000 ;
      RECT 2045.305000 -0.085000 2045.475000 0.085000 ;
      RECT 2045.305000  2.635000 2045.475000 2.805000 ;
      RECT 2045.305000  5.355000 2045.475000 5.525000 ;
      RECT 2045.765000 -0.085000 2045.935000 0.085000 ;
      RECT 2045.765000  2.635000 2045.935000 2.805000 ;
      RECT 2045.765000  5.355000 2045.935000 5.525000 ;
      RECT 2046.045000  2.140000 2046.215000 2.310000 ;
      RECT 2046.045000  3.130000 2046.215000 3.300000 ;
      RECT 2046.225000 -0.085000 2046.395000 0.085000 ;
      RECT 2046.225000  5.355000 2046.395000 5.525000 ;
      RECT 2046.525000  1.785000 2046.695000 1.955000 ;
      RECT 2046.525000  3.485000 2046.695000 3.655000 ;
      RECT 2046.685000 -0.085000 2046.855000 0.085000 ;
      RECT 2046.685000  5.355000 2046.855000 5.525000 ;
      RECT 2046.995000  2.140000 2047.165000 2.310000 ;
      RECT 2046.995000  3.130000 2047.165000 3.300000 ;
      RECT 2047.145000 -0.085000 2047.315000 0.085000 ;
      RECT 2047.145000  5.355000 2047.315000 5.525000 ;
      RECT 2047.465000  1.785000 2047.635000 1.955000 ;
      RECT 2047.465000  3.485000 2047.635000 3.655000 ;
      RECT 2047.605000 -0.085000 2047.775000 0.085000 ;
      RECT 2047.605000  5.355000 2047.775000 5.525000 ;
      RECT 2047.945000  2.140000 2048.115000 2.310000 ;
      RECT 2047.945000  3.130000 2048.115000 3.300000 ;
      RECT 2048.065000 -0.085000 2048.235000 0.085000 ;
      RECT 2048.065000  2.635000 2048.235000 2.805000 ;
      RECT 2048.065000  5.355000 2048.235000 5.525000 ;
      RECT 2048.525000 -0.085000 2048.695000 0.085000 ;
      RECT 2048.525000  2.635000 2048.695000 2.805000 ;
      RECT 2048.525000  5.355000 2048.695000 5.525000 ;
      RECT 2048.925000  2.140000 2049.095000 2.310000 ;
      RECT 2048.925000  3.130000 2049.095000 3.300000 ;
      RECT 2048.985000 -0.085000 2049.155000 0.085000 ;
      RECT 2048.985000  2.635000 2049.155000 2.805000 ;
      RECT 2048.985000  5.355000 2049.155000 5.525000 ;
      RECT 2049.445000 -0.085000 2049.615000 0.085000 ;
      RECT 2049.445000  2.635000 2049.615000 2.805000 ;
      RECT 2049.445000  5.355000 2049.615000 5.525000 ;
      RECT 2049.865000  2.140000 2050.035000 2.310000 ;
      RECT 2049.865000  3.130000 2050.035000 3.300000 ;
      RECT 2049.905000 -0.085000 2050.075000 0.085000 ;
      RECT 2049.905000  2.635000 2050.075000 2.805000 ;
      RECT 2049.905000  5.355000 2050.075000 5.525000 ;
      RECT 2050.365000 -0.085000 2050.535000 0.085000 ;
      RECT 2050.365000  2.635000 2050.535000 2.805000 ;
      RECT 2050.365000  5.355000 2050.535000 5.525000 ;
      RECT 2050.825000 -0.085000 2050.995000 0.085000 ;
      RECT 2050.825000  2.635000 2050.995000 2.805000 ;
      RECT 2050.825000  5.355000 2050.995000 5.525000 ;
      RECT 2051.285000 -0.085000 2051.455000 0.085000 ;
      RECT 2051.285000  2.635000 2051.455000 2.805000 ;
      RECT 2051.285000  5.355000 2051.455000 5.525000 ;
      RECT 2051.325000  2.140000 2051.495000 2.310000 ;
      RECT 2051.325000  3.130000 2051.495000 3.300000 ;
      RECT 2051.745000 -0.085000 2051.915000 0.085000 ;
      RECT 2051.745000  2.635000 2051.915000 2.805000 ;
      RECT 2051.745000  5.355000 2051.915000 5.525000 ;
      RECT 2052.205000 -0.085000 2052.375000 0.085000 ;
      RECT 2052.205000  2.635000 2052.375000 2.805000 ;
      RECT 2052.205000  5.355000 2052.375000 5.525000 ;
      RECT 2052.265000  2.140000 2052.435000 2.310000 ;
      RECT 2052.265000  3.130000 2052.435000 3.300000 ;
      RECT 2052.665000 -0.085000 2052.835000 0.085000 ;
      RECT 2052.665000  2.635000 2052.835000 2.805000 ;
      RECT 2052.665000  5.355000 2052.835000 5.525000 ;
      RECT 2053.125000 -0.085000 2053.295000 0.085000 ;
      RECT 2053.125000  2.635000 2053.295000 2.805000 ;
      RECT 2053.125000  5.355000 2053.295000 5.525000 ;
      RECT 2053.245000  2.140000 2053.415000 2.310000 ;
      RECT 2053.245000  3.130000 2053.415000 3.300000 ;
      RECT 2053.585000 -0.085000 2053.755000 0.085000 ;
      RECT 2053.585000  5.355000 2053.755000 5.525000 ;
      RECT 2053.725000  1.785000 2053.895000 1.955000 ;
      RECT 2053.725000  3.485000 2053.895000 3.655000 ;
      RECT 2054.045000 -0.085000 2054.215000 0.085000 ;
      RECT 2054.045000  5.355000 2054.215000 5.525000 ;
      RECT 2054.195000  2.140000 2054.365000 2.310000 ;
      RECT 2054.195000  3.130000 2054.365000 3.300000 ;
      RECT 2054.505000 -0.085000 2054.675000 0.085000 ;
      RECT 2054.505000  5.355000 2054.675000 5.525000 ;
      RECT 2054.665000  1.785000 2054.835000 1.955000 ;
      RECT 2054.665000  3.485000 2054.835000 3.655000 ;
      RECT 2054.965000 -0.085000 2055.135000 0.085000 ;
      RECT 2054.965000  5.355000 2055.135000 5.525000 ;
      RECT 2055.145000  2.140000 2055.315000 2.310000 ;
      RECT 2055.145000  3.130000 2055.315000 3.300000 ;
      RECT 2055.425000 -0.085000 2055.595000 0.085000 ;
      RECT 2055.425000  2.635000 2055.595000 2.805000 ;
      RECT 2055.425000  5.355000 2055.595000 5.525000 ;
      RECT 2055.885000 -0.085000 2056.055000 0.085000 ;
      RECT 2055.885000  2.635000 2056.055000 2.805000 ;
      RECT 2055.885000  5.355000 2056.055000 5.525000 ;
      RECT 2056.345000 -0.085000 2056.515000 0.085000 ;
      RECT 2056.345000  2.635000 2056.515000 2.805000 ;
      RECT 2056.345000  5.355000 2056.515000 5.525000 ;
      RECT 2056.805000 -0.085000 2056.975000 0.085000 ;
      RECT 2056.805000  2.635000 2056.975000 2.805000 ;
      RECT 2056.805000  5.355000 2056.975000 5.525000 ;
      RECT 2057.265000 -0.085000 2057.435000 0.085000 ;
      RECT 2057.265000  2.635000 2057.435000 2.805000 ;
      RECT 2057.265000  5.355000 2057.435000 5.525000 ;
      RECT 2057.725000 -0.085000 2057.895000 0.085000 ;
      RECT 2057.725000  2.635000 2057.895000 2.805000 ;
      RECT 2057.725000  5.355000 2057.895000 5.525000 ;
      RECT 2058.185000 -0.085000 2058.355000 0.085000 ;
      RECT 2058.185000  2.635000 2058.355000 2.805000 ;
      RECT 2058.185000  5.355000 2058.355000 5.525000 ;
      RECT 2058.645000 -0.085000 2058.815000 0.085000 ;
      RECT 2058.645000  2.635000 2058.815000 2.805000 ;
      RECT 2058.645000  5.355000 2058.815000 5.525000 ;
      RECT 2058.925000  2.140000 2059.095000 2.310000 ;
      RECT 2058.925000  3.130000 2059.095000 3.300000 ;
      RECT 2059.105000 -0.085000 2059.275000 0.085000 ;
      RECT 2059.105000  5.355000 2059.275000 5.525000 ;
      RECT 2059.405000  1.785000 2059.575000 1.955000 ;
      RECT 2059.405000  3.485000 2059.575000 3.655000 ;
      RECT 2059.565000 -0.085000 2059.735000 0.085000 ;
      RECT 2059.565000  5.355000 2059.735000 5.525000 ;
      RECT 2059.875000  2.140000 2060.045000 2.310000 ;
      RECT 2059.875000  3.130000 2060.045000 3.300000 ;
      RECT 2060.025000 -0.085000 2060.195000 0.085000 ;
      RECT 2060.025000  5.355000 2060.195000 5.525000 ;
      RECT 2060.345000  1.785000 2060.515000 1.955000 ;
      RECT 2060.345000  3.485000 2060.515000 3.655000 ;
      RECT 2060.485000 -0.085000 2060.655000 0.085000 ;
      RECT 2060.485000  5.355000 2060.655000 5.525000 ;
      RECT 2060.825000  2.140000 2060.995000 2.310000 ;
      RECT 2060.825000  3.130000 2060.995000 3.300000 ;
      RECT 2060.945000 -0.085000 2061.115000 0.085000 ;
      RECT 2060.945000  2.635000 2061.115000 2.805000 ;
      RECT 2060.945000  5.355000 2061.115000 5.525000 ;
      RECT 2061.405000 -0.085000 2061.575000 0.085000 ;
      RECT 2061.405000  2.635000 2061.575000 2.805000 ;
      RECT 2061.405000  5.355000 2061.575000 5.525000 ;
      RECT 2061.805000  2.140000 2061.975000 2.310000 ;
      RECT 2061.805000  3.130000 2061.975000 3.300000 ;
      RECT 2061.865000 -0.085000 2062.035000 0.085000 ;
      RECT 2061.865000  2.635000 2062.035000 2.805000 ;
      RECT 2061.865000  5.355000 2062.035000 5.525000 ;
      RECT 2062.325000 -0.085000 2062.495000 0.085000 ;
      RECT 2062.325000  2.635000 2062.495000 2.805000 ;
      RECT 2062.325000  5.355000 2062.495000 5.525000 ;
      RECT 2062.745000  2.140000 2062.915000 2.310000 ;
      RECT 2062.745000  3.130000 2062.915000 3.300000 ;
      RECT 2062.785000 -0.085000 2062.955000 0.085000 ;
      RECT 2062.785000  2.635000 2062.955000 2.805000 ;
      RECT 2062.785000  5.355000 2062.955000 5.525000 ;
      RECT 2063.245000 -0.085000 2063.415000 0.085000 ;
      RECT 2063.245000  2.635000 2063.415000 2.805000 ;
      RECT 2063.245000  5.355000 2063.415000 5.525000 ;
      RECT 2063.705000 -0.085000 2063.875000 0.085000 ;
      RECT 2063.705000  2.635000 2063.875000 2.805000 ;
      RECT 2063.705000  5.355000 2063.875000 5.525000 ;
    LAYER met1 ;
      RECT   -0.380000 -0.070000 2064.400000  0.070000 ;
      RECT   -0.380000  0.070000   -0.240000  5.370000 ;
      RECT   -0.380000  5.370000  234.600000  5.510000 ;
      RECT    0.000000 -0.240000 2064.020000 -0.070000 ;
      RECT    0.000000  0.070000 2064.020000  0.240000 ;
      RECT    0.000000  2.480000 2064.020000  2.960000 ;
      RECT    0.000000  5.200000  234.600000  5.370000 ;
      RECT    0.000000  5.510000  234.600000  5.680000 ;
      RECT   29.525000  1.415000   29.815000  1.460000 ;
      RECT   29.525000  1.460000   32.870000  1.600000 ;
      RECT   29.525000  1.600000   29.815000  1.645000 ;
      RECT   32.580000  1.415000   32.870000  1.460000 ;
      RECT   32.580000  1.600000   32.870000  1.645000 ;
      RECT   52.095000  4.815000   52.385000  4.860000 ;
      RECT   52.095000  4.860000   61.885000  5.000000 ;
      RECT   52.095000  5.000000   52.385000  5.045000 ;
      RECT   52.565000  3.455000   52.855000  3.500000 ;
      RECT   52.565000  3.500000   59.015000  3.640000 ;
      RECT   52.565000  3.640000   52.855000  3.685000 ;
      RECT   53.505000  3.455000   53.795000  3.500000 ;
      RECT   53.505000  3.640000   53.795000  3.685000 ;
      RECT   54.965000  3.115000   55.255000  3.160000 ;
      RECT   54.965000  3.160000   59.640000  3.300000 ;
      RECT   54.965000  3.300000   55.255000  3.345000 ;
      RECT   55.905000  3.115000   56.195000  3.160000 ;
      RECT   55.905000  3.300000   56.195000  3.345000 ;
      RECT   57.785000  3.455000   58.075000  3.500000 ;
      RECT   57.785000  3.640000   58.075000  3.685000 ;
      RECT   58.725000  3.455000   59.015000  3.500000 ;
      RECT   58.725000  3.640000   59.015000  3.685000 ;
      RECT   59.500000  3.300000   59.640000  3.500000 ;
      RECT   59.500000  3.500000   61.415000  3.640000 ;
      RECT   60.185000  3.455000   60.475000  3.500000 ;
      RECT   60.185000  3.640000   60.475000  3.685000 ;
      RECT   61.125000  3.455000   61.415000  3.500000 ;
      RECT   61.125000  3.640000   61.415000  3.685000 ;
      RECT   61.595000  4.815000   61.885000  4.860000 ;
      RECT   61.595000  5.000000   61.885000  5.045000 ;
      RECT   69.115000  4.815000   69.405000  4.860000 ;
      RECT   69.115000  4.860000   78.905000  5.000000 ;
      RECT   69.115000  5.000000   69.405000  5.045000 ;
      RECT   69.585000  3.455000   69.875000  3.500000 ;
      RECT   69.585000  3.500000   76.035000  3.640000 ;
      RECT   69.585000  3.640000   69.875000  3.685000 ;
      RECT   70.525000  3.455000   70.815000  3.500000 ;
      RECT   70.525000  3.640000   70.815000  3.685000 ;
      RECT   71.985000  3.115000   72.275000  3.160000 ;
      RECT   71.985000  3.160000   76.660000  3.300000 ;
      RECT   71.985000  3.300000   72.275000  3.345000 ;
      RECT   72.925000  3.115000   73.215000  3.160000 ;
      RECT   72.925000  3.300000   73.215000  3.345000 ;
      RECT   74.805000  3.455000   75.095000  3.500000 ;
      RECT   74.805000  3.640000   75.095000  3.685000 ;
      RECT   75.745000  3.455000   76.035000  3.500000 ;
      RECT   75.745000  3.640000   76.035000  3.685000 ;
      RECT   76.520000  3.300000   76.660000  3.500000 ;
      RECT   76.520000  3.500000   78.435000  3.640000 ;
      RECT   77.205000  3.455000   77.495000  3.500000 ;
      RECT   77.205000  3.640000   77.495000  3.685000 ;
      RECT   78.145000  3.455000   78.435000  3.500000 ;
      RECT   78.145000  3.640000   78.435000  3.685000 ;
      RECT   78.615000  4.815000   78.905000  4.860000 ;
      RECT   78.615000  5.000000   78.905000  5.045000 ;
      RECT  156.185000  4.120000  156.825000  4.135000 ;
      RECT  156.185000  4.135000  157.870000  4.365000 ;
      RECT  156.185000  4.365000  156.825000  4.380000 ;
      RECT  166.145000  3.115000  166.435000  3.345000 ;
      RECT  166.220000  2.960000  166.360000  3.115000 ;
      RECT  166.605000  3.455000  166.895000  3.685000 ;
      RECT  166.680000  2.960000  166.820000  3.455000 ;
      RECT  167.780000  1.415000  168.120000  1.460000 ;
      RECT  167.780000  1.460000  171.100000  1.600000 ;
      RECT  167.780000  1.600000  168.120000  1.645000 ;
      RECT  170.810000  1.415000  171.100000  1.460000 ;
      RECT  170.810000  1.600000  171.100000  1.645000 ;
      RECT  175.440000  4.120000  176.080000  4.180000 ;
      RECT  175.440000  4.180000  178.315000  4.320000 ;
      RECT  175.440000  4.320000  176.080000  4.380000 ;
      RECT  177.665000  4.135000  178.315000  4.180000 ;
      RECT  177.665000  4.320000  178.315000  4.365000 ;
      RECT  180.435000  3.455000  180.725000  3.500000 ;
      RECT  180.435000  3.500000  183.370000  3.640000 ;
      RECT  180.435000  3.640000  180.725000  3.685000 ;
      RECT  180.895000  3.795000  181.185000  3.840000 ;
      RECT  180.895000  3.840000  182.815000  3.980000 ;
      RECT  180.895000  3.980000  181.185000  4.025000 ;
      RECT  182.525000  3.795000  182.815000  3.840000 ;
      RECT  182.525000  3.980000  182.815000  4.025000 ;
      RECT  183.080000  3.455000  183.370000  3.500000 ;
      RECT  183.080000  3.640000  183.370000  3.685000 ;
      RECT  187.305000  3.795000  187.595000  3.840000 ;
      RECT  187.305000  3.840000  189.715000  3.980000 ;
      RECT  187.305000  3.980000  187.595000  4.025000 ;
      RECT  187.815000  3.455000  188.105000  3.500000 ;
      RECT  187.815000  3.500000  190.270000  3.640000 ;
      RECT  187.815000  3.640000  188.105000  3.685000 ;
      RECT  189.425000  3.795000  189.715000  3.840000 ;
      RECT  189.425000  3.980000  189.715000  4.025000 ;
      RECT  189.980000  3.455000  190.270000  3.500000 ;
      RECT  189.980000  3.640000  190.270000  3.685000 ;
      RECT  194.235000  3.455000  194.525000  3.500000 ;
      RECT  194.235000  3.500000  197.170000  3.640000 ;
      RECT  194.235000  3.640000  194.525000  3.685000 ;
      RECT  194.695000  3.795000  194.985000  3.840000 ;
      RECT  194.695000  3.840000  196.615000  3.980000 ;
      RECT  194.695000  3.980000  194.985000  4.025000 ;
      RECT  196.325000  3.795000  196.615000  3.840000 ;
      RECT  196.325000  3.980000  196.615000  4.025000 ;
      RECT  196.880000  3.455000  197.170000  3.500000 ;
      RECT  196.880000  3.640000  197.170000  3.685000 ;
      RECT  201.565000  3.795000  201.855000  3.840000 ;
      RECT  201.565000  3.840000  203.975000  3.980000 ;
      RECT  201.565000  3.980000  201.855000  4.025000 ;
      RECT  202.075000  3.455000  202.365000  3.500000 ;
      RECT  202.075000  3.500000  204.530000  3.640000 ;
      RECT  202.075000  3.640000  202.365000  3.685000 ;
      RECT  203.685000  3.795000  203.975000  3.840000 ;
      RECT  203.685000  3.980000  203.975000  4.025000 ;
      RECT  204.240000  3.455000  204.530000  3.500000 ;
      RECT  204.240000  3.640000  204.530000  3.685000 ;
      RECT  208.955000  3.455000  209.245000  3.500000 ;
      RECT  208.955000  3.500000  211.890000  3.640000 ;
      RECT  208.955000  3.640000  209.245000  3.685000 ;
      RECT  209.415000  3.795000  209.705000  3.840000 ;
      RECT  209.415000  3.840000  211.335000  3.980000 ;
      RECT  209.415000  3.980000  209.705000  4.025000 ;
      RECT  211.045000  3.795000  211.335000  3.840000 ;
      RECT  211.045000  3.980000  211.335000  4.025000 ;
      RECT  211.600000  3.455000  211.890000  3.500000 ;
      RECT  211.600000  3.640000  211.890000  3.685000 ;
      RECT  217.205000  3.795000  217.495000  3.840000 ;
      RECT  217.205000  3.840000  219.615000  3.980000 ;
      RECT  217.205000  3.980000  217.495000  4.025000 ;
      RECT  217.715000  3.455000  218.005000  3.500000 ;
      RECT  217.715000  3.500000  220.170000  3.640000 ;
      RECT  217.715000  3.640000  218.005000  3.685000 ;
      RECT  219.325000  3.795000  219.615000  3.840000 ;
      RECT  219.325000  3.980000  219.615000  4.025000 ;
      RECT  219.880000  3.455000  220.170000  3.500000 ;
      RECT  219.880000  3.640000  220.170000  3.685000 ;
      RECT  475.415000  1.075000  476.215000  1.120000 ;
      RECT  475.415000  1.120000  484.935000  1.260000 ;
      RECT  475.415000  1.260000  476.215000  1.305000 ;
      RECT  484.085000  1.075000  484.935000  1.120000 ;
      RECT  484.085000  1.260000  484.935000  1.305000 ;
      RECT  508.440000  1.075000  508.730000  1.120000 ;
      RECT  508.440000  1.120000  514.090000  1.260000 ;
      RECT  508.440000  1.260000  508.730000  1.305000 ;
      RECT  508.845000  1.755000  509.185000  1.800000 ;
      RECT  508.845000  1.800000  514.540000  1.940000 ;
      RECT  508.845000  1.940000  509.185000  1.985000 ;
      RECT  510.260000  1.075000  510.550000  1.120000 ;
      RECT  510.260000  1.260000  510.550000  1.305000 ;
      RECT  510.505000  1.755000  510.795000  1.800000 ;
      RECT  510.505000  1.940000  510.795000  1.985000 ;
      RECT  511.835000  0.735000  512.585000  0.780000 ;
      RECT  511.835000  0.780000  515.705000  0.920000 ;
      RECT  511.835000  0.920000  512.585000  0.965000 ;
      RECT  513.800000  1.075000  514.090000  1.120000 ;
      RECT  513.800000  1.260000  514.090000  1.305000 ;
      RECT  514.250000  1.755000  514.540000  1.800000 ;
      RECT  514.250000  1.940000  514.540000  1.985000 ;
      RECT  515.415000  0.735000  515.705000  0.780000 ;
      RECT  515.415000  0.920000  515.705000  0.965000 ;
      RECT  518.560000  1.075000  518.850000  1.120000 ;
      RECT  518.560000  1.120000  524.210000  1.260000 ;
      RECT  518.560000  1.260000  518.850000  1.305000 ;
      RECT  518.965000  1.755000  519.305000  1.800000 ;
      RECT  518.965000  1.800000  524.660000  1.940000 ;
      RECT  518.965000  1.940000  519.305000  1.985000 ;
      RECT  520.380000  1.075000  520.670000  1.120000 ;
      RECT  520.380000  1.260000  520.670000  1.305000 ;
      RECT  520.625000  1.755000  520.915000  1.800000 ;
      RECT  520.625000  1.940000  520.915000  1.985000 ;
      RECT  521.955000  0.735000  522.705000  0.780000 ;
      RECT  521.955000  0.780000  525.825000  0.920000 ;
      RECT  521.955000  0.920000  522.705000  0.965000 ;
      RECT  523.920000  1.075000  524.210000  1.120000 ;
      RECT  523.920000  1.260000  524.210000  1.305000 ;
      RECT  524.370000  1.755000  524.660000  1.800000 ;
      RECT  524.370000  1.940000  524.660000  1.985000 ;
      RECT  525.535000  0.735000  525.825000  0.780000 ;
      RECT  525.535000  0.920000  525.825000  0.965000 ;
      RECT  529.140000  1.075000  529.430000  1.120000 ;
      RECT  529.140000  1.120000  535.345000  1.260000 ;
      RECT  529.140000  1.260000  529.430000  1.305000 ;
      RECT  529.545000  1.755000  529.885000  1.800000 ;
      RECT  529.545000  1.800000  535.345000  1.940000 ;
      RECT  529.545000  1.940000  529.885000  1.985000 ;
      RECT  531.075000  1.075000  531.365000  1.120000 ;
      RECT  531.075000  1.260000  531.365000  1.305000 ;
      RECT  531.585000  1.755000  531.875000  1.800000 ;
      RECT  531.585000  1.940000  531.875000  1.985000 ;
      RECT  532.715000  0.735000  533.465000  0.780000 ;
      RECT  532.715000  0.780000  536.935000  0.920000 ;
      RECT  532.715000  0.920000  533.465000  0.965000 ;
      RECT  535.005000  1.075000  535.345000  1.120000 ;
      RECT  535.005000  1.260000  535.345000  1.305000 ;
      RECT  535.005000  1.755000  535.345000  1.800000 ;
      RECT  535.005000  1.940000  535.345000  1.985000 ;
      RECT  536.350000  0.920000  536.935000  1.280000 ;
      RECT  536.645000  0.735000  536.935000  0.780000 ;
      RECT  541.105000  1.710000  541.395000  1.800000 ;
      RECT  541.105000  1.800000  546.435000  1.940000 ;
      RECT  541.605000  0.690000  541.895000  0.780000 ;
      RECT  541.605000  0.780000  543.885000  0.920000 ;
      RECT  543.085000  1.710000  543.375000  1.800000 ;
      RECT  543.595000  0.690000  543.885000  0.780000 ;
      RECT  543.670000  0.920000  543.885000  1.120000 ;
      RECT  543.670000  1.120000  546.455000  1.260000 ;
      RECT  544.720000  0.735000  545.010000  0.780000 ;
      RECT  544.720000  0.780000  548.235000  0.920000 ;
      RECT  544.720000  0.920000  545.010000  0.965000 ;
      RECT  546.145000  1.710000  546.435000  1.800000 ;
      RECT  546.165000  1.080000  546.455000  1.120000 ;
      RECT  546.165000  1.260000  546.455000  1.310000 ;
      RECT  547.945000  0.735000  548.235000  0.780000 ;
      RECT  547.945000  0.920000  548.235000  0.965000 ;
      RECT  551.685000  1.710000  551.975000  1.800000 ;
      RECT  551.685000  1.800000  557.015000  1.940000 ;
      RECT  552.185000  0.690000  552.475000  0.780000 ;
      RECT  552.185000  0.780000  554.465000  0.920000 ;
      RECT  553.665000  1.710000  553.955000  1.800000 ;
      RECT  554.175000  0.690000  554.465000  0.780000 ;
      RECT  554.250000  0.920000  554.465000  1.120000 ;
      RECT  554.250000  1.120000  557.035000  1.260000 ;
      RECT  555.300000  0.735000  555.590000  0.780000 ;
      RECT  555.300000  0.780000  558.815000  0.920000 ;
      RECT  555.300000  0.920000  555.590000  0.965000 ;
      RECT  556.725000  1.710000  557.015000  1.800000 ;
      RECT  556.745000  1.080000  557.035000  1.120000 ;
      RECT  556.745000  1.260000  557.035000  1.310000 ;
      RECT  558.525000  0.735000  558.815000  0.780000 ;
      RECT  558.525000  0.920000  558.815000  0.965000 ;
      RECT  562.725000  1.710000  563.015000  1.800000 ;
      RECT  562.725000  1.800000  568.055000  1.940000 ;
      RECT  563.225000  0.690000  563.515000  0.780000 ;
      RECT  563.225000  0.780000  565.505000  0.920000 ;
      RECT  564.705000  1.710000  564.995000  1.800000 ;
      RECT  565.215000  0.690000  565.505000  0.780000 ;
      RECT  565.290000  0.920000  565.505000  1.120000 ;
      RECT  565.290000  1.120000  568.075000  1.260000 ;
      RECT  566.340000  0.735000  566.630000  0.780000 ;
      RECT  566.340000  0.780000  569.855000  0.920000 ;
      RECT  566.340000  0.920000  566.630000  0.965000 ;
      RECT  567.765000  1.710000  568.055000  1.800000 ;
      RECT  567.785000  1.080000  568.075000  1.120000 ;
      RECT  567.785000  1.260000  568.075000  1.310000 ;
      RECT  569.565000  0.735000  569.855000  0.780000 ;
      RECT  569.565000  0.920000  569.855000  0.965000 ;
      RECT  575.140000  1.415000  575.430000  1.460000 ;
      RECT  575.140000  1.460000  577.945000  1.600000 ;
      RECT  575.140000  1.600000  575.430000  1.645000 ;
      RECT  575.650000  1.755000  575.940000  1.800000 ;
      RECT  575.650000  1.800000  577.440000  1.940000 ;
      RECT  575.650000  1.940000  575.940000  1.985000 ;
      RECT  577.150000  1.755000  577.440000  1.800000 ;
      RECT  577.150000  1.940000  577.440000  1.985000 ;
      RECT  577.655000  1.415000  577.945000  1.460000 ;
      RECT  577.655000  1.600000  577.945000  1.645000 ;
      RECT  581.580000  1.415000  581.870000  1.460000 ;
      RECT  581.580000  1.460000  584.385000  1.600000 ;
      RECT  581.580000  1.600000  581.870000  1.645000 ;
      RECT  582.090000  1.755000  582.380000  1.800000 ;
      RECT  582.090000  1.800000  583.880000  1.940000 ;
      RECT  582.090000  1.940000  582.380000  1.985000 ;
      RECT  583.590000  1.755000  583.880000  1.800000 ;
      RECT  583.590000  1.940000  583.880000  1.985000 ;
      RECT  584.095000  1.415000  584.385000  1.460000 ;
      RECT  584.095000  1.600000  584.385000  1.645000 ;
      RECT  588.480000  1.370000  588.770000  1.460000 ;
      RECT  588.480000  1.460000  591.290000  1.600000 ;
      RECT  588.935000  1.740000  589.225000  1.800000 ;
      RECT  588.935000  1.800000  590.780000  1.940000 ;
      RECT  588.935000  1.940000  589.225000  1.970000 ;
      RECT  590.490000  1.740000  590.780000  1.800000 ;
      RECT  590.490000  1.940000  590.780000  1.970000 ;
      RECT  590.995000  1.370000  591.290000  1.460000 ;
      RECT  611.425000  1.030000  611.720000  1.120000 ;
      RECT  611.425000  1.120000  615.250000  1.260000 ;
      RECT  614.910000  1.030000  615.250000  1.120000 ;
      RECT  616.485000  1.075000  616.780000  1.165000 ;
      RECT  616.485000  1.165000  621.340000  1.305000 ;
      RECT  621.050000  1.075000  621.340000  1.165000 ;
      RECT  623.845000  1.030000  624.185000  1.120000 ;
      RECT  623.845000  1.120000  631.160000  1.260000 ;
      RECT  630.820000  1.030000  631.160000  1.120000 ;
      RECT  734.180000  1.075000  734.520000  1.120000 ;
      RECT  734.180000  1.120000  738.675000  1.260000 ;
      RECT  734.180000  1.260000  734.520000  1.305000 ;
      RECT  734.670000  0.735000  734.960000  0.780000 ;
      RECT  734.670000  0.780000  737.990000  0.920000 ;
      RECT  734.670000  0.920000  734.960000  0.965000 ;
      RECT  735.670000  1.415000  735.960000  1.460000 ;
      RECT  735.670000  1.460000  739.595000  1.600000 ;
      RECT  735.670000  1.600000  735.960000  1.645000 ;
      RECT  737.650000  0.735000  737.990000  0.780000 ;
      RECT  737.650000  0.920000  737.990000  0.965000 ;
      RECT  738.325000  1.075000  738.675000  1.120000 ;
      RECT  738.325000  1.260000  738.675000  1.305000 ;
      RECT  739.305000  1.415000  739.595000  1.460000 ;
      RECT  739.305000  1.600000  739.595000  1.645000 ;
      RECT  746.310000  0.735000  746.600000  0.780000 ;
      RECT  746.310000  0.780000  749.680000  0.920000 ;
      RECT  746.310000  0.920000  746.600000  0.965000 ;
      RECT  749.340000  0.735000  749.680000  0.780000 ;
      RECT  749.340000  0.920000  749.680000  0.965000 ;
      RECT  752.800000  0.735000  753.090000  0.780000 ;
      RECT  752.800000  0.780000  758.210000  0.920000 ;
      RECT  752.800000  0.920000  753.090000  0.965000 ;
      RECT  757.870000  0.735000  758.210000  0.780000 ;
      RECT  757.870000  0.920000  758.210000  0.965000 ;
      RECT  867.740000  1.075000  870.025000  1.305000 ;
      RECT  875.275000  1.075000  875.565000  1.120000 ;
      RECT  875.275000  1.120000  878.115000  1.260000 ;
      RECT  875.275000  1.260000  875.565000  1.305000 ;
      RECT  877.775000  1.075000  878.115000  1.120000 ;
      RECT  877.775000  1.260000  878.115000  1.305000 ;
      RECT  926.775000  2.065000  927.120000  2.140000 ;
      RECT  926.775000  2.140000  930.180000  2.280000 ;
      RECT  926.775000  2.280000  927.120000  2.335000 ;
      RECT  929.835000  2.065000  930.180000  2.140000 ;
      RECT  929.835000  2.280000  930.180000  2.335000 ;
      RECT 1034.730000  0.395000 1035.020000  0.440000 ;
      RECT 1034.730000  0.440000 1042.170000  0.580000 ;
      RECT 1034.730000  0.580000 1035.020000  0.625000 ;
      RECT 1041.880000  0.395000 1042.170000  0.440000 ;
      RECT 1041.880000  0.580000 1042.170000  0.625000 ;
      RECT 1188.515000  1.385000 1188.855000  1.460000 ;
      RECT 1188.515000  1.460000 1191.840000  1.600000 ;
      RECT 1188.515000  1.600000 1188.855000  1.635000 ;
      RECT 1191.545000  1.395000 1191.840000  1.460000 ;
      RECT 1191.545000  1.600000 1191.840000  1.645000 ;
      RECT 1350.235000  1.755000 1350.525000  1.800000 ;
      RECT 1350.235000  1.800000 1359.045000  1.940000 ;
      RECT 1350.235000  1.940000 1350.525000  1.985000 ;
      RECT 1350.730000  0.735000 1351.020000  0.780000 ;
      RECT 1350.730000  0.780000 1355.525000  0.920000 ;
      RECT 1350.730000  0.920000 1351.020000  0.965000 ;
      RECT 1352.685000  1.075000 1352.975000  1.120000 ;
      RECT 1352.685000  1.120000 1354.515000  1.260000 ;
      RECT 1352.685000  1.260000 1352.975000  1.305000 ;
      RECT 1354.225000  1.075000 1354.515000  1.120000 ;
      RECT 1354.225000  1.260000 1354.515000  1.305000 ;
      RECT 1354.725000  1.755000 1355.015000  1.800000 ;
      RECT 1354.725000  1.940000 1355.015000  1.985000 ;
      RECT 1355.235000  0.735000 1355.525000  0.780000 ;
      RECT 1355.235000  0.920000 1355.525000  0.965000 ;
      RECT 1355.310000  0.965000 1355.525000  1.120000 ;
      RECT 1355.310000  1.120000 1359.045000  1.260000 ;
      RECT 1356.165000  0.735000 1356.455000  0.780000 ;
      RECT 1356.165000  0.780000 1360.585000  0.920000 ;
      RECT 1356.165000  0.920000 1356.455000  0.965000 ;
      RECT 1358.295000  1.415000 1358.585000  1.460000 ;
      RECT 1358.295000  1.460000 1362.035000  1.600000 ;
      RECT 1358.295000  1.600000 1358.585000  1.645000 ;
      RECT 1358.755000  1.075000 1359.045000  1.120000 ;
      RECT 1358.755000  1.260000 1359.045000  1.305000 ;
      RECT 1358.755000  1.755000 1359.045000  1.800000 ;
      RECT 1358.755000  1.940000 1359.045000  1.985000 ;
      RECT 1360.295000  0.735000 1360.585000  0.780000 ;
      RECT 1360.295000  0.920000 1360.585000  0.965000 ;
      RECT 1361.745000  1.415000 1362.035000  1.460000 ;
      RECT 1361.745000  1.600000 1362.035000  1.645000 ;
      RECT 1366.535000  1.075000 1366.825000  1.120000 ;
      RECT 1366.535000  1.120000 1375.205000  1.260000 ;
      RECT 1366.535000  1.260000 1366.825000  1.305000 ;
      RECT 1366.810000  1.755000 1367.110000  1.800000 ;
      RECT 1366.810000  1.800000 1375.535000  1.940000 ;
      RECT 1366.810000  1.940000 1367.110000  1.985000 ;
      RECT 1371.160000  1.075000 1371.450000  1.120000 ;
      RECT 1371.160000  1.260000 1371.450000  1.305000 ;
      RECT 1371.630000  1.755000 1371.920000  1.800000 ;
      RECT 1371.630000  1.940000 1371.920000  1.985000 ;
      RECT 1372.885000  0.735000 1373.640000  0.780000 ;
      RECT 1372.885000  0.780000 1377.145000  0.920000 ;
      RECT 1372.885000  0.920000 1373.640000  0.965000 ;
      RECT 1374.895000  1.075000 1375.205000  1.120000 ;
      RECT 1374.895000  1.260000 1375.205000  1.305000 ;
      RECT 1375.240000  1.755000 1375.535000  1.800000 ;
      RECT 1375.240000  1.940000 1375.535000  1.985000 ;
      RECT 1376.855000  0.735000 1377.145000  0.780000 ;
      RECT 1376.855000  0.920000 1377.145000  0.965000 ;
      RECT 1381.255000  1.075000 1381.545000  1.120000 ;
      RECT 1381.255000  1.120000 1389.925000  1.260000 ;
      RECT 1381.255000  1.260000 1381.545000  1.305000 ;
      RECT 1381.530000  1.755000 1381.830000  1.800000 ;
      RECT 1381.530000  1.800000 1390.255000  1.940000 ;
      RECT 1381.530000  1.940000 1381.830000  1.985000 ;
      RECT 1385.880000  1.075000 1386.170000  1.120000 ;
      RECT 1385.880000  1.260000 1386.170000  1.305000 ;
      RECT 1386.350000  1.755000 1386.640000  1.800000 ;
      RECT 1386.350000  1.940000 1386.640000  1.985000 ;
      RECT 1387.605000  0.735000 1388.360000  0.780000 ;
      RECT 1387.605000  0.780000 1391.865000  0.920000 ;
      RECT 1387.605000  0.920000 1388.360000  0.965000 ;
      RECT 1389.615000  1.075000 1389.925000  1.120000 ;
      RECT 1389.615000  1.260000 1389.925000  1.305000 ;
      RECT 1389.960000  1.755000 1390.255000  1.800000 ;
      RECT 1389.960000  1.940000 1390.255000  1.985000 ;
      RECT 1391.575000  0.735000 1391.865000  0.780000 ;
      RECT 1391.575000  0.920000 1391.865000  0.965000 ;
      RECT 1396.300000  1.755000 1396.600000  1.800000 ;
      RECT 1396.300000  1.800000 1405.435000  1.940000 ;
      RECT 1396.300000  1.940000 1396.600000  1.985000 ;
      RECT 1396.775000  1.075000 1397.065000  1.120000 ;
      RECT 1396.775000  1.120000 1405.105000  1.260000 ;
      RECT 1396.775000  1.260000 1397.065000  1.305000 ;
      RECT 1401.060000  1.075000 1401.350000  1.120000 ;
      RECT 1401.060000  1.260000 1401.350000  1.305000 ;
      RECT 1401.530000  1.755000 1401.820000  1.800000 ;
      RECT 1401.530000  1.940000 1401.820000  1.985000 ;
      RECT 1402.785000  0.735000 1403.540000  0.780000 ;
      RECT 1402.785000  0.780000 1407.045000  0.920000 ;
      RECT 1402.785000  0.920000 1403.540000  0.965000 ;
      RECT 1404.795000  1.075000 1405.105000  1.120000 ;
      RECT 1404.795000  1.260000 1405.105000  1.305000 ;
      RECT 1405.140000  1.755000 1405.435000  1.800000 ;
      RECT 1405.140000  1.940000 1405.435000  1.985000 ;
      RECT 1406.755000  0.735000 1407.045000  0.780000 ;
      RECT 1406.755000  0.920000 1407.045000  0.965000 ;
      RECT 1409.775000  1.075000 1410.065000  1.120000 ;
      RECT 1409.775000  1.120000 1418.445000  1.260000 ;
      RECT 1409.775000  1.260000 1410.065000  1.305000 ;
      RECT 1410.050000  1.755000 1410.350000  1.800000 ;
      RECT 1410.050000  1.800000 1418.775000  1.940000 ;
      RECT 1410.050000  1.940000 1410.350000  1.985000 ;
      RECT 1414.400000  1.075000 1414.690000  1.120000 ;
      RECT 1414.400000  1.260000 1414.690000  1.305000 ;
      RECT 1414.870000  1.755000 1415.160000  1.800000 ;
      RECT 1414.870000  1.940000 1415.160000  1.985000 ;
      RECT 1416.125000  0.735000 1416.880000  0.780000 ;
      RECT 1416.125000  0.780000 1420.385000  0.920000 ;
      RECT 1416.125000  0.920000 1416.880000  0.965000 ;
      RECT 1418.135000  1.075000 1418.445000  1.120000 ;
      RECT 1418.135000  1.260000 1418.445000  1.305000 ;
      RECT 1418.480000  1.755000 1418.775000  1.800000 ;
      RECT 1418.480000  1.940000 1418.775000  1.985000 ;
      RECT 1420.095000  0.735000 1420.385000  0.780000 ;
      RECT 1420.095000  0.920000 1420.385000  0.965000 ;
      RECT 1423.115000  1.075000 1423.405000  1.120000 ;
      RECT 1423.115000  1.120000 1431.785000  1.260000 ;
      RECT 1423.115000  1.260000 1423.405000  1.305000 ;
      RECT 1423.390000  1.755000 1423.690000  1.800000 ;
      RECT 1423.390000  1.800000 1432.115000  1.940000 ;
      RECT 1423.390000  1.940000 1423.690000  1.985000 ;
      RECT 1427.740000  1.075000 1428.030000  1.120000 ;
      RECT 1427.740000  1.260000 1428.030000  1.305000 ;
      RECT 1428.210000  1.755000 1428.500000  1.800000 ;
      RECT 1428.210000  1.940000 1428.500000  1.985000 ;
      RECT 1429.465000  0.735000 1430.220000  0.780000 ;
      RECT 1429.465000  0.780000 1433.690000  0.920000 ;
      RECT 1429.465000  0.920000 1430.220000  0.965000 ;
      RECT 1431.475000  1.075000 1431.785000  1.120000 ;
      RECT 1431.475000  1.260000 1431.785000  1.305000 ;
      RECT 1431.820000  1.755000 1432.115000  1.800000 ;
      RECT 1431.820000  1.940000 1432.115000  1.985000 ;
      RECT 1433.400000  0.735000 1433.690000  0.780000 ;
      RECT 1433.400000  0.920000 1433.690000  0.965000 ;
      RECT 1436.690000  1.075000 1436.980000  1.120000 ;
      RECT 1436.690000  1.120000 1438.995000  1.260000 ;
      RECT 1436.690000  1.260000 1436.980000  1.305000 ;
      RECT 1437.735000  1.415000 1438.075000  1.460000 ;
      RECT 1437.735000  1.460000 1441.360000  1.600000 ;
      RECT 1437.735000  1.600000 1438.075000  1.645000 ;
      RECT 1438.705000  1.075000 1438.995000  1.120000 ;
      RECT 1438.705000  1.260000 1438.995000  1.305000 ;
      RECT 1440.185000  1.755000 1440.525000  1.800000 ;
      RECT 1440.185000  1.800000 1444.555000  1.940000 ;
      RECT 1440.185000  1.940000 1440.525000  1.985000 ;
      RECT 1440.645000  1.075000 1440.935000  1.120000 ;
      RECT 1440.645000  1.120000 1445.575000  1.260000 ;
      RECT 1440.645000  1.260000 1440.935000  1.305000 ;
      RECT 1441.070000  1.415000 1441.360000  1.460000 ;
      RECT 1441.070000  1.600000 1441.360000  1.645000 ;
      RECT 1441.665000  1.755000 1442.005000  1.800000 ;
      RECT 1441.665000  1.940000 1442.005000  1.985000 ;
      RECT 1443.505000  1.415000 1443.845000  1.460000 ;
      RECT 1443.505000  1.460000 1446.085000  1.600000 ;
      RECT 1443.505000  1.600000 1443.845000  1.645000 ;
      RECT 1444.265000  1.755000 1444.555000  1.800000 ;
      RECT 1444.265000  1.940000 1444.555000  1.985000 ;
      RECT 1445.235000  1.075000 1445.575000  1.120000 ;
      RECT 1445.235000  1.260000 1445.575000  1.305000 ;
      RECT 1445.795000  1.415000 1446.085000  1.460000 ;
      RECT 1445.795000  1.600000 1446.085000  1.645000 ;
      RECT 1451.870000  1.075000 1452.160000  1.120000 ;
      RECT 1451.870000  1.120000 1454.175000  1.260000 ;
      RECT 1451.870000  1.260000 1452.160000  1.305000 ;
      RECT 1452.915000  1.415000 1453.255000  1.460000 ;
      RECT 1452.915000  1.460000 1456.540000  1.600000 ;
      RECT 1452.915000  1.600000 1453.255000  1.645000 ;
      RECT 1453.885000  1.075000 1454.175000  1.120000 ;
      RECT 1453.885000  1.260000 1454.175000  1.305000 ;
      RECT 1455.365000  1.755000 1455.705000  1.800000 ;
      RECT 1455.365000  1.800000 1459.735000  1.940000 ;
      RECT 1455.365000  1.940000 1455.705000  1.985000 ;
      RECT 1455.825000  1.075000 1456.115000  1.120000 ;
      RECT 1455.825000  1.120000 1460.755000  1.260000 ;
      RECT 1455.825000  1.260000 1456.115000  1.305000 ;
      RECT 1456.250000  1.415000 1456.540000  1.460000 ;
      RECT 1456.250000  1.600000 1456.540000  1.645000 ;
      RECT 1456.845000  1.755000 1457.185000  1.800000 ;
      RECT 1456.845000  1.940000 1457.185000  1.985000 ;
      RECT 1458.685000  1.415000 1459.025000  1.460000 ;
      RECT 1458.685000  1.460000 1461.265000  1.600000 ;
      RECT 1458.685000  1.600000 1459.025000  1.645000 ;
      RECT 1459.445000  1.755000 1459.735000  1.800000 ;
      RECT 1459.445000  1.940000 1459.735000  1.985000 ;
      RECT 1460.415000  1.075000 1460.755000  1.120000 ;
      RECT 1460.415000  1.260000 1460.755000  1.305000 ;
      RECT 1460.975000  1.415000 1461.265000  1.460000 ;
      RECT 1460.975000  1.600000 1461.265000  1.645000 ;
      RECT 1467.980000  1.075000 1468.270000  1.120000 ;
      RECT 1467.980000  1.120000 1470.275000  1.260000 ;
      RECT 1467.980000  1.260000 1468.270000  1.305000 ;
      RECT 1469.015000  1.415000 1469.355000  1.460000 ;
      RECT 1469.015000  1.460000 1472.640000  1.600000 ;
      RECT 1469.015000  1.600000 1469.355000  1.645000 ;
      RECT 1469.985000  1.075000 1470.275000  1.120000 ;
      RECT 1469.985000  1.260000 1470.275000  1.305000 ;
      RECT 1471.465000  1.755000 1471.805000  1.800000 ;
      RECT 1471.465000  1.800000 1475.890000  1.940000 ;
      RECT 1471.465000  1.940000 1471.805000  1.985000 ;
      RECT 1471.975000  1.070000 1472.265000  1.120000 ;
      RECT 1471.975000  1.120000 1476.730000  1.260000 ;
      RECT 1471.975000  1.260000 1472.265000  1.300000 ;
      RECT 1472.350000  1.415000 1472.640000  1.460000 ;
      RECT 1472.350000  1.600000 1472.640000  1.645000 ;
      RECT 1472.945000  1.755000 1473.285000  1.800000 ;
      RECT 1472.945000  1.940000 1473.285000  1.985000 ;
      RECT 1474.775000  1.415000 1475.115000  1.460000 ;
      RECT 1474.775000  1.460000 1477.305000  1.600000 ;
      RECT 1474.775000  1.600000 1475.115000  1.645000 ;
      RECT 1475.550000  1.755000 1475.890000  1.800000 ;
      RECT 1475.550000  1.940000 1475.890000  1.985000 ;
      RECT 1476.340000  1.075000 1476.730000  1.120000 ;
      RECT 1476.340000  1.260000 1476.730000  1.305000 ;
      RECT 1476.965000  1.415000 1477.305000  1.460000 ;
      RECT 1476.965000  1.600000 1477.305000  1.645000 ;
      RECT 1481.780000  1.075000 1482.070000  1.120000 ;
      RECT 1481.780000  1.120000 1484.075000  1.260000 ;
      RECT 1481.780000  1.260000 1482.070000  1.305000 ;
      RECT 1482.815000  1.415000 1483.155000  1.460000 ;
      RECT 1482.815000  1.460000 1486.440000  1.600000 ;
      RECT 1482.815000  1.600000 1483.155000  1.645000 ;
      RECT 1483.785000  1.075000 1484.075000  1.120000 ;
      RECT 1483.785000  1.260000 1484.075000  1.305000 ;
      RECT 1485.265000  1.755000 1485.605000  1.800000 ;
      RECT 1485.265000  1.800000 1489.690000  1.940000 ;
      RECT 1485.265000  1.940000 1485.605000  1.985000 ;
      RECT 1485.775000  1.070000 1486.065000  1.120000 ;
      RECT 1485.775000  1.120000 1490.760000  1.260000 ;
      RECT 1485.775000  1.260000 1486.065000  1.300000 ;
      RECT 1486.150000  1.415000 1486.440000  1.460000 ;
      RECT 1486.150000  1.600000 1486.440000  1.645000 ;
      RECT 1486.745000  1.755000 1487.085000  1.800000 ;
      RECT 1486.745000  1.940000 1487.085000  1.985000 ;
      RECT 1488.575000  1.415000 1488.915000  1.460000 ;
      RECT 1488.575000  1.460000 1491.270000  1.600000 ;
      RECT 1488.575000  1.600000 1488.915000  1.645000 ;
      RECT 1489.350000  1.755000 1489.690000  1.800000 ;
      RECT 1489.350000  1.940000 1489.690000  1.985000 ;
      RECT 1490.370000  1.075000 1490.760000  1.120000 ;
      RECT 1490.370000  1.260000 1490.760000  1.305000 ;
      RECT 1490.930000  1.415000 1491.270000  1.460000 ;
      RECT 1490.930000  1.600000 1491.270000  1.645000 ;
      RECT 1496.500000  1.075000 1496.790000  1.120000 ;
      RECT 1496.500000  1.120000 1498.795000  1.260000 ;
      RECT 1496.500000  1.260000 1496.790000  1.305000 ;
      RECT 1497.535000  1.415000 1497.875000  1.460000 ;
      RECT 1497.535000  1.460000 1501.160000  1.600000 ;
      RECT 1497.535000  1.600000 1497.875000  1.645000 ;
      RECT 1498.505000  1.075000 1498.795000  1.120000 ;
      RECT 1498.505000  1.260000 1498.795000  1.305000 ;
      RECT 1499.985000  1.755000 1500.325000  1.800000 ;
      RECT 1499.985000  1.800000 1504.410000  1.940000 ;
      RECT 1499.985000  1.940000 1500.325000  1.985000 ;
      RECT 1500.495000  1.070000 1500.785000  1.120000 ;
      RECT 1500.495000  1.120000 1505.480000  1.260000 ;
      RECT 1500.495000  1.260000 1500.785000  1.300000 ;
      RECT 1500.870000  1.415000 1501.160000  1.460000 ;
      RECT 1500.870000  1.600000 1501.160000  1.645000 ;
      RECT 1501.465000  1.755000 1501.805000  1.800000 ;
      RECT 1501.465000  1.940000 1501.805000  1.985000 ;
      RECT 1503.295000  1.415000 1503.635000  1.460000 ;
      RECT 1503.295000  1.460000 1505.990000  1.600000 ;
      RECT 1503.295000  1.600000 1503.635000  1.645000 ;
      RECT 1504.070000  1.755000 1504.410000  1.800000 ;
      RECT 1504.070000  1.940000 1504.410000  1.985000 ;
      RECT 1505.090000  1.075000 1505.480000  1.120000 ;
      RECT 1505.090000  1.260000 1505.480000  1.305000 ;
      RECT 1505.650000  1.415000 1505.990000  1.460000 ;
      RECT 1505.650000  1.600000 1505.990000  1.645000 ;
      RECT 1512.195000  1.755000 1512.485000  1.800000 ;
      RECT 1512.195000  1.800000 1518.965000  1.940000 ;
      RECT 1512.195000  1.940000 1512.485000  1.985000 ;
      RECT 1512.565000  0.395000 1512.905000  0.440000 ;
      RECT 1512.565000  0.440000 1516.845000  0.580000 ;
      RECT 1512.565000  0.580000 1512.905000  0.625000 ;
      RECT 1516.705000  0.580000 1516.845000  0.735000 ;
      RECT 1516.705000  0.735000 1516.995000  0.780000 ;
      RECT 1516.705000  0.780000 1518.975000  0.920000 ;
      RECT 1516.705000  0.920000 1516.995000  0.965000 ;
      RECT 1517.115000  1.755000 1517.405000  1.800000 ;
      RECT 1517.115000  1.940000 1517.405000  1.985000 ;
      RECT 1518.675000  1.755000 1518.965000  1.800000 ;
      RECT 1518.675000  1.940000 1518.965000  1.985000 ;
      RECT 1518.685000  0.735000 1518.975000  0.780000 ;
      RECT 1518.685000  0.920000 1518.975000  0.965000 ;
      RECT 1524.615000  1.755000 1524.905000  1.800000 ;
      RECT 1524.615000  1.800000 1531.385000  1.940000 ;
      RECT 1524.615000  1.940000 1524.905000  1.985000 ;
      RECT 1524.985000  0.395000 1525.325000  0.440000 ;
      RECT 1524.985000  0.440000 1529.205000  0.580000 ;
      RECT 1524.985000  0.580000 1525.325000  0.625000 ;
      RECT 1529.065000  0.580000 1529.205000  0.735000 ;
      RECT 1529.065000  0.735000 1529.355000  0.780000 ;
      RECT 1529.065000  0.780000 1531.395000  0.920000 ;
      RECT 1529.065000  0.920000 1529.355000  0.965000 ;
      RECT 1529.535000  1.755000 1529.825000  1.800000 ;
      RECT 1529.535000  1.940000 1529.825000  1.985000 ;
      RECT 1531.095000  1.755000 1531.385000  1.800000 ;
      RECT 1531.095000  1.940000 1531.385000  1.985000 ;
      RECT 1531.105000  0.735000 1531.395000  0.780000 ;
      RECT 1531.105000  0.920000 1531.395000  0.965000 ;
      RECT 1538.385000  1.710000 1538.675000  1.800000 ;
      RECT 1538.385000  1.800000 1545.250000  1.940000 ;
      RECT 1538.875000  0.690000 1539.165000  0.780000 ;
      RECT 1538.875000  0.780000 1545.320000  0.920000 ;
      RECT 1542.825000  0.690000 1543.165000  0.780000 ;
      RECT 1543.335000  1.710000 1543.675000  1.800000 ;
      RECT 1544.910000  1.710000 1545.250000  1.800000 ;
      RECT 1545.010000  0.690000 1545.320000  0.780000 ;
      RECT 1549.425000  1.710000 1549.715000  1.800000 ;
      RECT 1549.425000  1.800000 1556.275000  1.940000 ;
      RECT 1549.915000  0.690000 1550.205000  0.780000 ;
      RECT 1549.915000  0.780000 1556.275000  0.920000 ;
      RECT 1553.865000  0.690000 1554.205000  0.780000 ;
      RECT 1554.375000  1.710000 1554.715000  1.800000 ;
      RECT 1555.935000  0.690000 1556.275000  0.780000 ;
      RECT 1555.935000  1.710000 1556.275000  1.800000 ;
      RECT 1560.925000  1.710000 1561.215000  1.800000 ;
      RECT 1560.925000  1.800000 1567.775000  1.940000 ;
      RECT 1561.415000  0.690000 1561.705000  0.780000 ;
      RECT 1561.415000  0.780000 1567.775000  0.920000 ;
      RECT 1565.365000  0.690000 1565.705000  0.780000 ;
      RECT 1565.875000  1.710000 1566.215000  1.800000 ;
      RECT 1567.435000  0.690000 1567.775000  0.780000 ;
      RECT 1567.435000  1.710000 1567.775000  1.800000 ;
      RECT 1574.305000  1.415000 1574.595000  1.460000 ;
      RECT 1574.305000  1.460000 1577.335000  1.600000 ;
      RECT 1574.305000  1.600000 1574.595000  1.645000 ;
      RECT 1574.815000  0.735000 1575.105000  0.780000 ;
      RECT 1574.815000  0.780000 1576.770000  0.920000 ;
      RECT 1574.815000  0.920000 1575.105000  0.965000 ;
      RECT 1576.480000  0.735000 1576.770000  0.780000 ;
      RECT 1576.480000  0.920000 1576.770000  0.965000 ;
      RECT 1577.045000  1.415000 1577.335000  1.460000 ;
      RECT 1577.045000  1.600000 1577.335000  1.645000 ;
      RECT 1577.485000  1.075000 1577.775000  1.120000 ;
      RECT 1577.485000  1.120000 1578.970000  1.260000 ;
      RECT 1577.485000  1.260000 1577.775000  1.305000 ;
      RECT 1578.680000  1.075000 1578.970000  1.120000 ;
      RECT 1578.680000  1.260000 1578.970000  1.305000 ;
      RECT 1582.125000  1.415000 1582.415000  1.460000 ;
      RECT 1582.125000  1.460000 1585.290000  1.600000 ;
      RECT 1582.125000  1.600000 1582.415000  1.645000 ;
      RECT 1582.635000  0.735000 1582.925000  0.780000 ;
      RECT 1582.635000  0.780000 1584.780000  0.920000 ;
      RECT 1582.635000  0.920000 1582.925000  0.965000 ;
      RECT 1584.490000  0.735000 1584.780000  0.780000 ;
      RECT 1584.490000  0.920000 1584.780000  0.965000 ;
      RECT 1585.000000  1.415000 1585.290000  1.460000 ;
      RECT 1585.000000  1.600000 1585.290000  1.645000 ;
      RECT 1585.510000  1.075000 1585.800000  1.120000 ;
      RECT 1585.510000  1.120000 1586.790000  1.260000 ;
      RECT 1585.510000  1.260000 1585.800000  1.305000 ;
      RECT 1586.500000  1.075000 1586.790000  1.120000 ;
      RECT 1586.500000  1.260000 1586.790000  1.305000 ;
      RECT 1590.460000  1.415000 1590.750000  1.460000 ;
      RECT 1590.460000  1.460000 1593.730000  1.600000 ;
      RECT 1590.460000  1.600000 1590.750000  1.645000 ;
      RECT 1590.970000  0.735000 1591.260000  0.780000 ;
      RECT 1590.970000  0.780000 1593.220000  0.920000 ;
      RECT 1590.970000  0.920000 1591.260000  0.965000 ;
      RECT 1592.930000  0.735000 1593.220000  0.780000 ;
      RECT 1592.930000  0.920000 1593.220000  0.965000 ;
      RECT 1593.440000  1.415000 1593.730000  1.460000 ;
      RECT 1593.440000  1.600000 1593.730000  1.645000 ;
      RECT 1593.895000  1.075000 1594.185000  1.120000 ;
      RECT 1593.895000  1.120000 1595.230000  1.260000 ;
      RECT 1593.895000  1.260000 1594.185000  1.305000 ;
      RECT 1594.940000  1.075000 1595.230000  1.120000 ;
      RECT 1594.940000  1.260000 1595.230000  1.305000 ;
      RECT 1599.125000  1.755000 1599.415000  1.800000 ;
      RECT 1599.125000  1.800000 1609.915000  1.940000 ;
      RECT 1599.125000  1.940000 1599.415000  1.985000 ;
      RECT 1599.505000  1.415000 1599.845000  1.460000 ;
      RECT 1599.505000  1.460000 1610.385000  1.600000 ;
      RECT 1599.505000  1.600000 1599.845000  1.645000 ;
      RECT 1599.895000  0.395000 1603.265000  0.580000 ;
      RECT 1599.895000  0.580000 1600.185000  0.625000 ;
      RECT 1602.545000  0.735000 1602.835000  0.780000 ;
      RECT 1602.545000  0.780000 1612.430000  0.920000 ;
      RECT 1602.545000  0.920000 1602.835000  0.965000 ;
      RECT 1602.925000  0.580000 1603.265000  0.625000 ;
      RECT 1603.405000  0.395000 1606.045000  0.580000 ;
      RECT 1603.405000  0.580000 1603.745000  0.625000 ;
      RECT 1605.705000  0.580000 1606.045000  0.625000 ;
      RECT 1606.325000  1.415000 1606.665000  1.460000 ;
      RECT 1606.325000  1.600000 1606.665000  1.645000 ;
      RECT 1606.785000  1.755000 1607.125000  1.800000 ;
      RECT 1606.785000  1.940000 1607.125000  1.985000 ;
      RECT 1609.575000  1.755000 1609.915000  1.800000 ;
      RECT 1609.575000  1.940000 1609.915000  1.985000 ;
      RECT 1610.045000  1.415000 1610.385000  1.460000 ;
      RECT 1610.045000  1.600000 1610.385000  1.645000 ;
      RECT 1610.605000  1.075000 1610.895000  1.120000 ;
      RECT 1610.605000  1.120000 1612.925000  1.260000 ;
      RECT 1610.605000  1.260000 1610.895000  1.305000 ;
      RECT 1612.140000  0.735000 1612.430000  0.780000 ;
      RECT 1612.140000  0.920000 1612.430000  0.965000 ;
      RECT 1612.635000  1.075000 1612.925000  1.120000 ;
      RECT 1612.635000  1.260000 1612.925000  1.305000 ;
      RECT 1614.765000  1.755000 1615.055000  1.800000 ;
      RECT 1614.765000  1.800000 1625.555000  1.940000 ;
      RECT 1614.765000  1.940000 1615.055000  1.985000 ;
      RECT 1615.145000  1.415000 1615.485000  1.460000 ;
      RECT 1615.145000  1.460000 1626.025000  1.600000 ;
      RECT 1615.145000  1.600000 1615.485000  1.645000 ;
      RECT 1615.535000  0.395000 1618.905000  0.580000 ;
      RECT 1615.535000  0.580000 1615.825000  0.625000 ;
      RECT 1618.185000  0.735000 1618.475000  0.780000 ;
      RECT 1618.185000  0.780000 1628.815000  0.920000 ;
      RECT 1618.185000  0.920000 1618.475000  0.965000 ;
      RECT 1618.565000  0.580000 1618.905000  0.625000 ;
      RECT 1619.045000  0.395000 1621.685000  0.580000 ;
      RECT 1619.045000  0.580000 1619.385000  0.625000 ;
      RECT 1621.345000  0.580000 1621.685000  0.625000 ;
      RECT 1621.965000  1.415000 1622.305000  1.460000 ;
      RECT 1621.965000  1.600000 1622.305000  1.645000 ;
      RECT 1622.425000  1.755000 1622.765000  1.800000 ;
      RECT 1622.425000  1.940000 1622.765000  1.985000 ;
      RECT 1625.215000  1.755000 1625.555000  1.800000 ;
      RECT 1625.215000  1.940000 1625.555000  1.985000 ;
      RECT 1625.685000  1.415000 1626.025000  1.460000 ;
      RECT 1625.685000  1.600000 1626.025000  1.645000 ;
      RECT 1626.245000  1.755000 1626.535000  1.800000 ;
      RECT 1626.245000  1.800000 1628.355000  1.940000 ;
      RECT 1626.245000  1.940000 1626.535000  1.985000 ;
      RECT 1628.065000  1.755000 1628.355000  1.800000 ;
      RECT 1628.065000  1.940000 1628.355000  1.985000 ;
      RECT 1628.525000  0.735000 1628.815000  0.780000 ;
      RECT 1628.525000  0.920000 1628.815000  0.965000 ;
      RECT 1637.905000  2.095000 1638.195000  2.140000 ;
      RECT 1637.905000  2.140000 1639.215000  2.280000 ;
      RECT 1637.905000  2.280000 1638.195000  2.325000 ;
      RECT 1638.925000  2.095000 1639.215000  2.140000 ;
      RECT 1638.925000  2.280000 1639.215000  2.325000 ;
      RECT 1643.255000  1.415000 1643.595000  1.460000 ;
      RECT 1643.255000  1.460000 1649.205000  1.600000 ;
      RECT 1643.255000  1.600000 1643.595000  1.645000 ;
      RECT 1648.855000  1.415000 1649.205000  1.460000 ;
      RECT 1648.855000  1.600000 1649.205000  1.645000 ;
      RECT 1656.745000  1.415000 1657.035000  1.460000 ;
      RECT 1656.745000  1.460000 1659.485000  1.600000 ;
      RECT 1656.745000  1.600000 1657.035000  1.645000 ;
      RECT 1657.715000  0.735000 1658.005000  0.780000 ;
      RECT 1657.715000  0.780000 1660.965000  0.920000 ;
      RECT 1657.715000  0.920000 1658.005000  0.965000 ;
      RECT 1658.225000  0.395000 1658.515000  0.440000 ;
      RECT 1658.225000  0.440000 1661.475000  0.580000 ;
      RECT 1658.225000  0.580000 1658.515000  0.625000 ;
      RECT 1659.195000  0.735000 1659.485000  0.780000 ;
      RECT 1659.195000  0.920000 1659.485000  0.965000 ;
      RECT 1659.195000  1.415000 1659.485000  1.460000 ;
      RECT 1659.195000  1.600000 1659.485000  1.645000 ;
      RECT 1660.675000  0.735000 1660.965000  0.780000 ;
      RECT 1660.675000  0.920000 1660.965000  0.965000 ;
      RECT 1661.185000  0.395000 1661.475000  0.440000 ;
      RECT 1661.185000  0.580000 1661.475000  0.625000 ;
      RECT 1666.915000  1.415000 1667.205000  1.460000 ;
      RECT 1666.915000  1.460000 1669.655000  1.600000 ;
      RECT 1666.915000  1.600000 1667.205000  1.645000 ;
      RECT 1667.885000  0.735000 1668.175000  0.780000 ;
      RECT 1667.885000  0.780000 1671.135000  0.920000 ;
      RECT 1667.885000  0.920000 1668.175000  0.965000 ;
      RECT 1668.395000  0.395000 1668.685000  0.440000 ;
      RECT 1668.395000  0.440000 1671.645000  0.580000 ;
      RECT 1668.395000  0.580000 1668.685000  0.625000 ;
      RECT 1669.365000  0.735000 1669.655000  0.780000 ;
      RECT 1669.365000  0.920000 1669.655000  0.965000 ;
      RECT 1669.365000  1.415000 1669.655000  1.460000 ;
      RECT 1669.365000  1.600000 1669.655000  1.645000 ;
      RECT 1670.845000  0.735000 1671.135000  0.780000 ;
      RECT 1670.845000  0.920000 1671.135000  0.965000 ;
      RECT 1671.355000  0.395000 1671.645000  0.440000 ;
      RECT 1671.355000  0.580000 1671.645000  0.625000 ;
      RECT 1678.055000  1.415000 1678.345000  1.460000 ;
      RECT 1678.055000  1.460000 1680.795000  1.600000 ;
      RECT 1678.055000  1.600000 1678.345000  1.645000 ;
      RECT 1679.025000  0.735000 1679.315000  0.780000 ;
      RECT 1679.025000  0.780000 1682.275000  0.920000 ;
      RECT 1679.025000  0.920000 1679.315000  0.965000 ;
      RECT 1679.495000  0.395000 1679.795000  0.440000 ;
      RECT 1679.495000  0.440000 1682.785000  0.580000 ;
      RECT 1679.495000  0.580000 1679.795000  0.625000 ;
      RECT 1680.505000  0.735000 1680.795000  0.780000 ;
      RECT 1680.505000  0.920000 1680.795000  0.965000 ;
      RECT 1680.505000  1.415000 1680.795000  1.460000 ;
      RECT 1680.505000  1.600000 1680.795000  1.645000 ;
      RECT 1681.985000  0.735000 1682.275000  0.780000 ;
      RECT 1681.985000  0.920000 1682.275000  0.965000 ;
      RECT 1682.495000  0.395000 1682.785000  0.440000 ;
      RECT 1682.495000  0.580000 1682.785000  0.625000 ;
      RECT 1688.745000  2.095000 1689.035000  2.140000 ;
      RECT 1688.745000  2.140000 1690.055000  2.280000 ;
      RECT 1688.745000  2.280000 1689.035000  2.325000 ;
      RECT 1689.765000  1.075000 1690.055000  1.120000 ;
      RECT 1689.765000  1.120000 1692.715000  1.260000 ;
      RECT 1689.765000  1.260000 1690.055000  1.305000 ;
      RECT 1689.765000  2.095000 1690.055000  2.140000 ;
      RECT 1689.765000  2.280000 1690.055000  2.325000 ;
      RECT 1692.425000  1.075000 1692.715000  1.120000 ;
      RECT 1692.425000  1.260000 1692.715000  1.305000 ;
      RECT 1697.685000  1.415000 1697.975000  1.460000 ;
      RECT 1697.685000  1.460000 1704.095000  1.600000 ;
      RECT 1697.685000  1.600000 1697.975000  1.645000 ;
      RECT 1701.205000  0.695000 1701.495000  0.780000 ;
      RECT 1701.205000  0.780000 1704.555000  0.925000 ;
      RECT 1703.805000  1.415000 1704.095000  1.460000 ;
      RECT 1703.805000  1.600000 1704.095000  1.645000 ;
      RECT 1704.265000  0.695000 1704.555000  0.780000 ;
      RECT 1710.565000  1.415000 1710.855000  1.460000 ;
      RECT 1710.565000  1.460000 1713.305000  1.600000 ;
      RECT 1710.565000  1.600000 1710.855000  1.645000 ;
      RECT 1711.535000  0.735000 1711.825000  0.780000 ;
      RECT 1711.535000  0.780000 1714.785000  0.920000 ;
      RECT 1711.535000  0.920000 1711.825000  0.965000 ;
      RECT 1712.045000  0.395000 1712.335000  0.440000 ;
      RECT 1712.045000  0.440000 1715.295000  0.580000 ;
      RECT 1712.045000  0.580000 1712.335000  0.625000 ;
      RECT 1713.015000  0.735000 1713.305000  0.780000 ;
      RECT 1713.015000  0.920000 1713.305000  0.965000 ;
      RECT 1713.015000  1.415000 1713.305000  1.460000 ;
      RECT 1713.015000  1.600000 1713.305000  1.645000 ;
      RECT 1714.495000  0.735000 1714.785000  0.780000 ;
      RECT 1714.495000  0.920000 1714.785000  0.965000 ;
      RECT 1715.005000  0.395000 1715.295000  0.440000 ;
      RECT 1715.005000  0.580000 1715.295000  0.625000 ;
      RECT 1720.980000  1.415000 1721.270000  1.460000 ;
      RECT 1720.980000  1.460000 1723.720000  1.600000 ;
      RECT 1720.980000  1.600000 1721.270000  1.645000 ;
      RECT 1721.950000  0.735000 1722.240000  0.780000 ;
      RECT 1721.950000  0.780000 1725.200000  0.920000 ;
      RECT 1721.950000  0.920000 1722.240000  0.965000 ;
      RECT 1722.460000  0.395000 1722.750000  0.440000 ;
      RECT 1722.460000  0.440000 1725.710000  0.580000 ;
      RECT 1722.460000  0.580000 1722.750000  0.625000 ;
      RECT 1723.430000  0.735000 1723.720000  0.780000 ;
      RECT 1723.430000  0.920000 1723.720000  0.965000 ;
      RECT 1723.430000  1.415000 1723.720000  1.460000 ;
      RECT 1723.430000  1.600000 1723.720000  1.645000 ;
      RECT 1724.910000  0.735000 1725.200000  0.780000 ;
      RECT 1724.910000  0.920000 1725.200000  0.965000 ;
      RECT 1725.420000  0.395000 1725.710000  0.440000 ;
      RECT 1725.420000  0.580000 1725.710000  0.625000 ;
      RECT 1731.975000  1.415000 1732.265000  1.460000 ;
      RECT 1731.975000  1.460000 1734.715000  1.600000 ;
      RECT 1731.975000  1.600000 1732.265000  1.645000 ;
      RECT 1732.945000  0.735000 1733.285000  0.780000 ;
      RECT 1732.945000  0.780000 1736.195000  0.920000 ;
      RECT 1732.945000  0.920000 1733.285000  0.965000 ;
      RECT 1733.455000  0.395000 1733.745000  0.440000 ;
      RECT 1733.455000  0.440000 1736.705000  0.580000 ;
      RECT 1733.455000  0.580000 1733.745000  0.625000 ;
      RECT 1734.425000  0.735000 1734.715000  0.780000 ;
      RECT 1734.425000  0.920000 1734.715000  0.965000 ;
      RECT 1734.425000  1.415000 1734.715000  1.460000 ;
      RECT 1734.425000  1.600000 1734.715000  1.645000 ;
      RECT 1735.905000  0.735000 1736.195000  0.780000 ;
      RECT 1735.905000  0.920000 1736.195000  0.965000 ;
      RECT 1736.415000  0.395000 1736.705000  0.440000 ;
      RECT 1736.415000  0.580000 1736.705000  0.625000 ;
      RECT 1739.135000  1.075000 1739.425000  1.120000 ;
      RECT 1739.135000  1.120000 1747.805000  1.260000 ;
      RECT 1739.135000  1.260000 1739.425000  1.305000 ;
      RECT 1739.410000  1.755000 1739.710000  1.800000 ;
      RECT 1739.410000  1.800000 1748.135000  1.940000 ;
      RECT 1739.410000  1.940000 1739.710000  1.985000 ;
      RECT 1743.760000  1.075000 1744.050000  1.120000 ;
      RECT 1743.760000  1.260000 1744.050000  1.305000 ;
      RECT 1744.230000  1.755000 1744.520000  1.800000 ;
      RECT 1744.230000  1.940000 1744.520000  1.985000 ;
      RECT 1745.485000  0.735000 1746.240000  0.780000 ;
      RECT 1745.485000  0.780000 1749.745000  0.920000 ;
      RECT 1745.485000  0.920000 1746.240000  0.965000 ;
      RECT 1747.495000  1.075000 1747.805000  1.120000 ;
      RECT 1747.495000  1.260000 1747.805000  1.305000 ;
      RECT 1747.840000  1.755000 1748.135000  1.800000 ;
      RECT 1747.840000  1.940000 1748.135000  1.985000 ;
      RECT 1749.115000  0.920000 1749.745000  0.965000 ;
      RECT 1749.115000  0.965000 1749.405000  1.310000 ;
      RECT 1749.455000  0.735000 1749.745000  0.780000 ;
      RECT 1834.105000  1.755000 1834.395000  1.800000 ;
      RECT 1834.105000  1.800000 1840.835000  1.940000 ;
      RECT 1834.105000  1.940000 1834.395000  1.985000 ;
      RECT 1836.405000  1.755000 1836.695000  1.800000 ;
      RECT 1836.405000  1.940000 1836.695000  1.985000 ;
      RECT 1838.245000  1.755000 1838.535000  1.800000 ;
      RECT 1838.245000  1.940000 1838.535000  1.985000 ;
      RECT 1840.545000  1.755000 1840.835000  1.800000 ;
      RECT 1840.545000  1.940000 1840.835000  1.985000 ;
      RECT 1843.765000  1.755000 1844.055000  1.800000 ;
      RECT 1843.765000  1.800000 1853.715000  1.940000 ;
      RECT 1843.765000  1.940000 1844.055000  1.985000 ;
      RECT 1846.985000  1.755000 1847.275000  1.800000 ;
      RECT 1846.985000  1.940000 1847.275000  1.985000 ;
      RECT 1850.205000  1.755000 1850.495000  1.800000 ;
      RECT 1850.205000  1.940000 1850.495000  1.985000 ;
      RECT 1853.425000  1.755000 1853.715000  1.800000 ;
      RECT 1853.425000  1.940000 1853.715000  1.985000 ;
      RECT 1858.625000  1.755000 1858.915000  1.800000 ;
      RECT 1858.625000  1.800000 1878.415000  1.940000 ;
      RECT 1858.625000  1.940000 1858.915000  1.985000 ;
      RECT 1859.565000  1.755000 1859.855000  1.800000 ;
      RECT 1859.565000  1.940000 1859.855000  1.985000 ;
      RECT 1864.305000  1.755000 1864.595000  1.800000 ;
      RECT 1864.305000  1.940000 1864.595000  1.985000 ;
      RECT 1865.245000  1.755000 1865.535000  1.800000 ;
      RECT 1865.245000  1.940000 1865.535000  1.985000 ;
      RECT 1871.505000  1.755000 1871.795000  1.800000 ;
      RECT 1871.505000  1.940000 1871.795000  1.985000 ;
      RECT 1872.445000  1.755000 1872.735000  1.800000 ;
      RECT 1872.445000  1.940000 1872.735000  1.985000 ;
      RECT 1877.185000  1.755000 1877.475000  1.800000 ;
      RECT 1877.185000  1.940000 1877.475000  1.985000 ;
      RECT 1878.125000  1.755000 1878.415000  1.800000 ;
      RECT 1878.125000  1.940000 1878.415000  1.985000 ;
      RECT 1882.865000  1.755000 1883.155000  1.800000 ;
      RECT 1882.865000  1.800000 1897.875000  1.940000 ;
      RECT 1882.865000  1.940000 1883.155000  1.985000 ;
      RECT 1885.165000  1.755000 1885.455000  1.800000 ;
      RECT 1885.165000  1.940000 1885.455000  1.985000 ;
      RECT 1887.005000  1.755000 1887.295000  1.800000 ;
      RECT 1887.005000  1.940000 1887.295000  1.985000 ;
      RECT 1889.305000  1.755000 1889.595000  1.800000 ;
      RECT 1889.305000  1.940000 1889.595000  1.985000 ;
      RECT 1891.145000  1.755000 1891.435000  1.800000 ;
      RECT 1891.145000  1.940000 1891.435000  1.985000 ;
      RECT 1893.445000  1.755000 1893.735000  1.800000 ;
      RECT 1893.445000  1.940000 1893.735000  1.985000 ;
      RECT 1895.285000  1.755000 1895.575000  1.800000 ;
      RECT 1895.285000  1.940000 1895.575000  1.985000 ;
      RECT 1897.585000  1.755000 1897.875000  1.800000 ;
      RECT 1897.585000  1.940000 1897.875000  1.985000 ;
      RECT 1900.805000  1.755000 1901.095000  1.800000 ;
      RECT 1900.805000  1.800000 1923.635000  1.940000 ;
      RECT 1900.805000  1.940000 1901.095000  1.985000 ;
      RECT 1904.025000  1.755000 1904.315000  1.800000 ;
      RECT 1904.025000  1.940000 1904.315000  1.985000 ;
      RECT 1907.245000  1.755000 1907.535000  1.800000 ;
      RECT 1907.245000  1.940000 1907.535000  1.985000 ;
      RECT 1910.465000  1.755000 1910.755000  1.800000 ;
      RECT 1910.465000  1.940000 1910.755000  1.985000 ;
      RECT 1913.685000  1.755000 1913.975000  1.800000 ;
      RECT 1913.685000  1.940000 1913.975000  1.985000 ;
      RECT 1916.905000  1.755000 1917.195000  1.800000 ;
      RECT 1916.905000  1.940000 1917.195000  1.985000 ;
      RECT 1920.125000  1.755000 1920.415000  1.800000 ;
      RECT 1920.125000  1.940000 1920.415000  1.985000 ;
      RECT 1923.345000  1.755000 1923.635000  1.800000 ;
      RECT 1923.345000  1.940000 1923.635000  1.985000 ;
      RECT 1942.120000  5.200000 2064.020000  5.370000 ;
      RECT 1942.120000  5.370000 2064.400000  5.510000 ;
      RECT 1942.120000  5.510000 2064.020000  5.680000 ;
      RECT 1944.325000  2.110000 1944.615000  2.155000 ;
      RECT 1944.325000  2.155000 1948.435000  2.295000 ;
      RECT 1944.325000  2.295000 1944.615000  2.340000 ;
      RECT 1944.325000  3.100000 1944.615000  3.145000 ;
      RECT 1944.325000  3.145000 1948.435000  3.285000 ;
      RECT 1944.325000  3.285000 1944.615000  3.330000 ;
      RECT 1944.805000  1.755000 1945.095000  1.800000 ;
      RECT 1944.805000  1.800000 1965.195000  1.940000 ;
      RECT 1944.805000  1.940000 1945.095000  1.985000 ;
      RECT 1944.805000  3.455000 1945.095000  3.500000 ;
      RECT 1944.805000  3.500000 1965.195000  3.640000 ;
      RECT 1944.805000  3.640000 1945.095000  3.685000 ;
      RECT 1945.275000  2.110000 1945.565000  2.155000 ;
      RECT 1945.275000  2.295000 1945.565000  2.340000 ;
      RECT 1945.275000  3.100000 1945.565000  3.145000 ;
      RECT 1945.275000  3.285000 1945.565000  3.330000 ;
      RECT 1945.745000  1.755000 1946.035000  1.800000 ;
      RECT 1945.745000  1.940000 1946.035000  1.985000 ;
      RECT 1945.745000  3.455000 1946.035000  3.500000 ;
      RECT 1945.745000  3.640000 1946.035000  3.685000 ;
      RECT 1946.225000  2.110000 1946.515000  2.155000 ;
      RECT 1946.225000  2.295000 1946.515000  2.340000 ;
      RECT 1946.225000  3.100000 1946.515000  3.145000 ;
      RECT 1946.225000  3.285000 1946.515000  3.330000 ;
      RECT 1947.205000  2.110000 1947.495000  2.155000 ;
      RECT 1947.205000  2.295000 1947.495000  2.340000 ;
      RECT 1947.205000  3.100000 1947.495000  3.145000 ;
      RECT 1947.205000  3.285000 1947.495000  3.330000 ;
      RECT 1948.145000  2.110000 1948.435000  2.155000 ;
      RECT 1948.145000  2.295000 1948.435000  2.340000 ;
      RECT 1948.145000  3.100000 1948.435000  3.145000 ;
      RECT 1948.145000  3.285000 1948.435000  3.330000 ;
      RECT 1949.145000  2.110000 1949.435000  2.155000 ;
      RECT 1949.145000  2.155000 1953.255000  2.295000 ;
      RECT 1949.145000  2.295000 1949.435000  2.340000 ;
      RECT 1949.145000  3.100000 1949.435000  3.145000 ;
      RECT 1949.145000  3.145000 1953.255000  3.285000 ;
      RECT 1949.145000  3.285000 1949.435000  3.330000 ;
      RECT 1950.085000  2.110000 1950.375000  2.155000 ;
      RECT 1950.085000  2.295000 1950.375000  2.340000 ;
      RECT 1950.085000  3.100000 1950.375000  3.145000 ;
      RECT 1950.085000  3.285000 1950.375000  3.330000 ;
      RECT 1951.065000  2.110000 1951.355000  2.155000 ;
      RECT 1951.065000  2.295000 1951.355000  2.340000 ;
      RECT 1951.065000  3.100000 1951.355000  3.145000 ;
      RECT 1951.065000  3.285000 1951.355000  3.330000 ;
      RECT 1951.545000  1.755000 1951.835000  1.800000 ;
      RECT 1951.545000  1.940000 1951.835000  1.985000 ;
      RECT 1951.545000  3.455000 1951.835000  3.500000 ;
      RECT 1951.545000  3.640000 1951.835000  3.685000 ;
      RECT 1952.015000  2.110000 1952.305000  2.155000 ;
      RECT 1952.015000  2.295000 1952.305000  2.340000 ;
      RECT 1952.015000  3.100000 1952.305000  3.145000 ;
      RECT 1952.015000  3.285000 1952.305000  3.330000 ;
      RECT 1952.485000  1.755000 1952.775000  1.800000 ;
      RECT 1952.485000  1.940000 1952.775000  1.985000 ;
      RECT 1952.485000  3.455000 1952.775000  3.500000 ;
      RECT 1952.485000  3.640000 1952.775000  3.685000 ;
      RECT 1952.965000  2.110000 1953.255000  2.155000 ;
      RECT 1952.965000  2.295000 1953.255000  2.340000 ;
      RECT 1952.965000  3.100000 1953.255000  3.145000 ;
      RECT 1952.965000  3.285000 1953.255000  3.330000 ;
      RECT 1956.745000  2.110000 1957.035000  2.155000 ;
      RECT 1956.745000  2.155000 1960.855000  2.295000 ;
      RECT 1956.745000  2.295000 1957.035000  2.340000 ;
      RECT 1956.745000  3.100000 1957.035000  3.145000 ;
      RECT 1956.745000  3.145000 1960.855000  3.285000 ;
      RECT 1956.745000  3.285000 1957.035000  3.330000 ;
      RECT 1957.225000  1.755000 1957.515000  1.800000 ;
      RECT 1957.225000  1.940000 1957.515000  1.985000 ;
      RECT 1957.225000  3.455000 1957.515000  3.500000 ;
      RECT 1957.225000  3.640000 1957.515000  3.685000 ;
      RECT 1957.695000  2.110000 1957.985000  2.155000 ;
      RECT 1957.695000  2.295000 1957.985000  2.340000 ;
      RECT 1957.695000  3.100000 1957.985000  3.145000 ;
      RECT 1957.695000  3.285000 1957.985000  3.330000 ;
      RECT 1958.165000  1.755000 1958.455000  1.800000 ;
      RECT 1958.165000  1.940000 1958.455000  1.985000 ;
      RECT 1958.165000  3.455000 1958.455000  3.500000 ;
      RECT 1958.165000  3.640000 1958.455000  3.685000 ;
      RECT 1958.645000  2.110000 1958.935000  2.155000 ;
      RECT 1958.645000  2.295000 1958.935000  2.340000 ;
      RECT 1958.645000  3.100000 1958.935000  3.145000 ;
      RECT 1958.645000  3.285000 1958.935000  3.330000 ;
      RECT 1959.625000  2.110000 1959.915000  2.155000 ;
      RECT 1959.625000  2.295000 1959.915000  2.340000 ;
      RECT 1959.625000  3.100000 1959.915000  3.145000 ;
      RECT 1959.625000  3.285000 1959.915000  3.330000 ;
      RECT 1960.565000  2.110000 1960.855000  2.155000 ;
      RECT 1960.565000  2.295000 1960.855000  2.340000 ;
      RECT 1960.565000  3.100000 1960.855000  3.145000 ;
      RECT 1960.565000  3.285000 1960.855000  3.330000 ;
      RECT 1961.565000  2.110000 1961.855000  2.155000 ;
      RECT 1961.565000  2.155000 1965.675000  2.295000 ;
      RECT 1961.565000  2.295000 1961.855000  2.340000 ;
      RECT 1961.565000  3.100000 1961.855000  3.145000 ;
      RECT 1961.565000  3.145000 1965.675000  3.285000 ;
      RECT 1961.565000  3.285000 1961.855000  3.330000 ;
      RECT 1962.505000  2.110000 1962.795000  2.155000 ;
      RECT 1962.505000  2.295000 1962.795000  2.340000 ;
      RECT 1962.505000  3.100000 1962.795000  3.145000 ;
      RECT 1962.505000  3.285000 1962.795000  3.330000 ;
      RECT 1963.485000  2.110000 1963.775000  2.155000 ;
      RECT 1963.485000  2.295000 1963.775000  2.340000 ;
      RECT 1963.485000  3.100000 1963.775000  3.145000 ;
      RECT 1963.485000  3.285000 1963.775000  3.330000 ;
      RECT 1963.965000  1.755000 1964.255000  1.800000 ;
      RECT 1963.965000  1.940000 1964.255000  1.985000 ;
      RECT 1963.965000  3.455000 1964.255000  3.500000 ;
      RECT 1963.965000  3.640000 1964.255000  3.685000 ;
      RECT 1964.435000  2.110000 1964.725000  2.155000 ;
      RECT 1964.435000  2.295000 1964.725000  2.340000 ;
      RECT 1964.435000  3.100000 1964.725000  3.145000 ;
      RECT 1964.435000  3.285000 1964.725000  3.330000 ;
      RECT 1964.905000  1.755000 1965.195000  1.800000 ;
      RECT 1964.905000  1.940000 1965.195000  1.985000 ;
      RECT 1964.905000  3.455000 1965.195000  3.500000 ;
      RECT 1964.905000  3.640000 1965.195000  3.685000 ;
      RECT 1965.385000  2.110000 1965.675000  2.155000 ;
      RECT 1965.385000  2.295000 1965.675000  2.340000 ;
      RECT 1965.385000  3.100000 1965.675000  3.145000 ;
      RECT 1965.385000  3.285000 1965.675000  3.330000 ;
      RECT 1968.885000  1.755000 1969.175000  1.800000 ;
      RECT 1968.885000  1.800000 1983.895000  1.940000 ;
      RECT 1968.885000  1.940000 1969.175000  1.985000 ;
      RECT 1968.885000  3.455000 1969.175000  3.500000 ;
      RECT 1968.885000  3.500000 1983.895000  3.640000 ;
      RECT 1968.885000  3.640000 1969.175000  3.685000 ;
      RECT 1971.185000  1.755000 1971.475000  1.800000 ;
      RECT 1971.185000  1.940000 1971.475000  1.985000 ;
      RECT 1971.185000  3.455000 1971.475000  3.500000 ;
      RECT 1971.185000  3.640000 1971.475000  3.685000 ;
      RECT 1973.025000  1.755000 1973.315000  1.800000 ;
      RECT 1973.025000  1.940000 1973.315000  1.985000 ;
      RECT 1973.025000  3.455000 1973.315000  3.500000 ;
      RECT 1973.025000  3.640000 1973.315000  3.685000 ;
      RECT 1975.325000  1.755000 1975.615000  1.800000 ;
      RECT 1975.325000  1.940000 1975.615000  1.985000 ;
      RECT 1975.325000  3.455000 1975.615000  3.500000 ;
      RECT 1975.325000  3.640000 1975.615000  3.685000 ;
      RECT 1977.165000  1.755000 1977.455000  1.800000 ;
      RECT 1977.165000  1.940000 1977.455000  1.985000 ;
      RECT 1977.165000  3.455000 1977.455000  3.500000 ;
      RECT 1977.165000  3.640000 1977.455000  3.685000 ;
      RECT 1979.465000  1.755000 1979.755000  1.800000 ;
      RECT 1979.465000  1.940000 1979.755000  1.985000 ;
      RECT 1979.465000  3.455000 1979.755000  3.500000 ;
      RECT 1979.465000  3.640000 1979.755000  3.685000 ;
      RECT 1981.305000  1.755000 1981.595000  1.800000 ;
      RECT 1981.305000  1.940000 1981.595000  1.985000 ;
      RECT 1981.305000  3.455000 1981.595000  3.500000 ;
      RECT 1981.305000  3.640000 1981.595000  3.685000 ;
      RECT 1983.605000  1.755000 1983.895000  1.800000 ;
      RECT 1983.605000  1.940000 1983.895000  1.985000 ;
      RECT 1983.605000  3.455000 1983.895000  3.500000 ;
      RECT 1983.605000  3.640000 1983.895000  3.685000 ;
      RECT 1985.475000  2.110000 1985.765000  2.155000 ;
      RECT 1985.475000  2.155000 1987.700000  2.295000 ;
      RECT 1985.475000  2.295000 1985.765000  2.340000 ;
      RECT 1985.475000  3.100000 1985.765000  3.145000 ;
      RECT 1985.475000  3.145000 1987.700000  3.285000 ;
      RECT 1985.475000  3.285000 1985.765000  3.330000 ;
      RECT 1986.415000  2.110000 1986.705000  2.155000 ;
      RECT 1986.415000  2.295000 1986.705000  2.340000 ;
      RECT 1986.415000  3.100000 1986.705000  3.145000 ;
      RECT 1986.415000  3.285000 1986.705000  3.330000 ;
      RECT 1986.825000  1.755000 1987.115000  1.800000 ;
      RECT 1986.825000  1.800000 2009.655000  1.940000 ;
      RECT 1986.825000  1.940000 1987.115000  1.985000 ;
      RECT 1986.825000  3.455000 1987.115000  3.500000 ;
      RECT 1986.825000  3.500000 2009.655000  3.640000 ;
      RECT 1986.825000  3.640000 1987.115000  3.685000 ;
      RECT 1987.410000  2.110000 1987.700000  2.155000 ;
      RECT 1987.410000  2.295000 1987.700000  2.340000 ;
      RECT 1987.410000  3.100000 1987.700000  3.145000 ;
      RECT 1987.410000  3.285000 1987.700000  3.330000 ;
      RECT 1989.460000  2.110000 1989.750000  2.155000 ;
      RECT 1989.460000  2.155000 1991.685000  2.295000 ;
      RECT 1989.460000  2.295000 1989.750000  2.340000 ;
      RECT 1989.460000  3.100000 1989.750000  3.145000 ;
      RECT 1989.460000  3.145000 1991.685000  3.285000 ;
      RECT 1989.460000  3.285000 1989.750000  3.330000 ;
      RECT 1990.045000  1.755000 1990.335000  1.800000 ;
      RECT 1990.045000  1.940000 1990.335000  1.985000 ;
      RECT 1990.045000  3.455000 1990.335000  3.500000 ;
      RECT 1990.045000  3.640000 1990.335000  3.685000 ;
      RECT 1990.455000  2.110000 1990.745000  2.155000 ;
      RECT 1990.455000  2.295000 1990.745000  2.340000 ;
      RECT 1990.455000  3.100000 1990.745000  3.145000 ;
      RECT 1990.455000  3.285000 1990.745000  3.330000 ;
      RECT 1991.395000  2.110000 1991.685000  2.155000 ;
      RECT 1991.395000  2.295000 1991.685000  2.340000 ;
      RECT 1991.395000  3.100000 1991.685000  3.145000 ;
      RECT 1991.395000  3.285000 1991.685000  3.330000 ;
      RECT 1991.915000  2.110000 1992.205000  2.155000 ;
      RECT 1991.915000  2.155000 1994.140000  2.295000 ;
      RECT 1991.915000  2.295000 1992.205000  2.340000 ;
      RECT 1991.915000  3.100000 1992.205000  3.145000 ;
      RECT 1991.915000  3.145000 1994.140000  3.285000 ;
      RECT 1991.915000  3.285000 1992.205000  3.330000 ;
      RECT 1992.855000  2.110000 1993.145000  2.155000 ;
      RECT 1992.855000  2.295000 1993.145000  2.340000 ;
      RECT 1992.855000  3.100000 1993.145000  3.145000 ;
      RECT 1992.855000  3.285000 1993.145000  3.330000 ;
      RECT 1993.265000  1.755000 1993.555000  1.800000 ;
      RECT 1993.265000  1.940000 1993.555000  1.985000 ;
      RECT 1993.265000  3.455000 1993.555000  3.500000 ;
      RECT 1993.265000  3.640000 1993.555000  3.685000 ;
      RECT 1993.850000  2.110000 1994.140000  2.155000 ;
      RECT 1993.850000  2.295000 1994.140000  2.340000 ;
      RECT 1993.850000  3.100000 1994.140000  3.145000 ;
      RECT 1993.850000  3.285000 1994.140000  3.330000 ;
      RECT 1995.900000  2.110000 1996.190000  2.155000 ;
      RECT 1995.900000  2.155000 1998.125000  2.295000 ;
      RECT 1995.900000  2.295000 1996.190000  2.340000 ;
      RECT 1995.900000  3.100000 1996.190000  3.145000 ;
      RECT 1995.900000  3.145000 1998.125000  3.285000 ;
      RECT 1995.900000  3.285000 1996.190000  3.330000 ;
      RECT 1996.485000  1.755000 1996.775000  1.800000 ;
      RECT 1996.485000  1.940000 1996.775000  1.985000 ;
      RECT 1996.485000  3.455000 1996.775000  3.500000 ;
      RECT 1996.485000  3.640000 1996.775000  3.685000 ;
      RECT 1996.895000  2.110000 1997.185000  2.155000 ;
      RECT 1996.895000  2.295000 1997.185000  2.340000 ;
      RECT 1996.895000  3.100000 1997.185000  3.145000 ;
      RECT 1996.895000  3.285000 1997.185000  3.330000 ;
      RECT 1997.835000  2.110000 1998.125000  2.155000 ;
      RECT 1997.835000  2.295000 1998.125000  2.340000 ;
      RECT 1997.835000  3.100000 1998.125000  3.145000 ;
      RECT 1997.835000  3.285000 1998.125000  3.330000 ;
      RECT 1998.355000  2.110000 1998.645000  2.155000 ;
      RECT 1998.355000  2.155000 2000.580000  2.295000 ;
      RECT 1998.355000  2.295000 1998.645000  2.340000 ;
      RECT 1998.355000  3.100000 1998.645000  3.145000 ;
      RECT 1998.355000  3.145000 2000.580000  3.285000 ;
      RECT 1998.355000  3.285000 1998.645000  3.330000 ;
      RECT 1999.295000  2.110000 1999.585000  2.155000 ;
      RECT 1999.295000  2.295000 1999.585000  2.340000 ;
      RECT 1999.295000  3.100000 1999.585000  3.145000 ;
      RECT 1999.295000  3.285000 1999.585000  3.330000 ;
      RECT 1999.705000  1.755000 1999.995000  1.800000 ;
      RECT 1999.705000  1.940000 1999.995000  1.985000 ;
      RECT 1999.705000  3.455000 1999.995000  3.500000 ;
      RECT 1999.705000  3.640000 1999.995000  3.685000 ;
      RECT 2000.290000  2.110000 2000.580000  2.155000 ;
      RECT 2000.290000  2.295000 2000.580000  2.340000 ;
      RECT 2000.290000  3.100000 2000.580000  3.145000 ;
      RECT 2000.290000  3.285000 2000.580000  3.330000 ;
      RECT 2002.340000  2.110000 2002.630000  2.155000 ;
      RECT 2002.340000  2.155000 2004.565000  2.295000 ;
      RECT 2002.340000  2.295000 2002.630000  2.340000 ;
      RECT 2002.340000  3.100000 2002.630000  3.145000 ;
      RECT 2002.340000  3.145000 2004.565000  3.285000 ;
      RECT 2002.340000  3.285000 2002.630000  3.330000 ;
      RECT 2002.925000  1.755000 2003.215000  1.800000 ;
      RECT 2002.925000  1.940000 2003.215000  1.985000 ;
      RECT 2002.925000  3.455000 2003.215000  3.500000 ;
      RECT 2002.925000  3.640000 2003.215000  3.685000 ;
      RECT 2003.335000  2.110000 2003.625000  2.155000 ;
      RECT 2003.335000  2.295000 2003.625000  2.340000 ;
      RECT 2003.335000  3.100000 2003.625000  3.145000 ;
      RECT 2003.335000  3.285000 2003.625000  3.330000 ;
      RECT 2004.275000  2.110000 2004.565000  2.155000 ;
      RECT 2004.275000  2.295000 2004.565000  2.340000 ;
      RECT 2004.275000  3.100000 2004.565000  3.145000 ;
      RECT 2004.275000  3.285000 2004.565000  3.330000 ;
      RECT 2004.795000  2.110000 2005.085000  2.155000 ;
      RECT 2004.795000  2.155000 2007.020000  2.295000 ;
      RECT 2004.795000  2.295000 2005.085000  2.340000 ;
      RECT 2004.795000  3.100000 2005.085000  3.145000 ;
      RECT 2004.795000  3.145000 2007.020000  3.285000 ;
      RECT 2004.795000  3.285000 2005.085000  3.330000 ;
      RECT 2005.735000  2.110000 2006.025000  2.155000 ;
      RECT 2005.735000  2.295000 2006.025000  2.340000 ;
      RECT 2005.735000  3.100000 2006.025000  3.145000 ;
      RECT 2005.735000  3.285000 2006.025000  3.330000 ;
      RECT 2006.145000  1.755000 2006.435000  1.800000 ;
      RECT 2006.145000  1.940000 2006.435000  1.985000 ;
      RECT 2006.145000  3.455000 2006.435000  3.500000 ;
      RECT 2006.145000  3.640000 2006.435000  3.685000 ;
      RECT 2006.730000  2.110000 2007.020000  2.155000 ;
      RECT 2006.730000  2.295000 2007.020000  2.340000 ;
      RECT 2006.730000  3.100000 2007.020000  3.145000 ;
      RECT 2006.730000  3.285000 2007.020000  3.330000 ;
      RECT 2008.780000  2.110000 2009.070000  2.155000 ;
      RECT 2008.780000  2.155000 2011.005000  2.295000 ;
      RECT 2008.780000  2.295000 2009.070000  2.340000 ;
      RECT 2008.780000  3.100000 2009.070000  3.145000 ;
      RECT 2008.780000  3.145000 2011.005000  3.285000 ;
      RECT 2008.780000  3.285000 2009.070000  3.330000 ;
      RECT 2009.365000  1.755000 2009.655000  1.800000 ;
      RECT 2009.365000  1.940000 2009.655000  1.985000 ;
      RECT 2009.365000  3.455000 2009.655000  3.500000 ;
      RECT 2009.365000  3.640000 2009.655000  3.685000 ;
      RECT 2009.775000  2.110000 2010.065000  2.155000 ;
      RECT 2009.775000  2.295000 2010.065000  2.340000 ;
      RECT 2009.775000  3.100000 2010.065000  3.145000 ;
      RECT 2009.775000  3.285000 2010.065000  3.330000 ;
      RECT 2010.715000  2.110000 2011.005000  2.155000 ;
      RECT 2010.715000  2.295000 2011.005000  2.340000 ;
      RECT 2010.715000  3.100000 2011.005000  3.145000 ;
      RECT 2010.715000  3.285000 2011.005000  3.330000 ;
      RECT 2012.165000  2.110000 2012.455000  2.155000 ;
      RECT 2012.165000  2.155000 2016.275000  2.295000 ;
      RECT 2012.165000  2.295000 2012.455000  2.340000 ;
      RECT 2012.165000  3.100000 2012.455000  3.145000 ;
      RECT 2012.165000  3.145000 2016.275000  3.285000 ;
      RECT 2012.165000  3.285000 2012.455000  3.330000 ;
      RECT 2013.105000  2.110000 2013.395000  2.155000 ;
      RECT 2013.105000  2.295000 2013.395000  2.340000 ;
      RECT 2013.105000  3.100000 2013.395000  3.145000 ;
      RECT 2013.105000  3.285000 2013.395000  3.330000 ;
      RECT 2014.085000  2.110000 2014.375000  2.155000 ;
      RECT 2014.085000  2.295000 2014.375000  2.340000 ;
      RECT 2014.085000  3.100000 2014.375000  3.145000 ;
      RECT 2014.085000  3.285000 2014.375000  3.330000 ;
      RECT 2014.565000  1.755000 2014.855000  1.800000 ;
      RECT 2014.565000  1.800000 2060.575000  1.940000 ;
      RECT 2014.565000  1.940000 2014.855000  1.985000 ;
      RECT 2014.565000  3.455000 2014.855000  3.500000 ;
      RECT 2014.565000  3.500000 2060.575000  3.640000 ;
      RECT 2014.565000  3.640000 2014.855000  3.685000 ;
      RECT 2015.035000  2.110000 2015.325000  2.155000 ;
      RECT 2015.035000  2.295000 2015.325000  2.340000 ;
      RECT 2015.035000  3.100000 2015.325000  3.145000 ;
      RECT 2015.035000  3.285000 2015.325000  3.330000 ;
      RECT 2015.505000  1.755000 2015.795000  1.800000 ;
      RECT 2015.505000  1.940000 2015.795000  1.985000 ;
      RECT 2015.505000  3.455000 2015.795000  3.500000 ;
      RECT 2015.505000  3.640000 2015.795000  3.685000 ;
      RECT 2015.985000  2.110000 2016.275000  2.155000 ;
      RECT 2015.985000  2.295000 2016.275000  2.340000 ;
      RECT 2015.985000  3.100000 2016.275000  3.145000 ;
      RECT 2015.985000  3.285000 2016.275000  3.330000 ;
      RECT 2019.765000  2.110000 2020.055000  2.155000 ;
      RECT 2019.765000  2.155000 2023.875000  2.295000 ;
      RECT 2019.765000  2.295000 2020.055000  2.340000 ;
      RECT 2019.765000  3.100000 2020.055000  3.145000 ;
      RECT 2019.765000  3.145000 2023.875000  3.285000 ;
      RECT 2019.765000  3.285000 2020.055000  3.330000 ;
      RECT 2020.245000  1.755000 2020.535000  1.800000 ;
      RECT 2020.245000  1.940000 2020.535000  1.985000 ;
      RECT 2020.245000  3.455000 2020.535000  3.500000 ;
      RECT 2020.245000  3.640000 2020.535000  3.685000 ;
      RECT 2020.715000  2.110000 2021.005000  2.155000 ;
      RECT 2020.715000  2.295000 2021.005000  2.340000 ;
      RECT 2020.715000  3.100000 2021.005000  3.145000 ;
      RECT 2020.715000  3.285000 2021.005000  3.330000 ;
      RECT 2021.185000  1.755000 2021.475000  1.800000 ;
      RECT 2021.185000  1.940000 2021.475000  1.985000 ;
      RECT 2021.185000  3.455000 2021.475000  3.500000 ;
      RECT 2021.185000  3.640000 2021.475000  3.685000 ;
      RECT 2021.665000  2.110000 2021.955000  2.155000 ;
      RECT 2021.665000  2.295000 2021.955000  2.340000 ;
      RECT 2021.665000  3.100000 2021.955000  3.145000 ;
      RECT 2021.665000  3.285000 2021.955000  3.330000 ;
      RECT 2022.645000  2.110000 2022.935000  2.155000 ;
      RECT 2022.645000  2.295000 2022.935000  2.340000 ;
      RECT 2022.645000  3.100000 2022.935000  3.145000 ;
      RECT 2022.645000  3.285000 2022.935000  3.330000 ;
      RECT 2023.585000  2.110000 2023.875000  2.155000 ;
      RECT 2023.585000  2.295000 2023.875000  2.340000 ;
      RECT 2023.585000  3.100000 2023.875000  3.145000 ;
      RECT 2023.585000  3.285000 2023.875000  3.330000 ;
      RECT 2025.045000  2.110000 2025.335000  2.155000 ;
      RECT 2025.045000  2.155000 2029.155000  2.295000 ;
      RECT 2025.045000  2.295000 2025.335000  2.340000 ;
      RECT 2025.045000  3.100000 2025.335000  3.145000 ;
      RECT 2025.045000  3.145000 2029.155000  3.285000 ;
      RECT 2025.045000  3.285000 2025.335000  3.330000 ;
      RECT 2025.985000  2.110000 2026.275000  2.155000 ;
      RECT 2025.985000  2.295000 2026.275000  2.340000 ;
      RECT 2025.985000  3.100000 2026.275000  3.145000 ;
      RECT 2025.985000  3.285000 2026.275000  3.330000 ;
      RECT 2026.965000  2.110000 2027.255000  2.155000 ;
      RECT 2026.965000  2.295000 2027.255000  2.340000 ;
      RECT 2026.965000  3.100000 2027.255000  3.145000 ;
      RECT 2026.965000  3.285000 2027.255000  3.330000 ;
      RECT 2027.445000  1.755000 2027.735000  1.800000 ;
      RECT 2027.445000  1.940000 2027.735000  1.985000 ;
      RECT 2027.445000  3.455000 2027.735000  3.500000 ;
      RECT 2027.445000  3.640000 2027.735000  3.685000 ;
      RECT 2027.915000  2.110000 2028.205000  2.155000 ;
      RECT 2027.915000  2.295000 2028.205000  2.340000 ;
      RECT 2027.915000  3.100000 2028.205000  3.145000 ;
      RECT 2027.915000  3.285000 2028.205000  3.330000 ;
      RECT 2028.385000  1.755000 2028.675000  1.800000 ;
      RECT 2028.385000  1.940000 2028.675000  1.985000 ;
      RECT 2028.385000  3.455000 2028.675000  3.500000 ;
      RECT 2028.385000  3.640000 2028.675000  3.685000 ;
      RECT 2028.865000  2.110000 2029.155000  2.155000 ;
      RECT 2028.865000  2.295000 2029.155000  2.340000 ;
      RECT 2028.865000  3.100000 2029.155000  3.145000 ;
      RECT 2028.865000  3.285000 2029.155000  3.330000 ;
      RECT 2032.645000  2.110000 2032.935000  2.155000 ;
      RECT 2032.645000  2.155000 2036.755000  2.295000 ;
      RECT 2032.645000  2.295000 2032.935000  2.340000 ;
      RECT 2032.645000  3.100000 2032.935000  3.145000 ;
      RECT 2032.645000  3.145000 2036.755000  3.285000 ;
      RECT 2032.645000  3.285000 2032.935000  3.330000 ;
      RECT 2033.125000  1.755000 2033.415000  1.800000 ;
      RECT 2033.125000  1.940000 2033.415000  1.985000 ;
      RECT 2033.125000  3.455000 2033.415000  3.500000 ;
      RECT 2033.125000  3.640000 2033.415000  3.685000 ;
      RECT 2033.595000  2.110000 2033.885000  2.155000 ;
      RECT 2033.595000  2.295000 2033.885000  2.340000 ;
      RECT 2033.595000  3.100000 2033.885000  3.145000 ;
      RECT 2033.595000  3.285000 2033.885000  3.330000 ;
      RECT 2034.065000  1.755000 2034.355000  1.800000 ;
      RECT 2034.065000  1.940000 2034.355000  1.985000 ;
      RECT 2034.065000  3.455000 2034.355000  3.500000 ;
      RECT 2034.065000  3.640000 2034.355000  3.685000 ;
      RECT 2034.545000  2.110000 2034.835000  2.155000 ;
      RECT 2034.545000  2.295000 2034.835000  2.340000 ;
      RECT 2034.545000  3.100000 2034.835000  3.145000 ;
      RECT 2034.545000  3.285000 2034.835000  3.330000 ;
      RECT 2035.525000  2.110000 2035.815000  2.155000 ;
      RECT 2035.525000  2.295000 2035.815000  2.340000 ;
      RECT 2035.525000  3.100000 2035.815000  3.145000 ;
      RECT 2035.525000  3.285000 2035.815000  3.330000 ;
      RECT 2036.465000  2.110000 2036.755000  2.155000 ;
      RECT 2036.465000  2.295000 2036.755000  2.340000 ;
      RECT 2036.465000  3.100000 2036.755000  3.145000 ;
      RECT 2036.465000  3.285000 2036.755000  3.330000 ;
      RECT 2038.385000  2.110000 2038.675000  2.155000 ;
      RECT 2038.385000  2.155000 2042.495000  2.295000 ;
      RECT 2038.385000  2.295000 2038.675000  2.340000 ;
      RECT 2038.385000  3.100000 2038.675000  3.145000 ;
      RECT 2038.385000  3.145000 2042.495000  3.285000 ;
      RECT 2038.385000  3.285000 2038.675000  3.330000 ;
      RECT 2039.325000  2.110000 2039.615000  2.155000 ;
      RECT 2039.325000  2.295000 2039.615000  2.340000 ;
      RECT 2039.325000  3.100000 2039.615000  3.145000 ;
      RECT 2039.325000  3.285000 2039.615000  3.330000 ;
      RECT 2040.305000  2.110000 2040.595000  2.155000 ;
      RECT 2040.305000  2.295000 2040.595000  2.340000 ;
      RECT 2040.305000  3.100000 2040.595000  3.145000 ;
      RECT 2040.305000  3.285000 2040.595000  3.330000 ;
      RECT 2040.785000  1.755000 2041.075000  1.800000 ;
      RECT 2040.785000  1.940000 2041.075000  1.985000 ;
      RECT 2040.785000  3.455000 2041.075000  3.500000 ;
      RECT 2040.785000  3.640000 2041.075000  3.685000 ;
      RECT 2041.255000  2.110000 2041.545000  2.155000 ;
      RECT 2041.255000  2.295000 2041.545000  2.340000 ;
      RECT 2041.255000  3.100000 2041.545000  3.145000 ;
      RECT 2041.255000  3.285000 2041.545000  3.330000 ;
      RECT 2041.725000  1.755000 2042.015000  1.800000 ;
      RECT 2041.725000  1.940000 2042.015000  1.985000 ;
      RECT 2041.725000  3.455000 2042.015000  3.500000 ;
      RECT 2041.725000  3.640000 2042.015000  3.685000 ;
      RECT 2042.205000  2.110000 2042.495000  2.155000 ;
      RECT 2042.205000  2.295000 2042.495000  2.340000 ;
      RECT 2042.205000  3.100000 2042.495000  3.145000 ;
      RECT 2042.205000  3.285000 2042.495000  3.330000 ;
      RECT 2045.985000  2.110000 2046.275000  2.155000 ;
      RECT 2045.985000  2.155000 2050.095000  2.295000 ;
      RECT 2045.985000  2.295000 2046.275000  2.340000 ;
      RECT 2045.985000  3.100000 2046.275000  3.145000 ;
      RECT 2045.985000  3.145000 2050.095000  3.285000 ;
      RECT 2045.985000  3.285000 2046.275000  3.330000 ;
      RECT 2046.465000  1.755000 2046.755000  1.800000 ;
      RECT 2046.465000  1.940000 2046.755000  1.985000 ;
      RECT 2046.465000  3.455000 2046.755000  3.500000 ;
      RECT 2046.465000  3.640000 2046.755000  3.685000 ;
      RECT 2046.935000  2.110000 2047.225000  2.155000 ;
      RECT 2046.935000  2.295000 2047.225000  2.340000 ;
      RECT 2046.935000  3.100000 2047.225000  3.145000 ;
      RECT 2046.935000  3.285000 2047.225000  3.330000 ;
      RECT 2047.405000  1.755000 2047.695000  1.800000 ;
      RECT 2047.405000  1.940000 2047.695000  1.985000 ;
      RECT 2047.405000  3.455000 2047.695000  3.500000 ;
      RECT 2047.405000  3.640000 2047.695000  3.685000 ;
      RECT 2047.885000  2.110000 2048.175000  2.155000 ;
      RECT 2047.885000  2.295000 2048.175000  2.340000 ;
      RECT 2047.885000  3.100000 2048.175000  3.145000 ;
      RECT 2047.885000  3.285000 2048.175000  3.330000 ;
      RECT 2048.865000  2.110000 2049.155000  2.155000 ;
      RECT 2048.865000  2.295000 2049.155000  2.340000 ;
      RECT 2048.865000  3.100000 2049.155000  3.145000 ;
      RECT 2048.865000  3.285000 2049.155000  3.330000 ;
      RECT 2049.805000  2.110000 2050.095000  2.155000 ;
      RECT 2049.805000  2.295000 2050.095000  2.340000 ;
      RECT 2049.805000  3.100000 2050.095000  3.145000 ;
      RECT 2049.805000  3.285000 2050.095000  3.330000 ;
      RECT 2051.265000  2.110000 2051.555000  2.155000 ;
      RECT 2051.265000  2.155000 2055.375000  2.295000 ;
      RECT 2051.265000  2.295000 2051.555000  2.340000 ;
      RECT 2051.265000  3.100000 2051.555000  3.145000 ;
      RECT 2051.265000  3.145000 2055.375000  3.285000 ;
      RECT 2051.265000  3.285000 2051.555000  3.330000 ;
      RECT 2052.205000  2.110000 2052.495000  2.155000 ;
      RECT 2052.205000  2.295000 2052.495000  2.340000 ;
      RECT 2052.205000  3.100000 2052.495000  3.145000 ;
      RECT 2052.205000  3.285000 2052.495000  3.330000 ;
      RECT 2053.185000  2.110000 2053.475000  2.155000 ;
      RECT 2053.185000  2.295000 2053.475000  2.340000 ;
      RECT 2053.185000  3.100000 2053.475000  3.145000 ;
      RECT 2053.185000  3.285000 2053.475000  3.330000 ;
      RECT 2053.665000  1.755000 2053.955000  1.800000 ;
      RECT 2053.665000  1.940000 2053.955000  1.985000 ;
      RECT 2053.665000  3.455000 2053.955000  3.500000 ;
      RECT 2053.665000  3.640000 2053.955000  3.685000 ;
      RECT 2054.135000  2.110000 2054.425000  2.155000 ;
      RECT 2054.135000  2.295000 2054.425000  2.340000 ;
      RECT 2054.135000  3.100000 2054.425000  3.145000 ;
      RECT 2054.135000  3.285000 2054.425000  3.330000 ;
      RECT 2054.605000  1.755000 2054.895000  1.800000 ;
      RECT 2054.605000  1.940000 2054.895000  1.985000 ;
      RECT 2054.605000  3.455000 2054.895000  3.500000 ;
      RECT 2054.605000  3.640000 2054.895000  3.685000 ;
      RECT 2055.085000  2.110000 2055.375000  2.155000 ;
      RECT 2055.085000  2.295000 2055.375000  2.340000 ;
      RECT 2055.085000  3.100000 2055.375000  3.145000 ;
      RECT 2055.085000  3.285000 2055.375000  3.330000 ;
      RECT 2058.865000  2.110000 2059.155000  2.155000 ;
      RECT 2058.865000  2.155000 2062.975000  2.295000 ;
      RECT 2058.865000  2.295000 2059.155000  2.340000 ;
      RECT 2058.865000  3.100000 2059.155000  3.145000 ;
      RECT 2058.865000  3.145000 2062.975000  3.285000 ;
      RECT 2058.865000  3.285000 2059.155000  3.330000 ;
      RECT 2059.345000  1.755000 2059.635000  1.800000 ;
      RECT 2059.345000  1.940000 2059.635000  1.985000 ;
      RECT 2059.345000  3.455000 2059.635000  3.500000 ;
      RECT 2059.345000  3.640000 2059.635000  3.685000 ;
      RECT 2059.815000  2.110000 2060.105000  2.155000 ;
      RECT 2059.815000  2.295000 2060.105000  2.340000 ;
      RECT 2059.815000  3.100000 2060.105000  3.145000 ;
      RECT 2059.815000  3.285000 2060.105000  3.330000 ;
      RECT 2060.285000  1.755000 2060.575000  1.800000 ;
      RECT 2060.285000  1.940000 2060.575000  1.985000 ;
      RECT 2060.285000  3.455000 2060.575000  3.500000 ;
      RECT 2060.285000  3.640000 2060.575000  3.685000 ;
      RECT 2060.765000  2.110000 2061.055000  2.155000 ;
      RECT 2060.765000  2.295000 2061.055000  2.340000 ;
      RECT 2060.765000  3.100000 2061.055000  3.145000 ;
      RECT 2060.765000  3.285000 2061.055000  3.330000 ;
      RECT 2061.745000  2.110000 2062.035000  2.155000 ;
      RECT 2061.745000  2.295000 2062.035000  2.340000 ;
      RECT 2061.745000  3.100000 2062.035000  3.145000 ;
      RECT 2061.745000  3.285000 2062.035000  3.330000 ;
      RECT 2062.685000  2.110000 2062.975000  2.155000 ;
      RECT 2062.685000  2.295000 2062.975000  2.340000 ;
      RECT 2062.685000  3.100000 2062.975000  3.145000 ;
      RECT 2062.685000  3.285000 2062.975000  3.330000 ;
      RECT 2064.260000  0.070000 2064.400000  5.370000 ;
    LAYER met2 ;
      RECT 156.165000 4.065000 156.845000 4.435000 ;
      RECT 175.310000 4.110000 176.080000 4.390000 ;
      RECT 178.555000 2.580000 179.325000 2.860000 ;
      RECT 178.555000 5.300000 179.325000 5.580000 ;
    LAYER met3 ;
      RECT 156.115000 4.085000 156.895000 4.415000 ;
      RECT 172.705000 4.090000 173.485000 4.410000 ;
      RECT 175.305000 4.085000 176.085000 4.415000 ;
      RECT 178.550000 2.555000 179.330000 2.885000 ;
      RECT 178.550000 5.275000 179.330000 5.605000 ;
    LAYER met4 ;
      RECT 154.090000 3.580000 156.870000 4.760000 ;
      RECT 172.280000 3.490000 173.460000 4.670000 ;
      RECT 174.880000 3.490000 176.060000 4.670000 ;
      RECT 178.350000 1.825000 179.530000 3.005000 ;
      RECT 178.350000 5.155000 179.530000 6.335000 ;
    LAYER met5 ;
      RECT 153.970000 3.280000 156.990000 3.490000 ;
      RECT 153.970000 3.495000 156.990000 4.880000 ;
      RECT 172.160000 3.280000 174.480000 4.880000 ;
      RECT 174.580000 1.615000 176.180000 6.545000 ;
      RECT 177.780000 2.365000 177.880000 2.465000 ;
      RECT 177.780000 5.695000 177.880000 5.795000 ;
    LAYER via ;
      RECT 156.215000 4.120000 156.475000 4.380000 ;
      RECT 156.535000 4.120000 156.795000 4.380000 ;
      RECT 175.470000 4.120000 175.730000 4.380000 ;
      RECT 175.790000 4.120000 176.050000 4.380000 ;
      RECT 178.650000 2.590000 178.910000 2.850000 ;
      RECT 178.650000 5.310000 178.910000 5.570000 ;
      RECT 178.970000 2.590000 179.230000 2.850000 ;
      RECT 178.970000 5.310000 179.230000 5.570000 ;
    LAYER via2 ;
      RECT 156.165000 4.110000 156.445000 4.390000 ;
      RECT 156.565000 4.110000 156.845000 4.390000 ;
      RECT 175.355000 4.110000 175.635000 4.390000 ;
      RECT 175.755000 4.110000 176.035000 4.390000 ;
      RECT 178.600000 2.580000 178.880000 2.860000 ;
      RECT 178.600000 5.300000 178.880000 5.580000 ;
      RECT 179.000000 2.580000 179.280000 2.860000 ;
      RECT 179.000000 5.300000 179.280000 5.580000 ;
    LAYER via3 ;
      RECT 156.145000 4.090000 156.465000 4.410000 ;
      RECT 156.545000 4.090000 156.865000 4.410000 ;
      RECT 172.735000 4.090000 173.055000 4.410000 ;
      RECT 173.135000 4.090000 173.455000 4.410000 ;
      RECT 175.335000 4.090000 175.655000 4.410000 ;
      RECT 175.735000 4.090000 176.055000 4.410000 ;
      RECT 178.580000 2.560000 178.900000 2.880000 ;
      RECT 178.580000 5.280000 178.900000 5.600000 ;
      RECT 178.980000 2.560000 179.300000 2.880000 ;
      RECT 178.980000 5.280000 179.300000 5.600000 ;
    LAYER via4 ;
      RECT 155.690000 3.580000 156.870000 4.760000 ;
  END
END sky130_fd_sc_hdll__tap
END LIBRARY
