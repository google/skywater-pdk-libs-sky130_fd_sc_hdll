* File: sky130_fd_sc_hdll__dlxtn_1.pex.spice
* Created: Wed Sep  2 08:29:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__DLXTN_1%GATE_N 4 5 7 8 10 13 19 20 24 26
c41 19 0 2.67999e-20 $X=0.23 $Y=1.19
c42 13 0 2.71124e-20 $X=0.52 $Y=0.805
r43 24 27 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r44 24 26 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r45 19 20 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r46 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r47 11 13 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.52 $Y2=0.805
r48 8 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.805
r49 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.445
r50 5 15 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.495 $Y=1.665
+ $X2=0.305 $Y2=1.665
r51 5 7 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.74
+ $X2=0.495 $Y2=2.135
r52 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r53 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r54 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r55 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_1%A_27_47# 1 2 8 9 11 14 18 19 21 24 28 29
+ 30 38 42 45 47 52 54 56 57 60 63 64 69 72 77
c163 8 0 2.67999e-20 $X=0.965 $Y=1.64
r164 68 69 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.235
+ $X2=0.99 $Y2=1.235
r165 64 77 6.77715 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=3.34 $Y=1.53
+ $X2=3.34 $Y2=1.415
r166 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.26 $Y=1.53
+ $X2=3.26 $Y2=1.53
r167 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.745 $Y=1.53
+ $X2=0.745 $Y2=1.53
r168 57 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.89 $Y=1.53
+ $X2=0.745 $Y2=1.53
r169 56 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.115 $Y=1.53
+ $X2=3.26 $Y2=1.53
r170 56 57 2.75371 $w=1.4e-07 $l=2.225e-06 $layer=MET1_cond $X=3.115 $Y=1.53
+ $X2=0.89 $Y2=1.53
r171 52 72 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.97 $Y=0.87
+ $X2=2.97 $Y2=0.705
r172 51 54 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.97 $Y=0.87
+ $X2=3.255 $Y2=0.87
r173 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.97
+ $Y=0.87 $X2=2.97 $Y2=0.87
r174 49 60 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.745 $Y=1.795
+ $X2=0.745 $Y2=1.53
r175 48 60 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.745 $Y=1.4
+ $X2=0.745 $Y2=1.53
r176 46 68 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=0.805 $Y=1.235
+ $X2=0.965 $Y2=1.235
r177 45 48 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.775 $Y=1.235
+ $X2=0.775 $Y2=1.4
r178 45 47 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.775 $Y=1.235
+ $X2=0.775 $Y2=1.07
r179 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.805
+ $Y=1.235 $X2=0.805 $Y2=1.235
r180 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.425
+ $Y=1.74 $X2=3.425 $Y2=1.74
r181 36 64 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=3.34 $Y=1.585
+ $X2=3.34 $Y2=1.53
r182 36 38 5.25378 $w=3.38e-07 $l=1.55e-07 $layer=LI1_cond $X=3.34 $Y=1.585
+ $X2=3.34 $Y2=1.74
r183 34 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=1.035
+ $X2=3.255 $Y2=0.87
r184 34 77 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.255 $Y=1.035
+ $X2=3.255 $Y2=1.415
r185 32 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.745 $Y=0.805
+ $X2=0.745 $Y2=1.07
r186 31 42 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r187 30 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.66 $Y=1.88
+ $X2=0.745 $Y2=1.795
r188 30 31 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.66 $Y=1.88
+ $X2=0.345 $Y2=1.88
r189 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.66 $Y=0.72
+ $X2=0.745 $Y2=0.805
r190 28 29 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.66 $Y=0.72
+ $X2=0.345 $Y2=0.72
r191 22 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r192 22 24 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r193 19 39 48.3784 $w=2.91e-07 $l=2.80624e-07 $layer=POLY_cond $X=3.49 $Y=1.99
+ $X2=3.425 $Y2=1.74
r194 19 21 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.49 $Y=1.99
+ $X2=3.49 $Y2=2.275
r195 18 72 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.96 $Y=0.415
+ $X2=2.96 $Y2=0.705
r196 12 69 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=1.235
r197 12 14 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=0.445
r198 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.965 $Y=1.74
+ $X2=0.965 $Y2=2.135
r199 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.64 $X2=0.965
+ $Y2=1.74
r200 7 68 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=0.965 $Y=1.37
+ $X2=0.965 $Y2=1.235
r201 7 8 89.5258 $w=2e-07 $l=2.7e-07 $layer=POLY_cond $X=0.965 $Y=1.37 $X2=0.965
+ $Y2=1.64
r202 2 42 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r203 1 24 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_1%D 2 3 5 8 10 14 17
c43 14 0 1.08116e-19 $X=1.725 $Y=1.04
r44 16 17 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.955 $Y=1.04
+ $X2=1.98 $Y2=1.04
r45 13 16 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=1.725 $Y=1.04
+ $X2=1.955 $Y2=1.04
r46 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.725
+ $Y=1.04 $X2=1.725 $Y2=1.04
r47 10 14 4.06745 $w=4.23e-07 $l=1.5e-07 $layer=LI1_cond $X=1.677 $Y=1.19
+ $X2=1.677 $Y2=1.04
r48 6 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.98 $Y=0.875
+ $X2=1.98 $Y2=1.04
r49 6 8 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.98 $Y=0.875 $X2=1.98
+ $Y2=0.445
r50 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.955 $Y=1.77
+ $X2=1.955 $Y2=2.165
r51 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.955 $Y=1.67 $X2=1.955
+ $Y2=1.77
r52 1 16 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.955 $Y=1.205
+ $X2=1.955 $Y2=1.04
r53 1 2 154.183 $w=2e-07 $l=4.65e-07 $layer=POLY_cond $X=1.955 $Y=1.205
+ $X2=1.955 $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_1%A_319_47# 1 2 8 9 11 14 17 19 21 22 23 24
+ 26 33 35
c88 33 0 2.1121e-19 $X=2.405 $Y=0.93
c89 19 0 7.13094e-20 $X=2.12 $Y=0.7
r90 33 36 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=0.93
+ $X2=2.405 $Y2=1.095
r91 33 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=0.93
+ $X2=2.405 $Y2=0.765
r92 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.405
+ $Y=0.93 $X2=2.405 $Y2=0.93
r93 26 28 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.72 $Y=0.51
+ $X2=1.72 $Y2=0.7
r94 23 32 8.96999 $w=3.41e-07 $l=2.18746e-07 $layer=LI1_cond $X=2.205 $Y=1.095
+ $X2=2.33 $Y2=0.93
r95 23 24 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.205 $Y=1.095
+ $X2=2.205 $Y2=1.495
r96 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.12 $Y=1.58
+ $X2=2.205 $Y2=1.495
r97 21 22 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.12 $Y=1.58
+ $X2=1.885 $Y2=1.58
r98 20 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.805 $Y=0.7
+ $X2=1.72 $Y2=0.7
r99 19 32 8.22874 $w=3.41e-07 $l=3.18119e-07 $layer=LI1_cond $X=2.12 $Y=0.7
+ $X2=2.33 $Y2=0.93
r100 19 20 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.12 $Y=0.7
+ $X2=1.805 $Y2=0.7
r101 15 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.72 $Y=1.665
+ $X2=1.885 $Y2=1.58
r102 15 17 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.72 $Y=1.665
+ $X2=1.72 $Y2=1.99
r103 14 35 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.42 $Y=0.445
+ $X2=2.42 $Y2=0.765
r104 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.425 $Y=1.77
+ $X2=2.425 $Y2=2.165
r105 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.425 $Y=1.67 $X2=2.425
+ $Y2=1.77
r106 8 36 190.657 $w=2e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=1.67
+ $X2=2.425 $Y2=1.095
r107 2 17 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.595
+ $Y=1.845 $X2=1.72 $Y2=1.99
r108 1 26 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.72 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_1%A_211_363# 1 2 7 8 9 11 12 16 20 22 24 25
+ 28 31 37
c110 8 0 1.86795e-19 $X=2.95 $Y=1.89
r111 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.87
+ $Y=1.52 $X2=2.87 $Y2=1.52
r112 34 36 33.8246 $w=2.85e-07 $l=2e-07 $layer=POLY_cond $X=2.892 $Y=1.32
+ $X2=2.892 $Y2=1.52
r113 32 37 14.1528 $w=2.83e-07 $l=3.5e-07 $layer=LI1_cond $X=2.812 $Y=1.87
+ $X2=2.812 $Y2=1.52
r114 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.755 $Y=1.87
+ $X2=2.755 $Y2=1.87
r115 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.255 $Y=1.87
+ $X2=1.255 $Y2=1.87
r116 25 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.4 $Y=1.87
+ $X2=1.255 $Y2=1.87
r117 24 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.61 $Y=1.87
+ $X2=2.755 $Y2=1.87
r118 24 25 1.49752 $w=1.4e-07 $l=1.21e-06 $layer=MET1_cond $X=2.61 $Y=1.87
+ $X2=1.4 $Y2=1.87
r119 22 28 3.73904 $w=2.23e-07 $l=7.3e-08 $layer=LI1_cond $X=1.227 $Y=1.797
+ $X2=1.227 $Y2=1.87
r120 22 23 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.227 $Y=1.797
+ $X2=1.227 $Y2=1.685
r121 20 23 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.2 $Y=0.51
+ $X2=1.2 $Y2=1.685
r122 14 16 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.4 $Y=1.245
+ $X2=3.4 $Y2=0.415
r123 13 34 17.7656 $w=1.5e-07 $l=1.58e-07 $layer=POLY_cond $X=3.05 $Y=1.32
+ $X2=2.892 $Y2=1.32
r124 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.325 $Y=1.32
+ $X2=3.4 $Y2=1.245
r125 12 13 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=3.325 $Y=1.32
+ $X2=3.05 $Y2=1.32
r126 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.95 $Y=1.99
+ $X2=2.95 $Y2=2.275
r127 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.95 $Y=1.89 $X2=2.95
+ $Y2=1.99
r128 7 36 32.2493 $w=2.85e-07 $l=1.9182e-07 $layer=POLY_cond $X=2.95 $Y=1.685
+ $X2=2.892 $Y2=1.52
r129 7 8 67.9733 $w=2e-07 $l=2.05e-07 $layer=POLY_cond $X=2.95 $Y=1.685 $X2=2.95
+ $Y2=1.89
r130 2 28 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.815 $X2=1.2 $Y2=1.96
r131 1 20 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_1%A_760_21# 1 2 9 11 13 14 16 17 19 20 27 31
+ 34 36 39 42 44 45
r70 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.335
+ $Y=1.16 $X2=5.335 $Y2=1.16
r71 37 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.79 $Y=1.16
+ $X2=4.705 $Y2=1.16
r72 37 39 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=4.79 $Y=1.16
+ $X2=5.335 $Y2=1.16
r73 36 44 7.80489 $w=1.95e-07 $l=1.77059e-07 $layer=LI1_cond $X=4.705 $Y=1.535
+ $X2=4.68 $Y2=1.7
r74 35 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=1.325
+ $X2=4.705 $Y2=1.16
r75 35 36 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.705 $Y=1.325
+ $X2=4.705 $Y2=1.535
r76 34 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=0.995
+ $X2=4.705 $Y2=1.16
r77 34 42 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.705 $Y=0.995
+ $X2=4.705 $Y2=0.825
r78 29 44 7.80489 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=4.68 $Y=1.865
+ $X2=4.68 $Y2=1.7
r79 29 31 21.2154 $w=2.18e-07 $l=4.05e-07 $layer=LI1_cond $X=4.68 $Y=1.865
+ $X2=4.68 $Y2=2.27
r80 25 42 6.3875 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=4.68 $Y=0.715
+ $X2=4.68 $Y2=0.825
r81 25 27 7.07181 $w=2.18e-07 $l=1.35e-07 $layer=LI1_cond $X=4.68 $Y=0.715
+ $X2=4.68 $Y2=0.58
r82 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.155
+ $Y=1.7 $X2=4.155 $Y2=1.7
r83 20 44 0.463323 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.57 $Y=1.7 $X2=4.68
+ $Y2=1.7
r84 20 22 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=4.57 $Y=1.7
+ $X2=4.155 $Y2=1.7
r85 17 40 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=5.395 $Y=0.995
+ $X2=5.335 $Y2=1.16
r86 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.395 $Y=0.995
+ $X2=5.395 $Y2=0.56
r87 14 40 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=5.37 $Y=1.41
+ $X2=5.335 $Y2=1.16
r88 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.37 $Y=1.41
+ $X2=5.37 $Y2=1.985
r89 11 23 49.5109 $w=4.1e-07 $l=3.55176e-07 $layer=POLY_cond $X=3.9 $Y=1.99
+ $X2=4.045 $Y2=1.7
r90 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.9 $Y=1.99 $X2=3.9
+ $Y2=2.275
r91 7 23 39.7867 $w=4.1e-07 $l=2.38642e-07 $layer=POLY_cond $X=3.875 $Y=1.535
+ $X2=4.045 $Y2=1.7
r92 7 9 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.875 $Y=1.535
+ $X2=3.875 $Y2=0.445
r93 2 44 600 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=1 $X=4.53
+ $Y=1.485 $X2=4.655 $Y2=1.755
r94 2 31 600 $w=1.7e-07 $l=8.45192e-07 $layer=licon1_PDIFF $count=1 $X=4.53
+ $Y=1.485 $X2=4.655 $Y2=2.27
r95 1 27 182 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_NDIFF $count=1 $X=4.53
+ $Y=0.235 $X2=4.655 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_1%A_607_47# 1 2 7 9 10 12 13 14 15 19 24 26
+ 29 32
c82 32 0 1.58879e-19 $X=3.765 $Y=1.16
r83 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.345
+ $Y=1.16 $X2=4.345 $Y2=1.16
r84 27 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=1.16
+ $X2=3.765 $Y2=1.16
r85 27 29 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.85 $Y=1.16
+ $X2=4.345 $Y2=1.16
r86 25 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.765 $Y=1.325
+ $X2=3.765 $Y2=1.16
r87 25 26 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.765 $Y=1.325
+ $X2=3.765 $Y2=2.255
r88 24 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.765 $Y=0.995
+ $X2=3.765 $Y2=1.16
r89 23 24 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.765 $Y=0.535
+ $X2=3.765 $Y2=0.995
r90 19 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.68 $Y=2.34
+ $X2=3.765 $Y2=2.255
r91 19 21 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.68 $Y=2.34
+ $X2=3.185 $Y2=2.34
r92 15 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.68 $Y=0.45
+ $X2=3.765 $Y2=0.535
r93 15 17 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.68 $Y=0.45
+ $X2=3.17 $Y2=0.45
r94 13 30 77.8133 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=4.79 $Y=1.16
+ $X2=4.345 $Y2=1.16
r95 13 14 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=4.79 $Y=1.16
+ $X2=4.89 $Y2=1.202
r96 10 14 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=4.915 $Y=0.995
+ $X2=4.89 $Y2=1.202
r97 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.915 $Y=0.995
+ $X2=4.915 $Y2=0.56
r98 7 14 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=4.89 $Y=1.41
+ $X2=4.89 $Y2=1.202
r99 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.89 $Y=1.41 $X2=4.89
+ $Y2=1.985
r100 2 21 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=2.065 $X2=3.185 $Y2=2.34
r101 1 17 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=3.035
+ $Y=0.235 $X2=3.17 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_1%VPWR 1 2 3 4 15 19 23 27 30 31 33 34 36 37
+ 38 40 62 63 66
c87 19 0 1.86795e-19 $X=2.19 $Y=2
r88 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r89 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r90 60 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r91 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r92 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r93 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r94 54 57 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r95 53 56 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r96 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r97 51 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r98 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r99 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r100 48 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r101 47 50 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r102 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r103 45 66 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r104 45 47 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r105 40 66 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r106 40 42 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r107 38 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r108 38 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r109 36 59 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.02 $Y=2.72
+ $X2=4.83 $Y2=2.72
r110 36 37 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.02 $Y=2.72
+ $X2=5.155 $Y2=2.72
r111 35 62 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r112 35 37 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=5.155 $Y2=2.72
r113 33 56 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.05 $Y=2.72
+ $X2=3.91 $Y2=2.72
r114 33 34 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.05 $Y=2.72 $X2=4.2
+ $Y2=2.72
r115 32 59 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.35 $Y=2.72
+ $X2=4.83 $Y2=2.72
r116 32 34 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.35 $Y=2.72 $X2=4.2
+ $Y2=2.72
r117 30 50 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.07 $Y2=2.72
r118 30 31 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.262 $Y2=2.72
r119 29 53 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.42 $Y=2.72
+ $X2=2.53 $Y2=2.72
r120 29 31 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.42 $Y=2.72
+ $X2=2.262 $Y2=2.72
r121 25 37 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=2.635
+ $X2=5.155 $Y2=2.72
r122 25 27 38.4148 $w=2.68e-07 $l=9e-07 $layer=LI1_cond $X=5.155 $Y=2.635
+ $X2=5.155 $Y2=1.735
r123 21 34 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.2 $Y=2.635 $X2=4.2
+ $Y2=2.72
r124 21 23 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=4.2 $Y=2.635
+ $X2=4.2 $Y2=2.3
r125 17 31 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.262 $Y=2.635
+ $X2=2.262 $Y2=2.72
r126 17 19 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=2.262 $Y=2.635
+ $X2=2.262 $Y2=2
r127 13 66 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r128 13 15 12.5859 $w=3.78e-07 $l=4.15e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.22
r129 4 27 300 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_PDIFF $count=2 $X=4.98
+ $Y=1.485 $X2=5.125 $Y2=1.735
r130 3 23 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=2.065 $X2=4.135 $Y2=2.3
r131 2 19 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=1.845 $X2=2.19 $Y2=2
r132 1 15 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.815 $X2=0.73 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_1%Q 1 2 7 8 9
r12 8 9 15.1637 $w=2.83e-07 $l=3.75e-07 $layer=LI1_cond $X=5.732 $Y=1.835
+ $X2=5.732 $Y2=2.21
r13 7 8 53.5785 $w=2.83e-07 $l=1.325e-06 $layer=LI1_cond $X=5.732 $Y=0.51
+ $X2=5.732 $Y2=1.835
r14 2 8 300 $w=1.7e-07 $l=4.44691e-07 $layer=licon1_PDIFF $count=2 $X=5.46
+ $Y=1.485 $X2=5.675 $Y2=1.835
r15 1 7 182 $w=1.7e-07 $l=4.35603e-07 $layer=licon1_NDIFF $count=1 $X=5.47
+ $Y=0.235 $X2=5.675 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_1%VGND 1 2 3 4 15 19 22 23 25 26 27 29 34 50
+ 51 55 62
c88 62 0 1.03094e-19 $X=2.07 $Y=0
c89 51 0 2.71124e-20 $X=5.75 $Y=0
c90 2 0 7.13094e-20 $X=2.055 $Y=0.235
r91 62 65 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=2.165 $Y=0 $X2=2.165
+ $Y2=0.36
r92 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r93 55 58 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0 $X2=0.705
+ $Y2=0.38
r94 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r95 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r96 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r97 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r98 45 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r99 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r100 42 45 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.91 $Y2=0
r101 42 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r102 41 44 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r103 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r104 39 62 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.165
+ $Y2=0
r105 39 41 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.355 $Y=0
+ $X2=2.53 $Y2=0
r106 38 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r107 38 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r108 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r109 35 55 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r110 35 37 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.61 $Y2=0
r111 34 62 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=2.165
+ $Y2=0
r112 34 37 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.975 $Y=0
+ $X2=1.61 $Y2=0
r113 29 55 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r114 29 31 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r115 27 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r116 27 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r117 25 47 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.02 $Y=0 $X2=4.83
+ $Y2=0
r118 25 26 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.02 $Y=0 $X2=5.155
+ $Y2=0
r119 24 50 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r120 24 26 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.29 $Y=0 $X2=5.155
+ $Y2=0
r121 22 44 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.02 $Y=0 $X2=3.91
+ $Y2=0
r122 22 23 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.02 $Y=0 $X2=4.16
+ $Y2=0
r123 21 47 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.3 $Y=0 $X2=4.83
+ $Y2=0
r124 21 23 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.3 $Y=0 $X2=4.16
+ $Y2=0
r125 17 26 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=0.085
+ $X2=5.155 $Y2=0
r126 17 19 19.8476 $w=2.68e-07 $l=4.65e-07 $layer=LI1_cond $X=5.155 $Y=0.085
+ $X2=5.155 $Y2=0.55
r127 13 23 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.16 $Y=0.085
+ $X2=4.16 $Y2=0
r128 13 15 14.8171 $w=2.78e-07 $l=3.6e-07 $layer=LI1_cond $X=4.16 $Y=0.085
+ $X2=4.16 $Y2=0.445
r129 4 19 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=4.99
+ $Y=0.235 $X2=5.125 $Y2=0.55
r130 3 15 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=3.95
+ $Y=0.235 $X2=4.135 $Y2=0.445
r131 2 65 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.055
+ $Y=0.235 $X2=2.19 $Y2=0.36
r132 1 58 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

