* File: sky130_fd_sc_hdll__sdfbbp_1.spice
* Created: Wed Sep  2 08:50:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__sdfbbp_1.pex.spice"
.subckt sky130_fd_sc_hdll__sdfbbp_1  VNB VPB CLK SCD SCE D SET_B RESET_B VPWR
+ Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* D	D
* SCE	SCE
* SCD	SCD
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1033 N_VGND_M1033_d N_CLK_M1033_g N_A_27_47#_M1033_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_A_211_363#_M1001_d N_A_27_47#_M1001_g N_VGND_M1033_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0672 PD=1.36 PS=0.74 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 A_411_47# N_SCD_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1302 PD=0.63 PS=1.46 NRD=14.28 NRS=12.852 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1024 N_A_483_47#_M1024_d N_SCE_M1024_g A_411_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1449 AS=0.0441 PD=1.53 PS=0.63 NRD=22.848 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_SCE_M1003_g N_A_453_315#_M1003_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0798 AS=0.1365 PD=0.8 PS=1.49 NRD=15.708 NRS=17.136 M=1 R=2.8
+ SA=75000.2 SB=75003.9 A=0.063 P=1.14 MULT=1
MM1045 A_824_47# N_A_453_315#_M1045_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0546 AS=0.0798 PD=0.68 PS=0.8 NRD=21.42 NRS=12.852 M=1 R=2.8 SA=75000.8
+ SB=75003.4 A=0.063 P=1.14 MULT=1
MM1035 N_A_483_47#_M1035_d N_D_M1035_g A_824_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0730154 AS=0.0546 PD=0.813077 PS=0.68 NRD=17.136 NRS=21.42 M=1 R=2.8
+ SA=75001.2 SB=75003 A=0.063 P=1.14 MULT=1
MM1027 N_A_1003_47#_M1027_d N_A_27_47#_M1027_g N_A_483_47#_M1035_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0792 AS=0.0625846 PD=0.8 PS=0.696923 NRD=36.66 NRS=0 M=1
+ R=2.4 SA=75001.7 SB=75003 A=0.054 P=1.02 MULT=1
MM1019 A_1121_47# N_A_211_363#_M1019_g N_A_1003_47#_M1027_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0702 AS=0.0792 PD=0.738462 PS=0.8 NRD=46.656 NRS=16.656 M=1 R=2.4
+ SA=75002.3 SB=75002.4 A=0.054 P=1.02 MULT=1
MM1025 N_VGND_M1025_d N_A_1197_21#_M1025_g A_1121_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1008 AS=0.0819 PD=0.9 PS=0.861538 NRD=55.704 NRS=39.996 M=1 R=2.8
+ SA=75002.4 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1009 N_A_1353_47#_M1009_d N_SET_B_M1009_g N_VGND_M1025_d VNB NSHORT L=0.15
+ W=0.42 AD=0.101553 AS=0.1008 PD=0.855849 PS=0.9 NRD=9.996 NRS=1.428 M=1 R=2.8
+ SA=75003.1 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1013 N_A_1197_21#_M1013_d N_A_1003_47#_M1013_g N_A_1353_47#_M1009_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.0864 AS=0.154747 PD=0.91 PS=1.30415 NRD=0 NRS=23.436 M=1
+ R=4.26667 SA=75002.5 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1021 N_A_1353_47#_M1021_d N_A_1525_21#_M1021_g N_A_1197_21#_M1013_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.0864 PD=1.85 PS=0.91 NRD=3.744 NRS=0 M=1
+ R=4.26667 SA=75002.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1037 A_1769_47# N_A_1197_21#_M1037_g N_VGND_M1037_s VNB NSHORT L=0.15 W=0.64
+ AD=0.11968 AS=0.2336 PD=1.2352 PS=2.01 NRD=24.744 NRS=18.744 M=1 R=4.26667
+ SA=75000.3 SB=75002 A=0.096 P=1.58 MULT=1
MM1010 N_A_1864_47#_M1010_d N_A_211_363#_M1010_g A_1769_47# VNB NSHORT L=0.15
+ W=0.36 AD=0.0882 AS=0.06732 PD=0.85 PS=0.6948 NRD=39.996 NRS=43.992 M=1 R=2.4
+ SA=75000.8 SB=75002.9 A=0.054 P=1.02 MULT=1
MM1046 A_1992_47# N_A_27_47#_M1046_g N_A_1864_47#_M1010_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0618923 AS=0.0882 PD=0.692308 PS=0.85 NRD=38.964 NRS=30 M=1 R=2.4
+ SA=75001.4 SB=75002.3 A=0.054 P=1.02 MULT=1
MM1014 N_VGND_M1014_d N_A_2058_21#_M1014_g A_1992_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1029 AS=0.0722077 PD=0.91 PS=0.807692 NRD=15.708 NRS=33.396 M=1 R=2.8
+ SA=75001.6 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1000 N_A_2216_47#_M1000_d N_SET_B_M1000_g N_VGND_M1014_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0898245 AS=0.1029 PD=0.808302 PS=0.91 NRD=0 NRS=44.28 M=1 R=2.8
+ SA=75002.3 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1040 N_A_2058_21#_M1040_d N_A_1864_47#_M1040_g N_A_2216_47#_M1000_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1008 AS=0.136875 PD=0.955 PS=1.2317 NRD=0 NRS=19.68 M=1
+ R=4.26667 SA=75001.9 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1007 N_A_2216_47#_M1007_d N_A_1525_21#_M1007_g N_A_2058_21#_M1040_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1664 AS=0.1008 PD=1.8 PS=0.955 NRD=0 NRS=6.552 M=1
+ R=4.26667 SA=75002.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1028 N_VGND_M1028_d N_RESET_B_M1028_g N_A_1525_21#_M1028_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0914579 AS=0.1302 PD=0.812523 PS=1.46 NRD=17.856 NRS=12.852 M=1
+ R=2.8 SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1005 N_Q_N_M1005_d N_A_2058_21#_M1005_g N_VGND_M1028_d VNB NSHORT L=0.15
+ W=0.65 AD=0.23075 AS=0.141542 PD=2.01 PS=1.25748 NRD=16.608 NRS=8.304 M=1
+ R=4.33333 SA=75000.6 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1043 N_VGND_M1043_d N_A_2058_21#_M1043_g N_A_2845_47#_M1043_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0889065 AS=0.1302 PD=0.804673 PS=1.46 NRD=14.28 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1047 N_Q_M1047_d N_A_2845_47#_M1047_g N_VGND_M1043_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.137593 PD=1.82 PS=1.24533 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_VPWR_M1008_d N_CLK_M1008_g N_A_27_47#_M1008_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1038 N_A_211_363#_M1038_d N_A_27_47#_M1038_g N_VPWR_M1008_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1018 A_409_363# N_SCD_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0736 AS=0.1728 PD=0.87 PS=1.82 NRD=18.4589 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1022 N_A_483_47#_M1022_d N_A_453_315#_M1022_g A_409_363# VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.0736 PD=1.82 PS=0.87 NRD=1.5366 NRS=18.4589 M=1
+ R=3.55556 SA=90000.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1011 N_VPWR_M1011_d N_SCE_M1011_g N_A_453_315#_M1011_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0609 AS=0.1449 PD=0.71 PS=1.53 NRD=2.3443 NRS=37.5088 M=1
+ R=2.33333 SA=90000.3 SB=90008.6 A=0.0756 P=1.2 MULT=1
MM1004 A_810_413# N_SCE_M1004_g N_VPWR_M1011_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0609 AS=0.0609 PD=0.71 PS=0.71 NRD=42.1974 NRS=2.3443 M=1 R=2.33333
+ SA=90000.7 SB=90008.1 A=0.0756 P=1.2 MULT=1
MM1044 N_A_483_47#_M1044_d N_D_M1044_g A_810_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.07455 AS=0.0609 PD=0.775 PS=0.71 NRD=32.8202 NRS=42.1974 M=1 R=2.33333
+ SA=90001.2 SB=90007.7 A=0.0756 P=1.2 MULT=1
MM1020 N_A_1003_47#_M1020_d N_A_211_363#_M1020_g N_A_483_47#_M1044_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.0609 AS=0.07455 PD=0.71 PS=0.775 NRD=2.3443 NRS=2.3443 M=1
+ R=2.33333 SA=90001.7 SB=90007.1 A=0.0756 P=1.2 MULT=1
MM1006 A_1105_413# N_A_27_47#_M1006_g N_A_1003_47#_M1020_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0987 AS=0.0609 PD=0.89 PS=0.71 NRD=84.4145 NRS=2.3443 M=1
+ R=2.33333 SA=90002.2 SB=90006.7 A=0.0756 P=1.2 MULT=1
MM1015 N_VPWR_M1015_d N_A_1197_21#_M1015_g A_1105_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.084 AS=0.0987 PD=0.82 PS=0.89 NRD=25.7873 NRS=84.4145 M=1 R=2.33333
+ SA=90002.8 SB=90006 A=0.0756 P=1.2 MULT=1
MM1012 N_A_1197_21#_M1012_d N_SET_B_M1012_g N_VPWR_M1015_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1022 AS=0.084 PD=0.833333 PS=0.82 NRD=58.6272 NRS=30.4759 M=1
+ R=2.33333 SA=90003.4 SB=90005.4 A=0.0756 P=1.2 MULT=1
MM1031 A_1469_329# N_A_1003_47#_M1031_g N_A_1197_21#_M1012_d VPB PHIGHVT L=0.18
+ W=0.84 AD=0.1218 AS=0.2044 PD=1.13 PS=1.66667 NRD=21.0987 NRS=1.1623 M=1
+ R=4.66667 SA=90002.1 SB=90003.1 A=0.1512 P=2.04 MULT=1
MM1026 N_VPWR_M1026_d N_A_1525_21#_M1026_g A_1469_329# VPB PHIGHVT L=0.18 W=0.84
+ AD=0.2331 AS=0.1218 PD=1.395 PS=1.13 NRD=8.1952 NRS=21.0987 M=1 R=4.66667
+ SA=90002.6 SB=90002.7 A=0.1512 P=2.04 MULT=1
MM1041 A_1710_329# N_A_1197_21#_M1041_g N_VPWR_M1026_d VPB PHIGHVT L=0.18 W=0.84
+ AD=0.2688 AS=0.2331 PD=1.97333 PS=1.395 NRD=62.1338 NRS=56.2829 M=1 R=4.66667
+ SA=90003.3 SB=90001.9 A=0.1512 P=2.04 MULT=1
MM1042 N_A_1864_47#_M1042_d N_A_27_47#_M1042_g A_1710_329# VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0609 AS=0.1344 PD=0.71 PS=0.986667 NRD=2.3443 NRS=124.287 M=1
+ R=2.33333 SA=90006 SB=90002.8 A=0.0756 P=1.2 MULT=1
MM1032 A_1968_413# N_A_211_363#_M1032_g N_A_1864_47#_M1042_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0966 AS=0.0609 PD=0.88 PS=0.71 NRD=82.0702 NRS=2.3443 M=1
+ R=2.33333 SA=90006.5 SB=90002.3 A=0.0756 P=1.2 MULT=1
MM1029 N_VPWR_M1029_d N_A_2058_21#_M1029_g A_1968_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0861 AS=0.0966 PD=0.83 PS=0.88 NRD=30.4759 NRS=82.0702 M=1 R=2.33333
+ SA=90007.2 SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1002 N_A_2058_21#_M1002_d N_SET_B_M1002_g N_VPWR_M1029_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0861 AS=0.0861 PD=0.793333 PS=0.83 NRD=30.4759 NRS=30.4759 M=1
+ R=2.33333 SA=90007.7 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1034 A_2320_329# N_A_1864_47#_M1034_g N_A_2058_21#_M1002_d VPB PHIGHVT L=0.18
+ W=0.84 AD=0.0966 AS=0.1722 PD=1.07 PS=1.58667 NRD=14.0658 NRS=1.1623 M=1
+ R=4.66667 SA=90004.2 SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1036 N_VPWR_M1036_d N_A_1525_21#_M1036_g A_2320_329# VPB PHIGHVT L=0.18 W=0.84
+ AD=0.2268 AS=0.0966 PD=2.22 PS=1.07 NRD=1.1623 NRS=14.0658 M=1 R=4.66667
+ SA=90004.6 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1017 N_VPWR_M1017_d N_RESET_B_M1017_g N_A_1525_21#_M1017_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.126517 AS=0.1728 PD=1.05756 PS=1.82 NRD=43.9113 NRS=1.5366 M=1
+ R=3.55556 SA=90000.2 SB=90000.8 A=0.1152 P=1.64 MULT=1
MM1039 N_Q_N_M1039_d N_A_2058_21#_M1039_g N_VPWR_M1017_d VPB PHIGHVT L=0.18 W=1
+ AD=0.365 AS=0.197683 PD=2.73 PS=1.65244 NRD=19.7 NRS=0.9653 M=1 R=5.55556
+ SA=90000.5 SB=90000.3 A=0.18 P=2.36 MULT=1
MM1030 N_VPWR_M1030_d N_A_2058_21#_M1030_g N_A_2845_47#_M1030_s VPB PHIGHVT
+ L=0.18 W=0.64 AD=0.122693 AS=0.1728 PD=1.04976 PS=1.82 NRD=18.4589 NRS=1.5366
+ M=1 R=3.55556 SA=90000.2 SB=90000.7 A=0.1152 P=1.64 MULT=1
MM1016 N_Q_M1016_d N_A_2845_47#_M1016_g N_VPWR_M1030_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.191707 PD=2.54 PS=1.64024 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.5 SB=90000.2 A=0.18 P=2.36 MULT=1
DX48_noxref VNB VPB NWDIODE A=25.7121 P=35.25
c_147 VNB 0 4.38175e-20 $X=0.145 $Y=-0.085
c_291 VPB 0 1.98844e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__sdfbbp_1.pxi.spice"
*
.ends
*
*
