* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 VPWR A1 a_425_297# VPB phighvt w=1e+06u l=180000u
+  ad=6.607e+11p pd=5.42e+06u as=2.8e+11p ps=2.56e+06u
M1001 a_425_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.2e+11p ps=2.64e+06u
M1002 a_105_352# B1_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=3.615e+11p ps=3.5e+06u
M1003 VGND A2 a_327_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.965e+11p ps=3.82e+06u
M1004 a_327_47# a_105_352# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1005 a_327_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR B1_N a_105_352# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1007 Y a_105_352# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
