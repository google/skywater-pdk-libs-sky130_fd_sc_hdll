* File: sky130_fd_sc_hdll__and4bb_1.pex.spice
* Created: Thu Aug 27 18:59:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND4BB_1%A_N 3 5 7 8 12
c31 3 0 1.51173e-19 $X=0.53 $Y=0.445
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.745 $X2=0.59 $Y2=1.745
r33 8 12 2.95498 $w=3.88e-07 $l=1e-07 $layer=LI1_cond $X=0.62 $Y=1.845 $X2=0.62
+ $Y2=1.745
r34 5 11 50.4353 $w=2.56e-07 $l=2.61916e-07 $layer=POLY_cond $X=0.555 $Y=1.99
+ $X2=0.59 $Y2=1.745
r35 5 7 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.555 $Y=1.99
+ $X2=0.555 $Y2=2.275
r36 1 11 39.2615 $w=2.56e-07 $l=1.92678e-07 $layer=POLY_cond $X=0.53 $Y=1.58
+ $X2=0.59 $Y2=1.745
r37 1 3 581.989 $w=1.5e-07 $l=1.135e-06 $layer=POLY_cond $X=0.53 $Y=1.58
+ $X2=0.53 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_1%B_N 2 3 5 8 12 13 15
c42 12 0 1.51173e-19 $X=1 $Y=1.03
c43 2 0 1.84374e-19 $X=1.035 $Y=1.89
r44 15 23 7.97845 $w=2.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.655 $Y=0.85
+ $X2=0.655 $Y2=1.03
r45 13 19 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.03 $X2=1
+ $Y2=1.195
r46 13 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.03 $X2=1
+ $Y2=0.865
r47 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.03
+ $X2=1 $Y2=1.03
r48 10 23 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.785 $Y=1.03
+ $X2=0.655 $Y2=1.03
r49 10 12 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.785 $Y=1.03 $X2=1
+ $Y2=1.03
r50 8 18 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.06 $Y=0.445
+ $X2=1.06 $Y2=0.865
r51 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.035 $Y=1.99
+ $X2=1.035 $Y2=2.275
r52 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.035 $Y=1.89 $X2=1.035
+ $Y2=1.99
r53 2 19 230.446 $w=2e-07 $l=6.95e-07 $layer=POLY_cond $X=1.035 $Y=1.89
+ $X2=1.035 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_1%A_27_47# 1 2 7 9 12 14 15 17 19 20 24 30
+ 32 36 38
c85 24 0 1.84374e-19 $X=1.48 $Y=1.66
r86 38 40 15.1913 $w=2.18e-07 $l=2.9e-07 $layer=LI1_cond $X=1.125 $Y=1.37
+ $X2=1.125 $Y2=1.66
r87 33 36 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.17 $Y=2.3 $X2=0.26
+ $Y2=2.3
r88 27 30 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.17 $Y=0.42 $X2=0.26
+ $Y2=0.42
r89 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.48
+ $Y=1.66 $X2=1.48 $Y2=1.66
r90 22 40 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.235 $Y=1.66
+ $X2=1.125 $Y2=1.66
r91 22 24 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.235 $Y=1.66
+ $X2=1.48 $Y2=1.66
r92 21 32 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.255 $Y=1.37
+ $X2=0.17 $Y2=1.37
r93 20 38 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.015 $Y=1.37
+ $X2=1.125 $Y2=1.37
r94 20 21 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=1.015 $Y=1.37
+ $X2=0.255 $Y2=1.37
r95 19 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=2.135
+ $X2=0.17 $Y2=2.3
r96 18 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.17 $Y=1.455
+ $X2=0.17 $Y2=1.37
r97 18 19 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.17 $Y=1.455
+ $X2=0.17 $Y2=2.135
r98 17 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.17 $Y=1.285
+ $X2=0.17 $Y2=1.37
r99 16 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.17 $Y2=0.42
r100 16 17 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.17 $Y2=1.285
r101 14 25 77.8133 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=1.925 $Y=1.66
+ $X2=1.48 $Y2=1.66
r102 14 15 3.90195 $w=3.3e-07 $l=1.34907e-07 $layer=POLY_cond $X=1.925 $Y=1.66
+ $X2=2.025 $Y2=1.742
r103 10 15 34.7346 $w=1.65e-07 $l=2.59199e-07 $layer=POLY_cond $X=2.05 $Y=1.495
+ $X2=2.025 $Y2=1.742
r104 10 12 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.05 $Y=1.495
+ $X2=2.05 $Y2=0.675
r105 7 15 34.7346 $w=1.65e-07 $l=2.48e-07 $layer=POLY_cond $X=2.025 $Y=1.99
+ $X2=2.025 $Y2=1.742
r106 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.025 $Y=1.99
+ $X2=2.025 $Y2=2.275
r107 2 36 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
r108 1 30 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_1%A_225_413# 1 2 9 11 12 14 17 19 20 22 23
+ 25 26 28 31 32 34 40
r101 37 38 13.5455 $w=3.98e-07 $l=3.35e-07 $layer=LI1_cond $X=1.385 $Y=0.42
+ $X2=1.385 $Y2=0.755
r102 34 37 2.30489 $w=3.98e-07 $l=8e-08 $layer=LI1_cond $X=1.385 $Y=0.34
+ $X2=1.385 $Y2=0.42
r103 32 41 37.9622 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.56 $Y=1.16
+ $X2=2.56 $Y2=1.325
r104 32 40 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.56 $Y=1.16
+ $X2=2.56 $Y2=0.995
r105 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.58
+ $Y=1.16 $X2=2.58 $Y2=1.16
r106 29 31 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.58 $Y=0.425
+ $X2=2.58 $Y2=1.16
r107 27 28 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.9 $Y=1.405
+ $X2=1.9 $Y2=1.915
r108 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.815 $Y=1.32
+ $X2=1.9 $Y2=1.405
r109 25 26 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.815 $Y=1.32
+ $X2=1.585 $Y2=1.32
r110 24 34 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=1.585 $Y=0.34
+ $X2=1.385 $Y2=0.34
r111 23 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.495 $Y=0.34
+ $X2=2.58 $Y2=0.425
r112 23 24 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=2.495 $Y=0.34
+ $X2=1.585 $Y2=0.34
r113 22 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.5 $Y=1.235
+ $X2=1.585 $Y2=1.32
r114 22 38 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.5 $Y=1.235
+ $X2=1.5 $Y2=0.755
r115 19 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.815 $Y=2
+ $X2=1.9 $Y2=1.915
r116 19 20 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=1.815 $Y=2
+ $X2=1.375 $Y2=2
r117 15 20 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.27 $Y=2.085
+ $X2=1.375 $Y2=2
r118 15 17 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.27 $Y=2.085
+ $X2=1.27 $Y2=2.3
r119 12 14 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.505 $Y=1.99
+ $X2=2.505 $Y2=2.275
r120 11 12 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.505 $Y=1.89 $X2=2.505
+ $Y2=1.99
r121 11 41 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=2.505 $Y=1.89
+ $X2=2.505 $Y2=1.325
r122 9 40 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.48 $Y=0.675
+ $X2=2.48 $Y2=0.995
r123 2 17 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=2.065 $X2=1.27 $Y2=2.3
r124 1 37 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.135
+ $Y=0.235 $X2=1.27 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_1%C 3 5 6 8 9 10 11 12 18 20
c43 9 0 1.48364e-19 $X=3 $Y=0.51
r44 18 21 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.06 $Y=1.16
+ $X2=3.06 $Y2=1.325
r45 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.06 $Y=1.16
+ $X2=3.06 $Y2=0.995
r46 11 12 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.025 $Y=1.16
+ $X2=3.025 $Y2=1.53
r47 11 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.06
+ $Y=1.16 $X2=3.06 $Y2=1.16
r48 10 11 11.9086 $w=2.98e-07 $l=3.1e-07 $layer=LI1_cond $X=3.025 $Y=0.85
+ $X2=3.025 $Y2=1.16
r49 9 10 13.061 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=3.025 $Y=0.51
+ $X2=3.025 $Y2=0.85
r50 6 8 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.025 $Y=1.99
+ $X2=3.025 $Y2=2.275
r51 5 6 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.025 $Y=1.89 $X2=3.025
+ $Y2=1.99
r52 5 21 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=3.025 $Y=1.89
+ $X2=3.025 $Y2=1.325
r53 3 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3 $Y=0.675 $X2=3
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_1%D 2 3 5 8 9 10 11 12 18 20
r44 18 21 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.54 $Y=1.16
+ $X2=3.54 $Y2=1.325
r45 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.54 $Y=1.16
+ $X2=3.54 $Y2=0.995
r46 11 12 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=3.492 $Y=1.16
+ $X2=3.492 $Y2=1.53
r47 11 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.54
+ $Y=1.16 $X2=3.54 $Y2=1.16
r48 10 11 12.1104 $w=2.93e-07 $l=3.1e-07 $layer=LI1_cond $X=3.492 $Y=0.85
+ $X2=3.492 $Y2=1.16
r49 9 10 13.2824 $w=2.93e-07 $l=3.4e-07 $layer=LI1_cond $X=3.492 $Y=0.51
+ $X2=3.492 $Y2=0.85
r50 8 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.6 $Y=0.675 $X2=3.6
+ $Y2=0.995
r51 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.575 $Y=1.99
+ $X2=3.575 $Y2=2.275
r52 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.575 $Y=1.89 $X2=3.575
+ $Y2=1.99
r53 2 21 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=3.575 $Y=1.89
+ $X2=3.575 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_1%A_339_93# 1 2 3 10 12 13 15 16 21 24 26
+ 30 32 35 36 37 41
r89 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.02
+ $Y=1.16 $X2=4.02 $Y2=1.16
r90 38 41 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.895 $Y=1.16
+ $X2=4.02 $Y2=1.16
r91 34 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.895 $Y=1.325
+ $X2=3.895 $Y2=1.16
r92 34 35 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.895 $Y=1.325
+ $X2=3.895 $Y2=1.915
r93 33 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.38 $Y=2 $X2=3.295
+ $Y2=2
r94 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.81 $Y=2
+ $X2=3.895 $Y2=1.915
r95 32 33 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.81 $Y=2 $X2=3.38
+ $Y2=2
r96 28 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.295 $Y=2.085
+ $X2=3.295 $Y2=2
r97 28 30 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.295 $Y=2.085
+ $X2=3.295 $Y2=2.3
r98 27 36 1.34256 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.355 $Y=2 $X2=2.255
+ $Y2=2
r99 26 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=2 $X2=3.295
+ $Y2=2
r100 26 27 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=3.21 $Y=2
+ $X2=2.355 $Y2=2
r101 22 36 5.16603 $w=1.7e-07 $l=9.21954e-08 $layer=LI1_cond $X=2.27 $Y=2.085
+ $X2=2.255 $Y2=2
r102 22 24 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.27 $Y=2.085
+ $X2=2.27 $Y2=2.3
r103 21 36 5.16603 $w=1.7e-07 $l=9.21954e-08 $layer=LI1_cond $X=2.24 $Y=1.915
+ $X2=2.255 $Y2=2
r104 20 21 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=2.24 $Y=0.925
+ $X2=2.24 $Y2=1.915
r105 16 20 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.155 $Y=0.76
+ $X2=2.24 $Y2=0.925
r106 16 18 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.155 $Y=0.76
+ $X2=1.84 $Y2=0.76
r107 13 42 38.6072 $w=2.91e-07 $l=2.02287e-07 $layer=POLY_cond $X=4.125 $Y=0.995
+ $X2=4.042 $Y2=1.16
r108 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.125 $Y=0.995
+ $X2=4.125 $Y2=0.56
r109 10 42 48.3784 $w=2.91e-07 $l=2.77489e-07 $layer=POLY_cond $X=4.1 $Y=1.41
+ $X2=4.042 $Y2=1.16
r110 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.1 $Y=1.41
+ $X2=4.1 $Y2=1.985
r111 3 30 600 $w=1.7e-07 $l=3.1229e-07 $layer=licon1_PDIFF $count=1 $X=3.115
+ $Y=2.065 $X2=3.295 $Y2=2.3
r112 2 24 600 $w=1.7e-07 $l=3.02738e-07 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=2.065 $X2=2.27 $Y2=2.3
r113 1 18 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=1.695
+ $Y=0.465 $X2=1.84 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_1%VPWR 1 2 3 4 15 19 22 23 25 28 31 33 45
+ 51 52 55 62
r79 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r80 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r81 55 58 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.765 $Y=2.34
+ $X2=0.765 $Y2=2.72
r82 52 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r83 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r84 49 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.03 $Y=2.72
+ $X2=3.865 $Y2=2.72
r85 49 51 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.03 $Y=2.72
+ $X2=4.37 $Y2=2.72
r86 48 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r87 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r88 45 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.7 $Y=2.72
+ $X2=3.865 $Y2=2.72
r89 45 47 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.7 $Y=2.72 $X2=3.45
+ $Y2=2.72
r90 44 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r91 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r92 41 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r93 41 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r94 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r95 38 58 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.955 $Y=2.72
+ $X2=0.765 $Y2=2.72
r96 38 40 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r97 33 58 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.765 $Y2=2.72
r98 33 35 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.23 $Y2=2.72
r99 31 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r100 31 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r101 29 47 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.93 $Y=2.72
+ $X2=3.45 $Y2=2.72
r102 28 43 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=2.55 $Y=2.72 $X2=2.53
+ $Y2=2.72
r103 27 29 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.74 $Y=2.72
+ $X2=2.93 $Y2=2.72
r104 27 28 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.74 $Y=2.72
+ $X2=2.55 $Y2=2.72
r105 25 27 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=2.74 $Y=2.34
+ $X2=2.74 $Y2=2.72
r106 22 40 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.625 $Y=2.72
+ $X2=1.61 $Y2=2.72
r107 22 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.625 $Y=2.72
+ $X2=1.79 $Y2=2.72
r108 21 43 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.53 $Y2=2.72
r109 21 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.79 $Y2=2.72
r110 17 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.865 $Y=2.635
+ $X2=3.865 $Y2=2.72
r111 17 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.865 $Y=2.635
+ $X2=3.865 $Y2=2.34
r112 13 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.79 $Y=2.635
+ $X2=1.79 $Y2=2.72
r113 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.79 $Y=2.635
+ $X2=1.79 $Y2=2.34
r114 4 19 600 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=1 $X=3.665
+ $Y=2.065 $X2=3.865 $Y2=2.34
r115 3 25 600 $w=1.7e-07 $l=3.49821e-07 $layer=licon1_PDIFF $count=1 $X=2.595
+ $Y=2.065 $X2=2.765 $Y2=2.34
r116 2 15 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=1.665
+ $Y=2.065 $X2=1.79 $Y2=2.34
r117 1 55 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.645
+ $Y=2.065 $X2=0.79 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_1%X 1 2 7 8 9 10 11 22 40 46
r19 25 46 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=4.38 $Y=1.575
+ $X2=4.38 $Y2=1.53
r20 20 40 0.664871 $w=2.58e-07 $l=1.5e-08 $layer=LI1_cond $X=4.38 $Y=0.695
+ $X2=4.38 $Y2=0.71
r21 11 42 18.6952 $w=2.23e-07 $l=3.65e-07 $layer=LI1_cond $X=4.397 $Y=1.19
+ $X2=4.397 $Y2=0.825
r22 10 30 11.0812 $w=2.58e-07 $l=2.5e-07 $layer=LI1_cond $X=4.38 $Y=2.21
+ $X2=4.38 $Y2=1.96
r23 9 30 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=4.38 $Y=1.87 $X2=4.38
+ $Y2=1.96
r24 8 46 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=4.38 $Y=1.51 $X2=4.38
+ $Y2=1.53
r25 8 11 9.60685 $w=3.83e-07 $l=2.55e-07 $layer=LI1_cond $X=4.397 $Y=1.445
+ $X2=4.397 $Y2=1.19
r26 8 9 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=4.38 $Y=1.595
+ $X2=4.38 $Y2=1.87
r27 8 25 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=4.38 $Y=1.595 $X2=4.38
+ $Y2=1.575
r28 7 42 3.78622 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=4.38 $Y=0.745 $X2=4.38
+ $Y2=0.825
r29 7 40 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=4.38 $Y=0.745
+ $X2=4.38 $Y2=0.71
r30 7 20 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=4.38 $Y=0.66 $X2=4.38
+ $Y2=0.695
r31 7 22 10.6379 $w=2.58e-07 $l=2.4e-07 $layer=LI1_cond $X=4.38 $Y=0.66 $X2=4.38
+ $Y2=0.42
r32 2 30 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.19
+ $Y=1.485 $X2=4.335 $Y2=1.96
r33 1 22 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.2
+ $Y=0.235 $X2=4.335 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_1%VGND 1 2 9 12 13 14 16 29 30 34
c49 9 0 1.48364e-19 $X=3.895 $Y=0.38
r50 34 37 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.765
+ $Y2=0.38
r51 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r52 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r53 27 30 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r54 26 27 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r55 24 27 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r56 24 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r57 23 26 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r58 23 24 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r59 21 34 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.765
+ $Y2=0
r60 21 23 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.15
+ $Y2=0
r61 16 34 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.765
+ $Y2=0
r62 16 18 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.23
+ $Y2=0
r63 14 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r64 14 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r65 12 26 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.81 $Y=0 $X2=3.45
+ $Y2=0
r66 12 13 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.81 $Y=0 $X2=3.895
+ $Y2=0
r67 11 29 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.98 $Y=0 $X2=4.37
+ $Y2=0
r68 11 13 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.98 $Y=0 $X2=3.895
+ $Y2=0
r69 7 13 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.895 $Y=0.085
+ $X2=3.895 $Y2=0
r70 7 9 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.895 $Y=0.085
+ $X2=3.895 $Y2=0.38
r71 2 9 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=3.675
+ $Y=0.465 $X2=3.895 $Y2=0.38
r72 1 37 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.605
+ $Y=0.235 $X2=0.79 $Y2=0.38
.ends

