# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a2bb2o_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445000 0.995000 1.815000 1.615000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.995000 2.335000 1.375000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.080000 0.765000 4.455000 1.655000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.300000 1.050000 3.760000 1.655000 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.600000 0.085000 ;
        RECT 0.185000  0.085000 0.355000 0.930000 ;
        RECT 1.000000  0.085000 1.480000 0.530000 ;
        RECT 2.155000  0.085000 2.890000 0.485000 ;
        RECT 3.905000  0.085000 4.355000 0.595000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 4.600000 2.805000 ;
        RECT 0.185000 1.445000 0.355000 2.635000 ;
        RECT 1.000000 2.235000 1.380000 2.635000 ;
        RECT 3.675000 2.175000 3.925000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 0.255000 0.830000 0.810000 ;
        RECT 0.525000 0.810000 0.745000 1.525000 ;
        RECT 0.525000 1.525000 0.830000 2.465000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.915000 0.995000 1.220000 1.325000 ;
      RECT 1.000000 1.325000 1.220000 1.805000 ;
      RECT 1.000000 1.805000 1.860000 1.975000 ;
      RECT 1.640000 1.975000 1.860000 2.200000 ;
      RECT 1.640000 2.200000 2.870000 2.370000 ;
      RECT 1.765000 0.255000 1.935000 0.655000 ;
      RECT 1.765000 0.655000 2.710000 0.825000 ;
      RECT 2.175000 1.545000 2.710000 1.715000 ;
      RECT 2.175000 1.715000 2.345000 1.905000 ;
      RECT 2.540000 0.825000 2.710000 1.545000 ;
      RECT 2.640000 1.895000 3.100000 2.065000 ;
      RECT 2.640000 2.065000 2.870000 2.200000 ;
      RECT 2.700000 2.370000 2.870000 2.465000 ;
      RECT 2.880000 0.700000 3.280000 0.870000 ;
      RECT 2.880000 0.870000 3.100000 1.895000 ;
      RECT 3.110000 0.255000 3.280000 0.700000 ;
      RECT 3.125000 2.255000 3.455000 2.425000 ;
      RECT 3.285000 1.835000 4.315000 2.005000 ;
      RECT 3.285000 2.005000 3.455000 2.255000 ;
      RECT 4.145000 2.005000 4.315000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a2bb2o_2
END LIBRARY
