* File: sky130_fd_sc_hdll__o21a_2.spice
* Created: Wed Sep  2 08:43:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o21a_2.pex.spice"
.subckt sky130_fd_sc_hdll__o21a_2  VNB VPB B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1005 N_X_M1005_d N_A_79_21#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.105625 AS=0.169 PD=0.975 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1005_d N_A_79_21#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.105625 AS=0.20475 PD=0.975 PS=1.93 NRD=0 NRS=9.228 M=1 R=4.33333
+ SA=75000.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_414_47#_M1002_d N_B1_M1002_g N_A_79_21#_M1002_s VNB NSHORT L=0.15
+ W=0.65 AD=0.091 AS=0.20475 PD=0.93 PS=1.93 NRD=0 NRS=9.228 M=1 R=4.33333
+ SA=75000.2 SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g N_A_414_47#_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.091 PD=1.18 PS=0.93 NRD=12.912 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1003 N_A_414_47#_M1003_d N_A1_M1003_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.20475 AS=0.17225 PD=1.93 PS=1.18 NRD=9.228 NRS=33.228 M=1 R=4.33333
+ SA=75001.3 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_X_M1001_d N_A_79_21#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1475 AS=0.27 PD=1.295 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.8 A=0.18 P=2.36 MULT=1
MM1006 N_X_M1001_d N_A_79_21#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1475 AS=0.41 PD=1.295 PS=1.82 NRD=1.9503 NRS=1.9503 M=1 R=5.55556
+ SA=90000.7 SB=90002.3 A=0.18 P=2.36 MULT=1
MM1000 N_A_79_21#_M1000_d N_B1_M1000_g N_VPWR_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.41 PD=1.3 PS=1.82 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.7
+ SB=90001.3 A=0.18 P=2.36 MULT=1
MM1007 A_508_297# N_A2_M1007_g N_A_79_21#_M1000_d VPB PHIGHVT L=0.18 W=1 AD=0.25
+ AS=0.15 PD=1.5 PS=1.3 NRD=38.3953 NRS=1.9503 M=1 R=5.55556 SA=90002.1
+ SB=90000.9 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g A_508_297# VPB PHIGHVT L=0.18 W=1 AD=0.275
+ AS=0.25 PD=2.55 PS=1.5 NRD=1.9503 NRS=38.3953 M=1 R=5.55556 SA=90002.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
pX11_noxref noxref_12 B1 B1 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o21a_2.pxi.spice"
*
.ends
*
*
