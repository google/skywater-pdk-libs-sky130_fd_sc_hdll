* File: sky130_fd_sc_hdll__or4bb_2.pex.spice
* Created: Thu Aug 27 19:25:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR4BB_2%C_N 2 3 5 8 9 10 14 15 16
c33 2 0 1.33125e-19 $X=0.495 $Y=1.875
r34 14 17 39.5599 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=0.547 $Y=1.16
+ $X2=0.547 $Y2=1.325
r35 14 16 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=0.547 $Y=1.16
+ $X2=0.547 $Y2=0.995
r36 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.16 $X2=0.53 $Y2=1.16
r37 9 10 9.79577 $w=3.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.63 $Y=1.19 $X2=0.63
+ $Y2=1.53
r38 9 15 0.864332 $w=3.98e-07 $l=3e-08 $layer=LI1_cond $X=0.63 $Y=1.19 $X2=0.63
+ $Y2=1.16
r39 8 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.56 $Y=0.675
+ $X2=0.56 $Y2=0.995
r40 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.975
+ $X2=0.495 $Y2=2.26
r41 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.875 $X2=0.495
+ $Y2=1.975
r42 2 17 182.367 $w=2e-07 $l=5.5e-07 $layer=POLY_cond $X=0.495 $Y=1.875
+ $X2=0.495 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_2%D_N 1 3 4 6 7 14
r34 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.085
+ $Y=1.16 $X2=1.085 $Y2=1.16
r35 7 14 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.255 $Y=1.16
+ $X2=1.085 $Y2=1.16
r36 4 10 46.2237 $w=3.35e-07 $l=2.89396e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.115 $Y2=1.16
r37 4 6 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.03 $Y=1.41 $X2=1.03
+ $Y2=1.695
r38 1 10 38.6365 $w=3.35e-07 $l=2.13014e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.115 $Y2=1.16
r39 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_2%A_216_93# 1 2 8 9 11 14 16 21 23 25 30 36
c69 16 0 1.33125e-19 $X=1.51 $Y=1.61
r70 35 36 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.04 $Y=1.16
+ $X2=2.065 $Y2=1.16
r71 31 35 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=1.77 $Y=1.16
+ $X2=2.04 $Y2=1.16
r72 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.77
+ $Y=1.16 $X2=1.77 $Y2=1.16
r73 27 30 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.605 $Y=1.16
+ $X2=1.77 $Y2=1.16
r74 25 26 17.5021 $w=2.37e-07 $l=3.4e-07 $layer=LI1_cond $X=1.265 $Y=0.655
+ $X2=1.605 $Y2=0.655
r75 22 27 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=1.245
+ $X2=1.605 $Y2=1.16
r76 22 23 16.3445 $w=1.88e-07 $l=2.8e-07 $layer=LI1_cond $X=1.605 $Y=1.245
+ $X2=1.605 $Y2=1.525
r77 21 27 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=1.075
+ $X2=1.605 $Y2=1.16
r78 20 26 2.03416 $w=1.9e-07 $l=1.7e-07 $layer=LI1_cond $X=1.605 $Y=0.825
+ $X2=1.605 $Y2=0.655
r79 20 21 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=1.605 $Y=0.825
+ $X2=1.605 $Y2=1.075
r80 16 23 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.51 $Y=1.61
+ $X2=1.605 $Y2=1.525
r81 16 18 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.51 $Y=1.61
+ $X2=1.265 $Y2=1.61
r82 12 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.065 $Y=0.995
+ $X2=2.065 $Y2=1.16
r83 12 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.065 $Y=0.995
+ $X2=2.065 $Y2=0.445
r84 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.04 $Y=1.99
+ $X2=2.04 $Y2=2.275
r85 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.04 $Y=1.89 $X2=2.04
+ $Y2=1.99
r86 7 35 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.04 $Y=1.325 $X2=2.04
+ $Y2=1.16
r87 7 8 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=2.04 $Y=1.325 $X2=2.04
+ $Y2=1.89
r88 2 18 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.485 $X2=1.265 $Y2=1.61
r89 1 25 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.465 $X2=1.265 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_2%A_27_410# 1 2 9 11 13 15 18 20 23 24 25 28
+ 34 36
c94 28 0 1.86536e-20 $X=2.485 $Y=1.16
r95 31 34 3.93367 $w=3.73e-07 $l=1.28e-07 $layer=LI1_cond $X=0.172 $Y=0.637
+ $X2=0.3 $Y2=0.637
r96 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.485
+ $Y=1.16 $X2=2.485 $Y2=1.16
r97 26 28 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.485 $Y=1.415
+ $X2=2.485 $Y2=1.16
r98 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.4 $Y=1.5
+ $X2=2.485 $Y2=1.415
r99 24 25 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.4 $Y=1.5 $X2=2.04
+ $Y2=1.5
r100 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.955 $Y=1.585
+ $X2=2.04 $Y2=1.5
r101 22 23 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.955 $Y=1.585
+ $X2=1.955 $Y2=1.865
r102 21 36 2.24312 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.95
+ $X2=0.215 $Y2=1.95
r103 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.87 $Y=1.95
+ $X2=1.955 $Y2=1.865
r104 20 21 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=1.87 $Y=1.95
+ $X2=0.345 $Y2=1.95
r105 16 36 4.18896 $w=2.17e-07 $l=8.5e-08 $layer=LI1_cond $X=0.215 $Y=2.035
+ $X2=0.215 $Y2=1.95
r106 16 18 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.215 $Y=2.035
+ $X2=0.215 $Y2=2.29
r107 15 36 4.18896 $w=2.17e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.172 $Y=1.865
+ $X2=0.215 $Y2=1.95
r108 14 31 5.2298 $w=1.75e-07 $l=1.88e-07 $layer=LI1_cond $X=0.172 $Y=0.825
+ $X2=0.172 $Y2=0.637
r109 14 15 65.9117 $w=1.73e-07 $l=1.04e-06 $layer=LI1_cond $X=0.172 $Y=0.825
+ $X2=0.172 $Y2=1.865
r110 11 29 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.57 $Y=1.41
+ $X2=2.51 $Y2=1.16
r111 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.57 $Y=1.41
+ $X2=2.57 $Y2=1.695
r112 7 29 38.578 $w=2.95e-07 $l=1.83916e-07 $layer=POLY_cond $X=2.55 $Y=0.995
+ $X2=2.51 $Y2=1.16
r113 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.55 $Y=0.995
+ $X2=2.55 $Y2=0.445
r114 2 18 600 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.05 $X2=0.26 $Y2=2.29
r115 1 34 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.465 $X2=0.3 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_2%B 1 2 3 4 6 9 10 11 17
c43 6 0 1.86536e-20 $X=2.98 $Y=1.695
c44 2 0 8.49032e-20 $X=2.98 $Y=1.31
c45 1 0 1.42379e-20 $X=2.98 $Y=0.86
r46 15 17 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=3.045 $Y=2.29
+ $X2=3.015 $Y2=2.29
r47 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.045
+ $Y=2.335 $X2=3.045 $Y2=2.335
r48 11 15 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=3.265 $Y=2.29
+ $X2=3.045 $Y2=2.29
r49 9 10 101.22 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=3.005 $Y=0.445
+ $X2=3.005 $Y2=0.76
r50 4 14 56.473 $w=2.93e-07 $l=3.3541e-07 $layer=POLY_cond $X=2.98 $Y=2.035
+ $X2=3.055 $Y2=2.335
r51 4 6 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=2.98 $Y=2.035 $X2=2.98
+ $Y2=1.695
r52 3 6 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.98 $Y=1.41 $X2=2.98
+ $Y2=1.695
r53 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.98 $Y=1.31 $X2=2.98
+ $Y2=1.41
r54 1 10 37.4512 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.98 $Y=0.86 $X2=2.98
+ $Y2=0.76
r55 1 2 149.21 $w=2e-07 $l=4.5e-07 $layer=POLY_cond $X=2.98 $Y=0.86 $X2=2.98
+ $Y2=1.31
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_2%A 1 3 6 8 12 14
c39 1 0 1.97843e-19 $X=3.465 $Y=1.41
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.425
+ $Y=1.16 $X2=3.425 $Y2=1.16
r41 8 12 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=3.265 $Y=1.16
+ $X2=3.425 $Y2=1.16
r42 8 14 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.265 $Y=1.16
+ $X2=3.015 $Y2=1.16
r43 4 11 38.578 $w=2.95e-07 $l=1.83916e-07 $layer=POLY_cond $X=3.49 $Y=0.995
+ $X2=3.45 $Y2=1.16
r44 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.49 $Y=0.995 $X2=3.49
+ $Y2=0.445
r45 1 11 48.1208 $w=2.95e-07 $l=2.57391e-07 $layer=POLY_cond $X=3.465 $Y=1.41
+ $X2=3.45 $Y2=1.16
r46 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.465 $Y=1.41
+ $X2=3.465 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_2%A_336_413# 1 2 3 10 12 13 15 16 18 19 21
+ 22 28 31 32 33 34 35 38 40 42 47 48 49 54 56 61
c129 54 0 1.14153e-19 $X=3.955 $Y=1.16
c130 47 0 1.07404e-19 $X=3.85 $Y=1.495
c131 34 0 1.97843e-19 $X=3.225 $Y=1.87
r132 61 62 3.21333 $w=3.75e-07 $l=2.5e-08 $layer=POLY_cond $X=4.475 $Y=1.202
+ $X2=4.5 $Y2=1.202
r133 60 61 57.1973 $w=3.75e-07 $l=4.45e-07 $layer=POLY_cond $X=4.03 $Y=1.202
+ $X2=4.475 $Y2=1.202
r134 59 60 3.21333 $w=3.75e-07 $l=2.5e-08 $layer=POLY_cond $X=4.005 $Y=1.202
+ $X2=4.03 $Y2=1.202
r135 55 59 6.42667 $w=3.75e-07 $l=5e-08 $layer=POLY_cond $X=3.955 $Y=1.202
+ $X2=4.005 $Y2=1.202
r136 54 57 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=3.902 $Y=1.16
+ $X2=3.902 $Y2=1.325
r137 54 56 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=3.902 $Y=1.16
+ $X2=3.902 $Y2=0.995
r138 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.955
+ $Y=1.16 $X2=3.955 $Y2=1.16
r139 49 51 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.31 $Y=1.58
+ $X2=3.31 $Y2=1.87
r140 47 57 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.85 $Y=1.495
+ $X2=3.85 $Y2=1.325
r141 44 56 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.85 $Y=0.825
+ $X2=3.85 $Y2=0.995
r142 43 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.395 $Y=1.58
+ $X2=3.31 $Y2=1.58
r143 42 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.765 $Y=1.58
+ $X2=3.85 $Y2=1.495
r144 42 43 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.765 $Y=1.58
+ $X2=3.395 $Y2=1.58
r145 41 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.315 $Y=0.74
+ $X2=3.23 $Y2=0.74
r146 40 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.765 $Y=0.74
+ $X2=3.85 $Y2=0.825
r147 40 41 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.765 $Y=0.74
+ $X2=3.315 $Y2=0.74
r148 36 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.23 $Y=0.655
+ $X2=3.23 $Y2=0.74
r149 36 38 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.23 $Y=0.655
+ $X2=3.23 $Y2=0.47
r150 34 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.225 $Y=1.87
+ $X2=3.31 $Y2=1.87
r151 34 35 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=3.225 $Y=1.87
+ $X2=2.43 $Y2=1.87
r152 32 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.145 $Y=0.74
+ $X2=3.23 $Y2=0.74
r153 32 33 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=3.145 $Y=0.74
+ $X2=2.36 $Y2=0.74
r154 30 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.345 $Y=1.955
+ $X2=2.43 $Y2=1.87
r155 30 31 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.345 $Y=1.955
+ $X2=2.345 $Y2=2.205
r156 26 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.275 $Y=0.655
+ $X2=2.36 $Y2=0.74
r157 26 28 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.275 $Y=0.655
+ $X2=2.275 $Y2=0.47
r158 22 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.26 $Y=2.29
+ $X2=2.345 $Y2=2.205
r159 22 24 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.26 $Y=2.29
+ $X2=1.805 $Y2=2.29
r160 19 62 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.5 $Y=0.995
+ $X2=4.5 $Y2=1.202
r161 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.5 $Y=0.995
+ $X2=4.5 $Y2=0.56
r162 16 61 19.9308 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.475 $Y=1.41
+ $X2=4.475 $Y2=1.202
r163 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.475 $Y=1.41
+ $X2=4.475 $Y2=1.985
r164 13 60 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.03 $Y=0.995
+ $X2=4.03 $Y2=1.202
r165 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.03 $Y=0.995
+ $X2=4.03 $Y2=0.56
r166 10 59 19.9308 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.005 $Y=1.41
+ $X2=4.005 $Y2=1.202
r167 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.005 $Y=1.41
+ $X2=4.005 $Y2=1.985
r168 3 24 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=1.68
+ $Y=2.065 $X2=1.805 $Y2=2.29
r169 2 38 182 $w=1.7e-07 $l=3.00791e-07 $layer=licon1_NDIFF $count=1 $X=3.08
+ $Y=0.235 $X2=3.23 $Y2=0.47
r170 1 28 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=2.14
+ $Y=0.235 $X2=2.275 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_2%VPWR 1 2 3 12 16 18 20 25 26 27 29 41 46
+ 50
c58 2 0 1.07404e-19 $X=3.555 $Y=1.485
r59 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r60 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 44 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r62 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r63 41 49 3.40825 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=4.65 $Y=2.72
+ $X2=4.855 $Y2=2.72
r64 41 43 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.65 $Y=2.72
+ $X2=4.37 $Y2=2.72
r65 40 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r66 39 40 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r67 37 40 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r68 37 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 36 39 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r70 36 37 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r71 34 46 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r72 34 36 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r73 29 46 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r74 29 31 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r75 27 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r76 27 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r77 25 39 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=2.72
+ $X2=3.45 $Y2=2.72
r78 25 26 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.615 $Y=2.72
+ $X2=3.755 $Y2=2.72
r79 24 43 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.895 $Y=2.72
+ $X2=4.37 $Y2=2.72
r80 24 26 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.895 $Y=2.72
+ $X2=3.755 $Y2=2.72
r81 20 23 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.735 $Y=1.66
+ $X2=4.735 $Y2=2.34
r82 18 49 3.40825 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=4.735 $Y=2.635
+ $X2=4.855 $Y2=2.72
r83 18 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.735 $Y=2.635
+ $X2=4.735 $Y2=2.34
r84 14 26 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.755 $Y=2.635
+ $X2=3.755 $Y2=2.72
r85 14 16 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=3.755 $Y=2.635
+ $X2=3.755 $Y2=2
r86 10 46 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r87 10 12 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.29
r88 3 23 400 $w=1.7e-07 $l=9.36149e-07 $layer=licon1_PDIFF $count=1 $X=4.565
+ $Y=1.485 $X2=4.735 $Y2=2.34
r89 3 20 400 $w=1.7e-07 $l=2.45713e-07 $layer=licon1_PDIFF $count=1 $X=4.565
+ $Y=1.485 $X2=4.735 $Y2=1.66
r90 2 16 300 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=2 $X=3.555
+ $Y=1.485 $X2=3.765 $Y2=2
r91 1 12 600 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.05 $X2=0.73 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_2%X 1 2 12 14 15 16
r26 14 16 7.68295 $w=2.98e-07 $l=2e-07 $layer=LI1_cond $X=4.305 $Y=1.645
+ $X2=4.305 $Y2=1.845
r27 14 15 7.17198 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=4.305 $Y=1.645
+ $X2=4.305 $Y2=1.495
r28 10 12 3.90828 $w=3.43e-07 $l=1.17e-07 $layer=LI1_cond $X=4.24 $Y=0.587
+ $X2=4.357 $Y2=0.587
r29 7 12 4.09374 $w=1.95e-07 $l=1.73e-07 $layer=LI1_cond $X=4.357 $Y=0.76
+ $X2=4.357 $Y2=0.587
r30 7 15 41.8042 $w=1.93e-07 $l=7.35e-07 $layer=LI1_cond $X=4.357 $Y=0.76
+ $X2=4.357 $Y2=1.495
r31 2 16 300 $w=1.7e-07 $l=4.2638e-07 $layer=licon1_PDIFF $count=2 $X=4.095
+ $Y=1.485 $X2=4.24 $Y2=1.845
r32 1 10 182 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_NDIFF $count=1 $X=4.105
+ $Y=0.235 $X2=4.24 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_2%VGND 1 2 3 4 5 18 20 24 28 30 32 34 35 37
+ 38 39 40 46 59 64 68 70
c77 40 0 1.42379e-20 $X=3.485 $Y=0
r78 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r79 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r80 62 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r81 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r82 59 67 3.40825 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=4.65 $Y=0 $X2=4.855
+ $Y2=0
r83 59 61 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.65 $Y=0 $X2=4.37
+ $Y2=0
r84 58 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r85 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r86 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r87 55 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r88 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r89 52 64 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=1.97 $Y=0 $X2=1.782
+ $Y2=0
r90 52 54 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.97 $Y=0 $X2=2.53
+ $Y2=0
r91 50 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r92 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r93 46 50 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r94 46 70 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r95 42 61 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.915 $Y=0 $X2=4.37
+ $Y2=0
r96 40 57 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.485 $Y=0 $X2=3.45
+ $Y2=0
r97 39 44 10.7204 $w=4.28e-07 $l=4e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.7
+ $Y2=0.4
r98 39 42 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.915
+ $Y2=0
r99 39 40 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.485
+ $Y2=0
r100 37 54 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.545 $Y=0 $X2=2.53
+ $Y2=0
r101 37 38 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.545 $Y=0 $X2=2.735
+ $Y2=0
r102 36 57 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.925 $Y=0
+ $X2=3.45 $Y2=0
r103 36 38 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=2.735
+ $Y2=0
r104 34 49 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=0.71 $Y=0 $X2=0.69
+ $Y2=0
r105 34 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0 $X2=0.795
+ $Y2=0
r106 30 67 3.40825 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=4.735 $Y=0.085
+ $X2=4.855 $Y2=0
r107 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.735 $Y=0.085
+ $X2=4.735 $Y2=0.39
r108 26 38 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=0.085
+ $X2=2.735 $Y2=0
r109 26 28 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.735 $Y=0.085
+ $X2=2.735 $Y2=0.4
r110 22 64 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.782 $Y=0.085
+ $X2=1.782 $Y2=0
r111 22 24 9.68052 $w=3.73e-07 $l=3.15e-07 $layer=LI1_cond $X=1.782 $Y=0.085
+ $X2=1.782 $Y2=0.4
r112 21 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.795
+ $Y2=0
r113 20 64 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=1.595 $Y=0
+ $X2=1.782 $Y2=0
r114 20 21 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.595 $Y=0
+ $X2=0.88 $Y2=0
r115 16 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0
r116 16 18 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0.66
r117 5 32 91 $w=1.7e-07 $l=2.24499e-07 $layer=licon1_NDIFF $count=2 $X=4.575
+ $Y=0.235 $X2=4.735 $Y2=0.39
r118 4 44 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.565
+ $Y=0.235 $X2=3.75 $Y2=0.4
r119 3 28 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.625
+ $Y=0.235 $X2=2.76 $Y2=0.4
r120 2 24 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=1.66
+ $Y=0.235 $X2=1.785 $Y2=0.4
r121 1 18 182 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_NDIFF $count=1 $X=0.635
+ $Y=0.465 $X2=0.795 $Y2=0.66
.ends

