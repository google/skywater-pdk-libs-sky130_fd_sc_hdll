* File: sky130_fd_sc_hdll__or4bb_1.pex.spice
* Created: Wed Sep  2 08:49:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR4BB_1%C_N 2 3 5 8 9 10 14 16
c33 2 0 1.38252e-19 $X=0.495 $Y=1.875
r34 14 17 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.16
+ $X2=0.53 $Y2=1.325
r35 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.16
+ $X2=0.53 $Y2=0.995
r36 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.16 $X2=0.53 $Y2=1.16
r37 9 10 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.617 $Y=1.53
+ $X2=0.617 $Y2=1.16
r38 8 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.555 $Y=0.675
+ $X2=0.555 $Y2=0.995
r39 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.975
+ $X2=0.495 $Y2=2.26
r40 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.875 $X2=0.495
+ $Y2=1.975
r41 2 17 182.367 $w=2e-07 $l=5.5e-07 $layer=POLY_cond $X=0.495 $Y=1.875
+ $X2=0.495 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_1%D_N 1 3 4 6 7 14
r34 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.065
+ $Y=1.16 $X2=1.065 $Y2=1.16
r35 7 14 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.25 $Y=1.16
+ $X2=1.065 $Y2=1.16
r36 4 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.065 $Y2=1.16
r37 4 6 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.03 $Y=1.41 $X2=1.03
+ $Y2=1.695
r38 1 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.065 $Y2=1.16
r39 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_1%A_216_93# 1 2 8 9 11 14 16 21 23 26 27 30
+ 32
c68 27 0 1.69441e-19 $X=1.97 $Y=1.16
c69 16 0 1.38252e-19 $X=1.505 $Y=1.61
r70 30 31 16.8452 $w=2.39e-07 $l=3.3e-07 $layer=LI1_cond $X=1.26 $Y=0.655
+ $X2=1.59 $Y2=0.655
r71 27 35 40.3353 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.975 $Y=1.16
+ $X2=1.975 $Y2=1.325
r72 27 34 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.975 $Y=1.16
+ $X2=1.975 $Y2=0.995
r73 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.97
+ $Y=1.16 $X2=1.97 $Y2=1.16
r74 24 32 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.675 $Y=1.16
+ $X2=1.59 $Y2=1.16
r75 24 26 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.675 $Y=1.16
+ $X2=1.97 $Y2=1.16
r76 22 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=1.245
+ $X2=1.59 $Y2=1.16
r77 22 23 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.59 $Y=1.245
+ $X2=1.59 $Y2=1.525
r78 21 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=1.075
+ $X2=1.59 $Y2=1.16
r79 20 31 2.73298 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.59 $Y=0.825
+ $X2=1.59 $Y2=0.655
r80 20 21 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.59 $Y=0.825
+ $X2=1.59 $Y2=1.075
r81 16 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.505 $Y=1.61
+ $X2=1.59 $Y2=1.525
r82 16 18 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.505 $Y=1.61
+ $X2=1.265 $Y2=1.61
r83 14 34 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.04 $Y=0.445
+ $X2=2.04 $Y2=0.995
r84 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.015 $Y=1.99
+ $X2=2.015 $Y2=2.275
r85 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.015 $Y=1.89 $X2=2.015
+ $Y2=1.99
r86 8 35 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=2.015 $Y=1.89
+ $X2=2.015 $Y2=1.325
r87 2 18 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.485 $X2=1.265 $Y2=1.61
r88 1 30 182 $w=1.7e-07 $l=2.70416e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.465 $X2=1.26 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_1%A_27_410# 1 2 9 11 13 15 18 20 23 24 25 28
+ 34 36
c92 28 0 1.86536e-20 $X=2.46 $Y=1.16
c93 20 0 1.69441e-19 $X=1.845 $Y=1.95
r94 31 34 3.84148 $w=3.73e-07 $l=1.25e-07 $layer=LI1_cond $X=0.17 $Y=0.637
+ $X2=0.295 $Y2=0.637
r95 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.46
+ $Y=1.16 $X2=2.46 $Y2=1.16
r96 26 28 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.46 $Y=1.415
+ $X2=2.46 $Y2=1.16
r97 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.375 $Y=1.5
+ $X2=2.46 $Y2=1.415
r98 24 25 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.375 $Y=1.5
+ $X2=2.015 $Y2=1.5
r99 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.93 $Y=1.585
+ $X2=2.015 $Y2=1.5
r100 22 23 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.93 $Y=1.585
+ $X2=1.93 $Y2=1.865
r101 21 36 2.20034 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.95
+ $X2=0.215 $Y2=1.95
r102 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.845 $Y=1.95
+ $X2=1.93 $Y2=1.865
r103 20 21 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=1.845 $Y=1.95
+ $X2=0.345 $Y2=1.95
r104 16 36 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.215 $Y=2.035
+ $X2=0.215 $Y2=1.95
r105 16 18 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.215 $Y=2.035
+ $X2=0.215 $Y2=2.29
r106 15 36 4.23118 $w=2.15e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.17 $Y=1.865
+ $X2=0.215 $Y2=1.95
r107 14 31 5.38787 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=0.637
r108 14 15 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=1.865
r109 11 29 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.545 $Y=1.41
+ $X2=2.485 $Y2=1.16
r110 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.545 $Y=1.41
+ $X2=2.545 $Y2=1.695
r111 7 29 38.578 $w=2.95e-07 $l=1.83916e-07 $layer=POLY_cond $X=2.525 $Y=0.995
+ $X2=2.485 $Y2=1.16
r112 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.525 $Y=0.995
+ $X2=2.525 $Y2=0.445
r113 2 18 600 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.05 $X2=0.26 $Y2=2.29
r114 1 34 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.465 $X2=0.295 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_1%B 1 2 3 4 6 9 10 11 17
c43 6 0 1.86536e-20 $X=2.955 $Y=1.695
c44 2 0 8.49032e-20 $X=2.955 $Y=1.31
c45 1 0 1.42379e-20 $X=2.955 $Y=0.86
r46 14 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=2.335 $X2=2.99 $Y2=2.335
r47 11 17 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.24 $Y=2.29
+ $X2=2.99 $Y2=2.29
r48 9 10 101.22 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=2.98 $Y=0.445
+ $X2=2.98 $Y2=0.76
r49 4 14 61.8547 $w=2.49e-07 $l=3.17017e-07 $layer=POLY_cond $X=2.955 $Y=2.035
+ $X2=2.99 $Y2=2.335
r50 4 6 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=2.955 $Y=2.035
+ $X2=2.955 $Y2=1.695
r51 3 6 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.955 $Y=1.41
+ $X2=2.955 $Y2=1.695
r52 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.955 $Y=1.31 $X2=2.955
+ $Y2=1.41
r53 1 10 37.4512 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.955 $Y=0.86 $X2=2.955
+ $Y2=0.76
r54 1 2 149.21 $w=2e-07 $l=4.5e-07 $layer=POLY_cond $X=2.955 $Y=0.86 $X2=2.955
+ $Y2=1.31
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_1%A 1 3 6 8 12 14
c38 1 0 1.97843e-19 $X=3.44 $Y=1.41
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.405
+ $Y=1.16 $X2=3.405 $Y2=1.16
r40 8 12 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.24 $Y=1.16
+ $X2=3.405 $Y2=1.16
r41 8 14 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.24 $Y=1.16 $X2=2.99
+ $Y2=1.16
r42 4 11 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.465 $Y=0.995
+ $X2=3.405 $Y2=1.16
r43 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.465 $Y=0.995
+ $X2=3.465 $Y2=0.445
r44 1 11 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.44 $Y=1.41
+ $X2=3.405 $Y2=1.16
r45 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.44 $Y=1.41 $X2=3.44
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_1%A_331_413# 1 2 3 10 12 13 15 16 22 25 26
+ 27 28 29 32 34 36 41 42 43 48 50
c110 48 0 1.16645e-19 $X=3.945 $Y=1.16
c111 41 0 1.07404e-19 $X=3.825 $Y=1.495
c112 28 0 1.97843e-19 $X=3.2 $Y=1.87
r113 48 51 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=1.16
+ $X2=3.885 $Y2=1.325
r114 48 50 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=1.16
+ $X2=3.885 $Y2=0.995
r115 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.945
+ $Y=1.16 $X2=3.945 $Y2=1.16
r116 43 45 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.285 $Y=1.58
+ $X2=3.285 $Y2=1.87
r117 41 51 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.825 $Y=1.495
+ $X2=3.825 $Y2=1.325
r118 38 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.825 $Y=0.825
+ $X2=3.825 $Y2=0.995
r119 37 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.37 $Y=1.58
+ $X2=3.285 $Y2=1.58
r120 36 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.74 $Y=1.58
+ $X2=3.825 $Y2=1.495
r121 36 37 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.74 $Y=1.58
+ $X2=3.37 $Y2=1.58
r122 35 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.29 $Y=0.74
+ $X2=3.205 $Y2=0.74
r123 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.74 $Y=0.74
+ $X2=3.825 $Y2=0.825
r124 34 35 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.74 $Y=0.74
+ $X2=3.29 $Y2=0.74
r125 30 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.205 $Y=0.655
+ $X2=3.205 $Y2=0.74
r126 30 32 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.205 $Y=0.655
+ $X2=3.205 $Y2=0.47
r127 28 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=1.87
+ $X2=3.285 $Y2=1.87
r128 28 29 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=3.2 $Y=1.87
+ $X2=2.405 $Y2=1.87
r129 26 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=0.74
+ $X2=3.205 $Y2=0.74
r130 26 27 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=3.12 $Y=0.74
+ $X2=2.335 $Y2=0.74
r131 24 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.32 $Y=1.955
+ $X2=2.405 $Y2=1.87
r132 24 25 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.32 $Y=1.955
+ $X2=2.32 $Y2=2.205
r133 20 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.25 $Y=0.655
+ $X2=2.335 $Y2=0.74
r134 20 22 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.25 $Y=0.655
+ $X2=2.25 $Y2=0.47
r135 16 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.235 $Y=2.29
+ $X2=2.32 $Y2=2.205
r136 16 18 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.235 $Y=2.29
+ $X2=1.78 $Y2=2.29
r137 13 49 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=4.005 $Y=0.995
+ $X2=3.945 $Y2=1.16
r138 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.005 $Y=0.995
+ $X2=4.005 $Y2=0.56
r139 10 49 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.98 $Y=1.41
+ $X2=3.945 $Y2=1.16
r140 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.98 $Y=1.41
+ $X2=3.98 $Y2=1.985
r141 3 18 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=1.655
+ $Y=2.065 $X2=1.78 $Y2=2.29
r142 2 32 182 $w=1.7e-07 $l=3.00791e-07 $layer=licon1_NDIFF $count=1 $X=3.055
+ $Y=0.235 $X2=3.205 $Y2=0.47
r143 1 22 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=2.115
+ $Y=0.235 $X2=2.25 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_1%VPWR 1 2 9 13 16 17 18 20 33 34 37
c50 2 0 1.07404e-19 $X=3.53 $Y=1.485
r51 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r53 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r54 30 31 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r55 28 31 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r56 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r57 27 30 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r58 27 28 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r59 25 37 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r60 25 27 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r61 20 37 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r62 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r63 18 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r64 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r65 16 30 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.59 $Y=2.72
+ $X2=3.45 $Y2=2.72
r66 16 17 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.59 $Y=2.72 $X2=3.73
+ $Y2=2.72
r67 15 33 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.87 $Y=2.72 $X2=4.37
+ $Y2=2.72
r68 15 17 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.87 $Y=2.72 $X2=3.73
+ $Y2=2.72
r69 11 17 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.73 $Y=2.635
+ $X2=3.73 $Y2=2.72
r70 11 13 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=3.73 $Y=2.635
+ $X2=3.73 $Y2=2
r71 7 37 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r72 7 9 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.29
r73 2 13 300 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=2 $X=3.53
+ $Y=1.485 $X2=3.74 $Y2=2
r74 1 9 600 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.05 $X2=0.73 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_1%X 1 2 10 13 14 15
r18 13 15 6.66644 $w=3.23e-07 $l=1.88e-07 $layer=LI1_cond $X=4.292 $Y=1.657
+ $X2=4.292 $Y2=1.845
r19 13 14 6.95351 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=4.292 $Y=1.657
+ $X2=4.292 $Y2=1.495
r20 12 14 38.5021 $w=2.18e-07 $l=7.35e-07 $layer=LI1_cond $X=4.345 $Y=0.76
+ $X2=4.345 $Y2=1.495
r21 10 12 7.23718 $w=3.23e-07 $l=1.7e-07 $layer=LI1_cond $X=4.292 $Y=0.59
+ $X2=4.292 $Y2=0.76
r22 2 15 300 $w=1.7e-07 $l=4.2638e-07 $layer=licon1_PDIFF $count=2 $X=4.07
+ $Y=1.485 $X2=4.215 $Y2=1.845
r23 1 10 182 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_NDIFF $count=1 $X=4.08
+ $Y=0.235 $X2=4.215 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_1%VGND 1 2 3 4 15 17 21 23 27 29 30 31 32 38
+ 49 50 53 56
c69 32 0 1.42379e-20 $X=3.46 $Y=0
r70 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r71 54 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r72 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r73 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r74 47 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r75 47 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r76 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r77 44 56 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.9 $Y=0 $X2=2.71
+ $Y2=0
r78 44 46 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.9 $Y=0 $X2=3.45
+ $Y2=0
r79 42 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r80 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r81 38 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r82 34 49 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=4.37
+ $Y2=0
r83 32 46 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=3.46 $Y=0 $X2=3.45
+ $Y2=0
r84 31 36 10.7204 $w=4.28e-07 $l=4e-07 $layer=LI1_cond $X=3.675 $Y=0 $X2=3.675
+ $Y2=0.4
r85 31 34 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=3.675 $Y=0 $X2=3.89
+ $Y2=0
r86 31 32 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=3.675 $Y=0 $X2=3.46
+ $Y2=0
r87 29 41 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.705 $Y=0 $X2=0.69
+ $Y2=0
r88 29 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0 $X2=0.79
+ $Y2=0
r89 25 56 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=0.085
+ $X2=2.71 $Y2=0
r90 25 27 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.71 $Y=0.085
+ $X2=2.71 $Y2=0.4
r91 24 53 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=1.757
+ $Y2=0
r92 23 56 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.52 $Y=0 $X2=2.71
+ $Y2=0
r93 23 24 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.52 $Y=0 $X2=1.945
+ $Y2=0
r94 19 53 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.757 $Y=0.085
+ $X2=1.757 $Y2=0
r95 19 21 9.68052 $w=3.73e-07 $l=3.15e-07 $layer=LI1_cond $X=1.757 $Y=0.085
+ $X2=1.757 $Y2=0.4
r96 18 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.79
+ $Y2=0
r97 17 53 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=1.57 $Y=0 $X2=1.757
+ $Y2=0
r98 17 18 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.57 $Y=0 $X2=0.875
+ $Y2=0
r99 13 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r100 13 15 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.66
r101 4 36 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.54
+ $Y=0.235 $X2=3.725 $Y2=0.4
r102 3 27 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.6
+ $Y=0.235 $X2=2.735 $Y2=0.4
r103 2 21 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=1.655
+ $Y=0.235 $X2=1.78 $Y2=0.4
r104 1 15 182 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_NDIFF $count=1 $X=0.63
+ $Y=0.465 $X2=0.79 $Y2=0.66
.ends

