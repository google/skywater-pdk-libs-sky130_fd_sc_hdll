* NGSPICE file created from sky130_fd_sc_hdll__mux2_8.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__mux2_8 A0 A1 S VGND VNB VPB VPWR X
M1000 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=2.16e+12p pd=1.832e+07u as=1.16e+12p ps=1.032e+07u
M1001 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_870_297# A0 a_79_21# VPB phighvt w=1e+06u l=180000u
+  ad=1.385e+12p pd=6.77e+06u as=5.8e+11p ps=5.16e+06u
M1003 a_79_21# A1 a_872_47# VNB nshort w=640000u l=150000u
+  ad=4.096e+11p pd=3.84e+06u as=9.568e+11p ps=5.55e+06u
M1004 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_872_47# A1 a_79_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=8.645e+11p pd=7.86e+06u as=1.5084e+12p ps=1.374e+07u
M1007 VGND S a_872_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_1369_199# a_1422_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.0464e+12p ps=5.83e+06u
M1012 a_79_21# A0 a_870_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_1369_199# a_1420_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.675e+12p ps=7.35e+06u
M1014 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1420_297# a_1369_199# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1420_297# A1 a_79_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_79_21# A0 a_1422_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1369_199# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1020 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_870_297# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_872_47# S VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_79_21# A1 a_1420_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1422_47# a_1369_199# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1422_47# A0 a_79_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1369_199# S VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=0p ps=0u
M1033 VPWR S a_870_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

