* File: sky130_fd_sc_hdll__muxb4to1_2.pxi.spice
* Created: Thu Aug 27 19:11:52 2020
* 
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%D[0] N_D[0]_M1002_g N_D[0]_M1013_g
+ N_D[0]_M1026_g N_D[0]_M1017_g D[0] N_D[0]_c_219_n N_D[0]_c_220_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%D[0]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_278_265# N_A_278_265#_M1021_s
+ N_A_278_265#_M1006_s N_A_278_265#_M1005_g N_A_278_265#_c_267_n
+ N_A_278_265#_c_268_n N_A_278_265#_M1009_g N_A_278_265#_c_262_n
+ N_A_278_265#_c_263_n N_A_278_265#_c_270_n N_A_278_265#_c_264_n
+ N_A_278_265#_c_265_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_278_265#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%S[0] N_S[0]_c_339_n N_S[0]_M1011_g
+ N_S[0]_c_340_n N_S[0]_c_341_n N_S[0]_c_342_n N_S[0]_M1014_g N_S[0]_c_343_n
+ N_S[0]_c_344_n N_S[0]_c_345_n N_S[0]_c_346_n N_S[0]_c_347_n N_S[0]_M1006_g
+ N_S[0]_c_348_n N_S[0]_M1021_g N_S[0]_c_349_n S[0]
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%S[0]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%S[1] N_S[1]_c_404_n N_S[1]_M1018_g
+ N_S[1]_c_405_n N_S[1]_M1022_g N_S[1]_c_406_n N_S[1]_c_407_n N_S[1]_c_408_n
+ N_S[1]_c_409_n N_S[1]_c_410_n N_S[1]_M1010_g N_S[1]_c_411_n N_S[1]_c_412_n
+ N_S[1]_M1012_g N_S[1]_c_413_n S[1] PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%S[1]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_701_47# N_A_701_47#_M1018_d
+ N_A_701_47#_M1022_d N_A_701_47#_M1020_g N_A_701_47#_c_471_n
+ N_A_701_47#_c_466_n N_A_701_47#_M1027_g N_A_701_47#_c_474_n
+ N_A_701_47#_c_467_n N_A_701_47#_c_468_n N_A_701_47#_c_469_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_701_47#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%D[1] N_D[1]_M1015_g N_D[1]_M1019_g
+ N_D[1]_M1024_g N_D[1]_M1023_g D[1] N_D[1]_c_545_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%D[1]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%D[2] N_D[2]_M1000_g N_D[2]_M1028_g
+ N_D[2]_M1033_g N_D[2]_M1030_g D[2] N_D[2]_c_597_n N_D[2]_c_598_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%D[2]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_1566_265# N_A_1566_265#_M1038_s
+ N_A_1566_265#_M1035_s N_A_1566_265#_M1003_g N_A_1566_265#_c_652_n
+ N_A_1566_265#_c_653_n N_A_1566_265#_M1031_g N_A_1566_265#_c_647_n
+ N_A_1566_265#_c_648_n N_A_1566_265#_c_655_n N_A_1566_265#_c_649_n
+ N_A_1566_265#_c_650_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_1566_265#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%S[2] N_S[2]_c_725_n N_S[2]_M1029_g
+ N_S[2]_c_726_n N_S[2]_c_727_n N_S[2]_c_728_n N_S[2]_M1037_g N_S[2]_c_729_n
+ N_S[2]_c_730_n N_S[2]_c_731_n N_S[2]_c_732_n N_S[2]_c_733_n N_S[2]_M1035_g
+ N_S[2]_c_734_n N_S[2]_M1038_g N_S[2]_c_735_n S[2]
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%S[2]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%S[3] N_S[3]_c_790_n N_S[3]_M1007_g
+ N_S[3]_c_791_n N_S[3]_M1016_g N_S[3]_c_792_n N_S[3]_c_793_n N_S[3]_c_794_n
+ N_S[3]_c_795_n N_S[3]_c_796_n N_S[3]_M1025_g N_S[3]_c_797_n N_S[3]_c_798_n
+ N_S[3]_M1034_g N_S[3]_c_799_n S[3] PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%S[3]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_1989_47# N_A_1989_47#_M1007_d
+ N_A_1989_47#_M1016_d N_A_1989_47#_M1004_g N_A_1989_47#_c_857_n
+ N_A_1989_47#_c_852_n N_A_1989_47#_M1032_g N_A_1989_47#_c_860_n
+ N_A_1989_47#_c_853_n N_A_1989_47#_c_854_n N_A_1989_47#_c_855_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_1989_47#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%D[3] N_D[3]_M1001_g N_D[3]_M1008_g
+ N_D[3]_M1039_g N_D[3]_M1036_g D[3] N_D[3]_c_930_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%D[3]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_27_297# N_A_27_297#_M1002_d
+ N_A_27_297#_M1017_d N_A_27_297#_M1009_d N_A_27_297#_c_971_n
+ N_A_27_297#_c_977_n N_A_27_297#_c_981_n N_A_27_297#_c_985_n
+ N_A_27_297#_c_993_p N_A_27_297#_c_972_n N_A_27_297#_c_973_n
+ N_A_27_297#_c_974_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%VPWR N_VPWR_M1002_s N_VPWR_M1006_d
+ N_VPWR_M1015_s N_VPWR_M1000_d N_VPWR_M1035_d N_VPWR_M1001_d N_VPWR_c_1019_n
+ N_VPWR_c_1020_n N_VPWR_c_1021_n N_VPWR_c_1022_n N_VPWR_c_1023_n
+ N_VPWR_c_1024_n N_VPWR_c_1041_n N_VPWR_c_1025_n N_VPWR_c_1026_n
+ N_VPWR_c_1077_n N_VPWR_c_1085_n N_VPWR_c_1027_n N_VPWR_c_1028_n
+ N_VPWR_c_1121_n VPWR VPWR VPWR VPWR N_VPWR_c_1030_n N_VPWR_c_1031_n
+ N_VPWR_c_1032_n N_VPWR_c_1033_n N_VPWR_c_1034_n N_VPWR_c_1035_n
+ N_VPWR_c_1036_n N_VPWR_c_1037_n N_VPWR_c_1038_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%VPWR
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%Z N_Z_M1011_s N_Z_M1010_s N_Z_M1029_d
+ N_Z_M1025_d N_Z_M1005_s N_Z_M1020_s N_Z_M1003_d N_Z_M1004_d N_Z_c_1200_n
+ N_Z_c_1201_n N_Z_c_1202_n N_Z_c_1203_n N_Z_c_1208_n N_Z_c_1226_n N_Z_c_1209_n
+ N_Z_c_1257_n N_Z_c_1210_n N_Z_c_1289_n Z Z Z Z N_Z_c_1227_n N_Z_c_1204_n
+ N_Z_c_1258_n N_Z_c_1205_n N_Z_c_1290_n N_Z_c_1206_n N_Z_c_1320_n N_Z_c_1207_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%Z
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_824_333# N_A_824_333#_M1020_d
+ N_A_824_333#_M1027_d N_A_824_333#_M1023_d N_A_824_333#_c_1428_n
+ N_A_824_333#_c_1436_n N_A_824_333#_c_1438_n N_A_824_333#_c_1439_n
+ N_A_824_333#_c_1442_n N_A_824_333#_c_1440_n N_A_824_333#_c_1429_n
+ N_A_824_333#_c_1430_n N_A_824_333#_c_1431_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_824_333#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_1315_297# N_A_1315_297#_M1000_s
+ N_A_1315_297#_M1030_s N_A_1315_297#_M1031_s N_A_1315_297#_c_1487_n
+ N_A_1315_297#_c_1493_n N_A_1315_297#_c_1497_n N_A_1315_297#_c_1501_n
+ N_A_1315_297#_c_1516_n N_A_1315_297#_c_1488_n N_A_1315_297#_c_1489_n
+ N_A_1315_297#_c_1490_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_1315_297#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_2112_333# N_A_2112_333#_M1004_s
+ N_A_2112_333#_M1032_s N_A_2112_333#_M1036_s N_A_2112_333#_c_1544_n
+ N_A_2112_333#_c_1552_n N_A_2112_333#_c_1554_n N_A_2112_333#_c_1555_n
+ N_A_2112_333#_c_1558_n N_A_2112_333#_c_1556_n N_A_2112_333#_c_1545_n
+ N_A_2112_333#_c_1546_n N_A_2112_333#_c_1547_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_2112_333#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_27_47# N_A_27_47#_M1013_d
+ N_A_27_47#_M1026_d N_A_27_47#_M1014_d N_A_27_47#_c_1596_n N_A_27_47#_c_1593_n
+ N_A_27_47#_c_1594_n N_A_27_47#_c_1625_p N_A_27_47#_c_1595_n
+ N_A_27_47#_c_1606_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%VGND N_VGND_M1013_s N_VGND_M1021_d
+ N_VGND_M1019_d N_VGND_M1028_s N_VGND_M1038_d N_VGND_M1008_s N_VGND_c_1635_n
+ N_VGND_c_1636_n N_VGND_c_1637_n N_VGND_c_1638_n N_VGND_c_1639_n
+ N_VGND_c_1640_n N_VGND_c_1641_n N_VGND_c_1642_n N_VGND_c_1643_n
+ N_VGND_c_1644_n N_VGND_c_1645_n N_VGND_c_1646_n N_VGND_c_1647_n VGND VGND VGND
+ VGND N_VGND_c_1649_n N_VGND_c_1650_n N_VGND_c_1651_n N_VGND_c_1652_n
+ N_VGND_c_1653_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%VGND
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_845_69# N_A_845_69#_M1010_d
+ N_A_845_69#_M1012_d N_A_845_69#_M1024_s N_A_845_69#_c_1782_n
+ N_A_845_69#_c_1778_n N_A_845_69#_c_1779_n N_A_845_69#_c_1815_n
+ N_A_845_69#_c_1780_n N_A_845_69#_c_1781_n N_A_845_69#_c_1800_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_845_69#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_1315_47# N_A_1315_47#_M1028_d
+ N_A_1315_47#_M1033_d N_A_1315_47#_M1037_s N_A_1315_47#_c_1829_n
+ N_A_1315_47#_c_1826_n N_A_1315_47#_c_1827_n N_A_1315_47#_c_1864_n
+ N_A_1315_47#_c_1828_n N_A_1315_47#_c_1839_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_1315_47#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_2133_69# N_A_2133_69#_M1025_s
+ N_A_2133_69#_M1034_s N_A_2133_69#_M1039_d N_A_2133_69#_c_1874_n
+ N_A_2133_69#_c_1870_n N_A_2133_69#_c_1871_n N_A_2133_69#_c_1907_n
+ N_A_2133_69#_c_1872_n N_A_2133_69#_c_1873_n N_A_2133_69#_c_1892_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_2133_69#
cc_1 VNB N_D[0]_M1002_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_2 VNB N_D[0]_M1013_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_3 VNB N_D[0]_M1026_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_4 VNB N_D[0]_M1017_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_5 VNB N_D[0]_c_219_n 0.0128835f $X=-0.19 $Y=-0.24 $X2=0.75 $Y2=1.16
cc_6 VNB N_D[0]_c_220_n 0.0571683f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_7 VNB N_A_278_265#_c_262_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_8 VNB N_A_278_265#_c_263_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_278_265#_c_264_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_10 VNB N_A_278_265#_c_265_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_S[0]_c_339_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_12 VNB N_S[0]_c_340_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_S[0]_c_341_n 0.0101495f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.025
cc_14 VNB N_S[0]_c_342_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_15 VNB N_S[0]_c_343_n 0.032124f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_16 VNB N_S[0]_c_344_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_S[0]_c_345_n 0.0222544f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_18 VNB N_S[0]_c_346_n 0.0073997f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_19 VNB N_S[0]_c_347_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_20 VNB N_S[0]_c_348_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_S[0]_c_349_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_22 VNB S[0] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_S[1]_c_404_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_24 VNB N_S[1]_c_405_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_S[1]_c_406_n 0.0296541f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_26 VNB N_S[1]_c_407_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_27 VNB N_S[1]_c_408_n 0.0214653f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_28 VNB N_S[1]_c_409_n 0.0106587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_S[1]_c_410_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_30 VNB N_S[1]_c_411_n 0.0254151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_S[1]_c_412_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_S[1]_c_413_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_33 VNB S[1] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_701_47#_c_466_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_701_47#_c_467_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_701_47#_c_468_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_37 VNB N_A_701_47#_c_469_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_38 VNB N_D[1]_M1015_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_39 VNB N_D[1]_M1019_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_40 VNB N_D[1]_M1024_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_41 VNB N_D[1]_M1023_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_42 VNB D[1] 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_43 VNB N_D[1]_c_545_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_44 VNB N_D[2]_M1000_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_45 VNB N_D[2]_M1028_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_46 VNB N_D[2]_M1033_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_47 VNB N_D[2]_M1030_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_48 VNB N_D[2]_c_597_n 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.75 $Y2=1.16
cc_49 VNB N_D[2]_c_598_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_50 VNB N_A_1566_265#_c_647_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.105
cc_51 VNB N_A_1566_265#_c_648_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_1566_265#_c_649_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_53 VNB N_A_1566_265#_c_650_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_S[2]_c_725_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_55 VNB N_S[2]_c_726_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_S[2]_c_727_n 0.0101495f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.025
cc_57 VNB N_S[2]_c_728_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_58 VNB N_S[2]_c_729_n 0.032124f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_59 VNB N_S[2]_c_730_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_S[2]_c_731_n 0.0222544f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_61 VNB N_S[2]_c_732_n 0.0073997f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_62 VNB N_S[2]_c_733_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_63 VNB N_S[2]_c_734_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_S[2]_c_735_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_65 VNB S[2] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_S[3]_c_790_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_67 VNB N_S[3]_c_791_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_S[3]_c_792_n 0.0296541f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_69 VNB N_S[3]_c_793_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_70 VNB N_S[3]_c_794_n 0.0214653f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_71 VNB N_S[3]_c_795_n 0.0106587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_S[3]_c_796_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_73 VNB N_S[3]_c_797_n 0.0254151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_S[3]_c_798_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_S[3]_c_799_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_76 VNB S[3] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1989_47#_c_852_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1989_47#_c_853_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_1989_47#_c_854_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_80 VNB N_A_1989_47#_c_855_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_81 VNB N_D[3]_M1001_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_82 VNB N_D[3]_M1008_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_83 VNB N_D[3]_M1039_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_84 VNB N_D[3]_M1036_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_85 VNB D[3] 0.0128835f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_86 VNB N_D[3]_c_930_n 0.0571683f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_87 VNB VPWR 0.535415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_Z_c_1200_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.19
cc_89 VNB N_Z_c_1201_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_Z_c_1202_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_Z_c_1203_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_Z_c_1204_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_Z_c_1205_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_Z_c_1206_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_Z_c_1207_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_A_27_47#_c_1593_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_97 VNB N_A_27_47#_c_1594_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_98 VNB N_A_27_47#_c_1595_n 0.0034739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1635_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_100 VNB N_VGND_c_1636_n 0.00516508f $X=-0.19 $Y=-0.24 $X2=0.75 $Y2=1.16
cc_101 VNB N_VGND_c_1637_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_102 VNB N_VGND_c_1638_n 0.0332577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1639_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1640_n 0.00516508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1641_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1642_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1643_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1644_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1645_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1646_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1647_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB VGND 0.60715f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1649_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1650_n 0.0188039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1651_n 0.0229085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1652_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1653_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_A_845_69#_c_1778_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_119 VNB N_A_845_69#_c_1779_n 0.00109213f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_120 VNB N_A_845_69#_c_1780_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_A_845_69#_c_1781_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_122 VNB N_A_1315_47#_c_1826_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_123 VNB N_A_1315_47#_c_1827_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_124 VNB N_A_1315_47#_c_1828_n 0.0034739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_A_2133_69#_c_1870_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_126 VNB N_A_2133_69#_c_1871_n 0.00109213f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_127 VNB N_A_2133_69#_c_1872_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_A_2133_69#_c_1873_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_129 VPB N_D[0]_M1002_g 0.0296461f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_130 VPB N_D[0]_M1017_g 0.0229174f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_131 VPB N_D[0]_c_219_n 0.00632455f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_132 VPB N_A_278_265#_M1005_g 0.0234575f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_133 VPB N_A_278_265#_c_267_n 0.0152663f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_134 VPB N_A_278_265#_c_268_n 0.0114291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_278_265#_M1009_g 0.0267037f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_136 VPB N_A_278_265#_c_270_n 0.0080424f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_137 VPB N_A_278_265#_c_264_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_138 VPB N_A_278_265#_c_265_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_S[0]_c_347_n 0.0295425f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_140 VPB N_S[1]_c_405_n 0.0295425f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_701_47#_M1020_g 0.0267037f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_142 VPB N_A_701_47#_c_471_n 0.0265655f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_143 VPB N_A_701_47#_c_466_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_701_47#_M1027_g 0.0234575f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_145 VPB N_A_701_47#_c_474_n 0.0080424f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_146 VPB N_A_701_47#_c_469_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_147 VPB N_D[1]_M1015_g 0.0229174f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_148 VPB N_D[1]_M1023_g 0.0296461f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_149 VPB D[1] 0.00525107f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_150 VPB N_D[2]_M1000_g 0.0296461f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_151 VPB N_D[2]_M1030_g 0.0229174f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_152 VPB N_D[2]_c_597_n 0.00525107f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_153 VPB N_A_1566_265#_M1003_g 0.0234575f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_154 VPB N_A_1566_265#_c_652_n 0.0152663f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_155 VPB N_A_1566_265#_c_653_n 0.0112992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_1566_265#_M1031_g 0.0267037f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_157 VPB N_A_1566_265#_c_655_n 0.0080424f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_158 VPB N_A_1566_265#_c_649_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_159 VPB N_A_1566_265#_c_650_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_S[2]_c_733_n 0.0295425f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_161 VPB N_S[3]_c_791_n 0.0295425f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_1989_47#_M1004_g 0.0267037f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_163 VPB N_A_1989_47#_c_857_n 0.0266954f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_164 VPB N_A_1989_47#_c_852_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_1989_47#_M1032_g 0.0234575f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_166 VPB N_A_1989_47#_c_860_n 0.0080424f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_167 VPB N_A_1989_47#_c_855_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_168 VPB N_D[3]_M1001_g 0.0229174f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_169 VPB N_D[3]_M1036_g 0.0296461f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_170 VPB D[3] 0.00632455f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_171 VPB N_A_27_297#_c_971_n 0.0075508f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_172 VPB N_A_27_297#_c_972_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_27_297#_c_973_n 0.0101553f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_174 VPB N_A_27_297#_c_974_n 0.0207852f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_175 VPB N_VPWR_c_1019_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1020_n 0.0147403f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_177 VPB N_VPWR_c_1021_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1022_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1023_n 0.0147403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1024_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1025_n 0.0531719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1026_n 0.00631862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1027_n 0.0531719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1028_n 0.00631862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB VPWR 0.0639365f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1030_n 0.0177253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1031_n 0.0531719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_1032_n 0.0311005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_1033_n 0.0531719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1034_n 0.0177253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1035_n 0.00455763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1036_n 0.00455763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1037_n 0.00455763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1038_n 0.00455763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_Z_c_1208_n 0.0098056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_Z_c_1209_n 0.00920862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_Z_c_1210_n 0.0098056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_Z_c_1204_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_Z_c_1205_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_Z_c_1206_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_Z_c_1207_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_A_824_333#_c_1428_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_A_824_333#_c_1429_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_A_824_333#_c_1430_n 0.00256593f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_205 VPB N_A_824_333#_c_1431_n 0.00433305f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_206 VPB N_A_1315_297#_c_1487_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=0.56
cc_207 VPB N_A_1315_297#_c_1488_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_A_1315_297#_c_1489_n 0.00256593f $X=-0.19 $Y=1.305 $X2=0.75
+ $Y2=1.16
cc_209 VPB N_A_1315_297#_c_1490_n 0.00433305f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=1.16
cc_210 VPB N_A_2112_333#_c_1544_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_A_2112_333#_c_1545_n 0.0075508f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_A_2112_333#_c_1546_n 0.0101553f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_213 VPB N_A_2112_333#_c_1547_n 0.0207852f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_214 N_D[0]_M1017_g N_A_278_265#_M1005_g 0.0232231f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_215 N_D[0]_M1017_g N_A_278_265#_c_268_n 0.00671996f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_216 N_D[0]_M1026_g N_S[0]_c_341_n 0.0165585f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_217 N_D[0]_c_219_n N_A_27_297#_c_971_n 0.0235932f $X=0.75 $Y=1.16 $X2=0 $Y2=0
cc_218 N_D[0]_c_220_n N_A_27_297#_c_971_n 9.6385e-19 $X=0.965 $Y=1.16 $X2=0
+ $Y2=0
cc_219 N_D[0]_M1002_g N_A_27_297#_c_977_n 0.0142998f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_220 N_D[0]_M1017_g N_A_27_297#_c_977_n 0.0174487f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_221 N_D[0]_c_219_n N_A_27_297#_c_977_n 0.0339353f $X=0.75 $Y=1.16 $X2=0 $Y2=0
cc_222 N_D[0]_c_220_n N_A_27_297#_c_977_n 7.13708e-19 $X=0.965 $Y=1.16 $X2=0
+ $Y2=0
cc_223 N_D[0]_M1017_g N_A_27_297#_c_981_n 0.00557487f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_224 N_D[0]_M1002_g N_A_27_297#_c_973_n 0.00329008f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_225 N_D[0]_M1002_g N_VPWR_c_1019_n 0.0031734f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_226 N_D[0]_M1017_g N_VPWR_c_1019_n 0.00919666f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_227 N_D[0]_M1002_g N_VPWR_c_1041_n 0.00363183f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_228 N_D[0]_M1017_g N_VPWR_c_1041_n 0.00343746f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_229 N_D[0]_M1017_g N_VPWR_c_1025_n 0.00622633f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_230 N_D[0]_M1002_g VPWR 0.0120316f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_231 N_D[0]_M1017_g VPWR 0.0105515f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_232 N_D[0]_M1002_g N_VPWR_c_1030_n 0.00652917f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_233 N_D[0]_M1026_g N_Z_c_1204_n 8.13311e-19 $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_234 N_D[0]_M1017_g N_Z_c_1204_n 0.00112534f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_235 N_D[0]_c_219_n N_Z_c_1204_n 0.00742792f $X=0.75 $Y=1.16 $X2=0 $Y2=0
cc_236 N_D[0]_c_220_n N_Z_c_1204_n 0.00583073f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_237 N_D[0]_M1013_g N_A_27_47#_c_1596_n 0.00633603f $X=0.52 $Y=0.56 $X2=0
+ $Y2=0
cc_238 N_D[0]_M1026_g N_A_27_47#_c_1596_n 5.29024e-19 $X=0.94 $Y=0.56 $X2=0
+ $Y2=0
cc_239 N_D[0]_M1013_g N_A_27_47#_c_1593_n 0.0084485f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_240 N_D[0]_M1026_g N_A_27_47#_c_1593_n 0.0125955f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_241 N_D[0]_c_219_n N_A_27_47#_c_1593_n 0.0274027f $X=0.75 $Y=1.16 $X2=0 $Y2=0
cc_242 N_D[0]_c_220_n N_A_27_47#_c_1593_n 0.00321151f $X=0.965 $Y=1.16 $X2=0
+ $Y2=0
cc_243 N_D[0]_M1013_g N_A_27_47#_c_1594_n 8.68782e-19 $X=0.52 $Y=0.56 $X2=0
+ $Y2=0
cc_244 N_D[0]_c_219_n N_A_27_47#_c_1594_n 0.024456f $X=0.75 $Y=1.16 $X2=0 $Y2=0
cc_245 N_D[0]_c_220_n N_A_27_47#_c_1594_n 0.00464565f $X=0.965 $Y=1.16 $X2=0
+ $Y2=0
cc_246 N_D[0]_M1013_g N_VGND_c_1635_n 0.0030929f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_247 N_D[0]_M1026_g N_VGND_c_1635_n 0.00300333f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_248 N_D[0]_M1026_g N_VGND_c_1642_n 0.00436487f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_249 N_D[0]_M1013_g VGND 0.00697949f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_250 N_D[0]_M1026_g VGND 0.00600262f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_251 N_D[0]_M1013_g N_VGND_c_1651_n 0.00430643f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_252 N_A_278_265#_c_268_n N_S[0]_c_339_n 0.00779314f $X=1.58 $Y=1.4 $X2=-0.19
+ $Y2=-0.24
cc_253 N_A_278_265#_c_267_n N_S[0]_c_342_n 0.00810157f $X=1.87 $Y=1.4 $X2=0
+ $Y2=0
cc_254 N_A_278_265#_c_263_n N_S[0]_c_342_n 7.04048e-19 $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_255 N_A_278_265#_c_262_n N_S[0]_c_344_n 0.0100587f $X=2.43 $Y=0.755 $X2=0
+ $Y2=0
cc_256 N_A_278_265#_c_263_n N_S[0]_c_344_n 0.00267287f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_257 N_A_278_265#_c_262_n N_S[0]_c_345_n 0.0105766f $X=2.43 $Y=0.755 $X2=0
+ $Y2=0
cc_258 N_A_278_265#_c_263_n N_S[0]_c_345_n 0.0090765f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_259 N_A_278_265#_c_264_n N_S[0]_c_345_n 0.00742826f $X=2.715 $Y=1.63 $X2=0
+ $Y2=0
cc_260 N_A_278_265#_c_263_n N_S[0]_c_346_n 0.00445422f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_261 N_A_278_265#_c_264_n N_S[0]_c_346_n 4.25171e-19 $X=2.715 $Y=1.63 $X2=0
+ $Y2=0
cc_262 N_A_278_265#_c_265_n N_S[0]_c_346_n 0.00920672f $X=1.96 $Y=1.34 $X2=0
+ $Y2=0
cc_263 N_A_278_265#_c_263_n N_S[0]_c_347_n 0.00205356f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_264 N_A_278_265#_c_270_n N_S[0]_c_347_n 0.00862444f $X=2.715 $Y=2.31 $X2=0
+ $Y2=0
cc_265 N_A_278_265#_c_264_n N_S[0]_c_347_n 0.00828481f $X=2.715 $Y=1.63 $X2=0
+ $Y2=0
cc_266 N_A_278_265#_c_265_n N_S[0]_c_347_n 0.00692516f $X=1.96 $Y=1.34 $X2=0
+ $Y2=0
cc_267 N_A_278_265#_c_263_n N_S[0]_c_348_n 0.00149517f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_268 N_A_278_265#_c_262_n S[0] 0.0061421f $X=2.43 $Y=0.755 $X2=0 $Y2=0
cc_269 N_A_278_265#_c_263_n S[0] 0.0101733f $X=2.43 $Y=1.205 $X2=0 $Y2=0
cc_270 N_A_278_265#_c_264_n S[0] 0.0127184f $X=2.715 $Y=1.63 $X2=0 $Y2=0
cc_271 N_A_278_265#_c_265_n S[0] 3.07062e-19 $X=1.96 $Y=1.34 $X2=0 $Y2=0
cc_272 N_A_278_265#_M1005_g N_A_27_297#_c_977_n 0.00176121f $X=1.49 $Y=2.075
+ $X2=0 $Y2=0
cc_273 N_A_278_265#_M1005_g N_A_27_297#_c_981_n 0.00736707f $X=1.49 $Y=2.075
+ $X2=0 $Y2=0
cc_274 N_A_278_265#_M1005_g N_A_27_297#_c_985_n 0.0128147f $X=1.49 $Y=2.075
+ $X2=0 $Y2=0
cc_275 N_A_278_265#_M1009_g N_A_27_297#_c_985_n 0.00971609f $X=1.96 $Y=2.075
+ $X2=0 $Y2=0
cc_276 N_A_278_265#_c_270_n N_A_27_297#_c_985_n 0.010563f $X=2.715 $Y=2.31 $X2=0
+ $Y2=0
cc_277 N_A_278_265#_M1009_g N_A_27_297#_c_972_n 0.00745341f $X=1.96 $Y=2.075
+ $X2=0 $Y2=0
cc_278 N_A_278_265#_c_270_n N_A_27_297#_c_972_n 0.0347621f $X=2.715 $Y=2.31
+ $X2=0 $Y2=0
cc_279 N_A_278_265#_c_264_n N_A_27_297#_c_972_n 0.0132748f $X=2.715 $Y=1.63
+ $X2=0 $Y2=0
cc_280 N_A_278_265#_c_265_n N_A_27_297#_c_972_n 0.00133381f $X=1.96 $Y=1.34
+ $X2=0 $Y2=0
cc_281 N_A_278_265#_M1005_g N_VPWR_c_1019_n 0.00107974f $X=1.49 $Y=2.075 $X2=0
+ $Y2=0
cc_282 N_A_278_265#_c_270_n N_VPWR_c_1020_n 0.0321301f $X=2.715 $Y=2.31 $X2=0
+ $Y2=0
cc_283 N_A_278_265#_c_264_n N_VPWR_c_1020_n 0.00732952f $X=2.715 $Y=1.63 $X2=0
+ $Y2=0
cc_284 N_A_278_265#_M1005_g N_VPWR_c_1025_n 0.00429453f $X=1.49 $Y=2.075 $X2=0
+ $Y2=0
cc_285 N_A_278_265#_M1009_g N_VPWR_c_1025_n 0.00429453f $X=1.96 $Y=2.075 $X2=0
+ $Y2=0
cc_286 N_A_278_265#_c_270_n N_VPWR_c_1025_n 0.0210596f $X=2.715 $Y=2.31 $X2=0
+ $Y2=0
cc_287 N_A_278_265#_M1006_s VPWR 0.00179197f $X=2.59 $Y=1.485 $X2=0 $Y2=0
cc_288 N_A_278_265#_M1005_g VPWR 0.00617598f $X=1.49 $Y=2.075 $X2=0 $Y2=0
cc_289 N_A_278_265#_M1009_g VPWR 0.00728421f $X=1.96 $Y=2.075 $X2=0 $Y2=0
cc_290 N_A_278_265#_c_270_n VPWR 0.00594162f $X=2.715 $Y=2.31 $X2=0 $Y2=0
cc_291 N_A_278_265#_c_267_n N_Z_c_1200_n 0.00168443f $X=1.87 $Y=1.4 $X2=0 $Y2=0
cc_292 N_A_278_265#_c_268_n N_Z_c_1200_n 0.00180308f $X=1.58 $Y=1.4 $X2=0 $Y2=0
cc_293 N_A_278_265#_c_263_n N_Z_c_1200_n 0.0033343f $X=2.43 $Y=1.205 $X2=0 $Y2=0
cc_294 N_A_278_265#_M1009_g N_Z_c_1208_n 0.00753886f $X=1.96 $Y=2.075 $X2=0
+ $Y2=0
cc_295 N_A_278_265#_c_270_n N_Z_c_1208_n 0.0308332f $X=2.715 $Y=2.31 $X2=0 $Y2=0
cc_296 N_A_278_265#_c_264_n N_Z_c_1208_n 0.0132841f $X=2.715 $Y=1.63 $X2=0 $Y2=0
cc_297 N_A_278_265#_c_265_n N_Z_c_1208_n 9.57301e-19 $X=1.96 $Y=1.34 $X2=0 $Y2=0
cc_298 N_A_278_265#_M1005_g N_Z_c_1226_n 0.00635853f $X=1.49 $Y=2.075 $X2=0
+ $Y2=0
cc_299 N_A_278_265#_M1005_g N_Z_c_1227_n 0.0105371f $X=1.49 $Y=2.075 $X2=0 $Y2=0
cc_300 N_A_278_265#_c_267_n N_Z_c_1227_n 8.37785e-19 $X=1.87 $Y=1.4 $X2=0 $Y2=0
cc_301 N_A_278_265#_M1009_g N_Z_c_1227_n 0.00635536f $X=1.96 $Y=2.075 $X2=0
+ $Y2=0
cc_302 N_A_278_265#_M1005_g N_Z_c_1204_n 0.00268051f $X=1.49 $Y=2.075 $X2=0
+ $Y2=0
cc_303 N_A_278_265#_c_267_n N_Z_c_1204_n 0.0140509f $X=1.87 $Y=1.4 $X2=0 $Y2=0
cc_304 N_A_278_265#_M1009_g N_Z_c_1204_n 0.00476154f $X=1.96 $Y=2.075 $X2=0
+ $Y2=0
cc_305 N_A_278_265#_c_263_n N_Z_c_1204_n 0.00967956f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_306 N_A_278_265#_c_264_n N_Z_c_1204_n 0.0117695f $X=2.715 $Y=1.63 $X2=0 $Y2=0
cc_307 N_A_278_265#_c_265_n N_Z_c_1204_n 7.26438e-19 $X=1.96 $Y=1.34 $X2=0 $Y2=0
cc_308 N_A_278_265#_c_262_n N_A_27_47#_c_1595_n 0.00358194f $X=2.43 $Y=0.755
+ $X2=0 $Y2=0
cc_309 N_A_278_265#_c_262_n N_A_27_47#_c_1606_n 0.0185512f $X=2.43 $Y=0.755
+ $X2=0 $Y2=0
cc_310 N_A_278_265#_c_263_n N_A_27_47#_c_1606_n 0.00101918f $X=2.43 $Y=1.205
+ $X2=0 $Y2=0
cc_311 N_A_278_265#_c_264_n N_A_27_47#_c_1606_n 0.00285813f $X=2.715 $Y=1.63
+ $X2=0 $Y2=0
cc_312 N_A_278_265#_c_265_n N_A_27_47#_c_1606_n 0.00308807f $X=1.96 $Y=1.34
+ $X2=0 $Y2=0
cc_313 N_A_278_265#_c_262_n N_VGND_c_1642_n 0.0173492f $X=2.43 $Y=0.755 $X2=0
+ $Y2=0
cc_314 N_A_278_265#_M1021_s VGND 0.00250855f $X=2.675 $Y=0.235 $X2=0 $Y2=0
cc_315 N_A_278_265#_c_262_n VGND 0.0186564f $X=2.43 $Y=0.755 $X2=0 $Y2=0
cc_316 N_S[0]_c_348_n N_S[1]_c_404_n 0.0133556f $X=3.01 $Y=0.845 $X2=-0.19
+ $Y2=-0.24
cc_317 N_S[0]_c_347_n N_S[1]_c_405_n 0.0418422f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_318 S[0] N_S[1]_c_405_n 8.74983e-19 $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_319 N_S[0]_c_347_n S[1] 8.74983e-19 $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_320 S[0] S[1] 0.0208489f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_321 N_S[0]_c_347_n N_VPWR_c_1020_n 0.00456891f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_322 S[0] N_VPWR_c_1020_n 0.00569857f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_323 N_S[0]_c_347_n N_VPWR_c_1025_n 0.00673617f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_324 N_S[0]_c_347_n VPWR 0.00852379f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_325 N_S[0]_c_339_n N_Z_c_1200_n 0.00413022f $X=1.46 $Y=0.255 $X2=0 $Y2=0
cc_326 N_S[0]_c_342_n N_Z_c_1200_n 0.00495983f $X=1.88 $Y=0.255 $X2=0 $Y2=0
cc_327 N_S[0]_c_344_n N_Z_c_1200_n 4.25992e-19 $X=2.365 $Y=0.845 $X2=0 $Y2=0
cc_328 N_S[0]_c_347_n N_Z_c_1208_n 0.00513674f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_329 S[0] N_Z_c_1208_n 0.00545567f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_330 N_S[0]_c_339_n N_Z_c_1204_n 0.00199103f $X=1.46 $Y=0.255 $X2=0 $Y2=0
cc_331 N_S[0]_c_342_n N_Z_c_1204_n 0.00133607f $X=1.88 $Y=0.255 $X2=0 $Y2=0
cc_332 N_S[0]_c_339_n N_A_27_47#_c_1593_n 0.00139422f $X=1.46 $Y=0.255 $X2=0
+ $Y2=0
cc_333 N_S[0]_c_339_n N_A_27_47#_c_1595_n 0.0132844f $X=1.46 $Y=0.255 $X2=0
+ $Y2=0
cc_334 N_S[0]_c_340_n N_A_27_47#_c_1595_n 0.00211351f $X=1.805 $Y=0.18 $X2=0
+ $Y2=0
cc_335 N_S[0]_c_342_n N_A_27_47#_c_1595_n 0.0126455f $X=1.88 $Y=0.255 $X2=0
+ $Y2=0
cc_336 N_S[0]_c_343_n N_A_27_47#_c_1595_n 0.00436105f $X=2.29 $Y=0.18 $X2=0
+ $Y2=0
cc_337 N_S[0]_c_344_n N_A_27_47#_c_1595_n 0.00349455f $X=2.365 $Y=0.845 $X2=0
+ $Y2=0
cc_338 N_S[0]_c_344_n N_A_27_47#_c_1606_n 0.00295202f $X=2.365 $Y=0.845 $X2=0
+ $Y2=0
cc_339 N_S[0]_c_348_n N_VGND_c_1636_n 0.00330937f $X=3.01 $Y=0.845 $X2=0 $Y2=0
cc_340 N_S[0]_c_341_n N_VGND_c_1642_n 0.0271255f $X=1.535 $Y=0.18 $X2=0 $Y2=0
cc_341 N_S[0]_c_348_n N_VGND_c_1642_n 0.00585385f $X=3.01 $Y=0.845 $X2=0 $Y2=0
cc_342 N_S[0]_c_340_n VGND 0.00642387f $X=1.805 $Y=0.18 $X2=0 $Y2=0
cc_343 N_S[0]_c_341_n VGND 0.00474746f $X=1.535 $Y=0.18 $X2=0 $Y2=0
cc_344 N_S[0]_c_343_n VGND 0.0193094f $X=2.29 $Y=0.18 $X2=0 $Y2=0
cc_345 N_S[0]_c_348_n VGND 0.0111218f $X=3.01 $Y=0.845 $X2=0 $Y2=0
cc_346 N_S[0]_c_349_n VGND 0.00366655f $X=1.88 $Y=0.18 $X2=0 $Y2=0
cc_347 N_S[1]_c_412_n N_A_701_47#_c_471_n 0.00779314f $X=4.98 $Y=0.255 $X2=0
+ $Y2=0
cc_348 N_S[1]_c_405_n N_A_701_47#_c_466_n 0.00692516f $X=3.49 $Y=1.41 $X2=0
+ $Y2=0
cc_349 N_S[1]_c_406_n N_A_701_47#_c_466_n 0.00920672f $X=4 $Y=0.92 $X2=0 $Y2=0
cc_350 N_S[1]_c_410_n N_A_701_47#_c_466_n 0.00810157f $X=4.56 $Y=0.255 $X2=0
+ $Y2=0
cc_351 S[1] N_A_701_47#_c_466_n 3.07062e-19 $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_352 N_S[1]_c_405_n N_A_701_47#_c_474_n 0.00862444f $X=3.49 $Y=1.41 $X2=0
+ $Y2=0
cc_353 N_S[1]_c_404_n N_A_701_47#_c_467_n 0.00149517f $X=3.43 $Y=0.845 $X2=0
+ $Y2=0
cc_354 N_S[1]_c_405_n N_A_701_47#_c_467_n 0.00205356f $X=3.49 $Y=1.41 $X2=0
+ $Y2=0
cc_355 N_S[1]_c_406_n N_A_701_47#_c_467_n 0.0135307f $X=4 $Y=0.92 $X2=0 $Y2=0
cc_356 N_S[1]_c_407_n N_A_701_47#_c_467_n 0.00267287f $X=4.075 $Y=0.845 $X2=0
+ $Y2=0
cc_357 N_S[1]_c_410_n N_A_701_47#_c_467_n 7.04048e-19 $X=4.56 $Y=0.255 $X2=0
+ $Y2=0
cc_358 S[1] N_A_701_47#_c_467_n 0.0101733f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_359 N_S[1]_c_405_n N_A_701_47#_c_468_n 0.0105766f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_360 N_S[1]_c_407_n N_A_701_47#_c_468_n 0.0100587f $X=4.075 $Y=0.845 $X2=0
+ $Y2=0
cc_361 S[1] N_A_701_47#_c_468_n 0.0061421f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_362 N_S[1]_c_405_n N_A_701_47#_c_469_n 0.00828481f $X=3.49 $Y=1.41 $X2=0
+ $Y2=0
cc_363 N_S[1]_c_406_n N_A_701_47#_c_469_n 0.00785343f $X=4 $Y=0.92 $X2=0 $Y2=0
cc_364 S[1] N_A_701_47#_c_469_n 0.0127184f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_365 N_S[1]_c_411_n N_D[1]_M1019_g 0.0165585f $X=4.905 $Y=0.18 $X2=0 $Y2=0
cc_366 N_S[1]_c_405_n N_VPWR_c_1020_n 0.00456891f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_367 S[1] N_VPWR_c_1020_n 0.00569857f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_368 N_S[1]_c_405_n VPWR 0.00852379f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_369 N_S[1]_c_405_n N_VPWR_c_1031_n 0.00673617f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_370 N_S[1]_c_407_n N_Z_c_1201_n 4.25992e-19 $X=4.075 $Y=0.845 $X2=0 $Y2=0
cc_371 N_S[1]_c_410_n N_Z_c_1201_n 0.00495983f $X=4.56 $Y=0.255 $X2=0 $Y2=0
cc_372 N_S[1]_c_412_n N_Z_c_1201_n 0.00413022f $X=4.98 $Y=0.255 $X2=0 $Y2=0
cc_373 N_S[1]_c_405_n N_Z_c_1208_n 0.00513674f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_374 S[1] N_Z_c_1208_n 0.00545567f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_375 N_S[1]_c_410_n N_Z_c_1205_n 0.00133607f $X=4.56 $Y=0.255 $X2=0 $Y2=0
cc_376 N_S[1]_c_412_n N_Z_c_1205_n 0.00199103f $X=4.98 $Y=0.255 $X2=0 $Y2=0
cc_377 N_S[1]_c_404_n N_VGND_c_1636_n 0.00330937f $X=3.43 $Y=0.845 $X2=0 $Y2=0
cc_378 N_S[1]_c_404_n VGND 0.0111218f $X=3.43 $Y=0.845 $X2=0 $Y2=0
cc_379 N_S[1]_c_408_n VGND 0.0119932f $X=4.485 $Y=0.18 $X2=0 $Y2=0
cc_380 N_S[1]_c_409_n VGND 0.00731624f $X=4.15 $Y=0.18 $X2=0 $Y2=0
cc_381 N_S[1]_c_411_n VGND 0.0111713f $X=4.905 $Y=0.18 $X2=0 $Y2=0
cc_382 N_S[1]_c_413_n VGND 0.00366655f $X=4.56 $Y=0.18 $X2=0 $Y2=0
cc_383 N_S[1]_c_404_n N_VGND_c_1649_n 0.00585385f $X=3.43 $Y=0.845 $X2=0 $Y2=0
cc_384 N_S[1]_c_409_n N_VGND_c_1649_n 0.0271255f $X=4.15 $Y=0.18 $X2=0 $Y2=0
cc_385 N_S[1]_c_407_n N_A_845_69#_c_1782_n 0.00295202f $X=4.075 $Y=0.845 $X2=0
+ $Y2=0
cc_386 N_S[1]_c_410_n N_A_845_69#_c_1778_n 0.0126455f $X=4.56 $Y=0.255 $X2=0
+ $Y2=0
cc_387 N_S[1]_c_411_n N_A_845_69#_c_1778_n 0.00211351f $X=4.905 $Y=0.18 $X2=0
+ $Y2=0
cc_388 N_S[1]_c_412_n N_A_845_69#_c_1778_n 0.0132844f $X=4.98 $Y=0.255 $X2=0
+ $Y2=0
cc_389 N_S[1]_c_407_n N_A_845_69#_c_1779_n 0.00349455f $X=4.075 $Y=0.845 $X2=0
+ $Y2=0
cc_390 N_S[1]_c_408_n N_A_845_69#_c_1779_n 0.00436105f $X=4.485 $Y=0.18 $X2=0
+ $Y2=0
cc_391 N_S[1]_c_412_n N_A_845_69#_c_1781_n 0.00139422f $X=4.98 $Y=0.255 $X2=0
+ $Y2=0
cc_392 N_A_701_47#_c_471_n N_D[1]_M1015_g 0.00671996f $X=4.86 $Y=1.4 $X2=0 $Y2=0
cc_393 N_A_701_47#_M1027_g N_D[1]_M1015_g 0.0241475f $X=4.95 $Y=2.075 $X2=0
+ $Y2=0
cc_394 N_A_701_47#_c_474_n N_VPWR_c_1020_n 0.0321301f $X=3.725 $Y=2.31 $X2=0
+ $Y2=0
cc_395 N_A_701_47#_c_469_n N_VPWR_c_1020_n 0.00732952f $X=4.01 $Y=1.42 $X2=0
+ $Y2=0
cc_396 N_A_701_47#_M1027_g N_VPWR_c_1021_n 0.00107974f $X=4.95 $Y=2.075 $X2=0
+ $Y2=0
cc_397 N_A_701_47#_M1022_d VPWR 0.00179197f $X=3.58 $Y=1.485 $X2=0 $Y2=0
cc_398 N_A_701_47#_M1020_g VPWR 0.00728421f $X=4.48 $Y=2.075 $X2=0 $Y2=0
cc_399 N_A_701_47#_M1027_g VPWR 0.00615305f $X=4.95 $Y=2.075 $X2=0 $Y2=0
cc_400 N_A_701_47#_c_474_n VPWR 0.00594162f $X=3.725 $Y=2.31 $X2=0 $Y2=0
cc_401 N_A_701_47#_M1020_g N_VPWR_c_1031_n 0.00429453f $X=4.48 $Y=2.075 $X2=0
+ $Y2=0
cc_402 N_A_701_47#_M1027_g N_VPWR_c_1031_n 0.00429453f $X=4.95 $Y=2.075 $X2=0
+ $Y2=0
cc_403 N_A_701_47#_c_474_n N_VPWR_c_1031_n 0.0210596f $X=3.725 $Y=2.31 $X2=0
+ $Y2=0
cc_404 N_A_701_47#_c_471_n N_Z_c_1201_n 0.00348752f $X=4.86 $Y=1.4 $X2=0 $Y2=0
cc_405 N_A_701_47#_c_467_n N_Z_c_1201_n 0.0033343f $X=4.01 $Y=1.205 $X2=0 $Y2=0
cc_406 N_A_701_47#_M1020_g N_Z_c_1208_n 0.00753886f $X=4.48 $Y=2.075 $X2=0 $Y2=0
cc_407 N_A_701_47#_c_466_n N_Z_c_1208_n 9.57301e-19 $X=4.57 $Y=1.4 $X2=0 $Y2=0
cc_408 N_A_701_47#_c_474_n N_Z_c_1208_n 0.0308332f $X=3.725 $Y=2.31 $X2=0 $Y2=0
cc_409 N_A_701_47#_c_469_n N_Z_c_1208_n 0.0132841f $X=4.01 $Y=1.42 $X2=0 $Y2=0
cc_410 N_A_701_47#_M1027_g N_Z_c_1209_n 0.00411531f $X=4.95 $Y=2.075 $X2=0 $Y2=0
cc_411 N_A_701_47#_M1027_g N_Z_c_1257_n 0.00513826f $X=4.95 $Y=2.075 $X2=0 $Y2=0
cc_412 N_A_701_47#_M1020_g N_Z_c_1258_n 0.00635536f $X=4.48 $Y=2.075 $X2=0 $Y2=0
cc_413 N_A_701_47#_c_471_n N_Z_c_1258_n 8.37785e-19 $X=4.86 $Y=1.4 $X2=0 $Y2=0
cc_414 N_A_701_47#_M1027_g N_Z_c_1258_n 0.0105371f $X=4.95 $Y=2.075 $X2=0 $Y2=0
cc_415 N_A_701_47#_M1020_g N_Z_c_1205_n 0.00476154f $X=4.48 $Y=2.075 $X2=0 $Y2=0
cc_416 N_A_701_47#_c_471_n N_Z_c_1205_n 0.0140509f $X=4.86 $Y=1.4 $X2=0 $Y2=0
cc_417 N_A_701_47#_c_466_n N_Z_c_1205_n 7.26438e-19 $X=4.57 $Y=1.4 $X2=0 $Y2=0
cc_418 N_A_701_47#_M1027_g N_Z_c_1205_n 0.00268051f $X=4.95 $Y=2.075 $X2=0 $Y2=0
cc_419 N_A_701_47#_c_467_n N_Z_c_1205_n 0.00967956f $X=4.01 $Y=1.205 $X2=0 $Y2=0
cc_420 N_A_701_47#_c_469_n N_Z_c_1205_n 0.0117695f $X=4.01 $Y=1.42 $X2=0 $Y2=0
cc_421 N_A_701_47#_M1020_g N_A_824_333#_c_1428_n 0.00745341f $X=4.48 $Y=2.075
+ $X2=0 $Y2=0
cc_422 N_A_701_47#_c_466_n N_A_824_333#_c_1428_n 0.00133381f $X=4.57 $Y=1.4
+ $X2=0 $Y2=0
cc_423 N_A_701_47#_c_474_n N_A_824_333#_c_1428_n 0.0347621f $X=3.725 $Y=2.31
+ $X2=0 $Y2=0
cc_424 N_A_701_47#_c_469_n N_A_824_333#_c_1428_n 0.0132748f $X=4.01 $Y=1.42
+ $X2=0 $Y2=0
cc_425 N_A_701_47#_M1020_g N_A_824_333#_c_1436_n 0.00971609f $X=4.48 $Y=2.075
+ $X2=0 $Y2=0
cc_426 N_A_701_47#_M1027_g N_A_824_333#_c_1436_n 0.0111338f $X=4.95 $Y=2.075
+ $X2=0 $Y2=0
cc_427 N_A_701_47#_c_474_n N_A_824_333#_c_1438_n 0.010563f $X=3.725 $Y=2.31
+ $X2=0 $Y2=0
cc_428 N_A_701_47#_M1027_g N_A_824_333#_c_1439_n 0.00717732f $X=4.95 $Y=2.075
+ $X2=0 $Y2=0
cc_429 N_A_701_47#_M1027_g N_A_824_333#_c_1440_n 0.00176121f $X=4.95 $Y=2.075
+ $X2=0 $Y2=0
cc_430 N_A_701_47#_M1018_d VGND 0.00250855f $X=3.505 $Y=0.235 $X2=0 $Y2=0
cc_431 N_A_701_47#_c_468_n VGND 0.0186564f $X=3.64 $Y=0.495 $X2=0 $Y2=0
cc_432 N_A_701_47#_c_468_n N_VGND_c_1649_n 0.0173492f $X=3.64 $Y=0.495 $X2=0
+ $Y2=0
cc_433 N_A_701_47#_c_466_n N_A_845_69#_c_1782_n 0.00308807f $X=4.57 $Y=1.4 $X2=0
+ $Y2=0
cc_434 N_A_701_47#_c_467_n N_A_845_69#_c_1782_n 0.00101918f $X=4.01 $Y=1.205
+ $X2=0 $Y2=0
cc_435 N_A_701_47#_c_468_n N_A_845_69#_c_1782_n 0.0185512f $X=3.64 $Y=0.495
+ $X2=0 $Y2=0
cc_436 N_A_701_47#_c_469_n N_A_845_69#_c_1782_n 0.00285813f $X=4.01 $Y=1.42
+ $X2=0 $Y2=0
cc_437 N_A_701_47#_c_468_n N_A_845_69#_c_1779_n 0.00358194f $X=3.64 $Y=0.495
+ $X2=0 $Y2=0
cc_438 D[1] N_D[2]_c_597_n 0.0231965f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_439 N_D[1]_c_545_n N_D[2]_c_597_n 7.85936e-19 $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_440 D[1] N_D[2]_c_598_n 7.85936e-19 $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_441 N_D[1]_c_545_n N_D[2]_c_598_n 0.00603597f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_442 N_D[1]_M1015_g N_VPWR_c_1021_n 0.00919666f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_443 N_D[1]_M1023_g N_VPWR_c_1021_n 0.0031734f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_444 N_D[1]_M1015_g N_VPWR_c_1077_n 0.00295119f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_445 N_D[1]_M1023_g N_VPWR_c_1077_n 0.00314707f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_446 N_D[1]_M1015_g VPWR 0.00588601f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_447 N_D[1]_M1023_g VPWR 0.00822554f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_448 N_D[1]_M1015_g N_VPWR_c_1031_n 0.00622633f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_449 N_D[1]_M1023_g N_VPWR_c_1032_n 0.00652917f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_450 N_D[1]_M1015_g N_Z_c_1209_n 0.00431834f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_451 N_D[1]_M1023_g N_Z_c_1209_n 0.00406261f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_452 D[1] N_Z_c_1209_n 0.00125914f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_453 N_D[1]_M1015_g N_Z_c_1205_n 0.00112534f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_454 N_D[1]_M1019_g N_Z_c_1205_n 8.13311e-19 $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_455 D[1] N_Z_c_1205_n 0.00742792f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_456 N_D[1]_c_545_n N_Z_c_1205_n 0.00583073f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_457 N_D[1]_M1015_g N_A_824_333#_c_1439_n 0.00541465f $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_458 N_D[1]_M1015_g N_A_824_333#_c_1442_n 0.0127833f $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_459 N_D[1]_M1023_g N_A_824_333#_c_1442_n 0.0101085f $X=5.945 $Y=1.985 $X2=0
+ $Y2=0
cc_460 D[1] N_A_824_333#_c_1442_n 0.0323774f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_461 N_D[1]_c_545_n N_A_824_333#_c_1442_n 7.13708e-19 $X=6.03 $Y=1.16 $X2=0
+ $Y2=0
cc_462 D[1] N_A_824_333#_c_1429_n 0.0226682f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_463 N_D[1]_c_545_n N_A_824_333#_c_1429_n 9.6385e-19 $X=6.03 $Y=1.16 $X2=0
+ $Y2=0
cc_464 N_D[1]_M1023_g N_A_824_333#_c_1430_n 0.00325722f $X=5.945 $Y=1.985 $X2=0
+ $Y2=0
cc_465 N_D[1]_M1019_g N_VGND_c_1637_n 0.00300333f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_466 N_D[1]_M1024_g N_VGND_c_1637_n 0.0030929f $X=5.92 $Y=0.56 $X2=0 $Y2=0
cc_467 N_D[1]_M1024_g N_VGND_c_1638_n 0.00430643f $X=5.92 $Y=0.56 $X2=0 $Y2=0
cc_468 N_D[1]_M1019_g VGND 0.00600262f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_469 N_D[1]_M1024_g VGND 0.00733187f $X=5.92 $Y=0.56 $X2=0 $Y2=0
cc_470 N_D[1]_M1019_g N_VGND_c_1649_n 0.00436487f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_471 N_D[1]_M1019_g N_A_845_69#_c_1780_n 0.0114493f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_472 N_D[1]_M1024_g N_A_845_69#_c_1780_n 0.00931728f $X=5.92 $Y=0.56 $X2=0
+ $Y2=0
cc_473 D[1] N_A_845_69#_c_1780_n 0.0518587f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_474 N_D[1]_c_545_n N_A_845_69#_c_1780_n 0.00665175f $X=6.03 $Y=1.16 $X2=0
+ $Y2=0
cc_475 N_D[1]_M1019_g N_A_845_69#_c_1781_n 0.00114614f $X=5.5 $Y=0.56 $X2=0
+ $Y2=0
cc_476 N_D[1]_c_545_n N_A_845_69#_c_1781_n 0.00120541f $X=6.03 $Y=1.16 $X2=0
+ $Y2=0
cc_477 N_D[1]_M1019_g N_A_845_69#_c_1800_n 5.29024e-19 $X=5.5 $Y=0.56 $X2=0
+ $Y2=0
cc_478 N_D[1]_M1024_g N_A_845_69#_c_1800_n 0.00633603f $X=5.92 $Y=0.56 $X2=0
+ $Y2=0
cc_479 N_D[2]_M1030_g N_A_1566_265#_M1003_g 0.0241475f $X=7.405 $Y=1.985 $X2=0
+ $Y2=0
cc_480 N_D[2]_M1030_g N_A_1566_265#_c_653_n 0.00671996f $X=7.405 $Y=1.985 $X2=0
+ $Y2=0
cc_481 N_D[2]_M1033_g N_S[2]_c_727_n 0.0165585f $X=7.38 $Y=0.56 $X2=0 $Y2=0
cc_482 N_D[2]_M1000_g N_VPWR_c_1022_n 0.0031734f $X=6.935 $Y=1.985 $X2=0 $Y2=0
cc_483 N_D[2]_M1030_g N_VPWR_c_1022_n 0.00919666f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_484 N_D[2]_M1000_g N_VPWR_c_1085_n 0.00314707f $X=6.935 $Y=1.985 $X2=0 $Y2=0
cc_485 N_D[2]_M1030_g N_VPWR_c_1085_n 0.00295119f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_486 N_D[2]_M1030_g N_VPWR_c_1027_n 0.00622633f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_487 N_D[2]_M1000_g VPWR 0.00822554f $X=6.935 $Y=1.985 $X2=0 $Y2=0
cc_488 N_D[2]_M1030_g VPWR 0.00588601f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_489 N_D[2]_M1000_g N_VPWR_c_1032_n 0.00652917f $X=6.935 $Y=1.985 $X2=0 $Y2=0
cc_490 N_D[2]_M1000_g N_Z_c_1209_n 0.00406261f $X=6.935 $Y=1.985 $X2=0 $Y2=0
cc_491 N_D[2]_M1030_g N_Z_c_1209_n 0.00431834f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_492 N_D[2]_c_597_n N_Z_c_1209_n 0.00125914f $X=7.19 $Y=1.16 $X2=0 $Y2=0
cc_493 N_D[2]_M1033_g N_Z_c_1206_n 8.13311e-19 $X=7.38 $Y=0.56 $X2=0 $Y2=0
cc_494 N_D[2]_M1030_g N_Z_c_1206_n 0.00112534f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_495 N_D[2]_c_597_n N_Z_c_1206_n 0.00742792f $X=7.19 $Y=1.16 $X2=0 $Y2=0
cc_496 N_D[2]_c_598_n N_Z_c_1206_n 0.00583073f $X=7.405 $Y=1.16 $X2=0 $Y2=0
cc_497 N_D[2]_c_597_n N_A_1315_297#_c_1487_n 0.0226682f $X=7.19 $Y=1.16 $X2=0
+ $Y2=0
cc_498 N_D[2]_c_598_n N_A_1315_297#_c_1487_n 9.6385e-19 $X=7.405 $Y=1.16 $X2=0
+ $Y2=0
cc_499 N_D[2]_M1000_g N_A_1315_297#_c_1493_n 0.0101085f $X=6.935 $Y=1.985 $X2=0
+ $Y2=0
cc_500 N_D[2]_M1030_g N_A_1315_297#_c_1493_n 0.0127833f $X=7.405 $Y=1.985 $X2=0
+ $Y2=0
cc_501 N_D[2]_c_597_n N_A_1315_297#_c_1493_n 0.0323774f $X=7.19 $Y=1.16 $X2=0
+ $Y2=0
cc_502 N_D[2]_c_598_n N_A_1315_297#_c_1493_n 7.13708e-19 $X=7.405 $Y=1.16 $X2=0
+ $Y2=0
cc_503 N_D[2]_M1030_g N_A_1315_297#_c_1497_n 0.00541465f $X=7.405 $Y=1.985 $X2=0
+ $Y2=0
cc_504 N_D[2]_M1000_g N_A_1315_297#_c_1489_n 0.00325722f $X=6.935 $Y=1.985 $X2=0
+ $Y2=0
cc_505 N_D[2]_M1028_g N_VGND_c_1638_n 0.00430643f $X=6.96 $Y=0.56 $X2=0 $Y2=0
cc_506 N_D[2]_M1028_g N_VGND_c_1639_n 0.0030929f $X=6.96 $Y=0.56 $X2=0 $Y2=0
cc_507 N_D[2]_M1033_g N_VGND_c_1639_n 0.00300333f $X=7.38 $Y=0.56 $X2=0 $Y2=0
cc_508 N_D[2]_M1033_g N_VGND_c_1644_n 0.00436487f $X=7.38 $Y=0.56 $X2=0 $Y2=0
cc_509 N_D[2]_M1028_g VGND 0.00733187f $X=6.96 $Y=0.56 $X2=0 $Y2=0
cc_510 N_D[2]_M1033_g VGND 0.00600262f $X=7.38 $Y=0.56 $X2=0 $Y2=0
cc_511 N_D[2]_M1028_g N_A_1315_47#_c_1829_n 0.00633603f $X=6.96 $Y=0.56 $X2=0
+ $Y2=0
cc_512 N_D[2]_M1033_g N_A_1315_47#_c_1829_n 5.29024e-19 $X=7.38 $Y=0.56 $X2=0
+ $Y2=0
cc_513 N_D[2]_M1028_g N_A_1315_47#_c_1826_n 0.0084485f $X=6.96 $Y=0.56 $X2=0
+ $Y2=0
cc_514 N_D[2]_M1033_g N_A_1315_47#_c_1826_n 0.0125955f $X=7.38 $Y=0.56 $X2=0
+ $Y2=0
cc_515 N_D[2]_c_597_n N_A_1315_47#_c_1826_n 0.0274027f $X=7.19 $Y=1.16 $X2=0
+ $Y2=0
cc_516 N_D[2]_c_598_n N_A_1315_47#_c_1826_n 0.00321151f $X=7.405 $Y=1.16 $X2=0
+ $Y2=0
cc_517 N_D[2]_M1028_g N_A_1315_47#_c_1827_n 8.68782e-19 $X=6.96 $Y=0.56 $X2=0
+ $Y2=0
cc_518 N_D[2]_c_597_n N_A_1315_47#_c_1827_n 0.024456f $X=7.19 $Y=1.16 $X2=0
+ $Y2=0
cc_519 N_D[2]_c_598_n N_A_1315_47#_c_1827_n 0.00464565f $X=7.405 $Y=1.16 $X2=0
+ $Y2=0
cc_520 N_A_1566_265#_c_653_n N_S[2]_c_725_n 0.00779314f $X=8.02 $Y=1.4 $X2=-0.19
+ $Y2=-0.24
cc_521 N_A_1566_265#_c_652_n N_S[2]_c_728_n 0.00810157f $X=8.31 $Y=1.4 $X2=0
+ $Y2=0
cc_522 N_A_1566_265#_c_648_n N_S[2]_c_728_n 7.04048e-19 $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_523 N_A_1566_265#_c_647_n N_S[2]_c_730_n 0.0100587f $X=8.87 $Y=0.755 $X2=0
+ $Y2=0
cc_524 N_A_1566_265#_c_648_n N_S[2]_c_730_n 0.00267287f $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_525 N_A_1566_265#_c_647_n N_S[2]_c_731_n 0.0105766f $X=8.87 $Y=0.755 $X2=0
+ $Y2=0
cc_526 N_A_1566_265#_c_648_n N_S[2]_c_731_n 0.0090765f $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_527 N_A_1566_265#_c_649_n N_S[2]_c_731_n 0.00742826f $X=9.155 $Y=1.63 $X2=0
+ $Y2=0
cc_528 N_A_1566_265#_c_648_n N_S[2]_c_732_n 0.00445422f $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_529 N_A_1566_265#_c_649_n N_S[2]_c_732_n 4.25171e-19 $X=9.155 $Y=1.63 $X2=0
+ $Y2=0
cc_530 N_A_1566_265#_c_650_n N_S[2]_c_732_n 0.00920672f $X=8.4 $Y=1.34 $X2=0
+ $Y2=0
cc_531 N_A_1566_265#_c_648_n N_S[2]_c_733_n 0.00205356f $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_532 N_A_1566_265#_c_655_n N_S[2]_c_733_n 0.00862444f $X=9.155 $Y=2.31 $X2=0
+ $Y2=0
cc_533 N_A_1566_265#_c_649_n N_S[2]_c_733_n 0.00828481f $X=9.155 $Y=1.63 $X2=0
+ $Y2=0
cc_534 N_A_1566_265#_c_650_n N_S[2]_c_733_n 0.00692516f $X=8.4 $Y=1.34 $X2=0
+ $Y2=0
cc_535 N_A_1566_265#_c_648_n N_S[2]_c_734_n 0.00149517f $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_536 N_A_1566_265#_c_647_n S[2] 0.0061421f $X=8.87 $Y=0.755 $X2=0 $Y2=0
cc_537 N_A_1566_265#_c_648_n S[2] 0.0101733f $X=8.87 $Y=1.205 $X2=0 $Y2=0
cc_538 N_A_1566_265#_c_649_n S[2] 0.0127184f $X=9.155 $Y=1.63 $X2=0 $Y2=0
cc_539 N_A_1566_265#_c_650_n S[2] 3.07062e-19 $X=8.4 $Y=1.34 $X2=0 $Y2=0
cc_540 N_A_1566_265#_M1003_g N_VPWR_c_1022_n 0.00107974f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_541 N_A_1566_265#_c_655_n N_VPWR_c_1023_n 0.0321301f $X=9.155 $Y=2.31 $X2=0
+ $Y2=0
cc_542 N_A_1566_265#_c_649_n N_VPWR_c_1023_n 0.00732952f $X=9.155 $Y=1.63 $X2=0
+ $Y2=0
cc_543 N_A_1566_265#_M1003_g N_VPWR_c_1027_n 0.00429453f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_544 N_A_1566_265#_M1031_g N_VPWR_c_1027_n 0.00429453f $X=8.4 $Y=2.075 $X2=0
+ $Y2=0
cc_545 N_A_1566_265#_c_655_n N_VPWR_c_1027_n 0.0210596f $X=9.155 $Y=2.31 $X2=0
+ $Y2=0
cc_546 N_A_1566_265#_M1035_s VPWR 0.00179197f $X=9.03 $Y=1.485 $X2=0 $Y2=0
cc_547 N_A_1566_265#_M1003_g VPWR 0.00615305f $X=7.93 $Y=2.075 $X2=0 $Y2=0
cc_548 N_A_1566_265#_M1031_g VPWR 0.00728421f $X=8.4 $Y=2.075 $X2=0 $Y2=0
cc_549 N_A_1566_265#_c_655_n VPWR 0.00594162f $X=9.155 $Y=2.31 $X2=0 $Y2=0
cc_550 N_A_1566_265#_c_652_n N_Z_c_1202_n 0.00168443f $X=8.31 $Y=1.4 $X2=0 $Y2=0
cc_551 N_A_1566_265#_c_653_n N_Z_c_1202_n 0.00180308f $X=8.02 $Y=1.4 $X2=0 $Y2=0
cc_552 N_A_1566_265#_c_648_n N_Z_c_1202_n 0.0033343f $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_553 N_A_1566_265#_M1003_g N_Z_c_1209_n 0.00411531f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_554 N_A_1566_265#_M1031_g N_Z_c_1210_n 0.00753886f $X=8.4 $Y=2.075 $X2=0
+ $Y2=0
cc_555 N_A_1566_265#_c_655_n N_Z_c_1210_n 0.0308332f $X=9.155 $Y=2.31 $X2=0
+ $Y2=0
cc_556 N_A_1566_265#_c_649_n N_Z_c_1210_n 0.0132841f $X=9.155 $Y=1.63 $X2=0
+ $Y2=0
cc_557 N_A_1566_265#_c_650_n N_Z_c_1210_n 9.57301e-19 $X=8.4 $Y=1.34 $X2=0 $Y2=0
cc_558 N_A_1566_265#_M1003_g N_Z_c_1289_n 0.00513826f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_559 N_A_1566_265#_M1003_g N_Z_c_1290_n 0.0105371f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_560 N_A_1566_265#_c_652_n N_Z_c_1290_n 8.37785e-19 $X=8.31 $Y=1.4 $X2=0 $Y2=0
cc_561 N_A_1566_265#_M1031_g N_Z_c_1290_n 0.00635536f $X=8.4 $Y=2.075 $X2=0
+ $Y2=0
cc_562 N_A_1566_265#_M1003_g N_Z_c_1206_n 0.00268051f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_563 N_A_1566_265#_c_652_n N_Z_c_1206_n 0.0140509f $X=8.31 $Y=1.4 $X2=0 $Y2=0
cc_564 N_A_1566_265#_M1031_g N_Z_c_1206_n 0.00476154f $X=8.4 $Y=2.075 $X2=0
+ $Y2=0
cc_565 N_A_1566_265#_c_648_n N_Z_c_1206_n 0.00967956f $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_566 N_A_1566_265#_c_649_n N_Z_c_1206_n 0.0117695f $X=9.155 $Y=1.63 $X2=0
+ $Y2=0
cc_567 N_A_1566_265#_c_650_n N_Z_c_1206_n 7.26438e-19 $X=8.4 $Y=1.34 $X2=0 $Y2=0
cc_568 N_A_1566_265#_M1003_g N_A_1315_297#_c_1493_n 0.00176121f $X=7.93 $Y=2.075
+ $X2=0 $Y2=0
cc_569 N_A_1566_265#_M1003_g N_A_1315_297#_c_1497_n 0.00717732f $X=7.93 $Y=2.075
+ $X2=0 $Y2=0
cc_570 N_A_1566_265#_M1003_g N_A_1315_297#_c_1501_n 0.0111338f $X=7.93 $Y=2.075
+ $X2=0 $Y2=0
cc_571 N_A_1566_265#_M1031_g N_A_1315_297#_c_1501_n 0.00971609f $X=8.4 $Y=2.075
+ $X2=0 $Y2=0
cc_572 N_A_1566_265#_c_655_n N_A_1315_297#_c_1501_n 0.010563f $X=9.155 $Y=2.31
+ $X2=0 $Y2=0
cc_573 N_A_1566_265#_M1031_g N_A_1315_297#_c_1488_n 0.00745341f $X=8.4 $Y=2.075
+ $X2=0 $Y2=0
cc_574 N_A_1566_265#_c_655_n N_A_1315_297#_c_1488_n 0.0347621f $X=9.155 $Y=2.31
+ $X2=0 $Y2=0
cc_575 N_A_1566_265#_c_649_n N_A_1315_297#_c_1488_n 0.0132748f $X=9.155 $Y=1.63
+ $X2=0 $Y2=0
cc_576 N_A_1566_265#_c_650_n N_A_1315_297#_c_1488_n 0.00133381f $X=8.4 $Y=1.34
+ $X2=0 $Y2=0
cc_577 N_A_1566_265#_c_647_n N_VGND_c_1644_n 0.0173492f $X=8.87 $Y=0.755 $X2=0
+ $Y2=0
cc_578 N_A_1566_265#_M1038_s VGND 0.00250855f $X=9.115 $Y=0.235 $X2=0 $Y2=0
cc_579 N_A_1566_265#_c_647_n VGND 0.0186564f $X=8.87 $Y=0.755 $X2=0 $Y2=0
cc_580 N_A_1566_265#_c_647_n N_A_1315_47#_c_1828_n 0.00358194f $X=8.87 $Y=0.755
+ $X2=0 $Y2=0
cc_581 N_A_1566_265#_c_647_n N_A_1315_47#_c_1839_n 0.0185512f $X=8.87 $Y=0.755
+ $X2=0 $Y2=0
cc_582 N_A_1566_265#_c_648_n N_A_1315_47#_c_1839_n 0.00101918f $X=8.87 $Y=1.205
+ $X2=0 $Y2=0
cc_583 N_A_1566_265#_c_649_n N_A_1315_47#_c_1839_n 0.00285813f $X=9.155 $Y=1.63
+ $X2=0 $Y2=0
cc_584 N_A_1566_265#_c_650_n N_A_1315_47#_c_1839_n 0.00308807f $X=8.4 $Y=1.34
+ $X2=0 $Y2=0
cc_585 N_S[2]_c_734_n N_S[3]_c_790_n 0.0133556f $X=9.45 $Y=0.845 $X2=-0.19
+ $Y2=-0.24
cc_586 N_S[2]_c_733_n N_S[3]_c_791_n 0.0418422f $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_587 S[2] N_S[3]_c_791_n 8.74983e-19 $X=9.345 $Y=1.105 $X2=0 $Y2=0
cc_588 N_S[2]_c_733_n S[3] 8.74983e-19 $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_589 S[2] S[3] 0.0208489f $X=9.345 $Y=1.105 $X2=0 $Y2=0
cc_590 N_S[2]_c_733_n N_VPWR_c_1023_n 0.00456891f $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_591 S[2] N_VPWR_c_1023_n 0.00569857f $X=9.345 $Y=1.105 $X2=0 $Y2=0
cc_592 N_S[2]_c_733_n N_VPWR_c_1027_n 0.00673617f $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_593 N_S[2]_c_733_n VPWR 0.00852379f $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_594 N_S[2]_c_725_n N_Z_c_1202_n 0.00413022f $X=7.9 $Y=0.255 $X2=0 $Y2=0
cc_595 N_S[2]_c_728_n N_Z_c_1202_n 0.00495983f $X=8.32 $Y=0.255 $X2=0 $Y2=0
cc_596 N_S[2]_c_730_n N_Z_c_1202_n 4.25992e-19 $X=8.805 $Y=0.845 $X2=0 $Y2=0
cc_597 N_S[2]_c_733_n N_Z_c_1210_n 0.00513674f $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_598 S[2] N_Z_c_1210_n 0.00545567f $X=9.345 $Y=1.105 $X2=0 $Y2=0
cc_599 N_S[2]_c_725_n N_Z_c_1206_n 0.00199103f $X=7.9 $Y=0.255 $X2=0 $Y2=0
cc_600 N_S[2]_c_728_n N_Z_c_1206_n 0.00133607f $X=8.32 $Y=0.255 $X2=0 $Y2=0
cc_601 N_S[2]_c_734_n N_VGND_c_1640_n 0.00330937f $X=9.45 $Y=0.845 $X2=0 $Y2=0
cc_602 N_S[2]_c_727_n N_VGND_c_1644_n 0.0271255f $X=7.975 $Y=0.18 $X2=0 $Y2=0
cc_603 N_S[2]_c_734_n N_VGND_c_1644_n 0.00585385f $X=9.45 $Y=0.845 $X2=0 $Y2=0
cc_604 N_S[2]_c_726_n VGND 0.00642387f $X=8.245 $Y=0.18 $X2=0 $Y2=0
cc_605 N_S[2]_c_727_n VGND 0.00474746f $X=7.975 $Y=0.18 $X2=0 $Y2=0
cc_606 N_S[2]_c_729_n VGND 0.0193094f $X=8.73 $Y=0.18 $X2=0 $Y2=0
cc_607 N_S[2]_c_734_n VGND 0.0111218f $X=9.45 $Y=0.845 $X2=0 $Y2=0
cc_608 N_S[2]_c_735_n VGND 0.00366655f $X=8.32 $Y=0.18 $X2=0 $Y2=0
cc_609 N_S[2]_c_725_n N_A_1315_47#_c_1826_n 0.00139422f $X=7.9 $Y=0.255 $X2=0
+ $Y2=0
cc_610 N_S[2]_c_725_n N_A_1315_47#_c_1828_n 0.0132844f $X=7.9 $Y=0.255 $X2=0
+ $Y2=0
cc_611 N_S[2]_c_726_n N_A_1315_47#_c_1828_n 0.00211351f $X=8.245 $Y=0.18 $X2=0
+ $Y2=0
cc_612 N_S[2]_c_728_n N_A_1315_47#_c_1828_n 0.0126455f $X=8.32 $Y=0.255 $X2=0
+ $Y2=0
cc_613 N_S[2]_c_729_n N_A_1315_47#_c_1828_n 0.00436105f $X=8.73 $Y=0.18 $X2=0
+ $Y2=0
cc_614 N_S[2]_c_730_n N_A_1315_47#_c_1828_n 0.00349455f $X=8.805 $Y=0.845 $X2=0
+ $Y2=0
cc_615 N_S[2]_c_730_n N_A_1315_47#_c_1839_n 0.00295202f $X=8.805 $Y=0.845 $X2=0
+ $Y2=0
cc_616 N_S[3]_c_798_n N_A_1989_47#_c_857_n 0.00779314f $X=11.42 $Y=0.255 $X2=0
+ $Y2=0
cc_617 N_S[3]_c_791_n N_A_1989_47#_c_852_n 0.00692516f $X=9.93 $Y=1.41 $X2=0
+ $Y2=0
cc_618 N_S[3]_c_792_n N_A_1989_47#_c_852_n 0.00920672f $X=10.44 $Y=0.92 $X2=0
+ $Y2=0
cc_619 N_S[3]_c_796_n N_A_1989_47#_c_852_n 0.00810157f $X=11 $Y=0.255 $X2=0
+ $Y2=0
cc_620 S[3] N_A_1989_47#_c_852_n 3.07062e-19 $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_621 N_S[3]_c_791_n N_A_1989_47#_c_860_n 0.00862444f $X=9.93 $Y=1.41 $X2=0
+ $Y2=0
cc_622 N_S[3]_c_790_n N_A_1989_47#_c_853_n 0.00149517f $X=9.87 $Y=0.845 $X2=0
+ $Y2=0
cc_623 N_S[3]_c_791_n N_A_1989_47#_c_853_n 0.00205356f $X=9.93 $Y=1.41 $X2=0
+ $Y2=0
cc_624 N_S[3]_c_792_n N_A_1989_47#_c_853_n 0.0135307f $X=10.44 $Y=0.92 $X2=0
+ $Y2=0
cc_625 N_S[3]_c_793_n N_A_1989_47#_c_853_n 0.00267287f $X=10.515 $Y=0.845 $X2=0
+ $Y2=0
cc_626 N_S[3]_c_796_n N_A_1989_47#_c_853_n 7.04048e-19 $X=11 $Y=0.255 $X2=0
+ $Y2=0
cc_627 S[3] N_A_1989_47#_c_853_n 0.0101733f $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_628 N_S[3]_c_791_n N_A_1989_47#_c_854_n 0.0105766f $X=9.93 $Y=1.41 $X2=0
+ $Y2=0
cc_629 N_S[3]_c_793_n N_A_1989_47#_c_854_n 0.0100587f $X=10.515 $Y=0.845 $X2=0
+ $Y2=0
cc_630 S[3] N_A_1989_47#_c_854_n 0.0061421f $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_631 N_S[3]_c_791_n N_A_1989_47#_c_855_n 0.00828481f $X=9.93 $Y=1.41 $X2=0
+ $Y2=0
cc_632 N_S[3]_c_792_n N_A_1989_47#_c_855_n 0.00785343f $X=10.44 $Y=0.92 $X2=0
+ $Y2=0
cc_633 S[3] N_A_1989_47#_c_855_n 0.0127184f $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_634 N_S[3]_c_797_n N_D[3]_M1008_g 0.0165585f $X=11.345 $Y=0.18 $X2=0 $Y2=0
cc_635 N_S[3]_c_791_n N_VPWR_c_1023_n 0.00456891f $X=9.93 $Y=1.41 $X2=0 $Y2=0
cc_636 S[3] N_VPWR_c_1023_n 0.00569857f $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_637 N_S[3]_c_791_n VPWR 0.00852379f $X=9.93 $Y=1.41 $X2=0 $Y2=0
cc_638 N_S[3]_c_791_n N_VPWR_c_1033_n 0.00673617f $X=9.93 $Y=1.41 $X2=0 $Y2=0
cc_639 N_S[3]_c_793_n N_Z_c_1203_n 4.25992e-19 $X=10.515 $Y=0.845 $X2=0 $Y2=0
cc_640 N_S[3]_c_796_n N_Z_c_1203_n 0.00495983f $X=11 $Y=0.255 $X2=0 $Y2=0
cc_641 N_S[3]_c_798_n N_Z_c_1203_n 0.00413022f $X=11.42 $Y=0.255 $X2=0 $Y2=0
cc_642 N_S[3]_c_791_n N_Z_c_1210_n 0.00513674f $X=9.93 $Y=1.41 $X2=0 $Y2=0
cc_643 S[3] N_Z_c_1210_n 0.00545567f $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_644 N_S[3]_c_796_n N_Z_c_1207_n 0.00133607f $X=11 $Y=0.255 $X2=0 $Y2=0
cc_645 N_S[3]_c_798_n N_Z_c_1207_n 0.00199103f $X=11.42 $Y=0.255 $X2=0 $Y2=0
cc_646 N_S[3]_c_790_n N_VGND_c_1640_n 0.00330937f $X=9.87 $Y=0.845 $X2=0 $Y2=0
cc_647 N_S[3]_c_790_n N_VGND_c_1646_n 0.00585385f $X=9.87 $Y=0.845 $X2=0 $Y2=0
cc_648 N_S[3]_c_795_n N_VGND_c_1646_n 0.0271255f $X=10.59 $Y=0.18 $X2=0 $Y2=0
cc_649 N_S[3]_c_790_n VGND 0.0111218f $X=9.87 $Y=0.845 $X2=0 $Y2=0
cc_650 N_S[3]_c_794_n VGND 0.0119932f $X=10.925 $Y=0.18 $X2=0 $Y2=0
cc_651 N_S[3]_c_795_n VGND 0.00731624f $X=10.59 $Y=0.18 $X2=0 $Y2=0
cc_652 N_S[3]_c_797_n VGND 0.0111713f $X=11.345 $Y=0.18 $X2=0 $Y2=0
cc_653 N_S[3]_c_799_n VGND 0.00366655f $X=11 $Y=0.18 $X2=0 $Y2=0
cc_654 N_S[3]_c_793_n N_A_2133_69#_c_1874_n 0.00295202f $X=10.515 $Y=0.845 $X2=0
+ $Y2=0
cc_655 N_S[3]_c_796_n N_A_2133_69#_c_1870_n 0.0126455f $X=11 $Y=0.255 $X2=0
+ $Y2=0
cc_656 N_S[3]_c_797_n N_A_2133_69#_c_1870_n 0.00211351f $X=11.345 $Y=0.18 $X2=0
+ $Y2=0
cc_657 N_S[3]_c_798_n N_A_2133_69#_c_1870_n 0.0132844f $X=11.42 $Y=0.255 $X2=0
+ $Y2=0
cc_658 N_S[3]_c_793_n N_A_2133_69#_c_1871_n 0.00349455f $X=10.515 $Y=0.845 $X2=0
+ $Y2=0
cc_659 N_S[3]_c_794_n N_A_2133_69#_c_1871_n 0.00436105f $X=10.925 $Y=0.18 $X2=0
+ $Y2=0
cc_660 N_S[3]_c_798_n N_A_2133_69#_c_1873_n 0.00139422f $X=11.42 $Y=0.255 $X2=0
+ $Y2=0
cc_661 N_A_1989_47#_c_857_n N_D[3]_M1001_g 0.00671996f $X=11.3 $Y=1.4 $X2=0
+ $Y2=0
cc_662 N_A_1989_47#_M1032_g N_D[3]_M1001_g 0.0232231f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_663 N_A_1989_47#_c_860_n N_VPWR_c_1023_n 0.0321301f $X=10.165 $Y=2.31 $X2=0
+ $Y2=0
cc_664 N_A_1989_47#_c_855_n N_VPWR_c_1023_n 0.00732952f $X=10.45 $Y=1.42 $X2=0
+ $Y2=0
cc_665 N_A_1989_47#_M1032_g N_VPWR_c_1024_n 0.00107974f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_666 N_A_1989_47#_M1016_d VPWR 0.00179197f $X=10.02 $Y=1.485 $X2=0 $Y2=0
cc_667 N_A_1989_47#_M1004_g VPWR 0.00728421f $X=10.92 $Y=2.075 $X2=0 $Y2=0
cc_668 N_A_1989_47#_M1032_g VPWR 0.00617598f $X=11.39 $Y=2.075 $X2=0 $Y2=0
cc_669 N_A_1989_47#_c_860_n VPWR 0.00594162f $X=10.165 $Y=2.31 $X2=0 $Y2=0
cc_670 N_A_1989_47#_M1004_g N_VPWR_c_1033_n 0.00429453f $X=10.92 $Y=2.075 $X2=0
+ $Y2=0
cc_671 N_A_1989_47#_M1032_g N_VPWR_c_1033_n 0.00429453f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_672 N_A_1989_47#_c_860_n N_VPWR_c_1033_n 0.0210596f $X=10.165 $Y=2.31 $X2=0
+ $Y2=0
cc_673 N_A_1989_47#_c_857_n N_Z_c_1203_n 0.00348752f $X=11.3 $Y=1.4 $X2=0 $Y2=0
cc_674 N_A_1989_47#_c_853_n N_Z_c_1203_n 0.0033343f $X=10.45 $Y=1.205 $X2=0
+ $Y2=0
cc_675 N_A_1989_47#_M1004_g N_Z_c_1210_n 0.00753886f $X=10.92 $Y=2.075 $X2=0
+ $Y2=0
cc_676 N_A_1989_47#_c_852_n N_Z_c_1210_n 9.57301e-19 $X=11.01 $Y=1.4 $X2=0 $Y2=0
cc_677 N_A_1989_47#_c_860_n N_Z_c_1210_n 0.0308332f $X=10.165 $Y=2.31 $X2=0
+ $Y2=0
cc_678 N_A_1989_47#_c_855_n N_Z_c_1210_n 0.0132841f $X=10.45 $Y=1.42 $X2=0 $Y2=0
cc_679 N_A_1989_47#_M1032_g Z 0.00635853f $X=11.39 $Y=2.075 $X2=0 $Y2=0
cc_680 N_A_1989_47#_M1004_g N_Z_c_1320_n 0.00635536f $X=10.92 $Y=2.075 $X2=0
+ $Y2=0
cc_681 N_A_1989_47#_c_857_n N_Z_c_1320_n 8.37785e-19 $X=11.3 $Y=1.4 $X2=0 $Y2=0
cc_682 N_A_1989_47#_M1032_g N_Z_c_1320_n 0.0105371f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_683 N_A_1989_47#_M1004_g N_Z_c_1207_n 0.00476154f $X=10.92 $Y=2.075 $X2=0
+ $Y2=0
cc_684 N_A_1989_47#_c_857_n N_Z_c_1207_n 0.0140509f $X=11.3 $Y=1.4 $X2=0 $Y2=0
cc_685 N_A_1989_47#_c_852_n N_Z_c_1207_n 7.26438e-19 $X=11.01 $Y=1.4 $X2=0 $Y2=0
cc_686 N_A_1989_47#_M1032_g N_Z_c_1207_n 0.00268051f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_687 N_A_1989_47#_c_853_n N_Z_c_1207_n 0.00967956f $X=10.45 $Y=1.205 $X2=0
+ $Y2=0
cc_688 N_A_1989_47#_c_855_n N_Z_c_1207_n 0.0117695f $X=10.45 $Y=1.42 $X2=0 $Y2=0
cc_689 N_A_1989_47#_M1004_g N_A_2112_333#_c_1544_n 0.00745341f $X=10.92 $Y=2.075
+ $X2=0 $Y2=0
cc_690 N_A_1989_47#_c_852_n N_A_2112_333#_c_1544_n 0.00133381f $X=11.01 $Y=1.4
+ $X2=0 $Y2=0
cc_691 N_A_1989_47#_c_860_n N_A_2112_333#_c_1544_n 0.0347621f $X=10.165 $Y=2.31
+ $X2=0 $Y2=0
cc_692 N_A_1989_47#_c_855_n N_A_2112_333#_c_1544_n 0.0132748f $X=10.45 $Y=1.42
+ $X2=0 $Y2=0
cc_693 N_A_1989_47#_M1004_g N_A_2112_333#_c_1552_n 0.00971609f $X=10.92 $Y=2.075
+ $X2=0 $Y2=0
cc_694 N_A_1989_47#_M1032_g N_A_2112_333#_c_1552_n 0.0128147f $X=11.39 $Y=2.075
+ $X2=0 $Y2=0
cc_695 N_A_1989_47#_c_860_n N_A_2112_333#_c_1554_n 0.010563f $X=10.165 $Y=2.31
+ $X2=0 $Y2=0
cc_696 N_A_1989_47#_M1032_g N_A_2112_333#_c_1555_n 0.00736707f $X=11.39 $Y=2.075
+ $X2=0 $Y2=0
cc_697 N_A_1989_47#_M1032_g N_A_2112_333#_c_1556_n 0.00176121f $X=11.39 $Y=2.075
+ $X2=0 $Y2=0
cc_698 N_A_1989_47#_c_854_n N_VGND_c_1646_n 0.0173492f $X=10.08 $Y=0.495 $X2=0
+ $Y2=0
cc_699 N_A_1989_47#_M1007_d VGND 0.00250855f $X=9.945 $Y=0.235 $X2=0 $Y2=0
cc_700 N_A_1989_47#_c_854_n VGND 0.0186564f $X=10.08 $Y=0.495 $X2=0 $Y2=0
cc_701 N_A_1989_47#_c_852_n N_A_2133_69#_c_1874_n 0.00308807f $X=11.01 $Y=1.4
+ $X2=0 $Y2=0
cc_702 N_A_1989_47#_c_853_n N_A_2133_69#_c_1874_n 0.00101918f $X=10.45 $Y=1.205
+ $X2=0 $Y2=0
cc_703 N_A_1989_47#_c_854_n N_A_2133_69#_c_1874_n 0.0185512f $X=10.08 $Y=0.495
+ $X2=0 $Y2=0
cc_704 N_A_1989_47#_c_855_n N_A_2133_69#_c_1874_n 0.00285813f $X=10.45 $Y=1.42
+ $X2=0 $Y2=0
cc_705 N_A_1989_47#_c_854_n N_A_2133_69#_c_1871_n 0.00358194f $X=10.08 $Y=0.495
+ $X2=0 $Y2=0
cc_706 N_D[3]_M1001_g N_VPWR_c_1024_n 0.00919666f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_707 N_D[3]_M1036_g N_VPWR_c_1024_n 0.0031734f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_708 N_D[3]_M1001_g N_VPWR_c_1121_n 0.00343746f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_709 N_D[3]_M1036_g N_VPWR_c_1121_n 0.00363183f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_710 N_D[3]_M1001_g VPWR 0.0105515f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_711 N_D[3]_M1036_g VPWR 0.0120316f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_712 N_D[3]_M1001_g N_VPWR_c_1033_n 0.00622633f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_713 N_D[3]_M1036_g N_VPWR_c_1034_n 0.00652917f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_714 N_D[3]_M1001_g N_Z_c_1207_n 0.00112534f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_715 N_D[3]_M1008_g N_Z_c_1207_n 8.13311e-19 $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_716 D[3] N_Z_c_1207_n 0.00742792f $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_717 N_D[3]_c_930_n N_Z_c_1207_n 0.00583073f $X=12.47 $Y=1.16 $X2=0 $Y2=0
cc_718 N_D[3]_M1001_g N_A_2112_333#_c_1555_n 0.00557487f $X=11.915 $Y=1.985
+ $X2=0 $Y2=0
cc_719 N_D[3]_M1001_g N_A_2112_333#_c_1558_n 0.0174487f $X=11.915 $Y=1.985 $X2=0
+ $Y2=0
cc_720 N_D[3]_M1036_g N_A_2112_333#_c_1558_n 0.0142998f $X=12.385 $Y=1.985 $X2=0
+ $Y2=0
cc_721 D[3] N_A_2112_333#_c_1558_n 0.0339353f $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_722 N_D[3]_c_930_n N_A_2112_333#_c_1558_n 7.13708e-19 $X=12.47 $Y=1.16 $X2=0
+ $Y2=0
cc_723 D[3] N_A_2112_333#_c_1545_n 0.0235932f $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_724 N_D[3]_c_930_n N_A_2112_333#_c_1545_n 9.6385e-19 $X=12.47 $Y=1.16 $X2=0
+ $Y2=0
cc_725 N_D[3]_M1036_g N_A_2112_333#_c_1546_n 0.00329008f $X=12.385 $Y=1.985
+ $X2=0 $Y2=0
cc_726 N_D[3]_M1008_g N_VGND_c_1641_n 0.00300333f $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_727 N_D[3]_M1039_g N_VGND_c_1641_n 0.0030929f $X=12.36 $Y=0.56 $X2=0 $Y2=0
cc_728 N_D[3]_M1008_g N_VGND_c_1646_n 0.00436487f $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_729 N_D[3]_M1008_g VGND 0.00600262f $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_730 N_D[3]_M1039_g VGND 0.00697949f $X=12.36 $Y=0.56 $X2=0 $Y2=0
cc_731 N_D[3]_M1039_g N_VGND_c_1650_n 0.00430643f $X=12.36 $Y=0.56 $X2=0 $Y2=0
cc_732 N_D[3]_M1008_g N_A_2133_69#_c_1872_n 0.0114493f $X=11.94 $Y=0.56 $X2=0
+ $Y2=0
cc_733 N_D[3]_M1039_g N_A_2133_69#_c_1872_n 0.00931728f $X=12.36 $Y=0.56 $X2=0
+ $Y2=0
cc_734 D[3] N_A_2133_69#_c_1872_n 0.0518587f $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_735 N_D[3]_c_930_n N_A_2133_69#_c_1872_n 0.00665175f $X=12.47 $Y=1.16 $X2=0
+ $Y2=0
cc_736 N_D[3]_M1008_g N_A_2133_69#_c_1873_n 0.00114614f $X=11.94 $Y=0.56 $X2=0
+ $Y2=0
cc_737 N_D[3]_c_930_n N_A_2133_69#_c_1873_n 0.00120541f $X=12.47 $Y=1.16 $X2=0
+ $Y2=0
cc_738 N_D[3]_M1008_g N_A_2133_69#_c_1892_n 5.29024e-19 $X=11.94 $Y=0.56 $X2=0
+ $Y2=0
cc_739 N_D[3]_M1039_g N_A_2133_69#_c_1892_n 0.00633603f $X=12.36 $Y=0.56 $X2=0
+ $Y2=0
cc_740 N_A_27_297#_c_977_n N_VPWR_M1002_s 0.00350459f $X=1.115 $Y=1.58 $X2=-0.19
+ $Y2=1.305
cc_741 N_A_27_297#_c_993_p N_VPWR_c_1019_n 0.0114322f $X=1.285 $Y=2.38 $X2=0
+ $Y2=0
cc_742 N_A_27_297#_c_977_n N_VPWR_c_1041_n 0.0170301f $X=1.115 $Y=1.58 $X2=0
+ $Y2=0
cc_743 N_A_27_297#_c_981_n N_VPWR_c_1041_n 0.0272234f $X=1.2 $Y=1.78 $X2=0 $Y2=0
cc_744 N_A_27_297#_c_985_n N_VPWR_c_1025_n 0.0569572f $X=2.11 $Y=2.38 $X2=0
+ $Y2=0
cc_745 N_A_27_297#_c_993_p N_VPWR_c_1025_n 0.0119545f $X=1.285 $Y=2.38 $X2=0
+ $Y2=0
cc_746 N_A_27_297#_M1002_d VPWR 0.00217517f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_747 N_A_27_297#_M1017_d VPWR 0.00481062f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_748 N_A_27_297#_M1009_d VPWR 0.00210318f $X=2.05 $Y=1.665 $X2=0 $Y2=0
cc_749 N_A_27_297#_c_985_n VPWR 0.0196248f $X=2.11 $Y=2.38 $X2=0 $Y2=0
cc_750 N_A_27_297#_c_993_p VPWR 0.006547f $X=1.285 $Y=2.38 $X2=0 $Y2=0
cc_751 N_A_27_297#_c_973_n VPWR 0.0124483f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_752 N_A_27_297#_c_973_n N_VPWR_c_1030_n 0.020978f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_753 N_A_27_297#_c_985_n N_Z_M1005_s 0.00341588f $X=2.11 $Y=2.38 $X2=0 $Y2=0
cc_754 N_A_27_297#_M1009_d N_Z_c_1208_n 0.00237684f $X=2.05 $Y=1.665 $X2=0 $Y2=0
cc_755 N_A_27_297#_c_985_n N_Z_c_1208_n 0.00494997f $X=2.11 $Y=2.38 $X2=0 $Y2=0
cc_756 N_A_27_297#_c_972_n N_Z_c_1208_n 0.0132602f $X=2.195 $Y=1.81 $X2=0 $Y2=0
cc_757 N_A_27_297#_c_981_n N_Z_c_1226_n 0.0062686f $X=1.2 $Y=1.78 $X2=0 $Y2=0
cc_758 N_A_27_297#_c_985_n N_Z_c_1226_n 8.66896e-19 $X=2.11 $Y=2.38 $X2=0 $Y2=0
cc_759 N_A_27_297#_c_972_n N_Z_c_1226_n 4.86317e-19 $X=2.195 $Y=1.81 $X2=0 $Y2=0
cc_760 N_A_27_297#_c_981_n N_Z_c_1227_n 0.0235305f $X=1.2 $Y=1.78 $X2=0 $Y2=0
cc_761 N_A_27_297#_c_985_n N_Z_c_1227_n 0.0211175f $X=2.11 $Y=2.38 $X2=0 $Y2=0
cc_762 N_A_27_297#_c_972_n N_Z_c_1227_n 0.0212802f $X=2.195 $Y=1.81 $X2=0 $Y2=0
cc_763 N_A_27_297#_c_977_n N_Z_c_1204_n 0.00930189f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_764 N_A_27_297#_c_972_n N_Z_c_1204_n 0.00468052f $X=2.195 $Y=1.81 $X2=0 $Y2=0
cc_765 N_A_27_297#_c_977_n N_A_27_47#_c_1593_n 0.0110288f $X=1.115 $Y=1.58 $X2=0
+ $Y2=0
cc_766 VPWR N_Z_M1005_s 0.00187512f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_767 VPWR N_Z_M1020_s 0.00187512f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_768 VPWR N_Z_M1003_d 0.00187512f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_769 VPWR N_Z_M1004_d 0.00187512f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_770 N_VPWR_M1006_d N_Z_c_1208_n 5.82057e-19 $X=3.04 $Y=1.485 $X2=0 $Y2=0
cc_771 N_VPWR_c_1020_n N_Z_c_1208_n 0.0287846f $X=3.22 $Y=1.63 $X2=0 $Y2=0
cc_772 VPWR N_Z_c_1208_n 0.138617f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_773 VPWR N_Z_c_1226_n 0.0144354f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_774 N_VPWR_M1015_s N_Z_c_1209_n 0.00219731f $X=5.565 $Y=1.485 $X2=0 $Y2=0
cc_775 N_VPWR_M1000_d N_Z_c_1209_n 0.00219731f $X=7.025 $Y=1.485 $X2=0 $Y2=0
cc_776 N_VPWR_c_1077_n N_Z_c_1209_n 0.0159439f $X=5.71 $Y=1.94 $X2=0 $Y2=0
cc_777 N_VPWR_c_1085_n N_Z_c_1209_n 0.0159439f $X=7.17 $Y=1.94 $X2=0 $Y2=0
cc_778 VPWR N_Z_c_1209_n 0.136626f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_779 VPWR N_Z_c_1257_n 0.0144354f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_780 N_VPWR_M1035_d N_Z_c_1210_n 5.82057e-19 $X=9.48 $Y=1.485 $X2=0 $Y2=0
cc_781 N_VPWR_c_1023_n N_Z_c_1210_n 0.0287846f $X=9.66 $Y=1.63 $X2=0 $Y2=0
cc_782 VPWR N_Z_c_1210_n 0.138617f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_783 VPWR N_Z_c_1289_n 0.0144354f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_784 VPWR Z 0.0144354f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_785 VPWR N_A_824_333#_M1020_d 0.00210318f $X=12.565 $Y=2.635 $X2=-0.19
+ $Y2=-0.24
cc_786 VPWR N_A_824_333#_M1027_d 0.00273129f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_787 VPWR N_A_824_333#_M1023_d 0.00179197f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_788 N_VPWR_c_1021_n N_A_824_333#_c_1436_n 0.0114322f $X=5.71 $Y=2.34 $X2=0
+ $Y2=0
cc_789 VPWR N_A_824_333#_c_1436_n 0.0161639f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_790 N_VPWR_c_1031_n N_A_824_333#_c_1436_n 0.0570268f $X=5.545 $Y=2.72 $X2=0
+ $Y2=0
cc_791 VPWR N_A_824_333#_c_1438_n 0.0031082f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_792 N_VPWR_c_1031_n N_A_824_333#_c_1438_n 0.0118848f $X=5.545 $Y=2.72 $X2=0
+ $Y2=0
cc_793 N_VPWR_c_1077_n N_A_824_333#_c_1439_n 0.0265477f $X=5.71 $Y=1.94 $X2=0
+ $Y2=0
cc_794 N_VPWR_M1015_s N_A_824_333#_c_1442_n 0.00331615f $X=5.565 $Y=1.485 $X2=0
+ $Y2=0
cc_795 N_VPWR_c_1077_n N_A_824_333#_c_1442_n 0.0158304f $X=5.71 $Y=1.94 $X2=0
+ $Y2=0
cc_796 VPWR N_A_824_333#_c_1430_n 0.00591741f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_797 N_VPWR_c_1032_n N_A_824_333#_c_1430_n 0.020978f $X=7.035 $Y=2.72 $X2=0
+ $Y2=0
cc_798 N_VPWR_c_1077_n N_A_824_333#_c_1431_n 0.0115021f $X=5.71 $Y=1.94 $X2=0
+ $Y2=0
cc_799 VPWR N_A_1315_297#_M1000_s 0.00179197f $X=12.565 $Y=2.635 $X2=-0.19
+ $Y2=-0.24
cc_800 VPWR N_A_1315_297#_M1030_s 0.00273129f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_801 VPWR N_A_1315_297#_M1031_s 0.00210318f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_802 N_VPWR_M1000_d N_A_1315_297#_c_1493_n 0.00331615f $X=7.025 $Y=1.485 $X2=0
+ $Y2=0
cc_803 N_VPWR_c_1085_n N_A_1315_297#_c_1493_n 0.0158304f $X=7.17 $Y=1.94 $X2=0
+ $Y2=0
cc_804 N_VPWR_c_1085_n N_A_1315_297#_c_1497_n 0.0265477f $X=7.17 $Y=1.94 $X2=0
+ $Y2=0
cc_805 N_VPWR_c_1027_n N_A_1315_297#_c_1501_n 0.0569572f $X=9.495 $Y=2.72 $X2=0
+ $Y2=0
cc_806 VPWR N_A_1315_297#_c_1501_n 0.0161535f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_807 N_VPWR_c_1022_n N_A_1315_297#_c_1516_n 0.0114322f $X=7.17 $Y=2.34 $X2=0
+ $Y2=0
cc_808 N_VPWR_c_1027_n N_A_1315_297#_c_1516_n 0.0119545f $X=9.495 $Y=2.72 $X2=0
+ $Y2=0
cc_809 VPWR N_A_1315_297#_c_1516_n 0.00311866f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_810 VPWR N_A_1315_297#_c_1489_n 0.00591741f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_811 N_VPWR_c_1032_n N_A_1315_297#_c_1489_n 0.020978f $X=7.035 $Y=2.72 $X2=0
+ $Y2=0
cc_812 N_VPWR_c_1085_n N_A_1315_297#_c_1490_n 0.0115021f $X=7.17 $Y=1.94 $X2=0
+ $Y2=0
cc_813 VPWR N_A_2112_333#_M1004_s 0.00210318f $X=12.565 $Y=2.635 $X2=-0.19
+ $Y2=-0.24
cc_814 VPWR N_A_2112_333#_M1032_s 0.00481062f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_815 VPWR N_A_2112_333#_M1036_s 0.00217517f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_816 N_VPWR_c_1024_n N_A_2112_333#_c_1552_n 0.0114322f $X=12.15 $Y=2.34 $X2=0
+ $Y2=0
cc_817 VPWR N_A_2112_333#_c_1552_n 0.0230635f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_818 N_VPWR_c_1033_n N_A_2112_333#_c_1552_n 0.0570268f $X=11.985 $Y=2.72 $X2=0
+ $Y2=0
cc_819 VPWR N_A_2112_333#_c_1554_n 0.0031082f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_820 N_VPWR_c_1033_n N_A_2112_333#_c_1554_n 0.0118848f $X=11.985 $Y=2.72 $X2=0
+ $Y2=0
cc_821 N_VPWR_c_1121_n N_A_2112_333#_c_1555_n 0.0272234f $X=12.15 $Y=1.94 $X2=0
+ $Y2=0
cc_822 N_VPWR_M1001_d N_A_2112_333#_c_1558_n 0.00350459f $X=12.005 $Y=1.485
+ $X2=0 $Y2=0
cc_823 N_VPWR_c_1121_n N_A_2112_333#_c_1558_n 0.0170301f $X=12.15 $Y=1.94 $X2=0
+ $Y2=0
cc_824 VPWR N_A_2112_333#_c_1546_n 0.0124483f $X=12.565 $Y=2.635 $X2=0 $Y2=0
cc_825 N_VPWR_c_1034_n N_A_2112_333#_c_1546_n 0.020978f $X=12.65 $Y=2.72 $X2=0
+ $Y2=0
cc_826 N_Z_c_1208_n N_A_824_333#_M1020_d 0.00237684f $X=4.685 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_827 N_Z_c_1209_n N_A_824_333#_M1027_d 0.00645967f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_828 N_Z_c_1208_n N_A_824_333#_c_1428_n 0.0132602f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_829 N_Z_c_1257_n N_A_824_333#_c_1428_n 4.86317e-19 $X=4.975 $Y=1.87 $X2=0
+ $Y2=0
cc_830 N_Z_c_1258_n N_A_824_333#_c_1428_n 0.0212802f $X=4.83 $Y=1.87 $X2=0 $Y2=0
cc_831 N_Z_c_1205_n N_A_824_333#_c_1428_n 0.00468052f $X=4.76 $Y=1.755 $X2=0
+ $Y2=0
cc_832 N_Z_M1020_s N_A_824_333#_c_1436_n 0.00341588f $X=4.57 $Y=1.665 $X2=0
+ $Y2=0
cc_833 N_Z_c_1208_n N_A_824_333#_c_1436_n 0.00494997f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_834 N_Z_c_1209_n N_A_824_333#_c_1436_n 0.00415493f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_835 N_Z_c_1257_n N_A_824_333#_c_1436_n 8.66896e-19 $X=4.975 $Y=1.87 $X2=0
+ $Y2=0
cc_836 N_Z_c_1258_n N_A_824_333#_c_1436_n 0.0211175f $X=4.83 $Y=1.87 $X2=0 $Y2=0
cc_837 N_Z_c_1209_n N_A_824_333#_c_1439_n 0.0190087f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_838 N_Z_c_1257_n N_A_824_333#_c_1439_n 0.00221246f $X=4.975 $Y=1.87 $X2=0
+ $Y2=0
cc_839 N_Z_c_1258_n N_A_824_333#_c_1439_n 0.024193f $X=4.83 $Y=1.87 $X2=0 $Y2=0
cc_840 N_Z_c_1209_n N_A_824_333#_c_1442_n 0.0237468f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_841 N_Z_c_1205_n N_A_824_333#_c_1440_n 0.00930189f $X=4.76 $Y=1.755 $X2=0
+ $Y2=0
cc_842 N_Z_c_1209_n N_A_824_333#_c_1430_n 3.2447e-19 $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_843 N_Z_c_1209_n N_A_824_333#_c_1431_n 0.0219733f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_844 N_Z_c_1209_n N_A_1315_297#_M1030_s 0.00645967f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_845 N_Z_c_1210_n N_A_1315_297#_M1031_s 0.00237684f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_846 N_Z_c_1209_n N_A_1315_297#_c_1493_n 0.0237468f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_847 N_Z_c_1206_n N_A_1315_297#_c_1493_n 0.00930189f $X=8.12 $Y=1.755 $X2=0
+ $Y2=0
cc_848 N_Z_c_1209_n N_A_1315_297#_c_1497_n 0.0190087f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_849 N_Z_c_1289_n N_A_1315_297#_c_1497_n 0.00221246f $X=8.195 $Y=1.87 $X2=0
+ $Y2=0
cc_850 N_Z_c_1290_n N_A_1315_297#_c_1497_n 0.024193f $X=8.05 $Y=1.87 $X2=0 $Y2=0
cc_851 N_Z_M1003_d N_A_1315_297#_c_1501_n 0.00341588f $X=8.02 $Y=1.665 $X2=0
+ $Y2=0
cc_852 N_Z_c_1209_n N_A_1315_297#_c_1501_n 0.00415493f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_853 N_Z_c_1210_n N_A_1315_297#_c_1501_n 0.00494997f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_854 N_Z_c_1289_n N_A_1315_297#_c_1501_n 8.66896e-19 $X=8.195 $Y=1.87 $X2=0
+ $Y2=0
cc_855 N_Z_c_1290_n N_A_1315_297#_c_1501_n 0.0211175f $X=8.05 $Y=1.87 $X2=0
+ $Y2=0
cc_856 N_Z_c_1210_n N_A_1315_297#_c_1488_n 0.0132602f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_857 N_Z_c_1289_n N_A_1315_297#_c_1488_n 4.86317e-19 $X=8.195 $Y=1.87 $X2=0
+ $Y2=0
cc_858 N_Z_c_1290_n N_A_1315_297#_c_1488_n 0.0212802f $X=8.05 $Y=1.87 $X2=0
+ $Y2=0
cc_859 N_Z_c_1206_n N_A_1315_297#_c_1488_n 0.00468052f $X=8.12 $Y=1.755 $X2=0
+ $Y2=0
cc_860 N_Z_c_1209_n N_A_1315_297#_c_1489_n 3.2447e-19 $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_861 N_Z_c_1209_n N_A_1315_297#_c_1490_n 0.0219733f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_862 N_Z_c_1210_n N_A_2112_333#_M1004_s 0.00237684f $X=11.125 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_863 N_Z_c_1210_n N_A_2112_333#_c_1544_n 0.0132602f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_864 Z N_A_2112_333#_c_1544_n 4.86317e-19 $X=11.185 $Y=1.785 $X2=0 $Y2=0
cc_865 N_Z_c_1320_n N_A_2112_333#_c_1544_n 0.0212802f $X=11.27 $Y=1.87 $X2=0
+ $Y2=0
cc_866 N_Z_c_1207_n N_A_2112_333#_c_1544_n 0.00468052f $X=11.2 $Y=1.755 $X2=0
+ $Y2=0
cc_867 N_Z_M1004_d N_A_2112_333#_c_1552_n 0.00341588f $X=11.01 $Y=1.665 $X2=0
+ $Y2=0
cc_868 N_Z_c_1210_n N_A_2112_333#_c_1552_n 0.00494997f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_869 Z N_A_2112_333#_c_1552_n 8.66896e-19 $X=11.185 $Y=1.785 $X2=0 $Y2=0
cc_870 N_Z_c_1320_n N_A_2112_333#_c_1552_n 0.0211175f $X=11.27 $Y=1.87 $X2=0
+ $Y2=0
cc_871 Z N_A_2112_333#_c_1555_n 0.0062686f $X=11.185 $Y=1.785 $X2=0 $Y2=0
cc_872 N_Z_c_1320_n N_A_2112_333#_c_1555_n 0.0235305f $X=11.27 $Y=1.87 $X2=0
+ $Y2=0
cc_873 N_Z_c_1207_n N_A_2112_333#_c_1556_n 0.00930189f $X=11.2 $Y=1.755 $X2=0
+ $Y2=0
cc_874 N_Z_c_1200_n N_A_27_47#_c_1593_n 0.00729487f $X=1.67 $Y=0.68 $X2=0 $Y2=0
cc_875 N_Z_c_1204_n N_A_27_47#_c_1593_n 0.00238404f $X=1.68 $Y=1.755 $X2=0 $Y2=0
cc_876 N_Z_M1011_s N_A_27_47#_c_1595_n 0.00165831f $X=1.535 $Y=0.345 $X2=0 $Y2=0
cc_877 N_Z_c_1200_n N_A_27_47#_c_1595_n 0.0156951f $X=1.67 $Y=0.68 $X2=0 $Y2=0
cc_878 N_Z_M1010_s N_A_845_69#_c_1778_n 0.00165831f $X=4.635 $Y=0.345 $X2=0
+ $Y2=0
cc_879 N_Z_c_1201_n N_A_845_69#_c_1778_n 0.0156951f $X=4.77 $Y=0.68 $X2=0 $Y2=0
cc_880 N_Z_c_1201_n N_A_845_69#_c_1781_n 0.00729487f $X=4.77 $Y=0.68 $X2=0 $Y2=0
cc_881 N_Z_c_1205_n N_A_845_69#_c_1781_n 0.00238404f $X=4.76 $Y=1.755 $X2=0
+ $Y2=0
cc_882 N_Z_c_1202_n N_A_1315_47#_c_1826_n 0.00729487f $X=8.11 $Y=0.68 $X2=0
+ $Y2=0
cc_883 N_Z_c_1206_n N_A_1315_47#_c_1826_n 0.00238404f $X=8.12 $Y=1.755 $X2=0
+ $Y2=0
cc_884 N_Z_M1029_d N_A_1315_47#_c_1828_n 0.00165831f $X=7.975 $Y=0.345 $X2=0
+ $Y2=0
cc_885 N_Z_c_1202_n N_A_1315_47#_c_1828_n 0.0156951f $X=8.11 $Y=0.68 $X2=0 $Y2=0
cc_886 N_Z_M1025_d N_A_2133_69#_c_1870_n 0.00165831f $X=11.075 $Y=0.345 $X2=0
+ $Y2=0
cc_887 N_Z_c_1203_n N_A_2133_69#_c_1870_n 0.0156951f $X=11.21 $Y=0.68 $X2=0
+ $Y2=0
cc_888 N_Z_c_1203_n N_A_2133_69#_c_1873_n 0.00729487f $X=11.21 $Y=0.68 $X2=0
+ $Y2=0
cc_889 N_Z_c_1207_n N_A_2133_69#_c_1873_n 0.00238404f $X=11.2 $Y=1.755 $X2=0
+ $Y2=0
cc_890 N_A_824_333#_c_1429_n N_A_1315_297#_c_1487_n 0.0147157f $X=6.195 $Y=1.665
+ $X2=0 $Y2=0
cc_891 N_A_824_333#_c_1430_n N_A_1315_297#_c_1489_n 0.0296136f $X=6.18 $Y=2.34
+ $X2=0 $Y2=0
cc_892 N_A_824_333#_c_1431_n N_A_1315_297#_c_1490_n 0.0296136f $X=6.18 $Y=2.21
+ $X2=0 $Y2=0
cc_893 N_A_824_333#_c_1442_n N_A_845_69#_c_1780_n 0.00251701f $X=6.045 $Y=1.58
+ $X2=0 $Y2=0
cc_894 N_A_824_333#_c_1442_n N_A_845_69#_c_1781_n 0.00200781f $X=6.045 $Y=1.58
+ $X2=0 $Y2=0
cc_895 N_A_824_333#_c_1440_n N_A_845_69#_c_1781_n 0.00650395f $X=5.325 $Y=1.58
+ $X2=0 $Y2=0
cc_896 N_A_1315_297#_c_1493_n N_A_1315_47#_c_1826_n 0.0110288f $X=7.555 $Y=1.58
+ $X2=0 $Y2=0
cc_897 N_A_2112_333#_c_1558_n N_A_2133_69#_c_1872_n 0.00251701f $X=12.485
+ $Y=1.58 $X2=0 $Y2=0
cc_898 N_A_2112_333#_c_1558_n N_A_2133_69#_c_1873_n 0.00200781f $X=12.485
+ $Y=1.58 $X2=0 $Y2=0
cc_899 N_A_2112_333#_c_1556_n N_A_2133_69#_c_1873_n 0.00650395f $X=11.765
+ $Y=1.58 $X2=0 $Y2=0
cc_900 N_A_27_47#_c_1593_n N_VGND_M1013_s 0.00306532f $X=1.03 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_901 N_A_27_47#_c_1593_n N_VGND_c_1635_n 0.012179f $X=1.03 $Y=0.8 $X2=0 $Y2=0
cc_902 N_A_27_47#_c_1593_n N_VGND_c_1642_n 0.00219745f $X=1.03 $Y=0.8 $X2=0
+ $Y2=0
cc_903 N_A_27_47#_c_1625_p N_VGND_c_1642_n 0.0199987f $X=1.182 $Y=0.425 $X2=0
+ $Y2=0
cc_904 N_A_27_47#_c_1595_n N_VGND_c_1642_n 0.0535945f $X=2.005 $Y=0.34 $X2=0
+ $Y2=0
cc_905 N_A_27_47#_M1013_d VGND 0.00288496f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_906 N_A_27_47#_M1026_d VGND 0.0024283f $X=1.015 $Y=0.235 $X2=0 $Y2=0
cc_907 N_A_27_47#_c_1596_n VGND 0.0124017f $X=0.31 $Y=0.38 $X2=0 $Y2=0
cc_908 N_A_27_47#_c_1593_n VGND 0.00838939f $X=1.03 $Y=0.8 $X2=0 $Y2=0
cc_909 N_A_27_47#_c_1625_p VGND 0.0117415f $X=1.182 $Y=0.425 $X2=0 $Y2=0
cc_910 N_A_27_47#_c_1595_n VGND 0.0279432f $X=2.005 $Y=0.34 $X2=0 $Y2=0
cc_911 N_A_27_47#_c_1596_n N_VGND_c_1651_n 0.020879f $X=0.31 $Y=0.38 $X2=0 $Y2=0
cc_912 N_A_27_47#_c_1593_n N_VGND_c_1651_n 0.0020257f $X=1.03 $Y=0.8 $X2=0 $Y2=0
cc_913 VGND N_A_845_69#_M1012_d 0.0024283f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_914 VGND N_A_845_69#_M1024_s 0.00288496f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_915 VGND N_A_845_69#_c_1778_n 0.0222193f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_916 N_VGND_c_1649_n N_A_845_69#_c_1778_n 0.0422314f $X=5.58 $Y=0 $X2=0 $Y2=0
cc_917 VGND N_A_845_69#_c_1779_n 0.00572388f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_918 N_VGND_c_1649_n N_A_845_69#_c_1779_n 0.0113631f $X=5.58 $Y=0 $X2=0 $Y2=0
cc_919 VGND N_A_845_69#_c_1815_n 0.0117415f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_920 N_VGND_c_1649_n N_A_845_69#_c_1815_n 0.0199987f $X=5.58 $Y=0 $X2=0 $Y2=0
cc_921 N_VGND_M1019_d N_A_845_69#_c_1780_n 0.00306532f $X=5.575 $Y=0.235 $X2=0
+ $Y2=0
cc_922 N_VGND_c_1637_n N_A_845_69#_c_1780_n 0.012179f $X=5.71 $Y=0.38 $X2=0
+ $Y2=0
cc_923 N_VGND_c_1638_n N_A_845_69#_c_1780_n 0.0020257f $X=7.085 $Y=0 $X2=0 $Y2=0
cc_924 VGND N_A_845_69#_c_1780_n 0.00838939f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_925 N_VGND_c_1649_n N_A_845_69#_c_1780_n 0.00219745f $X=5.58 $Y=0 $X2=0 $Y2=0
cc_926 N_VGND_c_1638_n N_A_845_69#_c_1800_n 0.020879f $X=7.085 $Y=0 $X2=0 $Y2=0
cc_927 VGND N_A_845_69#_c_1800_n 0.0124017f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_928 VGND N_A_1315_47#_M1028_d 0.00288496f $X=12.565 $Y=-0.085 $X2=-0.19
+ $Y2=-0.24
cc_929 VGND N_A_1315_47#_M1033_d 0.0024283f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_930 N_VGND_c_1638_n N_A_1315_47#_c_1829_n 0.020879f $X=7.085 $Y=0 $X2=0 $Y2=0
cc_931 VGND N_A_1315_47#_c_1829_n 0.0124017f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_932 N_VGND_M1028_s N_A_1315_47#_c_1826_n 0.00306532f $X=7.035 $Y=0.235 $X2=0
+ $Y2=0
cc_933 N_VGND_c_1638_n N_A_1315_47#_c_1826_n 0.0020257f $X=7.085 $Y=0 $X2=0
+ $Y2=0
cc_934 N_VGND_c_1639_n N_A_1315_47#_c_1826_n 0.012179f $X=7.17 $Y=0.38 $X2=0
+ $Y2=0
cc_935 N_VGND_c_1644_n N_A_1315_47#_c_1826_n 0.00219745f $X=9.535 $Y=0 $X2=0
+ $Y2=0
cc_936 VGND N_A_1315_47#_c_1826_n 0.00838939f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_937 N_VGND_c_1644_n N_A_1315_47#_c_1864_n 0.0199987f $X=9.535 $Y=0 $X2=0
+ $Y2=0
cc_938 VGND N_A_1315_47#_c_1864_n 0.0117415f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_939 N_VGND_c_1644_n N_A_1315_47#_c_1828_n 0.0535945f $X=9.535 $Y=0 $X2=0
+ $Y2=0
cc_940 VGND N_A_1315_47#_c_1828_n 0.0279432f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_941 VGND N_A_2133_69#_M1034_s 0.0024283f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_942 VGND N_A_2133_69#_M1039_d 0.00288496f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_943 N_VGND_c_1646_n N_A_2133_69#_c_1870_n 0.0422314f $X=12.02 $Y=0 $X2=0
+ $Y2=0
cc_944 VGND N_A_2133_69#_c_1870_n 0.0222193f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_945 N_VGND_c_1646_n N_A_2133_69#_c_1871_n 0.0113631f $X=12.02 $Y=0 $X2=0
+ $Y2=0
cc_946 VGND N_A_2133_69#_c_1871_n 0.00572388f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_947 N_VGND_c_1646_n N_A_2133_69#_c_1907_n 0.0199987f $X=12.02 $Y=0 $X2=0
+ $Y2=0
cc_948 VGND N_A_2133_69#_c_1907_n 0.0117415f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_949 N_VGND_M1008_s N_A_2133_69#_c_1872_n 0.00306532f $X=12.015 $Y=0.235 $X2=0
+ $Y2=0
cc_950 N_VGND_c_1641_n N_A_2133_69#_c_1872_n 0.012179f $X=12.15 $Y=0.38 $X2=0
+ $Y2=0
cc_951 N_VGND_c_1646_n N_A_2133_69#_c_1872_n 0.00219745f $X=12.02 $Y=0 $X2=0
+ $Y2=0
cc_952 VGND N_A_2133_69#_c_1872_n 0.00838939f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_953 N_VGND_c_1650_n N_A_2133_69#_c_1872_n 0.0020257f $X=12.65 $Y=0 $X2=0
+ $Y2=0
cc_954 VGND N_A_2133_69#_c_1892_n 0.0124017f $X=12.565 $Y=-0.085 $X2=0 $Y2=0
cc_955 N_VGND_c_1650_n N_A_2133_69#_c_1892_n 0.020879f $X=12.65 $Y=0 $X2=0 $Y2=0
cc_956 N_A_845_69#_c_1800_n N_A_1315_47#_c_1829_n 0.0248576f $X=6.13 $Y=0.38
+ $X2=0 $Y2=0
cc_957 N_A_845_69#_c_1780_n N_A_1315_47#_c_1827_n 0.0103099f $X=5.965 $Y=0.8
+ $X2=0 $Y2=0
