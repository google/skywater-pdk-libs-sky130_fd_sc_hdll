* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
X0 a_27_297# B a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_883_297# a_1311_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_1311_21# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 Y a_1311_21# a_883_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 Y a_1311_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y a_1311_21# a_883_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_493_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 a_493_297# C a_883_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_883_297# a_1311_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_493_297# C a_883_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 a_1311_21# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_27_297# B a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 a_883_297# C a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 Y a_1311_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 VGND a_1311_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_883_297# C a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X31 VGND a_1311_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 a_493_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
