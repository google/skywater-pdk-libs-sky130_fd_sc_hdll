* NGSPICE file created from sky130_fd_sc_hdll__xor2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__xor2_2 A B VGND VNB VPB VPWR X
M1000 X B a_510_47# VNB nshort w=650000u l=150000u
+  ad=5.1675e+11p pd=4.19e+06u as=5.785e+11p ps=5.68e+06u
M1001 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=9.25e+11p pd=7.85e+06u as=8.45e+11p ps=7.69e+06u
M1002 VGND A a_112_47# VNB nshort w=650000u l=150000u
+  ad=1.06925e+12p pd=1.109e+07u as=4.485e+11p ps=3.98e+06u
M1003 VGND A a_510_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_510_47# B X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_510_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.39e+12p pd=1.278e+07u as=0p ps=0u
M1006 a_27_297# B a_112_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1007 a_510_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_112_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_112_47# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B a_510_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_510_297# a_112_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1012 X a_112_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_112_47# a_510_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_112_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B a_112_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_112_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_510_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A a_510_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

