* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__or3b_1 A B C_N VGND VNB VPB VPWR X
X0 a_225_53# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_225_53# a_117_297# a_315_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X2 VPWR C_N a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X3 VGND B a_225_53# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND a_225_53# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_315_297# B a_399_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X6 VGND C_N a_117_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR a_225_53# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 a_225_53# a_117_297# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_399_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
.ends
