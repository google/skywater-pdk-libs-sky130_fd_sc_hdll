* File: sky130_fd_sc_hdll__nand2_1.pex.spice
* Created: Wed Sep  2 08:36:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND2_1%B 1 3 4 6 7 12
r24 12 13 3.31956 $w=3.63e-07 $l=2.5e-08 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.54 $Y2=1.202
r25 10 12 33.1956 $w=3.63e-07 $l=2.5e-07 $layer=POLY_cond $X=0.265 $Y=1.202
+ $X2=0.515 $Y2=1.202
r26 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.265
+ $Y=1.16 $X2=0.265 $Y2=1.16
r27 4 13 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.54 $Y2=1.202
r28 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.54 $Y=0.995 $X2=0.54
+ $Y2=0.56
r29 1 12 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r30 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_1%A 1 3 4 6 7
r22 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.205
+ $Y=1.16 $X2=1.205 $Y2=1.16
r23 4 10 44.7166 $w=4.3e-07 $l=3.14245e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=1.13 $Y2=1.16
r24 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r25 1 10 40.2182 $w=4.3e-07 $l=2.38642e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=1.13 $Y2=1.16
r26 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.96 $Y=0.995 $X2=0.96
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_1%VPWR 1 2 7 9 13 17 21 25 26 32
r24 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r25 26 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r26 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r27 23 32 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.395 $Y=2.72
+ $X2=1.265 $Y2=2.72
r28 23 25 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.395 $Y=2.72
+ $X2=1.61 $Y2=2.72
r29 21 33 0.263201 $w=4.8e-07 $l=9.25e-07 $layer=MET1_cond $X=0.225 $Y=2.72
+ $X2=1.15 $Y2=2.72
r30 21 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r31 17 20 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.265 $Y=1.66
+ $X2=1.265 $Y2=2.34
r32 15 32 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=2.635
+ $X2=1.265 $Y2=2.72
r33 15 20 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=1.265 $Y=2.635
+ $X2=1.265 $Y2=2.34
r34 14 29 4.33083 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=2.72
+ $X2=0.182 $Y2=2.72
r35 13 32 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.135 $Y=2.72
+ $X2=1.265 $Y2=2.72
r36 13 14 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=2.72
+ $X2=0.365 $Y2=2.72
r37 9 12 27.9879 $w=2.78e-07 $l=6.8e-07 $layer=LI1_cond $X=0.225 $Y=1.66
+ $X2=0.225 $Y2=2.34
r38 7 29 3.02922 $w=2.8e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.225 $Y=2.635
+ $X2=0.182 $Y2=2.72
r39 7 12 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=0.225 $Y=2.635
+ $X2=0.225 $Y2=2.34
r40 2 20 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.34
r41 2 17 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.66
r42 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.485 $X2=0.28 $Y2=2.34
r43 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.485 $X2=0.28 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_1%Y 1 2 7 8 9 24 32 35
r28 29 32 7.40429 $w=6.28e-07 $l=3.9e-07 $layer=LI1_cond $X=0.735 $Y=0.57
+ $X2=1.125 $Y2=0.57
r29 24 25 5.99336 $w=3.78e-07 $l=8e-08 $layer=LI1_cond $X=0.725 $Y=1.565
+ $X2=0.725 $Y2=1.485
r30 17 28 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=0.725 $Y=1.675
+ $X2=0.725 $Y2=1.66
r31 14 29 8.63246 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=0.735 $Y=0.885
+ $X2=0.735 $Y2=0.57
r32 9 35 1.4239 $w=6.28e-07 $l=7.5e-08 $layer=LI1_cond $X=1.145 $Y=0.57 $X2=1.22
+ $Y2=0.57
r33 9 32 0.379707 $w=6.28e-07 $l=2e-08 $layer=LI1_cond $X=1.145 $Y=0.57
+ $X2=1.125 $Y2=0.57
r34 8 21 13.1924 $w=3.78e-07 $l=4.35e-07 $layer=LI1_cond $X=0.725 $Y=1.905
+ $X2=0.725 $Y2=2.34
r35 8 17 6.97531 $w=3.78e-07 $l=2.3e-07 $layer=LI1_cond $X=0.725 $Y=1.905
+ $X2=0.725 $Y2=1.675
r36 7 28 2.82045 $w=3.78e-07 $l=9.3e-08 $layer=LI1_cond $X=0.725 $Y=1.567
+ $X2=0.725 $Y2=1.66
r37 7 24 0.0606549 $w=3.78e-07 $l=2e-09 $layer=LI1_cond $X=0.725 $Y=1.567
+ $X2=0.725 $Y2=1.565
r38 7 25 0.195722 $w=1.68e-07 $l=3e-09 $layer=LI1_cond $X=0.735 $Y=1.482
+ $X2=0.735 $Y2=1.485
r39 7 14 38.9487 $w=1.68e-07 $l=5.97e-07 $layer=LI1_cond $X=0.735 $Y=1.482
+ $X2=0.735 $Y2=0.885
r40 2 28 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=1.66
r41 2 21 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=2.34
r42 1 35 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=1.035
+ $Y=0.235 $X2=1.22 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_1%VGND 1 4 6 8 15 16 24
r16 19 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r17 15 16 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r18 13 16 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r19 13 24 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r20 12 15 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r21 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r22 10 19 4.61546 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.197
+ $Y2=0
r23 10 12 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.69
+ $Y2=0
r24 8 24 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=0 $X2=0.23
+ $Y2=0
r25 4 19 2.98373 $w=3.1e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.197 $Y2=0
r26 4 6 10.9668 $w=3.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.38
r27 1 6 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.235 $X2=0.28 $Y2=0.38
.ends

