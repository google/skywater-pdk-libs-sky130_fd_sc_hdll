* File: sky130_fd_sc_hdll__bufbuf_16.pex.spice
* Created: Wed Sep  2 08:24:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__BUFBUF_16%A 1 3 4 6 7
r23 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r24 4 10 40.1292 $w=4.26e-07 $l=2.36525e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.352 $Y2=1.16
r25 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r26 1 10 44.7281 $w=4.26e-07 $l=3.13449e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.352 $Y2=1.16
r27 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFBUF_16%A_117_297# 1 2 9 11 13 16 18 20 21 23 26
+ 30 34 37 42 45 47 48 49 55
c97 42 0 1.39726e-19 $X=2.06 $Y=1.16
c98 26 0 1.25206e-19 $X=2.45 $Y=0.56
c99 21 0 1.26528e-19 $X=2.425 $Y=1.41
r100 55 56 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.425 $Y=1.217
+ $X2=2.45 $Y2=1.217
r101 52 53 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.93 $Y=1.217
+ $X2=1.955 $Y2=1.217
r102 51 52 64.997 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=1.485 $Y=1.217
+ $X2=1.93 $Y2=1.217
r103 50 51 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.46 $Y=1.217
+ $X2=1.485 $Y2=1.217
r104 47 48 7.27811 $w=3.78e-07 $l=1.85e-07 $layer=LI1_cond $X=0.705 $Y=1.63
+ $X2=0.705 $Y2=1.445
r105 43 55 53.3121 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=2.06 $Y=1.217
+ $X2=2.425 $Y2=1.217
r106 43 53 15.3364 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=2.06 $Y=1.217
+ $X2=1.955 $Y2=1.217
r107 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.06
+ $Y=1.16 $X2=2.06 $Y2=1.16
r108 40 49 1.92922 $w=2e-07 $l=1.18e-07 $layer=LI1_cond $X=0.895 $Y=1.175
+ $X2=0.777 $Y2=1.175
r109 40 42 64.6045 $w=1.98e-07 $l=1.165e-06 $layer=LI1_cond $X=0.895 $Y=1.175
+ $X2=2.06 $Y2=1.175
r110 38 49 4.50812 $w=2.35e-07 $l=1e-07 $layer=LI1_cond $X=0.777 $Y=1.275
+ $X2=0.777 $Y2=1.175
r111 38 48 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=0.777 $Y=1.275
+ $X2=0.777 $Y2=1.445
r112 37 49 4.50812 $w=2.35e-07 $l=1e-07 $layer=LI1_cond $X=0.777 $Y=1.075
+ $X2=0.777 $Y2=1.175
r113 37 45 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=0.777 $Y=1.075
+ $X2=0.777 $Y2=0.905
r114 32 47 0.151637 $w=3.78e-07 $l=5e-09 $layer=LI1_cond $X=0.705 $Y=1.635
+ $X2=0.705 $Y2=1.63
r115 32 34 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.705 $Y=1.635
+ $X2=0.705 $Y2=2.31
r116 28 45 7.42975 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=0.705 $Y=0.715
+ $X2=0.705 $Y2=0.905
r117 28 30 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.705 $Y=0.715
+ $X2=0.705 $Y2=0.4
r118 24 56 21.2229 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.45 $Y=1.025
+ $X2=2.45 $Y2=1.217
r119 24 26 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.45 $Y=1.025
+ $X2=2.45 $Y2=0.56
r120 21 55 16.9318 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.217
r121 21 23 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.985
r122 18 53 16.9318 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.217
r123 18 20 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.985
r124 14 52 21.2229 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=1.217
r125 14 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=0.56
r126 11 51 16.9318 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.217
r127 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.985
r128 7 50 21.2229 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=1.217
r129 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=0.56
r130 2 47 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.63
r131 2 34 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.31
r132 1 30 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFBUF_16%A_225_47# 1 2 3 4 15 17 19 22 24 26 29
+ 31 33 36 38 40 43 45 47 48 50 53 57 61 65 66 67 68 71 75 79 81 84 86 92 95 96
+ 97 110
c214 110 0 1.39726e-19 $X=5.245 $Y=1.217
c215 92 0 1.34672e-19 $X=4.9 $Y=1.16
c216 53 0 1.25206e-19 $X=5.27 $Y=0.56
c217 48 0 1.26528e-19 $X=5.245 $Y=1.41
r218 110 111 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=5.245 $Y=1.217
+ $X2=5.27 $Y2=1.217
r219 107 108 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=4.75 $Y=1.217
+ $X2=4.775 $Y2=1.217
r220 106 107 66.2006 $w=3.24e-07 $l=4.45e-07 $layer=POLY_cond $X=4.305 $Y=1.217
+ $X2=4.75 $Y2=1.217
r221 105 106 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=4.28 $Y=1.217
+ $X2=4.305 $Y2=1.217
r222 104 105 66.2006 $w=3.24e-07 $l=4.45e-07 $layer=POLY_cond $X=3.835 $Y=1.217
+ $X2=4.28 $Y2=1.217
r223 103 104 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=3.81 $Y=1.217
+ $X2=3.835 $Y2=1.217
r224 102 103 66.2006 $w=3.24e-07 $l=4.45e-07 $layer=POLY_cond $X=3.365 $Y=1.217
+ $X2=3.81 $Y2=1.217
r225 101 102 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=3.34 $Y=1.217
+ $X2=3.365 $Y2=1.217
r226 98 99 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=2.87 $Y=1.217
+ $X2=2.895 $Y2=1.217
r227 93 110 51.3241 $w=3.24e-07 $l=3.45e-07 $layer=POLY_cond $X=4.9 $Y=1.217
+ $X2=5.245 $Y2=1.217
r228 93 108 18.5957 $w=3.24e-07 $l=1.25e-07 $layer=POLY_cond $X=4.9 $Y=1.217
+ $X2=4.775 $Y2=1.217
r229 92 93 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=4.9
+ $Y=1.16 $X2=4.9 $Y2=1.16
r230 90 101 50.5802 $w=3.24e-07 $l=3.4e-07 $layer=POLY_cond $X=3 $Y=1.217
+ $X2=3.34 $Y2=1.217
r231 90 99 15.6204 $w=3.24e-07 $l=1.05e-07 $layer=POLY_cond $X=3 $Y=1.217
+ $X2=2.895 $Y2=1.217
r232 89 92 105.364 $w=1.98e-07 $l=1.9e-06 $layer=LI1_cond $X=3 $Y=1.175 $X2=4.9
+ $Y2=1.175
r233 89 90 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3
+ $Y=1.16 $X2=3 $Y2=1.16
r234 87 97 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=1.175
+ $X2=2.66 $Y2=1.175
r235 87 89 14.1409 $w=1.98e-07 $l=2.55e-07 $layer=LI1_cond $X=2.745 $Y=1.175
+ $X2=3 $Y2=1.175
r236 85 97 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.66 $Y=1.275 $X2=2.66
+ $Y2=1.175
r237 85 86 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.66 $Y=1.275
+ $X2=2.66 $Y2=1.445
r238 84 97 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.66 $Y=1.075 $X2=2.66
+ $Y2=1.175
r239 83 84 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.66 $Y=0.905
+ $X2=2.66 $Y2=1.075
r240 82 96 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.355 $Y=1.53
+ $X2=2.165 $Y2=1.53
r241 81 86 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.575 $Y=1.53
+ $X2=2.66 $Y2=1.445
r242 81 82 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.575 $Y=1.53
+ $X2=2.355 $Y2=1.53
r243 80 95 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.355 $Y=0.82
+ $X2=2.165 $Y2=0.82
r244 79 83 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.575 $Y=0.82
+ $X2=2.66 $Y2=0.905
r245 79 80 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.575 $Y=0.82
+ $X2=2.355 $Y2=0.82
r246 75 77 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=2.165 $Y=1.63
+ $X2=2.165 $Y2=2.31
r247 73 96 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=1.615
+ $X2=2.165 $Y2=1.53
r248 73 75 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=2.165 $Y=1.615
+ $X2=2.165 $Y2=1.63
r249 69 95 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=0.735
+ $X2=2.165 $Y2=0.82
r250 69 71 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.165 $Y=0.735
+ $X2=2.165 $Y2=0.4
r251 67 96 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.975 $Y=1.53
+ $X2=2.165 $Y2=1.53
r252 67 68 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.975 $Y=1.53
+ $X2=1.415 $Y2=1.53
r253 65 95 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.975 $Y=0.82
+ $X2=2.165 $Y2=0.82
r254 65 66 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.975 $Y=0.82
+ $X2=1.415 $Y2=0.82
r255 61 63 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.25 $Y=1.63
+ $X2=1.25 $Y2=2.31
r256 59 68 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.25 $Y=1.615
+ $X2=1.415 $Y2=1.53
r257 59 61 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.25 $Y=1.615
+ $X2=1.25 $Y2=1.63
r258 55 66 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.25 $Y=0.735
+ $X2=1.415 $Y2=0.82
r259 55 57 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.25 $Y=0.735
+ $X2=1.25 $Y2=0.4
r260 51 111 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.27 $Y=1.025
+ $X2=5.27 $Y2=1.217
r261 51 53 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.27 $Y=1.025
+ $X2=5.27 $Y2=0.56
r262 48 110 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.217
r263 48 50 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.985
r264 45 108 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.217
r265 45 47 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
r266 41 107 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.75 $Y=1.025
+ $X2=4.75 $Y2=1.217
r267 41 43 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.75 $Y=1.025
+ $X2=4.75 $Y2=0.56
r268 38 106 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.217
r269 38 40 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.985
r270 34 105 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.28 $Y=1.025
+ $X2=4.28 $Y2=1.217
r271 34 36 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.28 $Y=1.025
+ $X2=4.28 $Y2=0.56
r272 31 104 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.217
r273 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.985
r274 27 103 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.81 $Y=1.025
+ $X2=3.81 $Y2=1.217
r275 27 29 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.81 $Y=1.025
+ $X2=3.81 $Y2=0.56
r276 24 102 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.217
r277 24 26 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.985
r278 20 101 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.34 $Y=1.025
+ $X2=3.34 $Y2=1.217
r279 20 22 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.34 $Y=1.025
+ $X2=3.34 $Y2=0.56
r280 17 99 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.217
r281 17 19 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.985
r282 13 98 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.87 $Y=1.025
+ $X2=2.87 $Y2=1.217
r283 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.87 $Y=1.025
+ $X2=2.87 $Y2=0.56
r284 4 77 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.485 $X2=2.19 $Y2=2.31
r285 4 75 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.485 $X2=2.19 $Y2=1.63
r286 3 63 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.25 $Y2=2.31
r287 3 61 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.25 $Y2=1.63
r288 2 71 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=2.005
+ $Y=0.235 $X2=2.19 $Y2=0.4
r289 1 57 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=1.125
+ $Y=0.235 $X2=1.25 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFBUF_16%A_589_47# 1 2 3 4 5 6 21 23 25 28 30 32
+ 35 37 39 42 44 46 49 51 53 56 58 60 63 65 67 70 72 74 77 79 81 84 86 88 91 93
+ 95 98 100 102 105 107 109 112 114 116 119 121 123 124 126 129 133 137 141 142
+ 143 144 147 151 155 157 161 165 169 171 174 176 182 185 186 187 188 189 222
c462 222 0 1.34672e-19 $X=12.765 $Y=1.217
c463 144 0 1.26528e-19 $X=3.295 $Y=1.53
c464 142 0 1.25206e-19 $X=3.295 $Y=0.82
r465 222 223 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=12.765 $Y=1.217
+ $X2=12.79 $Y2=1.217
r466 221 222 70.7937 $w=3.2e-07 $l=4.7e-07 $layer=POLY_cond $X=12.295 $Y=1.217
+ $X2=12.765 $Y2=1.217
r467 218 219 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=11.825 $Y=1.217
+ $X2=12.27 $Y2=1.217
r468 217 218 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=11.8 $Y=1.217
+ $X2=11.825 $Y2=1.217
r469 216 217 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=11.355 $Y=1.217
+ $X2=11.8 $Y2=1.217
r470 215 216 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=11.33 $Y=1.217
+ $X2=11.355 $Y2=1.217
r471 214 215 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=10.885 $Y=1.217
+ $X2=11.33 $Y2=1.217
r472 213 214 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=10.86 $Y=1.217
+ $X2=10.885 $Y2=1.217
r473 212 213 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=10.415 $Y=1.217
+ $X2=10.86 $Y2=1.217
r474 211 212 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=10.39 $Y=1.217
+ $X2=10.415 $Y2=1.217
r475 210 211 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=9.945 $Y=1.217
+ $X2=10.39 $Y2=1.217
r476 209 210 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=9.92 $Y=1.217
+ $X2=9.945 $Y2=1.217
r477 208 209 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=9.475 $Y=1.217
+ $X2=9.92 $Y2=1.217
r478 207 208 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=9.45 $Y=1.217
+ $X2=9.475 $Y2=1.217
r479 206 207 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=9.005 $Y=1.217
+ $X2=9.45 $Y2=1.217
r480 205 206 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=8.98 $Y=1.217
+ $X2=9.005 $Y2=1.217
r481 204 205 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=8.535 $Y=1.217
+ $X2=8.98 $Y2=1.217
r482 203 204 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=8.51 $Y=1.217
+ $X2=8.535 $Y2=1.217
r483 202 203 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=8.065 $Y=1.217
+ $X2=8.51 $Y2=1.217
r484 201 202 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=8.04 $Y=1.217
+ $X2=8.065 $Y2=1.217
r485 200 201 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=7.595 $Y=1.217
+ $X2=8.04 $Y2=1.217
r486 199 200 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=7.57 $Y=1.217
+ $X2=7.595 $Y2=1.217
r487 198 199 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=7.125 $Y=1.217
+ $X2=7.57 $Y2=1.217
r488 197 198 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=7.1 $Y=1.217
+ $X2=7.125 $Y2=1.217
r489 196 197 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=6.655 $Y=1.217
+ $X2=7.1 $Y2=1.217
r490 195 196 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=6.63 $Y=1.217
+ $X2=6.655 $Y2=1.217
r491 194 195 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=6.185 $Y=1.217
+ $X2=6.63 $Y2=1.217
r492 193 194 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=6.16 $Y=1.217
+ $X2=6.185 $Y2=1.217
r493 190 191 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=5.69 $Y=1.217
+ $X2=5.715 $Y2=1.217
r494 183 221 2.25938 $w=3.2e-07 $l=1.5e-08 $layer=POLY_cond $X=12.28 $Y=1.217
+ $X2=12.295 $Y2=1.217
r495 183 219 1.50625 $w=3.2e-07 $l=1e-08 $layer=POLY_cond $X=12.28 $Y=1.217
+ $X2=12.27 $Y2=1.217
r496 182 183 16.1422 $w=1.7e-07 $l=1.53e-06 $layer=licon1_POLY $count=9 $X=12.28
+ $Y=1.16 $X2=12.28 $Y2=1.16
r497 180 193 54.225 $w=3.2e-07 $l=3.6e-07 $layer=POLY_cond $X=5.8 $Y=1.217
+ $X2=6.16 $Y2=1.217
r498 180 191 12.8031 $w=3.2e-07 $l=8.5e-08 $layer=POLY_cond $X=5.8 $Y=1.217
+ $X2=5.715 $Y2=1.217
r499 179 182 359.345 $w=1.98e-07 $l=6.48e-06 $layer=LI1_cond $X=5.8 $Y=1.175
+ $X2=12.28 $Y2=1.175
r500 179 180 16.1422 $w=1.7e-07 $l=1.53e-06 $layer=licon1_POLY $count=9 $X=5.8
+ $Y=1.16 $X2=5.8 $Y2=1.16
r501 177 189 0.866423 $w=2e-07 $l=8.8e-08 $layer=LI1_cond $X=5.565 $Y=1.175
+ $X2=5.477 $Y2=1.175
r502 177 179 13.0318 $w=1.98e-07 $l=2.35e-07 $layer=LI1_cond $X=5.565 $Y=1.175
+ $X2=5.8 $Y2=1.175
r503 175 189 5.7647 $w=1.75e-07 $l=1e-07 $layer=LI1_cond $X=5.477 $Y=1.275
+ $X2=5.477 $Y2=1.175
r504 175 176 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=5.477 $Y=1.275
+ $X2=5.477 $Y2=1.445
r505 174 189 5.7647 $w=1.75e-07 $l=1e-07 $layer=LI1_cond $X=5.477 $Y=1.075
+ $X2=5.477 $Y2=1.175
r506 173 174 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=5.477 $Y=0.905
+ $X2=5.477 $Y2=1.075
r507 172 188 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.175 $Y=1.53
+ $X2=4.985 $Y2=1.53
r508 171 176 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=5.39 $Y=1.53
+ $X2=5.477 $Y2=1.445
r509 171 172 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.39 $Y=1.53
+ $X2=5.175 $Y2=1.53
r510 170 187 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.175 $Y=0.82
+ $X2=4.985 $Y2=0.82
r511 169 173 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=5.39 $Y=0.82
+ $X2=5.477 $Y2=0.905
r512 169 170 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.39 $Y=0.82
+ $X2=5.175 $Y2=0.82
r513 165 167 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=4.985 $Y=1.63
+ $X2=4.985 $Y2=2.31
r514 163 188 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.985 $Y=1.615
+ $X2=4.985 $Y2=1.53
r515 163 165 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=4.985 $Y=1.615
+ $X2=4.985 $Y2=1.63
r516 159 187 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.985 $Y=0.735
+ $X2=4.985 $Y2=0.82
r517 159 161 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.985 $Y=0.735
+ $X2=4.985 $Y2=0.4
r518 158 186 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.235 $Y=1.53
+ $X2=4.045 $Y2=1.53
r519 157 188 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.795 $Y=1.53
+ $X2=4.985 $Y2=1.53
r520 157 158 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.795 $Y=1.53
+ $X2=4.235 $Y2=1.53
r521 156 185 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.235 $Y=0.82
+ $X2=4.045 $Y2=0.82
r522 155 187 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.795 $Y=0.82
+ $X2=4.985 $Y2=0.82
r523 155 156 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.795 $Y=0.82
+ $X2=4.235 $Y2=0.82
r524 151 153 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=4.045 $Y=1.63
+ $X2=4.045 $Y2=2.31
r525 149 186 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=1.615
+ $X2=4.045 $Y2=1.53
r526 149 151 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=4.045 $Y=1.615
+ $X2=4.045 $Y2=1.63
r527 145 185 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=0.735
+ $X2=4.045 $Y2=0.82
r528 145 147 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.045 $Y=0.735
+ $X2=4.045 $Y2=0.4
r529 143 186 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.855 $Y=1.53
+ $X2=4.045 $Y2=1.53
r530 143 144 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.855 $Y=1.53
+ $X2=3.295 $Y2=1.53
r531 141 185 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.855 $Y=0.82
+ $X2=4.045 $Y2=0.82
r532 141 142 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.855 $Y=0.82
+ $X2=3.295 $Y2=0.82
r533 137 139 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=3.105 $Y=1.63
+ $X2=3.105 $Y2=2.31
r534 135 144 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=3.105 $Y=1.615
+ $X2=3.295 $Y2=1.53
r535 135 137 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=3.105 $Y=1.615
+ $X2=3.105 $Y2=1.63
r536 131 142 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=3.105 $Y=0.735
+ $X2=3.295 $Y2=0.82
r537 131 133 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.105 $Y=0.735
+ $X2=3.105 $Y2=0.4
r538 127 223 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=12.79 $Y=1.025
+ $X2=12.79 $Y2=1.217
r539 127 129 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=12.79 $Y=1.025
+ $X2=12.79 $Y2=0.56
r540 124 222 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=12.765 $Y=1.41
+ $X2=12.765 $Y2=1.217
r541 124 126 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.765 $Y=1.41
+ $X2=12.765 $Y2=1.985
r542 121 221 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=12.295 $Y=1.41
+ $X2=12.295 $Y2=1.217
r543 121 123 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.295 $Y=1.41
+ $X2=12.295 $Y2=1.985
r544 117 219 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=12.27 $Y=1.025
+ $X2=12.27 $Y2=1.217
r545 117 119 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=12.27 $Y=1.025
+ $X2=12.27 $Y2=0.56
r546 114 218 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=11.825 $Y=1.41
+ $X2=11.825 $Y2=1.217
r547 114 116 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.825 $Y=1.41
+ $X2=11.825 $Y2=1.985
r548 110 217 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=11.8 $Y=1.025
+ $X2=11.8 $Y2=1.217
r549 110 112 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.8 $Y=1.025
+ $X2=11.8 $Y2=0.56
r550 107 216 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=11.355 $Y=1.41
+ $X2=11.355 $Y2=1.217
r551 107 109 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.355 $Y=1.41
+ $X2=11.355 $Y2=1.985
r552 103 215 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=11.33 $Y=1.025
+ $X2=11.33 $Y2=1.217
r553 103 105 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.33 $Y=1.025
+ $X2=11.33 $Y2=0.56
r554 100 214 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=10.885 $Y=1.41
+ $X2=10.885 $Y2=1.217
r555 100 102 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.885 $Y=1.41
+ $X2=10.885 $Y2=1.985
r556 96 213 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=10.86 $Y=1.025
+ $X2=10.86 $Y2=1.217
r557 96 98 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=10.86 $Y=1.025
+ $X2=10.86 $Y2=0.56
r558 93 212 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=10.415 $Y=1.41
+ $X2=10.415 $Y2=1.217
r559 93 95 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.415 $Y=1.41
+ $X2=10.415 $Y2=1.985
r560 89 211 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=10.39 $Y=1.025
+ $X2=10.39 $Y2=1.217
r561 89 91 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=10.39 $Y=1.025
+ $X2=10.39 $Y2=0.56
r562 86 210 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=9.945 $Y=1.41
+ $X2=9.945 $Y2=1.217
r563 86 88 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.945 $Y=1.41
+ $X2=9.945 $Y2=1.985
r564 82 209 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=9.92 $Y=1.025
+ $X2=9.92 $Y2=1.217
r565 82 84 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.92 $Y=1.025
+ $X2=9.92 $Y2=0.56
r566 79 208 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=9.475 $Y=1.41
+ $X2=9.475 $Y2=1.217
r567 79 81 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.475 $Y=1.41
+ $X2=9.475 $Y2=1.985
r568 75 207 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=9.45 $Y=1.025
+ $X2=9.45 $Y2=1.217
r569 75 77 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.45 $Y=1.025
+ $X2=9.45 $Y2=0.56
r570 72 206 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=9.005 $Y=1.41
+ $X2=9.005 $Y2=1.217
r571 72 74 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.005 $Y=1.41
+ $X2=9.005 $Y2=1.985
r572 68 205 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=8.98 $Y=1.025
+ $X2=8.98 $Y2=1.217
r573 68 70 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.98 $Y=1.025
+ $X2=8.98 $Y2=0.56
r574 65 204 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=8.535 $Y=1.41
+ $X2=8.535 $Y2=1.217
r575 65 67 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.535 $Y=1.41
+ $X2=8.535 $Y2=1.985
r576 61 203 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=8.51 $Y=1.025
+ $X2=8.51 $Y2=1.217
r577 61 63 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.51 $Y=1.025
+ $X2=8.51 $Y2=0.56
r578 58 202 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=8.065 $Y=1.41
+ $X2=8.065 $Y2=1.217
r579 58 60 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.065 $Y=1.41
+ $X2=8.065 $Y2=1.985
r580 54 201 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=8.04 $Y=1.025
+ $X2=8.04 $Y2=1.217
r581 54 56 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.04 $Y=1.025
+ $X2=8.04 $Y2=0.56
r582 51 200 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.595 $Y=1.41
+ $X2=7.595 $Y2=1.217
r583 51 53 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.595 $Y=1.41
+ $X2=7.595 $Y2=1.985
r584 47 199 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.57 $Y=1.025
+ $X2=7.57 $Y2=1.217
r585 47 49 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.57 $Y=1.025
+ $X2=7.57 $Y2=0.56
r586 44 198 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.217
r587 44 46 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.985
r588 40 197 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.1 $Y=1.025
+ $X2=7.1 $Y2=1.217
r589 40 42 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.1 $Y=1.025
+ $X2=7.1 $Y2=0.56
r590 37 196 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.217
r591 37 39 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.985
r592 33 195 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.63 $Y=1.025
+ $X2=6.63 $Y2=1.217
r593 33 35 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.63 $Y=1.025
+ $X2=6.63 $Y2=0.56
r594 30 194 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.217
r595 30 32 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.985
r596 26 193 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.16 $Y=1.025
+ $X2=6.16 $Y2=1.217
r597 26 28 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.16 $Y=1.025
+ $X2=6.16 $Y2=0.56
r598 23 191 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.217
r599 23 25 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.985
r600 19 190 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.69 $Y=1.025
+ $X2=5.69 $Y2=1.217
r601 19 21 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.69 $Y=1.025
+ $X2=5.69 $Y2=0.56
r602 6 167 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=2.31
r603 6 165 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=1.63
r604 5 153 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=2.31
r605 5 151 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=1.63
r606 4 139 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=2.985
+ $Y=1.485 $X2=3.13 $Y2=2.31
r607 4 137 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.985
+ $Y=1.485 $X2=3.13 $Y2=1.63
r608 3 161 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=4.825
+ $Y=0.235 $X2=5.01 $Y2=0.4
r609 2 147 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=3.885
+ $Y=0.235 $X2=4.07 $Y2=0.4
r610 1 133 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=2.945
+ $Y=0.235 $X2=3.13 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFBUF_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 14 43
+ 45 51 55 59 63 67 71 75 79 83 87 91 95 97 99 102 103 105 106 108 109 111 112
+ 114 115 117 118 120 121 123 124 126 127 129 130 132 133 135 136 137 179 188
+ 191
r217 187 188 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r218 184 191 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r219 182 188 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=13.11 $Y2=2.72
r220 181 182 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r221 179 187 3.40825 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=12.915 $Y=2.72
+ $X2=13.127 $Y2=2.72
r222 179 181 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=12.915 $Y=2.72
+ $X2=12.65 $Y2=2.72
r223 178 182 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=12.65 $Y2=2.72
r224 177 178 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r225 175 178 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.73 $Y2=2.72
r226 174 175 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r227 172 175 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.81 $Y2=2.72
r228 171 172 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r229 169 172 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r230 168 169 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r231 166 169 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r232 165 166 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r233 163 166 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r234 162 163 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r235 160 163 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r236 159 160 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r237 157 160 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r238 156 157 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r239 154 157 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r240 153 154 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r241 151 154 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r242 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r243 148 151 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r244 147 148 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r245 145 148 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r246 144 145 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r247 142 145 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r248 141 144 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r249 141 142 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r250 139 184 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r251 139 141 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r252 137 142 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r253 137 191 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r254 135 177 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=11.975 $Y=2.72
+ $X2=11.73 $Y2=2.72
r255 135 136 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.975 $Y=2.72
+ $X2=12.06 $Y2=2.72
r256 134 181 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=12.145 $Y=2.72
+ $X2=12.65 $Y2=2.72
r257 134 136 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.145 $Y=2.72
+ $X2=12.06 $Y2=2.72
r258 132 174 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=11.035 $Y=2.72
+ $X2=10.81 $Y2=2.72
r259 132 133 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.035 $Y=2.72
+ $X2=11.12 $Y2=2.72
r260 131 177 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=11.205 $Y=2.72
+ $X2=11.73 $Y2=2.72
r261 131 133 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.205 $Y=2.72
+ $X2=11.12 $Y2=2.72
r262 129 171 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=10.095 $Y=2.72
+ $X2=9.89 $Y2=2.72
r263 129 130 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.095 $Y=2.72
+ $X2=10.18 $Y2=2.72
r264 128 174 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=10.265 $Y=2.72
+ $X2=10.81 $Y2=2.72
r265 128 130 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.265 $Y=2.72
+ $X2=10.18 $Y2=2.72
r266 126 168 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=9.155 $Y=2.72
+ $X2=8.97 $Y2=2.72
r267 126 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.155 $Y=2.72
+ $X2=9.24 $Y2=2.72
r268 125 171 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=9.325 $Y=2.72
+ $X2=9.89 $Y2=2.72
r269 125 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.325 $Y=2.72
+ $X2=9.24 $Y2=2.72
r270 123 165 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.215 $Y=2.72
+ $X2=8.05 $Y2=2.72
r271 123 124 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.215 $Y=2.72
+ $X2=8.3 $Y2=2.72
r272 122 168 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=8.385 $Y=2.72
+ $X2=8.97 $Y2=2.72
r273 122 124 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.385 $Y=2.72
+ $X2=8.3 $Y2=2.72
r274 120 162 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.275 $Y=2.72
+ $X2=7.13 $Y2=2.72
r275 120 121 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.275 $Y=2.72
+ $X2=7.36 $Y2=2.72
r276 119 165 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=7.445 $Y=2.72
+ $X2=8.05 $Y2=2.72
r277 119 121 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.445 $Y=2.72
+ $X2=7.36 $Y2=2.72
r278 117 159 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.335 $Y=2.72
+ $X2=6.21 $Y2=2.72
r279 117 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.335 $Y=2.72
+ $X2=6.42 $Y2=2.72
r280 116 162 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=6.505 $Y=2.72
+ $X2=7.13 $Y2=2.72
r281 116 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.505 $Y=2.72
+ $X2=6.42 $Y2=2.72
r282 114 156 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=5.395 $Y=2.72
+ $X2=5.29 $Y2=2.72
r283 114 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=2.72
+ $X2=5.48 $Y2=2.72
r284 113 159 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=5.565 $Y=2.72
+ $X2=6.21 $Y2=2.72
r285 113 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=2.72
+ $X2=5.48 $Y2=2.72
r286 111 153 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=2.72
+ $X2=4.37 $Y2=2.72
r287 111 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=2.72
+ $X2=4.54 $Y2=2.72
r288 110 156 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=5.29 $Y2=2.72
r289 110 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=4.54 $Y2=2.72
r290 108 150 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.515 $Y=2.72
+ $X2=3.45 $Y2=2.72
r291 108 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=2.72
+ $X2=3.6 $Y2=2.72
r292 107 153 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=4.37 $Y2=2.72
r293 107 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=3.6 $Y2=2.72
r294 105 147 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.575 $Y=2.72
+ $X2=2.53 $Y2=2.72
r295 105 106 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.575 $Y=2.72
+ $X2=2.66 $Y2=2.72
r296 104 150 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.745 $Y=2.72
+ $X2=3.45 $Y2=2.72
r297 104 106 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=2.72
+ $X2=2.66 $Y2=2.72
r298 102 144 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.635 $Y=2.72
+ $X2=1.61 $Y2=2.72
r299 102 103 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=2.72
+ $X2=1.72 $Y2=2.72
r300 101 147 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=2.53 $Y2=2.72
r301 101 103 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=1.72 $Y2=2.72
r302 97 187 3.40825 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=13 $Y=2.635
+ $X2=13.127 $Y2=2.72
r303 97 99 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=13 $Y=2.635 $X2=13
+ $Y2=2
r304 93 136 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.06 $Y=2.635
+ $X2=12.06 $Y2=2.72
r305 93 95 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=12.06 $Y=2.635
+ $X2=12.06 $Y2=2
r306 89 133 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.12 $Y=2.635
+ $X2=11.12 $Y2=2.72
r307 89 91 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=11.12 $Y=2.635
+ $X2=11.12 $Y2=2
r308 85 130 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.18 $Y=2.635
+ $X2=10.18 $Y2=2.72
r309 85 87 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=10.18 $Y=2.635
+ $X2=10.18 $Y2=2
r310 81 127 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.24 $Y=2.635
+ $X2=9.24 $Y2=2.72
r311 81 83 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=9.24 $Y=2.635
+ $X2=9.24 $Y2=2
r312 77 124 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.3 $Y=2.635
+ $X2=8.3 $Y2=2.72
r313 77 79 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.3 $Y=2.635
+ $X2=8.3 $Y2=2
r314 73 121 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=2.635
+ $X2=7.36 $Y2=2.72
r315 73 75 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.36 $Y=2.635
+ $X2=7.36 $Y2=2
r316 69 118 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=2.72
r317 69 71 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=2
r318 65 115 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2.72
r319 65 67 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2
r320 61 112 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=2.635
+ $X2=4.54 $Y2=2.72
r321 61 63 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.54 $Y=2.635
+ $X2=4.54 $Y2=2
r322 57 109 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=2.635
+ $X2=3.6 $Y2=2.72
r323 57 59 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.6 $Y=2.635
+ $X2=3.6 $Y2=2
r324 53 106 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=2.635
+ $X2=2.66 $Y2=2.72
r325 53 55 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.66 $Y=2.635
+ $X2=2.66 $Y2=2
r326 49 103 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=2.635
+ $X2=1.72 $Y2=2.72
r327 49 51 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.72 $Y=2.635
+ $X2=1.72 $Y2=2
r328 45 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r329 43 184 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.172 $Y2=2.72
r330 43 48 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r331 14 99 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=12.855
+ $Y=1.485 $X2=13 $Y2=2
r332 13 95 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=11.915
+ $Y=1.485 $X2=12.06 $Y2=2
r333 12 91 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=10.975
+ $Y=1.485 $X2=11.12 $Y2=2
r334 11 87 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=10.035
+ $Y=1.485 $X2=10.18 $Y2=2
r335 10 83 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=9.095
+ $Y=1.485 $X2=9.24 $Y2=2
r336 9 79 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=8.155
+ $Y=1.485 $X2=8.3 $Y2=2
r337 8 75 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=7.215
+ $Y=1.485 $X2=7.36 $Y2=2
r338 7 71 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.275
+ $Y=1.485 $X2=6.42 $Y2=2
r339 6 67 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=2
r340 5 63 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.395
+ $Y=1.485 $X2=4.54 $Y2=2
r341 4 59 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.455
+ $Y=1.485 $X2=3.6 $Y2=2
r342 3 55 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.515
+ $Y=1.485 $X2=2.66 $Y2=2
r343 2 51 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.575
+ $Y=1.485 $X2=1.72 $Y2=2
r344 1 48 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r345 1 45 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFBUF_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 49 50 53 57 58 59 60 61 62 65 69 71 73 74 77 81 83 87 91 95 97 101 105 109 111
+ 115 119 123 125 129 133 137 139 143 147 151 153 159 160 163 164 165 166 167
+ 168 169 170 171 172 173 174 176 177
c363 60 0 1.26528e-19 $X=6.115 $Y=1.53
c364 58 0 1.25206e-19 $X=6.115 $Y=0.82
r365 176 177 8.04866 $w=4.68e-07 $l=2.55e-07 $layer=LI1_cond $X=13.07 $Y=1.19
+ $X2=13.07 $Y2=1.445
r366 175 176 10.9482 $w=2.98e-07 $l=2.85e-07 $layer=LI1_cond $X=13.07 $Y=0.905
+ $X2=13.07 $Y2=1.19
r367 154 174 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=12.695 $Y=1.53
+ $X2=12.505 $Y2=1.53
r368 153 177 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=12.92 $Y=1.53
+ $X2=13.07 $Y2=1.53
r369 153 154 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=12.92 $Y=1.53
+ $X2=12.695 $Y2=1.53
r370 152 173 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=12.695 $Y=0.82
+ $X2=12.505 $Y2=0.82
r371 151 175 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=12.92 $Y=0.82
+ $X2=13.07 $Y2=0.905
r372 151 152 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=12.92 $Y=0.82
+ $X2=12.695 $Y2=0.82
r373 147 149 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=12.505 $Y=1.63
+ $X2=12.505 $Y2=2.31
r374 145 174 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=12.505 $Y=1.615
+ $X2=12.505 $Y2=1.53
r375 145 147 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=12.505 $Y=1.615
+ $X2=12.505 $Y2=1.63
r376 141 173 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=12.505 $Y=0.735
+ $X2=12.505 $Y2=0.82
r377 141 143 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=12.505 $Y=0.735
+ $X2=12.505 $Y2=0.4
r378 140 172 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.755 $Y=1.53
+ $X2=11.565 $Y2=1.53
r379 139 174 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=12.315 $Y=1.53
+ $X2=12.505 $Y2=1.53
r380 139 140 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=12.315 $Y=1.53
+ $X2=11.755 $Y2=1.53
r381 138 171 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.755 $Y=0.82
+ $X2=11.565 $Y2=0.82
r382 137 173 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=12.315 $Y=0.82
+ $X2=12.505 $Y2=0.82
r383 137 138 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=12.315 $Y=0.82
+ $X2=11.755 $Y2=0.82
r384 133 135 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=11.565 $Y=1.63
+ $X2=11.565 $Y2=2.31
r385 131 172 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=11.565 $Y=1.615
+ $X2=11.565 $Y2=1.53
r386 131 133 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=11.565 $Y=1.615
+ $X2=11.565 $Y2=1.63
r387 127 171 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=11.565 $Y=0.735
+ $X2=11.565 $Y2=0.82
r388 127 129 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=11.565 $Y=0.735
+ $X2=11.565 $Y2=0.4
r389 126 170 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.815 $Y=1.53
+ $X2=10.625 $Y2=1.53
r390 125 172 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.375 $Y=1.53
+ $X2=11.565 $Y2=1.53
r391 125 126 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=11.375 $Y=1.53
+ $X2=10.815 $Y2=1.53
r392 124 169 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.815 $Y=0.82
+ $X2=10.625 $Y2=0.82
r393 123 171 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.375 $Y=0.82
+ $X2=11.565 $Y2=0.82
r394 123 124 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=11.375 $Y=0.82
+ $X2=10.815 $Y2=0.82
r395 119 121 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=10.625 $Y=1.63
+ $X2=10.625 $Y2=2.31
r396 117 170 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=10.625 $Y=1.615
+ $X2=10.625 $Y2=1.53
r397 117 119 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=10.625 $Y=1.615
+ $X2=10.625 $Y2=1.63
r398 113 169 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=10.625 $Y=0.735
+ $X2=10.625 $Y2=0.82
r399 113 115 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=10.625 $Y=0.735
+ $X2=10.625 $Y2=0.4
r400 112 168 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.875 $Y=1.53
+ $X2=9.685 $Y2=1.53
r401 111 170 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.435 $Y=1.53
+ $X2=10.625 $Y2=1.53
r402 111 112 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=10.435 $Y=1.53
+ $X2=9.875 $Y2=1.53
r403 110 167 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.875 $Y=0.82
+ $X2=9.685 $Y2=0.82
r404 109 169 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.435 $Y=0.82
+ $X2=10.625 $Y2=0.82
r405 109 110 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=10.435 $Y=0.82
+ $X2=9.875 $Y2=0.82
r406 105 107 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=9.685 $Y=1.63
+ $X2=9.685 $Y2=2.31
r407 103 168 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.685 $Y=1.615
+ $X2=9.685 $Y2=1.53
r408 103 105 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=9.685 $Y=1.615
+ $X2=9.685 $Y2=1.63
r409 99 167 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.685 $Y=0.735
+ $X2=9.685 $Y2=0.82
r410 99 101 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=9.685 $Y=0.735
+ $X2=9.685 $Y2=0.4
r411 98 166 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.935 $Y=1.53
+ $X2=8.745 $Y2=1.53
r412 97 168 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.495 $Y=1.53
+ $X2=9.685 $Y2=1.53
r413 97 98 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=9.495 $Y=1.53
+ $X2=8.935 $Y2=1.53
r414 96 165 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.935 $Y=0.82
+ $X2=8.745 $Y2=0.82
r415 95 167 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.495 $Y=0.82
+ $X2=9.685 $Y2=0.82
r416 95 96 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=9.495 $Y=0.82
+ $X2=8.935 $Y2=0.82
r417 91 93 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=8.745 $Y=1.63
+ $X2=8.745 $Y2=2.31
r418 89 166 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.745 $Y=1.615
+ $X2=8.745 $Y2=1.53
r419 89 91 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=8.745 $Y=1.615
+ $X2=8.745 $Y2=1.63
r420 85 165 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.745 $Y=0.735
+ $X2=8.745 $Y2=0.82
r421 85 87 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=8.745 $Y=0.735
+ $X2=8.745 $Y2=0.4
r422 84 164 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.995 $Y=1.53
+ $X2=7.805 $Y2=1.53
r423 83 166 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.555 $Y=1.53
+ $X2=8.745 $Y2=1.53
r424 83 84 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.555 $Y=1.53
+ $X2=7.995 $Y2=1.53
r425 82 163 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.995 $Y=0.82
+ $X2=7.805 $Y2=0.82
r426 81 165 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.555 $Y=0.82
+ $X2=8.745 $Y2=0.82
r427 81 82 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.555 $Y=0.82
+ $X2=7.995 $Y2=0.82
r428 77 79 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=7.805 $Y=1.63
+ $X2=7.805 $Y2=2.31
r429 75 164 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.805 $Y=1.615
+ $X2=7.805 $Y2=1.53
r430 75 77 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=7.805 $Y=1.615
+ $X2=7.805 $Y2=1.63
r431 74 163 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.805 $Y=0.735
+ $X2=7.805 $Y2=0.82
r432 73 162 1.60526 $w=3.8e-07 $l=5e-08 $layer=LI1_cond $X=7.805 $Y=0.45
+ $X2=7.805 $Y2=0.4
r433 73 74 8.64332 $w=3.78e-07 $l=2.85e-07 $layer=LI1_cond $X=7.805 $Y=0.45
+ $X2=7.805 $Y2=0.735
r434 72 160 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.055 $Y=1.53
+ $X2=6.865 $Y2=1.53
r435 71 164 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.615 $Y=1.53
+ $X2=7.805 $Y2=1.53
r436 71 72 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.615 $Y=1.53
+ $X2=7.055 $Y2=1.53
r437 70 159 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.055 $Y=0.82
+ $X2=6.865 $Y2=0.82
r438 69 163 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.615 $Y=0.82
+ $X2=7.805 $Y2=0.82
r439 69 70 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.615 $Y=0.82
+ $X2=7.055 $Y2=0.82
r440 65 67 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=6.865 $Y=1.63
+ $X2=6.865 $Y2=2.31
r441 63 160 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.865 $Y=1.615
+ $X2=6.865 $Y2=1.53
r442 63 65 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=6.865 $Y=1.615
+ $X2=6.865 $Y2=1.63
r443 62 159 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.865 $Y=0.735
+ $X2=6.865 $Y2=0.82
r444 61 158 1.60526 $w=3.8e-07 $l=5e-08 $layer=LI1_cond $X=6.865 $Y=0.45
+ $X2=6.865 $Y2=0.4
r445 61 62 8.64332 $w=3.78e-07 $l=2.85e-07 $layer=LI1_cond $X=6.865 $Y=0.45
+ $X2=6.865 $Y2=0.735
r446 59 160 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.675 $Y=1.53
+ $X2=6.865 $Y2=1.53
r447 59 60 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.675 $Y=1.53
+ $X2=6.115 $Y2=1.53
r448 57 159 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.675 $Y=0.82
+ $X2=6.865 $Y2=0.82
r449 57 58 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.675 $Y=0.82
+ $X2=6.115 $Y2=0.82
r450 53 55 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=5.925 $Y=1.63
+ $X2=5.925 $Y2=2.31
r451 51 60 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=5.925 $Y=1.615
+ $X2=6.115 $Y2=1.53
r452 51 53 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=5.925 $Y=1.615
+ $X2=5.925 $Y2=1.63
r453 50 58 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=5.925 $Y=0.735
+ $X2=6.115 $Y2=0.82
r454 49 156 1.60526 $w=3.8e-07 $l=5e-08 $layer=LI1_cond $X=5.925 $Y=0.45
+ $X2=5.925 $Y2=0.4
r455 49 50 8.64332 $w=3.78e-07 $l=2.85e-07 $layer=LI1_cond $X=5.925 $Y=0.45
+ $X2=5.925 $Y2=0.735
r456 16 149 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=12.385
+ $Y=1.485 $X2=12.53 $Y2=2.31
r457 16 147 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=12.385
+ $Y=1.485 $X2=12.53 $Y2=1.63
r458 15 135 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=11.445
+ $Y=1.485 $X2=11.59 $Y2=2.31
r459 15 133 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=11.445
+ $Y=1.485 $X2=11.59 $Y2=1.63
r460 14 121 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=10.505
+ $Y=1.485 $X2=10.65 $Y2=2.31
r461 14 119 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.505
+ $Y=1.485 $X2=10.65 $Y2=1.63
r462 13 107 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=9.565
+ $Y=1.485 $X2=9.71 $Y2=2.31
r463 13 105 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=9.565
+ $Y=1.485 $X2=9.71 $Y2=1.63
r464 12 93 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=8.625
+ $Y=1.485 $X2=8.77 $Y2=2.31
r465 12 91 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=8.625
+ $Y=1.485 $X2=8.77 $Y2=1.63
r466 11 79 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=7.685
+ $Y=1.485 $X2=7.83 $Y2=2.31
r467 11 77 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.685
+ $Y=1.485 $X2=7.83 $Y2=1.63
r468 10 67 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=2.31
r469 10 65 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=1.63
r470 9 55 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=2.31
r471 9 53 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=1.63
r472 8 143 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=12.345
+ $Y=0.235 $X2=12.53 $Y2=0.4
r473 7 129 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=11.405
+ $Y=0.235 $X2=11.59 $Y2=0.4
r474 6 115 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=10.465
+ $Y=0.235 $X2=10.65 $Y2=0.4
r475 5 101 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=9.525
+ $Y=0.235 $X2=9.71 $Y2=0.4
r476 4 87 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=8.585
+ $Y=0.235 $X2=8.77 $Y2=0.4
r477 3 162 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=7.645
+ $Y=0.235 $X2=7.83 $Y2=0.4
r478 2 158 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=6.705
+ $Y=0.235 $X2=6.89 $Y2=0.4
r479 1 156 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=5.765
+ $Y=0.235 $X2=5.95 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFBUF_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 14 43
+ 45 49 53 57 61 65 69 73 77 81 85 89 93 95 97 100 101 103 104 106 107 109 110
+ 112 113 115 116 118 119 121 122 124 125 127 128 130 131 133 134 135 177 186
+ 189
r241 185 186 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r242 182 189 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r243 180 186 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.11 $Y2=0
r244 179 180 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r245 177 185 3.40825 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=12.915 $Y=0
+ $X2=13.127 $Y2=0
r246 177 179 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=12.915 $Y=0
+ $X2=12.65 $Y2=0
r247 176 180 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.65 $Y2=0
r248 175 176 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r249 173 176 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.73 $Y2=0
r250 172 173 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r251 170 173 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.81 $Y2=0
r252 169 170 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r253 167 170 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.89 $Y2=0
r254 166 167 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r255 164 167 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.97 $Y2=0
r256 163 164 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r257 161 164 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r258 160 161 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r259 158 161 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.13 $Y2=0
r260 157 158 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r261 155 158 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.21 $Y2=0
r262 154 155 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r263 152 155 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.29 $Y2=0
r264 151 152 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r265 149 152 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.37 $Y2=0
r266 148 149 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r267 146 149 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.45 $Y2=0
r268 145 146 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r269 143 146 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.53 $Y2=0
r270 142 143 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r271 140 143 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.61 $Y2=0
r272 139 142 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0
+ $X2=1.61 $Y2=0
r273 139 140 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r274 137 182 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r275 137 139 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.69 $Y2=0
r276 135 140 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r277 135 189 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r278 133 175 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=11.975 $Y=0
+ $X2=11.73 $Y2=0
r279 133 134 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.975 $Y=0
+ $X2=12.06 $Y2=0
r280 132 179 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=12.145 $Y=0
+ $X2=12.65 $Y2=0
r281 132 134 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.145 $Y=0
+ $X2=12.06 $Y2=0
r282 130 172 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=11.035 $Y=0
+ $X2=10.81 $Y2=0
r283 130 131 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.035 $Y=0
+ $X2=11.12 $Y2=0
r284 129 175 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=11.205 $Y=0
+ $X2=11.73 $Y2=0
r285 129 131 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.205 $Y=0
+ $X2=11.12 $Y2=0
r286 127 169 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=10.095 $Y=0
+ $X2=9.89 $Y2=0
r287 127 128 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.095 $Y=0
+ $X2=10.18 $Y2=0
r288 126 172 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=10.265 $Y=0
+ $X2=10.81 $Y2=0
r289 126 128 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.265 $Y=0
+ $X2=10.18 $Y2=0
r290 124 166 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=9.155 $Y=0
+ $X2=8.97 $Y2=0
r291 124 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.155 $Y=0
+ $X2=9.24 $Y2=0
r292 123 169 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=9.325 $Y=0
+ $X2=9.89 $Y2=0
r293 123 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.325 $Y=0
+ $X2=9.24 $Y2=0
r294 121 163 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.215 $Y=0
+ $X2=8.05 $Y2=0
r295 121 122 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.215 $Y=0 $X2=8.3
+ $Y2=0
r296 120 166 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=8.385 $Y=0
+ $X2=8.97 $Y2=0
r297 120 122 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.385 $Y=0 $X2=8.3
+ $Y2=0
r298 118 160 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.275 $Y=0
+ $X2=7.13 $Y2=0
r299 118 119 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.275 $Y=0
+ $X2=7.36 $Y2=0
r300 117 163 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=7.445 $Y=0
+ $X2=8.05 $Y2=0
r301 117 119 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.445 $Y=0
+ $X2=7.36 $Y2=0
r302 115 157 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.335 $Y=0
+ $X2=6.21 $Y2=0
r303 115 116 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.335 $Y=0
+ $X2=6.42 $Y2=0
r304 114 160 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=6.505 $Y=0
+ $X2=7.13 $Y2=0
r305 114 116 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.505 $Y=0
+ $X2=6.42 $Y2=0
r306 112 154 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=5.395 $Y=0
+ $X2=5.29 $Y2=0
r307 112 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=0
+ $X2=5.48 $Y2=0
r308 111 157 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=5.565 $Y=0
+ $X2=6.21 $Y2=0
r309 111 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=0
+ $X2=5.48 $Y2=0
r310 109 151 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=0
+ $X2=4.37 $Y2=0
r311 109 110 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=0
+ $X2=4.54 $Y2=0
r312 108 154 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.625 $Y=0
+ $X2=5.29 $Y2=0
r313 108 110 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=0
+ $X2=4.54 $Y2=0
r314 106 148 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.515 $Y=0
+ $X2=3.45 $Y2=0
r315 106 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=0 $X2=3.6
+ $Y2=0
r316 105 151 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.685 $Y=0
+ $X2=4.37 $Y2=0
r317 105 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.6
+ $Y2=0
r318 103 145 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.575 $Y=0
+ $X2=2.53 $Y2=0
r319 103 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.575 $Y=0
+ $X2=2.66 $Y2=0
r320 102 148 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.745 $Y=0
+ $X2=3.45 $Y2=0
r321 102 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=0
+ $X2=2.66 $Y2=0
r322 100 142 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.635 $Y=0
+ $X2=1.61 $Y2=0
r323 100 101 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=0
+ $X2=1.72 $Y2=0
r324 99 145 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.805 $Y=0
+ $X2=2.53 $Y2=0
r325 99 101 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.805 $Y=0 $X2=1.72
+ $Y2=0
r326 95 185 3.40825 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=13 $Y=0.085
+ $X2=13.127 $Y2=0
r327 95 97 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=13 $Y=0.085 $X2=13
+ $Y2=0.4
r328 91 134 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.06 $Y=0.085
+ $X2=12.06 $Y2=0
r329 91 93 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.06 $Y=0.085
+ $X2=12.06 $Y2=0.4
r330 87 131 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.12 $Y=0.085
+ $X2=11.12 $Y2=0
r331 87 89 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=11.12 $Y=0.085
+ $X2=11.12 $Y2=0.4
r332 83 128 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.18 $Y=0.085
+ $X2=10.18 $Y2=0
r333 83 85 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.18 $Y=0.085
+ $X2=10.18 $Y2=0.4
r334 79 125 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.24 $Y=0.085
+ $X2=9.24 $Y2=0
r335 79 81 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.24 $Y=0.085
+ $X2=9.24 $Y2=0.4
r336 75 122 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.3 $Y=0.085
+ $X2=8.3 $Y2=0
r337 75 77 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.3 $Y=0.085
+ $X2=8.3 $Y2=0.4
r338 71 119 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0
r339 71 73 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0.4
r340 67 116 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0
r341 67 69 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0.4
r342 63 113 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0
r343 63 65 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.4
r344 59 110 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0
r345 59 61 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0.4
r346 55 107 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=0.085
+ $X2=3.6 $Y2=0
r347 55 57 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.6 $Y=0.085
+ $X2=3.6 $Y2=0.4
r348 51 104 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=0.085
+ $X2=2.66 $Y2=0
r349 51 53 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.66 $Y=0.085
+ $X2=2.66 $Y2=0.4
r350 47 101 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=0.085
+ $X2=1.72 $Y2=0
r351 47 49 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.72 $Y=0.085
+ $X2=1.72 $Y2=0.4
r352 43 182 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r353 43 45 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.4
r354 14 97 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=12.865
+ $Y=0.235 $X2=13 $Y2=0.4
r355 13 93 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=11.875
+ $Y=0.235 $X2=12.06 $Y2=0.4
r356 12 89 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=10.935
+ $Y=0.235 $X2=11.12 $Y2=0.4
r357 11 85 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=9.995
+ $Y=0.235 $X2=10.18 $Y2=0.4
r358 10 81 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=9.055
+ $Y=0.235 $X2=9.24 $Y2=0.4
r359 9 77 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=8.115
+ $Y=0.235 $X2=8.3 $Y2=0.4
r360 8 73 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=7.175
+ $Y=0.235 $X2=7.36 $Y2=0.4
r361 7 69 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=6.235
+ $Y=0.235 $X2=6.42 $Y2=0.4
r362 6 65 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.345
+ $Y=0.235 $X2=5.48 $Y2=0.4
r363 5 61 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=4.355
+ $Y=0.235 $X2=4.54 $Y2=0.4
r364 4 57 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.235 $X2=3.6 $Y2=0.4
r365 3 53 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.525
+ $Y=0.235 $X2=2.66 $Y2=0.4
r366 2 49 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.72 $Y2=0.4
r367 1 45 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

