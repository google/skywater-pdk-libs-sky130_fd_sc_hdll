* File: sky130_fd_sc_hdll__xor3_2.pxi.spice
* Created: Thu Aug 27 19:30:14 2020
* 
x_PM_SKY130_FD_SC_HDLL__XOR3_2%A_81_21# N_A_81_21#_M1002_d N_A_81_21#_M1013_d
+ N_A_81_21#_c_165_n N_A_81_21#_M1001_g N_A_81_21#_c_172_n N_A_81_21#_M1007_g
+ N_A_81_21#_c_173_n N_A_81_21#_M1022_g N_A_81_21#_c_166_n N_A_81_21#_M1016_g
+ N_A_81_21#_c_167_n N_A_81_21#_c_175_n N_A_81_21#_c_182_p N_A_81_21#_c_187_p
+ N_A_81_21#_c_218_p N_A_81_21#_c_168_n N_A_81_21#_c_176_n N_A_81_21#_c_169_n
+ N_A_81_21#_c_177_n N_A_81_21#_c_178_n N_A_81_21#_c_192_p N_A_81_21#_c_170_n
+ N_A_81_21#_c_171_n PM_SKY130_FD_SC_HDLL__XOR3_2%A_81_21#
x_PM_SKY130_FD_SC_HDLL__XOR3_2%C N_C_c_291_n N_C_M1008_g N_C_M1012_g N_C_c_292_n
+ N_C_c_293_n N_C_M1013_g N_C_c_294_n N_C_M1002_g N_C_c_295_n C N_C_c_296_n
+ PM_SKY130_FD_SC_HDLL__XOR3_2%C
x_PM_SKY130_FD_SC_HDLL__XOR3_2%A_335_93# N_A_335_93#_M1008_d N_A_335_93#_M1012_d
+ N_A_335_93#_c_356_n N_A_335_93#_M1003_g N_A_335_93#_c_357_n
+ N_A_335_93#_M1019_g N_A_335_93#_c_372_n N_A_335_93#_c_358_n
+ N_A_335_93#_c_362_n N_A_335_93#_c_363_n N_A_335_93#_c_364_n
+ N_A_335_93#_c_359_n PM_SKY130_FD_SC_HDLL__XOR3_2%A_335_93#
x_PM_SKY130_FD_SC_HDLL__XOR3_2%A_934_297# N_A_934_297#_M1018_d
+ N_A_934_297#_M1004_d N_A_934_297#_c_445_n N_A_934_297#_M1017_g
+ N_A_934_297#_M1011_g N_A_934_297#_c_432_n N_A_934_297#_c_433_n
+ N_A_934_297#_c_447_n N_A_934_297#_M1010_g N_A_934_297#_c_434_n
+ N_A_934_297#_M1015_g N_A_934_297#_c_435_n N_A_934_297#_c_436_n
+ N_A_934_297#_c_450_n N_A_934_297#_c_437_n N_A_934_297#_c_438_n
+ N_A_934_297#_c_454_p N_A_934_297#_c_439_n N_A_934_297#_c_440_n
+ N_A_934_297#_c_441_n N_A_934_297#_c_442_n N_A_934_297#_c_443_n
+ N_A_934_297#_c_444_n PM_SKY130_FD_SC_HDLL__XOR3_2%A_934_297#
x_PM_SKY130_FD_SC_HDLL__XOR3_2%B N_B_c_619_n N_B_M1004_g N_B_M1018_g N_B_c_612_n
+ N_B_c_613_n N_B_M1021_g N_B_M1009_g N_B_c_622_n N_B_c_623_n N_B_M1005_g
+ N_B_c_624_n N_B_c_625_n N_B_M1014_g N_B_c_615_n B N_B_c_616_n N_B_c_617_n
+ N_B_c_618_n N_B_c_631_n PM_SKY130_FD_SC_HDLL__XOR3_2%B
x_PM_SKY130_FD_SC_HDLL__XOR3_2%A N_A_c_746_n N_A_M1000_g N_A_c_747_n N_A_M1006_g
+ A A PM_SKY130_FD_SC_HDLL__XOR3_2%A
x_PM_SKY130_FD_SC_HDLL__XOR3_2%A_1050_365# N_A_1050_365#_M1009_s
+ N_A_1050_365#_M1015_d N_A_1050_365#_M1021_s N_A_1050_365#_M1010_d
+ N_A_1050_365#_c_784_n N_A_1050_365#_M1020_g N_A_1050_365#_c_785_n
+ N_A_1050_365#_M1023_g N_A_1050_365#_c_786_n N_A_1050_365#_c_794_n
+ N_A_1050_365#_c_787_n N_A_1050_365#_c_788_n N_A_1050_365#_c_789_n
+ N_A_1050_365#_c_796_n N_A_1050_365#_c_806_n N_A_1050_365#_c_790_n
+ N_A_1050_365#_c_791_n N_A_1050_365#_c_819_n N_A_1050_365#_c_820_n
+ PM_SKY130_FD_SC_HDLL__XOR3_2%A_1050_365#
x_PM_SKY130_FD_SC_HDLL__XOR3_2%VPWR N_VPWR_M1007_s N_VPWR_M1022_s N_VPWR_M1004_s
+ N_VPWR_M1000_d N_VPWR_c_915_n N_VPWR_c_916_n N_VPWR_c_917_n N_VPWR_c_918_n
+ N_VPWR_c_919_n N_VPWR_c_920_n N_VPWR_c_921_n VPWR N_VPWR_c_922_n
+ N_VPWR_c_923_n N_VPWR_c_914_n N_VPWR_c_925_n N_VPWR_c_926_n
+ PM_SKY130_FD_SC_HDLL__XOR3_2%VPWR
x_PM_SKY130_FD_SC_HDLL__XOR3_2%X N_X_M1001_d N_X_M1007_d N_X_c_1025_n
+ N_X_c_1021_n N_X_c_1031_n X N_X_c_1023_n N_X_c_1022_n
+ PM_SKY130_FD_SC_HDLL__XOR3_2%X
x_PM_SKY130_FD_SC_HDLL__XOR3_2%A_465_325# N_A_465_325#_M1019_d
+ N_A_465_325#_M1005_d N_A_465_325#_M1013_s N_A_465_325#_M1021_d
+ N_A_465_325#_c_1068_n N_A_465_325#_c_1088_n N_A_465_325#_c_1066_n
+ N_A_465_325#_c_1070_n N_A_465_325#_c_1105_n N_A_465_325#_c_1071_n
+ N_A_465_325#_c_1067_n N_A_465_325#_c_1199_p N_A_465_325#_c_1118_n
+ N_A_465_325#_c_1119_n N_A_465_325#_c_1140_n N_A_465_325#_c_1073_n
+ N_A_465_325#_c_1074_n N_A_465_325#_c_1075_n N_A_465_325#_c_1076_n
+ PM_SKY130_FD_SC_HDLL__XOR3_2%A_465_325#
x_PM_SKY130_FD_SC_HDLL__XOR3_2%A_483_49# N_A_483_49#_M1002_s N_A_483_49#_M1009_d
+ N_A_483_49#_M1003_d N_A_483_49#_M1014_d N_A_483_49#_c_1213_n
+ N_A_483_49#_c_1237_n N_A_483_49#_c_1214_n N_A_483_49#_c_1238_n
+ N_A_483_49#_c_1220_n N_A_483_49#_c_1221_n N_A_483_49#_c_1222_n
+ N_A_483_49#_c_1215_n N_A_483_49#_c_1216_n N_A_483_49#_c_1224_n
+ N_A_483_49#_c_1225_n N_A_483_49#_c_1226_n N_A_483_49#_c_1227_n
+ N_A_483_49#_c_1217_n N_A_483_49#_c_1229_n N_A_483_49#_c_1274_n
+ N_A_483_49#_c_1230_n N_A_483_49#_c_1218_n N_A_483_49#_c_1231_n
+ N_A_483_49#_c_1219_n N_A_483_49#_c_1232_n
+ PM_SKY130_FD_SC_HDLL__XOR3_2%A_483_49#
x_PM_SKY130_FD_SC_HDLL__XOR3_2%A_1335_297# N_A_1335_297#_M1011_d
+ N_A_1335_297#_M1023_d N_A_1335_297#_M1017_d N_A_1335_297#_M1020_d
+ N_A_1335_297#_c_1400_n N_A_1335_297#_c_1412_n N_A_1335_297#_c_1404_n
+ N_A_1335_297#_c_1401_n N_A_1335_297#_c_1413_n N_A_1335_297#_c_1406_n
+ N_A_1335_297#_c_1402_n PM_SKY130_FD_SC_HDLL__XOR3_2%A_1335_297#
x_PM_SKY130_FD_SC_HDLL__XOR3_2%VGND N_VGND_M1001_s N_VGND_M1016_s N_VGND_M1018_s
+ N_VGND_M1006_d N_VGND_c_1466_n N_VGND_c_1467_n N_VGND_c_1468_n N_VGND_c_1469_n
+ N_VGND_c_1470_n N_VGND_c_1471_n N_VGND_c_1472_n N_VGND_c_1473_n
+ N_VGND_c_1474_n N_VGND_c_1475_n VGND N_VGND_c_1476_n N_VGND_c_1477_n
+ N_VGND_c_1478_n PM_SKY130_FD_SC_HDLL__XOR3_2%VGND
cc_1 VNB N_A_81_21#_c_165_n 0.0192601f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.995
cc_2 VNB N_A_81_21#_c_166_n 0.0200609f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=0.995
cc_3 VNB N_A_81_21#_c_167_n 0.00256933f $X=-0.19 $Y=-0.24 $X2=1.21 $Y2=1.325
cc_4 VNB N_A_81_21#_c_168_n 0.00138296f $X=-0.19 $Y=-0.24 $X2=1.635 $Y2=0.695
cc_5 VNB N_A_81_21#_c_169_n 0.00282518f $X=-0.19 $Y=-0.24 $X2=1.745 $Y2=0.34
cc_6 VNB N_A_81_21#_c_170_n 0.0162334f $X=-0.19 $Y=-0.24 $X2=2.785 $Y2=0.355
cc_7 VNB N_A_81_21#_c_171_n 0.0565738f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=1.202
cc_8 VNB N_C_c_291_n 0.0197204f $X=-0.19 $Y=-0.24 $X2=2.89 $Y2=0.245
cc_9 VNB N_C_c_292_n 0.0564636f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.56
cc_10 VNB N_C_c_293_n 0.0122497f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.41
cc_11 VNB N_C_c_294_n 0.022726f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.41
cc_12 VNB N_C_c_295_n 0.011844f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=0.995
cc_13 VNB N_C_c_296_n 0.00674928f $X=-0.19 $Y=-0.24 $X2=1.295 $Y2=0.78
cc_14 VNB N_A_335_93#_c_356_n 0.0267993f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.995
cc_15 VNB N_A_335_93#_c_357_n 0.0219005f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.41
cc_16 VNB N_A_335_93#_c_358_n 0.00270846f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=0.56
cc_17 VNB N_A_335_93#_c_359_n 0.00243033f $X=-0.19 $Y=-0.24 $X2=1.755 $Y2=2.235
cc_18 VNB N_A_934_297#_M1011_g 0.0360507f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.985
cc_19 VNB N_A_934_297#_c_432_n 0.0291121f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.985
cc_20 VNB N_A_934_297#_c_433_n 0.00143998f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.985
cc_21 VNB N_A_934_297#_c_434_n 0.0195477f $X=-0.19 $Y=-0.24 $X2=1.21 $Y2=1.325
cc_22 VNB N_A_934_297#_c_435_n 0.0291447f $X=-0.19 $Y=-0.24 $X2=1.295 $Y2=0.78
cc_23 VNB N_A_934_297#_c_436_n 0.0176862f $X=-0.19 $Y=-0.24 $X2=1.645 $Y2=1.96
cc_24 VNB N_A_934_297#_c_437_n 0.00235412f $X=-0.19 $Y=-0.24 $X2=1.195 $Y2=0.78
cc_25 VNB N_A_934_297#_c_438_n 0.00793619f $X=-0.19 $Y=-0.24 $X2=1.18 $Y2=1.16
cc_26 VNB N_A_934_297#_c_439_n 0.0128101f $X=-0.19 $Y=-0.24 $X2=3.025 $Y2=0.355
cc_27 VNB N_A_934_297#_c_440_n 0.00135073f $X=-0.19 $Y=-0.24 $X2=3.025 $Y2=0.37
cc_28 VNB N_A_934_297#_c_441_n 0.00305701f $X=-0.19 $Y=-0.24 $X2=1.18 $Y2=1.202
cc_29 VNB N_A_934_297#_c_442_n 0.00216739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_934_297#_c_443_n 0.00623207f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_934_297#_c_444_n 0.00257621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_B_M1018_g 0.0300394f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_B_c_612_n 0.0593593f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.56
cc_34 VNB N_B_c_613_n 0.0270966f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.56
cc_35 VNB N_B_M1009_g 0.0287687f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=0.995
cc_36 VNB N_B_c_615_n 0.0103656f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=2.32
cc_37 VNB N_B_c_616_n 0.0278248f $X=-0.19 $Y=-0.24 $X2=1.18 $Y2=1.16
cc_38 VNB N_B_c_617_n 0.00131358f $X=-0.19 $Y=-0.24 $X2=3.025 $Y2=0.355
cc_39 VNB N_B_c_618_n 0.0212564f $X=-0.19 $Y=-0.24 $X2=3.025 $Y2=0.37
cc_40 VNB N_A_c_746_n 0.0230527f $X=-0.19 $Y=-0.24 $X2=2.89 $Y2=0.245
cc_41 VNB N_A_c_747_n 0.0182219f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB A 0.00404679f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.995
cc_43 VNB N_A_1050_365#_c_784_n 0.0267203f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.41
cc_44 VNB N_A_1050_365#_c_785_n 0.0198808f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=0.995
cc_45 VNB N_A_1050_365#_c_786_n 0.00641545f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.78
cc_46 VNB N_A_1050_365#_c_787_n 0.00275527f $X=-0.19 $Y=-0.24 $X2=1.755
+ $Y2=2.045
cc_47 VNB N_A_1050_365#_c_788_n 0.0020163f $X=-0.19 $Y=-0.24 $X2=1.755 $Y2=2.235
cc_48 VNB N_A_1050_365#_c_789_n 0.00350271f $X=-0.19 $Y=-0.24 $X2=2.785 $Y2=0.34
cc_49 VNB N_A_1050_365#_c_790_n 0.00203513f $X=-0.19 $Y=-0.24 $X2=1.18 $Y2=1.16
cc_50 VNB N_A_1050_365#_c_791_n 0.0051341f $X=-0.19 $Y=-0.24 $X2=3.025 $Y2=0.37
cc_51 VNB N_VPWR_c_914_n 0.402575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_X_c_1021_n 0.0041685f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.41
cc_53 VNB N_X_c_1022_n 0.0155504f $X=-0.19 $Y=-0.24 $X2=1.635 $Y2=0.425
cc_54 VNB N_A_465_325#_c_1066_n 0.00971866f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.78
cc_55 VNB N_A_465_325#_c_1067_n 0.0097913f $X=-0.19 $Y=-0.24 $X2=1.745 $Y2=0.34
cc_56 VNB N_A_483_49#_c_1213_n 0.0026438f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.41
cc_57 VNB N_A_483_49#_c_1214_n 0.00847369f $X=-0.19 $Y=-0.24 $X2=1.21 $Y2=1.325
cc_58 VNB N_A_483_49#_c_1215_n 0.0139223f $X=-0.19 $Y=-0.24 $X2=1.635 $Y2=0.695
cc_59 VNB N_A_483_49#_c_1216_n 0.00304946f $X=-0.19 $Y=-0.24 $X2=1.755 $Y2=2.235
cc_60 VNB N_A_483_49#_c_1217_n 0.00223545f $X=-0.19 $Y=-0.24 $X2=1.195 $Y2=1.16
cc_61 VNB N_A_483_49#_c_1218_n 0.0107774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_483_49#_c_1219_n 3.37974e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1335_297#_c_1400_n 0.00788636f $X=-0.19 $Y=-0.24 $X2=0.975
+ $Y2=1.985
cc_64 VNB N_A_1335_297#_c_1401_n 0.0311231f $X=-0.19 $Y=-0.24 $X2=1.635
+ $Y2=0.695
cc_65 VNB N_A_1335_297#_c_1402_n 0.0140863f $X=-0.19 $Y=-0.24 $X2=1.195 $Y2=1.16
cc_66 VNB N_VGND_c_1466_n 0.010622f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.41
cc_67 VNB N_VGND_c_1467_n 0.0125979f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.985
cc_68 VNB N_VGND_c_1468_n 0.0172244f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=0.56
cc_69 VNB N_VGND_c_1469_n 0.00462216f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.78
cc_70 VNB N_VGND_c_1470_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=1.635 $Y2=0.425
cc_71 VNB N_VGND_c_1471_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=2.785 $Y2=0.34
cc_72 VNB N_VGND_c_1472_n 0.071878f $X=-0.19 $Y=-0.24 $X2=3.025 $Y2=2.32
cc_73 VNB N_VGND_c_1473_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=3.025 $Y2=2.32
cc_74 VNB N_VGND_c_1474_n 0.109008f $X=-0.19 $Y=-0.24 $X2=1.195 $Y2=0.78
cc_75 VNB N_VGND_c_1475_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=1.195 $Y2=1.16
cc_76 VNB N_VGND_c_1476_n 0.0213733f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1477_n 0.484822f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1478_n 0.00478003f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VPB N_A_81_21#_c_172_n 0.0184001f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.41
cc_80 VPB N_A_81_21#_c_173_n 0.0191601f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.41
cc_81 VPB N_A_81_21#_c_167_n 0.00111888f $X=-0.19 $Y=1.305 $X2=1.21 $Y2=1.325
cc_82 VPB N_A_81_21#_c_175_n 0.0027789f $X=-0.19 $Y=1.305 $X2=1.21 $Y2=1.875
cc_83 VPB N_A_81_21#_c_176_n 0.0038652f $X=-0.19 $Y=1.305 $X2=1.755 $Y2=2.235
cc_84 VPB N_A_81_21#_c_177_n 0.00112766f $X=-0.19 $Y=1.305 $X2=1.865 $Y2=2.32
cc_85 VPB N_A_81_21#_c_178_n 0.0127396f $X=-0.19 $Y=1.305 $X2=3.025 $Y2=2.32
cc_86 VPB N_A_81_21#_c_171_n 0.0290227f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.202
cc_87 VPB N_C_M1012_g 0.0323013f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.995
cc_88 VPB N_C_c_292_n 0.0268393f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.56
cc_89 VPB N_C_c_293_n 0.0395822f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.41
cc_90 VPB N_C_c_295_n 0.00718175f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=0.995
cc_91 VPB N_C_c_296_n 0.00448796f $X=-0.19 $Y=1.305 $X2=1.295 $Y2=0.78
cc_92 VPB N_A_335_93#_c_356_n 0.0399465f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.995
cc_93 VPB N_A_335_93#_c_358_n 0.00446988f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=0.56
cc_94 VPB N_A_335_93#_c_362_n 0.0160888f $X=-0.19 $Y=1.305 $X2=1.21 $Y2=1.875
cc_95 VPB N_A_335_93#_c_363_n 0.00230347f $X=-0.19 $Y=1.305 $X2=1.645 $Y2=1.96
cc_96 VPB N_A_335_93#_c_364_n 0.00173244f $X=-0.19 $Y=1.305 $X2=1.295 $Y2=1.96
cc_97 VPB N_A_335_93#_c_359_n 2.7219e-19 $X=-0.19 $Y=1.305 $X2=1.755 $Y2=2.235
cc_98 VPB N_A_934_297#_c_445_n 0.0204741f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.995
cc_99 VPB N_A_934_297#_c_433_n 0.0104902f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.985
cc_100 VPB N_A_934_297#_c_447_n 0.0239536f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=0.995
cc_101 VPB N_A_934_297#_c_435_n 0.0105828f $X=-0.19 $Y=1.305 $X2=1.295 $Y2=0.78
cc_102 VPB N_A_934_297#_c_436_n 0.00766961f $X=-0.19 $Y=1.305 $X2=1.645 $Y2=1.96
cc_103 VPB N_A_934_297#_c_450_n 0.00591035f $X=-0.19 $Y=1.305 $X2=1.755
+ $Y2=2.045
cc_104 VPB N_A_934_297#_c_444_n 0.0032041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_B_c_619_n 0.0216572f $X=-0.19 $Y=1.305 $X2=2.89 $Y2=0.245
cc_106 VPB N_B_c_613_n 0.00747973f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.56
cc_107 VPB N_B_M1021_g 0.0155329f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.41
cc_108 VPB N_B_c_622_n 0.12486f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=0.56
cc_109 VPB N_B_c_623_n 0.0170126f $X=-0.19 $Y=1.305 $X2=1.21 $Y2=1.325
cc_110 VPB N_B_c_624_n 0.0101708f $X=-0.19 $Y=1.305 $X2=1.295 $Y2=1.96
cc_111 VPB N_B_c_625_n 0.00717497f $X=-0.19 $Y=1.305 $X2=1.635 $Y2=0.425
cc_112 VPB N_B_M1014_g 0.0130358f $X=-0.19 $Y=1.305 $X2=1.755 $Y2=2.235
cc_113 VPB N_B_c_615_n 0.0087608f $X=-0.19 $Y=1.305 $X2=1.865 $Y2=2.32
cc_114 VPB B 0.00185689f $X=-0.19 $Y=1.305 $X2=3.025 $Y2=2.32
cc_115 VPB N_B_c_616_n 0.00425314f $X=-0.19 $Y=1.305 $X2=1.18 $Y2=1.16
cc_116 VPB N_B_c_617_n 9.77983e-19 $X=-0.19 $Y=1.305 $X2=3.025 $Y2=0.355
cc_117 VPB N_B_c_631_n 0.00411193f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_c_746_n 0.02697f $X=-0.19 $Y=1.305 $X2=2.89 $Y2=0.245
cc_119 VPB A 0.00142645f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.995
cc_120 VPB N_A_1050_365#_c_784_n 0.0291085f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.41
cc_121 VPB N_A_1050_365#_c_786_n 0.00273235f $X=-0.19 $Y=1.305 $X2=1.525
+ $Y2=0.78
cc_122 VPB N_A_1050_365#_c_794_n 0.00176559f $X=-0.19 $Y=1.305 $X2=1.645
+ $Y2=1.96
cc_123 VPB N_A_1050_365#_c_789_n 2.7046e-19 $X=-0.19 $Y=1.305 $X2=2.785 $Y2=0.34
cc_124 VPB N_A_1050_365#_c_796_n 0.00156472f $X=-0.19 $Y=1.305 $X2=1.745
+ $Y2=0.34
cc_125 VPB N_VPWR_c_915_n 0.0106835f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.41
cc_126 VPB N_VPWR_c_916_n 0.0147646f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.985
cc_127 VPB N_VPWR_c_917_n 0.0174747f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=0.56
cc_128 VPB N_VPWR_c_918_n 0.00957549f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=0.78
cc_129 VPB N_VPWR_c_919_n 0.00804433f $X=-0.19 $Y=1.305 $X2=1.635 $Y2=0.425
cc_130 VPB N_VPWR_c_920_n 0.00563188f $X=-0.19 $Y=1.305 $X2=1.755 $Y2=2.235
cc_131 VPB N_VPWR_c_921_n 0.0960902f $X=-0.19 $Y=1.305 $X2=1.865 $Y2=2.32
cc_132 VPB N_VPWR_c_922_n 0.0663405f $X=-0.19 $Y=1.305 $X2=1.195 $Y2=1.16
cc_133 VPB N_VPWR_c_923_n 0.0172188f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_914_n 0.0731114f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_925_n 0.00641289f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_926_n 0.00513206f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_X_c_1023_n 0.00324118f $X=-0.19 $Y=1.305 $X2=1.295 $Y2=1.96
cc_138 VPB N_X_c_1022_n 0.00602721f $X=-0.19 $Y=1.305 $X2=1.635 $Y2=0.425
cc_139 VPB N_A_465_325#_c_1068_n 0.00306017f $X=-0.19 $Y=1.305 $X2=0.975
+ $Y2=1.41
cc_140 VPB N_A_465_325#_c_1066_n 0.00164253f $X=-0.19 $Y=1.305 $X2=1.525
+ $Y2=0.78
cc_141 VPB N_A_465_325#_c_1070_n 0.00270715f $X=-0.19 $Y=1.305 $X2=1.645
+ $Y2=1.96
cc_142 VPB N_A_465_325#_c_1071_n 8.62277e-19 $X=-0.19 $Y=1.305 $X2=1.755
+ $Y2=2.045
cc_143 VPB N_A_465_325#_c_1067_n 0.0021572f $X=-0.19 $Y=1.305 $X2=1.745 $Y2=0.34
cc_144 VPB N_A_465_325#_c_1073_n 0.0148089f $X=-0.19 $Y=1.305 $X2=1.18 $Y2=1.16
cc_145 VPB N_A_465_325#_c_1074_n 0.00318502f $X=-0.19 $Y=1.305 $X2=3.025
+ $Y2=0.355
cc_146 VPB N_A_465_325#_c_1075_n 0.0015478f $X=-0.19 $Y=1.305 $X2=0.975
+ $Y2=1.202
cc_147 VPB N_A_465_325#_c_1076_n 0.0215932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_483_49#_c_1220_n 0.0026444f $X=-0.19 $Y=1.305 $X2=1.295 $Y2=0.78
cc_149 VPB N_A_483_49#_c_1221_n 0.00579762f $X=-0.19 $Y=1.305 $X2=1.645 $Y2=1.96
cc_150 VPB N_A_483_49#_c_1222_n 8.62166e-19 $X=-0.19 $Y=1.305 $X2=1.295 $Y2=1.96
cc_151 VPB N_A_483_49#_c_1216_n 0.00847729f $X=-0.19 $Y=1.305 $X2=1.755
+ $Y2=2.235
cc_152 VPB N_A_483_49#_c_1224_n 0.00306425f $X=-0.19 $Y=1.305 $X2=2.785 $Y2=0.34
cc_153 VPB N_A_483_49#_c_1225_n 0.00298222f $X=-0.19 $Y=1.305 $X2=3.025 $Y2=2.32
cc_154 VPB N_A_483_49#_c_1226_n 0.0103424f $X=-0.19 $Y=1.305 $X2=3.025 $Y2=2.32
cc_155 VPB N_A_483_49#_c_1227_n 0.00185607f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_483_49#_c_1217_n 0.00149669f $X=-0.19 $Y=1.305 $X2=1.195 $Y2=1.16
cc_157 VPB N_A_483_49#_c_1229_n 0.024688f $X=-0.19 $Y=1.305 $X2=3.025 $Y2=0.355
cc_158 VPB N_A_483_49#_c_1230_n 0.00221665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_483_49#_c_1231_n 2.86933e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_483_49#_c_1232_n 3.79061e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_1335_297#_c_1400_n 0.00457449f $X=-0.19 $Y=1.305 $X2=0.975
+ $Y2=1.985
cc_162 VPB N_A_1335_297#_c_1404_n 0.015197f $X=-0.19 $Y=1.305 $X2=1.645 $Y2=1.96
cc_163 VPB N_A_1335_297#_c_1401_n 0.0233363f $X=-0.19 $Y=1.305 $X2=1.635
+ $Y2=0.695
cc_164 VPB N_A_1335_297#_c_1406_n 0.0103928f $X=-0.19 $Y=1.305 $X2=1.865
+ $Y2=2.32
cc_165 N_A_81_21#_c_166_n N_C_c_291_n 0.0122002f $X=0.98 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_166 N_A_81_21#_c_167_n N_C_c_291_n 0.00138795f $X=1.21 $Y=1.325 $X2=-0.19
+ $Y2=-0.24
cc_167 N_A_81_21#_c_182_p N_C_c_291_n 0.0123036f $X=1.525 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_168 N_A_81_21#_c_168_n N_C_c_291_n 0.010641f $X=1.635 $Y=0.695 $X2=-0.19
+ $Y2=-0.24
cc_169 N_A_81_21#_c_169_n N_C_c_291_n 0.00580453f $X=1.745 $Y=0.34 $X2=-0.19
+ $Y2=-0.24
cc_170 N_A_81_21#_c_173_n N_C_M1012_g 0.0186648f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_81_21#_c_175_n N_C_M1012_g 0.00553088f $X=1.21 $Y=1.875 $X2=0 $Y2=0
cc_172 N_A_81_21#_c_187_p N_C_M1012_g 0.0133197f $X=1.645 $Y=1.96 $X2=0 $Y2=0
cc_173 N_A_81_21#_c_176_n N_C_M1012_g 0.00763977f $X=1.755 $Y=2.235 $X2=0 $Y2=0
cc_174 N_A_81_21#_c_177_n N_C_M1012_g 0.00747755f $X=1.865 $Y=2.32 $X2=0 $Y2=0
cc_175 N_A_81_21#_c_170_n N_C_c_292_n 0.00948274f $X=2.785 $Y=0.355 $X2=0 $Y2=0
cc_176 N_A_81_21#_c_178_n N_C_c_293_n 0.0112964f $X=3.025 $Y=2.32 $X2=0 $Y2=0
cc_177 N_A_81_21#_c_192_p N_C_c_294_n 0.00558632f $X=3.025 $Y=0.37 $X2=0 $Y2=0
cc_178 N_A_81_21#_c_170_n N_C_c_294_n 0.00582901f $X=2.785 $Y=0.355 $X2=0 $Y2=0
cc_179 N_A_81_21#_c_167_n N_C_c_295_n 0.00158401f $X=1.21 $Y=1.325 $X2=0 $Y2=0
cc_180 N_A_81_21#_c_175_n N_C_c_295_n 9.13902e-19 $X=1.21 $Y=1.875 $X2=0 $Y2=0
cc_181 N_A_81_21#_c_171_n N_C_c_295_n 0.0257806f $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_182 N_A_81_21#_c_170_n N_C_c_296_n 0.0032871f $X=2.785 $Y=0.355 $X2=0 $Y2=0
cc_183 N_A_81_21#_c_182_p N_A_335_93#_M1008_d 0.00214557f $X=1.525 $Y=0.78
+ $X2=-0.19 $Y2=-0.24
cc_184 N_A_81_21#_c_168_n N_A_335_93#_M1008_d 0.00618081f $X=1.635 $Y=0.695
+ $X2=-0.19 $Y2=-0.24
cc_185 N_A_81_21#_c_187_p N_A_335_93#_M1012_d 0.00436734f $X=1.645 $Y=1.96 $X2=0
+ $Y2=0
cc_186 N_A_81_21#_c_176_n N_A_335_93#_M1012_d 0.00269214f $X=1.755 $Y=2.235
+ $X2=0 $Y2=0
cc_187 N_A_81_21#_c_178_n N_A_335_93#_c_356_n 0.00841967f $X=3.025 $Y=2.32 $X2=0
+ $Y2=0
cc_188 N_A_81_21#_c_192_p N_A_335_93#_c_357_n 0.00165819f $X=3.025 $Y=0.37 $X2=0
+ $Y2=0
cc_189 N_A_81_21#_c_182_p N_A_335_93#_c_372_n 0.00402121f $X=1.525 $Y=0.78 $X2=0
+ $Y2=0
cc_190 N_A_81_21#_c_187_p N_A_335_93#_c_372_n 0.0200253f $X=1.645 $Y=1.96 $X2=0
+ $Y2=0
cc_191 N_A_81_21#_c_178_n N_A_335_93#_c_372_n 0.00160427f $X=3.025 $Y=2.32 $X2=0
+ $Y2=0
cc_192 N_A_81_21#_c_167_n N_A_335_93#_c_358_n 0.0116338f $X=1.21 $Y=1.325 $X2=0
+ $Y2=0
cc_193 N_A_81_21#_c_175_n N_A_335_93#_c_358_n 0.00617983f $X=1.21 $Y=1.875 $X2=0
+ $Y2=0
cc_194 N_A_81_21#_c_182_p N_A_335_93#_c_358_n 0.013727f $X=1.525 $Y=0.78 $X2=0
+ $Y2=0
cc_195 N_A_81_21#_c_168_n N_A_335_93#_c_358_n 0.00736858f $X=1.635 $Y=0.695
+ $X2=0 $Y2=0
cc_196 N_A_81_21#_c_170_n N_A_335_93#_c_358_n 0.0130244f $X=2.785 $Y=0.355 $X2=0
+ $Y2=0
cc_197 N_A_81_21#_c_171_n N_A_335_93#_c_358_n 7.48596e-19 $X=0.98 $Y=1.202 $X2=0
+ $Y2=0
cc_198 N_A_81_21#_M1013_d N_A_335_93#_c_362_n 0.00327687f $X=2.835 $Y=1.625
+ $X2=0 $Y2=0
cc_199 N_A_81_21#_c_178_n N_A_335_93#_c_362_n 0.00614909f $X=3.025 $Y=2.32 $X2=0
+ $Y2=0
cc_200 N_A_81_21#_c_178_n N_A_335_93#_c_364_n 0.00632099f $X=3.025 $Y=2.32 $X2=0
+ $Y2=0
cc_201 N_A_81_21#_c_175_n N_VPWR_M1022_s 0.011386f $X=1.21 $Y=1.875 $X2=0 $Y2=0
cc_202 N_A_81_21#_c_187_p N_VPWR_M1022_s 0.00908042f $X=1.645 $Y=1.96 $X2=0
+ $Y2=0
cc_203 N_A_81_21#_c_218_p N_VPWR_M1022_s 0.00499482f $X=1.295 $Y=1.96 $X2=0
+ $Y2=0
cc_204 N_A_81_21#_c_172_n N_VPWR_c_916_n 0.00934006f $X=0.505 $Y=1.41 $X2=0
+ $Y2=0
cc_205 N_A_81_21#_c_173_n N_VPWR_c_916_n 9.95344e-19 $X=0.975 $Y=1.41 $X2=0
+ $Y2=0
cc_206 N_A_81_21#_c_172_n N_VPWR_c_917_n 0.00458723f $X=0.505 $Y=1.41 $X2=0
+ $Y2=0
cc_207 N_A_81_21#_c_173_n N_VPWR_c_917_n 0.00673617f $X=0.975 $Y=1.41 $X2=0
+ $Y2=0
cc_208 N_A_81_21#_c_173_n N_VPWR_c_918_n 0.0086641f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A_81_21#_c_187_p N_VPWR_c_918_n 0.0126462f $X=1.645 $Y=1.96 $X2=0 $Y2=0
cc_210 N_A_81_21#_c_218_p N_VPWR_c_918_n 0.0143755f $X=1.295 $Y=1.96 $X2=0 $Y2=0
cc_211 N_A_81_21#_c_176_n N_VPWR_c_918_n 0.00141178f $X=1.755 $Y=2.235 $X2=0
+ $Y2=0
cc_212 N_A_81_21#_c_177_n N_VPWR_c_918_n 0.0133539f $X=1.865 $Y=2.32 $X2=0 $Y2=0
cc_213 N_A_81_21#_c_187_p N_VPWR_c_922_n 0.00241968f $X=1.645 $Y=1.96 $X2=0
+ $Y2=0
cc_214 N_A_81_21#_c_177_n N_VPWR_c_922_n 0.0109705f $X=1.865 $Y=2.32 $X2=0 $Y2=0
cc_215 N_A_81_21#_c_178_n N_VPWR_c_922_n 0.0642605f $X=3.025 $Y=2.32 $X2=0 $Y2=0
cc_216 N_A_81_21#_c_172_n N_VPWR_c_914_n 0.00523894f $X=0.505 $Y=1.41 $X2=0
+ $Y2=0
cc_217 N_A_81_21#_c_173_n N_VPWR_c_914_n 0.0132531f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A_81_21#_c_187_p N_VPWR_c_914_n 0.00567317f $X=1.645 $Y=1.96 $X2=0
+ $Y2=0
cc_219 N_A_81_21#_c_218_p N_VPWR_c_914_n 7.91584e-19 $X=1.295 $Y=1.96 $X2=0
+ $Y2=0
cc_220 N_A_81_21#_c_177_n N_VPWR_c_914_n 0.00809357f $X=1.865 $Y=2.32 $X2=0
+ $Y2=0
cc_221 N_A_81_21#_c_178_n N_VPWR_c_914_n 0.0515593f $X=3.025 $Y=2.32 $X2=0 $Y2=0
cc_222 N_A_81_21#_c_173_n N_X_c_1025_n 0.00667442f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A_81_21#_c_165_n N_X_c_1021_n 0.0153207f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A_81_21#_c_166_n N_X_c_1021_n 0.00683169f $X=0.98 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A_81_21#_c_167_n N_X_c_1021_n 0.017335f $X=1.21 $Y=1.325 $X2=0 $Y2=0
cc_226 N_A_81_21#_c_168_n N_X_c_1021_n 9.11008e-19 $X=1.635 $Y=0.695 $X2=0 $Y2=0
cc_227 N_A_81_21#_c_171_n N_X_c_1021_n 0.00406447f $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_228 N_A_81_21#_c_165_n N_X_c_1031_n 0.00567701f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A_81_21#_c_166_n N_X_c_1031_n 0.00499441f $X=0.98 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A_81_21#_c_168_n N_X_c_1031_n 0.00341331f $X=1.635 $Y=0.695 $X2=0 $Y2=0
cc_231 N_A_81_21#_c_172_n N_X_c_1023_n 0.0244282f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_232 N_A_81_21#_c_173_n N_X_c_1023_n 0.00822531f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_233 N_A_81_21#_c_175_n N_X_c_1023_n 0.027545f $X=1.21 $Y=1.875 $X2=0 $Y2=0
cc_234 N_A_81_21#_c_218_p N_X_c_1023_n 0.0119692f $X=1.295 $Y=1.96 $X2=0 $Y2=0
cc_235 N_A_81_21#_c_171_n N_X_c_1023_n 0.00612148f $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_236 N_A_81_21#_c_165_n N_X_c_1022_n 0.00312365f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A_81_21#_c_172_n N_X_c_1022_n 0.00109528f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_238 N_A_81_21#_c_173_n N_X_c_1022_n 2.66476e-19 $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_239 N_A_81_21#_c_166_n N_X_c_1022_n 6.4569e-19 $X=0.98 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A_81_21#_c_167_n N_X_c_1022_n 0.0150382f $X=1.21 $Y=1.325 $X2=0 $Y2=0
cc_241 N_A_81_21#_c_175_n N_X_c_1022_n 0.00477144f $X=1.21 $Y=1.875 $X2=0 $Y2=0
cc_242 N_A_81_21#_c_171_n N_X_c_1022_n 0.0292276f $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_243 N_A_81_21#_c_178_n N_A_465_325#_M1013_s 0.00721138f $X=3.025 $Y=2.32
+ $X2=0 $Y2=0
cc_244 N_A_81_21#_M1013_d N_A_465_325#_c_1068_n 0.00649326f $X=2.835 $Y=1.625
+ $X2=0 $Y2=0
cc_245 N_A_81_21#_c_187_p N_A_465_325#_c_1068_n 0.00740552f $X=1.645 $Y=1.96
+ $X2=0 $Y2=0
cc_246 N_A_81_21#_c_176_n N_A_465_325#_c_1068_n 8.52135e-19 $X=1.755 $Y=2.235
+ $X2=0 $Y2=0
cc_247 N_A_81_21#_c_178_n N_A_465_325#_c_1068_n 0.0612998f $X=3.025 $Y=2.32
+ $X2=0 $Y2=0
cc_248 N_A_81_21#_c_170_n N_A_483_49#_M1002_s 0.00684027f $X=2.785 $Y=0.355
+ $X2=-0.19 $Y2=-0.24
cc_249 N_A_81_21#_M1002_d N_A_483_49#_c_1213_n 0.0127352f $X=2.89 $Y=0.245 $X2=0
+ $Y2=0
cc_250 N_A_81_21#_c_192_p N_A_483_49#_c_1213_n 0.0206573f $X=3.025 $Y=0.37 $X2=0
+ $Y2=0
cc_251 N_A_81_21#_c_170_n N_A_483_49#_c_1213_n 0.0191269f $X=2.785 $Y=0.355
+ $X2=0 $Y2=0
cc_252 N_A_81_21#_c_192_p N_A_483_49#_c_1237_n 0.00219372f $X=3.025 $Y=0.37
+ $X2=0 $Y2=0
cc_253 N_A_81_21#_c_192_p N_A_483_49#_c_1238_n 0.0147713f $X=3.025 $Y=0.37 $X2=0
+ $Y2=0
cc_254 N_A_81_21#_c_178_n N_A_483_49#_c_1230_n 0.0100105f $X=3.025 $Y=2.32 $X2=0
+ $Y2=0
cc_255 N_A_81_21#_c_167_n N_VGND_M1016_s 0.00493665f $X=1.21 $Y=1.325 $X2=0
+ $Y2=0
cc_256 N_A_81_21#_c_182_p N_VGND_M1016_s 0.00907954f $X=1.525 $Y=0.78 $X2=0
+ $Y2=0
cc_257 N_A_81_21#_c_165_n N_VGND_c_1467_n 0.00929407f $X=0.48 $Y=0.995 $X2=0
+ $Y2=0
cc_258 N_A_81_21#_c_166_n N_VGND_c_1467_n 8.51748e-19 $X=0.98 $Y=0.995 $X2=0
+ $Y2=0
cc_259 N_A_81_21#_c_165_n N_VGND_c_1468_n 0.00342263f $X=0.48 $Y=0.995 $X2=0
+ $Y2=0
cc_260 N_A_81_21#_c_166_n N_VGND_c_1468_n 0.0055096f $X=0.98 $Y=0.995 $X2=0
+ $Y2=0
cc_261 N_A_81_21#_c_166_n N_VGND_c_1469_n 0.00637763f $X=0.98 $Y=0.995 $X2=0
+ $Y2=0
cc_262 N_A_81_21#_c_167_n N_VGND_c_1469_n 0.0151684f $X=1.21 $Y=1.325 $X2=0
+ $Y2=0
cc_263 N_A_81_21#_c_182_p N_VGND_c_1469_n 0.00454809f $X=1.525 $Y=0.78 $X2=0
+ $Y2=0
cc_264 N_A_81_21#_c_168_n N_VGND_c_1469_n 0.00733827f $X=1.635 $Y=0.695 $X2=0
+ $Y2=0
cc_265 N_A_81_21#_c_169_n N_VGND_c_1469_n 0.0140929f $X=1.745 $Y=0.34 $X2=0
+ $Y2=0
cc_266 N_A_81_21#_c_171_n N_VGND_c_1469_n 7.93989e-19 $X=0.98 $Y=1.202 $X2=0
+ $Y2=0
cc_267 N_A_81_21#_c_182_p N_VGND_c_1472_n 0.0022086f $X=1.525 $Y=0.78 $X2=0
+ $Y2=0
cc_268 N_A_81_21#_c_169_n N_VGND_c_1472_n 0.0156439f $X=1.745 $Y=0.34 $X2=0
+ $Y2=0
cc_269 N_A_81_21#_c_170_n N_VGND_c_1472_n 0.088963f $X=2.785 $Y=0.355 $X2=0
+ $Y2=0
cc_270 N_A_81_21#_c_165_n N_VGND_c_1477_n 0.00424115f $X=0.48 $Y=0.995 $X2=0
+ $Y2=0
cc_271 N_A_81_21#_c_166_n N_VGND_c_1477_n 0.0113468f $X=0.98 $Y=0.995 $X2=0
+ $Y2=0
cc_272 N_A_81_21#_c_167_n N_VGND_c_1477_n 7.71903e-19 $X=1.21 $Y=1.325 $X2=0
+ $Y2=0
cc_273 N_A_81_21#_c_182_p N_VGND_c_1477_n 0.00486519f $X=1.525 $Y=0.78 $X2=0
+ $Y2=0
cc_274 N_A_81_21#_c_169_n N_VGND_c_1477_n 0.00844855f $X=1.745 $Y=0.34 $X2=0
+ $Y2=0
cc_275 N_A_81_21#_c_170_n N_VGND_c_1477_n 0.0531745f $X=2.785 $Y=0.355 $X2=0
+ $Y2=0
cc_276 N_C_c_293_n N_A_335_93#_c_356_n 0.049491f $X=2.745 $Y=1.55 $X2=0 $Y2=0
cc_277 N_C_c_296_n N_A_335_93#_c_356_n 0.00113464f $X=2.705 $Y=1.16 $X2=0 $Y2=0
cc_278 N_C_c_294_n N_A_335_93#_c_357_n 0.0200603f $X=2.815 $Y=0.995 $X2=0 $Y2=0
cc_279 N_C_M1012_g N_A_335_93#_c_372_n 0.0115705f $X=1.625 $Y=1.805 $X2=0 $Y2=0
cc_280 N_C_c_292_n N_A_335_93#_c_372_n 0.00616727f $X=2.645 $Y=1.16 $X2=0 $Y2=0
cc_281 N_C_c_291_n N_A_335_93#_c_358_n 0.00440057f $X=1.6 $Y=0.995 $X2=0 $Y2=0
cc_282 N_C_M1012_g N_A_335_93#_c_358_n 0.00204947f $X=1.625 $Y=1.805 $X2=0 $Y2=0
cc_283 N_C_c_292_n N_A_335_93#_c_358_n 0.024155f $X=2.645 $Y=1.16 $X2=0 $Y2=0
cc_284 N_C_c_293_n N_A_335_93#_c_358_n 0.00495404f $X=2.745 $Y=1.55 $X2=0 $Y2=0
cc_285 N_C_c_294_n N_A_335_93#_c_358_n 0.00291386f $X=2.815 $Y=0.995 $X2=0 $Y2=0
cc_286 N_C_c_295_n N_A_335_93#_c_358_n 0.00205064f $X=1.625 $Y=1.202 $X2=0 $Y2=0
cc_287 N_C_c_296_n N_A_335_93#_c_358_n 0.0250283f $X=2.705 $Y=1.16 $X2=0 $Y2=0
cc_288 N_C_c_292_n N_A_335_93#_c_362_n 0.00875365f $X=2.645 $Y=1.16 $X2=0 $Y2=0
cc_289 N_C_c_293_n N_A_335_93#_c_362_n 0.0166592f $X=2.745 $Y=1.55 $X2=0 $Y2=0
cc_290 N_C_c_296_n N_A_335_93#_c_362_n 0.0433923f $X=2.705 $Y=1.16 $X2=0 $Y2=0
cc_291 N_C_c_293_n N_A_335_93#_c_363_n 0.00411747f $X=2.745 $Y=1.55 $X2=0 $Y2=0
cc_292 N_C_c_293_n N_A_335_93#_c_359_n 0.00100598f $X=2.745 $Y=1.55 $X2=0 $Y2=0
cc_293 N_C_c_296_n N_A_335_93#_c_359_n 0.028998f $X=2.705 $Y=1.16 $X2=0 $Y2=0
cc_294 N_C_M1012_g N_VPWR_c_918_n 0.00220316f $X=1.625 $Y=1.805 $X2=0 $Y2=0
cc_295 N_C_M1012_g N_VPWR_c_922_n 0.00514356f $X=1.625 $Y=1.805 $X2=0 $Y2=0
cc_296 N_C_c_293_n N_VPWR_c_922_n 0.00427564f $X=2.745 $Y=1.55 $X2=0 $Y2=0
cc_297 N_C_M1012_g N_VPWR_c_914_n 0.00682402f $X=1.625 $Y=1.805 $X2=0 $Y2=0
cc_298 N_C_c_293_n N_VPWR_c_914_n 0.00728509f $X=2.745 $Y=1.55 $X2=0 $Y2=0
cc_299 N_C_c_291_n N_X_c_1021_n 2.13275e-19 $X=1.6 $Y=0.995 $X2=0 $Y2=0
cc_300 N_C_c_291_n N_X_c_1031_n 4.30151e-19 $X=1.6 $Y=0.995 $X2=0 $Y2=0
cc_301 N_C_M1012_g N_X_c_1023_n 8.85562e-19 $X=1.625 $Y=1.805 $X2=0 $Y2=0
cc_302 N_C_M1012_g N_A_465_325#_c_1068_n 9.28125e-19 $X=1.625 $Y=1.805 $X2=0
+ $Y2=0
cc_303 N_C_c_293_n N_A_465_325#_c_1068_n 0.0104309f $X=2.745 $Y=1.55 $X2=0 $Y2=0
cc_304 N_C_c_292_n N_A_483_49#_c_1213_n 0.00200392f $X=2.645 $Y=1.16 $X2=0 $Y2=0
cc_305 N_C_c_294_n N_A_483_49#_c_1213_n 0.00938851f $X=2.815 $Y=0.995 $X2=0
+ $Y2=0
cc_306 N_C_c_296_n N_A_483_49#_c_1213_n 0.0385625f $X=2.705 $Y=1.16 $X2=0 $Y2=0
cc_307 N_C_c_294_n N_A_483_49#_c_1237_n 7.49049e-19 $X=2.815 $Y=0.995 $X2=0
+ $Y2=0
cc_308 N_C_c_291_n N_VGND_c_1469_n 0.00111462f $X=1.6 $Y=0.995 $X2=0 $Y2=0
cc_309 N_C_c_291_n N_VGND_c_1472_n 7.72982e-19 $X=1.6 $Y=0.995 $X2=0 $Y2=0
cc_310 N_C_c_294_n N_VGND_c_1472_n 0.00357877f $X=2.815 $Y=0.995 $X2=0 $Y2=0
cc_311 N_C_c_294_n N_VGND_c_1477_n 0.00705439f $X=2.815 $Y=0.995 $X2=0 $Y2=0
cc_312 N_A_335_93#_c_356_n N_VPWR_c_922_n 0.00455111f $X=3.325 $Y=1.55 $X2=0
+ $Y2=0
cc_313 N_A_335_93#_c_356_n N_VPWR_c_914_n 0.00760152f $X=3.325 $Y=1.55 $X2=0
+ $Y2=0
cc_314 N_A_335_93#_c_362_n N_A_465_325#_M1013_s 0.00366147f $X=3.11 $Y=1.62
+ $X2=0 $Y2=0
cc_315 N_A_335_93#_c_356_n N_A_465_325#_c_1068_n 0.0173326f $X=3.325 $Y=1.55
+ $X2=0 $Y2=0
cc_316 N_A_335_93#_c_362_n N_A_465_325#_c_1068_n 0.0559645f $X=3.11 $Y=1.62
+ $X2=0 $Y2=0
cc_317 N_A_335_93#_c_359_n N_A_465_325#_c_1068_n 0.00386917f $X=3.3 $Y=1.16
+ $X2=0 $Y2=0
cc_318 N_A_335_93#_c_356_n N_A_465_325#_c_1088_n 0.00748858f $X=3.325 $Y=1.55
+ $X2=0 $Y2=0
cc_319 N_A_335_93#_c_362_n N_A_465_325#_c_1088_n 6.13389e-19 $X=3.11 $Y=1.62
+ $X2=0 $Y2=0
cc_320 N_A_335_93#_c_356_n N_A_465_325#_c_1066_n 9.67237e-19 $X=3.325 $Y=1.55
+ $X2=0 $Y2=0
cc_321 N_A_335_93#_c_357_n N_A_465_325#_c_1066_n 0.0136697f $X=3.41 $Y=0.995
+ $X2=0 $Y2=0
cc_322 N_A_335_93#_c_363_n N_A_465_325#_c_1066_n 0.00166649f $X=3.195 $Y=1.535
+ $X2=0 $Y2=0
cc_323 N_A_335_93#_c_359_n N_A_465_325#_c_1066_n 0.015773f $X=3.3 $Y=1.16 $X2=0
+ $Y2=0
cc_324 N_A_335_93#_c_362_n N_A_465_325#_c_1074_n 4.56942e-19 $X=3.11 $Y=1.62
+ $X2=0 $Y2=0
cc_325 N_A_335_93#_c_363_n N_A_465_325#_c_1074_n 6.00479e-19 $X=3.195 $Y=1.535
+ $X2=0 $Y2=0
cc_326 N_A_335_93#_c_356_n N_A_465_325#_c_1076_n 0.00700676f $X=3.325 $Y=1.55
+ $X2=0 $Y2=0
cc_327 N_A_335_93#_c_362_n N_A_465_325#_c_1076_n 0.0109044f $X=3.11 $Y=1.62
+ $X2=0 $Y2=0
cc_328 N_A_335_93#_c_363_n N_A_465_325#_c_1076_n 0.00528578f $X=3.195 $Y=1.535
+ $X2=0 $Y2=0
cc_329 N_A_335_93#_c_356_n N_A_483_49#_c_1213_n 0.0041059f $X=3.325 $Y=1.55
+ $X2=0 $Y2=0
cc_330 N_A_335_93#_c_357_n N_A_483_49#_c_1213_n 0.0122193f $X=3.41 $Y=0.995
+ $X2=0 $Y2=0
cc_331 N_A_335_93#_c_358_n N_A_483_49#_c_1213_n 0.00977033f $X=2 $Y=0.76 $X2=0
+ $Y2=0
cc_332 N_A_335_93#_c_359_n N_A_483_49#_c_1213_n 0.0224243f $X=3.3 $Y=1.16 $X2=0
+ $Y2=0
cc_333 N_A_335_93#_c_357_n N_A_483_49#_c_1237_n 0.00958879f $X=3.41 $Y=0.995
+ $X2=0 $Y2=0
cc_334 N_A_335_93#_c_357_n N_A_483_49#_c_1238_n 0.00805112f $X=3.41 $Y=0.995
+ $X2=0 $Y2=0
cc_335 N_A_335_93#_c_356_n N_A_483_49#_c_1220_n 0.00452598f $X=3.325 $Y=1.55
+ $X2=0 $Y2=0
cc_336 N_A_335_93#_c_356_n N_A_483_49#_c_1222_n 7.6183e-19 $X=3.325 $Y=1.55
+ $X2=0 $Y2=0
cc_337 N_A_335_93#_c_357_n N_A_483_49#_c_1215_n 0.00103799f $X=3.41 $Y=0.995
+ $X2=0 $Y2=0
cc_338 N_A_335_93#_c_356_n N_A_483_49#_c_1230_n 0.00354471f $X=3.325 $Y=1.55
+ $X2=0 $Y2=0
cc_339 N_A_335_93#_c_357_n N_VGND_c_1472_n 0.00369393f $X=3.41 $Y=0.995 $X2=0
+ $Y2=0
cc_340 N_A_335_93#_c_357_n N_VGND_c_1477_n 0.0071645f $X=3.41 $Y=0.995 $X2=0
+ $Y2=0
cc_341 N_A_934_297#_c_450_n N_B_c_619_n 0.00851867f $X=4.97 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_342 N_A_934_297#_c_444_n N_B_c_619_n 8.21886e-19 $X=5.03 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_343 N_A_934_297#_c_454_p N_B_M1018_g 0.00372557f $X=5.06 $Y=0.85 $X2=0 $Y2=0
cc_344 N_A_934_297#_c_444_n N_B_M1018_g 0.0147084f $X=5.03 $Y=0.72 $X2=0 $Y2=0
cc_345 N_A_934_297#_c_438_n N_B_c_612_n 0.00502253f $X=6.25 $Y=0.85 $X2=0 $Y2=0
cc_346 N_A_934_297#_c_444_n N_B_c_612_n 0.0151314f $X=5.03 $Y=0.72 $X2=0 $Y2=0
cc_347 N_A_934_297#_c_450_n N_B_c_613_n 0.00767064f $X=4.97 $Y=1.58 $X2=0 $Y2=0
cc_348 N_A_934_297#_c_444_n N_B_c_613_n 0.00790646f $X=5.03 $Y=0.72 $X2=0 $Y2=0
cc_349 N_A_934_297#_c_445_n N_B_M1021_g 0.0117988f $X=6.585 $Y=1.41 $X2=0 $Y2=0
cc_350 N_A_934_297#_M1011_g N_B_M1009_g 0.0101671f $X=6.61 $Y=0.455 $X2=0 $Y2=0
cc_351 N_A_934_297#_c_435_n N_B_M1009_g 0.0212291f $X=6.485 $Y=1.16 $X2=0 $Y2=0
cc_352 N_A_934_297#_c_437_n N_B_M1009_g 0.00190447f $X=6.372 $Y=0.995 $X2=0
+ $Y2=0
cc_353 N_A_934_297#_c_438_n N_B_M1009_g 0.00156951f $X=6.25 $Y=0.85 $X2=0 $Y2=0
cc_354 N_A_934_297#_c_440_n N_B_M1009_g 6.73467e-19 $X=6.54 $Y=0.85 $X2=0 $Y2=0
cc_355 N_A_934_297#_c_441_n N_B_M1009_g 0.00123519f $X=6.395 $Y=0.85 $X2=0 $Y2=0
cc_356 N_A_934_297#_c_445_n N_B_c_622_n 0.0105804f $X=6.585 $Y=1.41 $X2=0 $Y2=0
cc_357 N_A_934_297#_c_447_n N_B_c_622_n 0.00616735f $X=8.075 $Y=1.57 $X2=0 $Y2=0
cc_358 N_A_934_297#_c_433_n N_B_c_624_n 0.00325476f $X=8.075 $Y=1.47 $X2=0 $Y2=0
cc_359 N_A_934_297#_c_447_n N_B_c_625_n 0.00325476f $X=8.075 $Y=1.57 $X2=0 $Y2=0
cc_360 N_A_934_297#_c_447_n N_B_M1014_g 0.0247105f $X=8.075 $Y=1.57 $X2=0 $Y2=0
cc_361 N_A_934_297#_c_436_n N_B_c_615_n 0.00179713f $X=6.585 $Y=1.202 $X2=0
+ $Y2=0
cc_362 N_A_934_297#_c_432_n N_B_c_616_n 0.0163648f $X=8.075 $Y=1.28 $X2=0 $Y2=0
cc_363 N_A_934_297#_c_436_n N_B_c_616_n 0.00773064f $X=6.585 $Y=1.202 $X2=0
+ $Y2=0
cc_364 N_A_934_297#_c_439_n N_B_c_616_n 3.11817e-19 $X=7.73 $Y=0.85 $X2=0 $Y2=0
cc_365 N_A_934_297#_c_443_n N_B_c_616_n 0.00175431f $X=7.875 $Y=0.85 $X2=0 $Y2=0
cc_366 N_A_934_297#_c_432_n N_B_c_617_n 0.00130403f $X=8.075 $Y=1.28 $X2=0 $Y2=0
cc_367 N_A_934_297#_c_439_n N_B_c_617_n 0.00735182f $X=7.73 $Y=0.85 $X2=0 $Y2=0
cc_368 N_A_934_297#_c_443_n N_B_c_617_n 0.0215777f $X=7.875 $Y=0.85 $X2=0 $Y2=0
cc_369 N_A_934_297#_M1011_g N_B_c_618_n 0.00773064f $X=6.61 $Y=0.455 $X2=0 $Y2=0
cc_370 N_A_934_297#_c_432_n N_B_c_618_n 0.00130645f $X=8.075 $Y=1.28 $X2=0 $Y2=0
cc_371 N_A_934_297#_c_434_n N_B_c_618_n 0.0134808f $X=8.105 $Y=0.945 $X2=0 $Y2=0
cc_372 N_A_934_297#_c_439_n N_B_c_618_n 0.00740121f $X=7.73 $Y=0.85 $X2=0 $Y2=0
cc_373 N_A_934_297#_c_442_n N_B_c_618_n 0.00141363f $X=7.875 $Y=0.85 $X2=0 $Y2=0
cc_374 N_A_934_297#_c_443_n N_B_c_618_n 0.00207916f $X=7.875 $Y=0.85 $X2=0 $Y2=0
cc_375 N_A_934_297#_c_432_n N_B_c_631_n 7.54224e-19 $X=8.075 $Y=1.28 $X2=0 $Y2=0
cc_376 N_A_934_297#_c_433_n N_B_c_631_n 0.00133812f $X=8.075 $Y=1.47 $X2=0 $Y2=0
cc_377 N_A_934_297#_c_447_n N_B_c_631_n 0.00617464f $X=8.075 $Y=1.57 $X2=0 $Y2=0
cc_378 N_A_934_297#_c_439_n N_B_c_631_n 0.00425555f $X=7.73 $Y=0.85 $X2=0 $Y2=0
cc_379 N_A_934_297#_c_442_n N_B_c_631_n 0.00240844f $X=7.875 $Y=0.85 $X2=0 $Y2=0
cc_380 N_A_934_297#_c_443_n N_B_c_631_n 0.0187117f $X=7.875 $Y=0.85 $X2=0 $Y2=0
cc_381 N_A_934_297#_c_432_n N_A_c_746_n 0.0181438f $X=8.075 $Y=1.28 $X2=-0.19
+ $Y2=-0.24
cc_382 N_A_934_297#_c_433_n N_A_c_746_n 0.0102542f $X=8.075 $Y=1.47 $X2=-0.19
+ $Y2=-0.24
cc_383 N_A_934_297#_c_447_n N_A_c_746_n 0.0315533f $X=8.075 $Y=1.57 $X2=-0.19
+ $Y2=-0.24
cc_384 N_A_934_297#_c_443_n N_A_c_746_n 6.56395e-19 $X=7.875 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_385 N_A_934_297#_c_434_n N_A_c_747_n 0.0188491f $X=8.105 $Y=0.945 $X2=0 $Y2=0
cc_386 N_A_934_297#_c_443_n N_A_c_747_n 2.42574e-19 $X=7.875 $Y=0.85 $X2=0 $Y2=0
cc_387 N_A_934_297#_c_432_n A 0.00153195f $X=8.075 $Y=1.28 $X2=0 $Y2=0
cc_388 N_A_934_297#_c_433_n A 0.00114147f $X=8.075 $Y=1.47 $X2=0 $Y2=0
cc_389 N_A_934_297#_c_443_n A 0.0138914f $X=7.875 $Y=0.85 $X2=0 $Y2=0
cc_390 N_A_934_297#_c_438_n N_A_1050_365#_M1009_s 8.50051e-19 $X=6.25 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_391 N_A_934_297#_c_450_n N_A_1050_365#_c_786_n 0.0199218f $X=4.97 $Y=1.58
+ $X2=0 $Y2=0
cc_392 N_A_934_297#_c_438_n N_A_1050_365#_c_786_n 0.0123662f $X=6.25 $Y=0.85
+ $X2=0 $Y2=0
cc_393 N_A_934_297#_c_454_p N_A_1050_365#_c_786_n 5.85147e-19 $X=5.06 $Y=0.85
+ $X2=0 $Y2=0
cc_394 N_A_934_297#_c_444_n N_A_1050_365#_c_786_n 0.0617744f $X=5.03 $Y=0.72
+ $X2=0 $Y2=0
cc_395 N_A_934_297#_c_447_n N_A_1050_365#_c_794_n 0.0030488f $X=8.075 $Y=1.57
+ $X2=0 $Y2=0
cc_396 N_A_934_297#_c_434_n N_A_1050_365#_c_788_n 0.00187335f $X=8.105 $Y=0.945
+ $X2=0 $Y2=0
cc_397 N_A_934_297#_c_442_n N_A_1050_365#_c_788_n 0.00537182f $X=7.875 $Y=0.85
+ $X2=0 $Y2=0
cc_398 N_A_934_297#_c_443_n N_A_1050_365#_c_788_n 0.00520032f $X=7.875 $Y=0.85
+ $X2=0 $Y2=0
cc_399 N_A_934_297#_M1011_g N_A_1050_365#_c_806_n 0.00614563f $X=6.61 $Y=0.455
+ $X2=0 $Y2=0
cc_400 N_A_934_297#_c_434_n N_A_1050_365#_c_806_n 0.00849993f $X=8.105 $Y=0.945
+ $X2=0 $Y2=0
cc_401 N_A_934_297#_c_437_n N_A_1050_365#_c_806_n 3.7129e-19 $X=6.372 $Y=0.995
+ $X2=0 $Y2=0
cc_402 N_A_934_297#_c_438_n N_A_1050_365#_c_806_n 0.0529545f $X=6.25 $Y=0.85
+ $X2=0 $Y2=0
cc_403 N_A_934_297#_c_439_n N_A_1050_365#_c_806_n 0.0955498f $X=7.73 $Y=0.85
+ $X2=0 $Y2=0
cc_404 N_A_934_297#_c_440_n N_A_1050_365#_c_806_n 0.0266362f $X=6.54 $Y=0.85
+ $X2=0 $Y2=0
cc_405 N_A_934_297#_c_441_n N_A_1050_365#_c_806_n 0.00318096f $X=6.395 $Y=0.85
+ $X2=0 $Y2=0
cc_406 N_A_934_297#_c_442_n N_A_1050_365#_c_806_n 0.0266136f $X=7.875 $Y=0.85
+ $X2=0 $Y2=0
cc_407 N_A_934_297#_c_443_n N_A_1050_365#_c_806_n 0.00508187f $X=7.875 $Y=0.85
+ $X2=0 $Y2=0
cc_408 N_A_934_297#_c_438_n N_A_1050_365#_c_790_n 0.0261136f $X=6.25 $Y=0.85
+ $X2=0 $Y2=0
cc_409 N_A_934_297#_c_444_n N_A_1050_365#_c_790_n 0.00677952f $X=5.03 $Y=0.72
+ $X2=0 $Y2=0
cc_410 N_A_934_297#_c_438_n N_A_1050_365#_c_791_n 0.00110106f $X=6.25 $Y=0.85
+ $X2=0 $Y2=0
cc_411 N_A_934_297#_c_444_n N_A_1050_365#_c_791_n 0.0118823f $X=5.03 $Y=0.72
+ $X2=0 $Y2=0
cc_412 N_A_934_297#_c_434_n N_A_1050_365#_c_819_n 0.00156626f $X=8.105 $Y=0.945
+ $X2=0 $Y2=0
cc_413 N_A_934_297#_c_434_n N_A_1050_365#_c_820_n 0.00809859f $X=8.105 $Y=0.945
+ $X2=0 $Y2=0
cc_414 N_A_934_297#_c_447_n N_VPWR_c_920_n 0.00129998f $X=8.075 $Y=1.57 $X2=0
+ $Y2=0
cc_415 N_A_934_297#_c_447_n N_VPWR_c_921_n 0.00434439f $X=8.075 $Y=1.57 $X2=0
+ $Y2=0
cc_416 N_A_934_297#_M1004_d N_VPWR_c_914_n 0.00359518f $X=4.67 $Y=1.485 $X2=0
+ $Y2=0
cc_417 N_A_934_297#_c_447_n N_VPWR_c_914_n 0.00650675f $X=8.075 $Y=1.57 $X2=0
+ $Y2=0
cc_418 N_A_934_297#_c_439_n N_A_465_325#_M1005_d 0.00140408f $X=7.73 $Y=0.85
+ $X2=0 $Y2=0
cc_419 N_A_934_297#_c_442_n N_A_465_325#_M1005_d 0.00214439f $X=7.875 $Y=0.85
+ $X2=0 $Y2=0
cc_420 N_A_934_297#_c_443_n N_A_465_325#_M1005_d 0.00513165f $X=7.875 $Y=0.85
+ $X2=0 $Y2=0
cc_421 N_A_934_297#_c_435_n N_A_465_325#_c_1070_n 0.00894291f $X=6.485 $Y=1.16
+ $X2=0 $Y2=0
cc_422 N_A_934_297#_c_437_n N_A_465_325#_c_1070_n 0.0270839f $X=6.372 $Y=0.995
+ $X2=0 $Y2=0
cc_423 N_A_934_297#_c_438_n N_A_465_325#_c_1070_n 5.63647e-19 $X=6.25 $Y=0.85
+ $X2=0 $Y2=0
cc_424 N_A_934_297#_c_445_n N_A_465_325#_c_1105_n 0.00385601f $X=6.585 $Y=1.41
+ $X2=0 $Y2=0
cc_425 N_A_934_297#_c_445_n N_A_465_325#_c_1071_n 0.0175866f $X=6.585 $Y=1.41
+ $X2=0 $Y2=0
cc_426 N_A_934_297#_c_435_n N_A_465_325#_c_1071_n 7.42472e-19 $X=6.485 $Y=1.16
+ $X2=0 $Y2=0
cc_427 N_A_934_297#_c_436_n N_A_465_325#_c_1071_n 9.0109e-19 $X=6.585 $Y=1.202
+ $X2=0 $Y2=0
cc_428 N_A_934_297#_c_437_n N_A_465_325#_c_1071_n 0.00152864f $X=6.372 $Y=0.995
+ $X2=0 $Y2=0
cc_429 N_A_934_297#_c_439_n N_A_465_325#_c_1071_n 0.00419686f $X=7.73 $Y=0.85
+ $X2=0 $Y2=0
cc_430 N_A_934_297#_c_440_n N_A_465_325#_c_1071_n 6.55203e-19 $X=6.54 $Y=0.85
+ $X2=0 $Y2=0
cc_431 N_A_934_297#_c_445_n N_A_465_325#_c_1067_n 0.00139259f $X=6.585 $Y=1.41
+ $X2=0 $Y2=0
cc_432 N_A_934_297#_M1011_g N_A_465_325#_c_1067_n 0.0164123f $X=6.61 $Y=0.455
+ $X2=0 $Y2=0
cc_433 N_A_934_297#_c_437_n N_A_465_325#_c_1067_n 0.0173003f $X=6.372 $Y=0.995
+ $X2=0 $Y2=0
cc_434 N_A_934_297#_c_439_n N_A_465_325#_c_1067_n 0.0173494f $X=7.73 $Y=0.85
+ $X2=0 $Y2=0
cc_435 N_A_934_297#_c_440_n N_A_465_325#_c_1067_n 0.00232583f $X=6.54 $Y=0.85
+ $X2=0 $Y2=0
cc_436 N_A_934_297#_c_441_n N_A_465_325#_c_1067_n 0.0185429f $X=6.395 $Y=0.85
+ $X2=0 $Y2=0
cc_437 N_A_934_297#_c_439_n N_A_465_325#_c_1118_n 0.00166303f $X=7.73 $Y=0.85
+ $X2=0 $Y2=0
cc_438 N_A_934_297#_c_434_n N_A_465_325#_c_1119_n 0.00333256f $X=8.105 $Y=0.945
+ $X2=0 $Y2=0
cc_439 N_A_934_297#_c_442_n N_A_465_325#_c_1119_n 3.55136e-19 $X=7.875 $Y=0.85
+ $X2=0 $Y2=0
cc_440 N_A_934_297#_c_443_n N_A_465_325#_c_1119_n 0.00528249f $X=7.875 $Y=0.85
+ $X2=0 $Y2=0
cc_441 N_A_934_297#_c_450_n N_A_465_325#_c_1073_n 0.0271848f $X=4.97 $Y=1.58
+ $X2=0 $Y2=0
cc_442 N_A_934_297#_c_437_n N_A_465_325#_c_1073_n 8.37577e-19 $X=6.372 $Y=0.995
+ $X2=0 $Y2=0
cc_443 N_A_934_297#_c_438_n N_A_465_325#_c_1073_n 0.0525503f $X=6.25 $Y=0.85
+ $X2=0 $Y2=0
cc_444 N_A_934_297#_c_454_p N_A_465_325#_c_1073_n 0.0124517f $X=5.06 $Y=0.85
+ $X2=0 $Y2=0
cc_445 N_A_934_297#_c_444_n N_A_465_325#_c_1073_n 0.00234408f $X=5.03 $Y=0.72
+ $X2=0 $Y2=0
cc_446 N_A_934_297#_c_445_n N_A_465_325#_c_1075_n 0.00348597f $X=6.585 $Y=1.41
+ $X2=0 $Y2=0
cc_447 N_A_934_297#_c_435_n N_A_465_325#_c_1075_n 0.00431105f $X=6.485 $Y=1.16
+ $X2=0 $Y2=0
cc_448 N_A_934_297#_c_436_n N_A_465_325#_c_1075_n 2.0806e-19 $X=6.585 $Y=1.202
+ $X2=0 $Y2=0
cc_449 N_A_934_297#_c_437_n N_A_465_325#_c_1075_n 0.00243787f $X=6.372 $Y=0.995
+ $X2=0 $Y2=0
cc_450 N_A_934_297#_c_440_n N_A_465_325#_c_1075_n 0.0154521f $X=6.54 $Y=0.85
+ $X2=0 $Y2=0
cc_451 N_A_934_297#_c_438_n N_A_483_49#_M1009_d 0.00139415f $X=6.25 $Y=0.85
+ $X2=0 $Y2=0
cc_452 N_A_934_297#_c_440_n N_A_483_49#_M1009_d 5.07779e-19 $X=6.54 $Y=0.85
+ $X2=0 $Y2=0
cc_453 N_A_934_297#_c_441_n N_A_483_49#_M1009_d 0.00662486f $X=6.395 $Y=0.85
+ $X2=0 $Y2=0
cc_454 N_A_934_297#_c_454_p N_A_483_49#_c_1215_n 0.00233211f $X=5.06 $Y=0.85
+ $X2=0 $Y2=0
cc_455 N_A_934_297#_c_444_n N_A_483_49#_c_1215_n 0.00358858f $X=5.03 $Y=0.72
+ $X2=0 $Y2=0
cc_456 N_A_934_297#_c_450_n N_A_483_49#_c_1216_n 0.0144112f $X=4.97 $Y=1.58
+ $X2=0 $Y2=0
cc_457 N_A_934_297#_c_444_n N_A_483_49#_c_1216_n 0.00935491f $X=5.03 $Y=0.72
+ $X2=0 $Y2=0
cc_458 N_A_934_297#_M1004_d N_A_483_49#_c_1224_n 0.0074794f $X=4.67 $Y=1.485
+ $X2=0 $Y2=0
cc_459 N_A_934_297#_c_450_n N_A_483_49#_c_1224_n 0.0314935f $X=4.97 $Y=1.58
+ $X2=0 $Y2=0
cc_460 N_A_934_297#_M1004_d N_A_483_49#_c_1225_n 0.00302314f $X=4.67 $Y=1.485
+ $X2=0 $Y2=0
cc_461 N_A_934_297#_M1004_d N_A_483_49#_c_1227_n 0.00298868f $X=4.67 $Y=1.485
+ $X2=0 $Y2=0
cc_462 N_A_934_297#_c_445_n N_A_483_49#_c_1217_n 0.00130504f $X=6.585 $Y=1.41
+ $X2=0 $Y2=0
cc_463 N_A_934_297#_c_435_n N_A_483_49#_c_1217_n 6.50075e-19 $X=6.485 $Y=1.16
+ $X2=0 $Y2=0
cc_464 N_A_934_297#_c_436_n N_A_483_49#_c_1217_n 3.92684e-19 $X=6.585 $Y=1.202
+ $X2=0 $Y2=0
cc_465 N_A_934_297#_c_437_n N_A_483_49#_c_1217_n 0.0156137f $X=6.372 $Y=0.995
+ $X2=0 $Y2=0
cc_466 N_A_934_297#_c_438_n N_A_483_49#_c_1217_n 0.00605333f $X=6.25 $Y=0.85
+ $X2=0 $Y2=0
cc_467 N_A_934_297#_c_440_n N_A_483_49#_c_1217_n 0.00104191f $X=6.54 $Y=0.85
+ $X2=0 $Y2=0
cc_468 N_A_934_297#_c_441_n N_A_483_49#_c_1217_n 0.00261896f $X=6.395 $Y=0.85
+ $X2=0 $Y2=0
cc_469 N_A_934_297#_c_445_n N_A_483_49#_c_1229_n 0.00258134f $X=6.585 $Y=1.41
+ $X2=0 $Y2=0
cc_470 N_A_934_297#_c_447_n N_A_483_49#_c_1229_n 0.00822576f $X=8.075 $Y=1.57
+ $X2=0 $Y2=0
cc_471 N_A_934_297#_M1011_g N_A_483_49#_c_1274_n 0.0022242f $X=6.61 $Y=0.455
+ $X2=0 $Y2=0
cc_472 N_A_934_297#_c_441_n N_A_483_49#_c_1274_n 0.00181204f $X=6.395 $Y=0.85
+ $X2=0 $Y2=0
cc_473 N_A_934_297#_c_444_n N_A_483_49#_c_1218_n 0.00622437f $X=5.03 $Y=0.72
+ $X2=0 $Y2=0
cc_474 N_A_934_297#_c_435_n N_A_483_49#_c_1219_n 2.22283e-19 $X=6.485 $Y=1.16
+ $X2=0 $Y2=0
cc_475 N_A_934_297#_c_437_n N_A_483_49#_c_1219_n 0.00265833f $X=6.372 $Y=0.995
+ $X2=0 $Y2=0
cc_476 N_A_934_297#_c_438_n N_A_483_49#_c_1219_n 0.0174471f $X=6.25 $Y=0.85
+ $X2=0 $Y2=0
cc_477 N_A_934_297#_c_440_n N_A_483_49#_c_1219_n 0.00133974f $X=6.54 $Y=0.85
+ $X2=0 $Y2=0
cc_478 N_A_934_297#_c_441_n N_A_483_49#_c_1219_n 0.0142042f $X=6.395 $Y=0.85
+ $X2=0 $Y2=0
cc_479 N_A_934_297#_c_439_n N_A_1335_297#_M1011_d 0.00166227f $X=7.73 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_480 N_A_934_297#_c_445_n N_A_1335_297#_c_1400_n 0.00686704f $X=6.585 $Y=1.41
+ $X2=0 $Y2=0
cc_481 N_A_934_297#_c_439_n N_A_1335_297#_c_1400_n 0.0181022f $X=7.73 $Y=0.85
+ $X2=0 $Y2=0
cc_482 N_A_934_297#_c_442_n N_A_1335_297#_c_1400_n 0.0020738f $X=7.875 $Y=0.85
+ $X2=0 $Y2=0
cc_483 N_A_934_297#_c_443_n N_A_1335_297#_c_1400_n 0.00517617f $X=7.875 $Y=0.85
+ $X2=0 $Y2=0
cc_484 N_A_934_297#_c_445_n N_A_1335_297#_c_1412_n 0.00431165f $X=6.585 $Y=1.41
+ $X2=0 $Y2=0
cc_485 N_A_934_297#_c_447_n N_A_1335_297#_c_1413_n 0.0163037f $X=8.075 $Y=1.57
+ $X2=0 $Y2=0
cc_486 N_A_934_297#_c_443_n N_A_1335_297#_c_1413_n 0.00184512f $X=7.875 $Y=0.85
+ $X2=0 $Y2=0
cc_487 N_A_934_297#_c_454_p N_VGND_c_1470_n 0.00369072f $X=5.06 $Y=0.85 $X2=0
+ $Y2=0
cc_488 N_A_934_297#_c_444_n N_VGND_c_1470_n 0.0242502f $X=5.03 $Y=0.72 $X2=0
+ $Y2=0
cc_489 N_A_934_297#_M1011_g N_VGND_c_1474_n 0.00575161f $X=6.61 $Y=0.455 $X2=0
+ $Y2=0
cc_490 N_A_934_297#_c_434_n N_VGND_c_1474_n 0.00585385f $X=8.105 $Y=0.945 $X2=0
+ $Y2=0
cc_491 N_A_934_297#_c_441_n N_VGND_c_1474_n 0.00348958f $X=6.395 $Y=0.85 $X2=0
+ $Y2=0
cc_492 N_A_934_297#_c_443_n N_VGND_c_1474_n 0.00104987f $X=7.875 $Y=0.85 $X2=0
+ $Y2=0
cc_493 N_A_934_297#_c_444_n N_VGND_c_1474_n 0.00893636f $X=5.03 $Y=0.72 $X2=0
+ $Y2=0
cc_494 N_A_934_297#_M1018_d N_VGND_c_1477_n 0.00234122f $X=4.845 $Y=0.235 $X2=0
+ $Y2=0
cc_495 N_A_934_297#_M1011_g N_VGND_c_1477_n 0.00669445f $X=6.61 $Y=0.455 $X2=0
+ $Y2=0
cc_496 N_A_934_297#_c_434_n N_VGND_c_1477_n 0.00635456f $X=8.105 $Y=0.945 $X2=0
+ $Y2=0
cc_497 N_A_934_297#_c_438_n N_VGND_c_1477_n 0.0112971f $X=6.25 $Y=0.85 $X2=0
+ $Y2=0
cc_498 N_A_934_297#_c_454_p N_VGND_c_1477_n 0.0148507f $X=5.06 $Y=0.85 $X2=0
+ $Y2=0
cc_499 N_A_934_297#_c_444_n N_VGND_c_1477_n 0.0045943f $X=5.03 $Y=0.72 $X2=0
+ $Y2=0
cc_500 N_B_c_619_n N_A_1050_365#_c_786_n 0.00363086f $X=4.58 $Y=1.41 $X2=0 $Y2=0
cc_501 N_B_M1018_g N_A_1050_365#_c_786_n 0.0010898f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_502 N_B_c_612_n N_A_1050_365#_c_786_n 0.0145436f $X=5.675 $Y=1.16 $X2=0 $Y2=0
cc_503 N_B_M1021_g N_A_1050_365#_c_786_n 0.00419529f $X=5.775 $Y=1.905 $X2=0
+ $Y2=0
cc_504 N_B_M1009_g N_A_1050_365#_c_786_n 0.00351927f $X=5.8 $Y=0.565 $X2=0 $Y2=0
cc_505 N_B_c_615_n N_A_1050_365#_c_786_n 0.00110014f $X=5.775 $Y=1.16 $X2=0
+ $Y2=0
cc_506 N_B_c_631_n N_A_1050_365#_c_794_n 0.0121884f $X=7.6 $Y=1.555 $X2=0 $Y2=0
cc_507 N_B_M1009_g N_A_1050_365#_c_806_n 0.00201366f $X=5.8 $Y=0.565 $X2=0 $Y2=0
cc_508 N_B_c_618_n N_A_1050_365#_c_806_n 0.00325658f $X=7.47 $Y=0.995 $X2=0
+ $Y2=0
cc_509 N_B_M1018_g N_A_1050_365#_c_790_n 4.07878e-19 $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_510 N_B_M1009_g N_A_1050_365#_c_790_n 9.1979e-19 $X=5.8 $Y=0.565 $X2=0 $Y2=0
cc_511 N_B_M1018_g N_A_1050_365#_c_791_n 0.00461232f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_512 N_B_c_612_n N_A_1050_365#_c_791_n 0.00313752f $X=5.675 $Y=1.16 $X2=0
+ $Y2=0
cc_513 N_B_c_619_n N_VPWR_c_919_n 0.0113699f $X=4.58 $Y=1.41 $X2=0 $Y2=0
cc_514 N_B_c_619_n N_VPWR_c_921_n 0.00455828f $X=4.58 $Y=1.41 $X2=0 $Y2=0
cc_515 N_B_c_623_n N_VPWR_c_921_n 0.0408109f $X=5.875 $Y=2.54 $X2=0 $Y2=0
cc_516 N_B_c_619_n N_VPWR_c_914_n 0.00656627f $X=4.58 $Y=1.41 $X2=0 $Y2=0
cc_517 N_B_c_622_n N_VPWR_c_914_n 0.0413158f $X=7.41 $Y=2.54 $X2=0 $Y2=0
cc_518 N_B_c_623_n N_VPWR_c_914_n 0.00712081f $X=5.875 $Y=2.54 $X2=0 $Y2=0
cc_519 N_B_c_613_n N_A_465_325#_c_1066_n 4.45781e-19 $X=4.845 $Y=1.16 $X2=0
+ $Y2=0
cc_520 N_B_M1021_g N_A_465_325#_c_1070_n 0.00146463f $X=5.775 $Y=1.905 $X2=0
+ $Y2=0
cc_521 N_B_M1021_g N_A_465_325#_c_1105_n 0.0044998f $X=5.775 $Y=1.905 $X2=0
+ $Y2=0
cc_522 N_B_c_618_n N_A_465_325#_c_1067_n 0.0026019f $X=7.47 $Y=0.995 $X2=0 $Y2=0
cc_523 N_B_c_616_n N_A_465_325#_c_1118_n 4.30216e-19 $X=7.465 $Y=1.16 $X2=0
+ $Y2=0
cc_524 N_B_c_617_n N_A_465_325#_c_1118_n 0.00294555f $X=7.465 $Y=1.16 $X2=0
+ $Y2=0
cc_525 N_B_c_618_n N_A_465_325#_c_1118_n 0.00498906f $X=7.47 $Y=0.995 $X2=0
+ $Y2=0
cc_526 N_B_c_616_n N_A_465_325#_c_1119_n 2.55873e-19 $X=7.465 $Y=1.16 $X2=0
+ $Y2=0
cc_527 N_B_c_618_n N_A_465_325#_c_1140_n 0.00521263f $X=7.47 $Y=0.995 $X2=0
+ $Y2=0
cc_528 N_B_c_619_n N_A_465_325#_c_1073_n 0.00484975f $X=4.58 $Y=1.41 $X2=0 $Y2=0
cc_529 N_B_c_612_n N_A_465_325#_c_1073_n 0.00478884f $X=5.675 $Y=1.16 $X2=0
+ $Y2=0
cc_530 N_B_c_613_n N_A_465_325#_c_1073_n 2.58451e-19 $X=4.845 $Y=1.16 $X2=0
+ $Y2=0
cc_531 N_B_M1021_g N_A_465_325#_c_1073_n 0.00508939f $X=5.775 $Y=1.905 $X2=0
+ $Y2=0
cc_532 N_B_c_615_n N_A_465_325#_c_1073_n 2.29578e-19 $X=5.775 $Y=1.16 $X2=0
+ $Y2=0
cc_533 N_B_M1021_g N_A_465_325#_c_1075_n 4.47596e-19 $X=5.775 $Y=1.905 $X2=0
+ $Y2=0
cc_534 N_B_c_631_n N_A_483_49#_M1014_d 0.00358887f $X=7.6 $Y=1.555 $X2=0 $Y2=0
cc_535 N_B_c_619_n N_A_483_49#_c_1220_n 0.00287893f $X=4.58 $Y=1.41 $X2=0 $Y2=0
cc_536 N_B_M1018_g N_A_483_49#_c_1215_n 0.00315172f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_537 N_B_c_619_n N_A_483_49#_c_1216_n 0.0127864f $X=4.58 $Y=1.41 $X2=0 $Y2=0
cc_538 N_B_c_613_n N_A_483_49#_c_1216_n 0.00534802f $X=4.845 $Y=1.16 $X2=0 $Y2=0
cc_539 N_B_c_619_n N_A_483_49#_c_1224_n 0.0174362f $X=4.58 $Y=1.41 $X2=0 $Y2=0
cc_540 N_B_c_619_n N_A_483_49#_c_1225_n 0.00608631f $X=4.58 $Y=1.41 $X2=0 $Y2=0
cc_541 N_B_M1021_g N_A_483_49#_c_1225_n 8.91158e-19 $X=5.775 $Y=1.905 $X2=0
+ $Y2=0
cc_542 N_B_c_619_n N_A_483_49#_c_1227_n 0.00366198f $X=4.58 $Y=1.41 $X2=0 $Y2=0
cc_543 N_B_c_612_n N_A_483_49#_c_1217_n 0.00364094f $X=5.675 $Y=1.16 $X2=0 $Y2=0
cc_544 N_B_M1021_g N_A_483_49#_c_1217_n 0.0315702f $X=5.775 $Y=1.905 $X2=0 $Y2=0
cc_545 N_B_M1009_g N_A_483_49#_c_1217_n 0.00650642f $X=5.8 $Y=0.565 $X2=0 $Y2=0
cc_546 N_B_c_615_n N_A_483_49#_c_1217_n 0.0104909f $X=5.775 $Y=1.16 $X2=0 $Y2=0
cc_547 N_B_M1021_g N_A_483_49#_c_1229_n 0.00851955f $X=5.775 $Y=1.905 $X2=0
+ $Y2=0
cc_548 N_B_c_622_n N_A_483_49#_c_1229_n 0.0365765f $X=7.41 $Y=2.54 $X2=0 $Y2=0
cc_549 N_B_c_623_n N_A_483_49#_c_1229_n 2.38151e-19 $X=5.875 $Y=2.54 $X2=0 $Y2=0
cc_550 N_B_M1014_g N_A_483_49#_c_1229_n 0.0102069f $X=7.51 $Y=1.965 $X2=0 $Y2=0
cc_551 N_B_M1009_g N_A_483_49#_c_1274_n 5.72667e-19 $X=5.8 $Y=0.565 $X2=0 $Y2=0
cc_552 N_B_M1018_g N_A_483_49#_c_1218_n 9.0609e-19 $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_553 N_B_c_613_n N_A_483_49#_c_1218_n 0.00386142f $X=4.845 $Y=1.16 $X2=0 $Y2=0
cc_554 N_B_M1009_g N_A_483_49#_c_1219_n 0.013823f $X=5.8 $Y=0.565 $X2=0 $Y2=0
cc_555 N_B_M1021_g N_A_483_49#_c_1232_n 0.00703655f $X=5.775 $Y=1.905 $X2=0
+ $Y2=0
cc_556 N_B_c_623_n N_A_483_49#_c_1232_n 2.51585e-19 $X=5.875 $Y=2.54 $X2=0 $Y2=0
cc_557 N_B_c_624_n N_A_1335_297#_c_1400_n 0.00160527f $X=7.51 $Y=1.47 $X2=0
+ $Y2=0
cc_558 N_B_M1014_g N_A_1335_297#_c_1400_n 0.00776798f $X=7.51 $Y=1.965 $X2=0
+ $Y2=0
cc_559 B N_A_1335_297#_c_1400_n 0.0174669f $X=7.51 $Y=1.445 $X2=0 $Y2=0
cc_560 N_B_c_617_n N_A_1335_297#_c_1400_n 0.0332296f $X=7.465 $Y=1.16 $X2=0
+ $Y2=0
cc_561 N_B_c_618_n N_A_1335_297#_c_1400_n 0.0104618f $X=7.47 $Y=0.995 $X2=0
+ $Y2=0
cc_562 N_B_M1014_g N_A_1335_297#_c_1413_n 0.0108967f $X=7.51 $Y=1.965 $X2=0
+ $Y2=0
cc_563 B N_A_1335_297#_c_1413_n 0.0094226f $X=7.51 $Y=1.445 $X2=0 $Y2=0
cc_564 N_B_c_616_n N_A_1335_297#_c_1413_n 0.00114355f $X=7.465 $Y=1.16 $X2=0
+ $Y2=0
cc_565 N_B_c_631_n N_A_1335_297#_c_1413_n 0.0154733f $X=7.6 $Y=1.555 $X2=0 $Y2=0
cc_566 N_B_M1018_g N_VGND_c_1470_n 0.00883459f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_567 N_B_c_613_n N_VGND_c_1470_n 0.00518895f $X=4.845 $Y=1.16 $X2=0 $Y2=0
cc_568 N_B_M1018_g N_VGND_c_1474_n 0.00560495f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_569 N_B_M1009_g N_VGND_c_1474_n 0.00427876f $X=5.8 $Y=0.565 $X2=0 $Y2=0
cc_570 N_B_c_618_n N_VGND_c_1474_n 0.00357877f $X=7.47 $Y=0.995 $X2=0 $Y2=0
cc_571 N_B_M1018_g N_VGND_c_1477_n 0.0110582f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_572 N_B_M1009_g N_VGND_c_1477_n 0.00718941f $X=5.8 $Y=0.565 $X2=0 $Y2=0
cc_573 N_B_c_618_n N_VGND_c_1477_n 0.00613199f $X=7.47 $Y=0.995 $X2=0 $Y2=0
cc_574 N_A_c_746_n N_A_1050_365#_c_784_n 0.0637929f $X=8.63 $Y=1.41 $X2=0 $Y2=0
cc_575 A N_A_1050_365#_c_784_n 8.4217e-19 $X=8.43 $Y=1.105 $X2=0 $Y2=0
cc_576 N_A_c_747_n N_A_1050_365#_c_785_n 0.0202318f $X=8.655 $Y=0.995 $X2=0
+ $Y2=0
cc_577 N_A_c_746_n N_A_1050_365#_c_794_n 0.0144336f $X=8.63 $Y=1.41 $X2=0 $Y2=0
cc_578 A N_A_1050_365#_c_794_n 0.0301432f $X=8.43 $Y=1.105 $X2=0 $Y2=0
cc_579 N_A_c_746_n N_A_1050_365#_c_787_n 5.76324e-19 $X=8.63 $Y=1.41 $X2=0 $Y2=0
cc_580 N_A_c_747_n N_A_1050_365#_c_787_n 0.0114592f $X=8.655 $Y=0.995 $X2=0
+ $Y2=0
cc_581 A N_A_1050_365#_c_787_n 0.0142387f $X=8.43 $Y=1.105 $X2=0 $Y2=0
cc_582 N_A_c_746_n N_A_1050_365#_c_788_n 0.00444032f $X=8.63 $Y=1.41 $X2=0 $Y2=0
cc_583 A N_A_1050_365#_c_788_n 0.0205785f $X=8.43 $Y=1.105 $X2=0 $Y2=0
cc_584 N_A_c_746_n N_A_1050_365#_c_789_n 7.33895e-19 $X=8.63 $Y=1.41 $X2=0 $Y2=0
cc_585 N_A_c_747_n N_A_1050_365#_c_789_n 0.00359979f $X=8.655 $Y=0.995 $X2=0
+ $Y2=0
cc_586 A N_A_1050_365#_c_789_n 0.021115f $X=8.43 $Y=1.105 $X2=0 $Y2=0
cc_587 N_A_c_746_n N_A_1050_365#_c_796_n 0.00336141f $X=8.63 $Y=1.41 $X2=0 $Y2=0
cc_588 A N_A_1050_365#_c_819_n 9.51454e-19 $X=8.43 $Y=1.105 $X2=0 $Y2=0
cc_589 N_A_c_746_n N_VPWR_c_920_n 0.0113659f $X=8.63 $Y=1.41 $X2=0 $Y2=0
cc_590 N_A_c_746_n N_VPWR_c_921_n 0.00309549f $X=8.63 $Y=1.41 $X2=0 $Y2=0
cc_591 N_A_c_746_n N_VPWR_c_914_n 0.00394227f $X=8.63 $Y=1.41 $X2=0 $Y2=0
cc_592 N_A_c_746_n N_A_483_49#_c_1229_n 0.00147672f $X=8.63 $Y=1.41 $X2=0 $Y2=0
cc_593 N_A_c_746_n N_A_1335_297#_c_1413_n 0.0136104f $X=8.63 $Y=1.41 $X2=0 $Y2=0
cc_594 N_A_c_746_n N_A_1335_297#_c_1406_n 3.68126e-19 $X=8.63 $Y=1.41 $X2=0
+ $Y2=0
cc_595 N_A_c_747_n N_VGND_c_1471_n 0.00276126f $X=8.655 $Y=0.995 $X2=0 $Y2=0
cc_596 N_A_c_747_n N_VGND_c_1474_n 0.00439206f $X=8.655 $Y=0.995 $X2=0 $Y2=0
cc_597 N_A_c_747_n N_VGND_c_1477_n 0.00642697f $X=8.655 $Y=0.995 $X2=0 $Y2=0
cc_598 N_A_1050_365#_c_794_n N_VPWR_M1000_d 0.00495492f $X=8.93 $Y=1.6 $X2=0
+ $Y2=0
cc_599 N_A_1050_365#_c_784_n N_VPWR_c_920_n 0.00837545f $X=9.1 $Y=1.41 $X2=0
+ $Y2=0
cc_600 N_A_1050_365#_c_784_n N_VPWR_c_923_n 0.00436183f $X=9.1 $Y=1.41 $X2=0
+ $Y2=0
cc_601 N_A_1050_365#_M1010_d N_VPWR_c_914_n 0.00402227f $X=8.165 $Y=1.645 $X2=0
+ $Y2=0
cc_602 N_A_1050_365#_c_784_n N_VPWR_c_914_n 0.00591185f $X=9.1 $Y=1.41 $X2=0
+ $Y2=0
cc_603 N_A_1050_365#_c_806_n N_A_465_325#_M1005_d 0.00432974f $X=8.24 $Y=0.51
+ $X2=0 $Y2=0
cc_604 N_A_1050_365#_c_806_n N_A_465_325#_c_1067_n 0.014738f $X=8.24 $Y=0.51
+ $X2=0 $Y2=0
cc_605 N_A_1050_365#_c_806_n N_A_465_325#_c_1118_n 0.00610486f $X=8.24 $Y=0.51
+ $X2=0 $Y2=0
cc_606 N_A_1050_365#_c_806_n N_A_465_325#_c_1119_n 0.00980954f $X=8.24 $Y=0.51
+ $X2=0 $Y2=0
cc_607 N_A_1050_365#_c_819_n N_A_465_325#_c_1119_n 0.0012274f $X=8.385 $Y=0.51
+ $X2=0 $Y2=0
cc_608 N_A_1050_365#_c_820_n N_A_465_325#_c_1119_n 0.00676874f $X=8.385 $Y=0.51
+ $X2=0 $Y2=0
cc_609 N_A_1050_365#_c_806_n N_A_465_325#_c_1140_n 0.0119237f $X=8.24 $Y=0.51
+ $X2=0 $Y2=0
cc_610 N_A_1050_365#_M1021_s N_A_465_325#_c_1073_n 0.00764502f $X=5.25 $Y=1.825
+ $X2=0 $Y2=0
cc_611 N_A_1050_365#_c_786_n N_A_465_325#_c_1073_n 0.0182772f $X=5.375 $Y=1.94
+ $X2=0 $Y2=0
cc_612 N_A_1050_365#_c_806_n N_A_483_49#_M1009_d 0.00606718f $X=8.24 $Y=0.51
+ $X2=0 $Y2=0
cc_613 N_A_1050_365#_c_786_n N_A_483_49#_c_1224_n 0.0138372f $X=5.375 $Y=1.94
+ $X2=0 $Y2=0
cc_614 N_A_1050_365#_c_786_n N_A_483_49#_c_1225_n 0.0028603f $X=5.375 $Y=1.94
+ $X2=0 $Y2=0
cc_615 N_A_1050_365#_M1021_s N_A_483_49#_c_1226_n 0.0104901f $X=5.25 $Y=1.825
+ $X2=0 $Y2=0
cc_616 N_A_1050_365#_c_786_n N_A_483_49#_c_1226_n 0.0128549f $X=5.375 $Y=1.94
+ $X2=0 $Y2=0
cc_617 N_A_1050_365#_c_786_n N_A_483_49#_c_1217_n 0.067594f $X=5.375 $Y=1.94
+ $X2=0 $Y2=0
cc_618 N_A_1050_365#_M1010_d N_A_483_49#_c_1229_n 0.00261136f $X=8.165 $Y=1.645
+ $X2=0 $Y2=0
cc_619 N_A_1050_365#_c_806_n N_A_483_49#_c_1274_n 0.0125744f $X=8.24 $Y=0.51
+ $X2=0 $Y2=0
cc_620 N_A_1050_365#_c_790_n N_A_483_49#_c_1274_n 0.00143452f $X=5.57 $Y=0.51
+ $X2=0 $Y2=0
cc_621 N_A_1050_365#_c_791_n N_A_483_49#_c_1274_n 0.00335094f $X=5.425 $Y=0.51
+ $X2=0 $Y2=0
cc_622 N_A_1050_365#_M1009_s N_A_483_49#_c_1219_n 0.00157756f $X=5.415 $Y=0.245
+ $X2=0 $Y2=0
cc_623 N_A_1050_365#_c_786_n N_A_483_49#_c_1219_n 0.0123139f $X=5.375 $Y=1.94
+ $X2=0 $Y2=0
cc_624 N_A_1050_365#_c_806_n N_A_483_49#_c_1219_n 0.00370418f $X=8.24 $Y=0.51
+ $X2=0 $Y2=0
cc_625 N_A_1050_365#_c_791_n N_A_483_49#_c_1219_n 0.0020377f $X=5.425 $Y=0.51
+ $X2=0 $Y2=0
cc_626 N_A_1050_365#_c_806_n N_A_1335_297#_M1011_d 0.00653094f $X=8.24 $Y=0.51
+ $X2=-0.19 $Y2=-0.24
cc_627 N_A_1050_365#_c_806_n N_A_1335_297#_c_1400_n 0.00162336f $X=8.24 $Y=0.51
+ $X2=0 $Y2=0
cc_628 N_A_1050_365#_c_784_n N_A_1335_297#_c_1401_n 0.0195627f $X=9.1 $Y=1.41
+ $X2=0 $Y2=0
cc_629 N_A_1050_365#_c_785_n N_A_1335_297#_c_1401_n 0.0097849f $X=9.125 $Y=0.995
+ $X2=0 $Y2=0
cc_630 N_A_1050_365#_c_794_n N_A_1335_297#_c_1401_n 0.0112214f $X=8.93 $Y=1.6
+ $X2=0 $Y2=0
cc_631 N_A_1050_365#_c_789_n N_A_1335_297#_c_1401_n 0.0381742f $X=9.015 $Y=1.325
+ $X2=0 $Y2=0
cc_632 N_A_1050_365#_c_796_n N_A_1335_297#_c_1401_n 0.00830381f $X=9.015
+ $Y=1.495 $X2=0 $Y2=0
cc_633 N_A_1050_365#_M1010_d N_A_1335_297#_c_1413_n 0.00774465f $X=8.165
+ $Y=1.645 $X2=0 $Y2=0
cc_634 N_A_1050_365#_c_784_n N_A_1335_297#_c_1413_n 0.00221849f $X=9.1 $Y=1.41
+ $X2=0 $Y2=0
cc_635 N_A_1050_365#_c_794_n N_A_1335_297#_c_1413_n 0.0353842f $X=8.93 $Y=1.6
+ $X2=0 $Y2=0
cc_636 N_A_1050_365#_c_784_n N_A_1335_297#_c_1406_n 0.0126341f $X=9.1 $Y=1.41
+ $X2=0 $Y2=0
cc_637 N_A_1050_365#_c_794_n N_A_1335_297#_c_1406_n 0.00653478f $X=8.93 $Y=1.6
+ $X2=0 $Y2=0
cc_638 N_A_1050_365#_c_789_n N_A_1335_297#_c_1406_n 0.00278512f $X=9.015
+ $Y=1.325 $X2=0 $Y2=0
cc_639 N_A_1050_365#_c_784_n N_A_1335_297#_c_1402_n 2.03932e-19 $X=9.1 $Y=1.41
+ $X2=0 $Y2=0
cc_640 N_A_1050_365#_c_787_n N_VGND_M1006_d 0.00147467f $X=8.93 $Y=0.82 $X2=0
+ $Y2=0
cc_641 N_A_1050_365#_c_789_n N_VGND_M1006_d 0.00108061f $X=9.015 $Y=1.325 $X2=0
+ $Y2=0
cc_642 N_A_1050_365#_c_785_n N_VGND_c_1471_n 0.00414899f $X=9.125 $Y=0.995 $X2=0
+ $Y2=0
cc_643 N_A_1050_365#_c_787_n N_VGND_c_1471_n 0.0111874f $X=8.93 $Y=0.82 $X2=0
+ $Y2=0
cc_644 N_A_1050_365#_c_789_n N_VGND_c_1471_n 0.00164729f $X=9.015 $Y=1.325 $X2=0
+ $Y2=0
cc_645 N_A_1050_365#_c_819_n N_VGND_c_1471_n 0.00112928f $X=8.385 $Y=0.51 $X2=0
+ $Y2=0
cc_646 N_A_1050_365#_c_787_n N_VGND_c_1474_n 0.00248202f $X=8.93 $Y=0.82 $X2=0
+ $Y2=0
cc_647 N_A_1050_365#_c_806_n N_VGND_c_1474_n 0.00575847f $X=8.24 $Y=0.51 $X2=0
+ $Y2=0
cc_648 N_A_1050_365#_c_790_n N_VGND_c_1474_n 2.49898e-19 $X=5.57 $Y=0.51 $X2=0
+ $Y2=0
cc_649 N_A_1050_365#_c_791_n N_VGND_c_1474_n 0.0254286f $X=5.425 $Y=0.51 $X2=0
+ $Y2=0
cc_650 N_A_1050_365#_c_819_n N_VGND_c_1474_n 3.63685e-19 $X=8.385 $Y=0.51 $X2=0
+ $Y2=0
cc_651 N_A_1050_365#_c_820_n N_VGND_c_1474_n 0.0149689f $X=8.385 $Y=0.51 $X2=0
+ $Y2=0
cc_652 N_A_1050_365#_c_785_n N_VGND_c_1476_n 0.00536613f $X=9.125 $Y=0.995 $X2=0
+ $Y2=0
cc_653 N_A_1050_365#_c_789_n N_VGND_c_1476_n 0.00182428f $X=9.015 $Y=1.325 $X2=0
+ $Y2=0
cc_654 N_A_1050_365#_M1015_d N_VGND_c_1477_n 0.00240207f $X=8.18 $Y=0.235 $X2=0
+ $Y2=0
cc_655 N_A_1050_365#_c_785_n N_VGND_c_1477_n 0.010284f $X=9.125 $Y=0.995 $X2=0
+ $Y2=0
cc_656 N_A_1050_365#_c_787_n N_VGND_c_1477_n 0.00552122f $X=8.93 $Y=0.82 $X2=0
+ $Y2=0
cc_657 N_A_1050_365#_c_789_n N_VGND_c_1477_n 0.00402105f $X=9.015 $Y=1.325 $X2=0
+ $Y2=0
cc_658 N_A_1050_365#_c_806_n N_VGND_c_1477_n 0.232956f $X=8.24 $Y=0.51 $X2=0
+ $Y2=0
cc_659 N_A_1050_365#_c_790_n N_VGND_c_1477_n 0.0285546f $X=5.57 $Y=0.51 $X2=0
+ $Y2=0
cc_660 N_A_1050_365#_c_791_n N_VGND_c_1477_n 0.00396297f $X=5.425 $Y=0.51 $X2=0
+ $Y2=0
cc_661 N_A_1050_365#_c_819_n N_VGND_c_1477_n 0.0285254f $X=8.385 $Y=0.51 $X2=0
+ $Y2=0
cc_662 N_A_1050_365#_c_820_n N_VGND_c_1477_n 0.0036194f $X=8.385 $Y=0.51 $X2=0
+ $Y2=0
cc_663 N_VPWR_c_914_n N_X_M1007_d 0.00255333f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_664 N_VPWR_c_916_n N_X_c_1025_n 0.0155816f $X=0.27 $Y=2.3 $X2=0 $Y2=0
cc_665 N_VPWR_c_917_n N_X_c_1025_n 0.0153803f $X=1.125 $Y=2.72 $X2=0 $Y2=0
cc_666 N_VPWR_c_918_n N_X_c_1025_n 0.0156188f $X=1.295 $Y=2.3 $X2=0 $Y2=0
cc_667 N_VPWR_c_914_n N_X_c_1025_n 0.00939158f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_668 N_VPWR_M1007_s N_X_c_1023_n 0.0250386f $X=0.145 $Y=1.485 $X2=0 $Y2=0
cc_669 N_VPWR_c_916_n N_X_c_1023_n 0.00378314f $X=0.27 $Y=2.3 $X2=0 $Y2=0
cc_670 N_VPWR_c_917_n N_X_c_1023_n 0.00316862f $X=1.125 $Y=2.72 $X2=0 $Y2=0
cc_671 N_VPWR_c_914_n N_X_c_1023_n 0.00606537f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_672 N_VPWR_c_922_n N_A_465_325#_c_1068_n 0.00407465f $X=4.18 $Y=2.72 $X2=0
+ $Y2=0
cc_673 N_VPWR_c_914_n N_A_465_325#_c_1068_n 0.0092333f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_674 N_VPWR_M1004_s N_A_465_325#_c_1073_n 0.00109947f $X=4.22 $Y=1.485 $X2=0
+ $Y2=0
cc_675 N_VPWR_c_914_n N_A_483_49#_M1014_d 0.00241089f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_676 N_VPWR_c_919_n N_A_483_49#_c_1221_n 0.00147971f $X=4.345 $Y=2.32 $X2=0
+ $Y2=0
cc_677 N_VPWR_c_922_n N_A_483_49#_c_1221_n 0.00296166f $X=4.18 $Y=2.72 $X2=0
+ $Y2=0
cc_678 N_VPWR_c_914_n N_A_483_49#_c_1221_n 0.00485654f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_679 N_VPWR_M1004_s N_A_483_49#_c_1216_n 0.00659923f $X=4.22 $Y=1.485 $X2=0
+ $Y2=0
cc_680 N_VPWR_M1004_s N_A_483_49#_c_1224_n 0.00155527f $X=4.22 $Y=1.485 $X2=0
+ $Y2=0
cc_681 N_VPWR_c_919_n N_A_483_49#_c_1224_n 0.00612755f $X=4.345 $Y=2.32 $X2=0
+ $Y2=0
cc_682 N_VPWR_c_921_n N_A_483_49#_c_1224_n 0.00666556f $X=8.65 $Y=2.72 $X2=0
+ $Y2=0
cc_683 N_VPWR_c_914_n N_A_483_49#_c_1224_n 0.0119497f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_684 N_VPWR_c_919_n N_A_483_49#_c_1225_n 0.00140976f $X=4.345 $Y=2.32 $X2=0
+ $Y2=0
cc_685 N_VPWR_c_921_n N_A_483_49#_c_1226_n 0.0294498f $X=8.65 $Y=2.72 $X2=0
+ $Y2=0
cc_686 N_VPWR_c_914_n N_A_483_49#_c_1226_n 0.0189426f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_687 N_VPWR_c_919_n N_A_483_49#_c_1227_n 0.00679194f $X=4.345 $Y=2.32 $X2=0
+ $Y2=0
cc_688 N_VPWR_c_921_n N_A_483_49#_c_1227_n 0.0105745f $X=8.65 $Y=2.72 $X2=0
+ $Y2=0
cc_689 N_VPWR_c_914_n N_A_483_49#_c_1227_n 0.00644066f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_690 N_VPWR_c_920_n N_A_483_49#_c_1229_n 0.00711003f $X=8.865 $Y=2.36 $X2=0
+ $Y2=0
cc_691 N_VPWR_c_921_n N_A_483_49#_c_1229_n 0.135241f $X=8.65 $Y=2.72 $X2=0 $Y2=0
cc_692 N_VPWR_c_914_n N_A_483_49#_c_1229_n 0.0814431f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_693 N_VPWR_c_919_n N_A_483_49#_c_1230_n 0.0142739f $X=4.345 $Y=2.32 $X2=0
+ $Y2=0
cc_694 N_VPWR_c_922_n N_A_483_49#_c_1230_n 0.0186431f $X=4.18 $Y=2.72 $X2=0
+ $Y2=0
cc_695 N_VPWR_c_914_n N_A_483_49#_c_1230_n 0.0145279f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_696 N_VPWR_M1004_s N_A_483_49#_c_1231_n 0.00243878f $X=4.22 $Y=1.485 $X2=0
+ $Y2=0
cc_697 N_VPWR_c_919_n N_A_483_49#_c_1231_n 0.0143988f $X=4.345 $Y=2.32 $X2=0
+ $Y2=0
cc_698 N_VPWR_c_914_n N_A_483_49#_c_1231_n 8.22076e-19 $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_699 N_VPWR_c_921_n N_A_483_49#_c_1232_n 0.010368f $X=8.65 $Y=2.72 $X2=0 $Y2=0
cc_700 N_VPWR_c_914_n N_A_483_49#_c_1232_n 0.00590105f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_701 N_VPWR_c_914_n N_A_1335_297#_M1020_d 0.00243468f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_702 N_VPWR_c_920_n N_A_1335_297#_c_1404_n 0.0121318f $X=8.865 $Y=2.36 $X2=0
+ $Y2=0
cc_703 N_VPWR_c_923_n N_A_1335_297#_c_1404_n 0.0197866f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_704 N_VPWR_c_914_n N_A_1335_297#_c_1404_n 0.0111058f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_705 N_VPWR_M1000_d N_A_1335_297#_c_1413_n 0.00390782f $X=8.72 $Y=1.485 $X2=0
+ $Y2=0
cc_706 N_VPWR_c_920_n N_A_1335_297#_c_1413_n 0.0198562f $X=8.865 $Y=2.36 $X2=0
+ $Y2=0
cc_707 N_VPWR_c_921_n N_A_1335_297#_c_1413_n 0.00692236f $X=8.65 $Y=2.72 $X2=0
+ $Y2=0
cc_708 N_VPWR_c_914_n N_A_1335_297#_c_1413_n 0.0149452f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_709 N_VPWR_c_923_n N_A_1335_297#_c_1406_n 0.00346082f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_710 N_VPWR_c_914_n N_A_1335_297#_c_1406_n 0.00566025f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_711 N_X_c_1021_n N_VGND_M1001_s 0.0101527f $X=0.805 $Y=0.66 $X2=-0.19
+ $Y2=-0.24
cc_712 N_X_c_1021_n N_VGND_c_1467_n 0.00311128f $X=0.805 $Y=0.66 $X2=0 $Y2=0
cc_713 N_X_c_1031_n N_VGND_c_1467_n 0.00660118f $X=0.765 $Y=0.56 $X2=0 $Y2=0
cc_714 N_X_c_1021_n N_VGND_c_1468_n 0.00361536f $X=0.805 $Y=0.66 $X2=0 $Y2=0
cc_715 N_X_c_1031_n N_VGND_c_1468_n 0.00913811f $X=0.765 $Y=0.56 $X2=0 $Y2=0
cc_716 N_X_M1001_d N_VGND_c_1477_n 0.00339635f $X=0.555 $Y=0.235 $X2=0 $Y2=0
cc_717 N_X_c_1021_n N_VGND_c_1477_n 0.00689139f $X=0.805 $Y=0.66 $X2=0 $Y2=0
cc_718 N_X_c_1031_n N_VGND_c_1477_n 0.00873403f $X=0.765 $Y=0.56 $X2=0 $Y2=0
cc_719 N_A_465_325#_c_1068_n N_A_483_49#_M1003_d 0.00645539f $X=3.5 $Y=1.98
+ $X2=0 $Y2=0
cc_720 N_A_465_325#_c_1088_n N_A_483_49#_M1003_d 0.00677252f $X=3.585 $Y=1.895
+ $X2=0 $Y2=0
cc_721 N_A_465_325#_c_1076_n N_A_483_49#_M1003_d 0.00697789f $X=3.83 $Y=1.535
+ $X2=0 $Y2=0
cc_722 N_A_465_325#_M1019_d N_A_483_49#_c_1213_n 0.00334341f $X=3.485 $Y=0.245
+ $X2=0 $Y2=0
cc_723 N_A_465_325#_c_1066_n N_A_483_49#_c_1213_n 0.0138308f $X=3.83 $Y=0.76
+ $X2=0 $Y2=0
cc_724 N_A_465_325#_M1019_d N_A_483_49#_c_1237_n 0.00348392f $X=3.485 $Y=0.245
+ $X2=0 $Y2=0
cc_725 N_A_465_325#_c_1066_n N_A_483_49#_c_1237_n 0.00439841f $X=3.83 $Y=0.76
+ $X2=0 $Y2=0
cc_726 N_A_465_325#_M1019_d N_A_483_49#_c_1214_n 0.0175141f $X=3.485 $Y=0.245
+ $X2=0 $Y2=0
cc_727 N_A_465_325#_c_1066_n N_A_483_49#_c_1214_n 0.0128008f $X=3.83 $Y=0.76
+ $X2=0 $Y2=0
cc_728 N_A_465_325#_M1019_d N_A_483_49#_c_1238_n 3.2099e-19 $X=3.485 $Y=0.245
+ $X2=0 $Y2=0
cc_729 N_A_465_325#_c_1073_n N_A_483_49#_c_1221_n 0.00437461f $X=6.25 $Y=1.53
+ $X2=0 $Y2=0
cc_730 N_A_465_325#_c_1074_n N_A_483_49#_c_1221_n 0.00277011f $X=4.09 $Y=1.53
+ $X2=0 $Y2=0
cc_731 N_A_465_325#_c_1076_n N_A_483_49#_c_1221_n 0.00125154f $X=3.83 $Y=1.535
+ $X2=0 $Y2=0
cc_732 N_A_465_325#_c_1068_n N_A_483_49#_c_1222_n 0.0153275f $X=3.5 $Y=1.98
+ $X2=0 $Y2=0
cc_733 N_A_465_325#_c_1074_n N_A_483_49#_c_1222_n 0.00119193f $X=4.09 $Y=1.53
+ $X2=0 $Y2=0
cc_734 N_A_465_325#_c_1076_n N_A_483_49#_c_1222_n 0.0114314f $X=3.83 $Y=1.535
+ $X2=0 $Y2=0
cc_735 N_A_465_325#_c_1066_n N_A_483_49#_c_1215_n 0.0327455f $X=3.83 $Y=0.76
+ $X2=0 $Y2=0
cc_736 N_A_465_325#_c_1088_n N_A_483_49#_c_1216_n 0.00649967f $X=3.585 $Y=1.895
+ $X2=0 $Y2=0
cc_737 N_A_465_325#_c_1066_n N_A_483_49#_c_1216_n 0.00891656f $X=3.83 $Y=0.76
+ $X2=0 $Y2=0
cc_738 N_A_465_325#_c_1073_n N_A_483_49#_c_1216_n 0.0161183f $X=6.25 $Y=1.53
+ $X2=0 $Y2=0
cc_739 N_A_465_325#_c_1074_n N_A_483_49#_c_1216_n 0.00275249f $X=4.09 $Y=1.53
+ $X2=0 $Y2=0
cc_740 N_A_465_325#_c_1076_n N_A_483_49#_c_1216_n 0.0233325f $X=3.83 $Y=1.535
+ $X2=0 $Y2=0
cc_741 N_A_465_325#_c_1073_n N_A_483_49#_c_1224_n 0.011487f $X=6.25 $Y=1.53
+ $X2=0 $Y2=0
cc_742 N_A_465_325#_c_1070_n N_A_483_49#_c_1217_n 0.00833378f $X=6.247 $Y=1.615
+ $X2=0 $Y2=0
cc_743 N_A_465_325#_c_1105_n N_A_483_49#_c_1217_n 0.0247324f $X=6.215 $Y=1.62
+ $X2=0 $Y2=0
cc_744 N_A_465_325#_c_1073_n N_A_483_49#_c_1217_n 0.0194987f $X=6.25 $Y=1.53
+ $X2=0 $Y2=0
cc_745 N_A_465_325#_c_1075_n N_A_483_49#_c_1217_n 0.00126802f $X=6.395 $Y=1.53
+ $X2=0 $Y2=0
cc_746 N_A_465_325#_M1021_d N_A_483_49#_c_1229_n 0.0094538f $X=5.865 $Y=1.485
+ $X2=0 $Y2=0
cc_747 N_A_465_325#_c_1105_n N_A_483_49#_c_1229_n 0.0238103f $X=6.215 $Y=1.62
+ $X2=0 $Y2=0
cc_748 N_A_465_325#_c_1071_n N_A_483_49#_c_1229_n 0.0100462f $X=6.7 $Y=1.53
+ $X2=0 $Y2=0
cc_749 N_A_465_325#_c_1067_n N_A_483_49#_c_1274_n 0.00250545f $X=6.785 $Y=1.445
+ $X2=0 $Y2=0
cc_750 N_A_465_325#_c_1068_n N_A_483_49#_c_1230_n 0.0049241f $X=3.5 $Y=1.98
+ $X2=0 $Y2=0
cc_751 N_A_465_325#_c_1074_n N_A_483_49#_c_1230_n 2.48159e-19 $X=4.09 $Y=1.53
+ $X2=0 $Y2=0
cc_752 N_A_465_325#_c_1076_n N_A_483_49#_c_1230_n 0.00535873f $X=3.83 $Y=1.535
+ $X2=0 $Y2=0
cc_753 N_A_465_325#_c_1066_n N_A_483_49#_c_1218_n 0.0132287f $X=3.83 $Y=0.76
+ $X2=0 $Y2=0
cc_754 N_A_465_325#_c_1073_n N_A_483_49#_c_1218_n 0.0052436f $X=6.25 $Y=1.53
+ $X2=0 $Y2=0
cc_755 N_A_465_325#_c_1074_n N_A_483_49#_c_1218_n 2.29009e-19 $X=4.09 $Y=1.53
+ $X2=0 $Y2=0
cc_756 N_A_465_325#_c_1070_n N_A_483_49#_c_1219_n 2.53366e-19 $X=6.247 $Y=1.615
+ $X2=0 $Y2=0
cc_757 N_A_465_325#_c_1073_n N_A_483_49#_c_1219_n 9.70582e-19 $X=6.25 $Y=1.53
+ $X2=0 $Y2=0
cc_758 N_A_465_325#_c_1067_n N_A_1335_297#_M1011_d 0.00729398f $X=6.785 $Y=1.445
+ $X2=-0.19 $Y2=-0.24
cc_759 N_A_465_325#_c_1199_p N_A_1335_297#_M1011_d 0.0024562f $X=6.87 $Y=0.34
+ $X2=-0.19 $Y2=-0.24
cc_760 N_A_465_325#_c_1140_n N_A_1335_297#_M1011_d 0.0107136f $X=7.38 $Y=0.36
+ $X2=-0.19 $Y2=-0.24
cc_761 N_A_465_325#_c_1071_n N_A_1335_297#_M1017_d 0.00444096f $X=6.7 $Y=1.53
+ $X2=0 $Y2=0
cc_762 N_A_465_325#_c_1105_n N_A_1335_297#_c_1400_n 0.00453141f $X=6.215 $Y=1.62
+ $X2=0 $Y2=0
cc_763 N_A_465_325#_c_1071_n N_A_1335_297#_c_1400_n 0.013519f $X=6.7 $Y=1.53
+ $X2=0 $Y2=0
cc_764 N_A_465_325#_c_1067_n N_A_1335_297#_c_1400_n 0.062318f $X=6.785 $Y=1.445
+ $X2=0 $Y2=0
cc_765 N_A_465_325#_c_1140_n N_A_1335_297#_c_1400_n 0.0106102f $X=7.38 $Y=0.36
+ $X2=0 $Y2=0
cc_766 N_A_465_325#_c_1075_n N_A_1335_297#_c_1400_n 0.00130235f $X=6.395 $Y=1.53
+ $X2=0 $Y2=0
cc_767 N_A_465_325#_c_1073_n N_VGND_c_1470_n 0.00558664f $X=6.25 $Y=1.53 $X2=0
+ $Y2=0
cc_768 N_A_465_325#_c_1199_p N_VGND_c_1474_n 0.0104913f $X=6.87 $Y=0.34 $X2=0
+ $Y2=0
cc_769 N_A_465_325#_c_1140_n N_VGND_c_1474_n 0.0617902f $X=7.38 $Y=0.36 $X2=0
+ $Y2=0
cc_770 N_A_465_325#_M1005_d N_VGND_c_1477_n 0.00231474f $X=7.48 $Y=0.245 $X2=0
+ $Y2=0
cc_771 N_A_465_325#_c_1199_p N_VGND_c_1477_n 0.00184693f $X=6.87 $Y=0.34 $X2=0
+ $Y2=0
cc_772 N_A_465_325#_c_1140_n N_VGND_c_1477_n 0.00974346f $X=7.38 $Y=0.36 $X2=0
+ $Y2=0
cc_773 N_A_483_49#_c_1229_n N_A_1335_297#_M1017_d 0.00563686f $X=7.83 $Y=2.36
+ $X2=0 $Y2=0
cc_774 N_A_483_49#_c_1229_n N_A_1335_297#_c_1412_n 0.0129278f $X=7.83 $Y=2.36
+ $X2=0 $Y2=0
cc_775 N_A_483_49#_M1014_d N_A_1335_297#_c_1413_n 0.00649554f $X=7.6 $Y=1.645
+ $X2=0 $Y2=0
cc_776 N_A_483_49#_c_1229_n N_A_1335_297#_c_1413_n 0.0533312f $X=7.83 $Y=2.36
+ $X2=0 $Y2=0
cc_777 N_A_483_49#_c_1214_n N_VGND_c_1470_n 0.0141317f $X=4.085 $Y=0.34 $X2=0
+ $Y2=0
cc_778 N_A_483_49#_c_1215_n N_VGND_c_1470_n 0.0321793f $X=4.17 $Y=1.035 $X2=0
+ $Y2=0
cc_779 N_A_483_49#_c_1213_n N_VGND_c_1472_n 0.00238811f $X=3.36 $Y=0.74 $X2=0
+ $Y2=0
cc_780 N_A_483_49#_c_1214_n N_VGND_c_1472_n 0.0445697f $X=4.085 $Y=0.34 $X2=0
+ $Y2=0
cc_781 N_A_483_49#_c_1238_n N_VGND_c_1472_n 0.0127275f $X=3.575 $Y=0.34 $X2=0
+ $Y2=0
cc_782 N_A_483_49#_c_1274_n N_VGND_c_1474_n 0.00800682f $X=6.01 $Y=0.545 $X2=0
+ $Y2=0
cc_783 N_A_483_49#_c_1219_n N_VGND_c_1474_n 0.0028353f $X=5.715 $Y=0.772 $X2=0
+ $Y2=0
cc_784 N_A_483_49#_c_1213_n N_VGND_c_1477_n 0.00647697f $X=3.36 $Y=0.74 $X2=0
+ $Y2=0
cc_785 N_A_483_49#_c_1214_n N_VGND_c_1477_n 0.0255342f $X=4.085 $Y=0.34 $X2=0
+ $Y2=0
cc_786 N_A_483_49#_c_1238_n N_VGND_c_1477_n 0.0076707f $X=3.575 $Y=0.34 $X2=0
+ $Y2=0
cc_787 N_A_483_49#_c_1274_n N_VGND_c_1477_n 0.0018012f $X=6.01 $Y=0.545 $X2=0
+ $Y2=0
cc_788 N_A_1335_297#_c_1402_n N_VGND_c_1476_n 0.0197872f $X=9.465 $Y=0.42 $X2=0
+ $Y2=0
cc_789 N_A_1335_297#_M1023_d N_VGND_c_1477_n 0.00379446f $X=9.2 $Y=0.235 $X2=0
+ $Y2=0
cc_790 N_A_1335_297#_c_1402_n N_VGND_c_1477_n 0.0113402f $X=9.465 $Y=0.42 $X2=0
+ $Y2=0
