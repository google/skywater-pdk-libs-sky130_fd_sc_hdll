* File: sky130_fd_sc_hdll__and3b_4.pxi.spice
* Created: Wed Sep  2 08:22:46 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND3B_4%A_98_199# N_A_98_199#_M1013_d
+ N_A_98_199#_M1011_d N_A_98_199#_c_71_n N_A_98_199#_M1005_g N_A_98_199#_c_72_n
+ N_A_98_199#_M1009_g N_A_98_199#_c_76_n N_A_98_199#_c_77_n N_A_98_199#_c_105_p
+ N_A_98_199#_c_73_n N_A_98_199#_c_74_n PM_SKY130_FD_SC_HDLL__AND3B_4%A_98_199#
x_PM_SKY130_FD_SC_HDLL__AND3B_4%B N_B_c_146_n N_B_M1015_g N_B_c_147_n
+ N_B_M1014_g B B PM_SKY130_FD_SC_HDLL__AND3B_4%B
x_PM_SKY130_FD_SC_HDLL__AND3B_4%C N_C_c_180_n N_C_M1000_g N_C_c_181_n
+ N_C_M1003_g C C PM_SKY130_FD_SC_HDLL__AND3B_4%C
x_PM_SKY130_FD_SC_HDLL__AND3B_4%A_56_297# N_A_56_297#_M1009_s
+ N_A_56_297#_M1005_s N_A_56_297#_M1015_d N_A_56_297#_c_219_n
+ N_A_56_297#_M1004_g N_A_56_297#_c_228_n N_A_56_297#_M1001_g
+ N_A_56_297#_c_220_n N_A_56_297#_M1006_g N_A_56_297#_c_229_n
+ N_A_56_297#_M1002_g N_A_56_297#_c_221_n N_A_56_297#_M1008_g
+ N_A_56_297#_c_230_n N_A_56_297#_M1007_g N_A_56_297#_c_231_n
+ N_A_56_297#_M1012_g N_A_56_297#_c_222_n N_A_56_297#_M1010_g
+ N_A_56_297#_c_243_n N_A_56_297#_c_245_n N_A_56_297#_c_272_n
+ N_A_56_297#_c_223_n N_A_56_297#_c_232_n N_A_56_297#_c_233_n
+ N_A_56_297#_c_224_n N_A_56_297#_c_234_n N_A_56_297#_c_225_n
+ N_A_56_297#_c_264_n N_A_56_297#_c_226_n N_A_56_297#_c_227_n
+ PM_SKY130_FD_SC_HDLL__AND3B_4%A_56_297#
x_PM_SKY130_FD_SC_HDLL__AND3B_4%A_N N_A_N_c_370_n N_A_N_c_371_n N_A_N_M1011_g
+ N_A_N_M1013_g A_N A_N N_A_N_c_368_n N_A_N_c_369_n
+ PM_SKY130_FD_SC_HDLL__AND3B_4%A_N
x_PM_SKY130_FD_SC_HDLL__AND3B_4%VPWR N_VPWR_M1005_d N_VPWR_M1003_d
+ N_VPWR_M1002_d N_VPWR_M1012_d N_VPWR_c_409_n VPWR N_VPWR_c_410_n
+ N_VPWR_c_411_n N_VPWR_c_412_n N_VPWR_c_413_n N_VPWR_c_414_n N_VPWR_c_408_n
+ N_VPWR_c_416_n N_VPWR_c_417_n N_VPWR_c_418_n N_VPWR_c_419_n
+ PM_SKY130_FD_SC_HDLL__AND3B_4%VPWR
x_PM_SKY130_FD_SC_HDLL__AND3B_4%X N_X_M1004_d N_X_M1008_d N_X_M1001_s
+ N_X_M1007_s N_X_c_480_n N_X_c_487_n N_X_c_522_p N_X_c_490_n X X
+ PM_SKY130_FD_SC_HDLL__AND3B_4%X
x_PM_SKY130_FD_SC_HDLL__AND3B_4%VGND N_VGND_M1000_d N_VGND_M1006_s
+ N_VGND_M1010_s N_VGND_c_538_n N_VGND_c_539_n VGND N_VGND_c_540_n
+ N_VGND_c_541_n N_VGND_c_542_n N_VGND_c_543_n N_VGND_c_544_n N_VGND_c_545_n
+ N_VGND_c_546_n N_VGND_c_547_n PM_SKY130_FD_SC_HDLL__AND3B_4%VGND
cc_1 VNB N_A_98_199#_c_71_n 0.0253064f $X=-0.19 $Y=-0.24 $X2=0.71 $Y2=1.41
cc_2 VNB N_A_98_199#_c_72_n 0.0209699f $X=-0.19 $Y=-0.24 $X2=0.735 $Y2=0.995
cc_3 VNB N_A_98_199#_c_73_n 0.0432846f $X=-0.19 $Y=-0.24 $X2=4.71 $Y2=0.59
cc_4 VNB N_A_98_199#_c_74_n 0.00262888f $X=-0.19 $Y=-0.24 $X2=0.772 $Y2=1.16
cc_5 VNB N_B_c_146_n 0.0284279f $X=-0.19 $Y=-0.24 $X2=4.44 $Y2=0.465
cc_6 VNB N_B_c_147_n 0.0172191f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB B 0.00112907f $X=-0.19 $Y=-0.24 $X2=0.71 $Y2=1.41
cc_8 VNB N_C_c_180_n 0.0178196f $X=-0.19 $Y=-0.24 $X2=4.44 $Y2=0.465
cc_9 VNB N_C_c_181_n 0.0244294f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB C 0.00307439f $X=-0.19 $Y=-0.24 $X2=0.71 $Y2=1.41
cc_11 VNB N_A_56_297#_c_219_n 0.0172296f $X=-0.19 $Y=-0.24 $X2=0.735 $Y2=0.995
cc_12 VNB N_A_56_297#_c_220_n 0.016944f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=1.99
cc_13 VNB N_A_56_297#_c_221_n 0.0175501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_56_297#_c_222_n 0.017072f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_56_297#_c_223_n 0.00134716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_56_297#_c_224_n 0.0257406f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_56_297#_c_225_n 0.0246451f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_56_297#_c_226_n 0.00187039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_56_297#_c_227_n 0.0744908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB A_N 0.00459272f $X=-0.19 $Y=-0.24 $X2=0.735 $Y2=0.56
cc_21 VNB N_A_N_c_368_n 0.0301547f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=1.99
cc_22 VNB N_A_N_c_369_n 0.0373928f $X=-0.19 $Y=-0.24 $X2=4.58 $Y2=2.02
cc_23 VNB N_VPWR_c_408_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB X 0.00379684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_538_n 0.00279285f $X=-0.19 $Y=-0.24 $X2=0.735 $Y2=0.56
cc_26 VNB N_VGND_c_539_n 0.00226353f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=1.99
cc_27 VNB N_VGND_c_540_n 0.0497091f $X=-0.19 $Y=-0.24 $X2=4.765 $Y2=0.59
cc_28 VNB N_VGND_c_541_n 0.0145554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_542_n 0.0141785f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_543_n 0.0268989f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_544_n 0.273648f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_545_n 0.00512961f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_546_n 0.00548421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_547_n 0.0109624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VPB N_A_98_199#_c_71_n 0.0332573f $X=-0.19 $Y=1.305 $X2=0.71 $Y2=1.41
cc_36 VPB N_A_98_199#_c_76_n 0.00184405f $X=-0.19 $Y=1.305 $X2=0.772 $Y2=1.875
cc_37 VPB N_A_98_199#_c_77_n 0.0132138f $X=-0.19 $Y=1.305 $X2=4.625 $Y2=1.99
cc_38 VPB N_A_98_199#_c_73_n 0.0287383f $X=-0.19 $Y=1.305 $X2=4.71 $Y2=0.59
cc_39 VPB N_A_98_199#_c_74_n 2.68624e-19 $X=-0.19 $Y=1.305 $X2=0.772 $Y2=1.16
cc_40 VPB N_B_c_146_n 0.0293691f $X=-0.19 $Y=1.305 $X2=4.44 $Y2=0.465
cc_41 VPB B 0.00238893f $X=-0.19 $Y=1.305 $X2=0.71 $Y2=1.41
cc_42 VPB N_C_c_181_n 0.027818f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB C 0.00207389f $X=-0.19 $Y=1.305 $X2=0.71 $Y2=1.41
cc_44 VPB N_A_56_297#_c_228_n 0.0171871f $X=-0.19 $Y=1.305 $X2=0.772 $Y2=1.325
cc_45 VPB N_A_56_297#_c_229_n 0.0159445f $X=-0.19 $Y=1.305 $X2=4.765 $Y2=1.875
cc_46 VPB N_A_56_297#_c_230_n 0.0161547f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.16
cc_47 VPB N_A_56_297#_c_231_n 0.0158529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_56_297#_c_232_n 0.00240942f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_56_297#_c_233_n 0.00549531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_56_297#_c_234_n 0.029929f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_56_297#_c_225_n 0.0094273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_56_297#_c_226_n 9.41933e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_56_297#_c_227_n 0.0477681f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_N_c_370_n 0.0147995f $X=-0.19 $Y=1.305 $X2=4.43 $Y2=1.725
cc_55 VPB N_A_N_c_371_n 0.00710238f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_N_M1011_g 0.0522965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB A_N 0.00714049f $X=-0.19 $Y=1.305 $X2=0.735 $Y2=0.56
cc_58 VPB N_A_N_c_368_n 0.00534359f $X=-0.19 $Y=1.305 $X2=0.865 $Y2=1.99
cc_59 VPB N_VPWR_c_409_n 0.00449519f $X=-0.19 $Y=1.305 $X2=4.625 $Y2=1.99
cc_60 VPB N_VPWR_c_410_n 0.0222531f $X=-0.19 $Y=1.305 $X2=4.765 $Y2=1.875
cc_61 VPB N_VPWR_c_411_n 0.0170074f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.16
cc_62 VPB N_VPWR_c_412_n 0.0157834f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.16
cc_63 VPB N_VPWR_c_413_n 0.013534f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_414_n 0.0266718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_408_n 0.0554546f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_416_n 0.00747677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_417_n 0.00631318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_418_n 0.00544833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_419_n 0.0111148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB X 0.00272265f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 N_A_98_199#_c_71_n N_B_c_146_n 0.0527705f $X=0.71 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_72 N_A_98_199#_c_76_n N_B_c_146_n 0.00805253f $X=0.772 $Y=1.875 $X2=-0.19
+ $Y2=-0.24
cc_73 N_A_98_199#_c_77_n N_B_c_146_n 0.0201362f $X=4.625 $Y=1.99 $X2=-0.19
+ $Y2=-0.24
cc_74 N_A_98_199#_c_74_n N_B_c_146_n 0.00192593f $X=0.772 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_75 N_A_98_199#_c_72_n N_B_c_147_n 0.0240304f $X=0.735 $Y=0.995 $X2=0 $Y2=0
cc_76 N_A_98_199#_c_71_n B 4.05619e-19 $X=0.71 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A_98_199#_c_72_n B 0.0034087f $X=0.735 $Y=0.995 $X2=0 $Y2=0
cc_78 N_A_98_199#_c_76_n B 0.00117064f $X=0.772 $Y=1.875 $X2=0 $Y2=0
cc_79 N_A_98_199#_c_77_n B 0.00757915f $X=4.625 $Y=1.99 $X2=0 $Y2=0
cc_80 N_A_98_199#_c_74_n B 0.0255387f $X=0.772 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_98_199#_c_77_n N_C_c_181_n 0.016768f $X=4.625 $Y=1.99 $X2=0 $Y2=0
cc_82 N_A_98_199#_c_77_n N_A_56_297#_M1015_d 0.00576854f $X=4.625 $Y=1.99 $X2=0
+ $Y2=0
cc_83 N_A_98_199#_c_77_n N_A_56_297#_c_228_n 0.0181557f $X=4.625 $Y=1.99 $X2=0
+ $Y2=0
cc_84 N_A_98_199#_c_77_n N_A_56_297#_c_229_n 0.0154813f $X=4.625 $Y=1.99 $X2=0
+ $Y2=0
cc_85 N_A_98_199#_c_77_n N_A_56_297#_c_230_n 0.0158783f $X=4.625 $Y=1.99 $X2=0
+ $Y2=0
cc_86 N_A_98_199#_c_77_n N_A_56_297#_c_231_n 0.016054f $X=4.625 $Y=1.99 $X2=0
+ $Y2=0
cc_87 N_A_98_199#_c_72_n N_A_56_297#_c_243_n 0.0110637f $X=0.735 $Y=0.995 $X2=0
+ $Y2=0
cc_88 N_A_98_199#_c_74_n N_A_56_297#_c_243_n 0.00648713f $X=0.772 $Y=1.16 $X2=0
+ $Y2=0
cc_89 N_A_98_199#_c_76_n N_A_56_297#_c_245_n 0.0060585f $X=0.772 $Y=1.875 $X2=0
+ $Y2=0
cc_90 N_A_98_199#_c_77_n N_A_56_297#_c_245_n 0.0493521f $X=4.625 $Y=1.99 $X2=0
+ $Y2=0
cc_91 N_A_98_199#_c_77_n N_A_56_297#_c_233_n 0.00320895f $X=4.625 $Y=1.99 $X2=0
+ $Y2=0
cc_92 N_A_98_199#_c_71_n N_A_56_297#_c_224_n 0.00422384f $X=0.71 $Y=1.41 $X2=0
+ $Y2=0
cc_93 N_A_98_199#_c_74_n N_A_56_297#_c_224_n 0.00576156f $X=0.772 $Y=1.16 $X2=0
+ $Y2=0
cc_94 N_A_98_199#_c_71_n N_A_56_297#_c_234_n 8.36899e-19 $X=0.71 $Y=1.41 $X2=0
+ $Y2=0
cc_95 N_A_98_199#_c_76_n N_A_56_297#_c_234_n 0.0284101f $X=0.772 $Y=1.875 $X2=0
+ $Y2=0
cc_96 N_A_98_199#_c_105_p N_A_56_297#_c_234_n 0.0190739f $X=0.865 $Y=1.99 $X2=0
+ $Y2=0
cc_97 N_A_98_199#_c_71_n N_A_56_297#_c_225_n 0.0102445f $X=0.71 $Y=1.41 $X2=0
+ $Y2=0
cc_98 N_A_98_199#_c_72_n N_A_56_297#_c_225_n 0.00246901f $X=0.735 $Y=0.995 $X2=0
+ $Y2=0
cc_99 N_A_98_199#_c_76_n N_A_56_297#_c_225_n 0.00562124f $X=0.772 $Y=1.875 $X2=0
+ $Y2=0
cc_100 N_A_98_199#_c_74_n N_A_56_297#_c_225_n 0.0252377f $X=0.772 $Y=1.16 $X2=0
+ $Y2=0
cc_101 N_A_98_199#_c_77_n N_A_56_297#_c_226_n 0.00136874f $X=4.625 $Y=1.99 $X2=0
+ $Y2=0
cc_102 N_A_98_199#_c_77_n N_A_56_297#_c_227_n 4.58134e-19 $X=4.625 $Y=1.99 $X2=0
+ $Y2=0
cc_103 N_A_98_199#_c_77_n N_A_N_M1011_g 0.0136855f $X=4.625 $Y=1.99 $X2=0 $Y2=0
cc_104 N_A_98_199#_c_73_n N_A_N_M1011_g 0.00563209f $X=4.71 $Y=0.59 $X2=0 $Y2=0
cc_105 N_A_98_199#_c_77_n A_N 0.0200364f $X=4.625 $Y=1.99 $X2=0 $Y2=0
cc_106 N_A_98_199#_c_73_n A_N 0.0772936f $X=4.71 $Y=0.59 $X2=0 $Y2=0
cc_107 N_A_98_199#_c_77_n N_A_N_c_368_n 0.00151809f $X=4.625 $Y=1.99 $X2=0 $Y2=0
cc_108 N_A_98_199#_c_73_n N_A_N_c_369_n 0.0138293f $X=4.71 $Y=0.59 $X2=0 $Y2=0
cc_109 N_A_98_199#_c_76_n N_VPWR_M1005_d 0.00525334f $X=0.772 $Y=1.875 $X2=-0.19
+ $Y2=-0.24
cc_110 N_A_98_199#_c_77_n N_VPWR_M1005_d 0.0112495f $X=4.625 $Y=1.99 $X2=-0.19
+ $Y2=-0.24
cc_111 N_A_98_199#_c_77_n N_VPWR_M1003_d 0.00573323f $X=4.625 $Y=1.99 $X2=0
+ $Y2=0
cc_112 N_A_98_199#_c_77_n N_VPWR_M1002_d 0.00351756f $X=4.625 $Y=1.99 $X2=0
+ $Y2=0
cc_113 N_A_98_199#_c_77_n N_VPWR_M1012_d 0.00959635f $X=4.625 $Y=1.99 $X2=0
+ $Y2=0
cc_114 N_A_98_199#_c_77_n N_VPWR_c_409_n 0.0201796f $X=4.625 $Y=1.99 $X2=0 $Y2=0
cc_115 N_A_98_199#_c_71_n N_VPWR_c_410_n 0.00374808f $X=0.71 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A_98_199#_c_105_p N_VPWR_c_410_n 9.32307e-19 $X=0.865 $Y=1.99 $X2=0
+ $Y2=0
cc_117 N_A_98_199#_c_77_n N_VPWR_c_411_n 0.0108985f $X=4.625 $Y=1.99 $X2=0 $Y2=0
cc_118 N_A_98_199#_c_77_n N_VPWR_c_412_n 0.0100642f $X=4.625 $Y=1.99 $X2=0 $Y2=0
cc_119 N_A_98_199#_c_77_n N_VPWR_c_413_n 0.00945518f $X=4.625 $Y=1.99 $X2=0
+ $Y2=0
cc_120 N_A_98_199#_c_77_n N_VPWR_c_414_n 0.0128423f $X=4.625 $Y=1.99 $X2=0 $Y2=0
cc_121 N_A_98_199#_c_71_n N_VPWR_c_408_n 0.0068124f $X=0.71 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A_98_199#_c_77_n N_VPWR_c_408_n 0.0769402f $X=4.625 $Y=1.99 $X2=0 $Y2=0
cc_123 N_A_98_199#_c_105_p N_VPWR_c_408_n 0.00197308f $X=0.865 $Y=1.99 $X2=0
+ $Y2=0
cc_124 N_A_98_199#_c_71_n N_VPWR_c_416_n 0.0210123f $X=0.71 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A_98_199#_c_77_n N_VPWR_c_416_n 0.0234941f $X=4.625 $Y=1.99 $X2=0 $Y2=0
cc_126 N_A_98_199#_c_105_p N_VPWR_c_416_n 0.00605084f $X=0.865 $Y=1.99 $X2=0
+ $Y2=0
cc_127 N_A_98_199#_c_77_n N_VPWR_c_418_n 0.0202591f $X=4.625 $Y=1.99 $X2=0 $Y2=0
cc_128 N_A_98_199#_c_77_n N_VPWR_c_419_n 0.0244949f $X=4.625 $Y=1.99 $X2=0 $Y2=0
cc_129 N_A_98_199#_c_77_n N_X_M1001_s 0.00527586f $X=4.625 $Y=1.99 $X2=0 $Y2=0
cc_130 N_A_98_199#_c_77_n N_X_M1007_s 0.0049956f $X=4.625 $Y=1.99 $X2=0 $Y2=0
cc_131 N_A_98_199#_c_77_n N_X_c_480_n 0.0901969f $X=4.625 $Y=1.99 $X2=0 $Y2=0
cc_132 N_A_98_199#_c_72_n N_VGND_c_540_n 0.00377907f $X=0.735 $Y=0.995 $X2=0
+ $Y2=0
cc_133 N_A_98_199#_c_73_n N_VGND_c_543_n 0.00953624f $X=4.71 $Y=0.59 $X2=0 $Y2=0
cc_134 N_A_98_199#_c_72_n N_VGND_c_544_n 0.00679642f $X=0.735 $Y=0.995 $X2=0
+ $Y2=0
cc_135 N_A_98_199#_c_73_n N_VGND_c_544_n 0.0097021f $X=4.71 $Y=0.59 $X2=0 $Y2=0
cc_136 N_A_98_199#_c_73_n N_VGND_c_547_n 8.57e-19 $X=4.71 $Y=0.59 $X2=0 $Y2=0
cc_137 N_B_c_147_n N_C_c_180_n 0.0392074f $X=1.31 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_138 B N_C_c_180_n 0.00104185f $X=1.115 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_139 N_B_c_146_n N_C_c_181_n 0.0607746f $X=1.285 $Y=1.41 $X2=0 $Y2=0
cc_140 B N_C_c_181_n 3.05157e-19 $X=1.115 $Y=0.765 $X2=0 $Y2=0
cc_141 N_B_c_146_n C 0.00246475f $X=1.285 $Y=1.41 $X2=0 $Y2=0
cc_142 B C 0.0234699f $X=1.115 $Y=0.765 $X2=0 $Y2=0
cc_143 N_B_c_146_n N_A_56_297#_c_243_n 0.0011458f $X=1.285 $Y=1.41 $X2=0 $Y2=0
cc_144 N_B_c_147_n N_A_56_297#_c_243_n 0.0141361f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_145 B N_A_56_297#_c_243_n 0.0139459f $X=1.115 $Y=0.765 $X2=0 $Y2=0
cc_146 N_B_c_146_n N_A_56_297#_c_245_n 0.00575564f $X=1.285 $Y=1.41 $X2=0 $Y2=0
cc_147 B N_A_56_297#_c_225_n 0.00418341f $X=1.115 $Y=0.765 $X2=0 $Y2=0
cc_148 N_B_c_147_n N_A_56_297#_c_264_n 0.00471288f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_149 B N_A_56_297#_c_264_n 0.00452801f $X=1.115 $Y=0.765 $X2=0 $Y2=0
cc_150 N_B_c_146_n N_VPWR_c_411_n 0.00408042f $X=1.285 $Y=1.41 $X2=0 $Y2=0
cc_151 N_B_c_146_n N_VPWR_c_408_n 0.00480655f $X=1.285 $Y=1.41 $X2=0 $Y2=0
cc_152 N_B_c_146_n N_VPWR_c_416_n 0.00960995f $X=1.285 $Y=1.41 $X2=0 $Y2=0
cc_153 B A_162_47# 0.00374423f $X=1.115 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_154 N_B_c_147_n N_VGND_c_540_n 0.00377907f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_155 N_B_c_147_n N_VGND_c_544_n 0.00576005f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_156 N_C_c_180_n N_A_56_297#_c_219_n 0.0180204f $X=1.74 $Y=0.995 $X2=0 $Y2=0
cc_157 N_C_c_181_n N_A_56_297#_c_228_n 0.0286034f $X=1.785 $Y=1.41 $X2=0 $Y2=0
cc_158 N_C_c_180_n N_A_56_297#_c_243_n 2.11302e-19 $X=1.74 $Y=0.995 $X2=0 $Y2=0
cc_159 C N_A_56_297#_c_243_n 0.00118191f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_160 N_C_c_181_n N_A_56_297#_c_245_n 0.0108499f $X=1.785 $Y=1.41 $X2=0 $Y2=0
cc_161 C N_A_56_297#_c_245_n 0.0244555f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_162 N_C_c_180_n N_A_56_297#_c_272_n 0.00982684f $X=1.74 $Y=0.995 $X2=0 $Y2=0
cc_163 N_C_c_181_n N_A_56_297#_c_272_n 0.00297013f $X=1.785 $Y=1.41 $X2=0 $Y2=0
cc_164 C N_A_56_297#_c_272_n 0.00932874f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_165 N_C_c_180_n N_A_56_297#_c_223_n 0.00415545f $X=1.74 $Y=0.995 $X2=0 $Y2=0
cc_166 N_C_c_181_n N_A_56_297#_c_223_n 2.04075e-19 $X=1.785 $Y=1.41 $X2=0 $Y2=0
cc_167 C N_A_56_297#_c_223_n 0.00183337f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_168 N_C_c_181_n N_A_56_297#_c_232_n 0.0037292f $X=1.785 $Y=1.41 $X2=0 $Y2=0
cc_169 N_C_c_180_n N_A_56_297#_c_264_n 0.00987605f $X=1.74 $Y=0.995 $X2=0 $Y2=0
cc_170 N_C_c_181_n N_A_56_297#_c_264_n 0.00142506f $X=1.785 $Y=1.41 $X2=0 $Y2=0
cc_171 C N_A_56_297#_c_264_n 0.0110981f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_172 N_C_c_181_n N_A_56_297#_c_226_n 0.00312675f $X=1.785 $Y=1.41 $X2=0 $Y2=0
cc_173 C N_A_56_297#_c_226_n 0.0272693f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_174 N_C_c_181_n N_A_56_297#_c_227_n 0.0138413f $X=1.785 $Y=1.41 $X2=0 $Y2=0
cc_175 C N_A_56_297#_c_227_n 2.94805e-19 $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_176 N_C_c_181_n N_VPWR_c_409_n 0.0018504f $X=1.785 $Y=1.41 $X2=0 $Y2=0
cc_177 N_C_c_181_n N_VPWR_c_411_n 0.00506535f $X=1.785 $Y=1.41 $X2=0 $Y2=0
cc_178 N_C_c_181_n N_VPWR_c_408_n 0.00685329f $X=1.785 $Y=1.41 $X2=0 $Y2=0
cc_179 N_C_c_181_n N_VPWR_c_416_n 0.00109403f $X=1.785 $Y=1.41 $X2=0 $Y2=0
cc_180 N_C_c_180_n N_VGND_c_538_n 0.00669741f $X=1.74 $Y=0.995 $X2=0 $Y2=0
cc_181 N_C_c_180_n N_VGND_c_540_n 0.00413138f $X=1.74 $Y=0.995 $X2=0 $Y2=0
cc_182 N_C_c_180_n N_VGND_c_544_n 0.00613194f $X=1.74 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_56_297#_c_231_n N_A_N_c_370_n 0.00742728f $X=3.78 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A_56_297#_c_227_n N_A_N_c_370_n 0.00273253f $X=3.78 $Y=1.202 $X2=0
+ $Y2=0
cc_185 N_A_56_297#_c_231_n N_A_N_M1011_g 0.0267933f $X=3.78 $Y=1.41 $X2=0 $Y2=0
cc_186 N_A_56_297#_c_231_n A_N 8.10763e-19 $X=3.78 $Y=1.41 $X2=0 $Y2=0
cc_187 N_A_56_297#_c_222_n A_N 0.00109674f $X=3.805 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_56_297#_c_227_n A_N 5.44194e-19 $X=3.78 $Y=1.202 $X2=0 $Y2=0
cc_189 N_A_56_297#_c_227_n N_A_N_c_368_n 0.0177884f $X=3.78 $Y=1.202 $X2=0 $Y2=0
cc_190 N_A_56_297#_c_222_n N_A_N_c_369_n 0.0185935f $X=3.805 $Y=0.995 $X2=0
+ $Y2=0
cc_191 N_A_56_297#_c_245_n N_VPWR_M1003_d 0.00801422f $X=2.035 $Y=1.61 $X2=0
+ $Y2=0
cc_192 N_A_56_297#_c_232_n N_VPWR_M1003_d 4.49409e-19 $X=2.12 $Y=1.525 $X2=0
+ $Y2=0
cc_193 N_A_56_297#_c_228_n N_VPWR_c_409_n 0.00176848f $X=2.34 $Y=1.41 $X2=0
+ $Y2=0
cc_194 N_A_56_297#_c_234_n N_VPWR_c_410_n 0.00843196f $X=0.425 $Y=1.66 $X2=0
+ $Y2=0
cc_195 N_A_56_297#_c_228_n N_VPWR_c_412_n 0.00506535f $X=2.34 $Y=1.41 $X2=0
+ $Y2=0
cc_196 N_A_56_297#_c_229_n N_VPWR_c_412_n 0.00295479f $X=2.83 $Y=1.41 $X2=0
+ $Y2=0
cc_197 N_A_56_297#_c_230_n N_VPWR_c_413_n 0.00450253f $X=3.3 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_56_297#_c_231_n N_VPWR_c_413_n 0.0032362f $X=3.78 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A_56_297#_M1005_s N_VPWR_c_408_n 0.00718714f $X=0.28 $Y=1.485 $X2=0
+ $Y2=0
cc_200 N_A_56_297#_M1015_d N_VPWR_c_408_n 0.00364536f $X=1.375 $Y=1.485 $X2=0
+ $Y2=0
cc_201 N_A_56_297#_c_228_n N_VPWR_c_408_n 0.00681939f $X=2.34 $Y=1.41 $X2=0
+ $Y2=0
cc_202 N_A_56_297#_c_229_n N_VPWR_c_408_n 0.00363171f $X=2.83 $Y=1.41 $X2=0
+ $Y2=0
cc_203 N_A_56_297#_c_230_n N_VPWR_c_408_n 0.00515739f $X=3.3 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A_56_297#_c_231_n N_VPWR_c_408_n 0.00388795f $X=3.78 $Y=1.41 $X2=0
+ $Y2=0
cc_205 N_A_56_297#_c_234_n N_VPWR_c_408_n 0.0114138f $X=0.425 $Y=1.66 $X2=0
+ $Y2=0
cc_206 N_A_56_297#_c_228_n N_VPWR_c_418_n 0.00116474f $X=2.34 $Y=1.41 $X2=0
+ $Y2=0
cc_207 N_A_56_297#_c_229_n N_VPWR_c_418_n 0.0112572f $X=2.83 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A_56_297#_c_230_n N_VPWR_c_418_n 0.00792658f $X=3.3 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A_56_297#_c_231_n N_VPWR_c_418_n 0.00101406f $X=3.78 $Y=1.41 $X2=0
+ $Y2=0
cc_210 N_A_56_297#_c_230_n N_VPWR_c_419_n 0.00111658f $X=3.3 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A_56_297#_c_231_n N_VPWR_c_419_n 0.0104876f $X=3.78 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A_56_297#_c_228_n N_X_c_480_n 0.00379252f $X=2.34 $Y=1.41 $X2=0 $Y2=0
cc_213 N_A_56_297#_c_229_n N_X_c_480_n 0.00987265f $X=2.83 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A_56_297#_c_230_n N_X_c_480_n 0.00987265f $X=3.3 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A_56_297#_c_231_n N_X_c_480_n 0.0069504f $X=3.78 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A_56_297#_c_233_n N_X_c_480_n 0.0654351f $X=3.185 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A_56_297#_c_227_n N_X_c_480_n 0.00864539f $X=3.78 $Y=1.202 $X2=0 $Y2=0
cc_218 N_A_56_297#_c_220_n N_X_c_487_n 0.0115023f $X=2.795 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A_56_297#_c_221_n N_X_c_487_n 0.0116545f $X=3.275 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_56_297#_c_227_n N_X_c_487_n 0.00347757f $X=3.78 $Y=1.202 $X2=0 $Y2=0
cc_221 N_A_56_297#_c_272_n N_X_c_490_n 0.0134127f $X=2.035 $Y=0.71 $X2=0 $Y2=0
cc_222 N_A_56_297#_c_223_n N_X_c_490_n 0.00254669f $X=2.15 $Y=1.02 $X2=0 $Y2=0
cc_223 N_A_56_297#_c_233_n N_X_c_490_n 0.0576898f $X=3.185 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A_56_297#_c_227_n N_X_c_490_n 0.00339319f $X=3.78 $Y=1.202 $X2=0 $Y2=0
cc_225 N_A_56_297#_c_222_n X 0.00804171f $X=3.805 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A_56_297#_c_227_n X 0.00576108f $X=3.78 $Y=1.202 $X2=0 $Y2=0
cc_227 N_A_56_297#_c_221_n X 0.00345508f $X=3.275 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A_56_297#_c_230_n X 0.00289445f $X=3.3 $Y=1.41 $X2=0 $Y2=0
cc_229 N_A_56_297#_c_231_n X 0.00366454f $X=3.78 $Y=1.41 $X2=0 $Y2=0
cc_230 N_A_56_297#_c_222_n X 0.00449489f $X=3.805 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A_56_297#_c_233_n X 0.0271998f $X=3.185 $Y=1.16 $X2=0 $Y2=0
cc_232 N_A_56_297#_c_227_n X 0.0257182f $X=3.78 $Y=1.202 $X2=0 $Y2=0
cc_233 N_A_56_297#_c_243_n A_162_47# 0.0117741f $X=1.52 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_234 N_A_56_297#_c_243_n A_277_47# 0.00372133f $X=1.52 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_235 N_A_56_297#_c_264_n A_277_47# 0.00526977f $X=1.61 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_236 N_A_56_297#_c_272_n N_VGND_M1000_d 0.00939743f $X=2.035 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_237 N_A_56_297#_c_223_n N_VGND_M1000_d 0.001056f $X=2.15 $Y=1.02 $X2=-0.19
+ $Y2=-0.24
cc_238 N_A_56_297#_c_219_n N_VGND_c_538_n 0.00791459f $X=2.315 $Y=0.995 $X2=0
+ $Y2=0
cc_239 N_A_56_297#_c_220_n N_VGND_c_538_n 0.00104968f $X=2.795 $Y=0.995 $X2=0
+ $Y2=0
cc_240 N_A_56_297#_c_272_n N_VGND_c_538_n 0.0217515f $X=2.035 $Y=0.71 $X2=0
+ $Y2=0
cc_241 N_A_56_297#_c_264_n N_VGND_c_538_n 0.00530357f $X=1.61 $Y=0.45 $X2=0
+ $Y2=0
cc_242 N_A_56_297#_c_219_n N_VGND_c_539_n 0.00106188f $X=2.315 $Y=0.995 $X2=0
+ $Y2=0
cc_243 N_A_56_297#_c_220_n N_VGND_c_539_n 0.0079907f $X=2.795 $Y=0.995 $X2=0
+ $Y2=0
cc_244 N_A_56_297#_c_221_n N_VGND_c_539_n 0.00177289f $X=3.275 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_A_56_297#_c_243_n N_VGND_c_540_n 0.0307579f $X=1.52 $Y=0.45 $X2=0 $Y2=0
cc_246 N_A_56_297#_c_272_n N_VGND_c_540_n 0.00363298f $X=2.035 $Y=0.71 $X2=0
+ $Y2=0
cc_247 N_A_56_297#_c_224_n N_VGND_c_540_n 0.0328451f $X=0.47 $Y=0.38 $X2=0 $Y2=0
cc_248 N_A_56_297#_c_264_n N_VGND_c_540_n 0.00623502f $X=1.61 $Y=0.45 $X2=0
+ $Y2=0
cc_249 N_A_56_297#_c_219_n N_VGND_c_541_n 0.00501198f $X=2.315 $Y=0.995 $X2=0
+ $Y2=0
cc_250 N_A_56_297#_c_220_n N_VGND_c_541_n 0.00351072f $X=2.795 $Y=0.995 $X2=0
+ $Y2=0
cc_251 N_A_56_297#_c_221_n N_VGND_c_542_n 0.00422112f $X=3.275 $Y=0.995 $X2=0
+ $Y2=0
cc_252 N_A_56_297#_c_222_n N_VGND_c_542_n 0.00210981f $X=3.805 $Y=0.995 $X2=0
+ $Y2=0
cc_253 N_A_56_297#_M1009_s N_VGND_c_544_n 0.00287355f $X=0.305 $Y=0.235 $X2=0
+ $Y2=0
cc_254 N_A_56_297#_c_219_n N_VGND_c_544_n 0.00853927f $X=2.315 $Y=0.995 $X2=0
+ $Y2=0
cc_255 N_A_56_297#_c_220_n N_VGND_c_544_n 0.00424612f $X=2.795 $Y=0.995 $X2=0
+ $Y2=0
cc_256 N_A_56_297#_c_221_n N_VGND_c_544_n 0.00592301f $X=3.275 $Y=0.995 $X2=0
+ $Y2=0
cc_257 N_A_56_297#_c_222_n N_VGND_c_544_n 0.00295961f $X=3.805 $Y=0.995 $X2=0
+ $Y2=0
cc_258 N_A_56_297#_c_243_n N_VGND_c_544_n 0.0294947f $X=1.52 $Y=0.45 $X2=0 $Y2=0
cc_259 N_A_56_297#_c_272_n N_VGND_c_544_n 0.00792525f $X=2.035 $Y=0.71 $X2=0
+ $Y2=0
cc_260 N_A_56_297#_c_224_n N_VGND_c_544_n 0.0185454f $X=0.47 $Y=0.38 $X2=0 $Y2=0
cc_261 N_A_56_297#_c_264_n N_VGND_c_544_n 0.00624139f $X=1.61 $Y=0.45 $X2=0
+ $Y2=0
cc_262 N_A_56_297#_c_221_n N_VGND_c_547_n 5.24562e-19 $X=3.275 $Y=0.995 $X2=0
+ $Y2=0
cc_263 N_A_56_297#_c_222_n N_VGND_c_547_n 0.00963409f $X=3.805 $Y=0.995 $X2=0
+ $Y2=0
cc_264 N_A_N_M1011_g N_VPWR_c_414_n 0.00559072f $X=4.34 $Y=1.935 $X2=0 $Y2=0
cc_265 N_A_N_M1011_g N_VPWR_c_408_n 0.00851485f $X=4.34 $Y=1.935 $X2=0 $Y2=0
cc_266 N_A_N_M1011_g N_VPWR_c_419_n 0.00915693f $X=4.34 $Y=1.935 $X2=0 $Y2=0
cc_267 N_A_N_c_370_n N_X_c_480_n 4.09535e-19 $X=4.34 $Y=1.55 $X2=0 $Y2=0
cc_268 A_N N_X_c_480_n 0.0145986f $X=4.275 $Y=1.105 $X2=0 $Y2=0
cc_269 A_N X 0.0194104f $X=4.275 $Y=1.105 $X2=0 $Y2=0
cc_270 N_A_N_c_369_n X 7.5205e-19 $X=4.277 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A_N_c_370_n X 6.82363e-19 $X=4.34 $Y=1.55 $X2=0 $Y2=0
cc_272 A_N X 0.0563855f $X=4.275 $Y=1.105 $X2=0 $Y2=0
cc_273 N_A_N_c_368_n X 0.00222884f $X=4.25 $Y=1.16 $X2=0 $Y2=0
cc_274 N_A_N_c_369_n X 4.47201e-19 $X=4.277 $Y=0.995 $X2=0 $Y2=0
cc_275 A_N N_VGND_M1010_s 0.00344287f $X=4.275 $Y=1.105 $X2=0 $Y2=0
cc_276 A_N N_VGND_c_543_n 0.00452574f $X=4.275 $Y=1.105 $X2=0 $Y2=0
cc_277 N_A_N_c_369_n N_VGND_c_543_n 0.00397697f $X=4.277 $Y=0.995 $X2=0 $Y2=0
cc_278 A_N N_VGND_c_544_n 0.00758681f $X=4.275 $Y=1.105 $X2=0 $Y2=0
cc_279 N_A_N_c_369_n N_VGND_c_544_n 0.00667499f $X=4.277 $Y=0.995 $X2=0 $Y2=0
cc_280 A_N N_VGND_c_547_n 0.00153732f $X=4.275 $Y=1.105 $X2=0 $Y2=0
cc_281 N_A_N_c_368_n N_VGND_c_547_n 0.00153163f $X=4.25 $Y=1.16 $X2=0 $Y2=0
cc_282 N_A_N_c_369_n N_VGND_c_547_n 0.00760021f $X=4.277 $Y=0.995 $X2=0 $Y2=0
cc_283 N_VPWR_c_408_n N_X_M1001_s 0.00353144f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_284 N_VPWR_c_408_n N_X_M1007_s 0.00341753f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_285 N_VPWR_M1002_d N_X_c_480_n 0.00340229f $X=2.92 $Y=1.485 $X2=0 $Y2=0
cc_286 N_VPWR_M1012_d N_X_c_480_n 0.00226774f $X=3.87 $Y=1.485 $X2=0 $Y2=0
cc_287 N_VPWR_M1012_d X 4.33671e-19 $X=3.87 $Y=1.485 $X2=0 $Y2=0
cc_288 N_X_c_487_n N_VGND_M1006_s 0.00421224f $X=3.365 $Y=0.73 $X2=0 $Y2=0
cc_289 X N_VGND_M1010_s 0.00271653f $X=3.715 $Y=0.765 $X2=0 $Y2=0
cc_290 X N_VGND_M1010_s 3.52146e-19 $X=3.805 $Y=0.85 $X2=0 $Y2=0
cc_291 N_X_c_487_n N_VGND_c_539_n 0.0183972f $X=3.365 $Y=0.73 $X2=0 $Y2=0
cc_292 N_X_c_487_n N_VGND_c_541_n 0.00263122f $X=3.365 $Y=0.73 $X2=0 $Y2=0
cc_293 N_X_c_490_n N_VGND_c_541_n 0.00449666f $X=2.675 $Y=0.68 $X2=0 $Y2=0
cc_294 N_X_c_487_n N_VGND_c_542_n 0.00281024f $X=3.365 $Y=0.73 $X2=0 $Y2=0
cc_295 N_X_c_522_p N_VGND_c_542_n 0.0172992f $X=3.54 $Y=0.42 $X2=0 $Y2=0
cc_296 X N_VGND_c_542_n 0.00275941f $X=3.715 $Y=0.765 $X2=0 $Y2=0
cc_297 N_X_M1004_d N_VGND_c_544_n 0.00648119f $X=2.39 $Y=0.235 $X2=0 $Y2=0
cc_298 N_X_M1008_d N_VGND_c_544_n 0.00341057f $X=3.35 $Y=0.235 $X2=0 $Y2=0
cc_299 N_X_c_487_n N_VGND_c_544_n 0.0100686f $X=3.365 $Y=0.73 $X2=0 $Y2=0
cc_300 N_X_c_522_p N_VGND_c_544_n 0.0102921f $X=3.54 $Y=0.42 $X2=0 $Y2=0
cc_301 N_X_c_490_n N_VGND_c_544_n 0.00604783f $X=2.675 $Y=0.68 $X2=0 $Y2=0
cc_302 X N_VGND_c_544_n 0.00574715f $X=3.715 $Y=0.765 $X2=0 $Y2=0
cc_303 N_X_c_522_p N_VGND_c_547_n 0.0146794f $X=3.54 $Y=0.42 $X2=0 $Y2=0
cc_304 X N_VGND_c_547_n 0.0106295f $X=3.715 $Y=0.765 $X2=0 $Y2=0
cc_305 A_162_47# N_VGND_c_544_n 0.00359325f $X=0.81 $Y=0.235 $X2=0 $Y2=0
cc_306 A_277_47# N_VGND_c_544_n 0.00235072f $X=1.385 $Y=0.235 $X2=1.545 $Y2=1.61
