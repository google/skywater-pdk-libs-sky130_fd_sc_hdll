* File: sky130_fd_sc_hdll__clkinv_8.pxi.spice
* Created: Wed Sep  2 08:26:36 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKINV_8%A N_A_c_101_n N_A_M1001_g N_A_c_102_n
+ N_A_M1002_g N_A_c_103_n N_A_M1003_g N_A_M1000_g N_A_c_104_n N_A_M1006_g
+ N_A_M1004_g N_A_c_105_n N_A_M1008_g N_A_M1005_g N_A_c_106_n N_A_M1009_g
+ N_A_M1007_g N_A_c_107_n N_A_M1011_g N_A_M1010_g N_A_c_108_n N_A_M1013_g
+ N_A_M1012_g N_A_c_109_n N_A_M1014_g N_A_M1015_g N_A_c_110_n N_A_M1016_g
+ N_A_M1019_g N_A_c_111_n N_A_M1017_g N_A_c_112_n N_A_M1018_g A A A A A A A A A
+ N_A_c_100_n N_A_c_152_p A A A A A A A A A PM_SKY130_FD_SC_HDLL__CLKINV_8%A
x_PM_SKY130_FD_SC_HDLL__CLKINV_8%VPWR N_VPWR_M1001_d N_VPWR_M1002_d
+ N_VPWR_M1006_d N_VPWR_M1009_d N_VPWR_M1013_d N_VPWR_M1016_d N_VPWR_M1018_d
+ N_VPWR_c_263_n N_VPWR_c_264_n N_VPWR_c_265_n N_VPWR_c_266_n N_VPWR_c_267_n
+ N_VPWR_c_268_n N_VPWR_c_269_n N_VPWR_c_270_n N_VPWR_c_271_n N_VPWR_c_272_n
+ N_VPWR_c_273_n N_VPWR_c_274_n N_VPWR_c_275_n N_VPWR_c_276_n N_VPWR_c_277_n
+ VPWR N_VPWR_c_278_n N_VPWR_c_279_n N_VPWR_c_280_n N_VPWR_c_281_n
+ N_VPWR_c_282_n N_VPWR_c_262_n PM_SKY130_FD_SC_HDLL__CLKINV_8%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKINV_8%Y N_Y_M1000_s N_Y_M1005_s N_Y_M1010_s
+ N_Y_M1015_s N_Y_M1001_s N_Y_M1003_s N_Y_M1008_s N_Y_M1011_s N_Y_M1014_s
+ N_Y_M1017_s N_Y_c_356_n N_Y_c_357_n N_Y_c_358_n N_Y_c_370_n N_Y_c_371_n
+ N_Y_c_473_n N_Y_c_372_n N_Y_c_477_n N_Y_c_359_n N_Y_c_373_n N_Y_c_360_n
+ N_Y_c_481_n N_Y_c_361_n N_Y_c_374_n N_Y_c_362_n N_Y_c_485_n N_Y_c_363_n
+ N_Y_c_375_n N_Y_c_364_n N_Y_c_489_n N_Y_c_365_n N_Y_c_376_n N_Y_c_366_n
+ N_Y_c_493_n N_Y_c_377_n N_Y_c_378_n N_Y_c_379_n N_Y_c_444_n N_Y_c_380_n
+ N_Y_c_448_n N_Y_c_381_n N_Y_c_452_n N_Y_c_382_n N_Y_c_456_n N_Y_c_383_n Y Y Y
+ N_Y_c_368_n N_Y_c_385_n PM_SKY130_FD_SC_HDLL__CLKINV_8%Y
x_PM_SKY130_FD_SC_HDLL__CLKINV_8%VGND N_VGND_M1000_d N_VGND_M1004_d
+ N_VGND_M1007_d N_VGND_M1012_d N_VGND_M1019_d N_VGND_c_541_n N_VGND_c_542_n
+ N_VGND_c_543_n N_VGND_c_544_n N_VGND_c_545_n N_VGND_c_546_n N_VGND_c_547_n
+ N_VGND_c_548_n N_VGND_c_549_n N_VGND_c_550_n N_VGND_c_551_n VGND
+ N_VGND_c_552_n N_VGND_c_553_n N_VGND_c_554_n N_VGND_c_555_n N_VGND_c_556_n
+ N_VGND_c_557_n PM_SKY130_FD_SC_HDLL__CLKINV_8%VGND
cc_1 VNB N_A_M1000_g 0.0228043f $X=-0.19 $Y=-0.24 $X2=1.515 $Y2=0.445
cc_2 VNB N_A_M1004_g 0.0186127f $X=-0.19 $Y=-0.24 $X2=1.995 $Y2=0.445
cc_3 VNB N_A_M1005_g 0.0184098f $X=-0.19 $Y=-0.24 $X2=2.475 $Y2=0.445
cc_4 VNB N_A_M1007_g 0.0186127f $X=-0.19 $Y=-0.24 $X2=2.955 $Y2=0.445
cc_5 VNB N_A_M1010_g 0.0186255f $X=-0.19 $Y=-0.24 $X2=3.435 $Y2=0.445
cc_6 VNB N_A_M1012_g 0.0193943f $X=-0.19 $Y=-0.24 $X2=3.965 $Y2=0.445
cc_7 VNB N_A_M1015_g 0.0193943f $X=-0.19 $Y=-0.24 $X2=4.495 $Y2=0.445
cc_8 VNB N_A_M1019_g 0.0232992f $X=-0.19 $Y=-0.24 $X2=5.025 $Y2=0.445
cc_9 VNB N_A_c_100_n 0.402315f $X=-0.19 $Y=-0.24 $X2=5.35 $Y2=1.16
cc_10 VNB N_VPWR_c_262_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.11
cc_11 VNB N_Y_c_356_n 0.0204297f $X=-0.19 $Y=-0.24 $X2=2.955 $Y2=0.445
cc_12 VNB N_Y_c_357_n 0.0171399f $X=-0.19 $Y=-0.24 $X2=2.955 $Y2=0.445
cc_13 VNB N_Y_c_358_n 0.00997812f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_Y_c_359_n 7.13037e-19 $X=-0.19 $Y=-0.24 $X2=4.31 $Y2=1.41
cc_15 VNB N_Y_c_360_n 0.00481263f $X=-0.19 $Y=-0.24 $X2=4.495 $Y2=0.445
cc_16 VNB N_Y_c_361_n 7.13037e-19 $X=-0.19 $Y=-0.24 $X2=5.025 $Y2=0.445
cc_17 VNB N_Y_c_362_n 0.00481263f $X=-0.19 $Y=-0.24 $X2=5.35 $Y2=1.985
cc_18 VNB N_Y_c_363_n 7.27967e-19 $X=-0.19 $Y=-0.24 $X2=2.7 $Y2=1.105
cc_19 VNB N_Y_c_364_n 0.00579788f $X=-0.19 $Y=-0.24 $X2=4.75 $Y2=1.105
cc_20 VNB N_Y_c_365_n 7.27967e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_366_n 0.0143227f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_22 VNB Y 0.0241054f $X=-0.19 $Y=-0.24 $X2=5.025 $Y2=1.11
cc_23 VNB N_Y_c_368_n 0.0122224f $X=-0.19 $Y=-0.24 $X2=0.745 $Y2=1.162
cc_24 VNB N_VGND_c_541_n 0.0141301f $X=-0.19 $Y=-0.24 $X2=1.995 $Y2=0.445
cc_25 VNB N_VGND_c_542_n 0.00218451f $X=-0.19 $Y=-0.24 $X2=2.38 $Y2=1.985
cc_26 VNB N_VGND_c_543_n 0.00217674f $X=-0.19 $Y=-0.24 $X2=2.475 $Y2=0.445
cc_27 VNB N_VGND_c_544_n 4.44285e-19 $X=-0.19 $Y=-0.24 $X2=2.85 $Y2=1.985
cc_28 VNB N_VGND_c_545_n 0.0150351f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_546_n 0.0155007f $X=-0.19 $Y=-0.24 $X2=3.32 $Y2=1.985
cc_30 VNB N_VGND_c_547_n 0.00510476f $X=-0.19 $Y=-0.24 $X2=3.435 $Y2=0.81
cc_31 VNB N_VGND_c_548_n 0.0155007f $X=-0.19 $Y=-0.24 $X2=3.435 $Y2=0.445
cc_32 VNB N_VGND_c_549_n 0.00577004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_550_n 0.0130599f $X=-0.19 $Y=-0.24 $X2=3.79 $Y2=1.985
cc_34 VNB N_VGND_c_551_n 0.00581396f $X=-0.19 $Y=-0.24 $X2=3.79 $Y2=1.985
cc_35 VNB N_VGND_c_552_n 0.0342426f $X=-0.19 $Y=-0.24 $X2=3.965 $Y2=0.445
cc_36 VNB N_VGND_c_553_n 0.0144539f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_554_n 0.0286462f $X=-0.19 $Y=-0.24 $X2=5.82 $Y2=1.985
cc_38 VNB N_VGND_c_555_n 0.337769f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_39 VNB N_VGND_c_556_n 0.00510476f $X=-0.19 $Y=-0.24 $X2=2.19 $Y2=1.105
cc_40 VNB N_VGND_c_557_n 0.00702712f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=1.105
cc_41 VPB N_A_c_101_n 0.0191485f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_42 VPB N_A_c_102_n 0.0160387f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_43 VPB N_A_c_103_n 0.0160577f $X=-0.19 $Y=1.305 $X2=1.44 $Y2=1.41
cc_44 VPB N_A_c_104_n 0.0160165f $X=-0.19 $Y=1.305 $X2=1.91 $Y2=1.41
cc_45 VPB N_A_c_105_n 0.0160165f $X=-0.19 $Y=1.305 $X2=2.38 $Y2=1.41
cc_46 VPB N_A_c_106_n 0.0160165f $X=-0.19 $Y=1.305 $X2=2.85 $Y2=1.41
cc_47 VPB N_A_c_107_n 0.0160165f $X=-0.19 $Y=1.305 $X2=3.32 $Y2=1.41
cc_48 VPB N_A_c_108_n 0.0164113f $X=-0.19 $Y=1.305 $X2=3.79 $Y2=1.41
cc_49 VPB N_A_c_109_n 0.0168061f $X=-0.19 $Y=1.305 $X2=4.31 $Y2=1.41
cc_50 VPB N_A_c_110_n 0.0168061f $X=-0.19 $Y=1.305 $X2=4.83 $Y2=1.41
cc_51 VPB N_A_c_111_n 0.0163925f $X=-0.19 $Y=1.305 $X2=5.35 $Y2=1.41
cc_52 VPB N_A_c_112_n 0.0191643f $X=-0.19 $Y=1.305 $X2=5.82 $Y2=1.41
cc_53 VPB N_A_c_100_n 0.151575f $X=-0.19 $Y=1.305 $X2=5.35 $Y2=1.16
cc_54 VPB N_VPWR_c_263_n 0.0114824f $X=-0.19 $Y=1.305 $X2=2.38 $Y2=1.985
cc_55 VPB N_VPWR_c_264_n 0.00523594f $X=-0.19 $Y=1.305 $X2=2.475 $Y2=0.81
cc_56 VPB N_VPWR_c_265_n 0.0194638f $X=-0.19 $Y=1.305 $X2=2.475 $Y2=0.445
cc_57 VPB N_VPWR_c_266_n 0.00522194f $X=-0.19 $Y=1.305 $X2=2.85 $Y2=1.985
cc_58 VPB N_VPWR_c_267_n 0.0194638f $X=-0.19 $Y=1.305 $X2=2.955 $Y2=0.445
cc_59 VPB N_VPWR_c_268_n 0.00522176f $X=-0.19 $Y=1.305 $X2=3.32 $Y2=1.985
cc_60 VPB N_VPWR_c_269_n 0.0196933f $X=-0.19 $Y=1.305 $X2=3.435 $Y2=0.81
cc_61 VPB N_VPWR_c_270_n 0.00513784f $X=-0.19 $Y=1.305 $X2=3.79 $Y2=1.41
cc_62 VPB N_VPWR_c_271_n 0.0195785f $X=-0.19 $Y=1.305 $X2=3.79 $Y2=1.985
cc_63 VPB N_VPWR_c_272_n 0.00547479f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_273_n 0.00544692f $X=-0.19 $Y=1.305 $X2=4.495 $Y2=0.81
cc_65 VPB N_VPWR_c_274_n 0.0153735f $X=-0.19 $Y=1.305 $X2=4.495 $Y2=0.445
cc_66 VPB N_VPWR_c_275_n 0.00520797f $X=-0.19 $Y=1.305 $X2=4.83 $Y2=1.41
cc_67 VPB N_VPWR_c_276_n 0.0209555f $X=-0.19 $Y=1.305 $X2=5.025 $Y2=0.81
cc_68 VPB N_VPWR_c_277_n 0.00574453f $X=-0.19 $Y=1.305 $X2=5.025 $Y2=0.445
cc_69 VPB N_VPWR_c_278_n 0.0194638f $X=-0.19 $Y=1.305 $X2=5.82 $Y2=1.985
cc_70 VPB N_VPWR_c_279_n 0.00497514f $X=-0.19 $Y=1.305 $X2=3.81 $Y2=1.105
cc_71 VPB N_VPWR_c_280_n 0.00497514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_281_n 0.00468662f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_282_n 0.00584071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_262_n 0.0518596f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.11
cc_75 VPB N_Y_c_356_n 0.00734091f $X=-0.19 $Y=1.305 $X2=2.955 $Y2=0.445
cc_76 VPB N_Y_c_370_n 0.00178529f $X=-0.19 $Y=1.305 $X2=3.32 $Y2=1.41
cc_77 VPB N_Y_c_371_n 0.00790647f $X=-0.19 $Y=1.305 $X2=3.32 $Y2=1.985
cc_78 VPB N_Y_c_372_n 0.00196324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_Y_c_373_n 0.00196324f $X=-0.19 $Y=1.305 $X2=4.31 $Y2=1.985
cc_80 VPB N_Y_c_374_n 0.00185282f $X=-0.19 $Y=1.305 $X2=5.35 $Y2=1.41
cc_81 VPB N_Y_c_375_n 0.00222477f $X=-0.19 $Y=1.305 $X2=3.81 $Y2=1.105
cc_82 VPB N_Y_c_376_n 0.00217247f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.11
cc_83 VPB N_Y_c_377_n 0.00223462f $X=-0.19 $Y=1.305 $X2=1.995 $Y2=1.11
cc_84 VPB N_Y_c_378_n 0.00142578f $X=-0.19 $Y=1.305 $X2=2.475 $Y2=1.11
cc_85 VPB N_Y_c_379_n 0.00142578f $X=-0.19 $Y=1.305 $X2=2.85 $Y2=1.11
cc_86 VPB N_Y_c_380_n 0.00148519f $X=-0.19 $Y=1.305 $X2=3.32 $Y2=1.11
cc_87 VPB N_Y_c_381_n 0.00145548f $X=-0.19 $Y=1.305 $X2=3.79 $Y2=1.11
cc_88 VPB N_Y_c_382_n 0.00181193f $X=-0.19 $Y=1.305 $X2=4.31 $Y2=1.11
cc_89 VPB N_Y_c_383_n 0.00173161f $X=-0.19 $Y=1.305 $X2=4.83 $Y2=1.11
cc_90 VPB Y 0.00849939f $X=-0.19 $Y=1.305 $X2=5.025 $Y2=1.11
cc_91 VPB N_Y_c_385_n 0.0140184f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.162
cc_92 N_A_c_101_n N_VPWR_c_264_n 0.00488841f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_93 N_A_c_101_n N_VPWR_c_265_n 0.00702461f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_c_102_n N_VPWR_c_265_n 0.00702461f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A_c_102_n N_VPWR_c_266_n 0.00302761f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A_c_103_n N_VPWR_c_266_n 0.00305721f $X=1.44 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A_c_103_n N_VPWR_c_267_n 0.00702461f $X=1.44 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A_c_104_n N_VPWR_c_267_n 0.00702461f $X=1.91 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A_c_104_n N_VPWR_c_268_n 0.0030489f $X=1.91 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A_c_105_n N_VPWR_c_268_n 0.0030489f $X=2.38 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_c_105_n N_VPWR_c_269_n 0.00702461f $X=2.38 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_c_106_n N_VPWR_c_269_n 0.00702461f $X=2.85 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_c_106_n N_VPWR_c_270_n 0.00297226f $X=2.85 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_c_107_n N_VPWR_c_270_n 0.00300127f $X=3.32 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A_c_107_n N_VPWR_c_271_n 0.00702461f $X=3.32 $Y=1.41 $X2=0 $Y2=0
cc_106 N_A_c_108_n N_VPWR_c_271_n 0.00702461f $X=3.79 $Y=1.41 $X2=0 $Y2=0
cc_107 N_A_c_108_n N_VPWR_c_272_n 0.00318005f $X=3.79 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A_c_109_n N_VPWR_c_272_n 0.00314909f $X=4.31 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A_c_110_n N_VPWR_c_273_n 0.00311335f $X=4.83 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A_c_111_n N_VPWR_c_273_n 0.00317485f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A_c_112_n N_VPWR_c_275_n 0.00483954f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A_c_109_n N_VPWR_c_276_n 0.00702461f $X=4.31 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_c_110_n N_VPWR_c_276_n 0.00702461f $X=4.83 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_c_111_n N_VPWR_c_278_n 0.00702461f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A_c_112_n N_VPWR_c_278_n 0.00702461f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A_c_101_n N_VPWR_c_262_n 0.0133734f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A_c_102_n N_VPWR_c_262_n 0.0124998f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A_c_103_n N_VPWR_c_262_n 0.0124873f $X=1.44 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_c_104_n N_VPWR_c_262_n 0.0124745f $X=1.91 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_c_105_n N_VPWR_c_262_n 0.0124745f $X=2.38 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_c_106_n N_VPWR_c_262_n 0.0124996f $X=2.85 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A_c_107_n N_VPWR_c_262_n 0.0124871f $X=3.32 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A_c_108_n N_VPWR_c_262_n 0.0125967f $X=3.79 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A_c_109_n N_VPWR_c_262_n 0.0127361f $X=4.31 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A_c_110_n N_VPWR_c_262_n 0.0127487f $X=4.83 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A_c_111_n N_VPWR_c_262_n 0.0125967f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A_c_112_n N_VPWR_c_262_n 0.0134831f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A_c_101_n N_Y_c_356_n 0.00180824f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_c_100_n N_Y_c_356_n 0.0199029f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A_c_152_p N_Y_c_356_n 0.0202172f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_M1000_g N_Y_c_357_n 0.00925734f $X=1.515 $Y=0.445 $X2=0 $Y2=0
cc_132 N_A_c_100_n N_Y_c_357_n 0.0433368f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_c_152_p N_Y_c_357_n 0.0860157f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A_c_101_n N_Y_c_370_n 0.0193394f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_c_100_n N_Y_c_370_n 0.00119794f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_c_152_p N_Y_c_370_n 0.0112679f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_c_102_n N_Y_c_372_n 0.0174373f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_c_103_n N_Y_c_372_n 0.0174373f $X=1.44 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_c_100_n N_Y_c_372_n 0.00963258f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A_c_152_p N_Y_c_372_n 0.050166f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A_M1000_g N_Y_c_359_n 0.00432033f $X=1.515 $Y=0.445 $X2=0 $Y2=0
cc_142 N_A_M1004_g N_Y_c_359_n 0.0010475f $X=1.995 $Y=0.445 $X2=0 $Y2=0
cc_143 N_A_c_104_n N_Y_c_373_n 0.0174075f $X=1.91 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_105_n N_Y_c_373_n 0.0174075f $X=2.38 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_c_100_n N_Y_c_373_n 0.00984483f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A_c_152_p N_Y_c_373_n 0.050166f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_M1004_g N_Y_c_360_n 0.00836783f $X=1.995 $Y=0.445 $X2=0 $Y2=0
cc_148 N_A_M1005_g N_Y_c_360_n 0.00807876f $X=2.475 $Y=0.445 $X2=0 $Y2=0
cc_149 N_A_c_100_n N_Y_c_360_n 0.0169026f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A_c_152_p N_Y_c_360_n 0.0538007f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_M1005_g N_Y_c_361_n 0.00432033f $X=2.475 $Y=0.445 $X2=0 $Y2=0
cc_152 N_A_M1007_g N_Y_c_361_n 0.0010475f $X=2.955 $Y=0.445 $X2=0 $Y2=0
cc_153 N_A_c_106_n N_Y_c_374_n 0.0174075f $X=2.85 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_c_107_n N_Y_c_374_n 0.0174075f $X=3.32 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_c_100_n N_Y_c_374_n 0.00944307f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_c_152_p N_Y_c_374_n 0.0490606f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A_M1007_g N_Y_c_362_n 0.00836783f $X=2.955 $Y=0.445 $X2=0 $Y2=0
cc_158 N_A_M1010_g N_Y_c_362_n 0.0076973f $X=3.435 $Y=0.445 $X2=0 $Y2=0
cc_159 N_A_c_100_n N_Y_c_362_n 0.0169026f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_c_152_p N_Y_c_362_n 0.0538007f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A_M1010_g N_Y_c_363_n 0.0041822f $X=3.435 $Y=0.445 $X2=0 $Y2=0
cc_162 N_A_M1012_g N_Y_c_363_n 0.00435198f $X=3.965 $Y=0.445 $X2=0 $Y2=0
cc_163 N_A_c_108_n N_Y_c_375_n 0.0176882f $X=3.79 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_c_109_n N_Y_c_375_n 0.0179689f $X=4.31 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A_c_100_n N_Y_c_375_n 0.0112243f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_c_152_p N_Y_c_375_n 0.0534822f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_M1012_g N_Y_c_364_n 0.0084179f $X=3.965 $Y=0.445 $X2=0 $Y2=0
cc_168 N_A_M1015_g N_Y_c_364_n 0.0084179f $X=4.495 $Y=0.445 $X2=0 $Y2=0
cc_169 N_A_c_100_n N_Y_c_364_n 0.0196083f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_c_152_p N_Y_c_364_n 0.0607966f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_M1015_g N_Y_c_365_n 0.00435198f $X=4.495 $Y=0.445 $X2=0 $Y2=0
cc_172 N_A_M1019_g N_Y_c_365_n 0.00435198f $X=5.025 $Y=0.445 $X2=0 $Y2=0
cc_173 N_A_c_110_n N_Y_c_376_n 0.0179689f $X=4.83 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_c_111_n N_Y_c_376_n 0.0176882f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_c_100_n N_Y_c_376_n 0.0109653f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A_c_152_p N_Y_c_376_n 0.0531137f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_M1019_g N_Y_c_366_n 0.00942691f $X=5.025 $Y=0.445 $X2=0 $Y2=0
cc_178 N_A_c_100_n N_Y_c_366_n 0.0389759f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_c_152_p N_Y_c_366_n 0.049637f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_c_112_n N_Y_c_377_n 0.0213094f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_c_100_n N_Y_c_377_n 0.00118224f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_c_100_n N_Y_c_378_n 0.00700529f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A_c_152_p N_Y_c_378_n 0.0198869f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A_c_100_n N_Y_c_379_n 0.007173f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_c_152_p N_Y_c_379_n 0.0198869f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_c_100_n N_Y_c_444_n 0.00697087f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_c_152_p N_Y_c_444_n 0.0147099f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A_c_100_n N_Y_c_380_n 0.00749172f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_c_152_p N_Y_c_380_n 0.0207155f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_c_100_n N_Y_c_448_n 0.00697087f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A_c_152_p N_Y_c_448_n 0.0147099f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_c_100_n N_Y_c_381_n 0.00737931f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_c_152_p N_Y_c_381_n 0.0203012f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_c_100_n N_Y_c_452_n 0.00797286f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A_c_152_p N_Y_c_452_n 0.0147099f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A_c_100_n N_Y_c_382_n 0.00922455f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A_c_152_p N_Y_c_382_n 0.0252729f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A_c_100_n N_Y_c_456_n 0.00797286f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A_c_152_p N_Y_c_456_n 0.0147099f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A_c_100_n N_Y_c_383_n 0.00800417f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A_c_152_p N_Y_c_383_n 0.0082862f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_202 N_A_c_112_n Y 0.00184784f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A_c_100_n Y 0.0209145f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A_c_152_p Y 0.0092936f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A_M1000_g N_VGND_c_541_n 0.00889184f $X=1.515 $Y=0.445 $X2=0 $Y2=0
cc_206 N_A_M1004_g N_VGND_c_541_n 5.82735e-19 $X=1.995 $Y=0.445 $X2=0 $Y2=0
cc_207 N_A_c_100_n N_VGND_c_541_n 0.00163455f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_208 N_A_M1004_g N_VGND_c_542_n 0.0016992f $X=1.995 $Y=0.445 $X2=0 $Y2=0
cc_209 N_A_M1005_g N_VGND_c_542_n 0.00778241f $X=2.475 $Y=0.445 $X2=0 $Y2=0
cc_210 N_A_M1007_g N_VGND_c_542_n 5.82735e-19 $X=2.955 $Y=0.445 $X2=0 $Y2=0
cc_211 N_A_c_100_n N_VGND_c_542_n 8.73002e-19 $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_M1007_g N_VGND_c_543_n 0.00171872f $X=2.955 $Y=0.445 $X2=0 $Y2=0
cc_213 N_A_M1010_g N_VGND_c_543_n 0.0104606f $X=3.435 $Y=0.445 $X2=0 $Y2=0
cc_214 N_A_M1012_g N_VGND_c_543_n 5.80786e-19 $X=3.965 $Y=0.445 $X2=0 $Y2=0
cc_215 N_A_c_100_n N_VGND_c_543_n 8.72612e-19 $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A_M1010_g N_VGND_c_544_n 5.32087e-19 $X=3.435 $Y=0.445 $X2=0 $Y2=0
cc_217 N_A_M1012_g N_VGND_c_544_n 0.00814801f $X=3.965 $Y=0.445 $X2=0 $Y2=0
cc_218 N_A_M1015_g N_VGND_c_544_n 0.00827666f $X=4.495 $Y=0.445 $X2=0 $Y2=0
cc_219 N_A_M1019_g N_VGND_c_544_n 5.48915e-19 $X=5.025 $Y=0.445 $X2=0 $Y2=0
cc_220 N_A_c_100_n N_VGND_c_544_n 0.00116239f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A_M1015_g N_VGND_c_545_n 5.48915e-19 $X=4.495 $Y=0.445 $X2=0 $Y2=0
cc_222 N_A_M1019_g N_VGND_c_545_n 0.00909943f $X=5.025 $Y=0.445 $X2=0 $Y2=0
cc_223 N_A_c_100_n N_VGND_c_545_n 0.00221504f $X=5.35 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A_M1000_g N_VGND_c_546_n 0.00360664f $X=1.515 $Y=0.445 $X2=0 $Y2=0
cc_225 N_A_M1004_g N_VGND_c_546_n 0.00433717f $X=1.995 $Y=0.445 $X2=0 $Y2=0
cc_226 N_A_M1005_g N_VGND_c_548_n 0.00360664f $X=2.475 $Y=0.445 $X2=0 $Y2=0
cc_227 N_A_M1007_g N_VGND_c_548_n 0.00433717f $X=2.955 $Y=0.445 $X2=0 $Y2=0
cc_228 N_A_M1010_g N_VGND_c_550_n 0.00216092f $X=3.435 $Y=0.445 $X2=0 $Y2=0
cc_229 N_A_M1012_g N_VGND_c_550_n 0.00360664f $X=3.965 $Y=0.445 $X2=0 $Y2=0
cc_230 N_A_M1015_g N_VGND_c_553_n 0.00360664f $X=4.495 $Y=0.445 $X2=0 $Y2=0
cc_231 N_A_M1019_g N_VGND_c_553_n 0.00360664f $X=5.025 $Y=0.445 $X2=0 $Y2=0
cc_232 N_A_M1000_g N_VGND_c_555_n 0.00440982f $X=1.515 $Y=0.445 $X2=0 $Y2=0
cc_233 N_A_M1004_g N_VGND_c_555_n 0.00610209f $X=1.995 $Y=0.445 $X2=0 $Y2=0
cc_234 N_A_M1005_g N_VGND_c_555_n 0.00440982f $X=2.475 $Y=0.445 $X2=0 $Y2=0
cc_235 N_A_M1007_g N_VGND_c_555_n 0.00610209f $X=2.955 $Y=0.445 $X2=0 $Y2=0
cc_236 N_A_M1010_g N_VGND_c_555_n 0.00311213f $X=3.435 $Y=0.445 $X2=0 $Y2=0
cc_237 N_A_M1012_g N_VGND_c_555_n 0.00452732f $X=3.965 $Y=0.445 $X2=0 $Y2=0
cc_238 N_A_M1015_g N_VGND_c_555_n 0.00452732f $X=4.495 $Y=0.445 $X2=0 $Y2=0
cc_239 N_A_M1019_g N_VGND_c_555_n 0.00452732f $X=5.025 $Y=0.445 $X2=0 $Y2=0
cc_240 N_VPWR_c_262_n N_Y_M1001_s 0.00414718f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_241 N_VPWR_c_262_n N_Y_M1003_s 0.00414718f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_242 N_VPWR_c_262_n N_Y_M1008_s 0.00380058f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_243 N_VPWR_c_262_n N_Y_M1011_s 0.00397388f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_244 N_VPWR_c_262_n N_Y_M1014_s 0.00403157f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_245 N_VPWR_c_262_n N_Y_M1017_s 0.00414718f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_246 N_VPWR_M1001_d N_Y_c_370_n 6.59072e-19 $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_247 N_VPWR_c_264_n N_Y_c_370_n 0.00508911f $X=0.26 $Y=1.965 $X2=0 $Y2=0
cc_248 N_VPWR_M1001_d N_Y_c_371_n 0.00237119f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_249 N_VPWR_c_264_n N_Y_c_371_n 0.0134341f $X=0.26 $Y=1.965 $X2=0 $Y2=0
cc_250 N_VPWR_c_265_n N_Y_c_473_n 0.012244f $X=1.075 $Y=2.72 $X2=0 $Y2=0
cc_251 N_VPWR_c_262_n N_Y_c_473_n 0.00903178f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_252 N_VPWR_M1002_d N_Y_c_372_n 0.00192406f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_253 N_VPWR_c_266_n N_Y_c_372_n 0.0147259f $X=1.205 $Y=1.965 $X2=0 $Y2=0
cc_254 N_VPWR_c_267_n N_Y_c_477_n 0.012244f $X=2.015 $Y=2.72 $X2=0 $Y2=0
cc_255 N_VPWR_c_262_n N_Y_c_477_n 0.00903178f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_256 N_VPWR_M1006_d N_Y_c_373_n 0.00187091f $X=2 $Y=1.485 $X2=0 $Y2=0
cc_257 N_VPWR_c_268_n N_Y_c_373_n 0.0143191f $X=2.145 $Y=1.965 $X2=0 $Y2=0
cc_258 N_VPWR_c_269_n N_Y_c_481_n 0.0125459f $X=2.965 $Y=2.72 $X2=0 $Y2=0
cc_259 N_VPWR_c_262_n N_Y_c_481_n 0.00941127f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_260 N_VPWR_M1009_d N_Y_c_374_n 0.00187091f $X=2.94 $Y=1.485 $X2=0 $Y2=0
cc_261 N_VPWR_c_270_n N_Y_c_374_n 0.0143191f $X=3.085 $Y=1.965 $X2=0 $Y2=0
cc_262 N_VPWR_c_271_n N_Y_c_485_n 0.0123949f $X=3.895 $Y=2.72 $X2=0 $Y2=0
cc_263 N_VPWR_c_262_n N_Y_c_485_n 0.00922153f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_264 N_VPWR_M1013_d N_Y_c_375_n 0.00240242f $X=3.88 $Y=1.485 $X2=0 $Y2=0
cc_265 N_VPWR_c_272_n N_Y_c_375_n 0.018387f $X=4.025 $Y=1.965 $X2=0 $Y2=0
cc_266 N_VPWR_c_276_n N_Y_c_489_n 0.0156435f $X=4.945 $Y=2.72 $X2=0 $Y2=0
cc_267 N_VPWR_c_262_n N_Y_c_489_n 0.0114984f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_268 N_VPWR_M1016_d N_Y_c_376_n 0.00240242f $X=4.92 $Y=1.485 $X2=0 $Y2=0
cc_269 N_VPWR_c_273_n N_Y_c_376_n 0.018387f $X=5.065 $Y=1.965 $X2=0 $Y2=0
cc_270 N_VPWR_c_278_n N_Y_c_493_n 0.012244f $X=5.925 $Y=2.72 $X2=0 $Y2=0
cc_271 N_VPWR_c_262_n N_Y_c_493_n 0.00903178f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_272 N_VPWR_M1018_d N_Y_c_377_n 9.77978e-19 $X=5.91 $Y=1.485 $X2=0 $Y2=0
cc_273 N_VPWR_c_275_n N_Y_c_377_n 0.00752987f $X=6.055 $Y=1.965 $X2=0 $Y2=0
cc_274 N_VPWR_M1018_d N_Y_c_385_n 0.0020392f $X=5.91 $Y=1.485 $X2=0 $Y2=0
cc_275 N_VPWR_c_275_n N_Y_c_385_n 0.0107293f $X=6.055 $Y=1.965 $X2=0 $Y2=0
cc_276 N_Y_c_357_n N_VGND_c_541_n 0.0232314f $X=1.685 $Y=0.78 $X2=0 $Y2=0
cc_277 N_Y_c_359_n N_VGND_c_541_n 0.0149566f $X=1.78 $Y=0.445 $X2=0 $Y2=0
cc_278 N_Y_c_360_n N_VGND_c_542_n 0.021795f $X=2.645 $Y=0.78 $X2=0 $Y2=0
cc_279 N_Y_c_361_n N_VGND_c_542_n 0.0149566f $X=2.74 $Y=0.445 $X2=0 $Y2=0
cc_280 N_Y_c_362_n N_VGND_c_543_n 0.0254298f $X=3.605 $Y=0.78 $X2=0 $Y2=0
cc_281 N_Y_c_363_n N_VGND_c_543_n 0.0184403f $X=3.7 $Y=0.445 $X2=0 $Y2=0
cc_282 N_Y_c_363_n N_VGND_c_544_n 0.0152658f $X=3.7 $Y=0.445 $X2=0 $Y2=0
cc_283 N_Y_c_364_n N_VGND_c_544_n 0.0283446f $X=4.665 $Y=0.78 $X2=0 $Y2=0
cc_284 N_Y_c_365_n N_VGND_c_544_n 0.0152658f $X=4.76 $Y=0.445 $X2=0 $Y2=0
cc_285 N_Y_c_365_n N_VGND_c_545_n 0.0152658f $X=4.76 $Y=0.445 $X2=0 $Y2=0
cc_286 N_Y_c_366_n N_VGND_c_545_n 0.0311189f $X=6.06 $Y=0.78 $X2=0 $Y2=0
cc_287 N_Y_c_357_n N_VGND_c_546_n 0.00330521f $X=1.685 $Y=0.78 $X2=0 $Y2=0
cc_288 N_Y_c_359_n N_VGND_c_546_n 0.0109465f $X=1.78 $Y=0.445 $X2=0 $Y2=0
cc_289 N_Y_c_360_n N_VGND_c_546_n 0.00325846f $X=2.645 $Y=0.78 $X2=0 $Y2=0
cc_290 N_Y_c_360_n N_VGND_c_548_n 0.00330521f $X=2.645 $Y=0.78 $X2=0 $Y2=0
cc_291 N_Y_c_361_n N_VGND_c_548_n 0.0109465f $X=2.74 $Y=0.445 $X2=0 $Y2=0
cc_292 N_Y_c_362_n N_VGND_c_548_n 0.00325846f $X=3.605 $Y=0.78 $X2=0 $Y2=0
cc_293 N_Y_c_362_n N_VGND_c_550_n 0.00259073f $X=3.605 $Y=0.78 $X2=0 $Y2=0
cc_294 N_Y_c_363_n N_VGND_c_550_n 0.0112652f $X=3.7 $Y=0.445 $X2=0 $Y2=0
cc_295 N_Y_c_364_n N_VGND_c_550_n 0.00330521f $X=4.665 $Y=0.78 $X2=0 $Y2=0
cc_296 N_Y_c_357_n N_VGND_c_552_n 0.0137196f $X=1.685 $Y=0.78 $X2=0 $Y2=0
cc_297 N_Y_c_358_n N_VGND_c_552_n 0.0030627f $X=0.285 $Y=0.78 $X2=0 $Y2=0
cc_298 N_Y_c_364_n N_VGND_c_553_n 0.00330521f $X=4.665 $Y=0.78 $X2=0 $Y2=0
cc_299 N_Y_c_365_n N_VGND_c_553_n 0.0112652f $X=4.76 $Y=0.445 $X2=0 $Y2=0
cc_300 N_Y_c_366_n N_VGND_c_553_n 0.00330521f $X=6.06 $Y=0.78 $X2=0 $Y2=0
cc_301 N_Y_c_366_n N_VGND_c_554_n 0.00895251f $X=6.06 $Y=0.78 $X2=0 $Y2=0
cc_302 N_Y_c_368_n N_VGND_c_554_n 0.0048643f $X=6.195 $Y=0.865 $X2=0 $Y2=0
cc_303 N_Y_M1000_s N_VGND_c_555_n 0.00327545f $X=1.59 $Y=0.235 $X2=0 $Y2=0
cc_304 N_Y_M1005_s N_VGND_c_555_n 0.00327545f $X=2.55 $Y=0.235 $X2=0 $Y2=0
cc_305 N_Y_M1010_s N_VGND_c_555_n 0.00393282f $X=3.51 $Y=0.235 $X2=0 $Y2=0
cc_306 N_Y_M1015_s N_VGND_c_555_n 0.00390323f $X=4.57 $Y=0.235 $X2=0 $Y2=0
cc_307 N_Y_c_357_n N_VGND_c_555_n 0.0296764f $X=1.685 $Y=0.78 $X2=0 $Y2=0
cc_308 N_Y_c_358_n N_VGND_c_555_n 0.00489372f $X=0.285 $Y=0.78 $X2=0 $Y2=0
cc_309 N_Y_c_359_n N_VGND_c_555_n 0.00712214f $X=1.78 $Y=0.445 $X2=0 $Y2=0
cc_310 N_Y_c_360_n N_VGND_c_555_n 0.0118085f $X=2.645 $Y=0.78 $X2=0 $Y2=0
cc_311 N_Y_c_361_n N_VGND_c_555_n 0.00712214f $X=2.74 $Y=0.445 $X2=0 $Y2=0
cc_312 N_Y_c_362_n N_VGND_c_555_n 0.010888f $X=3.605 $Y=0.78 $X2=0 $Y2=0
cc_313 N_Y_c_363_n N_VGND_c_555_n 0.00712214f $X=3.7 $Y=0.445 $X2=0 $Y2=0
cc_314 N_Y_c_364_n N_VGND_c_555_n 0.0123994f $X=4.665 $Y=0.78 $X2=0 $Y2=0
cc_315 N_Y_c_365_n N_VGND_c_555_n 0.00712214f $X=4.76 $Y=0.445 $X2=0 $Y2=0
cc_316 N_Y_c_366_n N_VGND_c_555_n 0.0220982f $X=6.06 $Y=0.78 $X2=0 $Y2=0
cc_317 N_Y_c_368_n N_VGND_c_555_n 0.00777238f $X=6.195 $Y=0.865 $X2=0 $Y2=0
