* File: sky130_fd_sc_hdll__and4_1.pex.spice
* Created: Thu Aug 27 18:58:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND4_1%A 2 3 5 8 10 17
r34 16 17 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r35 13 16 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=0.24 $Y=1.16
+ $X2=0.495 $Y2=1.16
r36 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r37 6 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.16
r38 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r39 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r40 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.89 $X2=0.495
+ $Y2=1.99
r41 1 16 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r42 1 2 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_1%B 3 6 7 9 10 11 15
r38 15 18 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.16 $X2=1
+ $Y2=1.325
r39 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.16 $X2=1
+ $Y2=0.995
r40 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.16
+ $X2=1 $Y2=1.16
r41 11 16 9.40151 $w=3.78e-07 $l=3.1e-07 $layer=LI1_cond $X=1.045 $Y=0.85
+ $X2=1.045 $Y2=1.16
r42 10 11 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=1.045 $Y=0.51
+ $X2=1.045 $Y2=0.85
r43 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.965 $Y=1.99
+ $X2=0.965 $Y2=2.275
r44 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.89 $X2=0.965
+ $Y2=1.99
r45 6 18 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.965 $Y=1.89
+ $X2=0.965 $Y2=1.325
r46 3 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.94 $Y=0.445
+ $X2=0.94 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_1%C 3 6 7 9 10 11 12 17
c39 17 0 1.0356e-19 $X=1.49 $Y=1.16
c40 10 0 2.74744e-20 $X=1.44 $Y=0.51
r41 17 20 40.3353 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.485 $Y=1.16
+ $X2=1.485 $Y2=1.325
r42 17 19 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.485 $Y=1.16
+ $X2=1.485 $Y2=0.995
r43 12 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.49
+ $Y=1.16 $X2=1.49 $Y2=1.16
r44 11 12 12.3192 $w=2.88e-07 $l=3.1e-07 $layer=LI1_cond $X=1.55 $Y=0.85
+ $X2=1.55 $Y2=1.16
r45 10 11 13.5114 $w=2.88e-07 $l=3.4e-07 $layer=LI1_cond $X=1.55 $Y=0.51
+ $X2=1.55 $Y2=0.85
r46 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.445 $Y=1.99
+ $X2=1.445 $Y2=2.275
r47 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.445 $Y=1.89 $X2=1.445
+ $Y2=1.99
r48 6 20 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=1.445 $Y=1.89
+ $X2=1.445 $Y2=1.325
r49 3 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.42 $Y=0.445
+ $X2=1.42 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_1%D 3 6 7 9 10 13 18
c43 13 0 1.65736e-19 $X=1.97 $Y=1.16
r44 13 16 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.97 $Y=1.16
+ $X2=1.97 $Y2=1.325
r45 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.97 $Y=1.16
+ $X2=1.97 $Y2=0.995
r46 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.97
+ $Y=1.16 $X2=1.97 $Y2=1.16
r47 10 18 2.98039 $w=6.08e-07 $l=1.52e-07 $layer=LI1_cond $X=2.062 $Y=1.02
+ $X2=1.91 $Y2=1.02
r48 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.935 $Y=1.99
+ $X2=1.935 $Y2=2.275
r49 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.935 $Y=1.89 $X2=1.935
+ $Y2=1.99
r50 6 16 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=1.935 $Y=1.89
+ $X2=1.935 $Y2=1.325
r51 3 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.91 $Y=0.445
+ $X2=1.91 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_1%A_27_47# 1 2 3 10 12 13 15 17 20 22 26 28
+ 32 38 40 41
c84 32 0 1.45514e-19 $X=2.45 $Y=1.16
c85 22 0 1.0356e-19 $X=1.56 $Y=1.58
r86 36 38 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=0.26 $Y=0.42
+ $X2=0.59 $Y2=0.42
r87 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.45
+ $Y=1.16 $X2=2.45 $Y2=1.16
r88 30 32 18.5773 $w=1.98e-07 $l=3.35e-07 $layer=LI1_cond $X=2.435 $Y=1.495
+ $X2=2.435 $Y2=1.16
r89 29 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.81 $Y=1.58
+ $X2=1.685 $Y2=1.58
r90 28 30 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.335 $Y=1.58
+ $X2=2.435 $Y2=1.495
r91 28 29 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.335 $Y=1.58
+ $X2=1.81 $Y2=1.58
r92 24 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.685 $Y=1.665
+ $X2=1.685 $Y2=1.58
r93 24 26 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.685 $Y=1.665
+ $X2=1.685 $Y2=2.3
r94 23 40 2.28545 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.855 $Y=1.58
+ $X2=0.675 $Y2=1.58
r95 22 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.56 $Y=1.58
+ $X2=1.685 $Y2=1.58
r96 22 23 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=1.56 $Y=1.58
+ $X2=0.855 $Y2=1.58
r97 18 40 4.14756 $w=2.2e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.675 $Y2=1.58
r98 18 20 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=2.3
r99 17 40 4.14756 $w=2.2e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.59 $Y=1.495
+ $X2=0.675 $Y2=1.58
r100 16 38 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.59 $Y=0.585
+ $X2=0.59 $Y2=0.42
r101 16 17 53.1196 $w=1.88e-07 $l=9.1e-07 $layer=LI1_cond $X=0.59 $Y=0.585
+ $X2=0.59 $Y2=1.495
r102 13 33 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.51 $Y=0.995
+ $X2=2.45 $Y2=1.16
r103 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.51 $Y=0.995
+ $X2=2.51 $Y2=0.56
r104 10 33 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.485 $Y=1.41
+ $X2=2.45 $Y2=1.16
r105 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.485 $Y=1.41
+ $X2=2.485 $Y2=1.985
r106 3 26 600 $w=1.7e-07 $l=3.00791e-07 $layer=licon1_PDIFF $count=1 $X=1.535
+ $Y=2.065 $X2=1.685 $Y2=2.3
r107 2 20 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.065 $X2=0.73 $Y2=2.3
r108 1 36 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_1%VPWR 1 2 3 10 12 16 18 22 24 26 33 34 40 43
c49 3 0 1.18039e-19 $X=2.025 $Y=2.065
r50 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r51 41 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r52 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r53 34 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r54 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r55 31 43 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.375 $Y=2.72
+ $X2=2.19 $Y2=2.72
r56 31 33 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.375 $Y=2.72
+ $X2=2.99 $Y2=2.72
r57 30 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r58 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r59 27 37 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r60 27 29 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 26 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=1.2 $Y2=2.72
r62 26 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=0.69 $Y2=2.72
r63 24 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r64 24 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r65 20 43 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2.72
r66 20 22 19.7784 $w=3.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2
r67 19 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.2 $Y2=2.72
r68 18 43 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=2.19 $Y2=2.72
r69 18 19 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=1.365 $Y2=2.72
r70 14 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.72
r71 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.34
r72 10 37 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.212 $Y2=2.72
r73 10 12 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.257 $Y2=2.34
r74 3 22 300 $w=1.7e-07 $l=2.55441e-07 $layer=licon1_PDIFF $count=2 $X=2.025
+ $Y=2.065 $X2=2.25 $Y2=2
r75 2 16 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=2.065 $X2=1.2 $Y2=2.34
r76 1 12 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_1%X 1 2 7 8 9 10 11 12 24 36 43
r19 43 44 1.43124 $w=3.88e-07 $l=5e-09 $layer=LI1_cond $X=2.89 $Y=2.21 $X2=2.89
+ $Y2=2.205
r20 24 41 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=2.955 $Y=0.85
+ $X2=2.955 $Y2=0.805
r21 12 47 2.65948 $w=3.88e-07 $l=9e-08 $layer=LI1_cond $X=2.89 $Y=2.25 $X2=2.89
+ $Y2=2.34
r22 12 43 1.18199 $w=3.88e-07 $l=4e-08 $layer=LI1_cond $X=2.89 $Y=2.25 $X2=2.89
+ $Y2=2.21
r23 12 44 1.77299 $w=2.58e-07 $l=4e-08 $layer=LI1_cond $X=2.955 $Y=2.165
+ $X2=2.955 $Y2=2.205
r24 11 12 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=2.955 $Y=1.87
+ $X2=2.955 $Y2=2.165
r25 11 31 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=2.955 $Y=1.87
+ $X2=2.955 $Y2=1.66
r26 10 31 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=2.955 $Y=1.53
+ $X2=2.955 $Y2=1.66
r27 9 10 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=2.955 $Y=1.19
+ $X2=2.955 $Y2=1.53
r28 8 41 1.87449 $w=3.88e-07 $l=2e-08 $layer=LI1_cond $X=2.89 $Y=0.785 $X2=2.89
+ $Y2=0.805
r29 8 9 14.1839 $w=2.58e-07 $l=3.2e-07 $layer=LI1_cond $X=2.955 $Y=0.87
+ $X2=2.955 $Y2=1.19
r30 8 24 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=2.955 $Y=0.87
+ $X2=2.955 $Y2=0.85
r31 7 8 8.1262 $w=3.88e-07 $l=2.75e-07 $layer=LI1_cond $X=2.89 $Y=0.51 $X2=2.89
+ $Y2=0.785
r32 7 36 3.84148 $w=3.88e-07 $l=1.3e-07 $layer=LI1_cond $X=2.89 $Y=0.51 $X2=2.89
+ $Y2=0.38
r33 2 47 600 $w=1.7e-07 $l=1.00869e-06 $layer=licon1_PDIFF $count=1 $X=2.575
+ $Y=1.485 $X2=2.91 $Y2=2.34
r34 2 31 300 $w=1.7e-07 $l=4.1334e-07 $layer=licon1_PDIFF $count=2 $X=2.575
+ $Y=1.485 $X2=2.91 $Y2=1.66
r35 1 36 91 $w=1.7e-07 $l=3.90832e-07 $layer=licon1_NDIFF $count=2 $X=2.585
+ $Y=0.235 $X2=2.91 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_1%VGND 1 6 8 10 17 18 21
c38 6 0 1.65736e-19 $X=2.175 $Y=0.38
r39 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r40 18 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r41 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r42 15 21 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.2
+ $Y2=0
r43 15 17 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.99
+ $Y2=0
r44 10 21 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.065 $Y=0 $X2=2.2
+ $Y2=0
r45 10 12 119.717 $w=1.68e-07 $l=1.835e-06 $layer=LI1_cond $X=2.065 $Y=0
+ $X2=0.23 $Y2=0
r46 8 22 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r47 8 12 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r48 4 21 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=0.085 $X2=2.2
+ $Y2=0
r49 4 6 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.2 $Y=0.085 $X2=2.2
+ $Y2=0.38
r50 1 6 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=1.985
+ $Y=0.235 $X2=2.175 $Y2=0.38
.ends

