* File: sky130_fd_sc_hdll__or2_1.pxi.spice
* Created: Wed Sep  2 08:47:28 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR2_1%B N_B_M1002_g N_B_c_40_n N_B_M1001_g B B
+ N_B_c_39_n PM_SKY130_FD_SC_HDLL__OR2_1%B
x_PM_SKY130_FD_SC_HDLL__OR2_1%A N_A_M1004_g N_A_c_64_n N_A_M1000_g A A
+ PM_SKY130_FD_SC_HDLL__OR2_1%A
x_PM_SKY130_FD_SC_HDLL__OR2_1%A_38_297# N_A_38_297#_M1002_d N_A_38_297#_M1001_s
+ N_A_38_297#_c_96_n N_A_38_297#_M1003_g N_A_38_297#_c_97_n N_A_38_297#_M1005_g
+ N_A_38_297#_c_98_n N_A_38_297#_c_117_n N_A_38_297#_c_102_n N_A_38_297#_c_99_n
+ N_A_38_297#_c_110_n PM_SKY130_FD_SC_HDLL__OR2_1%A_38_297#
x_PM_SKY130_FD_SC_HDLL__OR2_1%VPWR N_VPWR_M1000_d N_VPWR_c_150_n VPWR
+ N_VPWR_c_151_n N_VPWR_c_152_n N_VPWR_c_149_n N_VPWR_c_154_n
+ PM_SKY130_FD_SC_HDLL__OR2_1%VPWR
x_PM_SKY130_FD_SC_HDLL__OR2_1%X N_X_M1003_d N_X_M1005_d N_X_c_170_n X X
+ PM_SKY130_FD_SC_HDLL__OR2_1%X
x_PM_SKY130_FD_SC_HDLL__OR2_1%VGND N_VGND_M1002_s N_VGND_M1004_d N_VGND_c_196_n
+ N_VGND_c_197_n N_VGND_c_198_n N_VGND_c_199_n VGND N_VGND_c_200_n
+ N_VGND_c_201_n N_VGND_c_202_n PM_SKY130_FD_SC_HDLL__OR2_1%VGND
cc_1 VNB N_B_M1002_g 0.037386f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.445
cc_2 VNB B 0.0239552f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_B_c_39_n 0.0428512f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.202
cc_4 VNB N_A_M1004_g 0.0299841f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.445
cc_5 VNB N_A_c_64_n 0.0237369f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.41
cc_6 VNB A 0.00537191f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_7 VNB N_A_38_297#_c_96_n 0.0208212f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.695
cc_8 VNB N_A_38_297#_c_97_n 0.03444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_38_297#_c_98_n 0.00738117f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.16
cc_10 VNB N_A_38_297#_c_99_n 0.00186823f $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=1.16
cc_11 VNB N_VPWR_c_149_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_X_c_170_n 0.0366543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB X 0.0273524f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.16
cc_14 VNB N_VGND_c_196_n 0.0102177f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.695
cc_15 VNB N_VGND_c_197_n 0.0185f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_16 VNB N_VGND_c_198_n 0.0225618f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_199_n 0.00493424f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.202
cc_18 VNB N_VGND_c_200_n 0.0258489f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_201_n 0.144632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_202_n 0.00410625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VPB N_B_c_40_n 0.0231143f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.41
cc_22 VPB B 0.00508419f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_23 VPB N_B_c_39_n 0.0190951f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.202
cc_24 VPB N_A_c_64_n 0.0283335f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.41
cc_25 VPB A 0.00222914f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_26 VPB N_A_38_297#_c_97_n 0.0367685f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_A_38_297#_c_98_n 0.00158333f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.16
cc_28 VPB N_A_38_297#_c_102_n 0.0175009f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.202
cc_29 VPB N_A_38_297#_c_99_n 0.00147642f $X=-0.19 $Y=1.305 $X2=0.262 $Y2=1.16
cc_30 VPB N_VPWR_c_150_n 0.0216266f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.695
cc_31 VPB N_VPWR_c_151_n 0.0369884f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_152_n 0.0235972f $X=-0.19 $Y=1.305 $X2=0.262 $Y2=0.85
cc_33 VPB N_VPWR_c_149_n 0.0783203f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_154_n 0.00513801f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB X 0.0266613f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.16
cc_36 VPB X 0.0331333f $X=-0.19 $Y=1.305 $X2=0.262 $Y2=1.16
cc_37 N_B_M1002_g N_A_M1004_g 0.0170057f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_38 N_B_c_40_n N_A_c_64_n 0.0356345f $X=0.55 $Y=1.41 $X2=0 $Y2=0
cc_39 N_B_c_39_n N_A_c_64_n 0.0254794f $X=0.475 $Y=1.202 $X2=0 $Y2=0
cc_40 N_B_c_39_n A 2.77328e-19 $X=0.475 $Y=1.202 $X2=0 $Y2=0
cc_41 N_B_c_40_n N_A_38_297#_c_98_n 0.00390549f $X=0.55 $Y=1.41 $X2=0 $Y2=0
cc_42 B N_A_38_297#_c_98_n 0.0410481f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_43 N_B_c_39_n N_A_38_297#_c_98_n 0.0126153f $X=0.475 $Y=1.202 $X2=0 $Y2=0
cc_44 N_B_c_40_n N_A_38_297#_c_102_n 0.0222674f $X=0.55 $Y=1.41 $X2=0 $Y2=0
cc_45 B N_A_38_297#_c_102_n 0.0247514f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_46 N_B_c_39_n N_A_38_297#_c_102_n 0.00227952f $X=0.475 $Y=1.202 $X2=0 $Y2=0
cc_47 N_B_M1002_g N_A_38_297#_c_110_n 0.00705638f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_48 N_B_c_40_n N_VPWR_c_151_n 0.00393512f $X=0.55 $Y=1.41 $X2=0 $Y2=0
cc_49 N_B_c_40_n N_VPWR_c_149_n 0.00500987f $X=0.55 $Y=1.41 $X2=0 $Y2=0
cc_50 B N_VGND_c_196_n 3.74763e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_51 N_B_M1002_g N_VGND_c_197_n 0.00448362f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_52 B N_VGND_c_197_n 0.0206591f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_53 N_B_c_39_n N_VGND_c_197_n 0.00110332f $X=0.475 $Y=1.202 $X2=0 $Y2=0
cc_54 N_B_M1002_g N_VGND_c_198_n 0.00585385f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_55 N_B_M1002_g N_VGND_c_201_n 0.0104494f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_56 B N_VGND_c_201_n 0.0049547f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_57 N_A_M1004_g N_A_38_297#_c_96_n 0.0188645f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_58 A N_A_38_297#_c_96_n 0.00544127f $X=0.965 $Y=0.765 $X2=0 $Y2=0
cc_59 N_A_c_64_n N_A_38_297#_c_97_n 0.0389854f $X=0.96 $Y=1.41 $X2=0 $Y2=0
cc_60 N_A_M1004_g N_A_38_297#_c_98_n 0.00943794f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_61 N_A_c_64_n N_A_38_297#_c_98_n 0.00187654f $X=0.96 $Y=1.41 $X2=0 $Y2=0
cc_62 A N_A_38_297#_c_98_n 0.0420938f $X=0.965 $Y=0.765 $X2=0 $Y2=0
cc_63 N_A_c_64_n N_A_38_297#_c_117_n 0.0198704f $X=0.96 $Y=1.41 $X2=0 $Y2=0
cc_64 A N_A_38_297#_c_117_n 0.0239052f $X=0.965 $Y=0.765 $X2=0 $Y2=0
cc_65 N_A_c_64_n N_A_38_297#_c_102_n 8.66262e-19 $X=0.96 $Y=1.41 $X2=0 $Y2=0
cc_66 N_A_c_64_n N_A_38_297#_c_99_n 0.00111368f $X=0.96 $Y=1.41 $X2=0 $Y2=0
cc_67 A N_A_38_297#_c_99_n 0.0196459f $X=0.965 $Y=0.765 $X2=0 $Y2=0
cc_68 N_A_c_64_n N_VPWR_c_150_n 0.0040866f $X=0.96 $Y=1.41 $X2=0 $Y2=0
cc_69 N_A_c_64_n N_VPWR_c_151_n 0.00393512f $X=0.96 $Y=1.41 $X2=0 $Y2=0
cc_70 N_A_c_64_n N_VPWR_c_149_n 0.00500987f $X=0.96 $Y=1.41 $X2=0 $Y2=0
cc_71 N_A_M1004_g N_X_c_170_n 9.07816e-19 $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_72 A N_X_c_170_n 0.00386092f $X=0.965 $Y=0.765 $X2=0 $Y2=0
cc_73 A X 0.00549322f $X=0.965 $Y=0.765 $X2=0 $Y2=0
cc_74 A N_VGND_M1004_d 0.00329186f $X=0.965 $Y=0.765 $X2=0 $Y2=0
cc_75 N_A_M1004_g N_VGND_c_198_n 0.00585385f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_76 N_A_M1004_g N_VGND_c_199_n 0.00614826f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_77 N_A_c_64_n N_VGND_c_199_n 2.29546e-19 $X=0.96 $Y=1.41 $X2=0 $Y2=0
cc_78 A N_VGND_c_199_n 0.0131845f $X=0.965 $Y=0.765 $X2=0 $Y2=0
cc_79 N_A_M1004_g N_VGND_c_201_n 0.00933759f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_80 A N_VGND_c_201_n 0.00754496f $X=0.965 $Y=0.765 $X2=0 $Y2=0
cc_81 N_A_38_297#_c_117_n A_128_297# 0.00244196f $X=1.525 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_82 N_A_38_297#_c_102_n A_128_297# 0.00369906f $X=0.78 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_83 N_A_38_297#_c_117_n N_VPWR_M1000_d 0.00671898f $X=1.525 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_84 N_A_38_297#_c_97_n N_VPWR_c_150_n 0.0152645f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A_38_297#_c_117_n N_VPWR_c_150_n 0.0210126f $X=1.525 $Y=1.58 $X2=0 $Y2=0
cc_86 N_A_38_297#_c_97_n N_VPWR_c_152_n 0.00622633f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_38_297#_c_97_n N_VPWR_c_149_n 0.0116202f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A_38_297#_c_117_n N_X_M1005_d 0.00299646f $X=1.525 $Y=1.58 $X2=0 $Y2=0
cc_89 N_A_38_297#_c_96_n N_X_c_170_n 0.00886008f $X=1.47 $Y=0.995 $X2=0 $Y2=0
cc_90 N_A_38_297#_c_97_n N_X_c_170_n 0.00486646f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_91 N_A_38_297#_c_117_n N_X_c_170_n 2.26545e-19 $X=1.525 $Y=1.58 $X2=0 $Y2=0
cc_92 N_A_38_297#_c_99_n N_X_c_170_n 0.0161052f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_38_297#_c_96_n X 0.00241364f $X=1.47 $Y=0.995 $X2=0 $Y2=0
cc_94 N_A_38_297#_c_97_n X 0.0159899f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A_38_297#_c_117_n X 0.0143811f $X=1.525 $Y=1.58 $X2=0 $Y2=0
cc_96 N_A_38_297#_c_99_n X 0.0387356f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_38_297#_c_97_n X 0.0179667f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A_38_297#_c_117_n X 0.00843954f $X=1.525 $Y=1.58 $X2=0 $Y2=0
cc_99 N_A_38_297#_c_110_n N_VGND_c_198_n 0.0141521f $X=0.725 $Y=0.43 $X2=0 $Y2=0
cc_100 N_A_38_297#_c_96_n N_VGND_c_199_n 0.00291856f $X=1.47 $Y=0.995 $X2=0
+ $Y2=0
cc_101 N_A_38_297#_c_96_n N_VGND_c_200_n 0.00539883f $X=1.47 $Y=0.995 $X2=0
+ $Y2=0
cc_102 N_A_38_297#_M1002_d N_VGND_c_201_n 0.00490627f $X=0.55 $Y=0.235 $X2=0
+ $Y2=0
cc_103 N_A_38_297#_c_96_n N_VGND_c_201_n 0.0110745f $X=1.47 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A_38_297#_c_110_n N_VGND_c_201_n 0.00907366f $X=0.725 $Y=0.43 $X2=0
+ $Y2=0
cc_105 N_VPWR_c_149_n N_X_M1005_d 0.0049567f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_106 N_VPWR_c_150_n X 3.20848e-19 $X=1.26 $Y=1.92 $X2=0 $Y2=0
cc_107 N_VPWR_c_150_n X 0.0412204f $X=1.26 $Y=1.92 $X2=0 $Y2=0
cc_108 N_VPWR_c_152_n X 0.0401981f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_109 N_VPWR_c_149_n X 0.0218496f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_110 N_X_c_170_n N_VGND_c_200_n 0.0467348f $X=2.065 $Y=0.54 $X2=0 $Y2=0
cc_111 N_X_M1003_d N_VGND_c_201_n 0.00250339f $X=1.545 $Y=0.235 $X2=0 $Y2=0
cc_112 N_X_c_170_n N_VGND_c_201_n 0.0266101f $X=2.065 $Y=0.54 $X2=0 $Y2=0
