* File: sky130_fd_sc_hdll__nand2b_2.pex.spice
* Created: Thu Aug 27 19:13:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND2B_2%A_N 1 3 4 6 7 15
r25 11 15 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=0.54 $Y=1.16
+ $X2=0.695 $Y2=1.16
r26 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.54
+ $Y=1.16 $X2=0.54 $Y2=1.16
r27 7 15 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=0.745 $Y=1.16 $X2=0.695
+ $Y2=1.16
r28 4 10 47.6478 $w=3.03e-07 $l=2.80624e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.56 $Y2=1.16
r29 4 6 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.695
r30 1 10 38.5416 $w=3.03e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.56 $Y2=1.16
r31 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2B_2%A_27_93# 1 2 7 9 12 14 16 19 22 23 27 31
+ 38 42
c59 27 0 9.4217e-20 $X=1.105 $Y=1.16
c60 19 0 1.56657e-19 $X=1.83 $Y=0.56
r61 42 43 40.2934 $w=3.17e-07 $l=2.65e-07 $layer=POLY_cond $X=1.565 $Y=1.217
+ $X2=1.83 $Y2=1.217
r62 41 42 23.5678 $w=3.17e-07 $l=1.55e-07 $layer=POLY_cond $X=1.41 $Y=1.217
+ $X2=1.565 $Y2=1.217
r63 37 38 8.0507 $w=3.63e-07 $l=1.5e-07 $layer=LI1_cond $X=0.26 $Y=1.677
+ $X2=0.41 $Y2=1.677
r64 31 33 8.99284 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=0.227 $Y=0.675
+ $X2=0.227 $Y2=0.84
r65 28 41 46.3754 $w=3.17e-07 $l=3.05e-07 $layer=POLY_cond $X=1.105 $Y=1.217
+ $X2=1.41 $Y2=1.217
r66 28 39 10.6435 $w=3.17e-07 $l=7e-08 $layer=POLY_cond $X=1.105 $Y=1.217
+ $X2=1.035 $Y2=1.217
r67 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.105
+ $Y=1.16 $X2=1.105 $Y2=1.16
r68 25 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.105 $Y=1.495
+ $X2=1.105 $Y2=1.16
r69 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.02 $Y=1.58
+ $X2=1.105 $Y2=1.495
r70 23 38 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.02 $Y=1.58
+ $X2=0.41 $Y2=1.58
r71 22 37 2.0523 $w=3.63e-07 $l=6.5e-08 $layer=LI1_cond $X=0.195 $Y=1.677
+ $X2=0.26 $Y2=1.677
r72 22 33 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.195 $Y=1.495
+ $X2=0.195 $Y2=0.84
r73 17 43 20.269 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.83 $Y=1.025
+ $X2=1.83 $Y2=1.217
r74 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.83 $Y=1.025
+ $X2=1.83 $Y2=0.56
r75 14 42 15.9969 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.565 $Y=1.41
+ $X2=1.565 $Y2=1.217
r76 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.565 $Y=1.41
+ $X2=1.565 $Y2=1.985
r77 10 41 20.269 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=1.217
r78 10 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=0.56
r79 7 39 15.9969 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.035 $Y=1.41
+ $X2=1.035 $Y2=1.217
r80 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.035 $Y=1.41
+ $X2=1.035 $Y2=1.985
r81 2 37 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.695
r82 1 31 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2B_2%B 1 3 6 8 10 13 15 16 17 28 32
r52 28 29 3.57567 $w=3.37e-07 $l=2.5e-08 $layer=POLY_cond $X=2.695 $Y=1.217
+ $X2=2.72 $Y2=1.217
r53 26 28 10.727 $w=3.37e-07 $l=7.5e-08 $layer=POLY_cond $X=2.62 $Y=1.217
+ $X2=2.695 $Y2=1.217
r54 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.62
+ $Y=1.16 $X2=2.62 $Y2=1.16
r55 24 26 52.9199 $w=3.37e-07 $l=3.7e-07 $layer=POLY_cond $X=2.25 $Y=1.217
+ $X2=2.62 $Y2=1.217
r56 23 24 5.00593 $w=3.37e-07 $l=3.5e-08 $layer=POLY_cond $X=2.215 $Y=1.217
+ $X2=2.25 $Y2=1.217
r57 16 17 10.7196 $w=3.58e-07 $l=2.55e-07 $layer=LI1_cond $X=3 $Y=1.275 $X2=3
+ $Y2=1.53
r58 16 27 11.2937 $w=3.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.905 $Y=1.175
+ $X2=2.62 $Y2=1.175
r59 15 27 5.82273 $w=1.98e-07 $l=1.05e-07 $layer=LI1_cond $X=2.515 $Y=1.175
+ $X2=2.62 $Y2=1.175
r60 15 32 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=2.515 $Y=1.175
+ $X2=2.5 $Y2=1.175
r61 11 29 21.7231 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.72 $Y=1.025
+ $X2=2.72 $Y2=1.217
r62 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.72 $Y=1.025
+ $X2=2.72 $Y2=0.56
r63 8 28 17.4215 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.695 $Y=1.41
+ $X2=2.695 $Y2=1.217
r64 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.695 $Y=1.41
+ $X2=2.695 $Y2=1.985
r65 4 24 21.7231 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.25 $Y=1.025
+ $X2=2.25 $Y2=1.217
r66 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.25 $Y=1.025
+ $X2=2.25 $Y2=0.56
r67 1 23 17.4215 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.215 $Y=1.41
+ $X2=2.215 $Y2=1.217
r68 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.215 $Y=1.41
+ $X2=2.215 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2B_2%VPWR 1 2 3 14 18 20 22 25 26 27 33 38 42
r44 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r46 36 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r47 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r48 33 41 3.40825 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=2.845 $Y=2.72
+ $X2=3.032 $Y2=2.72
r49 33 35 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.845 $Y=2.72
+ $X2=2.53 $Y2=2.72
r50 32 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r51 32 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r53 29 38 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.885 $Y=2.72
+ $X2=0.757 $Y2=2.72
r54 29 31 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=0.885 $Y=2.72
+ $X2=1.61 $Y2=2.72
r55 27 39 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r56 25 31 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.725 $Y=2.72
+ $X2=1.61 $Y2=2.72
r57 25 26 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=1.725 $Y=2.72
+ $X2=1.912 $Y2=2.72
r58 24 35 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.1 $Y=2.72 $X2=2.53
+ $Y2=2.72
r59 24 26 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=2.1 $Y=2.72
+ $X2=1.912 $Y2=2.72
r60 20 41 3.40825 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=2.93 $Y=2.635
+ $X2=3.032 $Y2=2.72
r61 20 22 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.93 $Y=2.635
+ $X2=2.93 $Y2=2
r62 16 26 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.912 $Y=2.635
+ $X2=1.912 $Y2=2.72
r63 16 18 9.06588 $w=3.73e-07 $l=2.95e-07 $layer=LI1_cond $X=1.912 $Y=2.635
+ $X2=1.912 $Y2=2.34
r64 12 38 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.757 $Y=2.635
+ $X2=0.757 $Y2=2.72
r65 12 14 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=0.757 $Y=2.635
+ $X2=0.757 $Y2=2
r66 3 22 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.785
+ $Y=1.485 $X2=2.93 $Y2=2
r67 2 18 600 $w=1.7e-07 $l=9.7857e-07 $layer=licon1_PDIFF $count=1 $X=1.655
+ $Y=1.485 $X2=1.92 $Y2=2.34
r68 1 14 300 $w=1.7e-07 $l=6.13148e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.8 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2B_2%Y 1 2 3 10 11 16 19 20 21 22 23 31 43
c44 31 0 1.95148e-19 $X=1.62 $Y=0.72
c45 2 0 9.4217e-20 $X=1.125 $Y=1.485
r46 41 43 9.08189 $w=4.03e-07 $l=4.17133e-07 $layer=LI1_cond $X=1.3 $Y=2.15
+ $X2=1.6 $Y2=1.87
r47 23 31 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=1.62 $Y=0.85
+ $X2=1.62 $Y2=0.72
r48 22 29 0.30273 $w=4.03e-07 $l=6.48074e-08 $layer=LI1_cond $X=1.61 $Y=1.895
+ $X2=1.62 $Y2=1.835
r49 22 43 0.30273 $w=4.03e-07 $l=2.95804e-08 $layer=LI1_cond $X=1.61 $Y=1.895
+ $X2=1.6 $Y2=1.87
r50 22 29 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=1.62 $Y=1.81
+ $X2=1.62 $Y2=1.835
r51 21 22 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.62 $Y=1.53 $X2=1.62
+ $Y2=1.81
r52 20 21 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.62 $Y=1.19
+ $X2=1.62 $Y2=1.53
r53 20 23 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.62 $Y=1.19
+ $X2=1.62 $Y2=0.85
r54 14 19 3.12539 $w=3.02e-07 $l=9.75705e-08 $layer=LI1_cond $X=2.477 $Y=1.835
+ $X2=2.45 $Y2=1.92
r55 14 16 7.33373 $w=2.73e-07 $l=1.75e-07 $layer=LI1_cond $X=2.477 $Y=1.835
+ $X2=2.477 $Y2=1.66
r56 11 29 9.1679 $w=4.03e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.785 $Y=1.92
+ $X2=1.62 $Y2=1.835
r57 10 19 3.47949 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=1.92
+ $X2=2.45 $Y2=1.92
r58 10 11 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.285 $Y=1.92
+ $X2=1.785 $Y2=1.92
r59 3 19 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.305
+ $Y=1.485 $X2=2.45 $Y2=2
r60 3 16 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.305
+ $Y=1.485 $X2=2.45 $Y2=1.66
r61 2 41 300 $w=1.7e-07 $l=5.96112e-07 $layer=licon1_PDIFF $count=2 $X=1.125
+ $Y=1.485 $X2=1.3 $Y2=2
r62 1 31 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.62 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2B_2%VGND 1 2 9 13 16 17 18 20 30 31 34
r44 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r45 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r46 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r47 28 35 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=0.69
+ $Y2=0
r48 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r49 25 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.68
+ $Y2=0
r50 25 27 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=0.765 $Y=0 $X2=2.07
+ $Y2=0
r51 20 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.68
+ $Y2=0
r52 20 22 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r53 18 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r54 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r55 16 27 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.07
+ $Y2=0
r56 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.51
+ $Y2=0
r57 15 30 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.595 $Y=0 $X2=2.99
+ $Y2=0
r58 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=0 $X2=2.51
+ $Y2=0
r59 11 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=0.085
+ $X2=2.51 $Y2=0
r60 11 13 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.51 $Y=0.085
+ $X2=2.51 $Y2=0.36
r61 7 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0
r62 7 9 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.61
r63 2 13 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.235 $X2=2.51 $Y2=0.36
r64 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.465 $X2=0.68 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2B_2%A_215_47# 1 2 3 10 14 15 16 20
c39 15 0 1.56657e-19 $X=2.08 $Y=0.695
r40 18 20 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.93 $Y=0.695
+ $X2=2.93 $Y2=0.38
r41 17 25 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.205 $Y=0.8
+ $X2=2.08 $Y2=0.8
r42 16 18 7.26367 $w=2.1e-07 $l=2.11069e-07 $layer=LI1_cond $X=2.765 $Y=0.8
+ $X2=2.93 $Y2=0.695
r43 16 17 29.5758 $w=2.08e-07 $l=5.6e-07 $layer=LI1_cond $X=2.765 $Y=0.8
+ $X2=2.205 $Y2=0.8
r44 15 25 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=2.08 $Y=0.695
+ $X2=2.08 $Y2=0.8
r45 14 23 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=2.08 $Y=0.465
+ $X2=2.08 $Y2=0.36
r46 14 15 10.6025 $w=2.48e-07 $l=2.3e-07 $layer=LI1_cond $X=2.08 $Y=0.465
+ $X2=2.08 $Y2=0.695
r47 10 23 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.955 $Y=0.36
+ $X2=2.08 $Y2=0.36
r48 10 12 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=1.955 $Y=0.36
+ $X2=1.2 $Y2=0.36
r49 3 20 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.795
+ $Y=0.235 $X2=2.93 $Y2=0.38
r50 2 25 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.72
r51 2 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.38
r52 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.38
.ends

