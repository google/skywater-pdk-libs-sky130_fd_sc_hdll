* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__bufbuf_16 A VGND VNB VPB VPWR X
M1000 X a_589_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.32e+12p pd=2.064e+07u as=4.02e+12p ps=3.604e+07u
M1001 VGND a_589_47# X VNB nshort w=650000u l=150000u
+  ad=2.8015e+12p pd=2.682e+07u as=1.6965e+12p ps=1.562e+07u
M1002 X a_589_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_589_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_589_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_225_47# a_589_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.7e+11p ps=7.74e+06u
M1006 VGND a_589_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_589_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_225_47# a_589_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_589_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_589_47# a_225_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_589_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_589_47# a_225_47# VGND VNB nshort w=650000u l=150000u
+  ad=6.565e+11p pd=5.92e+06u as=0p ps=0u
M1013 X a_589_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_225_47# a_589_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_589_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_589_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_589_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_589_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_589_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_117_297# a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.095e+11p ps=3.86e+06u
M1021 X a_589_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_117_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1023 VGND a_225_47# a_589_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_589_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_589_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 X a_589_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR a_117_297# a_225_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.6e+11p ps=5.12e+06u
M1028 VGND a_589_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_589_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 X a_589_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_589_47# a_225_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 X a_589_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_589_47# a_225_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 X a_589_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_225_47# a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 X a_589_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_117_297# A VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1038 a_225_47# a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR a_225_47# a_589_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VPWR a_589_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPWR a_589_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPWR a_117_297# a_225_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VGND a_589_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VPWR a_589_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_589_47# a_225_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 VPWR a_589_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VGND a_225_47# a_589_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 X a_589_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_589_47# a_225_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1050 VGND a_117_297# a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1051 VGND a_589_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
