# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__muxb16to1_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  25.76000 BY  5.440000 ;
  SITE unithd ;
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.055000 0.915000 1.325000 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.525000 1.055000 6.345000 1.325000 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.535000 1.055000 7.355000 1.325000 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.965000 1.055000 12.785000 1.325000 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.975000 1.055000 13.795000 1.325000 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.405000 1.055000 19.225000 1.325000 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.415000 1.055000 20.235000 1.325000 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 24.845000 1.055000 25.665000 1.325000 ;
    END
  END D[7]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 4.115000 0.915000 4.385000 ;
    END
  END D[8]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.525000 4.115000 6.345000 4.385000 ;
    END
  END D[9]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.535000 4.115000 7.355000 4.385000 ;
    END
  END D[10]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.965000 4.115000 12.785000 4.385000 ;
    END
  END D[11]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.975000 4.115000 13.795000 4.385000 ;
    END
  END D[12]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.405000 4.115000 19.225000 4.385000 ;
    END
  END D[13]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.415000 4.115000 20.235000 4.385000 ;
    END
  END D[14]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 24.845000 4.115000 25.665000 4.385000 ;
    END
  END D[15]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 1.025000 3.125000 1.295000 ;
    END
  END S[0]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 1.025000 3.650000 1.295000 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.230000 1.025000 9.565000 1.295000 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.755000 1.025000 10.090000 1.295000 ;
    END
  END S[3]
  PIN S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.670000 1.025000 16.005000 1.295000 ;
    END
  END S[4]
  PIN S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.195000 1.025000 16.530000 1.295000 ;
    END
  END S[5]
  PIN S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 22.110000 1.025000 22.445000 1.295000 ;
    END
  END S[6]
  PIN S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 22.635000 1.025000 22.970000 1.295000 ;
    END
  END S[7]
  PIN S[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 4.145000 3.125000 4.415000 ;
    END
  END S[8]
  PIN S[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 4.145000 3.650000 4.415000 ;
    END
  END S[9]
  PIN S[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.230000 4.145000 9.565000 4.415000 ;
    END
  END S[10]
  PIN S[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.755000 4.145000 10.090000 4.415000 ;
    END
  END S[11]
  PIN S[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.670000 4.145000 16.005000 4.415000 ;
    END
  END S[12]
  PIN S[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.195000 4.145000 16.530000 4.415000 ;
    END
  END S[13]
  PIN S[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 22.110000 4.145000 22.445000 4.415000 ;
    END
  END S[14]
  PIN S[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 22.635000 4.145000 22.970000 4.415000 ;
    END
  END S[15]
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 25.760000 0.240000 ;
        RECT 0.000000  5.200000 25.760000 5.680000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 25.760000 2.960000 ;
    END
  END VPWR
  PIN Z
    ANTENNADIFFAREA  1.992000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  1.465000 1.755000  1.755000 1.800000 ;
        RECT  1.465000 1.800000 24.295000 1.940000 ;
        RECT  1.465000 1.940000  1.755000 1.985000 ;
        RECT  1.465000 3.455000  1.755000 3.500000 ;
        RECT  1.465000 3.500000 24.295000 3.640000 ;
        RECT  1.465000 3.640000  1.755000 3.685000 ;
        RECT  4.685000 1.755000  4.975000 1.800000 ;
        RECT  4.685000 1.940000  4.975000 1.985000 ;
        RECT  4.685000 3.455000  4.975000 3.500000 ;
        RECT  4.685000 3.640000  4.975000 3.685000 ;
        RECT  7.905000 1.755000  8.195000 1.800000 ;
        RECT  7.905000 1.940000  8.195000 1.985000 ;
        RECT  7.905000 3.455000  8.195000 3.500000 ;
        RECT  7.905000 3.640000  8.195000 3.685000 ;
        RECT 11.125000 1.755000 11.415000 1.800000 ;
        RECT 11.125000 1.940000 11.415000 1.985000 ;
        RECT 11.125000 3.455000 11.415000 3.500000 ;
        RECT 11.125000 3.640000 11.415000 3.685000 ;
        RECT 14.345000 1.755000 14.635000 1.800000 ;
        RECT 14.345000 1.940000 14.635000 1.985000 ;
        RECT 14.345000 3.455000 14.635000 3.500000 ;
        RECT 14.345000 3.640000 14.635000 3.685000 ;
        RECT 17.565000 1.755000 17.855000 1.800000 ;
        RECT 17.565000 1.940000 17.855000 1.985000 ;
        RECT 17.565000 3.455000 17.855000 3.500000 ;
        RECT 17.565000 3.640000 17.855000 3.685000 ;
        RECT 20.785000 1.755000 21.075000 1.800000 ;
        RECT 20.785000 1.940000 21.075000 1.985000 ;
        RECT 20.785000 3.455000 21.075000 3.500000 ;
        RECT 20.785000 3.640000 21.075000 3.685000 ;
        RECT 24.005000 1.755000 24.295000 1.800000 ;
        RECT 24.005000 1.940000 24.295000 1.985000 ;
        RECT 24.005000 3.455000 24.295000 3.500000 ;
        RECT 24.005000 3.640000 24.295000 3.685000 ;
    END
  END Z
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 25.760000 0.085000 ;
      RECT  0.000000  2.635000  1.415000 2.805000 ;
      RECT  0.000000  5.355000 25.760000 5.525000 ;
      RECT  0.095000  1.495000  1.285000 1.665000 ;
      RECT  0.095000  1.665000  0.395000 2.210000 ;
      RECT  0.095000  2.210000  0.425000 2.465000 ;
      RECT  0.095000  2.975000  0.425000 3.230000 ;
      RECT  0.095000  3.230000  0.395000 3.775000 ;
      RECT  0.095000  3.775000  1.285000 3.945000 ;
      RECT  0.145000  0.255000  0.475000 0.715000 ;
      RECT  0.145000  0.715000  1.335000 0.885000 ;
      RECT  0.145000  4.555000  1.335000 4.725000 ;
      RECT  0.145000  4.725000  0.475000 5.185000 ;
      RECT  0.565000  1.835000  0.895000 2.105000 ;
      RECT  0.565000  3.335000  0.895000 3.605000 ;
      RECT  0.595000  2.105000  0.895000 2.635000 ;
      RECT  0.595000  2.805000  0.895000 3.335000 ;
      RECT  0.645000  0.085000  0.860000 0.545000 ;
      RECT  0.645000  4.895000  0.860000 5.355000 ;
      RECT  1.030000  0.255000  2.175000 0.425000 ;
      RECT  1.030000  0.425000  1.335000 0.715000 ;
      RECT  1.030000  0.885000  1.335000 0.925000 ;
      RECT  1.030000  4.515000  1.335000 4.555000 ;
      RECT  1.030000  4.725000  1.335000 5.015000 ;
      RECT  1.030000  5.015000  2.175000 5.185000 ;
      RECT  1.115000  1.665000  1.285000 2.295000 ;
      RECT  1.115000  2.295000  1.415000 2.465000 ;
      RECT  1.115000  2.975000  1.415000 3.145000 ;
      RECT  1.115000  3.145000  1.285000 3.775000 ;
      RECT  1.465000  1.755000  1.895000 2.125000 ;
      RECT  1.465000  3.315000  1.895000 3.685000 ;
      RECT  1.505000  0.595000  1.835000 0.885000 ;
      RECT  1.505000  4.555000  1.835000 4.845000 ;
      RECT  1.585000  0.885000  1.755000 1.755000 ;
      RECT  1.585000  2.125000  1.755000 3.315000 ;
      RECT  1.585000  3.685000  1.755000 4.555000 ;
      RECT  1.925000  2.295000  2.280000 2.465000 ;
      RECT  1.925000  2.635000  4.515000 2.805000 ;
      RECT  1.925000  2.975000  2.280000 3.145000 ;
      RECT  2.005000  0.425000  2.175000 0.770000 ;
      RECT  2.005000  4.670000  2.175000 5.015000 ;
      RECT  2.100000  1.205000  2.515000 1.305000 ;
      RECT  2.100000  1.305000  2.620000 1.465000 ;
      RECT  2.100000  1.465000  2.880000 1.475000 ;
      RECT  2.100000  3.965000  2.880000 3.975000 ;
      RECT  2.100000  3.975000  2.620000 4.135000 ;
      RECT  2.100000  4.135000  2.515000 4.235000 ;
      RECT  2.110000  1.645000  2.280000 2.295000 ;
      RECT  2.110000  3.145000  2.280000 3.795000 ;
      RECT  2.345000  0.585000  2.925000 0.755000 ;
      RECT  2.345000  0.755000  2.515000 1.205000 ;
      RECT  2.345000  4.235000  2.515000 4.685000 ;
      RECT  2.345000  4.685000  2.925000 4.855000 ;
      RECT  2.450000  1.475000  2.880000 1.635000 ;
      RECT  2.450000  3.805000  2.880000 3.965000 ;
      RECT  2.550000  1.635000  2.880000 2.465000 ;
      RECT  2.550000  2.975000  2.880000 3.805000 ;
      RECT  2.675000  0.330000  2.925000 0.585000 ;
      RECT  2.675000  4.855000  2.925000 5.110000 ;
      RECT  3.055000  1.465000  3.385000 2.635000 ;
      RECT  3.055000  2.805000  3.385000 3.975000 ;
      RECT  3.095000  0.085000  3.345000 0.660000 ;
      RECT  3.095000  4.780000  3.345000 5.355000 ;
      RECT  3.515000  0.330000  3.765000 0.585000 ;
      RECT  3.515000  0.585000  4.095000 0.755000 ;
      RECT  3.515000  4.685000  4.095000 4.855000 ;
      RECT  3.515000  4.855000  3.765000 5.110000 ;
      RECT  3.560000  1.465000  4.340000 1.475000 ;
      RECT  3.560000  1.475000  3.990000 1.635000 ;
      RECT  3.560000  1.635000  3.890000 2.465000 ;
      RECT  3.560000  2.975000  3.890000 3.805000 ;
      RECT  3.560000  3.805000  3.990000 3.965000 ;
      RECT  3.560000  3.965000  4.340000 3.975000 ;
      RECT  3.820000  1.305000  4.340000 1.465000 ;
      RECT  3.820000  3.975000  4.340000 4.135000 ;
      RECT  3.925000  0.755000  4.095000 1.205000 ;
      RECT  3.925000  1.205000  4.340000 1.305000 ;
      RECT  3.925000  4.135000  4.340000 4.235000 ;
      RECT  3.925000  4.235000  4.095000 4.685000 ;
      RECT  4.160000  1.645000  4.330000 2.295000 ;
      RECT  4.160000  2.295000  4.515000 2.465000 ;
      RECT  4.160000  2.975000  4.515000 3.145000 ;
      RECT  4.160000  3.145000  4.330000 3.795000 ;
      RECT  4.265000  0.255000  5.410000 0.425000 ;
      RECT  4.265000  0.425000  4.435000 0.770000 ;
      RECT  4.265000  4.670000  4.435000 5.015000 ;
      RECT  4.265000  5.015000  5.410000 5.185000 ;
      RECT  4.545000  1.755000  4.975000 2.125000 ;
      RECT  4.545000  3.315000  4.975000 3.685000 ;
      RECT  4.605000  0.595000  4.935000 0.885000 ;
      RECT  4.605000  4.555000  4.935000 4.845000 ;
      RECT  4.685000  0.885000  4.855000 1.755000 ;
      RECT  4.685000  2.125000  4.855000 3.315000 ;
      RECT  4.685000  3.685000  4.855000 4.555000 ;
      RECT  5.025000  2.295000  5.325000 2.465000 ;
      RECT  5.025000  2.635000  7.855000 2.805000 ;
      RECT  5.025000  2.975000  5.325000 3.145000 ;
      RECT  5.105000  0.425000  5.410000 0.715000 ;
      RECT  5.105000  0.715000  6.295000 0.885000 ;
      RECT  5.105000  0.885000  5.410000 0.925000 ;
      RECT  5.105000  4.515000  5.410000 4.555000 ;
      RECT  5.105000  4.555000  6.295000 4.725000 ;
      RECT  5.105000  4.725000  5.410000 5.015000 ;
      RECT  5.155000  1.495000  6.345000 1.665000 ;
      RECT  5.155000  1.665000  5.325000 2.295000 ;
      RECT  5.155000  3.145000  5.325000 3.775000 ;
      RECT  5.155000  3.775000  6.345000 3.945000 ;
      RECT  5.545000  1.835000  5.875000 2.105000 ;
      RECT  5.545000  2.105000  5.845000 2.635000 ;
      RECT  5.545000  2.805000  5.845000 3.335000 ;
      RECT  5.545000  3.335000  5.875000 3.605000 ;
      RECT  5.580000  0.085000  5.795000 0.545000 ;
      RECT  5.580000  4.895000  5.795000 5.355000 ;
      RECT  5.965000  0.255000  6.295000 0.715000 ;
      RECT  5.965000  4.725000  6.295000 5.185000 ;
      RECT  6.015000  2.210000  6.345000 2.465000 ;
      RECT  6.015000  2.975000  6.345000 3.230000 ;
      RECT  6.045000  1.665000  6.345000 2.210000 ;
      RECT  6.045000  3.230000  6.345000 3.775000 ;
      RECT  6.535000  1.495000  7.725000 1.665000 ;
      RECT  6.535000  1.665000  6.835000 2.210000 ;
      RECT  6.535000  2.210000  6.865000 2.465000 ;
      RECT  6.535000  2.975000  6.865000 3.230000 ;
      RECT  6.535000  3.230000  6.835000 3.775000 ;
      RECT  6.535000  3.775000  7.725000 3.945000 ;
      RECT  6.585000  0.255000  6.915000 0.715000 ;
      RECT  6.585000  0.715000  7.775000 0.885000 ;
      RECT  6.585000  4.555000  7.775000 4.725000 ;
      RECT  6.585000  4.725000  6.915000 5.185000 ;
      RECT  7.005000  1.835000  7.335000 2.105000 ;
      RECT  7.005000  3.335000  7.335000 3.605000 ;
      RECT  7.035000  2.105000  7.335000 2.635000 ;
      RECT  7.035000  2.805000  7.335000 3.335000 ;
      RECT  7.085000  0.085000  7.300000 0.545000 ;
      RECT  7.085000  4.895000  7.300000 5.355000 ;
      RECT  7.470000  0.255000  8.615000 0.425000 ;
      RECT  7.470000  0.425000  7.775000 0.715000 ;
      RECT  7.470000  0.885000  7.775000 0.925000 ;
      RECT  7.470000  4.515000  7.775000 4.555000 ;
      RECT  7.470000  4.725000  7.775000 5.015000 ;
      RECT  7.470000  5.015000  8.615000 5.185000 ;
      RECT  7.555000  1.665000  7.725000 2.295000 ;
      RECT  7.555000  2.295000  7.855000 2.465000 ;
      RECT  7.555000  2.975000  7.855000 3.145000 ;
      RECT  7.555000  3.145000  7.725000 3.775000 ;
      RECT  7.905000  1.755000  8.335000 2.125000 ;
      RECT  7.905000  3.315000  8.335000 3.685000 ;
      RECT  7.945000  0.595000  8.275000 0.885000 ;
      RECT  7.945000  4.555000  8.275000 4.845000 ;
      RECT  8.025000  0.885000  8.195000 1.755000 ;
      RECT  8.025000  2.125000  8.195000 3.315000 ;
      RECT  8.025000  3.685000  8.195000 4.555000 ;
      RECT  8.365000  2.295000  8.720000 2.465000 ;
      RECT  8.365000  2.635000 10.955000 2.805000 ;
      RECT  8.365000  2.975000  8.720000 3.145000 ;
      RECT  8.445000  0.425000  8.615000 0.770000 ;
      RECT  8.445000  4.670000  8.615000 5.015000 ;
      RECT  8.540000  1.205000  8.955000 1.305000 ;
      RECT  8.540000  1.305000  9.060000 1.465000 ;
      RECT  8.540000  1.465000  9.320000 1.475000 ;
      RECT  8.540000  3.965000  9.320000 3.975000 ;
      RECT  8.540000  3.975000  9.060000 4.135000 ;
      RECT  8.540000  4.135000  8.955000 4.235000 ;
      RECT  8.550000  1.645000  8.720000 2.295000 ;
      RECT  8.550000  3.145000  8.720000 3.795000 ;
      RECT  8.785000  0.585000  9.365000 0.755000 ;
      RECT  8.785000  0.755000  8.955000 1.205000 ;
      RECT  8.785000  4.235000  8.955000 4.685000 ;
      RECT  8.785000  4.685000  9.365000 4.855000 ;
      RECT  8.890000  1.475000  9.320000 1.635000 ;
      RECT  8.890000  3.805000  9.320000 3.965000 ;
      RECT  8.990000  1.635000  9.320000 2.465000 ;
      RECT  8.990000  2.975000  9.320000 3.805000 ;
      RECT  9.115000  0.330000  9.365000 0.585000 ;
      RECT  9.115000  4.855000  9.365000 5.110000 ;
      RECT  9.495000  1.465000  9.825000 2.635000 ;
      RECT  9.495000  2.805000  9.825000 3.975000 ;
      RECT  9.535000  0.085000  9.785000 0.660000 ;
      RECT  9.535000  4.780000  9.785000 5.355000 ;
      RECT  9.955000  0.330000 10.205000 0.585000 ;
      RECT  9.955000  0.585000 10.535000 0.755000 ;
      RECT  9.955000  4.685000 10.535000 4.855000 ;
      RECT  9.955000  4.855000 10.205000 5.110000 ;
      RECT 10.000000  1.465000 10.780000 1.475000 ;
      RECT 10.000000  1.475000 10.430000 1.635000 ;
      RECT 10.000000  1.635000 10.330000 2.465000 ;
      RECT 10.000000  2.975000 10.330000 3.805000 ;
      RECT 10.000000  3.805000 10.430000 3.965000 ;
      RECT 10.000000  3.965000 10.780000 3.975000 ;
      RECT 10.260000  1.305000 10.780000 1.465000 ;
      RECT 10.260000  3.975000 10.780000 4.135000 ;
      RECT 10.365000  0.755000 10.535000 1.205000 ;
      RECT 10.365000  1.205000 10.780000 1.305000 ;
      RECT 10.365000  4.135000 10.780000 4.235000 ;
      RECT 10.365000  4.235000 10.535000 4.685000 ;
      RECT 10.600000  1.645000 10.770000 2.295000 ;
      RECT 10.600000  2.295000 10.955000 2.465000 ;
      RECT 10.600000  2.975000 10.955000 3.145000 ;
      RECT 10.600000  3.145000 10.770000 3.795000 ;
      RECT 10.705000  0.255000 11.850000 0.425000 ;
      RECT 10.705000  0.425000 10.875000 0.770000 ;
      RECT 10.705000  4.670000 10.875000 5.015000 ;
      RECT 10.705000  5.015000 11.850000 5.185000 ;
      RECT 10.985000  1.755000 11.415000 2.125000 ;
      RECT 10.985000  3.315000 11.415000 3.685000 ;
      RECT 11.045000  0.595000 11.375000 0.885000 ;
      RECT 11.045000  4.555000 11.375000 4.845000 ;
      RECT 11.125000  0.885000 11.295000 1.755000 ;
      RECT 11.125000  2.125000 11.295000 3.315000 ;
      RECT 11.125000  3.685000 11.295000 4.555000 ;
      RECT 11.465000  2.295000 11.765000 2.465000 ;
      RECT 11.465000  2.635000 14.295000 2.805000 ;
      RECT 11.465000  2.975000 11.765000 3.145000 ;
      RECT 11.545000  0.425000 11.850000 0.715000 ;
      RECT 11.545000  0.715000 12.735000 0.885000 ;
      RECT 11.545000  0.885000 11.850000 0.925000 ;
      RECT 11.545000  4.515000 11.850000 4.555000 ;
      RECT 11.545000  4.555000 12.735000 4.725000 ;
      RECT 11.545000  4.725000 11.850000 5.015000 ;
      RECT 11.595000  1.495000 12.785000 1.665000 ;
      RECT 11.595000  1.665000 11.765000 2.295000 ;
      RECT 11.595000  3.145000 11.765000 3.775000 ;
      RECT 11.595000  3.775000 12.785000 3.945000 ;
      RECT 11.985000  1.835000 12.315000 2.105000 ;
      RECT 11.985000  2.105000 12.285000 2.635000 ;
      RECT 11.985000  2.805000 12.285000 3.335000 ;
      RECT 11.985000  3.335000 12.315000 3.605000 ;
      RECT 12.020000  0.085000 12.235000 0.545000 ;
      RECT 12.020000  4.895000 12.235000 5.355000 ;
      RECT 12.405000  0.255000 12.735000 0.715000 ;
      RECT 12.405000  4.725000 12.735000 5.185000 ;
      RECT 12.455000  2.210000 12.785000 2.465000 ;
      RECT 12.455000  2.975000 12.785000 3.230000 ;
      RECT 12.485000  1.665000 12.785000 2.210000 ;
      RECT 12.485000  3.230000 12.785000 3.775000 ;
      RECT 12.975000  1.495000 14.165000 1.665000 ;
      RECT 12.975000  1.665000 13.275000 2.210000 ;
      RECT 12.975000  2.210000 13.305000 2.465000 ;
      RECT 12.975000  2.975000 13.305000 3.230000 ;
      RECT 12.975000  3.230000 13.275000 3.775000 ;
      RECT 12.975000  3.775000 14.165000 3.945000 ;
      RECT 13.025000  0.255000 13.355000 0.715000 ;
      RECT 13.025000  0.715000 14.215000 0.885000 ;
      RECT 13.025000  4.555000 14.215000 4.725000 ;
      RECT 13.025000  4.725000 13.355000 5.185000 ;
      RECT 13.445000  1.835000 13.775000 2.105000 ;
      RECT 13.445000  3.335000 13.775000 3.605000 ;
      RECT 13.475000  2.105000 13.775000 2.635000 ;
      RECT 13.475000  2.805000 13.775000 3.335000 ;
      RECT 13.525000  0.085000 13.740000 0.545000 ;
      RECT 13.525000  4.895000 13.740000 5.355000 ;
      RECT 13.910000  0.255000 15.055000 0.425000 ;
      RECT 13.910000  0.425000 14.215000 0.715000 ;
      RECT 13.910000  0.885000 14.215000 0.925000 ;
      RECT 13.910000  4.515000 14.215000 4.555000 ;
      RECT 13.910000  4.725000 14.215000 5.015000 ;
      RECT 13.910000  5.015000 15.055000 5.185000 ;
      RECT 13.995000  1.665000 14.165000 2.295000 ;
      RECT 13.995000  2.295000 14.295000 2.465000 ;
      RECT 13.995000  2.975000 14.295000 3.145000 ;
      RECT 13.995000  3.145000 14.165000 3.775000 ;
      RECT 14.345000  1.755000 14.775000 2.125000 ;
      RECT 14.345000  3.315000 14.775000 3.685000 ;
      RECT 14.385000  0.595000 14.715000 0.885000 ;
      RECT 14.385000  4.555000 14.715000 4.845000 ;
      RECT 14.465000  0.885000 14.635000 1.755000 ;
      RECT 14.465000  2.125000 14.635000 3.315000 ;
      RECT 14.465000  3.685000 14.635000 4.555000 ;
      RECT 14.805000  2.295000 15.160000 2.465000 ;
      RECT 14.805000  2.635000 17.395000 2.805000 ;
      RECT 14.805000  2.975000 15.160000 3.145000 ;
      RECT 14.885000  0.425000 15.055000 0.770000 ;
      RECT 14.885000  4.670000 15.055000 5.015000 ;
      RECT 14.980000  1.205000 15.395000 1.305000 ;
      RECT 14.980000  1.305000 15.500000 1.465000 ;
      RECT 14.980000  1.465000 15.760000 1.475000 ;
      RECT 14.980000  3.965000 15.760000 3.975000 ;
      RECT 14.980000  3.975000 15.500000 4.135000 ;
      RECT 14.980000  4.135000 15.395000 4.235000 ;
      RECT 14.990000  1.645000 15.160000 2.295000 ;
      RECT 14.990000  3.145000 15.160000 3.795000 ;
      RECT 15.225000  0.585000 15.805000 0.755000 ;
      RECT 15.225000  0.755000 15.395000 1.205000 ;
      RECT 15.225000  4.235000 15.395000 4.685000 ;
      RECT 15.225000  4.685000 15.805000 4.855000 ;
      RECT 15.330000  1.475000 15.760000 1.635000 ;
      RECT 15.330000  3.805000 15.760000 3.965000 ;
      RECT 15.430000  1.635000 15.760000 2.465000 ;
      RECT 15.430000  2.975000 15.760000 3.805000 ;
      RECT 15.555000  0.330000 15.805000 0.585000 ;
      RECT 15.555000  4.855000 15.805000 5.110000 ;
      RECT 15.935000  1.465000 16.265000 2.635000 ;
      RECT 15.935000  2.805000 16.265000 3.975000 ;
      RECT 15.975000  0.085000 16.225000 0.660000 ;
      RECT 15.975000  4.780000 16.225000 5.355000 ;
      RECT 16.395000  0.330000 16.645000 0.585000 ;
      RECT 16.395000  0.585000 16.975000 0.755000 ;
      RECT 16.395000  4.685000 16.975000 4.855000 ;
      RECT 16.395000  4.855000 16.645000 5.110000 ;
      RECT 16.440000  1.465000 17.220000 1.475000 ;
      RECT 16.440000  1.475000 16.870000 1.635000 ;
      RECT 16.440000  1.635000 16.770000 2.465000 ;
      RECT 16.440000  2.975000 16.770000 3.805000 ;
      RECT 16.440000  3.805000 16.870000 3.965000 ;
      RECT 16.440000  3.965000 17.220000 3.975000 ;
      RECT 16.700000  1.305000 17.220000 1.465000 ;
      RECT 16.700000  3.975000 17.220000 4.135000 ;
      RECT 16.805000  0.755000 16.975000 1.205000 ;
      RECT 16.805000  1.205000 17.220000 1.305000 ;
      RECT 16.805000  4.135000 17.220000 4.235000 ;
      RECT 16.805000  4.235000 16.975000 4.685000 ;
      RECT 17.040000  1.645000 17.210000 2.295000 ;
      RECT 17.040000  2.295000 17.395000 2.465000 ;
      RECT 17.040000  2.975000 17.395000 3.145000 ;
      RECT 17.040000  3.145000 17.210000 3.795000 ;
      RECT 17.145000  0.255000 18.290000 0.425000 ;
      RECT 17.145000  0.425000 17.315000 0.770000 ;
      RECT 17.145000  4.670000 17.315000 5.015000 ;
      RECT 17.145000  5.015000 18.290000 5.185000 ;
      RECT 17.425000  1.755000 17.855000 2.125000 ;
      RECT 17.425000  3.315000 17.855000 3.685000 ;
      RECT 17.485000  0.595000 17.815000 0.885000 ;
      RECT 17.485000  4.555000 17.815000 4.845000 ;
      RECT 17.565000  0.885000 17.735000 1.755000 ;
      RECT 17.565000  2.125000 17.735000 3.315000 ;
      RECT 17.565000  3.685000 17.735000 4.555000 ;
      RECT 17.905000  2.295000 18.205000 2.465000 ;
      RECT 17.905000  2.635000 20.735000 2.805000 ;
      RECT 17.905000  2.975000 18.205000 3.145000 ;
      RECT 17.985000  0.425000 18.290000 0.715000 ;
      RECT 17.985000  0.715000 19.175000 0.885000 ;
      RECT 17.985000  0.885000 18.290000 0.925000 ;
      RECT 17.985000  4.515000 18.290000 4.555000 ;
      RECT 17.985000  4.555000 19.175000 4.725000 ;
      RECT 17.985000  4.725000 18.290000 5.015000 ;
      RECT 18.035000  1.495000 19.225000 1.665000 ;
      RECT 18.035000  1.665000 18.205000 2.295000 ;
      RECT 18.035000  3.145000 18.205000 3.775000 ;
      RECT 18.035000  3.775000 19.225000 3.945000 ;
      RECT 18.425000  1.835000 18.755000 2.105000 ;
      RECT 18.425000  2.105000 18.725000 2.635000 ;
      RECT 18.425000  2.805000 18.725000 3.335000 ;
      RECT 18.425000  3.335000 18.755000 3.605000 ;
      RECT 18.460000  0.085000 18.675000 0.545000 ;
      RECT 18.460000  4.895000 18.675000 5.355000 ;
      RECT 18.845000  0.255000 19.175000 0.715000 ;
      RECT 18.845000  4.725000 19.175000 5.185000 ;
      RECT 18.895000  2.210000 19.225000 2.465000 ;
      RECT 18.895000  2.975000 19.225000 3.230000 ;
      RECT 18.925000  1.665000 19.225000 2.210000 ;
      RECT 18.925000  3.230000 19.225000 3.775000 ;
      RECT 19.415000  1.495000 20.605000 1.665000 ;
      RECT 19.415000  1.665000 19.715000 2.210000 ;
      RECT 19.415000  2.210000 19.745000 2.465000 ;
      RECT 19.415000  2.975000 19.745000 3.230000 ;
      RECT 19.415000  3.230000 19.715000 3.775000 ;
      RECT 19.415000  3.775000 20.605000 3.945000 ;
      RECT 19.465000  0.255000 19.795000 0.715000 ;
      RECT 19.465000  0.715000 20.655000 0.885000 ;
      RECT 19.465000  4.555000 20.655000 4.725000 ;
      RECT 19.465000  4.725000 19.795000 5.185000 ;
      RECT 19.885000  1.835000 20.215000 2.105000 ;
      RECT 19.885000  3.335000 20.215000 3.605000 ;
      RECT 19.915000  2.105000 20.215000 2.635000 ;
      RECT 19.915000  2.805000 20.215000 3.335000 ;
      RECT 19.965000  0.085000 20.180000 0.545000 ;
      RECT 19.965000  4.895000 20.180000 5.355000 ;
      RECT 20.350000  0.255000 21.495000 0.425000 ;
      RECT 20.350000  0.425000 20.655000 0.715000 ;
      RECT 20.350000  0.885000 20.655000 0.925000 ;
      RECT 20.350000  4.515000 20.655000 4.555000 ;
      RECT 20.350000  4.725000 20.655000 5.015000 ;
      RECT 20.350000  5.015000 21.495000 5.185000 ;
      RECT 20.435000  1.665000 20.605000 2.295000 ;
      RECT 20.435000  2.295000 20.735000 2.465000 ;
      RECT 20.435000  2.975000 20.735000 3.145000 ;
      RECT 20.435000  3.145000 20.605000 3.775000 ;
      RECT 20.785000  1.755000 21.215000 2.125000 ;
      RECT 20.785000  3.315000 21.215000 3.685000 ;
      RECT 20.825000  0.595000 21.155000 0.885000 ;
      RECT 20.825000  4.555000 21.155000 4.845000 ;
      RECT 20.905000  0.885000 21.075000 1.755000 ;
      RECT 20.905000  2.125000 21.075000 3.315000 ;
      RECT 20.905000  3.685000 21.075000 4.555000 ;
      RECT 21.245000  2.295000 21.600000 2.465000 ;
      RECT 21.245000  2.635000 23.835000 2.805000 ;
      RECT 21.245000  2.975000 21.600000 3.145000 ;
      RECT 21.325000  0.425000 21.495000 0.770000 ;
      RECT 21.325000  4.670000 21.495000 5.015000 ;
      RECT 21.420000  1.205000 21.835000 1.305000 ;
      RECT 21.420000  1.305000 21.940000 1.465000 ;
      RECT 21.420000  1.465000 22.200000 1.475000 ;
      RECT 21.420000  3.965000 22.200000 3.975000 ;
      RECT 21.420000  3.975000 21.940000 4.135000 ;
      RECT 21.420000  4.135000 21.835000 4.235000 ;
      RECT 21.430000  1.645000 21.600000 2.295000 ;
      RECT 21.430000  3.145000 21.600000 3.795000 ;
      RECT 21.665000  0.585000 22.245000 0.755000 ;
      RECT 21.665000  0.755000 21.835000 1.205000 ;
      RECT 21.665000  4.235000 21.835000 4.685000 ;
      RECT 21.665000  4.685000 22.245000 4.855000 ;
      RECT 21.770000  1.475000 22.200000 1.635000 ;
      RECT 21.770000  3.805000 22.200000 3.965000 ;
      RECT 21.870000  1.635000 22.200000 2.465000 ;
      RECT 21.870000  2.975000 22.200000 3.805000 ;
      RECT 21.995000  0.330000 22.245000 0.585000 ;
      RECT 21.995000  4.855000 22.245000 5.110000 ;
      RECT 22.375000  1.465000 22.705000 2.635000 ;
      RECT 22.375000  2.805000 22.705000 3.975000 ;
      RECT 22.415000  0.085000 22.665000 0.660000 ;
      RECT 22.415000  4.780000 22.665000 5.355000 ;
      RECT 22.835000  0.330000 23.085000 0.585000 ;
      RECT 22.835000  0.585000 23.415000 0.755000 ;
      RECT 22.835000  4.685000 23.415000 4.855000 ;
      RECT 22.835000  4.855000 23.085000 5.110000 ;
      RECT 22.880000  1.465000 23.660000 1.475000 ;
      RECT 22.880000  1.475000 23.310000 1.635000 ;
      RECT 22.880000  1.635000 23.210000 2.465000 ;
      RECT 22.880000  2.975000 23.210000 3.805000 ;
      RECT 22.880000  3.805000 23.310000 3.965000 ;
      RECT 22.880000  3.965000 23.660000 3.975000 ;
      RECT 23.140000  1.305000 23.660000 1.465000 ;
      RECT 23.140000  3.975000 23.660000 4.135000 ;
      RECT 23.245000  0.755000 23.415000 1.205000 ;
      RECT 23.245000  1.205000 23.660000 1.305000 ;
      RECT 23.245000  4.135000 23.660000 4.235000 ;
      RECT 23.245000  4.235000 23.415000 4.685000 ;
      RECT 23.480000  1.645000 23.650000 2.295000 ;
      RECT 23.480000  2.295000 23.835000 2.465000 ;
      RECT 23.480000  2.975000 23.835000 3.145000 ;
      RECT 23.480000  3.145000 23.650000 3.795000 ;
      RECT 23.585000  0.255000 24.730000 0.425000 ;
      RECT 23.585000  0.425000 23.755000 0.770000 ;
      RECT 23.585000  4.670000 23.755000 5.015000 ;
      RECT 23.585000  5.015000 24.730000 5.185000 ;
      RECT 23.865000  1.755000 24.295000 2.125000 ;
      RECT 23.865000  3.315000 24.295000 3.685000 ;
      RECT 23.925000  0.595000 24.255000 0.885000 ;
      RECT 23.925000  4.555000 24.255000 4.845000 ;
      RECT 24.005000  0.885000 24.175000 1.755000 ;
      RECT 24.005000  2.125000 24.175000 3.315000 ;
      RECT 24.005000  3.685000 24.175000 4.555000 ;
      RECT 24.345000  2.295000 24.645000 2.465000 ;
      RECT 24.345000  2.635000 25.760000 2.805000 ;
      RECT 24.345000  2.975000 24.645000 3.145000 ;
      RECT 24.425000  0.425000 24.730000 0.715000 ;
      RECT 24.425000  0.715000 25.615000 0.885000 ;
      RECT 24.425000  0.885000 24.730000 0.925000 ;
      RECT 24.425000  4.515000 24.730000 4.555000 ;
      RECT 24.425000  4.555000 25.615000 4.725000 ;
      RECT 24.425000  4.725000 24.730000 5.015000 ;
      RECT 24.475000  1.495000 25.665000 1.665000 ;
      RECT 24.475000  1.665000 24.645000 2.295000 ;
      RECT 24.475000  3.145000 24.645000 3.775000 ;
      RECT 24.475000  3.775000 25.665000 3.945000 ;
      RECT 24.865000  1.835000 25.195000 2.105000 ;
      RECT 24.865000  2.105000 25.165000 2.635000 ;
      RECT 24.865000  2.805000 25.165000 3.335000 ;
      RECT 24.865000  3.335000 25.195000 3.605000 ;
      RECT 24.900000  0.085000 25.115000 0.545000 ;
      RECT 24.900000  4.895000 25.115000 5.355000 ;
      RECT 25.285000  0.255000 25.615000 0.715000 ;
      RECT 25.285000  4.725000 25.615000 5.185000 ;
      RECT 25.335000  2.210000 25.665000 2.465000 ;
      RECT 25.335000  2.975000 25.665000 3.230000 ;
      RECT 25.365000  1.665000 25.665000 2.210000 ;
      RECT 25.365000  3.230000 25.665000 3.775000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.145000  5.355000  0.315000 5.525000 ;
      RECT  0.175000  2.140000  0.345000 2.310000 ;
      RECT  0.175000  3.130000  0.345000 3.300000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.605000  5.355000  0.775000 5.525000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.065000  5.355000  1.235000 5.525000 ;
      RECT  1.115000  2.140000  1.285000 2.310000 ;
      RECT  1.115000  3.130000  1.285000 3.300000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  1.785000  1.695000 1.955000 ;
      RECT  1.525000  3.485000  1.695000 3.655000 ;
      RECT  1.525000  5.355000  1.695000 5.525000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  1.985000  5.355000  2.155000 5.525000 ;
      RECT  2.110000  2.140000  2.280000 2.310000 ;
      RECT  2.110000  3.130000  2.280000 3.300000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.445000  5.355000  2.615000 5.525000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  2.905000  5.355000  3.075000 5.525000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.365000  5.355000  3.535000 5.525000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  3.825000  5.355000  3.995000 5.525000 ;
      RECT  4.160000  2.140000  4.330000 2.310000 ;
      RECT  4.160000  3.130000  4.330000 3.300000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.285000  5.355000  4.455000 5.525000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.785000  4.915000 1.955000 ;
      RECT  4.745000  3.485000  4.915000 3.655000 ;
      RECT  4.745000  5.355000  4.915000 5.525000 ;
      RECT  5.155000  2.140000  5.325000 2.310000 ;
      RECT  5.155000  3.130000  5.325000 3.300000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.205000  5.355000  5.375000 5.525000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.665000  5.355000  5.835000 5.525000 ;
      RECT  6.095000  2.140000  6.265000 2.310000 ;
      RECT  6.095000  3.130000  6.265000 3.300000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.125000  5.355000  6.295000 5.525000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  6.585000  5.355000  6.755000 5.525000 ;
      RECT  6.615000  2.140000  6.785000 2.310000 ;
      RECT  6.615000  3.130000  6.785000 3.300000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.045000  5.355000  7.215000 5.525000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.505000  5.355000  7.675000 5.525000 ;
      RECT  7.555000  2.140000  7.725000 2.310000 ;
      RECT  7.555000  3.130000  7.725000 3.300000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  1.785000  8.135000 1.955000 ;
      RECT  7.965000  3.485000  8.135000 3.655000 ;
      RECT  7.965000  5.355000  8.135000 5.525000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.425000  5.355000  8.595000 5.525000 ;
      RECT  8.550000  2.140000  8.720000 2.310000 ;
      RECT  8.550000  3.130000  8.720000 3.300000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  8.885000  5.355000  9.055000 5.525000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.345000  5.355000  9.515000 5.525000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT  9.805000  5.355000  9.975000 5.525000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.265000  5.355000 10.435000 5.525000 ;
      RECT 10.600000  2.140000 10.770000 2.310000 ;
      RECT 10.600000  3.130000 10.770000 3.300000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 10.725000  5.355000 10.895000 5.525000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  1.785000 11.355000 1.955000 ;
      RECT 11.185000  3.485000 11.355000 3.655000 ;
      RECT 11.185000  5.355000 11.355000 5.525000 ;
      RECT 11.595000  2.140000 11.765000 2.310000 ;
      RECT 11.595000  3.130000 11.765000 3.300000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 11.645000  5.355000 11.815000 5.525000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.105000  5.355000 12.275000 5.525000 ;
      RECT 12.535000  2.140000 12.705000 2.310000 ;
      RECT 12.535000  3.130000 12.705000 3.300000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 12.565000  5.355000 12.735000 5.525000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.025000  5.355000 13.195000 5.525000 ;
      RECT 13.055000  2.140000 13.225000 2.310000 ;
      RECT 13.055000  3.130000 13.225000 3.300000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.485000  5.355000 13.655000 5.525000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 13.945000  5.355000 14.115000 5.525000 ;
      RECT 13.995000  2.140000 14.165000 2.310000 ;
      RECT 13.995000  3.130000 14.165000 3.300000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  1.785000 14.575000 1.955000 ;
      RECT 14.405000  3.485000 14.575000 3.655000 ;
      RECT 14.405000  5.355000 14.575000 5.525000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 14.865000  5.355000 15.035000 5.525000 ;
      RECT 14.990000  2.140000 15.160000 2.310000 ;
      RECT 14.990000  3.130000 15.160000 3.300000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.325000  5.355000 15.495000 5.525000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
      RECT 15.785000  5.355000 15.955000 5.525000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
      RECT 16.245000  5.355000 16.415000 5.525000 ;
      RECT 16.705000 -0.085000 16.875000 0.085000 ;
      RECT 16.705000  2.635000 16.875000 2.805000 ;
      RECT 16.705000  5.355000 16.875000 5.525000 ;
      RECT 17.040000  2.140000 17.210000 2.310000 ;
      RECT 17.040000  3.130000 17.210000 3.300000 ;
      RECT 17.165000 -0.085000 17.335000 0.085000 ;
      RECT 17.165000  2.635000 17.335000 2.805000 ;
      RECT 17.165000  5.355000 17.335000 5.525000 ;
      RECT 17.625000 -0.085000 17.795000 0.085000 ;
      RECT 17.625000  1.785000 17.795000 1.955000 ;
      RECT 17.625000  3.485000 17.795000 3.655000 ;
      RECT 17.625000  5.355000 17.795000 5.525000 ;
      RECT 18.035000  2.140000 18.205000 2.310000 ;
      RECT 18.035000  3.130000 18.205000 3.300000 ;
      RECT 18.085000 -0.085000 18.255000 0.085000 ;
      RECT 18.085000  2.635000 18.255000 2.805000 ;
      RECT 18.085000  5.355000 18.255000 5.525000 ;
      RECT 18.545000 -0.085000 18.715000 0.085000 ;
      RECT 18.545000  2.635000 18.715000 2.805000 ;
      RECT 18.545000  5.355000 18.715000 5.525000 ;
      RECT 18.975000  2.140000 19.145000 2.310000 ;
      RECT 18.975000  3.130000 19.145000 3.300000 ;
      RECT 19.005000 -0.085000 19.175000 0.085000 ;
      RECT 19.005000  2.635000 19.175000 2.805000 ;
      RECT 19.005000  5.355000 19.175000 5.525000 ;
      RECT 19.465000 -0.085000 19.635000 0.085000 ;
      RECT 19.465000  2.635000 19.635000 2.805000 ;
      RECT 19.465000  5.355000 19.635000 5.525000 ;
      RECT 19.495000  2.140000 19.665000 2.310000 ;
      RECT 19.495000  3.130000 19.665000 3.300000 ;
      RECT 19.925000 -0.085000 20.095000 0.085000 ;
      RECT 19.925000  2.635000 20.095000 2.805000 ;
      RECT 19.925000  5.355000 20.095000 5.525000 ;
      RECT 20.385000 -0.085000 20.555000 0.085000 ;
      RECT 20.385000  2.635000 20.555000 2.805000 ;
      RECT 20.385000  5.355000 20.555000 5.525000 ;
      RECT 20.435000  2.140000 20.605000 2.310000 ;
      RECT 20.435000  3.130000 20.605000 3.300000 ;
      RECT 20.845000 -0.085000 21.015000 0.085000 ;
      RECT 20.845000  1.785000 21.015000 1.955000 ;
      RECT 20.845000  3.485000 21.015000 3.655000 ;
      RECT 20.845000  5.355000 21.015000 5.525000 ;
      RECT 21.305000 -0.085000 21.475000 0.085000 ;
      RECT 21.305000  2.635000 21.475000 2.805000 ;
      RECT 21.305000  5.355000 21.475000 5.525000 ;
      RECT 21.430000  2.140000 21.600000 2.310000 ;
      RECT 21.430000  3.130000 21.600000 3.300000 ;
      RECT 21.765000 -0.085000 21.935000 0.085000 ;
      RECT 21.765000  2.635000 21.935000 2.805000 ;
      RECT 21.765000  5.355000 21.935000 5.525000 ;
      RECT 22.225000 -0.085000 22.395000 0.085000 ;
      RECT 22.225000  2.635000 22.395000 2.805000 ;
      RECT 22.225000  5.355000 22.395000 5.525000 ;
      RECT 22.685000 -0.085000 22.855000 0.085000 ;
      RECT 22.685000  2.635000 22.855000 2.805000 ;
      RECT 22.685000  5.355000 22.855000 5.525000 ;
      RECT 23.145000 -0.085000 23.315000 0.085000 ;
      RECT 23.145000  2.635000 23.315000 2.805000 ;
      RECT 23.145000  5.355000 23.315000 5.525000 ;
      RECT 23.480000  2.140000 23.650000 2.310000 ;
      RECT 23.480000  3.130000 23.650000 3.300000 ;
      RECT 23.605000 -0.085000 23.775000 0.085000 ;
      RECT 23.605000  2.635000 23.775000 2.805000 ;
      RECT 23.605000  5.355000 23.775000 5.525000 ;
      RECT 24.065000 -0.085000 24.235000 0.085000 ;
      RECT 24.065000  1.785000 24.235000 1.955000 ;
      RECT 24.065000  3.485000 24.235000 3.655000 ;
      RECT 24.065000  5.355000 24.235000 5.525000 ;
      RECT 24.475000  2.140000 24.645000 2.310000 ;
      RECT 24.475000  3.130000 24.645000 3.300000 ;
      RECT 24.525000 -0.085000 24.695000 0.085000 ;
      RECT 24.525000  2.635000 24.695000 2.805000 ;
      RECT 24.525000  5.355000 24.695000 5.525000 ;
      RECT 24.985000 -0.085000 25.155000 0.085000 ;
      RECT 24.985000  2.635000 25.155000 2.805000 ;
      RECT 24.985000  5.355000 25.155000 5.525000 ;
      RECT 25.415000  2.140000 25.585000 2.310000 ;
      RECT 25.415000  3.130000 25.585000 3.300000 ;
      RECT 25.445000 -0.085000 25.615000 0.085000 ;
      RECT 25.445000  2.635000 25.615000 2.805000 ;
      RECT 25.445000  5.355000 25.615000 5.525000 ;
    LAYER met1 ;
      RECT  0.115000 2.110000  0.405000 2.155000 ;
      RECT  0.115000 2.155000  2.340000 2.295000 ;
      RECT  0.115000 2.295000  0.405000 2.340000 ;
      RECT  0.115000 3.100000  0.405000 3.145000 ;
      RECT  0.115000 3.145000  2.340000 3.285000 ;
      RECT  0.115000 3.285000  0.405000 3.330000 ;
      RECT  1.055000 2.110000  1.345000 2.155000 ;
      RECT  1.055000 2.295000  1.345000 2.340000 ;
      RECT  1.055000 3.100000  1.345000 3.145000 ;
      RECT  1.055000 3.285000  1.345000 3.330000 ;
      RECT  2.050000 2.110000  2.340000 2.155000 ;
      RECT  2.050000 2.295000  2.340000 2.340000 ;
      RECT  2.050000 3.100000  2.340000 3.145000 ;
      RECT  2.050000 3.285000  2.340000 3.330000 ;
      RECT  4.100000 2.110000  4.390000 2.155000 ;
      RECT  4.100000 2.155000  6.325000 2.295000 ;
      RECT  4.100000 2.295000  4.390000 2.340000 ;
      RECT  4.100000 3.100000  4.390000 3.145000 ;
      RECT  4.100000 3.145000  6.325000 3.285000 ;
      RECT  4.100000 3.285000  4.390000 3.330000 ;
      RECT  5.095000 2.110000  5.385000 2.155000 ;
      RECT  5.095000 2.295000  5.385000 2.340000 ;
      RECT  5.095000 3.100000  5.385000 3.145000 ;
      RECT  5.095000 3.285000  5.385000 3.330000 ;
      RECT  6.035000 2.110000  6.325000 2.155000 ;
      RECT  6.035000 2.295000  6.325000 2.340000 ;
      RECT  6.035000 3.100000  6.325000 3.145000 ;
      RECT  6.035000 3.285000  6.325000 3.330000 ;
      RECT  6.555000 2.110000  6.845000 2.155000 ;
      RECT  6.555000 2.155000  8.780000 2.295000 ;
      RECT  6.555000 2.295000  6.845000 2.340000 ;
      RECT  6.555000 3.100000  6.845000 3.145000 ;
      RECT  6.555000 3.145000  8.780000 3.285000 ;
      RECT  6.555000 3.285000  6.845000 3.330000 ;
      RECT  7.495000 2.110000  7.785000 2.155000 ;
      RECT  7.495000 2.295000  7.785000 2.340000 ;
      RECT  7.495000 3.100000  7.785000 3.145000 ;
      RECT  7.495000 3.285000  7.785000 3.330000 ;
      RECT  8.490000 2.110000  8.780000 2.155000 ;
      RECT  8.490000 2.295000  8.780000 2.340000 ;
      RECT  8.490000 3.100000  8.780000 3.145000 ;
      RECT  8.490000 3.285000  8.780000 3.330000 ;
      RECT 10.540000 2.110000 10.830000 2.155000 ;
      RECT 10.540000 2.155000 12.765000 2.295000 ;
      RECT 10.540000 2.295000 10.830000 2.340000 ;
      RECT 10.540000 3.100000 10.830000 3.145000 ;
      RECT 10.540000 3.145000 12.765000 3.285000 ;
      RECT 10.540000 3.285000 10.830000 3.330000 ;
      RECT 11.535000 2.110000 11.825000 2.155000 ;
      RECT 11.535000 2.295000 11.825000 2.340000 ;
      RECT 11.535000 3.100000 11.825000 3.145000 ;
      RECT 11.535000 3.285000 11.825000 3.330000 ;
      RECT 12.475000 2.110000 12.765000 2.155000 ;
      RECT 12.475000 2.295000 12.765000 2.340000 ;
      RECT 12.475000 3.100000 12.765000 3.145000 ;
      RECT 12.475000 3.285000 12.765000 3.330000 ;
      RECT 12.995000 2.110000 13.285000 2.155000 ;
      RECT 12.995000 2.155000 15.220000 2.295000 ;
      RECT 12.995000 2.295000 13.285000 2.340000 ;
      RECT 12.995000 3.100000 13.285000 3.145000 ;
      RECT 12.995000 3.145000 15.220000 3.285000 ;
      RECT 12.995000 3.285000 13.285000 3.330000 ;
      RECT 13.935000 2.110000 14.225000 2.155000 ;
      RECT 13.935000 2.295000 14.225000 2.340000 ;
      RECT 13.935000 3.100000 14.225000 3.145000 ;
      RECT 13.935000 3.285000 14.225000 3.330000 ;
      RECT 14.930000 2.110000 15.220000 2.155000 ;
      RECT 14.930000 2.295000 15.220000 2.340000 ;
      RECT 14.930000 3.100000 15.220000 3.145000 ;
      RECT 14.930000 3.285000 15.220000 3.330000 ;
      RECT 16.980000 2.110000 17.270000 2.155000 ;
      RECT 16.980000 2.155000 19.205000 2.295000 ;
      RECT 16.980000 2.295000 17.270000 2.340000 ;
      RECT 16.980000 3.100000 17.270000 3.145000 ;
      RECT 16.980000 3.145000 19.205000 3.285000 ;
      RECT 16.980000 3.285000 17.270000 3.330000 ;
      RECT 17.975000 2.110000 18.265000 2.155000 ;
      RECT 17.975000 2.295000 18.265000 2.340000 ;
      RECT 17.975000 3.100000 18.265000 3.145000 ;
      RECT 17.975000 3.285000 18.265000 3.330000 ;
      RECT 18.915000 2.110000 19.205000 2.155000 ;
      RECT 18.915000 2.295000 19.205000 2.340000 ;
      RECT 18.915000 3.100000 19.205000 3.145000 ;
      RECT 18.915000 3.285000 19.205000 3.330000 ;
      RECT 19.435000 2.110000 19.725000 2.155000 ;
      RECT 19.435000 2.155000 21.660000 2.295000 ;
      RECT 19.435000 2.295000 19.725000 2.340000 ;
      RECT 19.435000 3.100000 19.725000 3.145000 ;
      RECT 19.435000 3.145000 21.660000 3.285000 ;
      RECT 19.435000 3.285000 19.725000 3.330000 ;
      RECT 20.375000 2.110000 20.665000 2.155000 ;
      RECT 20.375000 2.295000 20.665000 2.340000 ;
      RECT 20.375000 3.100000 20.665000 3.145000 ;
      RECT 20.375000 3.285000 20.665000 3.330000 ;
      RECT 21.370000 2.110000 21.660000 2.155000 ;
      RECT 21.370000 2.295000 21.660000 2.340000 ;
      RECT 21.370000 3.100000 21.660000 3.145000 ;
      RECT 21.370000 3.285000 21.660000 3.330000 ;
      RECT 23.420000 2.110000 23.710000 2.155000 ;
      RECT 23.420000 2.155000 25.645000 2.295000 ;
      RECT 23.420000 2.295000 23.710000 2.340000 ;
      RECT 23.420000 3.100000 23.710000 3.145000 ;
      RECT 23.420000 3.145000 25.645000 3.285000 ;
      RECT 23.420000 3.285000 23.710000 3.330000 ;
      RECT 24.415000 2.110000 24.705000 2.155000 ;
      RECT 24.415000 2.295000 24.705000 2.340000 ;
      RECT 24.415000 3.100000 24.705000 3.145000 ;
      RECT 24.415000 3.285000 24.705000 3.330000 ;
      RECT 25.355000 2.110000 25.645000 2.155000 ;
      RECT 25.355000 2.295000 25.645000 2.340000 ;
      RECT 25.355000 3.100000 25.645000 3.145000 ;
      RECT 25.355000 3.285000 25.645000 3.330000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb16to1_2
END LIBRARY
