# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__buf_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__buf_6 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.280000 1.075000 1.265000 1.315000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.526500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.845000 0.255000 2.015000 0.735000 ;
        RECT 1.845000 0.735000 3.895000 0.905000 ;
        RECT 1.845000 1.445000 3.895000 1.615000 ;
        RECT 1.845000 1.615000 2.015000 2.465000 ;
        RECT 2.410000 0.905000 3.895000 1.445000 ;
        RECT 2.785000 0.255000 2.955000 0.735000 ;
        RECT 2.785000 1.615000 2.955000 2.465000 ;
        RECT 3.725000 0.255000 3.895000 0.735000 ;
        RECT 3.725000 1.615000 3.895000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.600000 0.085000 ;
        RECT 0.435000  0.085000 0.605000 0.565000 ;
        RECT 1.375000  0.085000 1.545000 0.565000 ;
        RECT 2.185000  0.085000 2.565000 0.565000 ;
        RECT 3.125000  0.085000 3.505000 0.565000 ;
        RECT 4.065000  0.085000 4.445000 0.885000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 4.600000 2.805000 ;
        RECT 0.435000 1.485000 0.605000 2.635000 ;
        RECT 1.375000 1.835000 1.615000 2.635000 ;
        RECT 2.185000 1.835000 2.565000 2.635000 ;
        RECT 3.125000 1.835000 3.505000 2.635000 ;
        RECT 4.065000 1.485000 4.445000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.775000 0.255000 1.155000 0.735000 ;
      RECT 0.775000 0.735000 1.625000 0.905000 ;
      RECT 0.775000 1.485000 1.625000 1.655000 ;
      RECT 0.775000 1.655000 1.155000 2.465000 ;
      RECT 1.455000 0.905000 1.625000 1.075000 ;
      RECT 1.455000 1.075000 1.975000 1.245000 ;
      RECT 1.455000 1.245000 1.625000 1.485000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__buf_6
