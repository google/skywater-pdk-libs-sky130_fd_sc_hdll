* File: sky130_fd_sc_hdll__clkinvlp_2.pex.spice
* Created: Wed Sep  2 08:26:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKINVLP_2%A 5 7 9 10 14 16 18 19 20 21 25 26
r39 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.16 $X2=0.515 $Y2=1.16
r40 20 21 8.93773 $w=4.53e-07 $l=3.4e-07 $layer=LI1_cond $X=0.372 $Y=1.19
+ $X2=0.372 $Y2=1.53
r41 20 26 0.788623 $w=4.53e-07 $l=3e-08 $layer=LI1_cond $X=0.372 $Y=1.19
+ $X2=0.372 $Y2=1.16
r42 16 19 18.238 $w=2e-07 $l=1.09174e-07 $layer=POLY_cond $X=1.185 $Y=0.995
+ $X2=1.135 $Y2=1.082
r43 16 18 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.185 $Y=0.995
+ $X2=1.185 $Y2=0.61
r44 12 19 18.238 $w=2e-07 $l=8.8e-08 $layer=POLY_cond $X=1.135 $Y=1.17 $X2=1.135
+ $Y2=1.082
r45 12 14 202.49 $w=2.5e-07 $l=8.15e-07 $layer=POLY_cond $X=1.135 $Y=1.17
+ $X2=1.135 $Y2=1.985
r46 11 25 9.58664 $w=1.75e-07 $l=3.10467e-07 $layer=POLY_cond $X=0.75 $Y=1.082
+ $X2=0.48 $Y2=0.995
r47 10 19 7.22026 $w=1.75e-07 $l=1.25e-07 $layer=POLY_cond $X=1.01 $Y=1.082
+ $X2=1.135 $Y2=1.082
r48 10 11 103.952 $w=1.75e-07 $l=2.6e-07 $layer=POLY_cond $X=1.01 $Y=1.082
+ $X2=0.75 $Y2=1.082
r49 7 25 14.7117 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=0.675 $Y=0.995
+ $X2=0.48 $Y2=0.995
r50 7 9 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.675 $Y=0.995
+ $X2=0.675 $Y2=0.61
r51 3 25 14.7117 $w=2.5e-07 $l=3.77359e-07 $layer=POLY_cond $X=0.605 $Y=1.315
+ $X2=0.48 $Y2=0.995
r52 3 5 166.464 $w=2.5e-07 $l=6.7e-07 $layer=POLY_cond $X=0.605 $Y=1.315
+ $X2=0.605 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINVLP_2%VPWR 1 2 7 9 11 13 17 19 29
r21 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r22 23 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r23 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r24 20 25 4.39998 $w=1.8e-07 $l=2.78e-07 $layer=LI1_cond $X=0.555 $Y=2.715
+ $X2=0.277 $Y2=2.715
r25 20 22 36.6616 $w=1.78e-07 $l=5.95e-07 $layer=LI1_cond $X=0.555 $Y=2.715
+ $X2=1.15 $Y2=2.715
r26 19 28 3.91797 $w=1.8e-07 $l=2.17e-07 $layer=LI1_cond $X=1.405 $Y=2.715
+ $X2=1.622 $Y2=2.715
r27 19 22 15.7121 $w=1.78e-07 $l=2.55e-07 $layer=LI1_cond $X=1.405 $Y=2.715
+ $X2=1.15 $Y2=2.715
r28 17 23 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r29 17 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r30 13 16 31.4706 $w=2.58e-07 $l=7.1e-07 $layer=LI1_cond $X=1.535 $Y=1.63
+ $X2=1.535 $Y2=2.34
r31 11 28 3.19576 $w=2.6e-07 $l=1.26214e-07 $layer=LI1_cond $X=1.535 $Y=2.625
+ $X2=1.622 $Y2=2.715
r32 11 16 12.6325 $w=2.58e-07 $l=2.85e-07 $layer=LI1_cond $X=1.535 $Y=2.625
+ $X2=1.535 $Y2=2.34
r33 7 25 3.21294 $w=3.3e-07 $l=1.51456e-07 $layer=LI1_cond $X=0.39 $Y=2.625
+ $X2=0.277 $Y2=2.715
r34 7 9 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=0.39 $Y=2.625
+ $X2=0.39 $Y2=2
r35 2 16 400 $w=1.7e-07 $l=9.67587e-07 $layer=licon1_PDIFF $count=1 $X=1.26
+ $Y=1.485 $X2=1.5 $Y2=2.34
r36 2 13 400 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_PDIFF $count=1 $X=1.26
+ $Y=1.485 $X2=1.5 $Y2=1.63
r37 1 9 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.195
+ $Y=1.485 $X2=0.32 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINVLP_2%Y 1 2 7 8 9 25 27
r22 25 27 5.56352 $w=4.33e-07 $l=2.1e-07 $layer=LI1_cond $X=1.19 $Y=0.532
+ $X2=1.4 $Y2=0.532
r23 13 21 0.508694 $w=4.5e-07 $l=2.18e-07 $layer=LI1_cond $X=1.01 $Y=0.75
+ $X2=1.01 $Y2=0.532
r24 9 19 12.7582 $w=4.48e-07 $l=4.8e-07 $layer=LI1_cond $X=1.01 $Y=1.19 $X2=1.01
+ $Y2=1.67
r25 8 9 9.03704 $w=4.48e-07 $l=3.4e-07 $layer=LI1_cond $X=1.01 $Y=0.85 $X2=1.01
+ $Y2=1.19
r26 8 13 2.65795 $w=4.48e-07 $l=1e-07 $layer=LI1_cond $X=1.01 $Y=0.85 $X2=1.01
+ $Y2=0.75
r27 7 25 1.32465 $w=4.33e-07 $l=5e-08 $layer=LI1_cond $X=1.14 $Y=0.532 $X2=1.19
+ $Y2=0.532
r28 7 21 3.44408 $w=4.33e-07 $l=1.3e-07 $layer=LI1_cond $X=1.14 $Y=0.532
+ $X2=1.01 $Y2=0.532
r29 2 19 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=0.73
+ $Y=1.485 $X2=0.87 $Y2=1.67
r30 1 27 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.26
+ $Y=0.335 $X2=1.4 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINVLP_2%VGND 1 6 9 10 11 21 22
r16 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r17 19 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r18 18 21 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r19 18 19 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r20 11 19 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r21 11 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r22 9 14 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.295 $Y=0 $X2=0.23
+ $Y2=0
r23 9 10 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.295 $Y=0 $X2=0.455
+ $Y2=0
r24 8 18 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.69
+ $Y2=0
r25 8 10 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.455
+ $Y2=0
r26 4 10 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.455 $Y=0.085
+ $X2=0.455 $Y2=0
r27 4 6 17.8269 $w=3.18e-07 $l=4.95e-07 $layer=LI1_cond $X=0.455 $Y=0.085
+ $X2=0.455 $Y2=0.58
r28 1 6 182 $w=1.7e-07 $l=3.09112e-07 $layer=licon1_NDIFF $count=1 $X=0.315
+ $Y=0.335 $X2=0.46 $Y2=0.58
.ends

