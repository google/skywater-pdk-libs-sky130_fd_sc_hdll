* File: sky130_fd_sc_hdll__and4bb_2.spice
* Created: Thu Aug 27 18:59:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and4bb_2.pex.spice"
.subckt sky130_fd_sc_hdll__and4bb_2  VNB VPB A_N C D B_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B_N	B_N
* D	D
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_N_M1011_g N_A_27_47#_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.1302 PD=0.765421 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1011_d N_A_184_21#_M1012_g N_X_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.11785 AS=0.104 PD=1.18458 PS=0.97 NRD=9.228 NRS=8.304 M=1 R=4.33333
+ SA=75000.5 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_A_184_21#_M1013_g N_X_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.19175 AS=0.104 PD=1.89 PS=0.97 NRD=5.532 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 A_503_47# N_A_27_47#_M1000_g N_A_184_21#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.07245 AS=0.1092 PD=0.765 PS=1.36 NRD=33.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1004 A_602_47# N_A_545_280#_M1004_g A_503_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.07245 PD=0.755 PS=0.765 NRD=32.136 NRS=33.564 M=1 R=2.8
+ SA=75000.7 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1006 A_699_47# N_C_M1006_g A_602_47# VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.07035 PD=0.69 PS=0.755 NRD=22.848 NRS=32.136 M=1 R=2.8 SA=75001.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_D_M1005_g A_699_47# VNB NSHORT L=0.15 W=0.42 AD=0.1134
+ AS=0.0567 PD=0.96 PS=0.69 NRD=61.428 NRS=22.848 M=1 R=2.8 SA=75001.6
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1014 N_A_545_280#_M1014_d N_B_N_M1014_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.1134 PD=1.36 PS=0.96 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75002.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_N_M1002_g N_A_27_47#_M1002_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0874606 AS=0.1134 PD=0.795634 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90004.2 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1002_d N_A_184_21#_M1010_g N_X_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.208239 AS=0.145 PD=1.89437 PS=1.29 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90000.4 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1015 N_VPWR_M1015_d N_A_184_21#_M1015_g N_X_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.481761 AS=0.145 PD=2.45775 PS=1.29 NRD=16.7253 NRS=0.9653 M=1 R=5.55556
+ SA=90000.9 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1008 N_A_184_21#_M1008_d N_A_27_47#_M1008_g N_VPWR_M1015_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0672 AS=0.202339 PD=0.74 PS=1.03225 NRD=16.4101 NRS=18.7544 M=1
+ R=2.33333 SA=90002.1 SB=90002.3 A=0.0756 P=1.2 MULT=1
MM1009 N_VPWR_M1009_d N_A_545_280#_M1009_g N_A_184_21#_M1008_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.063 AS=0.0672 PD=0.72 PS=0.74 NRD=2.3443 NRS=2.3443 M=1
+ R=2.33333 SA=90002.6 SB=90001.8 A=0.0756 P=1.2 MULT=1
MM1003 N_A_184_21#_M1003_d N_C_M1003_g N_VPWR_M1009_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0609 AS=0.063 PD=0.71 PS=0.72 NRD=2.3443 NRS=7.0329 M=1 R=2.33333
+ SA=90003.1 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1001 N_VPWR_M1001_d N_D_M1001_g N_A_184_21#_M1003_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0966 AS=0.0609 PD=0.88 PS=0.71 NRD=82.0702 NRS=2.3443 M=1 R=2.33333
+ SA=90003.5 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1007 N_A_545_280#_M1007_d N_B_N_M1007_g N_VPWR_M1001_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.0966 PD=1.38 PS=0.88 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90004.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.7312 P=14.09
pX17_noxref noxref_16 X X PROBETYPE=1
pX18_noxref noxref_17 X X PROBETYPE=1
pX19_noxref noxref_18 X X PROBETYPE=1
*
.include "sky130_fd_sc_hdll__and4bb_2.pxi.spice"
*
.ends
*
*
