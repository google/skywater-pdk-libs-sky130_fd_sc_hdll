* File: sky130_fd_sc_hdll__nand2_8.pxi.spice
* Created: Wed Sep  2 08:37:04 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND2_8%B N_B_M1008_g N_B_c_120_n N_B_M1000_g
+ N_B_M1010_g N_B_c_121_n N_B_M1001_g N_B_M1011_g N_B_c_122_n N_B_M1003_g
+ N_B_M1015_g N_B_c_123_n N_B_M1009_g N_B_M1023_g N_B_c_124_n N_B_M1013_g
+ N_B_M1025_g N_B_c_125_n N_B_M1014_g N_B_M1027_g N_B_c_126_n N_B_M1020_g
+ N_B_c_127_n N_B_M1026_g N_B_M1028_g B B B B B B N_B_c_158_p N_B_c_119_n B B B
+ B B B PM_SKY130_FD_SC_HDLL__NAND2_8%B
x_PM_SKY130_FD_SC_HDLL__NAND2_8%A N_A_M1005_g N_A_c_284_n N_A_M1002_g
+ N_A_M1006_g N_A_c_285_n N_A_M1004_g N_A_M1012_g N_A_c_286_n N_A_M1007_g
+ N_A_M1016_g N_A_c_287_n N_A_M1017_g N_A_M1018_g N_A_c_288_n N_A_M1021_g
+ N_A_M1019_g N_A_c_289_n N_A_M1022_g N_A_M1029_g N_A_c_290_n N_A_M1024_g
+ N_A_c_291_n N_A_M1031_g N_A_M1030_g A A A A A N_A_c_334_p N_A_c_283_n A A A A
+ PM_SKY130_FD_SC_HDLL__NAND2_8%A
x_PM_SKY130_FD_SC_HDLL__NAND2_8%VPWR N_VPWR_M1000_d N_VPWR_M1001_d
+ N_VPWR_M1009_d N_VPWR_M1014_d N_VPWR_M1026_d N_VPWR_M1004_d N_VPWR_M1017_d
+ N_VPWR_M1022_d N_VPWR_M1031_d N_VPWR_c_408_n N_VPWR_c_409_n N_VPWR_c_410_n
+ N_VPWR_c_411_n N_VPWR_c_412_n N_VPWR_c_413_n N_VPWR_c_414_n N_VPWR_c_415_n
+ N_VPWR_c_416_n N_VPWR_c_417_n N_VPWR_c_418_n N_VPWR_c_419_n N_VPWR_c_420_n
+ N_VPWR_c_421_n N_VPWR_c_422_n N_VPWR_c_423_n N_VPWR_c_424_n N_VPWR_c_425_n
+ N_VPWR_c_426_n N_VPWR_c_427_n N_VPWR_c_428_n N_VPWR_c_429_n N_VPWR_c_430_n
+ VPWR N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_433_n N_VPWR_c_407_n
+ PM_SKY130_FD_SC_HDLL__NAND2_8%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND2_8%Y N_Y_M1005_s N_Y_M1012_s N_Y_M1018_s
+ N_Y_M1029_s N_Y_M1000_s N_Y_M1003_s N_Y_M1013_s N_Y_M1020_s N_Y_M1002_s
+ N_Y_M1007_s N_Y_M1021_s N_Y_M1024_s N_Y_c_547_n N_Y_c_567_n N_Y_c_548_n
+ N_Y_c_574_n N_Y_c_549_n N_Y_c_582_n N_Y_c_550_n N_Y_c_590_n N_Y_c_551_n
+ N_Y_c_613_n N_Y_c_543_n N_Y_c_596_n N_Y_c_544_n N_Y_c_552_n N_Y_c_545_n
+ N_Y_c_636_n N_Y_c_554_n N_Y_c_644_n N_Y_c_555_n N_Y_c_652_n N_Y_c_655_n
+ N_Y_c_546_n N_Y_c_557_n N_Y_c_558_n N_Y_c_559_n N_Y_c_560_n N_Y_c_561_n
+ N_Y_c_562_n Y PM_SKY130_FD_SC_HDLL__NAND2_8%Y
x_PM_SKY130_FD_SC_HDLL__NAND2_8%A_27_47# N_A_27_47#_M1008_s N_A_27_47#_M1010_s
+ N_A_27_47#_M1015_s N_A_27_47#_M1025_s N_A_27_47#_M1028_s N_A_27_47#_M1006_d
+ N_A_27_47#_M1016_d N_A_27_47#_M1019_d N_A_27_47#_M1030_d N_A_27_47#_c_751_n
+ N_A_27_47#_c_752_n N_A_27_47#_c_753_n N_A_27_47#_c_770_n N_A_27_47#_c_754_n
+ N_A_27_47#_c_778_n N_A_27_47#_c_755_n N_A_27_47#_c_786_n N_A_27_47#_c_756_n
+ N_A_27_47#_c_794_n N_A_27_47#_c_757_n N_A_27_47#_c_809_n N_A_27_47#_c_758_n
+ N_A_27_47#_c_759_n N_A_27_47#_c_760_n N_A_27_47#_c_761_n N_A_27_47#_c_762_n
+ PM_SKY130_FD_SC_HDLL__NAND2_8%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NAND2_8%VGND N_VGND_M1008_d N_VGND_M1011_d
+ N_VGND_M1023_d N_VGND_M1027_d N_VGND_c_886_n N_VGND_c_887_n N_VGND_c_888_n
+ N_VGND_c_889_n N_VGND_c_890_n N_VGND_c_891_n N_VGND_c_892_n N_VGND_c_893_n
+ VGND N_VGND_c_894_n N_VGND_c_895_n N_VGND_c_896_n N_VGND_c_897_n
+ N_VGND_c_898_n PM_SKY130_FD_SC_HDLL__NAND2_8%VGND
cc_1 VNB N_B_M1008_g 0.0244194f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_B_M1010_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_3 VNB N_B_M1011_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.56
cc_4 VNB N_B_M1015_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_5 VNB N_B_M1023_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=0.56
cc_6 VNB N_B_M1025_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=2.82 $Y2=0.56
cc_7 VNB N_B_M1027_g 0.0188821f $X=-0.19 $Y=-0.24 $X2=3.29 $Y2=0.56
cc_8 VNB N_B_M1028_g 0.0185931f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.56
cc_9 VNB N_B_c_119_n 0.195577f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.217
cc_10 VNB N_A_M1005_g 0.0177228f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_11 VNB N_A_M1006_g 0.0183212f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_12 VNB N_A_M1012_g 0.0183649f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.56
cc_13 VNB N_A_M1016_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_14 VNB N_A_M1018_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=0.56
cc_15 VNB N_A_M1019_g 0.0183665f $X=-0.19 $Y=-0.24 $X2=2.82 $Y2=0.56
cc_16 VNB N_A_M1029_g 0.0188028f $X=-0.19 $Y=-0.24 $X2=3.29 $Y2=0.56
cc_17 VNB N_A_M1030_g 0.0248318f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.56
cc_18 VNB N_A_c_283_n 0.197548f $X=-0.19 $Y=-0.24 $X2=3.55 $Y2=1.16
cc_19 VNB N_VPWR_c_407_n 0.345644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_543_n 0.00115644f $X=-0.19 $Y=-0.24 $X2=2.905 $Y2=1.105
cc_21 VNB N_Y_c_544_n 0.0144942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_Y_c_545_n 0.00328251f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.217
cc_23 VNB N_Y_c_546_n 0.00237253f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_751_n 0.0189842f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=0.56
cc_25 VNB N_A_27_47#_c_752_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_753_n 0.013432f $X=-0.19 $Y=-0.24 $X2=2.375 $Y2=1.41
cc_27 VNB N_A_27_47#_c_754_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=2.82 $Y2=0.56
cc_28 VNB N_A_27_47#_c_755_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=3.29 $Y2=0.56
cc_29 VNB N_A_27_47#_c_756_n 0.00289542f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.41
cc_30 VNB N_A_27_47#_c_757_n 0.00317367f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=1.025
cc_31 VNB N_A_27_47#_c_758_n 0.0100703f $X=-0.19 $Y=-0.24 $X2=2.905 $Y2=1.105
cc_32 VNB N_A_27_47#_c_759_n 0.0234324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_27_47#_c_760_n 0.00253093f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_27_47#_c_761_n 0.00253093f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_27_47#_c_762_n 0.00253093f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_886_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.56
cc_37 VNB N_VGND_c_887_n 0.0192031f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_38 VNB N_VGND_c_888_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_39 VNB N_VGND_c_889_n 0.0192031f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_890_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=1.025
cc_41 VNB N_VGND_c_891_n 0.00469188f $X=-0.19 $Y=-0.24 $X2=2.375 $Y2=1.41
cc_42 VNB N_VGND_c_892_n 0.0192031f $X=-0.19 $Y=-0.24 $X2=2.82 $Y2=1.025
cc_43 VNB N_VGND_c_893_n 0.00323954f $X=-0.19 $Y=-0.24 $X2=2.82 $Y2=0.56
cc_44 VNB N_VGND_c_894_n 0.108031f $X=-0.19 $Y=-0.24 $X2=3.315 $Y2=1.985
cc_45 VNB N_VGND_c_895_n 0.39537f $X=-0.19 $Y=-0.24 $X2=3.315 $Y2=1.985
cc_46 VNB N_VGND_c_896_n 0.0218366f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.985
cc_47 VNB N_VGND_c_897_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.56
cc_48 VNB N_VGND_c_898_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.105
cc_49 VPB N_B_c_120_n 0.0209831f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_50 VPB N_B_c_121_n 0.0160541f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_51 VPB N_B_c_122_n 0.0160541f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_52 VPB N_B_c_123_n 0.0160541f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_53 VPB N_B_c_124_n 0.0160541f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_54 VPB N_B_c_125_n 0.0160541f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_55 VPB N_B_c_126_n 0.0160532f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.41
cc_56 VPB N_B_c_127_n 0.0161676f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_57 VPB N_B_c_119_n 0.0542456f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.217
cc_58 VPB N_A_c_284_n 0.0156532f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_59 VPB N_A_c_285_n 0.016036f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_60 VPB N_A_c_286_n 0.0160344f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_61 VPB N_A_c_287_n 0.0160541f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_62 VPB N_A_c_288_n 0.0160541f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_63 VPB N_A_c_289_n 0.0160343f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_64 VPB N_A_c_290_n 0.0160359f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.41
cc_65 VPB N_A_c_291_n 0.020749f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_66 VPB N_A_c_283_n 0.0528029f $X=-0.19 $Y=1.305 $X2=3.55 $Y2=1.16
cc_67 VPB N_VPWR_c_408_n 0.00994749f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_68 VPB N_VPWR_c_409_n 0.043135f $X=-0.19 $Y=1.305 $X2=2.35 $Y2=0.56
cc_69 VPB N_VPWR_c_410_n 0.0206409f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.985
cc_70 VPB N_VPWR_c_411_n 0.00469739f $X=-0.19 $Y=1.305 $X2=2.82 $Y2=0.56
cc_71 VPB N_VPWR_c_412_n 0.0206409f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_72 VPB N_VPWR_c_413_n 0.00469739f $X=-0.19 $Y=1.305 $X2=3.29 $Y2=0.56
cc_73 VPB N_VPWR_c_414_n 0.00469739f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.985
cc_74 VPB N_VPWR_c_415_n 0.00469739f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.985
cc_75 VPB N_VPWR_c_416_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_417_n 0.00469739f $X=-0.19 $Y=1.305 $X2=1.985 $Y2=1.105
cc_77 VPB N_VPWR_c_418_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_419_n 0.0157021f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_420_n 0.0452122f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_421_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0.725 $Y2=1.16
cc_81 VPB N_VPWR_c_422_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.217
cc_82 VPB N_VPWR_c_423_n 0.0206409f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=1.217
cc_83 VPB N_VPWR_c_424_n 0.00324069f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.217
cc_84 VPB N_VPWR_c_425_n 0.0206409f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.217
cc_85 VPB N_VPWR_c_426_n 0.00324069f $X=-0.19 $Y=1.305 $X2=2.35 $Y2=1.217
cc_86 VPB N_VPWR_c_427_n 0.0206409f $X=-0.19 $Y=1.305 $X2=2.82 $Y2=1.217
cc_87 VPB N_VPWR_c_428_n 0.00324069f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.217
cc_88 VPB N_VPWR_c_429_n 0.0206409f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.217
cc_89 VPB N_VPWR_c_430_n 0.00324069f $X=-0.19 $Y=1.305 $X2=3.55 $Y2=1.217
cc_90 VPB N_VPWR_c_431_n 0.0212773f $X=-0.19 $Y=1.305 $X2=2.535 $Y2=1.185
cc_91 VPB N_VPWR_c_432_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_433_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_407_n 0.0482998f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_Y_c_547_n 0.00177608f $X=-0.19 $Y=1.305 $X2=2.82 $Y2=0.56
cc_95 VPB N_Y_c_548_n 0.00174278f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.985
cc_96 VPB N_Y_c_549_n 0.00174278f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.41
cc_97 VPB N_Y_c_550_n 0.00174278f $X=-0.19 $Y=1.305 $X2=3.81 $Y2=1.025
cc_98 VPB N_Y_c_551_n 0.00245746f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=1.105
cc_99 VPB N_Y_c_552_n 0.00180268f $X=-0.19 $Y=1.305 $X2=0.725 $Y2=1.16
cc_100 VPB N_Y_c_545_n 0.00395107f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.217
cc_101 VPB N_Y_c_554_n 0.00180268f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.217
cc_102 VPB N_Y_c_555_n 0.00180268f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.217
cc_103 VPB N_Y_c_546_n 0.00151358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_Y_c_557_n 0.00177608f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.185
cc_105 VPB N_Y_c_558_n 0.00177608f $X=-0.19 $Y=1.305 $X2=1.61 $Y2=1.185
cc_106 VPB N_Y_c_559_n 0.00177608f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=1.19
cc_107 VPB N_Y_c_560_n 0.00183791f $X=-0.19 $Y=1.305 $X2=2.53 $Y2=1.185
cc_108 VPB N_Y_c_561_n 0.00183791f $X=-0.19 $Y=1.305 $X2=2.535 $Y2=1.19
cc_109 VPB N_Y_c_562_n 4.86222e-19 $X=-0.19 $Y=1.305 $X2=2.995 $Y2=1.185
cc_110 N_B_M1028_g N_A_M1005_g 0.0159017f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_111 N_B_c_127_n N_A_c_284_n 0.0226885f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_112 N_B_c_119_n N_A_c_283_n 0.0159017f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_113 N_B_c_120_n N_VPWR_c_409_n 0.00777002f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_114 N_B_c_120_n N_VPWR_c_410_n 0.00597712f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_115 N_B_c_121_n N_VPWR_c_410_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_116 N_B_c_121_n N_VPWR_c_411_n 0.0052072f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_117 N_B_c_122_n N_VPWR_c_411_n 0.004751f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_118 N_B_c_122_n N_VPWR_c_412_n 0.00597712f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_119 N_B_c_123_n N_VPWR_c_412_n 0.00673617f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_120 N_B_c_123_n N_VPWR_c_413_n 0.0052072f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_121 N_B_c_124_n N_VPWR_c_413_n 0.004751f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_122 N_B_c_125_n N_VPWR_c_414_n 0.0052072f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_123 N_B_c_126_n N_VPWR_c_414_n 0.004751f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_124 N_B_c_127_n N_VPWR_c_415_n 0.0052072f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_125 N_B_c_124_n N_VPWR_c_421_n 0.00597712f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_126 N_B_c_125_n N_VPWR_c_421_n 0.00673617f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_127 N_B_c_126_n N_VPWR_c_423_n 0.00597712f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_128 N_B_c_127_n N_VPWR_c_423_n 0.00673617f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_129 N_B_c_120_n N_VPWR_c_407_n 0.010906f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_130 N_B_c_121_n N_VPWR_c_407_n 0.0118438f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_131 N_B_c_122_n N_VPWR_c_407_n 0.00999457f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_132 N_B_c_123_n N_VPWR_c_407_n 0.0118438f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_133 N_B_c_124_n N_VPWR_c_407_n 0.00999457f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_134 N_B_c_125_n N_VPWR_c_407_n 0.0118438f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_135 N_B_c_126_n N_VPWR_c_407_n 0.00999457f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_136 N_B_c_127_n N_VPWR_c_407_n 0.011869f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_137 N_B_c_120_n N_Y_c_547_n 0.00525563f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_138 N_B_c_121_n N_Y_c_547_n 8.83441e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_139 N_B_c_158_p N_Y_c_547_n 0.0307772f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_140 N_B_c_119_n N_Y_c_547_n 0.00730145f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_141 N_B_c_120_n N_Y_c_567_n 0.0121679f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_142 N_B_c_121_n N_Y_c_567_n 0.0106251f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_143 N_B_c_122_n N_Y_c_567_n 6.24674e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_144 N_B_c_121_n N_Y_c_548_n 0.0147591f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_145 N_B_c_122_n N_Y_c_548_n 0.0108841f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_146 N_B_c_158_p N_Y_c_548_n 0.0402453f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_147 N_B_c_119_n N_Y_c_548_n 0.00706727f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_148 N_B_c_121_n N_Y_c_574_n 6.48386e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_149 N_B_c_122_n N_Y_c_574_n 0.0130707f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_150 N_B_c_123_n N_Y_c_574_n 0.0106251f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_151 N_B_c_124_n N_Y_c_574_n 6.24674e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_152 N_B_c_123_n N_Y_c_549_n 0.0147591f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_153 N_B_c_124_n N_Y_c_549_n 0.0108841f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_154 N_B_c_158_p N_Y_c_549_n 0.0402453f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_155 N_B_c_119_n N_Y_c_549_n 0.00706727f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_156 N_B_c_123_n N_Y_c_582_n 6.48386e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_157 N_B_c_124_n N_Y_c_582_n 0.0130707f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_158 N_B_c_125_n N_Y_c_582_n 0.0106251f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_159 N_B_c_126_n N_Y_c_582_n 6.24674e-19 $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_160 N_B_c_125_n N_Y_c_550_n 0.0147591f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_161 N_B_c_126_n N_Y_c_550_n 0.0108841f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_162 N_B_c_158_p N_Y_c_550_n 0.0402453f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_163 N_B_c_119_n N_Y_c_550_n 0.00706727f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_164 N_B_c_125_n N_Y_c_590_n 6.48386e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_165 N_B_c_126_n N_Y_c_590_n 0.0130707f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_166 N_B_c_127_n N_Y_c_590_n 0.0106251f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_167 N_B_c_127_n N_Y_c_551_n 0.0167312f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_168 N_B_c_119_n N_Y_c_551_n 3.53895e-19 $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_169 N_B_M1028_g N_Y_c_543_n 8.77318e-19 $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_170 N_B_c_127_n N_Y_c_596_n 6.48386e-19 $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_171 N_B_c_127_n N_Y_c_545_n 0.00144378f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_172 N_B_c_158_p N_Y_c_545_n 0.0117073f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_173 N_B_c_119_n N_Y_c_545_n 0.00528509f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_174 N_B_c_122_n N_Y_c_557_n 0.00254988f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_175 N_B_c_123_n N_Y_c_557_n 8.83441e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_176 N_B_c_158_p N_Y_c_557_n 0.0307772f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_177 N_B_c_119_n N_Y_c_557_n 0.00730145f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_178 N_B_c_124_n N_Y_c_558_n 0.00254988f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_179 N_B_c_125_n N_Y_c_558_n 8.83441e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_180 N_B_c_158_p N_Y_c_558_n 0.0307772f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_181 N_B_c_119_n N_Y_c_558_n 0.00730145f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_182 N_B_c_126_n N_Y_c_559_n 0.00254988f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_183 N_B_c_127_n N_Y_c_559_n 8.83441e-19 $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_184 N_B_c_158_p N_Y_c_559_n 0.0307772f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_185 N_B_c_119_n N_Y_c_559_n 0.00705894f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_186 N_B_M1008_g N_A_27_47#_c_751_n 0.00698303f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_187 N_B_M1010_g N_A_27_47#_c_751_n 5.49487e-19 $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_188 N_B_M1008_g N_A_27_47#_c_752_n 0.0113635f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_189 N_B_M1010_g N_A_27_47#_c_752_n 0.00879805f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_190 N_B_c_158_p N_A_27_47#_c_752_n 0.0340131f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_191 N_B_c_119_n N_A_27_47#_c_752_n 0.0031956f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_192 N_B_M1008_g N_A_27_47#_c_753_n 0.00231729f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_193 N_B_M1008_g N_A_27_47#_c_770_n 5.27166e-19 $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_194 N_B_M1010_g N_A_27_47#_c_770_n 0.0066221f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_195 N_B_M1011_g N_A_27_47#_c_770_n 0.00698303f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_196 N_B_M1015_g N_A_27_47#_c_770_n 5.48764e-19 $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_197 N_B_M1011_g N_A_27_47#_c_754_n 0.00879805f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_198 N_B_M1015_g N_A_27_47#_c_754_n 0.00879805f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_199 N_B_c_158_p N_A_27_47#_c_754_n 0.0398571f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_200 N_B_c_119_n N_A_27_47#_c_754_n 0.0031956f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_201 N_B_M1011_g N_A_27_47#_c_778_n 5.27166e-19 $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_202 N_B_M1015_g N_A_27_47#_c_778_n 0.0066221f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_203 N_B_M1023_g N_A_27_47#_c_778_n 0.00698303f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_204 N_B_M1025_g N_A_27_47#_c_778_n 5.48764e-19 $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_205 N_B_M1023_g N_A_27_47#_c_755_n 0.00879805f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_206 N_B_M1025_g N_A_27_47#_c_755_n 0.00879805f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_207 N_B_c_158_p N_A_27_47#_c_755_n 0.0398571f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_208 N_B_c_119_n N_A_27_47#_c_755_n 0.0031956f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_209 N_B_M1023_g N_A_27_47#_c_786_n 5.27166e-19 $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_210 N_B_M1025_g N_A_27_47#_c_786_n 0.0066221f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_211 N_B_M1027_g N_A_27_47#_c_786_n 0.00705334f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_212 N_B_M1028_g N_A_27_47#_c_786_n 5.37075e-19 $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_213 N_B_M1027_g N_A_27_47#_c_756_n 0.00905701f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_214 N_B_M1028_g N_A_27_47#_c_756_n 0.00717326f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_215 N_B_c_158_p N_A_27_47#_c_756_n 0.0337791f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_216 N_B_c_119_n N_A_27_47#_c_756_n 0.00433688f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_217 N_B_M1028_g N_A_27_47#_c_794_n 0.00388968f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_218 N_B_M1027_g N_A_27_47#_c_757_n 5.13362e-19 $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_219 N_B_M1028_g N_A_27_47#_c_757_n 0.00845447f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_220 N_B_M1010_g N_A_27_47#_c_760_n 0.00113905f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_221 N_B_M1011_g N_A_27_47#_c_760_n 0.00113905f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_222 N_B_c_158_p N_A_27_47#_c_760_n 0.0307978f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_223 N_B_c_119_n N_A_27_47#_c_760_n 0.00332f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_224 N_B_M1015_g N_A_27_47#_c_761_n 0.00113905f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_225 N_B_M1023_g N_A_27_47#_c_761_n 0.00113905f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_226 N_B_c_158_p N_A_27_47#_c_761_n 0.0307978f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_227 N_B_c_119_n N_A_27_47#_c_761_n 0.00332f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_228 N_B_M1025_g N_A_27_47#_c_762_n 0.00113905f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_229 N_B_M1027_g N_A_27_47#_c_762_n 0.00113905f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_230 N_B_c_158_p N_A_27_47#_c_762_n 0.0307978f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_231 N_B_c_119_n N_A_27_47#_c_762_n 0.00332f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_232 N_B_M1008_g N_VGND_c_886_n 0.00382421f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_233 N_B_M1010_g N_VGND_c_886_n 0.00276126f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_234 N_B_M1010_g N_VGND_c_887_n 0.00424416f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_235 N_B_M1011_g N_VGND_c_887_n 0.00424416f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_236 N_B_M1011_g N_VGND_c_888_n 0.00382421f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_237 N_B_M1015_g N_VGND_c_888_n 0.00276126f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_238 N_B_M1015_g N_VGND_c_889_n 0.00424416f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_239 N_B_M1023_g N_VGND_c_889_n 0.00424416f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_240 N_B_M1023_g N_VGND_c_890_n 0.00382421f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_241 N_B_M1025_g N_VGND_c_890_n 0.00276126f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_242 N_B_M1027_g N_VGND_c_891_n 0.00388664f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_243 N_B_M1028_g N_VGND_c_891_n 0.00367616f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_244 N_B_M1025_g N_VGND_c_892_n 0.00424416f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_245 N_B_M1027_g N_VGND_c_892_n 0.00424416f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_246 N_B_M1028_g N_VGND_c_894_n 0.00395719f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_247 N_B_M1008_g N_VGND_c_895_n 0.00694001f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_248 N_B_M1010_g N_VGND_c_895_n 0.00599001f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_249 N_B_M1011_g N_VGND_c_895_n 0.00611278f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_250 N_B_M1015_g N_VGND_c_895_n 0.00599001f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_251 N_B_M1023_g N_VGND_c_895_n 0.00611278f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_252 N_B_M1025_g N_VGND_c_895_n 0.00599001f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_253 N_B_M1027_g N_VGND_c_895_n 0.00622812f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_254 N_B_M1028_g N_VGND_c_895_n 0.00585096f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_255 N_B_M1008_g N_VGND_c_896_n 0.00424416f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_256 N_A_c_284_n N_VPWR_c_415_n 0.004751f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_257 N_A_c_285_n N_VPWR_c_416_n 0.0052072f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_258 N_A_c_286_n N_VPWR_c_416_n 0.004751f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A_c_287_n N_VPWR_c_417_n 0.0052072f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A_c_288_n N_VPWR_c_417_n 0.004751f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A_c_289_n N_VPWR_c_418_n 0.0052072f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A_c_290_n N_VPWR_c_418_n 0.004751f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A_c_291_n N_VPWR_c_420_n 0.0281539f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A_c_284_n N_VPWR_c_425_n 0.00597712f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A_c_285_n N_VPWR_c_425_n 0.00673617f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A_c_286_n N_VPWR_c_427_n 0.00597712f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_267 N_A_c_287_n N_VPWR_c_427_n 0.00673617f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A_c_288_n N_VPWR_c_429_n 0.00597712f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A_c_289_n N_VPWR_c_429_n 0.00673617f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_270 N_A_c_290_n N_VPWR_c_431_n 0.00597712f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_271 N_A_c_291_n N_VPWR_c_431_n 0.00673617f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_272 N_A_c_284_n N_VPWR_c_407_n 0.0100198f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_273 N_A_c_285_n N_VPWR_c_407_n 0.0118438f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_274 N_A_c_286_n N_VPWR_c_407_n 0.00999457f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_275 N_A_c_287_n N_VPWR_c_407_n 0.0118438f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_276 N_A_c_288_n N_VPWR_c_407_n 0.00999457f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_277 N_A_c_289_n N_VPWR_c_407_n 0.0118438f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_278 N_A_c_290_n N_VPWR_c_407_n 0.00999457f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_279 N_A_c_291_n N_VPWR_c_407_n 0.0130834f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_280 N_A_c_284_n N_Y_c_590_n 6.24674e-19 $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_281 N_A_M1005_g N_Y_c_613_n 0.00328621f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_282 N_A_M1005_g N_Y_c_543_n 0.00343295f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_283 N_A_M1006_g N_Y_c_543_n 0.00321836f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_284 N_A_c_283_n N_Y_c_543_n 0.00738569f $X=7.545 $Y=1.217 $X2=0 $Y2=0
cc_285 N_A_c_284_n N_Y_c_596_n 0.0130707f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_286 N_A_c_285_n N_Y_c_596_n 0.0106251f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_287 N_A_c_286_n N_Y_c_596_n 6.24674e-19 $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_288 N_A_M1006_g N_Y_c_544_n 0.0125002f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_289 N_A_M1012_g N_Y_c_544_n 0.0111698f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_290 N_A_M1016_g N_Y_c_544_n 0.0111698f $X=5.64 $Y=0.56 $X2=0 $Y2=0
cc_291 N_A_M1018_g N_Y_c_544_n 0.0111698f $X=6.11 $Y=0.56 $X2=0 $Y2=0
cc_292 N_A_M1019_g N_Y_c_544_n 0.0111698f $X=6.58 $Y=0.56 $X2=0 $Y2=0
cc_293 N_A_M1029_g N_Y_c_544_n 0.0125717f $X=7.05 $Y=0.56 $X2=0 $Y2=0
cc_294 N_A_c_334_p N_Y_c_544_n 0.166476f $X=6.84 $Y=1.16 $X2=0 $Y2=0
cc_295 N_A_c_283_n N_Y_c_544_n 0.0164066f $X=7.545 $Y=1.217 $X2=0 $Y2=0
cc_296 N_A_c_285_n N_Y_c_552_n 0.0158169f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_297 N_A_c_286_n N_Y_c_552_n 0.0109733f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_298 N_A_c_334_p N_Y_c_552_n 0.0312905f $X=6.84 $Y=1.16 $X2=0 $Y2=0
cc_299 N_A_c_283_n N_Y_c_552_n 0.00713968f $X=7.545 $Y=1.217 $X2=0 $Y2=0
cc_300 N_A_c_284_n N_Y_c_545_n 0.013432f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_301 N_A_c_285_n N_Y_c_545_n 0.00273701f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_302 N_A_c_334_p N_Y_c_545_n 0.016449f $X=6.84 $Y=1.16 $X2=0 $Y2=0
cc_303 N_A_c_283_n N_Y_c_545_n 0.0325622f $X=7.545 $Y=1.217 $X2=0 $Y2=0
cc_304 N_A_c_285_n N_Y_c_636_n 6.48386e-19 $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_305 N_A_c_286_n N_Y_c_636_n 0.0130707f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_306 N_A_c_287_n N_Y_c_636_n 0.0106251f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_307 N_A_c_288_n N_Y_c_636_n 6.24674e-19 $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_308 N_A_c_287_n N_Y_c_554_n 0.0148893f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_309 N_A_c_288_n N_Y_c_554_n 0.0109733f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_310 N_A_c_334_p N_Y_c_554_n 0.0366623f $X=6.84 $Y=1.16 $X2=0 $Y2=0
cc_311 N_A_c_283_n N_Y_c_554_n 0.00713968f $X=7.545 $Y=1.217 $X2=0 $Y2=0
cc_312 N_A_c_287_n N_Y_c_644_n 6.48386e-19 $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_313 N_A_c_288_n N_Y_c_644_n 0.0130707f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_314 N_A_c_289_n N_Y_c_644_n 0.0106251f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_315 N_A_c_290_n N_Y_c_644_n 6.24674e-19 $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_316 N_A_c_289_n N_Y_c_555_n 0.0148893f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_317 N_A_c_290_n N_Y_c_555_n 0.0119562f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_318 N_A_c_334_p N_Y_c_555_n 0.0309726f $X=6.84 $Y=1.16 $X2=0 $Y2=0
cc_319 N_A_c_283_n N_Y_c_555_n 0.00713968f $X=7.545 $Y=1.217 $X2=0 $Y2=0
cc_320 N_A_c_289_n N_Y_c_652_n 6.48386e-19 $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_321 N_A_c_290_n N_Y_c_652_n 0.0130707f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_322 N_A_c_291_n N_Y_c_652_n 0.0104317f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_323 N_A_M1030_g N_Y_c_655_n 2.15189e-19 $X=7.57 $Y=0.56 $X2=0 $Y2=0
cc_324 N_A_M1029_g N_Y_c_546_n 0.00301547f $X=7.05 $Y=0.56 $X2=0 $Y2=0
cc_325 N_A_c_290_n N_Y_c_546_n 0.00139555f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_326 N_A_c_291_n N_Y_c_546_n 0.00272791f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_327 N_A_M1030_g N_Y_c_546_n 0.00334167f $X=7.57 $Y=0.56 $X2=0 $Y2=0
cc_328 N_A_c_334_p N_Y_c_546_n 0.0125942f $X=6.84 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A_c_283_n N_Y_c_546_n 0.0420707f $X=7.545 $Y=1.217 $X2=0 $Y2=0
cc_330 N_A_c_286_n N_Y_c_560_n 0.00261058f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_331 N_A_c_287_n N_Y_c_560_n 9.00783e-19 $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_332 N_A_c_334_p N_Y_c_560_n 0.028094f $X=6.84 $Y=1.16 $X2=0 $Y2=0
cc_333 N_A_c_283_n N_Y_c_560_n 0.00739893f $X=7.545 $Y=1.217 $X2=0 $Y2=0
cc_334 N_A_c_288_n N_Y_c_561_n 0.00261058f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_335 N_A_c_289_n N_Y_c_561_n 9.00783e-19 $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_336 N_A_c_334_p N_Y_c_561_n 0.028094f $X=6.84 $Y=1.16 $X2=0 $Y2=0
cc_337 N_A_c_283_n N_Y_c_561_n 0.00739893f $X=7.545 $Y=1.217 $X2=0 $Y2=0
cc_338 N_A_c_290_n N_Y_c_562_n 0.00332859f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_339 N_A_c_291_n N_Y_c_562_n 0.00384224f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_340 N_A_c_283_n N_Y_c_562_n 0.00197478f $X=7.545 $Y=1.217 $X2=0 $Y2=0
cc_341 N_A_M1005_g N_A_27_47#_c_809_n 0.0111995f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_342 N_A_M1006_g N_A_27_47#_c_809_n 0.00958923f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_343 N_A_M1012_g N_A_27_47#_c_809_n 0.00958923f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_344 N_A_M1016_g N_A_27_47#_c_809_n 0.00958923f $X=5.64 $Y=0.56 $X2=0 $Y2=0
cc_345 N_A_M1018_g N_A_27_47#_c_809_n 0.00958923f $X=6.11 $Y=0.56 $X2=0 $Y2=0
cc_346 N_A_M1019_g N_A_27_47#_c_809_n 0.00958923f $X=6.58 $Y=0.56 $X2=0 $Y2=0
cc_347 N_A_M1029_g N_A_27_47#_c_809_n 0.00994068f $X=7.05 $Y=0.56 $X2=0 $Y2=0
cc_348 N_A_M1030_g N_A_27_47#_c_809_n 0.0197404f $X=7.57 $Y=0.56 $X2=0 $Y2=0
cc_349 N_A_c_283_n N_A_27_47#_c_809_n 0.00108741f $X=7.545 $Y=1.217 $X2=0 $Y2=0
cc_350 N_A_M1030_g N_A_27_47#_c_759_n 0.00817004f $X=7.57 $Y=0.56 $X2=0 $Y2=0
cc_351 N_A_M1005_g N_VGND_c_894_n 0.00357877f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_352 N_A_M1006_g N_VGND_c_894_n 0.00357877f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_353 N_A_M1012_g N_VGND_c_894_n 0.00357877f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_354 N_A_M1016_g N_VGND_c_894_n 0.00357877f $X=5.64 $Y=0.56 $X2=0 $Y2=0
cc_355 N_A_M1018_g N_VGND_c_894_n 0.00357877f $X=6.11 $Y=0.56 $X2=0 $Y2=0
cc_356 N_A_M1019_g N_VGND_c_894_n 0.00357877f $X=6.58 $Y=0.56 $X2=0 $Y2=0
cc_357 N_A_M1029_g N_VGND_c_894_n 0.00357877f $X=7.05 $Y=0.56 $X2=0 $Y2=0
cc_358 N_A_M1030_g N_VGND_c_894_n 0.00357877f $X=7.57 $Y=0.56 $X2=0 $Y2=0
cc_359 N_A_M1005_g N_VGND_c_895_n 0.00538422f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_360 N_A_M1006_g N_VGND_c_895_n 0.00548399f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_361 N_A_M1012_g N_VGND_c_895_n 0.00548399f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_362 N_A_M1016_g N_VGND_c_895_n 0.00548399f $X=5.64 $Y=0.56 $X2=0 $Y2=0
cc_363 N_A_M1018_g N_VGND_c_895_n 0.00548399f $X=6.11 $Y=0.56 $X2=0 $Y2=0
cc_364 N_A_M1019_g N_VGND_c_895_n 0.00548399f $X=6.58 $Y=0.56 $X2=0 $Y2=0
cc_365 N_A_M1029_g N_VGND_c_895_n 0.00560377f $X=7.05 $Y=0.56 $X2=0 $Y2=0
cc_366 N_A_M1030_g N_VGND_c_895_n 0.00667694f $X=7.57 $Y=0.56 $X2=0 $Y2=0
cc_367 N_VPWR_c_407_n N_Y_M1000_s 0.00231261f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_368 N_VPWR_c_407_n N_Y_M1003_s 0.00231261f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_369 N_VPWR_c_407_n N_Y_M1013_s 0.00231261f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_370 N_VPWR_c_407_n N_Y_M1020_s 0.00231261f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_371 N_VPWR_c_407_n N_Y_M1002_s 0.00231261f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_372 N_VPWR_c_407_n N_Y_M1007_s 0.00231261f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_373 N_VPWR_c_407_n N_Y_M1021_s 0.00231261f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_374 N_VPWR_c_407_n N_Y_M1024_s 0.00231261f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_375 N_VPWR_c_409_n N_Y_c_547_n 0.0137498f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_376 N_VPWR_c_409_n N_Y_c_567_n 0.0615045f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_377 N_VPWR_c_410_n N_Y_c_567_n 0.0223557f $X=1.115 $Y=2.72 $X2=0 $Y2=0
cc_378 N_VPWR_c_411_n N_Y_c_567_n 0.0385613f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_379 N_VPWR_c_407_n N_Y_c_567_n 0.0140101f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_380 N_VPWR_M1001_d N_Y_c_548_n 0.00179485f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_381 N_VPWR_c_411_n N_Y_c_548_n 0.0138194f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_382 N_VPWR_c_411_n N_Y_c_574_n 0.0470327f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_383 N_VPWR_c_412_n N_Y_c_574_n 0.0223557f $X=2.055 $Y=2.72 $X2=0 $Y2=0
cc_384 N_VPWR_c_413_n N_Y_c_574_n 0.0385613f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_385 N_VPWR_c_407_n N_Y_c_574_n 0.0140101f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_386 N_VPWR_M1009_d N_Y_c_549_n 0.00179485f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_387 N_VPWR_c_413_n N_Y_c_549_n 0.0138194f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_388 N_VPWR_c_413_n N_Y_c_582_n 0.0470327f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_389 N_VPWR_c_414_n N_Y_c_582_n 0.0385613f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_390 N_VPWR_c_421_n N_Y_c_582_n 0.0223557f $X=2.995 $Y=2.72 $X2=0 $Y2=0
cc_391 N_VPWR_c_407_n N_Y_c_582_n 0.0140101f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_392 N_VPWR_M1014_d N_Y_c_550_n 0.00179485f $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_393 N_VPWR_c_414_n N_Y_c_550_n 0.0138194f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_394 N_VPWR_c_414_n N_Y_c_590_n 0.0470327f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_395 N_VPWR_c_415_n N_Y_c_590_n 0.0385613f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_396 N_VPWR_c_423_n N_Y_c_590_n 0.0223557f $X=3.935 $Y=2.72 $X2=0 $Y2=0
cc_397 N_VPWR_c_407_n N_Y_c_590_n 0.0140101f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_398 N_VPWR_M1026_d N_Y_c_551_n 0.00110041f $X=3.875 $Y=1.485 $X2=0 $Y2=0
cc_399 N_VPWR_c_415_n N_Y_c_551_n 0.00851749f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_400 N_VPWR_c_415_n N_Y_c_596_n 0.0470327f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_401 N_VPWR_c_416_n N_Y_c_596_n 0.0385613f $X=4.96 $Y=2 $X2=0 $Y2=0
cc_402 N_VPWR_c_425_n N_Y_c_596_n 0.0223557f $X=4.875 $Y=2.72 $X2=0 $Y2=0
cc_403 N_VPWR_c_407_n N_Y_c_596_n 0.0140101f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_404 N_VPWR_M1004_d N_Y_c_552_n 0.00179485f $X=4.815 $Y=1.485 $X2=0 $Y2=0
cc_405 N_VPWR_c_416_n N_Y_c_552_n 0.0138194f $X=4.96 $Y=2 $X2=0 $Y2=0
cc_406 N_VPWR_M1026_d N_Y_c_545_n 7.05179e-19 $X=3.875 $Y=1.485 $X2=0 $Y2=0
cc_407 N_VPWR_c_415_n N_Y_c_545_n 0.00571024f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_408 N_VPWR_c_416_n N_Y_c_636_n 0.0470327f $X=4.96 $Y=2 $X2=0 $Y2=0
cc_409 N_VPWR_c_417_n N_Y_c_636_n 0.0385613f $X=5.9 $Y=2 $X2=0 $Y2=0
cc_410 N_VPWR_c_427_n N_Y_c_636_n 0.0223557f $X=5.815 $Y=2.72 $X2=0 $Y2=0
cc_411 N_VPWR_c_407_n N_Y_c_636_n 0.0140101f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_412 N_VPWR_M1017_d N_Y_c_554_n 0.00179485f $X=5.755 $Y=1.485 $X2=0 $Y2=0
cc_413 N_VPWR_c_417_n N_Y_c_554_n 0.0138194f $X=5.9 $Y=2 $X2=0 $Y2=0
cc_414 N_VPWR_c_417_n N_Y_c_644_n 0.0470327f $X=5.9 $Y=2 $X2=0 $Y2=0
cc_415 N_VPWR_c_418_n N_Y_c_644_n 0.0385613f $X=6.84 $Y=2 $X2=0 $Y2=0
cc_416 N_VPWR_c_429_n N_Y_c_644_n 0.0223557f $X=6.755 $Y=2.72 $X2=0 $Y2=0
cc_417 N_VPWR_c_407_n N_Y_c_644_n 0.0140101f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_418 N_VPWR_M1022_d N_Y_c_555_n 0.00179485f $X=6.695 $Y=1.485 $X2=0 $Y2=0
cc_419 N_VPWR_c_418_n N_Y_c_555_n 0.0138194f $X=6.84 $Y=2 $X2=0 $Y2=0
cc_420 N_VPWR_c_418_n N_Y_c_652_n 0.0470327f $X=6.84 $Y=2 $X2=0 $Y2=0
cc_421 N_VPWR_c_420_n N_Y_c_652_n 0.0484009f $X=7.88 $Y=1.66 $X2=0 $Y2=0
cc_422 N_VPWR_c_431_n N_Y_c_652_n 0.0223557f $X=7.715 $Y=2.72 $X2=0 $Y2=0
cc_423 N_VPWR_c_407_n N_Y_c_652_n 0.0140101f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_424 N_VPWR_c_420_n N_Y_c_562_n 0.0107883f $X=7.88 $Y=1.66 $X2=0 $Y2=0
cc_425 N_VPWR_c_409_n N_A_27_47#_c_753_n 0.00949095f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_426 N_VPWR_c_420_n N_A_27_47#_c_759_n 0.0132088f $X=7.88 $Y=1.66 $X2=0 $Y2=0
cc_427 N_Y_c_544_n N_A_27_47#_M1006_d 0.00214463f $X=7.225 $Y=0.78 $X2=0 $Y2=0
cc_428 N_Y_c_544_n N_A_27_47#_M1016_d 0.00214463f $X=7.225 $Y=0.78 $X2=0 $Y2=0
cc_429 N_Y_c_544_n N_A_27_47#_M1019_d 0.00214463f $X=7.225 $Y=0.78 $X2=0 $Y2=0
cc_430 N_Y_c_551_n N_A_27_47#_c_756_n 0.00236731f $X=4.04 $Y=1.565 $X2=0 $Y2=0
cc_431 N_Y_c_551_n N_A_27_47#_c_757_n 0.0080681f $X=4.04 $Y=1.565 $X2=0 $Y2=0
cc_432 N_Y_c_613_n N_A_27_47#_c_757_n 0.00808483f $X=4.422 $Y=0.905 $X2=0 $Y2=0
cc_433 N_Y_c_545_n N_A_27_47#_c_757_n 0.00600544f $X=4.655 $Y=1.565 $X2=0 $Y2=0
cc_434 N_Y_M1005_s N_A_27_47#_c_809_n 0.00401256f $X=4.305 $Y=0.235 $X2=0 $Y2=0
cc_435 N_Y_M1012_s N_A_27_47#_c_809_n 0.00401739f $X=5.245 $Y=0.235 $X2=0 $Y2=0
cc_436 N_Y_M1018_s N_A_27_47#_c_809_n 0.00401739f $X=6.185 $Y=0.235 $X2=0 $Y2=0
cc_437 N_Y_M1029_s N_A_27_47#_c_809_n 0.00508688f $X=7.125 $Y=0.235 $X2=0 $Y2=0
cc_438 N_Y_c_613_n N_A_27_47#_c_809_n 0.0184116f $X=4.422 $Y=0.905 $X2=0 $Y2=0
cc_439 N_Y_c_544_n N_A_27_47#_c_809_n 0.138906f $X=7.225 $Y=0.78 $X2=0 $Y2=0
cc_440 N_Y_c_545_n N_A_27_47#_c_809_n 0.00423797f $X=4.655 $Y=1.565 $X2=0 $Y2=0
cc_441 N_Y_c_655_n N_A_27_47#_c_809_n 0.0167869f $X=7.35 $Y=0.905 $X2=0 $Y2=0
cc_442 N_Y_c_655_n N_A_27_47#_c_759_n 0.00141307f $X=7.35 $Y=0.905 $X2=0 $Y2=0
cc_443 N_Y_M1005_s N_VGND_c_895_n 0.00256987f $X=4.305 $Y=0.235 $X2=0 $Y2=0
cc_444 N_Y_M1012_s N_VGND_c_895_n 0.00256987f $X=5.245 $Y=0.235 $X2=0 $Y2=0
cc_445 N_Y_M1018_s N_VGND_c_895_n 0.00256987f $X=6.185 $Y=0.235 $X2=0 $Y2=0
cc_446 N_Y_M1029_s N_VGND_c_895_n 0.00297142f $X=7.125 $Y=0.235 $X2=0 $Y2=0
cc_447 N_A_27_47#_c_752_n N_VGND_M1008_d 0.00251598f $X=0.985 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_448 N_A_27_47#_c_754_n N_VGND_M1011_d 0.00251598f $X=1.925 $Y=0.82 $X2=0
+ $Y2=0
cc_449 N_A_27_47#_c_755_n N_VGND_M1023_d 0.00251598f $X=2.865 $Y=0.82 $X2=0
+ $Y2=0
cc_450 N_A_27_47#_c_756_n N_VGND_M1027_d 0.00349437f $X=3.805 $Y=0.82 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_c_751_n N_VGND_c_886_n 0.0187901f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_452 N_A_27_47#_c_752_n N_VGND_c_886_n 0.0127122f $X=0.985 $Y=0.82 $X2=0 $Y2=0
cc_453 N_A_27_47#_c_752_n N_VGND_c_887_n 0.00193763f $X=0.985 $Y=0.82 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_c_770_n N_VGND_c_887_n 0.0223596f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_455 N_A_27_47#_c_754_n N_VGND_c_887_n 0.00260082f $X=1.925 $Y=0.82 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_c_770_n N_VGND_c_888_n 0.0189749f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_457 N_A_27_47#_c_754_n N_VGND_c_888_n 0.0127122f $X=1.925 $Y=0.82 $X2=0 $Y2=0
cc_458 N_A_27_47#_c_754_n N_VGND_c_889_n 0.00193763f $X=1.925 $Y=0.82 $X2=0
+ $Y2=0
cc_459 N_A_27_47#_c_778_n N_VGND_c_889_n 0.0223596f $X=2.14 $Y=0.4 $X2=0 $Y2=0
cc_460 N_A_27_47#_c_755_n N_VGND_c_889_n 0.00260082f $X=2.865 $Y=0.82 $X2=0
+ $Y2=0
cc_461 N_A_27_47#_c_778_n N_VGND_c_890_n 0.0189749f $X=2.14 $Y=0.4 $X2=0 $Y2=0
cc_462 N_A_27_47#_c_755_n N_VGND_c_890_n 0.0127122f $X=2.865 $Y=0.82 $X2=0 $Y2=0
cc_463 N_A_27_47#_c_786_n N_VGND_c_891_n 0.0189749f $X=3.08 $Y=0.4 $X2=0 $Y2=0
cc_464 N_A_27_47#_c_756_n N_VGND_c_891_n 0.013183f $X=3.805 $Y=0.82 $X2=0 $Y2=0
cc_465 N_A_27_47#_c_794_n N_VGND_c_891_n 0.0180776f $X=3.955 $Y=0.485 $X2=0
+ $Y2=0
cc_466 N_A_27_47#_c_757_n N_VGND_c_891_n 0.00582645f $X=3.955 $Y=0.735 $X2=0
+ $Y2=0
cc_467 N_A_27_47#_c_755_n N_VGND_c_892_n 0.00193763f $X=2.865 $Y=0.82 $X2=0
+ $Y2=0
cc_468 N_A_27_47#_c_786_n N_VGND_c_892_n 0.0223596f $X=3.08 $Y=0.4 $X2=0 $Y2=0
cc_469 N_A_27_47#_c_756_n N_VGND_c_892_n 0.00260082f $X=3.805 $Y=0.82 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_c_756_n N_VGND_c_894_n 0.00194552f $X=3.805 $Y=0.82 $X2=0
+ $Y2=0
cc_471 N_A_27_47#_c_794_n N_VGND_c_894_n 0.0186086f $X=3.955 $Y=0.485 $X2=0
+ $Y2=0
cc_472 N_A_27_47#_c_809_n N_VGND_c_894_n 0.203322f $X=7.695 $Y=0.37 $X2=0 $Y2=0
cc_473 N_A_27_47#_c_758_n N_VGND_c_894_n 0.0261024f $X=7.882 $Y=0.485 $X2=0
+ $Y2=0
cc_474 N_A_27_47#_M1008_s N_VGND_c_895_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_475 N_A_27_47#_M1010_s N_VGND_c_895_n 0.0025535f $X=1.015 $Y=0.235 $X2=0
+ $Y2=0
cc_476 N_A_27_47#_M1015_s N_VGND_c_895_n 0.0025535f $X=1.955 $Y=0.235 $X2=0
+ $Y2=0
cc_477 N_A_27_47#_M1025_s N_VGND_c_895_n 0.0025535f $X=2.895 $Y=0.235 $X2=0
+ $Y2=0
cc_478 N_A_27_47#_M1028_s N_VGND_c_895_n 0.00215206f $X=3.885 $Y=0.235 $X2=0
+ $Y2=0
cc_479 N_A_27_47#_M1006_d N_VGND_c_895_n 0.00255381f $X=4.775 $Y=0.235 $X2=0
+ $Y2=0
cc_480 N_A_27_47#_M1016_d N_VGND_c_895_n 0.00255381f $X=5.715 $Y=0.235 $X2=0
+ $Y2=0
cc_481 N_A_27_47#_M1019_d N_VGND_c_895_n 0.00255381f $X=6.655 $Y=0.235 $X2=0
+ $Y2=0
cc_482 N_A_27_47#_M1030_d N_VGND_c_895_n 0.00308503f $X=7.645 $Y=0.235 $X2=0
+ $Y2=0
cc_483 N_A_27_47#_c_751_n N_VGND_c_895_n 0.0126042f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_484 N_A_27_47#_c_752_n N_VGND_c_895_n 0.00961016f $X=0.985 $Y=0.82 $X2=0
+ $Y2=0
cc_485 N_A_27_47#_c_770_n N_VGND_c_895_n 0.0141302f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_486 N_A_27_47#_c_754_n N_VGND_c_895_n 0.00961016f $X=1.925 $Y=0.82 $X2=0
+ $Y2=0
cc_487 N_A_27_47#_c_778_n N_VGND_c_895_n 0.0141302f $X=2.14 $Y=0.4 $X2=0 $Y2=0
cc_488 N_A_27_47#_c_755_n N_VGND_c_895_n 0.00961016f $X=2.865 $Y=0.82 $X2=0
+ $Y2=0
cc_489 N_A_27_47#_c_786_n N_VGND_c_895_n 0.0141302f $X=3.08 $Y=0.4 $X2=0 $Y2=0
cc_490 N_A_27_47#_c_756_n N_VGND_c_895_n 0.00990055f $X=3.805 $Y=0.82 $X2=0
+ $Y2=0
cc_491 N_A_27_47#_c_794_n N_VGND_c_895_n 0.0111017f $X=3.955 $Y=0.485 $X2=0
+ $Y2=0
cc_492 N_A_27_47#_c_809_n N_VGND_c_895_n 0.12862f $X=7.695 $Y=0.37 $X2=0 $Y2=0
cc_493 N_A_27_47#_c_758_n N_VGND_c_895_n 0.0144249f $X=7.882 $Y=0.485 $X2=0
+ $Y2=0
cc_494 N_A_27_47#_c_751_n N_VGND_c_896_n 0.0213324f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_495 N_A_27_47#_c_752_n N_VGND_c_896_n 0.00260082f $X=0.985 $Y=0.82 $X2=0
+ $Y2=0
