* File: sky130_fd_sc_hdll__a21bo_2.spice
* Created: Thu Aug 27 18:52:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a21bo_2.pex.spice"
.subckt sky130_fd_sc_hdll__a21bo_2  VNB VPB B1_N A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_79_21#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.1235 PD=1.82 PS=1.03 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75000.2
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1010_d N_A_79_21#_M1010_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.131671 AS=0.1235 PD=1.2271 PS=1.03 NRD=1.836 NRS=9.228 M=1 R=4.33333
+ SA=75000.7 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1006 N_A_317_93#_M1006_d N_B1_N_M1006_g N_VGND_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1302 AS=0.0850794 PD=1.46 PS=0.792897 NRD=12.852 NRS=17.136 M=1
+ R=2.8 SA=75001.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_79_21#_M1011_d N_A_317_93#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.10725 AS=0.2015 PD=0.98 PS=1.92 NRD=1.836 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1000 A_621_47# N_A1_M1000_g N_A_79_21#_M1011_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.10725 PD=0.92 PS=0.98 NRD=14.76 NRS=7.38 M=1 R=4.33333
+ SA=75000.7 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g A_621_47# VNB NSHORT L=0.15 W=0.65 AD=0.2015
+ AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=14.76 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1003_d N_A_79_21#_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.27 PD=1.3 PS=2.54 NRD=1.9503 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90001 A=0.18 P=2.36 MULT=1
MM1007 N_X_M1003_d N_A_79_21#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.265634 PD=1.3 PS=2.15493 NRD=1.9503 NRS=19.7 M=1 R=5.55556
+ SA=90000.7 SB=90000.5 A=0.18 P=2.36 MULT=1
MM1008 N_A_317_93#_M1008_d N_B1_N_M1008_g N_VPWR_M1007_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.111566 PD=1.38 PS=0.90507 NRD=2.3443 NRS=98.7955 M=1
+ R=2.33333 SA=90001.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1005 N_A_523_297#_M1005_d N_A_317_93#_M1005_g N_A_79_21#_M1005_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.15 AS=0.27 PD=1.3 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g N_A_523_297#_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.15 PD=1.29 PS=1.3 NRD=0.9653 NRS=2.9353 M=1 R=5.55556 SA=90000.7
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1009 N_A_523_297#_M1009_d N_A2_M1009_g N_VPWR_M1001_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
pX13_noxref noxref_13 B1_N B1_N PROBETYPE=1
c_36 VNB 0 6.51255e-20 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hdll__a21bo_2.pxi.spice"
*
.ends
*
*
