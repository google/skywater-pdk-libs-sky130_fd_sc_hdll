* File: sky130_fd_sc_hdll__or2_6.pex.spice
* Created: Thu Aug 27 19:23:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR2_6%A 1 3 4 6 7 9 10 12 13 19 20 25
c39 10 0 1.11304e-19 $X=0.985 $Y=1.41
r40 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.96 $Y=1.202
+ $X2=0.985 $Y2=1.202
r41 19 25 12.4773 $w=1.98e-07 $l=2.25e-07 $layer=LI1_cond $X=0.92 $Y=1.175
+ $X2=0.695 $Y2=1.175
r42 18 20 5.07368 $w=3.8e-07 $l=4e-08 $layer=POLY_cond $X=0.92 $Y=1.202 $X2=0.96
+ $Y2=1.202
r43 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.92
+ $Y=1.16 $X2=0.92 $Y2=1.16
r44 16 18 48.2 $w=3.8e-07 $l=3.8e-07 $layer=POLY_cond $X=0.54 $Y=1.202 $X2=0.92
+ $Y2=1.202
r45 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.54 $Y2=1.202
r46 13 25 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=0.69 $Y=1.175
+ $X2=0.695 $Y2=1.175
r47 10 21 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r48 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r49 7 20 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=0.96 $Y2=1.202
r50 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.96 $Y=0.995 $X2=0.96
+ $Y2=0.56
r51 4 16 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.54 $Y2=1.202
r52 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.54 $Y=0.995 $X2=0.54
+ $Y2=0.56
r53 1 15 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r54 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_6%B 1 3 4 6 7 9 10 12 13 19 20 25
r55 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.9 $Y=1.202
+ $X2=1.925 $Y2=1.202
r56 19 25 13.5864 $w=1.98e-07 $l=2.45e-07 $layer=LI1_cond $X=1.86 $Y=1.175
+ $X2=1.615 $Y2=1.175
r57 18 20 5.07368 $w=3.8e-07 $l=4e-08 $layer=POLY_cond $X=1.86 $Y=1.202 $X2=1.9
+ $Y2=1.202
r58 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.86
+ $Y=1.16 $X2=1.86 $Y2=1.16
r59 16 18 48.2 $w=3.8e-07 $l=3.8e-07 $layer=POLY_cond $X=1.48 $Y=1.202 $X2=1.86
+ $Y2=1.202
r60 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.48 $Y2=1.202
r61 13 25 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=1.61 $Y=1.175
+ $X2=1.615 $Y2=1.175
r62 10 21 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r63 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r64 7 20 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.9 $Y=0.995 $X2=1.9
+ $Y2=1.202
r65 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.9 $Y=0.995 $X2=1.9
+ $Y2=0.56
r66 4 16 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.48 $Y=0.995
+ $X2=1.48 $Y2=1.202
r67 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.48 $Y=0.995 $X2=1.48
+ $Y2=0.56
r68 1 15 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r69 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_6%A_123_47# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 39 40 42 43 45 48 50 51 54 58 60 63 65 71 74 76
+ 77 90
c182 76 0 1.11304e-19 $X=1.69 $Y=1.62
r183 90 91 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.24 $Y=1.202
+ $X2=5.265 $Y2=1.202
r184 89 90 54.7135 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.82 $Y=1.202
+ $X2=5.24 $Y2=1.202
r185 88 89 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=4.795 $Y=1.202
+ $X2=4.82 $Y2=1.202
r186 85 86 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=4.3 $Y=1.202
+ $X2=4.325 $Y2=1.202
r187 84 85 54.7135 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.88 $Y=1.202
+ $X2=4.3 $Y2=1.202
r188 83 84 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=3.855 $Y=1.202
+ $X2=3.88 $Y2=1.202
r189 82 83 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=3.385 $Y=1.202
+ $X2=3.855 $Y2=1.202
r190 81 82 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=3.36 $Y=1.202
+ $X2=3.385 $Y2=1.202
r191 78 79 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=2.915 $Y=1.202
+ $X2=2.94 $Y2=1.202
r192 72 88 14.9811 $w=3.7e-07 $l=1.15e-07 $layer=POLY_cond $X=4.68 $Y=1.202
+ $X2=4.795 $Y2=1.202
r193 72 86 46.2459 $w=3.7e-07 $l=3.55e-07 $layer=POLY_cond $X=4.68 $Y=1.202
+ $X2=4.325 $Y2=1.202
r194 71 72 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=4.68
+ $Y=1.16 $X2=4.68 $Y2=1.16
r195 69 81 49.5027 $w=3.7e-07 $l=3.8e-07 $layer=POLY_cond $X=2.98 $Y=1.202
+ $X2=3.36 $Y2=1.202
r196 69 79 5.21081 $w=3.7e-07 $l=4e-08 $layer=POLY_cond $X=2.98 $Y=1.202
+ $X2=2.94 $Y2=1.202
r197 68 71 94.2727 $w=1.98e-07 $l=1.7e-06 $layer=LI1_cond $X=2.98 $Y=1.175
+ $X2=4.68 $Y2=1.175
r198 68 69 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=2.98
+ $Y=1.16 $X2=2.98 $Y2=1.16
r199 66 77 0.966048 $w=2e-07 $l=9e-08 $layer=LI1_cond $X=2.375 $Y=1.175
+ $X2=2.285 $Y2=1.175
r200 66 68 33.55 $w=1.98e-07 $l=6.05e-07 $layer=LI1_cond $X=2.375 $Y=1.175
+ $X2=2.98 $Y2=1.175
r201 64 77 5.63431 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=2.285 $Y=1.275
+ $X2=2.285 $Y2=1.175
r202 64 65 10.4747 $w=1.78e-07 $l=1.7e-07 $layer=LI1_cond $X=2.285 $Y=1.275
+ $X2=2.285 $Y2=1.445
r203 63 77 5.63431 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=2.285 $Y=1.075
+ $X2=2.285 $Y2=1.175
r204 62 63 10.4747 $w=1.78e-07 $l=1.7e-07 $layer=LI1_cond $X=2.285 $Y=0.905
+ $X2=2.285 $Y2=1.075
r205 61 76 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=1.555
+ $X2=1.69 $Y2=1.555
r206 60 65 6.90553 $w=2.2e-07 $l=1.48324e-07 $layer=LI1_cond $X=2.195 $Y=1.555
+ $X2=2.285 $Y2=1.445
r207 60 61 17.8105 $w=2.18e-07 $l=3.4e-07 $layer=LI1_cond $X=2.195 $Y=1.555
+ $X2=1.855 $Y2=1.555
r208 59 74 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=1.855 $Y=0.82
+ $X2=1.69 $Y2=0.815
r209 58 62 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.195 $Y=0.82
+ $X2=2.285 $Y2=0.905
r210 58 59 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.195 $Y=0.82
+ $X2=1.855 $Y2=0.82
r211 52 74 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.69 $Y=0.725
+ $X2=1.69 $Y2=0.815
r212 52 54 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.69 $Y=0.725
+ $X2=1.69 $Y2=0.39
r213 50 74 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=1.525 $Y=0.815
+ $X2=1.69 $Y2=0.815
r214 50 51 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=1.525 $Y=0.815
+ $X2=0.915 $Y2=0.815
r215 46 51 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.75 $Y=0.725
+ $X2=0.915 $Y2=0.815
r216 46 48 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.75 $Y=0.725
+ $X2=0.75 $Y2=0.39
r217 43 91 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.265 $Y=1.41
+ $X2=5.265 $Y2=1.202
r218 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.265 $Y=1.41
+ $X2=5.265 $Y2=1.985
r219 40 90 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=1.202
r220 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=0.56
r221 37 89 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.82 $Y=0.995
+ $X2=4.82 $Y2=1.202
r222 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.82 $Y=0.995
+ $X2=4.82 $Y2=0.56
r223 34 88 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.795 $Y=1.41
+ $X2=4.795 $Y2=1.202
r224 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.795 $Y=1.41
+ $X2=4.795 $Y2=1.985
r225 31 86 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.325 $Y=1.41
+ $X2=4.325 $Y2=1.202
r226 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.325 $Y=1.41
+ $X2=4.325 $Y2=1.985
r227 28 85 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.3 $Y=0.995
+ $X2=4.3 $Y2=1.202
r228 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.3 $Y=0.995
+ $X2=4.3 $Y2=0.56
r229 25 84 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.88 $Y=0.995
+ $X2=3.88 $Y2=1.202
r230 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.88 $Y=0.995
+ $X2=3.88 $Y2=0.56
r231 22 83 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.855 $Y=1.41
+ $X2=3.855 $Y2=1.202
r232 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.855 $Y=1.41
+ $X2=3.855 $Y2=1.985
r233 19 82 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.385 $Y=1.41
+ $X2=3.385 $Y2=1.202
r234 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.385 $Y=1.41
+ $X2=3.385 $Y2=1.985
r235 16 81 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.36 $Y=0.995
+ $X2=3.36 $Y2=1.202
r236 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.36 $Y=0.995
+ $X2=3.36 $Y2=0.56
r237 13 79 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.94 $Y=0.995
+ $X2=2.94 $Y2=1.202
r238 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.94 $Y=0.995
+ $X2=2.94 $Y2=0.56
r239 10 78 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.915 $Y=1.41
+ $X2=2.915 $Y2=1.202
r240 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.915 $Y=1.41
+ $X2=2.915 $Y2=1.985
r241 3 76 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=1.62
r242 2 54 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.555
+ $Y=0.235 $X2=1.69 $Y2=0.39
r243 1 48 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.615
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_6%A_27_297# 1 2 3 10 12 14 16 17 18 22
r34 20 22 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=2.175 $Y=2.295
+ $X2=2.175 $Y2=2
r35 19 29 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.355 $Y=2.38
+ $X2=1.22 $Y2=2.38
r36 18 20 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.025 $Y=2.38
+ $X2=2.175 $Y2=2.295
r37 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.025 $Y=2.38
+ $X2=1.355 $Y2=2.38
r38 17 29 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=2.295
+ $X2=1.22 $Y2=2.38
r39 16 27 3.04322 $w=2.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.22 $Y=1.665
+ $X2=1.22 $Y2=1.56
r40 16 17 26.8903 $w=2.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.22 $Y=1.665
+ $X2=1.22 $Y2=2.295
r41 15 25 4.39997 $w=2.1e-07 $l=1.63e-07 $layer=LI1_cond $X=0.415 $Y=1.56
+ $X2=0.252 $Y2=1.56
r42 14 27 3.91272 $w=2.1e-07 $l=1.35e-07 $layer=LI1_cond $X=1.085 $Y=1.56
+ $X2=1.22 $Y2=1.56
r43 14 15 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=1.085 $Y=1.56
+ $X2=0.415 $Y2=1.56
r44 10 25 2.83434 $w=3.25e-07 $l=1.05e-07 $layer=LI1_cond $X=0.252 $Y=1.665
+ $X2=0.252 $Y2=1.56
r45 10 12 22.517 $w=3.23e-07 $l=6.35e-07 $layer=LI1_cond $X=0.252 $Y=1.665
+ $X2=0.252 $Y2=2.3
r46 3 22 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=2
r47 2 29 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.3
r48 2 27 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.62
r49 1 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r50 1 12 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_6%VPWR 1 2 3 4 5 18 22 28 32 36 39 40 42 43 45
+ 46 48 49 50 52 74 75 78
r79 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r80 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r81 72 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r82 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r83 69 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r84 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r85 66 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r86 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r87 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r88 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r89 60 63 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r90 60 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r91 59 62 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r92 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r93 57 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=2.72
+ $X2=0.75 $Y2=2.72
r94 57 59 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.915 $Y=2.72
+ $X2=1.15 $Y2=2.72
r95 52 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=2.72
+ $X2=0.75 $Y2=2.72
r96 52 54 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.585 $Y=2.72
+ $X2=0.23 $Y2=2.72
r97 50 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r98 50 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r99 48 71 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.365 $Y=2.72
+ $X2=5.29 $Y2=2.72
r100 48 49 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.365 $Y=2.72
+ $X2=5.5 $Y2=2.72
r101 47 74 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=5.635 $Y=2.72
+ $X2=5.75 $Y2=2.72
r102 47 49 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.635 $Y=2.72
+ $X2=5.5 $Y2=2.72
r103 45 68 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.425 $Y=2.72
+ $X2=4.37 $Y2=2.72
r104 45 46 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.425 $Y=2.72
+ $X2=4.56 $Y2=2.72
r105 44 71 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=4.695 $Y=2.72
+ $X2=5.29 $Y2=2.72
r106 44 46 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.695 $Y=2.72
+ $X2=4.56 $Y2=2.72
r107 42 65 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.485 $Y=2.72
+ $X2=3.45 $Y2=2.72
r108 42 43 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.485 $Y=2.72
+ $X2=3.62 $Y2=2.72
r109 41 68 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=4.37 $Y2=2.72
r110 41 43 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=3.62 $Y2=2.72
r111 39 62 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.53 $Y2=2.72
r112 39 40 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.68 $Y2=2.72
r113 38 65 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.815 $Y=2.72
+ $X2=3.45 $Y2=2.72
r114 38 40 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.815 $Y=2.72
+ $X2=2.68 $Y2=2.72
r115 34 49 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.5 $Y=2.635
+ $X2=5.5 $Y2=2.72
r116 34 36 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.5 $Y=2.635
+ $X2=5.5 $Y2=2
r117 30 46 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=2.635
+ $X2=4.56 $Y2=2.72
r118 30 32 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.56 $Y=2.635
+ $X2=4.56 $Y2=2
r119 26 43 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=2.635
+ $X2=3.62 $Y2=2.72
r120 26 28 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.62 $Y=2.635
+ $X2=3.62 $Y2=2
r121 22 25 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.68 $Y=1.66
+ $X2=2.68 $Y2=2.34
r122 20 40 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=2.635
+ $X2=2.68 $Y2=2.72
r123 20 25 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.68 $Y=2.635
+ $X2=2.68 $Y2=2.34
r124 16 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r125 16 18 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2
r126 5 36 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.355
+ $Y=1.485 $X2=5.5 $Y2=2
r127 4 32 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.415
+ $Y=1.485 $X2=4.56 $Y2=2
r128 3 28 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.475
+ $Y=1.485 $X2=3.62 $Y2=2
r129 2 25 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.555
+ $Y=1.485 $X2=2.68 $Y2=2.34
r130 2 22 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=2.555
+ $Y=1.485 $X2=2.68 $Y2=1.66
r131 1 18 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_6%X 1 2 3 4 5 6 21 23 25 27 28 29 33 37 39 41
+ 45 49 54 55 58 60 61
r101 59 61 8.21116 $w=3.98e-07 $l=2.85e-07 $layer=LI1_cond $X=5.215 $Y=0.905
+ $X2=5.215 $Y2=1.19
r102 59 60 3.0006 $w=3.35e-07 $l=1.16189e-07 $layer=LI1_cond $X=5.215 $Y=0.905
+ $X2=5.155 $Y2=0.815
r103 56 61 8.78738 $w=3.98e-07 $l=3.05e-07 $layer=LI1_cond $X=5.215 $Y=1.495
+ $X2=5.215 $Y2=1.19
r104 56 58 2.63236 $w=3.65e-07 $l=1.16619e-07 $layer=LI1_cond $X=5.215 $Y=1.495
+ $X2=5.14 $Y2=1.58
r105 47 60 3.0006 $w=3.35e-07 $l=1.63936e-07 $layer=LI1_cond $X=5.03 $Y=0.725
+ $X2=5.155 $Y2=0.815
r106 47 49 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.03 $Y=0.725
+ $X2=5.03 $Y2=0.42
r107 43 58 2.63236 $w=3.65e-07 $l=1.46458e-07 $layer=LI1_cond $X=5.03 $Y=1.665
+ $X2=5.14 $Y2=1.58
r108 43 45 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.03 $Y=1.665
+ $X2=5.03 $Y2=2.34
r109 42 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.255 $Y=1.58
+ $X2=4.09 $Y2=1.58
r110 41 58 4.19346 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=4.865 $Y=1.58
+ $X2=5.14 $Y2=1.58
r111 41 42 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.865 $Y=1.58
+ $X2=4.255 $Y2=1.58
r112 40 55 7.13466 $w=1.8e-07 $l=1.35e-07 $layer=LI1_cond $X=4.225 $Y=0.815
+ $X2=4.09 $Y2=0.815
r113 39 60 3.64962 $w=1.8e-07 $l=2.6e-07 $layer=LI1_cond $X=4.895 $Y=0.815
+ $X2=5.155 $Y2=0.815
r114 39 40 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=4.895 $Y=0.815
+ $X2=4.225 $Y2=0.815
r115 35 55 0.067832 $w=2.7e-07 $l=9e-08 $layer=LI1_cond $X=4.09 $Y=0.725
+ $X2=4.09 $Y2=0.815
r116 35 37 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.09 $Y=0.725
+ $X2=4.09 $Y2=0.42
r117 31 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.09 $Y=1.665
+ $X2=4.09 $Y2=1.58
r118 31 33 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.09 $Y=1.665
+ $X2=4.09 $Y2=2.34
r119 30 52 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.315 $Y=1.58
+ $X2=3.15 $Y2=1.58
r120 29 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.925 $Y=1.58
+ $X2=4.09 $Y2=1.58
r121 29 30 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.925 $Y=1.58
+ $X2=3.315 $Y2=1.58
r122 27 55 7.13466 $w=1.8e-07 $l=1.35e-07 $layer=LI1_cond $X=3.955 $Y=0.815
+ $X2=4.09 $Y2=0.815
r123 27 28 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=3.955 $Y=0.815
+ $X2=3.285 $Y2=0.815
r124 23 52 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.15 $Y=1.665
+ $X2=3.15 $Y2=1.58
r125 23 25 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.15 $Y=1.665
+ $X2=3.15 $Y2=2.34
r126 19 28 7.38573 $w=1.8e-07 $l=1.89737e-07 $layer=LI1_cond $X=3.135 $Y=0.725
+ $X2=3.285 $Y2=0.815
r127 19 21 11.7165 $w=2.98e-07 $l=3.05e-07 $layer=LI1_cond $X=3.135 $Y=0.725
+ $X2=3.135 $Y2=0.42
r128 6 58 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.885
+ $Y=1.485 $X2=5.03 $Y2=1.66
r129 6 45 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.885
+ $Y=1.485 $X2=5.03 $Y2=2.34
r130 5 54 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.945
+ $Y=1.485 $X2=4.09 $Y2=1.66
r131 5 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.945
+ $Y=1.485 $X2=4.09 $Y2=2.34
r132 4 52 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.005
+ $Y=1.485 $X2=3.15 $Y2=1.66
r133 4 25 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.005
+ $Y=1.485 $X2=3.15 $Y2=2.34
r134 3 49 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=4.895
+ $Y=0.235 $X2=5.03 $Y2=0.42
r135 2 37 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=3.955
+ $Y=0.235 $X2=4.09 $Y2=0.42
r136 1 21 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=3.015
+ $Y=0.235 $X2=3.15 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_6%VGND 1 2 3 4 5 6 19 21 23 27 33 37 41 45 48
+ 49 51 52 54 55 56 69 70 76 81 90
r95 89 90 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=0.235
+ $X2=2.815 $Y2=0.235
r96 87 89 0.934436 $w=6.38e-07 $l=5e-08 $layer=LI1_cond $X=2.68 $Y=0.235
+ $X2=2.73 $Y2=0.235
r97 85 87 2.80331 $w=6.38e-07 $l=1.5e-07 $layer=LI1_cond $X=2.53 $Y=0.235
+ $X2=2.68 $Y2=0.235
r98 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r99 83 85 7.84926 $w=6.38e-07 $l=4.2e-07 $layer=LI1_cond $X=2.11 $Y=0.235
+ $X2=2.53 $Y2=0.235
r100 80 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r101 79 83 0.747549 $w=6.38e-07 $l=4e-08 $layer=LI1_cond $X=2.07 $Y=0.235
+ $X2=2.11 $Y2=0.235
r102 79 81 8.17421 $w=6.38e-07 $l=4.5e-08 $layer=LI1_cond $X=2.07 $Y=0.235
+ $X2=2.025 $Y2=0.235
r103 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r104 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r105 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r106 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r107 67 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r108 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r109 64 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r110 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r111 61 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r112 61 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r113 60 90 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.45 $Y=0
+ $X2=2.815 $Y2=0
r114 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r115 56 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r116 56 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r117 54 66 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.29
+ $Y2=0
r118 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.5
+ $Y2=0
r119 53 69 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.665 $Y=0 $X2=5.75
+ $Y2=0
r120 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.665 $Y=0 $X2=5.5
+ $Y2=0
r121 51 63 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.395 $Y=0 $X2=4.37
+ $Y2=0
r122 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=0 $X2=4.56
+ $Y2=0
r123 50 66 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=4.725 $Y=0 $X2=5.29
+ $Y2=0
r124 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=0 $X2=4.56
+ $Y2=0
r125 48 60 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.455 $Y=0 $X2=3.45
+ $Y2=0
r126 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.455 $Y=0 $X2=3.62
+ $Y2=0
r127 47 63 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.785 $Y=0
+ $X2=4.37 $Y2=0
r128 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.785 $Y=0 $X2=3.62
+ $Y2=0
r129 43 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.5 $Y=0.085 $X2=5.5
+ $Y2=0
r130 43 45 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.5 $Y=0.085
+ $X2=5.5 $Y2=0.42
r131 39 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=0.085
+ $X2=4.56 $Y2=0
r132 39 41 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.56 $Y=0.085
+ $X2=4.56 $Y2=0.42
r133 35 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=0.085
+ $X2=3.62 $Y2=0
r134 35 37 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.62 $Y=0.085
+ $X2=3.62 $Y2=0.42
r135 31 87 5.8233 $w=2.7e-07 $l=3.2e-07 $layer=LI1_cond $X=2.68 $Y=0.555
+ $X2=2.68 $Y2=0.235
r136 31 33 7.89637 $w=2.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.68 $Y=0.555
+ $X2=2.68 $Y2=0.74
r137 30 76 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.22
+ $Y2=0
r138 30 81 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.355 $Y=0
+ $X2=2.025 $Y2=0
r139 25 76 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r140 25 27 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.39
r141 24 73 4.13993 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.415 $Y=0
+ $X2=0.207 $Y2=0
r142 23 76 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.085 $Y=0 $X2=1.22
+ $Y2=0
r143 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.085 $Y=0
+ $X2=0.415 $Y2=0
r144 19 73 3.14476 $w=2.7e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.207 $Y2=0
r145 19 21 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.39
r146 6 45 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=5.315
+ $Y=0.235 $X2=5.5 $Y2=0.42
r147 5 41 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=4.375
+ $Y=0.235 $X2=4.56 $Y2=0.42
r148 4 37 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=3.435
+ $Y=0.235 $X2=3.62 $Y2=0.42
r149 3 89 182 $w=1.7e-07 $l=8.24318e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.73 $Y2=0.38
r150 3 83 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.11 $Y2=0.39
r151 3 33 182 $w=1.7e-07 $l=9.75346e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.73 $Y2=0.74
r152 2 27 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.235 $X2=1.22 $Y2=0.39
r153 1 21 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

