* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_1449_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 VGND A2 a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_119_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_27_297# B1 a_869_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 Y A1 a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Y A1 a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 a_119_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 Y C1 a_869_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_27_297# B1 a_1057_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 a_869_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 VGND A2 a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_119_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_1057_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 Y C1 a_1449_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X26 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X27 a_869_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X30 a_119_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
