* File: sky130_fd_sc_hdll__a21oi_4.pxi.spice
* Created: Thu Aug 27 18:53:30 2020
* 
x_PM_SKY130_FD_SC_HDLL__A21OI_4%B1 N_B1_c_80_n N_B1_M1001_g N_B1_c_86_n
+ N_B1_M1006_g N_B1_c_87_n N_B1_M1009_g N_B1_c_81_n N_B1_M1003_g N_B1_c_88_n
+ N_B1_M1017_g N_B1_c_82_n N_B1_M1010_g N_B1_c_89_n N_B1_M1020_g N_B1_c_83_n
+ N_B1_M1013_g N_B1_c_84_n B1 N_B1_c_91_n N_B1_c_85_n B1
+ PM_SKY130_FD_SC_HDLL__A21OI_4%B1
x_PM_SKY130_FD_SC_HDLL__A21OI_4%A2 N_A2_c_155_n N_A2_M1005_g N_A2_c_156_n
+ N_A2_M1002_g N_A2_c_157_n N_A2_M1008_g N_A2_c_165_n N_A2_M1018_g N_A2_c_158_n
+ N_A2_M1011_g N_A2_c_166_n N_A2_M1021_g N_A2_c_159_n N_A2_M1014_g N_A2_c_167_n
+ N_A2_M1022_g N_A2_c_160_n N_A2_c_178_n N_A2_c_161_n N_A2_c_170_n A2
+ N_A2_c_162_n N_A2_c_163_n A2 PM_SKY130_FD_SC_HDLL__A21OI_4%A2
x_PM_SKY130_FD_SC_HDLL__A21OI_4%A1 N_A1_c_283_n N_A1_M1015_g N_A1_c_289_n
+ N_A1_M1000_g N_A1_c_284_n N_A1_M1016_g N_A1_c_290_n N_A1_M1004_g N_A1_c_285_n
+ N_A1_M1019_g N_A1_c_291_n N_A1_M1007_g N_A1_c_292_n N_A1_M1012_g N_A1_c_286_n
+ N_A1_M1023_g A1 N_A1_c_287_n N_A1_c_288_n A1 PM_SKY130_FD_SC_HDLL__A21OI_4%A1
x_PM_SKY130_FD_SC_HDLL__A21OI_4%A_28_297# N_A_28_297#_M1006_s
+ N_A_28_297#_M1009_s N_A_28_297#_M1020_s N_A_28_297#_M1000_s
+ N_A_28_297#_M1007_s N_A_28_297#_M1018_s N_A_28_297#_M1022_s
+ N_A_28_297#_c_411_p N_A_28_297#_c_356_n N_A_28_297#_c_358_n
+ N_A_28_297#_c_368_n N_A_28_297#_c_360_n N_A_28_297#_c_400_p
+ N_A_28_297#_c_373_n N_A_28_297#_c_404_p N_A_28_297#_c_374_n
+ N_A_28_297#_c_406_p N_A_28_297#_c_376_n N_A_28_297#_c_354_n
+ N_A_28_297#_c_355_n N_A_28_297#_c_382_n N_A_28_297#_c_383_n
+ N_A_28_297#_c_384_n PM_SKY130_FD_SC_HDLL__A21OI_4%A_28_297#
x_PM_SKY130_FD_SC_HDLL__A21OI_4%Y N_Y_M1001_s N_Y_M1010_s N_Y_M1015_d
+ N_Y_M1019_d N_Y_M1006_d N_Y_M1017_d N_Y_c_442_n N_Y_c_490_p N_Y_c_437_n
+ N_Y_c_438_n N_Y_c_439_n N_Y_c_452_n N_Y_c_456_n N_Y_c_459_n N_Y_c_440_n Y Y
+ PM_SKY130_FD_SC_HDLL__A21OI_4%Y
x_PM_SKY130_FD_SC_HDLL__A21OI_4%VPWR N_VPWR_M1002_d N_VPWR_M1004_d
+ N_VPWR_M1012_d N_VPWR_M1021_d N_VPWR_c_518_n N_VPWR_c_519_n N_VPWR_c_520_n
+ N_VPWR_c_521_n N_VPWR_c_522_n VPWR N_VPWR_c_523_n N_VPWR_c_524_n
+ N_VPWR_c_517_n N_VPWR_c_526_n N_VPWR_c_527_n
+ PM_SKY130_FD_SC_HDLL__A21OI_4%VPWR
x_PM_SKY130_FD_SC_HDLL__A21OI_4%VGND N_VGND_M1001_d N_VGND_M1003_d
+ N_VGND_M1013_d N_VGND_M1008_s N_VGND_M1014_s N_VGND_c_617_n N_VGND_c_618_n
+ N_VGND_c_619_n N_VGND_c_620_n N_VGND_c_621_n N_VGND_c_622_n N_VGND_c_623_n
+ N_VGND_c_624_n VGND N_VGND_c_625_n N_VGND_c_626_n N_VGND_c_627_n
+ N_VGND_c_628_n N_VGND_c_629_n N_VGND_c_630_n
+ PM_SKY130_FD_SC_HDLL__A21OI_4%VGND
x_PM_SKY130_FD_SC_HDLL__A21OI_4%A_502_47# N_A_502_47#_M1005_d
+ N_A_502_47#_M1016_s N_A_502_47#_M1023_s N_A_502_47#_M1011_d
+ N_A_502_47#_c_716_n N_A_502_47#_c_717_n N_A_502_47#_c_718_n
+ N_A_502_47#_c_714_n N_A_502_47#_c_715_n N_A_502_47#_c_729_n
+ PM_SKY130_FD_SC_HDLL__A21OI_4%A_502_47#
cc_1 VNB N_B1_c_80_n 0.0221271f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_2 VNB N_B1_c_81_n 0.0171082f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=0.995
cc_3 VNB N_B1_c_82_n 0.0171215f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=0.995
cc_4 VNB N_B1_c_83_n 0.0157109f $X=-0.19 $Y=-0.24 $X2=1.965 $Y2=0.995
cc_5 VNB N_B1_c_84_n 0.0126238f $X=-0.19 $Y=-0.24 $X2=0.4 $Y2=1.205
cc_6 VNB N_B1_c_85_n 0.094739f $X=-0.19 $Y=-0.24 $X2=1.94 $Y2=1.202
cc_7 VNB N_A2_c_155_n 0.0173014f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_8 VNB N_A2_c_156_n 0.0267126f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_9 VNB N_A2_c_157_n 0.0166784f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=1.41
cc_10 VNB N_A2_c_158_n 0.0169453f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.41
cc_11 VNB N_A2_c_159_n 0.0224545f $X=-0.19 $Y=-0.24 $X2=1.94 $Y2=1.41
cc_12 VNB N_A2_c_160_n 0.00160282f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_13 VNB N_A2_c_161_n 0.00246559f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A2_c_162_n 0.071595f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=1.225
cc_15 VNB N_A2_c_163_n 0.00961897f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A1_c_283_n 0.0169502f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_17 VNB N_A1_c_284_n 0.0167597f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=1.41
cc_18 VNB N_A1_c_285_n 0.0171831f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.41
cc_19 VNB N_A1_c_286_n 0.0170612f $X=-0.19 $Y=-0.24 $X2=1.965 $Y2=0.995
cc_20 VNB N_A1_c_287_n 0.00170867f $X=-0.19 $Y=-0.24 $X2=1.965 $Y2=1.202
cc_21 VNB N_A1_c_288_n 0.100305f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.225
cc_22 VNB N_Y_c_437_n 0.00435771f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.205
cc_23 VNB N_Y_c_438_n 4.39987e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_Y_c_439_n 0.0110362f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.202
cc_25 VNB N_Y_c_440_n 0.00656144f $X=-0.19 $Y=-0.24 $X2=1.94 $Y2=1.202
cc_26 VNB N_VPWR_c_517_n 0.269736f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.225
cc_27 VNB N_VGND_c_617_n 0.0103023f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=0.995
cc_28 VNB N_VGND_c_618_n 0.0252256f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=0.56
cc_29 VNB N_VGND_c_619_n 0.00253981f $X=-0.19 $Y=-0.24 $X2=1.965 $Y2=0.995
cc_30 VNB N_VGND_c_620_n 0.00479809f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.205
cc_31 VNB N_VGND_c_621_n 0.0140602f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_32 VNB N_VGND_c_622_n 0.0366224f $X=-0.19 $Y=-0.24 $X2=0.4 $Y2=1.205
cc_33 VNB N_VGND_c_623_n 0.0616803f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.202
cc_34 VNB N_VGND_c_624_n 0.00362451f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.202
cc_35 VNB N_VGND_c_625_n 0.0141146f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=1.202
cc_36 VNB N_VGND_c_626_n 0.0144566f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=1.202
cc_37 VNB N_VGND_c_627_n 0.020013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_628_n 0.00792098f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_629_n 0.00492389f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_630_n 0.318436f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_502_47#_c_714_n 0.00511141f $X=-0.19 $Y=-0.24 $X2=1.965 $Y2=0.56
cc_42 VNB N_A_502_47#_c_715_n 0.00336803f $X=-0.19 $Y=-0.24 $X2=1.965 $Y2=0.56
cc_43 VPB N_B1_c_86_n 0.0209716f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_44 VPB N_B1_c_87_n 0.0163179f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.41
cc_45 VPB N_B1_c_88_n 0.016301f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.41
cc_46 VPB N_B1_c_89_n 0.0159808f $X=-0.19 $Y=1.305 $X2=1.94 $Y2=1.41
cc_47 VPB N_B1_c_84_n 0.0114231f $X=-0.19 $Y=1.305 $X2=0.4 $Y2=1.205
cc_48 VPB N_B1_c_91_n 0.00789998f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.16
cc_49 VPB N_B1_c_85_n 0.056695f $X=-0.19 $Y=1.305 $X2=1.94 $Y2=1.202
cc_50 VPB N_A2_c_156_n 0.0268131f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_51 VPB N_A2_c_165_n 0.015572f $X=-0.19 $Y=1.305 $X2=1.005 $Y2=0.995
cc_52 VPB N_A2_c_166_n 0.0152827f $X=-0.19 $Y=1.305 $X2=1.485 $Y2=0.995
cc_53 VPB N_A2_c_167_n 0.0192237f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=0.995
cc_54 VPB N_A2_c_160_n 0.00278154f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_55 VPB N_A2_c_161_n 0.00198511f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A2_c_170_n 0.0124351f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.202
cc_57 VPB N_A2_c_162_n 0.0381099f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.225
cc_58 VPB N_A2_c_163_n 0.00733094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A1_c_289_n 0.0162831f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_60 VPB N_A1_c_290_n 0.0158207f $X=-0.19 $Y=1.305 $X2=1.005 $Y2=0.995
cc_61 VPB N_A1_c_291_n 0.0161f $X=-0.19 $Y=1.305 $X2=1.485 $Y2=0.995
cc_62 VPB N_A1_c_292_n 0.0159297f $X=-0.19 $Y=1.305 $X2=1.94 $Y2=1.41
cc_63 VPB N_A1_c_287_n 0.00799673f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=1.202
cc_64 VPB N_A1_c_288_n 0.0254225f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.225
cc_65 VPB N_A_28_297#_c_354_n 0.0112688f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.225
cc_66 VPB N_A_28_297#_c_355_n 0.0137952f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_Y_c_437_n 0.00239113f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.205
cc_68 VPB N_VPWR_c_518_n 0.0127542f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.41
cc_69 VPB N_VPWR_c_519_n 0.00538475f $X=-0.19 $Y=1.305 $X2=1.485 $Y2=0.995
cc_70 VPB N_VPWR_c_520_n 0.0127542f $X=-0.19 $Y=1.305 $X2=1.94 $Y2=1.41
cc_71 VPB N_VPWR_c_521_n 0.00547506f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=0.56
cc_72 VPB N_VPWR_c_522_n 0.012802f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.205
cc_73 VPB N_VPWR_c_523_n 0.0587039f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=1.105
cc_74 VPB N_VPWR_c_524_n 0.019782f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=1.202
cc_75 VPB N_VPWR_c_517_n 0.0511377f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.225
cc_76 VPB N_VPWR_c_526_n 0.00547506f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.225
cc_77 VPB N_VPWR_c_527_n 0.00538475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 N_B1_c_83_n N_A2_c_155_n 0.0219137f $X=1.965 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_79 N_B1_c_89_n N_A2_c_156_n 0.0303905f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_80 N_B1_c_85_n N_A2_c_156_n 0.0242965f $X=1.94 $Y=1.202 $X2=0 $Y2=0
cc_81 N_B1_c_89_n N_A2_c_160_n 2.30501e-19 $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_82 N_B1_c_85_n N_A2_c_160_n 5.82523e-19 $X=1.94 $Y=1.202 $X2=0 $Y2=0
cc_83 N_B1_c_89_n N_A2_c_178_n 8.31559e-19 $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_84 N_B1_c_84_n N_A_28_297#_c_356_n 0.00904145f $X=0.4 $Y=1.205 $X2=0 $Y2=0
cc_85 N_B1_c_85_n N_A_28_297#_c_356_n 0.00108268f $X=1.94 $Y=1.202 $X2=0 $Y2=0
cc_86 N_B1_c_86_n N_A_28_297#_c_358_n 0.0171395f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_87 N_B1_c_87_n N_A_28_297#_c_358_n 0.00835107f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_88 N_B1_c_87_n N_A_28_297#_c_360_n 0.00317151f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_89 N_B1_c_88_n N_A_28_297#_c_360_n 0.0116963f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_90 N_B1_c_89_n N_A_28_297#_c_360_n 0.0188757f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_91 N_B1_c_81_n N_Y_c_442_n 0.0126854f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_92 N_B1_c_82_n N_Y_c_442_n 0.012178f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_93 N_B1_c_91_n N_Y_c_442_n 0.0490888f $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_94 N_B1_c_85_n N_Y_c_442_n 0.0036769f $X=1.94 $Y=1.202 $X2=0 $Y2=0
cc_95 N_B1_c_88_n N_Y_c_437_n 0.00392192f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_96 N_B1_c_82_n N_Y_c_437_n 0.00232492f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_97 N_B1_c_89_n N_Y_c_437_n 0.00501647f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_98 N_B1_c_83_n N_Y_c_437_n 0.0026933f $X=1.965 $Y=0.995 $X2=0 $Y2=0
cc_99 N_B1_c_91_n N_Y_c_437_n 0.0309402f $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_100 N_B1_c_85_n N_Y_c_437_n 0.0223396f $X=1.94 $Y=1.202 $X2=0 $Y2=0
cc_101 N_B1_c_80_n N_Y_c_452_n 0.00328215f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_102 N_B1_c_81_n N_Y_c_452_n 2.56032e-19 $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_103 N_B1_c_91_n N_Y_c_452_n 0.0152916f $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_104 N_B1_c_85_n N_Y_c_452_n 0.00454554f $X=1.94 $Y=1.202 $X2=0 $Y2=0
cc_105 N_B1_c_82_n N_Y_c_456_n 7.47525e-19 $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_106 N_B1_c_83_n N_Y_c_456_n 0.00856383f $X=1.965 $Y=0.995 $X2=0 $Y2=0
cc_107 N_B1_c_85_n N_Y_c_456_n 0.00454735f $X=1.94 $Y=1.202 $X2=0 $Y2=0
cc_108 N_B1_c_87_n N_Y_c_459_n 0.0190823f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_109 N_B1_c_88_n N_Y_c_459_n 0.019681f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_110 N_B1_c_89_n N_Y_c_459_n 0.0142997f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_111 N_B1_c_91_n N_Y_c_459_n 0.0686865f $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_112 N_B1_c_85_n N_Y_c_459_n 0.0089946f $X=1.94 $Y=1.202 $X2=0 $Y2=0
cc_113 N_B1_c_86_n N_VPWR_c_523_n 0.00429453f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_114 N_B1_c_87_n N_VPWR_c_523_n 0.00429362f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_115 N_B1_c_88_n N_VPWR_c_523_n 0.00429201f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_116 N_B1_c_89_n N_VPWR_c_523_n 0.00429201f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_117 N_B1_c_86_n N_VPWR_c_517_n 0.00700742f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_118 N_B1_c_87_n N_VPWR_c_517_n 0.00611667f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_119 N_B1_c_88_n N_VPWR_c_517_n 0.00611655f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_120 N_B1_c_89_n N_VPWR_c_517_n 0.00620861f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_121 N_B1_c_89_n N_VPWR_c_526_n 0.00101785f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_122 N_B1_c_80_n N_VGND_c_618_n 0.0127302f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_123 N_B1_c_81_n N_VGND_c_618_n 8.03266e-19 $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_124 N_B1_c_84_n N_VGND_c_618_n 0.0216211f $X=0.4 $Y=1.205 $X2=0 $Y2=0
cc_125 N_B1_c_91_n N_VGND_c_618_n 0.00145496f $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_126 N_B1_c_85_n N_VGND_c_618_n 0.00650316f $X=1.94 $Y=1.202 $X2=0 $Y2=0
cc_127 N_B1_c_82_n N_VGND_c_619_n 5.59007e-19 $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_128 N_B1_c_83_n N_VGND_c_619_n 0.00908352f $X=1.965 $Y=0.995 $X2=0 $Y2=0
cc_129 N_B1_c_80_n N_VGND_c_625_n 0.00486043f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_130 N_B1_c_81_n N_VGND_c_625_n 0.00211056f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_131 N_B1_c_82_n N_VGND_c_626_n 0.00422112f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_132 N_B1_c_83_n N_VGND_c_626_n 0.00273834f $X=1.965 $Y=0.995 $X2=0 $Y2=0
cc_133 N_B1_c_80_n N_VGND_c_628_n 8.40243e-19 $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_134 N_B1_c_81_n N_VGND_c_628_n 0.0101283f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_135 N_B1_c_82_n N_VGND_c_628_n 0.00167859f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_136 N_B1_c_80_n N_VGND_c_630_n 0.00854904f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_137 N_B1_c_81_n N_VGND_c_630_n 0.00301339f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_138 N_B1_c_82_n N_VGND_c_630_n 0.00586009f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_139 N_B1_c_83_n N_VGND_c_630_n 0.00348353f $X=1.965 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A2_c_155_n N_A1_c_283_n 0.0204522f $X=2.435 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_141 N_A2_c_156_n N_A1_c_289_n 0.0360875f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A2_c_160_n N_A1_c_289_n 0.00164446f $X=2.415 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A2_c_170_n N_A1_c_289_n 0.0143516f $X=4.675 $Y=1.39 $X2=0 $Y2=0
cc_144 N_A2_c_170_n N_A1_c_290_n 0.0143377f $X=4.675 $Y=1.39 $X2=0 $Y2=0
cc_145 N_A2_c_170_n N_A1_c_291_n 0.0143377f $X=4.675 $Y=1.39 $X2=0 $Y2=0
cc_146 N_A2_c_165_n N_A1_c_292_n 0.0375476f $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A2_c_161_n N_A1_c_292_n 0.00187003f $X=4.99 $Y=1.39 $X2=0 $Y2=0
cc_148 N_A2_c_170_n N_A1_c_292_n 0.0165069f $X=4.675 $Y=1.39 $X2=0 $Y2=0
cc_149 N_A2_c_157_n N_A1_c_286_n 0.0159585f $X=4.835 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A2_c_156_n N_A1_c_287_n 8.87839e-19 $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A2_c_160_n N_A1_c_287_n 0.021768f $X=2.415 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A2_c_161_n N_A1_c_287_n 0.0144695f $X=4.99 $Y=1.39 $X2=0 $Y2=0
cc_153 N_A2_c_170_n N_A1_c_287_n 0.119955f $X=4.675 $Y=1.39 $X2=0 $Y2=0
cc_154 N_A2_c_162_n N_A1_c_287_n 2.91841e-19 $X=5.82 $Y=1.202 $X2=0 $Y2=0
cc_155 N_A2_c_156_n N_A1_c_288_n 0.0258418f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A2_c_160_n N_A1_c_288_n 0.00318127f $X=2.415 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A2_c_161_n N_A1_c_288_n 0.00481353f $X=4.99 $Y=1.39 $X2=0 $Y2=0
cc_158 N_A2_c_170_n N_A1_c_288_n 0.00833524f $X=4.675 $Y=1.39 $X2=0 $Y2=0
cc_159 N_A2_c_162_n N_A1_c_288_n 0.0159585f $X=5.82 $Y=1.202 $X2=0 $Y2=0
cc_160 N_A2_c_178_n N_A_28_297#_M1020_s 0.00251451f $X=2.645 $Y=1.592 $X2=0
+ $Y2=0
cc_161 N_A2_c_170_n N_A_28_297#_M1000_s 0.00199437f $X=4.675 $Y=1.39 $X2=0 $Y2=0
cc_162 N_A2_c_170_n N_A_28_297#_M1007_s 0.00199437f $X=4.675 $Y=1.39 $X2=0 $Y2=0
cc_163 N_A2_c_163_n N_A_28_297#_M1018_s 0.0020586f $X=5.855 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A2_c_163_n N_A_28_297#_M1022_s 0.0110191f $X=5.855 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A2_c_156_n N_A_28_297#_c_368_n 0.0153939f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A2_c_178_n N_A_28_297#_c_368_n 0.0179009f $X=2.645 $Y=1.592 $X2=0 $Y2=0
cc_167 N_A2_c_170_n N_A_28_297#_c_368_n 0.0239153f $X=4.675 $Y=1.39 $X2=0 $Y2=0
cc_168 N_A2_c_156_n N_A_28_297#_c_360_n 2.09297e-19 $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A2_c_178_n N_A_28_297#_c_360_n 0.00470781f $X=2.645 $Y=1.592 $X2=0
+ $Y2=0
cc_170 N_A2_c_170_n N_A_28_297#_c_373_n 0.0395601f $X=4.675 $Y=1.39 $X2=0 $Y2=0
cc_171 N_A2_c_165_n N_A_28_297#_c_374_n 0.0159406f $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A2_c_170_n N_A_28_297#_c_374_n 0.0408835f $X=4.675 $Y=1.39 $X2=0 $Y2=0
cc_173 N_A2_c_166_n N_A_28_297#_c_376_n 0.0155699f $X=5.34 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A2_c_167_n N_A_28_297#_c_376_n 0.0130581f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A2_c_162_n N_A_28_297#_c_376_n 9.2015e-19 $X=5.82 $Y=1.202 $X2=0 $Y2=0
cc_176 N_A2_c_163_n N_A_28_297#_c_376_n 0.0435578f $X=5.855 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A2_c_162_n N_A_28_297#_c_354_n 2.63297e-19 $X=5.82 $Y=1.202 $X2=0 $Y2=0
cc_178 N_A2_c_163_n N_A_28_297#_c_354_n 0.00909513f $X=5.855 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A2_c_170_n N_A_28_297#_c_382_n 0.0152498f $X=4.675 $Y=1.39 $X2=0 $Y2=0
cc_180 N_A2_c_170_n N_A_28_297#_c_383_n 0.0152498f $X=4.675 $Y=1.39 $X2=0 $Y2=0
cc_181 N_A2_c_162_n N_A_28_297#_c_384_n 6.34633e-19 $X=5.82 $Y=1.202 $X2=0 $Y2=0
cc_182 N_A2_c_163_n N_A_28_297#_c_384_n 0.0157187f $X=5.855 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A2_c_155_n N_Y_c_437_n 0.00207984f $X=2.435 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A2_c_156_n N_Y_c_437_n 0.0036557f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A2_c_160_n N_Y_c_437_n 0.0338869f $X=2.415 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A2_c_178_n N_Y_c_437_n 0.00488847f $X=2.645 $Y=1.592 $X2=0 $Y2=0
cc_187 N_A2_c_155_n N_Y_c_438_n 0.00502003f $X=2.435 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A2_c_156_n N_Y_c_438_n 0.00307593f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A2_c_170_n N_Y_c_439_n 0.00563538f $X=4.675 $Y=1.39 $X2=0 $Y2=0
cc_190 N_A2_c_156_n N_Y_c_459_n 9.28308e-19 $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_191 N_A2_c_155_n N_Y_c_440_n 0.00906787f $X=2.435 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A2_c_156_n N_Y_c_440_n 0.00271655f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A2_c_160_n N_Y_c_440_n 0.0311338f $X=2.415 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A2_c_178_n N_VPWR_M1002_d 5.2043e-19 $X=2.645 $Y=1.592 $X2=-0.19
+ $Y2=-0.24
cc_195 N_A2_c_170_n N_VPWR_M1002_d 0.00158005f $X=4.675 $Y=1.39 $X2=-0.19
+ $Y2=-0.24
cc_196 N_A2_c_170_n N_VPWR_M1004_d 0.00199924f $X=4.675 $Y=1.39 $X2=0 $Y2=0
cc_197 N_A2_c_161_n N_VPWR_M1012_d 4.21561e-19 $X=4.99 $Y=1.39 $X2=0 $Y2=0
cc_198 N_A2_c_170_n N_VPWR_M1012_d 0.00158005f $X=4.675 $Y=1.39 $X2=0 $Y2=0
cc_199 N_A2_c_163_n N_VPWR_M1021_d 0.00206343f $X=5.855 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A2_c_165_n N_VPWR_c_519_n 0.00633356f $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A2_c_166_n N_VPWR_c_519_n 4.76818e-19 $X=5.34 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A2_c_165_n N_VPWR_c_521_n 5.28045e-19 $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A2_c_166_n N_VPWR_c_521_n 0.00901119f $X=5.34 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A2_c_167_n N_VPWR_c_521_n 0.00787483f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A2_c_165_n N_VPWR_c_522_n 0.00464324f $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A2_c_166_n N_VPWR_c_522_n 0.0032362f $X=5.34 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A2_c_156_n N_VPWR_c_523_n 0.0035176f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A2_c_167_n N_VPWR_c_524_n 0.00464324f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A2_c_156_n N_VPWR_c_517_n 0.00421648f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A2_c_165_n N_VPWR_c_517_n 0.00525281f $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A2_c_166_n N_VPWR_c_517_n 0.00384231f $X=5.34 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A2_c_167_n N_VPWR_c_517_n 0.00623601f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_213 N_A2_c_156_n N_VPWR_c_526_n 0.00947287f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A2_c_155_n N_VGND_c_619_n 0.0029807f $X=2.435 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A2_c_157_n N_VGND_c_620_n 0.00393281f $X=4.835 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A2_c_158_n N_VGND_c_620_n 0.00283414f $X=5.315 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A2_c_159_n N_VGND_c_622_n 0.00676599f $X=5.795 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A2_c_162_n N_VGND_c_622_n 0.00188138f $X=5.82 $Y=1.202 $X2=0 $Y2=0
cc_219 N_A2_c_163_n N_VGND_c_622_n 0.00838944f $X=5.855 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A2_c_155_n N_VGND_c_623_n 0.00420889f $X=2.435 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A2_c_157_n N_VGND_c_623_n 0.00425616f $X=4.835 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A2_c_158_n N_VGND_c_627_n 0.00427134f $X=5.315 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A2_c_159_n N_VGND_c_627_n 0.0054895f $X=5.795 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A2_c_155_n N_VGND_c_630_n 0.00598901f $X=2.435 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A2_c_157_n N_VGND_c_630_n 0.00608935f $X=4.835 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A2_c_158_n N_VGND_c_630_n 0.00605404f $X=5.315 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A2_c_159_n N_VGND_c_630_n 0.0110352f $X=5.795 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A2_c_155_n N_A_502_47#_c_716_n 0.0030746f $X=2.435 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A2_c_157_n N_A_502_47#_c_717_n 0.00305602f $X=4.835 $Y=0.995 $X2=0
+ $Y2=0
cc_230 N_A2_c_157_n N_A_502_47#_c_718_n 0.00379892f $X=4.835 $Y=0.995 $X2=0
+ $Y2=0
cc_231 N_A2_c_158_n N_A_502_47#_c_718_n 4.67045e-19 $X=5.315 $Y=0.995 $X2=0
+ $Y2=0
cc_232 N_A2_c_157_n N_A_502_47#_c_714_n 0.0091282f $X=4.835 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A2_c_158_n N_A_502_47#_c_714_n 0.0100639f $X=5.315 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A2_c_159_n N_A_502_47#_c_714_n 0.00334971f $X=5.795 $Y=0.995 $X2=0
+ $Y2=0
cc_235 N_A2_c_161_n N_A_502_47#_c_714_n 0.0448084f $X=4.99 $Y=1.39 $X2=0 $Y2=0
cc_236 N_A2_c_162_n N_A_502_47#_c_714_n 0.00753606f $X=5.82 $Y=1.202 $X2=0 $Y2=0
cc_237 N_A2_c_163_n N_A_502_47#_c_714_n 0.0331939f $X=5.855 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A2_c_157_n N_A_502_47#_c_715_n 9.23859e-19 $X=4.835 $Y=0.995 $X2=0
+ $Y2=0
cc_239 N_A2_c_161_n N_A_502_47#_c_715_n 0.00994332f $X=4.99 $Y=1.39 $X2=0 $Y2=0
cc_240 N_A2_c_170_n N_A_502_47#_c_715_n 0.00548957f $X=4.675 $Y=1.39 $X2=0 $Y2=0
cc_241 N_A2_c_157_n N_A_502_47#_c_729_n 5.23745e-19 $X=4.835 $Y=0.995 $X2=0
+ $Y2=0
cc_242 N_A2_c_158_n N_A_502_47#_c_729_n 0.00648408f $X=5.315 $Y=0.995 $X2=0
+ $Y2=0
cc_243 N_A2_c_159_n N_A_502_47#_c_729_n 0.00592327f $X=5.795 $Y=0.995 $X2=0
+ $Y2=0
cc_244 N_A1_c_289_n N_A_28_297#_c_368_n 0.0130725f $X=2.94 $Y=1.41 $X2=0 $Y2=0
cc_245 N_A1_c_290_n N_A_28_297#_c_373_n 0.0126261f $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_246 N_A1_c_291_n N_A_28_297#_c_373_n 0.0130581f $X=3.9 $Y=1.41 $X2=0 $Y2=0
cc_247 N_A1_c_292_n N_A_28_297#_c_374_n 0.0125649f $X=4.38 $Y=1.41 $X2=0 $Y2=0
cc_248 N_A1_c_283_n N_Y_c_439_n 0.0101935f $X=2.915 $Y=0.99 $X2=0 $Y2=0
cc_249 N_A1_c_284_n N_Y_c_439_n 0.0102676f $X=3.395 $Y=0.99 $X2=0 $Y2=0
cc_250 N_A1_c_285_n N_Y_c_439_n 0.0102651f $X=3.875 $Y=0.99 $X2=0 $Y2=0
cc_251 N_A1_c_287_n N_Y_c_439_n 0.110088f $X=4.215 $Y=1.16 $X2=0 $Y2=0
cc_252 N_A1_c_288_n N_Y_c_439_n 0.0121329f $X=4.38 $Y=1.2 $X2=0 $Y2=0
cc_253 N_A1_c_289_n N_VPWR_c_518_n 0.00464324f $X=2.94 $Y=1.41 $X2=0 $Y2=0
cc_254 N_A1_c_290_n N_VPWR_c_518_n 0.0032362f $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_255 N_A1_c_291_n N_VPWR_c_519_n 5.25185e-19 $X=3.9 $Y=1.41 $X2=0 $Y2=0
cc_256 N_A1_c_292_n N_VPWR_c_519_n 0.00893271f $X=4.38 $Y=1.41 $X2=0 $Y2=0
cc_257 N_A1_c_291_n N_VPWR_c_520_n 0.00464324f $X=3.9 $Y=1.41 $X2=0 $Y2=0
cc_258 N_A1_c_292_n N_VPWR_c_520_n 0.0032362f $X=4.38 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A1_c_289_n N_VPWR_c_517_n 0.00525281f $X=2.94 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A1_c_290_n N_VPWR_c_517_n 0.00384231f $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A1_c_291_n N_VPWR_c_517_n 0.00525281f $X=3.9 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A1_c_292_n N_VPWR_c_517_n 0.00384231f $X=4.38 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A1_c_289_n N_VPWR_c_526_n 0.00637633f $X=2.94 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A1_c_290_n N_VPWR_c_526_n 4.76818e-19 $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A1_c_289_n N_VPWR_c_527_n 5.25185e-19 $X=2.94 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A1_c_290_n N_VPWR_c_527_n 0.00896733f $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_267 N_A1_c_291_n N_VPWR_c_527_n 0.00636819f $X=3.9 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A1_c_292_n N_VPWR_c_527_n 4.76818e-19 $X=4.38 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A1_c_283_n N_VGND_c_623_n 0.00357877f $X=2.915 $Y=0.99 $X2=0 $Y2=0
cc_270 N_A1_c_284_n N_VGND_c_623_n 0.00357877f $X=3.395 $Y=0.99 $X2=0 $Y2=0
cc_271 N_A1_c_285_n N_VGND_c_623_n 0.00357877f $X=3.875 $Y=0.99 $X2=0 $Y2=0
cc_272 N_A1_c_286_n N_VGND_c_623_n 0.00357877f $X=4.405 $Y=0.99 $X2=0 $Y2=0
cc_273 N_A1_c_283_n N_VGND_c_630_n 0.0055497f $X=2.915 $Y=0.99 $X2=0 $Y2=0
cc_274 N_A1_c_284_n N_VGND_c_630_n 0.00553284f $X=3.395 $Y=0.99 $X2=0 $Y2=0
cc_275 N_A1_c_285_n N_VGND_c_630_n 0.00565034f $X=3.875 $Y=0.99 $X2=0 $Y2=0
cc_276 N_A1_c_286_n N_VGND_c_630_n 0.00555112f $X=4.405 $Y=0.99 $X2=0 $Y2=0
cc_277 N_A1_c_283_n N_A_502_47#_c_716_n 0.0102247f $X=2.915 $Y=0.99 $X2=0 $Y2=0
cc_278 N_A1_c_284_n N_A_502_47#_c_716_n 0.0102247f $X=3.395 $Y=0.99 $X2=0 $Y2=0
cc_279 N_A1_c_285_n N_A_502_47#_c_716_n 0.0105968f $X=3.875 $Y=0.99 $X2=0 $Y2=0
cc_280 N_A1_c_286_n N_A_502_47#_c_716_n 0.0140518f $X=4.405 $Y=0.99 $X2=0 $Y2=0
cc_281 N_A1_c_287_n N_A_502_47#_c_716_n 0.00222247f $X=4.215 $Y=1.16 $X2=0 $Y2=0
cc_282 N_A1_c_286_n N_A_502_47#_c_715_n 4.30873e-19 $X=4.405 $Y=0.99 $X2=0 $Y2=0
cc_283 N_A_28_297#_c_358_n N_Y_M1006_d 0.00382218f $X=1.005 $Y=2.34 $X2=0 $Y2=0
cc_284 N_A_28_297#_c_360_n N_Y_M1017_d 0.00375826f $X=2.315 $Y=1.99 $X2=0 $Y2=0
cc_285 N_A_28_297#_M1009_s N_Y_c_459_n 0.0036356f $X=1.07 $Y=1.485 $X2=0 $Y2=0
cc_286 N_A_28_297#_c_358_n N_Y_c_459_n 0.0213875f $X=1.005 $Y=2.34 $X2=0 $Y2=0
cc_287 N_A_28_297#_c_360_n N_Y_c_459_n 0.0657293f $X=2.315 $Y=1.99 $X2=0 $Y2=0
cc_288 N_A_28_297#_c_368_n N_VPWR_M1002_d 0.00408766f $X=3.085 $Y=1.99 $X2=-0.19
+ $Y2=1.305
cc_289 N_A_28_297#_c_373_n N_VPWR_M1004_d 0.00373237f $X=4.045 $Y=1.99 $X2=0
+ $Y2=0
cc_290 N_A_28_297#_c_374_n N_VPWR_M1012_d 0.00391313f $X=5.005 $Y=1.99 $X2=0
+ $Y2=0
cc_291 N_A_28_297#_c_376_n N_VPWR_M1021_d 0.00371742f $X=5.965 $Y=1.99 $X2=0
+ $Y2=0
cc_292 N_A_28_297#_c_368_n N_VPWR_c_518_n 0.00344373f $X=3.085 $Y=1.99 $X2=0
+ $Y2=0
cc_293 N_A_28_297#_c_400_p N_VPWR_c_518_n 0.0130156f $X=3.18 $Y=2.3 $X2=0 $Y2=0
cc_294 N_A_28_297#_c_373_n N_VPWR_c_518_n 0.00256992f $X=4.045 $Y=1.99 $X2=0
+ $Y2=0
cc_295 N_A_28_297#_c_374_n N_VPWR_c_519_n 0.0199464f $X=5.005 $Y=1.99 $X2=0
+ $Y2=0
cc_296 N_A_28_297#_c_373_n N_VPWR_c_520_n 0.00344373f $X=4.045 $Y=1.99 $X2=0
+ $Y2=0
cc_297 N_A_28_297#_c_404_p N_VPWR_c_520_n 0.0130156f $X=4.14 $Y=2.3 $X2=0 $Y2=0
cc_298 N_A_28_297#_c_374_n N_VPWR_c_520_n 0.00256992f $X=5.005 $Y=1.99 $X2=0
+ $Y2=0
cc_299 N_A_28_297#_c_406_p N_VPWR_c_521_n 0.0136279f $X=5.1 $Y=2.3 $X2=0 $Y2=0
cc_300 N_A_28_297#_c_376_n N_VPWR_c_521_n 0.0199464f $X=5.965 $Y=1.99 $X2=0
+ $Y2=0
cc_301 N_A_28_297#_c_374_n N_VPWR_c_522_n 0.00345089f $X=5.005 $Y=1.99 $X2=0
+ $Y2=0
cc_302 N_A_28_297#_c_406_p N_VPWR_c_522_n 0.0123537f $X=5.1 $Y=2.3 $X2=0 $Y2=0
cc_303 N_A_28_297#_c_376_n N_VPWR_c_522_n 0.00273875f $X=5.965 $Y=1.99 $X2=0
+ $Y2=0
cc_304 N_A_28_297#_c_411_p N_VPWR_c_523_n 0.0129329f $X=0.277 $Y=2.215 $X2=0
+ $Y2=0
cc_305 N_A_28_297#_c_358_n N_VPWR_c_523_n 0.0359212f $X=1.005 $Y=2.34 $X2=0
+ $Y2=0
cc_306 N_A_28_297#_c_368_n N_VPWR_c_523_n 0.00264869f $X=3.085 $Y=1.99 $X2=0
+ $Y2=0
cc_307 N_A_28_297#_c_360_n N_VPWR_c_523_n 0.0768983f $X=2.315 $Y=1.99 $X2=0
+ $Y2=0
cc_308 N_A_28_297#_c_376_n N_VPWR_c_524_n 0.00344373f $X=5.965 $Y=1.99 $X2=0
+ $Y2=0
cc_309 N_A_28_297#_c_355_n N_VPWR_c_524_n 0.0179734f $X=6.06 $Y=2.3 $X2=0 $Y2=0
cc_310 N_A_28_297#_M1006_s N_VPWR_c_517_n 0.00356383f $X=0.14 $Y=1.485 $X2=0
+ $Y2=0
cc_311 N_A_28_297#_M1009_s N_VPWR_c_517_n 0.00239291f $X=1.07 $Y=1.485 $X2=0
+ $Y2=0
cc_312 N_A_28_297#_M1020_s N_VPWR_c_517_n 0.00278173f $X=2.03 $Y=1.485 $X2=0
+ $Y2=0
cc_313 N_A_28_297#_M1000_s N_VPWR_c_517_n 0.00273993f $X=3.03 $Y=1.485 $X2=0
+ $Y2=0
cc_314 N_A_28_297#_M1007_s N_VPWR_c_517_n 0.00273993f $X=3.99 $Y=1.485 $X2=0
+ $Y2=0
cc_315 N_A_28_297#_M1018_s N_VPWR_c_517_n 0.00277355f $X=4.95 $Y=1.485 $X2=0
+ $Y2=0
cc_316 N_A_28_297#_M1022_s N_VPWR_c_517_n 0.00238967f $X=5.91 $Y=1.485 $X2=0
+ $Y2=0
cc_317 N_A_28_297#_c_411_p N_VPWR_c_517_n 0.00750689f $X=0.277 $Y=2.215 $X2=0
+ $Y2=0
cc_318 N_A_28_297#_c_358_n N_VPWR_c_517_n 0.0222394f $X=1.005 $Y=2.34 $X2=0
+ $Y2=0
cc_319 N_A_28_297#_c_368_n N_VPWR_c_517_n 0.0116231f $X=3.085 $Y=1.99 $X2=0
+ $Y2=0
cc_320 N_A_28_297#_c_360_n N_VPWR_c_517_n 0.0472839f $X=2.315 $Y=1.99 $X2=0
+ $Y2=0
cc_321 N_A_28_297#_c_400_p N_VPWR_c_517_n 0.00720328f $X=3.18 $Y=2.3 $X2=0 $Y2=0
cc_322 N_A_28_297#_c_373_n N_VPWR_c_517_n 0.0116586f $X=4.045 $Y=1.99 $X2=0
+ $Y2=0
cc_323 N_A_28_297#_c_404_p N_VPWR_c_517_n 0.00720328f $X=4.14 $Y=2.3 $X2=0 $Y2=0
cc_324 N_A_28_297#_c_374_n N_VPWR_c_517_n 0.0116694f $X=5.005 $Y=1.99 $X2=0
+ $Y2=0
cc_325 N_A_28_297#_c_406_p N_VPWR_c_517_n 0.00682467f $X=5.1 $Y=2.3 $X2=0 $Y2=0
cc_326 N_A_28_297#_c_376_n N_VPWR_c_517_n 0.0119605f $X=5.965 $Y=1.99 $X2=0
+ $Y2=0
cc_327 N_A_28_297#_c_355_n N_VPWR_c_517_n 0.00989423f $X=6.06 $Y=2.3 $X2=0 $Y2=0
cc_328 N_A_28_297#_c_368_n N_VPWR_c_526_n 0.0199956f $X=3.085 $Y=1.99 $X2=0
+ $Y2=0
cc_329 N_A_28_297#_c_373_n N_VPWR_c_527_n 0.0199464f $X=4.045 $Y=1.99 $X2=0
+ $Y2=0
cc_330 N_Y_M1006_d N_VPWR_c_517_n 0.00240926f $X=0.59 $Y=1.485 $X2=0 $Y2=0
cc_331 N_Y_M1017_d N_VPWR_c_517_n 0.00240897f $X=1.55 $Y=1.485 $X2=0 $Y2=0
cc_332 N_Y_c_442_n N_VGND_M1003_d 0.00419317f $X=1.605 $Y=0.74 $X2=0 $Y2=0
cc_333 N_Y_c_440_n N_VGND_M1013_d 0.00213857f $X=2.475 $Y=0.785 $X2=0 $Y2=0
cc_334 N_Y_c_452_n N_VGND_c_618_n 0.0265863f $X=0.74 $Y=0.535 $X2=0 $Y2=0
cc_335 N_Y_c_490_p N_VGND_c_619_n 0.0184469f $X=1.7 $Y=0.42 $X2=0 $Y2=0
cc_336 N_Y_c_456_n N_VGND_c_619_n 0.00430695f $X=1.7 $Y=0.76 $X2=0 $Y2=0
cc_337 N_Y_c_440_n N_VGND_c_619_n 0.0161669f $X=2.475 $Y=0.785 $X2=0 $Y2=0
cc_338 N_Y_c_440_n N_VGND_c_623_n 0.00202288f $X=2.475 $Y=0.785 $X2=0 $Y2=0
cc_339 N_Y_c_442_n N_VGND_c_625_n 0.00261192f $X=1.605 $Y=0.74 $X2=0 $Y2=0
cc_340 N_Y_c_452_n N_VGND_c_625_n 0.00739218f $X=0.74 $Y=0.535 $X2=0 $Y2=0
cc_341 N_Y_c_442_n N_VGND_c_626_n 0.00335005f $X=1.605 $Y=0.74 $X2=0 $Y2=0
cc_342 N_Y_c_490_p N_VGND_c_626_n 0.012763f $X=1.7 $Y=0.42 $X2=0 $Y2=0
cc_343 N_Y_c_456_n N_VGND_c_626_n 0.00260458f $X=1.7 $Y=0.76 $X2=0 $Y2=0
cc_344 N_Y_c_442_n N_VGND_c_628_n 0.0221395f $X=1.605 $Y=0.74 $X2=0 $Y2=0
cc_345 N_Y_c_452_n N_VGND_c_628_n 0.00564498f $X=0.74 $Y=0.535 $X2=0 $Y2=0
cc_346 N_Y_M1001_s N_VGND_c_630_n 0.00681879f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_347 N_Y_M1010_s N_VGND_c_630_n 0.00321424f $X=1.56 $Y=0.235 $X2=0 $Y2=0
cc_348 N_Y_M1015_d N_VGND_c_630_n 0.00265018f $X=2.99 $Y=0.235 $X2=0 $Y2=0
cc_349 N_Y_M1019_d N_VGND_c_630_n 0.00305172f $X=3.95 $Y=0.235 $X2=0 $Y2=0
cc_350 N_Y_c_442_n N_VGND_c_630_n 0.0119527f $X=1.605 $Y=0.74 $X2=0 $Y2=0
cc_351 N_Y_c_490_p N_VGND_c_630_n 0.00722448f $X=1.7 $Y=0.42 $X2=0 $Y2=0
cc_352 N_Y_c_438_n N_VGND_c_630_n 0.00352838f $X=2.585 $Y=0.785 $X2=0 $Y2=0
cc_353 N_Y_c_452_n N_VGND_c_630_n 0.00672198f $X=0.74 $Y=0.535 $X2=0 $Y2=0
cc_354 N_Y_c_456_n N_VGND_c_630_n 0.00537059f $X=1.7 $Y=0.76 $X2=0 $Y2=0
cc_355 N_Y_c_440_n N_VGND_c_630_n 0.00467993f $X=2.475 $Y=0.785 $X2=0 $Y2=0
cc_356 N_Y_c_439_n N_A_502_47#_M1005_d 0.0020497f $X=4.14 $Y=0.76 $X2=-0.19
+ $Y2=-0.24
cc_357 N_Y_c_439_n N_A_502_47#_M1016_s 0.00224739f $X=4.14 $Y=0.76 $X2=0 $Y2=0
cc_358 N_Y_M1015_d N_A_502_47#_c_716_n 0.00419532f $X=2.99 $Y=0.235 $X2=0 $Y2=0
cc_359 N_Y_M1019_d N_A_502_47#_c_716_n 0.00542196f $X=3.95 $Y=0.235 $X2=0 $Y2=0
cc_360 N_Y_c_438_n N_A_502_47#_c_716_n 0.098658f $X=2.585 $Y=0.785 $X2=0 $Y2=0
cc_361 N_Y_c_439_n N_A_502_47#_c_715_n 6.23804e-19 $X=4.14 $Y=0.76 $X2=0 $Y2=0
cc_362 N_VGND_c_630_n N_A_502_47#_M1005_d 0.00263412f $X=6.21 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_363 N_VGND_c_630_n N_A_502_47#_M1016_s 0.00263412f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_364 N_VGND_c_630_n N_A_502_47#_M1023_s 0.00223235f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_365 N_VGND_c_630_n N_A_502_47#_M1011_d 0.0026338f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_366 N_VGND_c_623_n N_A_502_47#_c_716_n 0.116449f $X=5.005 $Y=0 $X2=0 $Y2=0
cc_367 N_VGND_c_630_n N_A_502_47#_c_716_n 0.0734159f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_368 N_VGND_c_620_n N_A_502_47#_c_717_n 0.0162142f $X=5.1 $Y=0.4 $X2=0 $Y2=0
cc_369 N_VGND_c_623_n N_A_502_47#_c_717_n 0.0157493f $X=5.005 $Y=0 $X2=0 $Y2=0
cc_370 N_VGND_c_630_n N_A_502_47#_c_717_n 0.00981451f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_371 N_VGND_c_620_n N_A_502_47#_c_718_n 0.0035677f $X=5.1 $Y=0.4 $X2=0 $Y2=0
cc_372 N_VGND_M1008_s N_A_502_47#_c_714_n 0.00257482f $X=4.91 $Y=0.235 $X2=0
+ $Y2=0
cc_373 N_VGND_c_620_n N_A_502_47#_c_714_n 0.0138893f $X=5.1 $Y=0.4 $X2=0 $Y2=0
cc_374 N_VGND_c_622_n N_A_502_47#_c_714_n 0.00994924f $X=6.06 $Y=0.38 $X2=0
+ $Y2=0
cc_375 N_VGND_c_623_n N_A_502_47#_c_714_n 0.00259539f $X=5.005 $Y=0 $X2=0 $Y2=0
cc_376 N_VGND_c_627_n N_A_502_47#_c_714_n 0.00196536f $X=5.965 $Y=0 $X2=0 $Y2=0
cc_377 N_VGND_c_630_n N_A_502_47#_c_714_n 0.00963523f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_378 N_VGND_c_622_n N_A_502_47#_c_729_n 0.0302955f $X=6.06 $Y=0.38 $X2=0 $Y2=0
cc_379 N_VGND_c_627_n N_A_502_47#_c_729_n 0.0223809f $X=5.965 $Y=0 $X2=0 $Y2=0
cc_380 N_VGND_c_630_n N_A_502_47#_c_729_n 0.014176f $X=6.21 $Y=0 $X2=0 $Y2=0
