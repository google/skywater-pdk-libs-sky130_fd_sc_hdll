* File: sky130_fd_sc_hdll__and3_1.pxi.spice
* Created: Wed Sep  2 08:22:11 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND3_1%A N_A_c_48_n N_A_M1002_g N_A_c_49_n N_A_M1006_g A
+ PM_SKY130_FD_SC_HDLL__AND3_1%A
x_PM_SKY130_FD_SC_HDLL__AND3_1%B N_B_c_76_n N_B_M1007_g N_B_M1001_g N_B_c_75_n B
+ B PM_SKY130_FD_SC_HDLL__AND3_1%B
x_PM_SKY130_FD_SC_HDLL__AND3_1%C N_C_c_109_n N_C_M1004_g N_C_M1003_g C
+ PM_SKY130_FD_SC_HDLL__AND3_1%C
x_PM_SKY130_FD_SC_HDLL__AND3_1%A_27_47# N_A_27_47#_M1006_s N_A_27_47#_M1002_s
+ N_A_27_47#_M1007_d N_A_27_47#_c_140_n N_A_27_47#_M1000_g N_A_27_47#_c_141_n
+ N_A_27_47#_M1005_g N_A_27_47#_c_142_n N_A_27_47#_c_149_n N_A_27_47#_c_143_n
+ N_A_27_47#_c_144_n N_A_27_47#_c_145_n N_A_27_47#_c_152_n N_A_27_47#_c_146_n
+ N_A_27_47#_c_147_n PM_SKY130_FD_SC_HDLL__AND3_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__AND3_1%VPWR N_VPWR_M1002_d N_VPWR_M1004_d N_VPWR_c_214_n
+ VPWR N_VPWR_c_215_n N_VPWR_c_216_n N_VPWR_c_213_n N_VPWR_c_218_n
+ N_VPWR_c_219_n PM_SKY130_FD_SC_HDLL__AND3_1%VPWR
x_PM_SKY130_FD_SC_HDLL__AND3_1%X N_X_M1005_d N_X_M1000_d N_X_c_247_n N_X_c_244_n
+ N_X_c_245_n X X N_X_c_249_n PM_SKY130_FD_SC_HDLL__AND3_1%X
x_PM_SKY130_FD_SC_HDLL__AND3_1%VGND N_VGND_M1003_d N_VGND_c_266_n N_VGND_c_267_n
+ N_VGND_c_268_n VGND N_VGND_c_269_n N_VGND_c_270_n
+ PM_SKY130_FD_SC_HDLL__AND3_1%VGND
cc_1 VNB N_A_c_48_n 0.0741603f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.425
cc_2 VNB N_A_c_49_n 0.0179045f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_3 VNB A 0.0193438f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_4 VNB N_B_M1001_g 0.0425745f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_5 VNB N_B_c_75_n 0.00266648f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=0.93
cc_6 VNB N_C_c_109_n 0.0326198f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.425
cc_7 VNB N_C_M1003_g 0.0278233f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_8 VNB C 0.0110412f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_140_n 0.0258391f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=0.93
cc_10 VNB N_A_27_47#_c_141_n 0.0208424f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_142_n 0.00795526f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_143_n 0.00665611f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_144_n 0.00504859f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_145_n 0.00872518f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_146_n 0.00149979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_147_n 0.00757968f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VPWR_c_213_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_X_c_244_n 0.0254418f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=0.93
cc_19 VNB N_X_c_245_n 0.00494099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB X 0.0136214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_266_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_22 VNB N_VGND_c_267_n 0.0518159f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=0.93
cc_23 VNB N_VGND_c_268_n 0.00324476f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=0.93
cc_24 VNB N_VGND_c_269_n 0.0207186f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_270_n 0.162264f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VPB N_A_c_48_n 0.0314212f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.425
cc_27 VPB N_B_c_76_n 0.0482929f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.71
cc_28 VPB N_B_M1007_g 0.0125327f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_29 VPB N_B_c_75_n 0.00701635f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=0.93
cc_30 VPB B 0.0145583f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_C_c_109_n 0.0279049f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.425
cc_32 VPB N_A_27_47#_c_140_n 0.0312009f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=0.93
cc_33 VPB N_A_27_47#_c_149_n 0.0186616f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_27_47#_c_143_n 0.00395347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_27_47#_c_144_n 0.00224001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_27_47#_c_152_n 0.0119586f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_27_47#_c_146_n 0.0139943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_27_47#_c_147_n 7.01983e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_214_n 0.00253836f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=0.93
cc_40 VPB N_VPWR_c_215_n 0.03159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_216_n 0.0174623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_213_n 0.0560549f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_218_n 0.0614238f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_219_n 0.00378547f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_X_c_247_n 0.00524127f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=0.93
cc_46 VPB N_X_c_244_n 0.018551f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=0.93
cc_47 VPB N_X_c_249_n 0.0218575f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 N_A_c_48_n N_B_c_76_n 0.00308179f $X=0.495 $Y=1.425 $X2=0 $Y2=0
cc_49 N_A_c_48_n N_B_M1007_g 0.0122821f $X=0.495 $Y=1.425 $X2=0 $Y2=0
cc_50 N_A_c_49_n N_B_M1001_g 0.0448847f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_51 A N_B_M1001_g 0.00133945f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_52 N_A_c_48_n N_B_c_75_n 0.0065818f $X=0.495 $Y=1.425 $X2=0 $Y2=0
cc_53 A N_A_27_47#_M1006_s 0.00265319f $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_54 N_A_c_48_n N_A_27_47#_c_142_n 0.00164355f $X=0.495 $Y=1.425 $X2=0 $Y2=0
cc_55 N_A_c_49_n N_A_27_47#_c_142_n 0.00812634f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_56 A N_A_27_47#_c_142_n 0.0349872f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_57 N_A_c_48_n N_A_27_47#_c_149_n 0.00826777f $X=0.495 $Y=1.425 $X2=0 $Y2=0
cc_58 N_A_c_48_n N_A_27_47#_c_143_n 0.0166216f $X=0.495 $Y=1.425 $X2=0 $Y2=0
cc_59 A N_A_27_47#_c_143_n 0.0253131f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_60 N_A_c_48_n N_A_27_47#_c_144_n 0.0104883f $X=0.495 $Y=1.425 $X2=0 $Y2=0
cc_61 A N_A_27_47#_c_144_n 0.0212009f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_62 N_A_c_48_n N_A_27_47#_c_145_n 0.00352274f $X=0.495 $Y=1.425 $X2=0 $Y2=0
cc_63 N_A_c_49_n N_A_27_47#_c_145_n 0.0044106f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_64 A N_A_27_47#_c_145_n 0.0325483f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_65 N_A_c_48_n N_A_27_47#_c_146_n 6.83901e-19 $X=0.495 $Y=1.425 $X2=0 $Y2=0
cc_66 N_A_c_48_n N_VPWR_c_218_n 0.0259744f $X=0.495 $Y=1.425 $X2=0 $Y2=0
cc_67 A A_119_47# 5.13426e-19 $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_68 N_A_c_49_n N_VGND_c_267_n 0.00366111f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_69 N_A_c_49_n N_VGND_c_270_n 0.00638996f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_70 N_B_M1007_g N_C_c_109_n 0.00962644f $X=0.965 $Y=1.71 $X2=-0.19 $Y2=-0.24
cc_71 N_B_M1001_g N_C_c_109_n 0.0112223f $X=0.99 $Y=0.445 $X2=-0.19 $Y2=-0.24
cc_72 N_B_c_75_n N_C_c_109_n 0.00254446f $X=0.97 $Y=1.425 $X2=-0.19 $Y2=-0.24
cc_73 N_B_M1001_g N_C_M1003_g 0.0154098f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_74 N_B_M1001_g C 0.00389195f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_75 B N_A_27_47#_c_140_n 9.58704e-19 $X=1.15 $Y=2.21 $X2=0 $Y2=0
cc_76 N_B_M1001_g N_A_27_47#_c_142_n 0.00750669f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_77 N_B_M1001_g N_A_27_47#_c_145_n 0.0193537f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_78 B N_A_27_47#_c_152_n 0.0048204f $X=1.15 $Y=2.21 $X2=0 $Y2=0
cc_79 N_B_c_76_n N_A_27_47#_c_146_n 5.18249e-19 $X=0.965 $Y=2.05 $X2=0 $Y2=0
cc_80 N_B_M1007_g N_A_27_47#_c_146_n 0.00957724f $X=0.965 $Y=1.71 $X2=0 $Y2=0
cc_81 N_B_M1001_g N_A_27_47#_c_146_n 0.00271577f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_82 N_B_c_75_n N_A_27_47#_c_146_n 0.0075143f $X=0.97 $Y=1.425 $X2=0 $Y2=0
cc_83 B N_A_27_47#_c_146_n 0.0225657f $X=1.15 $Y=2.21 $X2=0 $Y2=0
cc_84 B N_VPWR_c_214_n 0.0150617f $X=1.15 $Y=2.21 $X2=0 $Y2=0
cc_85 N_B_c_76_n N_VPWR_c_215_n 0.00358793f $X=0.965 $Y=2.05 $X2=0 $Y2=0
cc_86 B N_VPWR_c_215_n 0.039241f $X=1.15 $Y=2.21 $X2=0 $Y2=0
cc_87 N_B_c_76_n N_VPWR_c_213_n 0.00175718f $X=0.965 $Y=2.05 $X2=0 $Y2=0
cc_88 B N_VPWR_c_213_n 0.0219398f $X=1.15 $Y=2.21 $X2=0 $Y2=0
cc_89 N_B_c_76_n N_VPWR_c_218_n 0.010808f $X=0.965 $Y=2.05 $X2=0 $Y2=0
cc_90 N_B_M1007_g N_VPWR_c_218_n 0.00771022f $X=0.965 $Y=1.71 $X2=0 $Y2=0
cc_91 B N_VPWR_c_218_n 0.0290712f $X=1.15 $Y=2.21 $X2=0 $Y2=0
cc_92 N_B_M1001_g N_VGND_c_267_n 0.00365909f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_93 N_B_M1001_g N_VGND_c_270_n 0.00599788f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_94 N_C_c_109_n N_A_27_47#_c_140_n 0.0332094f $X=1.65 $Y=1.425 $X2=0 $Y2=0
cc_95 C N_A_27_47#_c_140_n 8.09068e-19 $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_96 N_C_M1003_g N_A_27_47#_c_141_n 0.0162279f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_97 C N_A_27_47#_c_141_n 0.00543816f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_98 N_C_c_109_n N_A_27_47#_c_145_n 9.00145e-19 $X=1.65 $Y=1.425 $X2=0 $Y2=0
cc_99 N_C_M1003_g N_A_27_47#_c_145_n 8.64849e-19 $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_100 C N_A_27_47#_c_145_n 0.0333075f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_101 N_C_c_109_n N_A_27_47#_c_152_n 0.0358638f $X=1.65 $Y=1.425 $X2=0 $Y2=0
cc_102 C N_A_27_47#_c_152_n 0.0289244f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_103 N_C_c_109_n N_A_27_47#_c_146_n 0.00378159f $X=1.65 $Y=1.425 $X2=0 $Y2=0
cc_104 C N_A_27_47#_c_146_n 0.00296658f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_105 N_C_c_109_n N_A_27_47#_c_147_n 0.00410686f $X=1.65 $Y=1.425 $X2=0 $Y2=0
cc_106 C N_A_27_47#_c_147_n 0.0121361f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_107 N_C_c_109_n N_VPWR_c_215_n 0.00400776f $X=1.65 $Y=1.425 $X2=0 $Y2=0
cc_108 N_C_c_109_n N_VPWR_c_213_n 0.00505391f $X=1.65 $Y=1.425 $X2=0 $Y2=0
cc_109 N_C_c_109_n N_VPWR_c_218_n 4.10482e-19 $X=1.65 $Y=1.425 $X2=0 $Y2=0
cc_110 C A_213_47# 0.00633506f $X=1.525 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_111 N_C_M1003_g N_VGND_c_266_n 0.00491616f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_112 N_C_M1003_g N_VGND_c_267_n 0.00367922f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_113 C N_VGND_c_267_n 0.0175747f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_114 N_C_M1003_g N_VGND_c_270_n 0.00627564f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_115 C N_VGND_c_270_n 0.0131109f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_116 N_A_27_47#_c_152_n N_VPWR_M1004_d 0.00602429f $X=2.04 $Y=1.627 $X2=0
+ $Y2=0
cc_117 N_A_27_47#_c_140_n N_VPWR_c_214_n 0.0111557f $X=2.25 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A_27_47#_c_152_n N_VPWR_c_214_n 0.0145116f $X=2.04 $Y=1.627 $X2=0 $Y2=0
cc_119 N_A_27_47#_c_140_n N_VPWR_c_216_n 0.00681171f $X=2.25 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_27_47#_c_140_n N_VPWR_c_213_n 0.0123611f $X=2.25 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_27_47#_c_152_n N_VPWR_c_213_n 0.0164006f $X=2.04 $Y=1.627 $X2=0 $Y2=0
cc_122 N_A_27_47#_c_149_n N_VPWR_c_218_n 0.031387f $X=0.26 $Y=1.645 $X2=0 $Y2=0
cc_123 N_A_27_47#_c_143_n N_VPWR_c_218_n 0.0182938f $X=0.855 $Y=1.275 $X2=0
+ $Y2=0
cc_124 N_A_27_47#_c_146_n N_VPWR_c_218_n 0.0118296f $X=1.417 $Y=1.627 $X2=0
+ $Y2=0
cc_125 N_A_27_47#_c_140_n N_X_c_244_n 0.00705961f $X=2.25 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A_27_47#_c_141_n N_X_c_244_n 0.0186399f $X=2.275 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_27_47#_c_152_n N_X_c_244_n 0.0225924f $X=2.04 $Y=1.627 $X2=0 $Y2=0
cc_128 N_A_27_47#_c_147_n N_X_c_244_n 0.0228547f $X=2.185 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A_27_47#_c_142_n A_119_47# 0.00889314f $X=0.855 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_130 N_A_27_47#_c_145_n A_119_47# 0.00234049f $X=0.965 $Y=1.19 $X2=-0.19
+ $Y2=-0.24
cc_131 N_A_27_47#_c_140_n N_VGND_c_266_n 3.47141e-19 $X=2.25 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A_27_47#_c_141_n N_VGND_c_266_n 0.00471604f $X=2.275 $Y=0.995 $X2=0
+ $Y2=0
cc_133 N_A_27_47#_c_147_n N_VGND_c_266_n 0.00308815f $X=2.185 $Y=1.16 $X2=0
+ $Y2=0
cc_134 N_A_27_47#_c_142_n N_VGND_c_267_n 0.0463657f $X=0.855 $Y=0.38 $X2=0 $Y2=0
cc_135 N_A_27_47#_c_141_n N_VGND_c_269_n 0.00585385f $X=2.275 $Y=0.995 $X2=0
+ $Y2=0
cc_136 N_A_27_47#_M1006_s N_VGND_c_270_n 0.00253093f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_137 N_A_27_47#_c_141_n N_VGND_c_270_n 0.0122398f $X=2.275 $Y=0.995 $X2=0
+ $Y2=0
cc_138 N_A_27_47#_c_142_n N_VGND_c_270_n 0.0348136f $X=0.855 $Y=0.38 $X2=0 $Y2=0
cc_139 N_VPWR_c_213_n N_X_M1000_d 0.00378012f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_140 N_VPWR_c_216_n N_X_c_249_n 0.0188956f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_141 N_VPWR_c_213_n N_X_c_249_n 0.0105168f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_142 X N_VGND_c_269_n 0.0178555f $X=2.43 $Y=0.425 $X2=0 $Y2=0
cc_143 N_X_M1005_d N_VGND_c_270_n 0.00387172f $X=2.35 $Y=0.235 $X2=0 $Y2=0
cc_144 X N_VGND_c_270_n 0.00990557f $X=2.43 $Y=0.425 $X2=0 $Y2=0
cc_145 A_119_47# N_VGND_c_270_n 0.00259819f $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_146 A_213_47# N_VGND_c_270_n 0.0153222f $X=1.065 $Y=0.235 $X2=0 $Y2=0
