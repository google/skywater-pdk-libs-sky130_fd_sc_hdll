* File: sky130_fd_sc_hdll__clkinv_2.pex.spice
* Created: Wed Sep  2 08:26:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKINV_2%A 1 3 4 6 9 11 12 13 15 18 20 21 22 23 41
+ 46
r52 34 35 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.05
+ $Y=1.16 $X2=1.05 $Y2=1.16
r53 32 34 1.46061 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=1.04 $Y=1.212 $X2=1.05
+ $Y2=1.212
r54 31 32 5.84242 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=1 $Y=1.212 $X2=1.04
+ $Y2=1.212
r55 30 31 70.1091 $w=3.3e-07 $l=4.8e-07 $layer=POLY_cond $X=0.52 $Y=1.212 $X2=1
+ $Y2=1.212
r56 29 41 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.32 $Y=1.177
+ $X2=0.69 $Y2=1.177
r57 28 30 29.2121 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.32 $Y=1.212 $X2=0.52
+ $Y2=1.212
r58 28 29 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=1.16 $X2=0.32 $Y2=1.16
r59 23 46 0.256098 $w=2.23e-07 $l=5e-09 $layer=LI1_cond $X=1.145 $Y=1.177
+ $X2=1.15 $Y2=1.177
r60 23 35 4.86587 $w=2.23e-07 $l=9.5e-08 $layer=LI1_cond $X=1.145 $Y=1.177
+ $X2=1.05 $Y2=1.177
r61 22 35 15.8781 $w=2.23e-07 $l=3.1e-07 $layer=LI1_cond $X=0.74 $Y=1.177
+ $X2=1.05 $Y2=1.177
r62 22 41 2.56098 $w=2.23e-07 $l=5e-08 $layer=LI1_cond $X=0.74 $Y=1.177 $X2=0.69
+ $Y2=1.177
r63 21 29 4.60977 $w=2.23e-07 $l=9e-08 $layer=LI1_cond $X=0.23 $Y=1.177 $X2=0.32
+ $Y2=1.177
r64 16 20 30.0832 $w=1.65e-07 $l=2.04118e-07 $layer=POLY_cond $X=1.52 $Y=1.025
+ $X2=1.495 $Y2=1.217
r65 16 18 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.52 $Y=1.025
+ $X2=1.52 $Y2=0.445
r66 13 20 30.0832 $w=1.65e-07 $l=1.93e-07 $layer=POLY_cond $X=1.495 $Y=1.41
+ $X2=1.495 $Y2=1.217
r67 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.495 $Y=1.41
+ $X2=1.495 $Y2=1.985
r68 12 34 11.2297 $w=3.3e-07 $l=8.72066e-08 $layer=POLY_cond $X=1.115 $Y=1.16
+ $X2=1.05 $Y2=1.212
r69 11 20 1.40033 $w=2.7e-07 $l=1.253e-07 $layer=POLY_cond $X=1.395 $Y=1.16
+ $X2=1.495 $Y2=1.217
r70 11 12 62.2086 $w=2.7e-07 $l=2.8e-07 $layer=POLY_cond $X=1.395 $Y=1.16
+ $X2=1.115 $Y2=1.16
r71 7 32 21.2229 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=1.04 $Y=1.015
+ $X2=1.04 $Y2=1.212
r72 7 9 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.04 $Y=1.015 $X2=1.04
+ $Y2=0.445
r73 4 31 16.9318 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=1 $Y=1.41 $X2=1
+ $Y2=1.212
r74 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1 $Y=1.41 $X2=1
+ $Y2=1.985
r75 1 30 16.9318 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=0.52 $Y=1.41
+ $X2=0.52 $Y2=1.212
r76 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.52 $Y=1.41 $X2=0.52
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_2%Y 1 2 3 12 14 15 18 22 24 25 26 32 42
r48 32 42 14.8096 $w=1.68e-07 $l=2.27e-07 $layer=LI1_cond $X=1.837 $Y=0.81
+ $X2=1.61 $Y2=0.81
r49 26 33 2.17804 $w=4.47e-07 $l=2.43824e-07 $layer=LI1_cond $X=1.632 $Y=1.545
+ $X2=1.837 $Y2=1.46
r50 26 33 0.150687 $w=6.33e-07 $l=8e-09 $layer=LI1_cond $X=1.837 $Y=1.452
+ $X2=1.837 $Y2=1.46
r51 25 26 4.935 $w=6.33e-07 $l=2.62e-07 $layer=LI1_cond $X=1.837 $Y=1.19
+ $X2=1.837 $Y2=1.452
r52 24 42 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.605 $Y=0.81
+ $X2=1.61 $Y2=0.81
r53 24 25 5.17987 $w=6.33e-07 $l=2.75e-07 $layer=LI1_cond $X=1.837 $Y=0.915
+ $X2=1.837 $Y2=1.19
r54 24 32 0.376718 $w=6.33e-07 $l=2e-08 $layer=LI1_cond $X=1.837 $Y=0.915
+ $X2=1.837 $Y2=0.895
r55 20 24 24.0086 $w=1.68e-07 $l=3.68e-07 $layer=LI1_cond $X=1.237 $Y=0.81
+ $X2=1.605 $Y2=0.81
r56 20 22 14.3415 $w=2.23e-07 $l=2.8e-07 $layer=LI1_cond $X=1.237 $Y=0.725
+ $X2=1.237 $Y2=0.445
r57 16 26 2.17804 $w=4.47e-07 $l=4.32416e-07 $layer=LI1_cond $X=1.24 $Y=1.63
+ $X2=1.632 $Y2=1.545
r58 16 18 8.86495 $w=2.58e-07 $l=2e-07 $layer=LI1_cond $X=1.24 $Y=1.63 $X2=1.24
+ $Y2=1.83
r59 14 26 4.97337 $w=1.7e-07 $l=5.22e-07 $layer=LI1_cond $X=1.11 $Y=1.545
+ $X2=1.632 $Y2=1.545
r60 14 15 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.11 $Y=1.545 $X2=0.41
+ $Y2=1.545
r61 10 15 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.282 $Y=1.63
+ $X2=0.41 $Y2=1.545
r62 10 12 9.03877 $w=2.53e-07 $l=2e-07 $layer=LI1_cond $X=0.282 $Y=1.63
+ $X2=0.282 $Y2=1.83
r63 3 18 300 $w=1.7e-07 $l=4.13249e-07 $layer=licon1_PDIFF $count=2 $X=1.09
+ $Y=1.485 $X2=1.24 $Y2=1.83
r64 2 12 300 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=2 $X=0.155
+ $Y=1.485 $X2=0.28 $Y2=1.83
r65 1 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.115
+ $Y=0.235 $X2=1.255 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_2%VPWR 1 2 11 13 17 19 23 24 27 30
r27 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r28 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r29 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r30 24 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r31 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r32 21 30 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.86 $Y=2.72
+ $X2=1.732 $Y2=2.72
r33 21 23 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.86 $Y=2.72
+ $X2=2.07 $Y2=2.72
r34 19 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r35 15 30 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.732 $Y=2.635
+ $X2=1.732 $Y2=2.72
r36 15 17 30.2799 $w=2.53e-07 $l=6.7e-07 $layer=LI1_cond $X=1.732 $Y=2.635
+ $X2=1.732 $Y2=1.965
r37 14 27 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.89 $Y=2.72 $X2=0.76
+ $Y2=2.72
r38 13 30 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=1.732 $Y2=2.72
r39 13 14 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=0.89 $Y2=2.72
r40 9 27 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=2.635
+ $X2=0.76 $Y2=2.72
r41 9 11 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=0.76 $Y=2.635
+ $X2=0.76 $Y2=1.965
r42 2 17 300 $w=1.7e-07 $l=5.49909e-07 $layer=licon1_PDIFF $count=2 $X=1.585
+ $Y=1.485 $X2=1.735 $Y2=1.965
r43 1 11 300 $w=1.7e-07 $l=5.49909e-07 $layer=licon1_PDIFF $count=2 $X=0.61
+ $Y=1.485 $X2=0.76 $Y2=1.965
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_2%VGND 1 2 9 13 15 17 22 29 30 33 36
r25 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r26 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r27 30 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r28 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r29 27 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.9 $Y=0 $X2=1.71
+ $Y2=0
r30 27 29 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.9 $Y=0 $X2=2.07
+ $Y2=0
r31 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r32 26 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r33 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r34 23 33 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.732
+ $Y2=0
r35 23 25 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.15
+ $Y2=0
r36 22 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.52 $Y=0 $X2=1.71
+ $Y2=0
r37 22 25 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.52 $Y=0 $X2=1.15
+ $Y2=0
r38 17 33 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.732
+ $Y2=0
r39 17 19 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.23
+ $Y2=0
r40 15 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r41 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r42 11 36 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0
r43 11 13 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0.39
r44 7 33 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=0.732 $Y=0.085
+ $X2=0.732 $Y2=0
r45 7 9 12.0255 $w=3.43e-07 $l=3.6e-07 $layer=LI1_cond $X=0.732 $Y=0.085
+ $X2=0.732 $Y2=0.445
r46 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.73 $Y2=0.39
r47 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.65
+ $Y=0.235 $X2=0.775 $Y2=0.445
.ends

