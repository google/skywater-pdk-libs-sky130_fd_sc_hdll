* NGSPICE file created from sky130_fd_sc_hdll__a211oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.99e+12p pd=1.798e+07u as=1.16e+12p ps=1.032e+07u
M1001 VGND C1 Y VNB nshort w=650000u l=150000u
+  ad=1.404e+12p pd=1.342e+07u as=1.365e+12p ps=1.2e+07u
M1002 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND A2 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.995e+11p ps=7.66e+06u
M1004 Y C1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_869_297# C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=6.2e+11p ps=5.24e+06u
M1007 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1057_297# B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.2e+11p pd=2.64e+06u as=0p ps=0u
M1010 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A2 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_119_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND C1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y C1 a_1057_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_297# B1 a_869_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y C1 a_869_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_119_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y C1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_869_297# B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y A1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1449_297# C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=3.3e+11p pd=2.66e+06u as=0p ps=0u
M1027 a_27_297# B1 a_1449_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_119_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y A1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_119_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

