* File: sky130_fd_sc_hdll__buf_1.spice
* Created: Wed Sep  2 08:24:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__buf_1.pex.spice"
.subckt sky130_fd_sc_hdll__buf_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_27_47#_M1002_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0884 AS=0.1612 PD=0.86 PS=1.66 NRD=0 NRS=10.38 M=1 R=3.46667 SA=75000.2
+ SB=75000.7 A=0.078 P=1.34 MULT=1
MM1003 N_X_M1003_d N_A_27_47#_M1003_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0884 PD=1.56 PS=0.86 NRD=0 NRS=14.988 M=1 R=3.46667 SA=75000.7
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_27_47#_M1000_s VPB PHIGHVT L=0.18 W=0.79
+ AD=0.12245 AS=0.2133 PD=1.1 PS=2.12 NRD=1.2411 NRS=1.2411 M=1 R=4.38889
+ SA=90000.2 SB=90000.7 A=0.1422 P=1.94 MULT=1
MM1001 N_X_M1001_d N_A_27_47#_M1001_g N_VPWR_M1000_d VPB PHIGHVT L=0.18 W=0.79
+ AD=0.2133 AS=0.12245 PD=2.12 PS=1.1 NRD=1.2411 NRS=6.2252 M=1 R=4.38889
+ SA=90000.7 SB=90000.2 A=0.1422 P=1.94 MULT=1
DX4_noxref VNB VPB NWDIODE A=3.5631 P=7.65
pX5_noxref noxref_8 X X PROBETYPE=1
pX6_noxref noxref_9 X X PROBETYPE=1
pX7_noxref noxref_10 X X PROBETYPE=1
*
.include "sky130_fd_sc_hdll__buf_1.pxi.spice"
*
.ends
*
*
