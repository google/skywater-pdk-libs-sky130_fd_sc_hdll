* File: sky130_fd_sc_hdll__a2bb2oi_2.spice
* Created: Wed Sep  2 08:19:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a2bb2oi_2.pex.spice"
.subckt sky130_fd_sc_hdll__a2bb2oi_2  VNB VPB B1 B2 A1_N A2_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2_N	A2_N
* A1_N	A1_N
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1010 N_A_119_47#_M1010_d N_B1_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75005 A=0.0975 P=1.6 MULT=1
MM1003 N_Y_M1003_d N_B2_M1003_g N_A_119_47#_M1010_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1019 N_Y_M1003_d N_B2_M1019_g N_A_119_47#_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75004 A=0.0975 P=1.6 MULT=1
MM1011 N_A_119_47#_M1019_s N_B1_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1011_s N_A_455_21#_M1014_g N_Y_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.1
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1015_d N_A_455_21#_M1015_g N_Y_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.273 AS=0.104 PD=1.49 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.5
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1004 N_A_455_21#_M1004_d N_A1_N_M1004_g N_VGND_M1015_d VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.273 PD=1.02 PS=1.49 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75003.5 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1013 N_A_455_21#_M1004_d N_A1_N_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75004 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1013_s N_A2_N_M1006_g N_A_455_21#_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75004.5 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1017_d N_A2_N_M1017_g N_A_455_21#_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.182 AS=0.12025 PD=1.86 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75005 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_B1_M1005_g N_A_27_297#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1000 N_A_27_297#_M1000_d N_B2_M1000_g N_VPWR_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1016 N_A_27_297#_M1000_d N_B2_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1016_s N_B1_M1009_g N_A_27_297#_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1002 N_A_27_297#_M1009_s N_A_455_21#_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1007 N_A_27_297#_M1007_d N_A_455_21#_M1007_g N_Y_M1002_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1012 N_A_695_297#_M1012_d N_A1_N_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1018 N_A_695_297#_M1018_d N_A1_N_M1018_g N_VPWR_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1001 N_A_695_297#_M1018_d N_A2_N_M1001_g N_A_455_21#_M1001_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1008 N_A_695_297#_M1008_d N_A2_N_M1008_g N_A_455_21#_M1001_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.29 AS=0.145 PD=2.58 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.4245 P=16.2
pX21_noxref noxref_14 A1_N A1_N PROBETYPE=1
*
.include "sky130_fd_sc_hdll__a2bb2oi_2.pxi.spice"
*
.ends
*
*
