* File: sky130_fd_sc_hdll__einvp_8.pex.spice
* Created: Thu Aug 27 19:08:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__EINVP_8%TE 1 3 4 6 7 9 11 12 14 16 17 19 21 22 24
+ 26 27 29 31 32 34 36 37 39 41 42 44 46 47 48 49 50 51 52 53 54 55
c139 53 0 1.15978e-19 $X=3.78 $Y=1.035
c140 52 0 1.15978e-19 $X=3.31 $Y=1.035
c141 51 0 1.15978e-19 $X=2.84 $Y=1.035
c142 50 0 1.15978e-19 $X=2.37 $Y=1.035
c143 49 0 1.15978e-19 $X=1.9 $Y=1.035
c144 48 0 1.15616e-19 $X=1.48 $Y=1.035
c145 42 0 6.61776e-19 $X=4.225 $Y=1.035
c146 32 0 3.93344e-19 $X=3.235 $Y=1.035
c147 22 0 3.93344e-19 $X=2.295 $Y=1.035
c148 12 0 1.96687e-19 $X=1.405 $Y=1.035
r149 58 60 14.7311 $w=4.09e-07 $l=1.25e-07 $layer=POLY_cond $X=0.352 $Y=1.035
+ $X2=0.352 $Y2=1.16
r150 54 55 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.207 $Y=1.16
+ $X2=0.207 $Y2=1.53
r151 54 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r152 44 46 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.3 $Y=0.96 $X2=4.3
+ $Y2=0.56
r153 43 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.855 $Y=1.035
+ $X2=3.78 $Y2=1.035
r154 42 44 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.225 $Y=1.035
+ $X2=4.3 $Y2=0.96
r155 42 43 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.225 $Y=1.035
+ $X2=3.855 $Y2=1.035
r156 39 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.78 $Y=0.96
+ $X2=3.78 $Y2=1.035
r157 39 41 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.78 $Y=0.96 $X2=3.78
+ $Y2=0.56
r158 38 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.385 $Y=1.035
+ $X2=3.31 $Y2=1.035
r159 37 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.705 $Y=1.035
+ $X2=3.78 $Y2=1.035
r160 37 38 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.705 $Y=1.035
+ $X2=3.385 $Y2=1.035
r161 34 52 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.31 $Y=0.96
+ $X2=3.31 $Y2=1.035
r162 34 36 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.31 $Y=0.96 $X2=3.31
+ $Y2=0.56
r163 33 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.915 $Y=1.035
+ $X2=2.84 $Y2=1.035
r164 32 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.235 $Y=1.035
+ $X2=3.31 $Y2=1.035
r165 32 33 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.235 $Y=1.035
+ $X2=2.915 $Y2=1.035
r166 29 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.84 $Y=0.96
+ $X2=2.84 $Y2=1.035
r167 29 31 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.84 $Y=0.96 $X2=2.84
+ $Y2=0.56
r168 28 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.445 $Y=1.035
+ $X2=2.37 $Y2=1.035
r169 27 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.765 $Y=1.035
+ $X2=2.84 $Y2=1.035
r170 27 28 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.765 $Y=1.035
+ $X2=2.445 $Y2=1.035
r171 24 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.37 $Y=0.96
+ $X2=2.37 $Y2=1.035
r172 24 26 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.37 $Y=0.96 $X2=2.37
+ $Y2=0.56
r173 23 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.975 $Y=1.035
+ $X2=1.9 $Y2=1.035
r174 22 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.295 $Y=1.035
+ $X2=2.37 $Y2=1.035
r175 22 23 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.295 $Y=1.035
+ $X2=1.975 $Y2=1.035
r176 19 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.9 $Y=0.96 $X2=1.9
+ $Y2=1.035
r177 19 21 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.9 $Y=0.96 $X2=1.9
+ $Y2=0.56
r178 18 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.555 $Y=1.035
+ $X2=1.48 $Y2=1.035
r179 17 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.825 $Y=1.035
+ $X2=1.9 $Y2=1.035
r180 17 18 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.825 $Y=1.035
+ $X2=1.555 $Y2=1.035
r181 14 48 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.48 $Y=0.96
+ $X2=1.48 $Y2=1.035
r182 14 16 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.48 $Y=0.96 $X2=1.48
+ $Y2=0.56
r183 13 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.065 $Y=1.035
+ $X2=0.99 $Y2=1.035
r184 12 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.405 $Y=1.035
+ $X2=1.48 $Y2=1.035
r185 12 13 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.405 $Y=1.035
+ $X2=1.065 $Y2=1.035
r186 9 47 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.99 $Y=0.96
+ $X2=0.99 $Y2=1.035
r187 9 11 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.99 $Y=0.96 $X2=0.99
+ $Y2=0.56
r188 8 58 26.4068 $w=1.5e-07 $l=2.43e-07 $layer=POLY_cond $X=0.595 $Y=1.035
+ $X2=0.352 $Y2=1.035
r189 7 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.915 $Y=1.035
+ $X2=0.99 $Y2=1.035
r190 7 8 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.915 $Y=1.035
+ $X2=0.595 $Y2=1.035
r191 4 60 44.8154 $w=4.09e-07 $l=3.13449e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.352 $Y2=1.16
r192 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r193 1 58 29.1598 $w=4.09e-07 $l=1.50911e-07 $layer=POLY_cond $X=0.47 $Y=0.96
+ $X2=0.352 $Y2=1.035
r194 1 3 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.47 $Y=0.96 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_8%A_27_47# 1 2 7 9 10 11 12 14 15 17 19 20
+ 22 24 25 27 29 30 32 34 35 37 39 40 42 44 45 46 47 48 49 50 52 55 59 61 62 64
+ 67 68 78
c177 78 0 1.9418e-19 $X=0.712 $Y=1.16
c178 52 0 1.46731e-19 $X=4.765 $Y=1.395
c179 49 0 6.62625e-20 $X=3.885 $Y=1.395
c180 48 0 1.65302e-19 $X=3.415 $Y=1.395
c181 47 0 1.64162e-19 $X=2.945 $Y=1.395
c182 46 0 1.65302e-19 $X=2.475 $Y=1.395
c183 45 0 1.64162e-19 $X=2.005 $Y=1.395
c184 42 0 1.79447e-19 $X=4.825 $Y=1.47
c185 35 0 1.40591e-19 $X=4.265 $Y=1.395
c186 30 0 7.37964e-20 $X=3.795 $Y=1.395
c187 25 0 7.37964e-20 $X=3.325 $Y=1.395
c188 20 0 7.37964e-20 $X=2.855 $Y=1.395
c189 15 0 7.37964e-20 $X=2.385 $Y=1.395
c190 10 0 7.37964e-20 $X=1.915 $Y=1.395
r191 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.74
+ $Y=1.16 $X2=4.74 $Y2=1.16
r192 65 78 1.39677 $w=3.3e-07 $l=2.13e-07 $layer=LI1_cond $X=0.925 $Y=1.16
+ $X2=0.712 $Y2=1.16
r193 65 67 133.229 $w=3.28e-07 $l=3.815e-06 $layer=LI1_cond $X=0.925 $Y=1.16
+ $X2=4.74 $Y2=1.16
r194 63 78 5.10169 $w=3.35e-07 $l=1.65e-07 $layer=LI1_cond $X=0.712 $Y=1.325
+ $X2=0.712 $Y2=1.16
r195 63 64 12.4735 $w=4.23e-07 $l=4.6e-07 $layer=LI1_cond $X=0.712 $Y=1.325
+ $X2=0.712 $Y2=1.785
r196 62 78 5.10169 $w=3.35e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.622 $Y=0.995
+ $X2=0.712 $Y2=1.16
r197 61 62 7.99654 $w=2.43e-07 $l=1.7e-07 $layer=LI1_cond $X=0.622 $Y=0.825
+ $X2=0.622 $Y2=0.995
r198 57 64 32.4246 $w=1.68e-07 $l=4.97e-07 $layer=LI1_cond $X=0.215 $Y=1.87
+ $X2=0.712 $Y2=1.87
r199 57 59 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=1.955
+ $X2=0.215 $Y2=2.165
r200 53 61 26.5529 $w=1.68e-07 $l=4.07e-07 $layer=LI1_cond $X=0.215 $Y=0.74
+ $X2=0.622 $Y2=0.74
r201 53 55 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.215 $Y2=0.445
r202 51 68 28.8521 $w=3.2e-07 $l=1.6e-07 $layer=POLY_cond $X=4.765 $Y=1.32
+ $X2=4.765 $Y2=1.16
r203 51 52 13.0992 $w=2.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.765 $Y=1.32
+ $X2=4.765 $Y2=1.395
r204 42 52 13.0992 $w=2.5e-07 $l=1.00623e-07 $layer=POLY_cond $X=4.825 $Y=1.47
+ $X2=4.765 $Y2=1.395
r205 42 44 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=4.825 $Y=1.47
+ $X2=4.825 $Y2=2.015
r206 41 50 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.445 $Y=1.395
+ $X2=4.355 $Y2=1.395
r207 40 52 12.7694 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=4.605 $Y=1.395
+ $X2=4.765 $Y2=1.395
r208 40 41 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=4.605 $Y=1.395
+ $X2=4.445 $Y2=1.395
r209 37 50 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.355 $Y=1.47
+ $X2=4.355 $Y2=1.395
r210 37 39 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=4.355 $Y=1.47
+ $X2=4.355 $Y2=2.015
r211 36 49 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.975 $Y=1.395
+ $X2=3.885 $Y2=1.395
r212 35 50 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.265 $Y=1.395
+ $X2=4.355 $Y2=1.395
r213 35 36 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.265 $Y=1.395
+ $X2=3.975 $Y2=1.395
r214 32 49 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.885 $Y=1.47
+ $X2=3.885 $Y2=1.395
r215 32 34 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=3.885 $Y=1.47
+ $X2=3.885 $Y2=2.015
r216 31 48 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.505 $Y=1.395
+ $X2=3.415 $Y2=1.395
r217 30 49 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.795 $Y=1.395
+ $X2=3.885 $Y2=1.395
r218 30 31 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.795 $Y=1.395
+ $X2=3.505 $Y2=1.395
r219 27 48 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.415 $Y=1.47
+ $X2=3.415 $Y2=1.395
r220 27 29 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=3.415 $Y=1.47
+ $X2=3.415 $Y2=2.015
r221 26 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.035 $Y=1.395
+ $X2=2.945 $Y2=1.395
r222 25 48 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.325 $Y=1.395
+ $X2=3.415 $Y2=1.395
r223 25 26 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.325 $Y=1.395
+ $X2=3.035 $Y2=1.395
r224 22 47 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.945 $Y=1.47
+ $X2=2.945 $Y2=1.395
r225 22 24 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.945 $Y=1.47
+ $X2=2.945 $Y2=2.015
r226 21 46 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.565 $Y=1.395
+ $X2=2.475 $Y2=1.395
r227 20 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.855 $Y=1.395
+ $X2=2.945 $Y2=1.395
r228 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.855 $Y=1.395
+ $X2=2.565 $Y2=1.395
r229 17 46 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.475 $Y=1.47
+ $X2=2.475 $Y2=1.395
r230 17 19 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.475 $Y=1.47
+ $X2=2.475 $Y2=2.015
r231 16 45 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.095 $Y=1.395
+ $X2=2.005 $Y2=1.395
r232 15 46 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.385 $Y=1.395
+ $X2=2.475 $Y2=1.395
r233 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.385 $Y=1.395
+ $X2=2.095 $Y2=1.395
r234 12 45 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.005 $Y=1.47
+ $X2=2.005 $Y2=1.395
r235 12 14 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.005 $Y=1.47
+ $X2=2.005 $Y2=2.015
r236 10 45 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.915 $Y=1.395
+ $X2=2.005 $Y2=1.395
r237 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.915 $Y=1.395
+ $X2=1.625 $Y2=1.395
r238 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.535 $Y=1.47
+ $X2=1.625 $Y2=1.395
r239 7 9 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=1.535 $Y=1.47
+ $X2=1.535 $Y2=2.015
r240 2 59 600 $w=1.7e-07 $l=7.39865e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.165
r241 1 55 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_8%A 1 3 4 6 7 9 10 12 15 17 19 22 24 26 27
+ 29 30 32 33 35 36 38 41 43 45 48 50 52 53 54 55 56 57 58 59 100 107 111 115
+ 118 121 126
c136 17 0 1.69667e-19 $X=6.29 $Y=1.41
r137 100 102 32.4701 $w=3.34e-07 $l=2.25e-07 $layer=POLY_cond $X=8.64 $Y=1.202
+ $X2=8.865 $Y2=1.202
r138 99 100 3.60778 $w=3.34e-07 $l=2.5e-08 $layer=POLY_cond $X=8.615 $Y=1.202
+ $X2=8.64 $Y2=1.202
r139 97 99 20.2036 $w=3.34e-07 $l=1.4e-07 $layer=POLY_cond $X=8.475 $Y=1.202
+ $X2=8.615 $Y2=1.202
r140 95 97 44.015 $w=3.34e-07 $l=3.05e-07 $layer=POLY_cond $X=8.17 $Y=1.202
+ $X2=8.475 $Y2=1.202
r141 94 95 3.60778 $w=3.34e-07 $l=2.5e-08 $layer=POLY_cond $X=8.145 $Y=1.202
+ $X2=8.17 $Y2=1.202
r142 92 94 8.65868 $w=3.34e-07 $l=6e-08 $layer=POLY_cond $X=8.085 $Y=1.202
+ $X2=8.145 $Y2=1.202
r143 92 121 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.085
+ $Y=1.16 $X2=8.085 $Y2=1.16
r144 90 92 55.5599 $w=3.34e-07 $l=3.85e-07 $layer=POLY_cond $X=7.7 $Y=1.202
+ $X2=8.085 $Y2=1.202
r145 88 90 0.721557 $w=3.34e-07 $l=5e-09 $layer=POLY_cond $X=7.695 $Y=1.202
+ $X2=7.7 $Y2=1.202
r146 88 118 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.695
+ $Y=1.16 $X2=7.695 $Y2=1.16
r147 86 88 2.88623 $w=3.34e-07 $l=2e-08 $layer=POLY_cond $X=7.675 $Y=1.202
+ $X2=7.695 $Y2=1.202
r148 85 86 64.2186 $w=3.34e-07 $l=4.45e-07 $layer=POLY_cond $X=7.23 $Y=1.202
+ $X2=7.675 $Y2=1.202
r149 84 85 3.60778 $w=3.34e-07 $l=2.5e-08 $layer=POLY_cond $X=7.205 $Y=1.202
+ $X2=7.23 $Y2=1.202
r150 83 111 12.2023 $w=2.53e-07 $l=2.7e-07 $layer=LI1_cond $X=6.965 $Y=1.147
+ $X2=6.695 $Y2=1.147
r151 82 84 34.6347 $w=3.34e-07 $l=2.4e-07 $layer=POLY_cond $X=6.965 $Y=1.202
+ $X2=7.205 $Y2=1.202
r152 82 83 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.965
+ $Y=1.16 $X2=6.965 $Y2=1.16
r153 80 82 29.5838 $w=3.34e-07 $l=2.05e-07 $layer=POLY_cond $X=6.76 $Y=1.202
+ $X2=6.965 $Y2=1.202
r154 79 80 3.60778 $w=3.34e-07 $l=2.5e-08 $layer=POLY_cond $X=6.735 $Y=1.202
+ $X2=6.76 $Y2=1.202
r155 78 107 15.3659 $w=2.53e-07 $l=3.4e-07 $layer=LI1_cond $X=6.575 $Y=1.147
+ $X2=6.235 $Y2=1.147
r156 77 79 23.0898 $w=3.34e-07 $l=1.6e-07 $layer=POLY_cond $X=6.575 $Y=1.202
+ $X2=6.735 $Y2=1.202
r157 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.575
+ $Y=1.16 $X2=6.575 $Y2=1.16
r158 75 77 41.1287 $w=3.34e-07 $l=2.85e-07 $layer=POLY_cond $X=6.29 $Y=1.202
+ $X2=6.575 $Y2=1.202
r159 74 75 3.60778 $w=3.34e-07 $l=2.5e-08 $layer=POLY_cond $X=6.265 $Y=1.202
+ $X2=6.29 $Y2=1.202
r160 72 74 11.5449 $w=3.34e-07 $l=8e-08 $layer=POLY_cond $X=6.185 $Y=1.202
+ $X2=6.265 $Y2=1.202
r161 70 72 52.6737 $w=3.34e-07 $l=3.65e-07 $layer=POLY_cond $X=5.82 $Y=1.202
+ $X2=6.185 $Y2=1.202
r162 69 70 3.60778 $w=3.34e-07 $l=2.5e-08 $layer=POLY_cond $X=5.795 $Y=1.202
+ $X2=5.82 $Y2=1.202
r163 68 69 64.2186 $w=3.34e-07 $l=4.45e-07 $layer=POLY_cond $X=5.35 $Y=1.202
+ $X2=5.795 $Y2=1.202
r164 67 68 3.60778 $w=3.34e-07 $l=2.5e-08 $layer=POLY_cond $X=5.325 $Y=1.202
+ $X2=5.35 $Y2=1.202
r165 59 126 3.38954 $w=2.53e-07 $l=7.5e-08 $layer=LI1_cond $X=8.865 $Y=1.147
+ $X2=8.94 $Y2=1.147
r166 59 102 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.865
+ $Y=1.16 $X2=8.865 $Y2=1.16
r167 58 59 17.6256 $w=2.53e-07 $l=3.9e-07 $layer=LI1_cond $X=8.475 $Y=1.147
+ $X2=8.865 $Y2=1.147
r168 58 121 18.0775 $w=2.53e-07 $l=4e-07 $layer=LI1_cond $X=8.475 $Y=1.147
+ $X2=8.075 $Y2=1.147
r169 58 97 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.475
+ $Y=1.16 $X2=8.475 $Y2=1.16
r170 57 121 0.677908 $w=2.53e-07 $l=1.5e-08 $layer=LI1_cond $X=8.06 $Y=1.147
+ $X2=8.075 $Y2=1.147
r171 57 118 20.1113 $w=2.53e-07 $l=4.45e-07 $layer=LI1_cond $X=8.06 $Y=1.147
+ $X2=7.615 $Y2=1.147
r172 56 118 0.451938 $w=2.53e-07 $l=1e-08 $layer=LI1_cond $X=7.605 $Y=1.147
+ $X2=7.615 $Y2=1.147
r173 56 115 20.3372 $w=2.53e-07 $l=4.5e-07 $layer=LI1_cond $X=7.605 $Y=1.147
+ $X2=7.155 $Y2=1.147
r174 55 115 1.58178 $w=2.53e-07 $l=3.5e-08 $layer=LI1_cond $X=7.12 $Y=1.147
+ $X2=7.155 $Y2=1.147
r175 55 83 7.00505 $w=2.53e-07 $l=1.55e-07 $layer=LI1_cond $X=7.12 $Y=1.147
+ $X2=6.965 $Y2=1.147
r176 54 111 1.12985 $w=2.53e-07 $l=2.5e-08 $layer=LI1_cond $X=6.67 $Y=1.147
+ $X2=6.695 $Y2=1.147
r177 54 78 4.29342 $w=2.53e-07 $l=9.5e-08 $layer=LI1_cond $X=6.67 $Y=1.147
+ $X2=6.575 $Y2=1.147
r178 53 107 2.25969 $w=2.53e-07 $l=5e-08 $layer=LI1_cond $X=6.185 $Y=1.147
+ $X2=6.235 $Y2=1.147
r179 53 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.185
+ $Y=1.16 $X2=6.185 $Y2=1.16
r180 50 100 17.2128 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.64 $Y=1.41
+ $X2=8.64 $Y2=1.202
r181 50 52 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.64 $Y=1.41
+ $X2=8.64 $Y2=1.985
r182 46 99 21.5099 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=8.615 $Y=1.015
+ $X2=8.615 $Y2=1.202
r183 46 48 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=8.615 $Y=1.015
+ $X2=8.615 $Y2=0.56
r184 43 95 17.2128 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.17 $Y=1.41
+ $X2=8.17 $Y2=1.202
r185 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.17 $Y=1.41
+ $X2=8.17 $Y2=1.985
r186 39 94 21.5099 $w=1.5e-07 $l=1.77e-07 $layer=POLY_cond $X=8.145 $Y=1.025
+ $X2=8.145 $Y2=1.202
r187 39 41 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.145 $Y=1.025
+ $X2=8.145 $Y2=0.56
r188 36 90 17.2128 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.7 $Y=1.41
+ $X2=7.7 $Y2=1.202
r189 36 38 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.7 $Y=1.41
+ $X2=7.7 $Y2=1.985
r190 33 86 21.5099 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.675 $Y=0.995
+ $X2=7.675 $Y2=1.202
r191 33 35 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.675 $Y=0.995
+ $X2=7.675 $Y2=0.56
r192 30 85 17.2128 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.23 $Y=1.41
+ $X2=7.23 $Y2=1.202
r193 30 32 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.23 $Y=1.41
+ $X2=7.23 $Y2=1.985
r194 27 84 21.5099 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.205 $Y=0.995
+ $X2=7.205 $Y2=1.202
r195 27 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.205 $Y=0.995
+ $X2=7.205 $Y2=0.56
r196 24 80 17.2128 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.76 $Y=1.41
+ $X2=6.76 $Y2=1.202
r197 24 26 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.76 $Y=1.41
+ $X2=6.76 $Y2=1.985
r198 20 79 21.5099 $w=1.5e-07 $l=1.77e-07 $layer=POLY_cond $X=6.735 $Y=1.025
+ $X2=6.735 $Y2=1.202
r199 20 22 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.735 $Y=1.025
+ $X2=6.735 $Y2=0.56
r200 17 75 17.2128 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.29 $Y=1.41
+ $X2=6.29 $Y2=1.202
r201 17 19 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.29 $Y=1.41
+ $X2=6.29 $Y2=1.985
r202 13 74 21.5099 $w=1.5e-07 $l=1.77e-07 $layer=POLY_cond $X=6.265 $Y=1.025
+ $X2=6.265 $Y2=1.202
r203 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.265 $Y=1.025
+ $X2=6.265 $Y2=0.56
r204 10 70 17.2128 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.82 $Y=1.41
+ $X2=5.82 $Y2=1.202
r205 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.82 $Y=1.41
+ $X2=5.82 $Y2=1.985
r206 7 69 21.5099 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.795 $Y=0.995
+ $X2=5.795 $Y2=1.202
r207 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.795 $Y=0.995
+ $X2=5.795 $Y2=0.56
r208 4 68 17.2128 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.35 $Y=1.41
+ $X2=5.35 $Y2=1.202
r209 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.35 $Y=1.41
+ $X2=5.35 $Y2=1.985
r210 1 67 21.5099 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.325 $Y=0.995
+ $X2=5.325 $Y2=1.202
r211 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.325 $Y=0.995
+ $X2=5.325 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_8%VPWR 1 2 3 4 5 18 20 24 28 32 36 39 40 42
+ 43 45 46 47 49 68 69 72 75
r131 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r132 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r133 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r134 68 69 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r135 66 69 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=8.97 $Y2=2.72
r136 65 68 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=8.97 $Y2=2.72
r137 65 66 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r138 63 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r139 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r140 60 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r141 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r142 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r143 57 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r144 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r145 54 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=2.72
+ $X2=1.77 $Y2=2.72
r146 54 56 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=1.935 $Y=2.72
+ $X2=2.53 $Y2=2.72
r147 49 72 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.72 $Y2=2.72
r148 49 51 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r149 47 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r150 47 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r151 45 62 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.425 $Y=2.72
+ $X2=4.37 $Y2=2.72
r152 45 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=2.72
+ $X2=4.59 $Y2=2.72
r153 44 65 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.755 $Y=2.72
+ $X2=4.83 $Y2=2.72
r154 44 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.755 $Y=2.72
+ $X2=4.59 $Y2=2.72
r155 42 59 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.485 $Y=2.72
+ $X2=3.45 $Y2=2.72
r156 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.485 $Y=2.72
+ $X2=3.65 $Y2=2.72
r157 41 62 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.815 $Y=2.72
+ $X2=4.37 $Y2=2.72
r158 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.815 $Y=2.72
+ $X2=3.65 $Y2=2.72
r159 39 56 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.53 $Y2=2.72
r160 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.71 $Y2=2.72
r161 38 59 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.875 $Y=2.72
+ $X2=3.45 $Y2=2.72
r162 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=2.72
+ $X2=2.71 $Y2=2.72
r163 34 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.59 $Y=2.635
+ $X2=4.59 $Y2=2.72
r164 34 36 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=4.59 $Y=2.635
+ $X2=4.59 $Y2=2.02
r165 30 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.65 $Y=2.635
+ $X2=3.65 $Y2=2.72
r166 30 32 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=3.65 $Y=2.635
+ $X2=3.65 $Y2=2.02
r167 26 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=2.635
+ $X2=2.71 $Y2=2.72
r168 26 28 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.71 $Y=2.635
+ $X2=2.71 $Y2=2.02
r169 22 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.77 $Y=2.635
+ $X2=1.77 $Y2=2.72
r170 22 24 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.77 $Y=2.635
+ $X2=1.77 $Y2=2.02
r171 21 72 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=0.72 $Y2=2.72
r172 20 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=1.77 $Y2=2.72
r173 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=0.925 $Y2=2.72
r174 16 72 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=2.635
+ $X2=0.72 $Y2=2.72
r175 16 18 8.29197 $w=4.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.72 $Y=2.635
+ $X2=0.72 $Y2=2.34
r176 5 36 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.445
+ $Y=1.545 $X2=4.59 $Y2=2.02
r177 4 32 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.505
+ $Y=1.545 $X2=3.65 $Y2=2.02
r178 3 28 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.565
+ $Y=1.545 $X2=2.71 $Y2=2.02
r179 2 24 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.625
+ $Y=1.545 $X2=1.77 $Y2=2.02
r180 1 18 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_8%A_235_309# 1 2 3 4 5 6 7 8 9 30 32 33 36
+ 38 42 44 48 50 55 56 57 60 62 66 68 72 74 76 79 80 81 82 83 84
c132 81 0 1.97563e-19 $X=4.12 $Y=1.64
c133 80 0 1.96656e-19 $X=3.18 $Y=1.64
c134 79 0 1.96656e-19 $X=2.24 $Y=1.64
c135 50 0 7.0838e-20 $X=4.975 $Y=1.64
c136 44 0 2.31955e-19 $X=4.035 $Y=1.64
c137 38 0 2.31955e-19 $X=3.095 $Y=1.64
c138 32 0 2.31593e-19 $X=2.155 $Y=1.64
r139 76 78 13.4 $w=3.05e-07 $l=3.35e-07 $layer=LI1_cond $X=8.942 $Y=2.295
+ $X2=8.942 $Y2=1.96
r140 75 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.02 $Y=2.38
+ $X2=7.935 $Y2=2.38
r141 74 76 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=8.79 $Y=2.38
+ $X2=8.942 $Y2=2.295
r142 74 75 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=8.79 $Y=2.38
+ $X2=8.02 $Y2=2.38
r143 70 84 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.935 $Y=2.295
+ $X2=7.935 $Y2=2.38
r144 70 72 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.935 $Y=2.295
+ $X2=7.935 $Y2=1.96
r145 69 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.08 $Y=2.38
+ $X2=6.995 $Y2=2.38
r146 68 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.85 $Y=2.38
+ $X2=7.935 $Y2=2.38
r147 68 69 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=7.85 $Y=2.38
+ $X2=7.08 $Y2=2.38
r148 64 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.995 $Y=2.295
+ $X2=6.995 $Y2=2.38
r149 64 66 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.995 $Y=2.295
+ $X2=6.995 $Y2=1.96
r150 63 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.14 $Y=2.38
+ $X2=6.055 $Y2=2.38
r151 62 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.91 $Y=2.38
+ $X2=6.995 $Y2=2.38
r152 62 63 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=6.91 $Y=2.38
+ $X2=6.14 $Y2=2.38
r153 58 82 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.055 $Y=2.295
+ $X2=6.055 $Y2=2.38
r154 58 60 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.055 $Y=2.295
+ $X2=6.055 $Y2=1.96
r155 56 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.97 $Y=2.38
+ $X2=6.055 $Y2=2.38
r156 56 57 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.97 $Y=2.38
+ $X2=5.2 $Y2=2.38
r157 53 57 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=5.087 $Y=2.295
+ $X2=5.2 $Y2=2.38
r158 53 55 17.1586 $w=2.23e-07 $l=3.35e-07 $layer=LI1_cond $X=5.087 $Y=2.295
+ $X2=5.087 $Y2=1.96
r159 52 55 12.0366 $w=2.23e-07 $l=2.35e-07 $layer=LI1_cond $X=5.087 $Y=1.725
+ $X2=5.087 $Y2=1.96
r160 51 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.205 $Y=1.64
+ $X2=4.12 $Y2=1.64
r161 50 52 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=4.975 $Y=1.64
+ $X2=5.087 $Y2=1.725
r162 50 51 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.975 $Y=1.64
+ $X2=4.205 $Y2=1.64
r163 46 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.12 $Y=1.725
+ $X2=4.12 $Y2=1.64
r164 46 48 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.12 $Y=1.725
+ $X2=4.12 $Y2=1.96
r165 45 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.265 $Y=1.64
+ $X2=3.18 $Y2=1.64
r166 44 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.035 $Y=1.64
+ $X2=4.12 $Y2=1.64
r167 44 45 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.035 $Y=1.64
+ $X2=3.265 $Y2=1.64
r168 40 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.18 $Y=1.725
+ $X2=3.18 $Y2=1.64
r169 40 42 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.18 $Y=1.725
+ $X2=3.18 $Y2=1.96
r170 39 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.325 $Y=1.64
+ $X2=2.24 $Y2=1.64
r171 38 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=1.64
+ $X2=3.18 $Y2=1.64
r172 38 39 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.095 $Y=1.64
+ $X2=2.325 $Y2=1.64
r173 34 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=1.725
+ $X2=2.24 $Y2=1.64
r174 34 36 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.24 $Y=1.725
+ $X2=2.24 $Y2=1.96
r175 32 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=1.64
+ $X2=2.24 $Y2=1.64
r176 32 33 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.155 $Y=1.64
+ $X2=1.385 $Y2=1.64
r177 28 33 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.28 $Y=1.725
+ $X2=1.385 $Y2=1.64
r178 28 30 27.1991 $w=2.08e-07 $l=5.15e-07 $layer=LI1_cond $X=1.28 $Y=1.725
+ $X2=1.28 $Y2=2.24
r179 9 78 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=8.73
+ $Y=1.485 $X2=8.875 $Y2=1.96
r180 8 72 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=7.79
+ $Y=1.485 $X2=7.935 $Y2=1.96
r181 7 66 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.85
+ $Y=1.485 $X2=6.995 $Y2=1.96
r182 6 60 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.91
+ $Y=1.485 $X2=6.055 $Y2=1.96
r183 5 55 300 $w=1.7e-07 $l=4.94823e-07 $layer=licon1_PDIFF $count=2 $X=4.915
+ $Y=1.545 $X2=5.09 $Y2=1.96
r184 4 48 300 $w=1.7e-07 $l=4.82079e-07 $layer=licon1_PDIFF $count=2 $X=3.975
+ $Y=1.545 $X2=4.12 $Y2=1.96
r185 3 42 300 $w=1.7e-07 $l=4.82079e-07 $layer=licon1_PDIFF $count=2 $X=3.035
+ $Y=1.545 $X2=3.18 $Y2=1.96
r186 2 36 300 $w=1.7e-07 $l=4.82079e-07 $layer=licon1_PDIFF $count=2 $X=2.095
+ $Y=1.545 $X2=2.24 $Y2=1.96
r187 1 30 600 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_PDIFF $count=1 $X=1.175
+ $Y=1.545 $X2=1.3 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_8%Z 1 2 3 4 5 6 7 8 31 33 36 37 38 39 40 41
+ 42 43 44 61 66 67 70 74 80 94 99
c112 94 0 1.79447e-19 $X=5.707 $Y=1.87
c113 36 0 3.16397e-19 $X=5.775 $Y=1.53
r114 96 99 3.16609 $w=5.08e-07 $l=1.35e-07 $layer=LI1_cond $X=6.5 $Y=1.87
+ $X2=6.635 $Y2=1.87
r115 96 97 2.46227 $w=3.8e-07 $l=2.55e-07 $layer=LI1_cond $X=6.5 $Y=1.87 $X2=6.5
+ $Y2=1.615
r116 91 94 3.44752 $w=5.08e-07 $l=1.47e-07 $layer=LI1_cond $X=5.56 $Y=1.87
+ $X2=5.707 $Y2=1.87
r117 91 92 2.46227 $w=3.8e-07 $l=2.55e-07 $layer=LI1_cond $X=5.56 $Y=1.87
+ $X2=5.56 $Y2=1.615
r118 68 70 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.69 $Y=1.53
+ $X2=6.695 $Y2=1.53
r119 67 74 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.25 $Y=1.53
+ $X2=7.155 $Y2=1.53
r120 61 66 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.31 $Y=1.53
+ $X2=6.235 $Y2=1.53
r121 43 80 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.38 $Y=1.53
+ $X2=8.19 $Y2=1.53
r122 43 44 6.69888 $w=5.48e-07 $l=2.55e-07 $layer=LI1_cond $X=8.38 $Y=1.615
+ $X2=8.38 $Y2=1.87
r123 42 80 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.985 $Y=1.53
+ $X2=8.19 $Y2=1.53
r124 42 81 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.985 $Y=1.53
+ $X2=7.63 $Y2=1.53
r125 40 67 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.44 $Y=1.53
+ $X2=7.25 $Y2=1.53
r126 40 81 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.44 $Y=1.53
+ $X2=7.63 $Y2=1.53
r127 40 41 6.69888 $w=5.48e-07 $l=2.55e-07 $layer=LI1_cond $X=7.44 $Y=1.615
+ $X2=7.44 $Y2=1.87
r128 39 74 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=7.135 $Y=1.53
+ $X2=7.155 $Y2=1.53
r129 38 97 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.5 $Y=1.53 $X2=6.5
+ $Y2=1.615
r130 38 61 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.5 $Y=1.53 $X2=6.31
+ $Y2=1.53
r131 38 68 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.5 $Y=1.53 $X2=6.69
+ $Y2=1.53
r132 38 99 10.1092 $w=1.1e-07 $l=2.55e-07 $layer=LI1_cond $X=6.635 $Y=1.615
+ $X2=6.635 $Y2=1.87
r133 38 39 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.72 $Y=1.53
+ $X2=7.135 $Y2=1.53
r134 38 70 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=6.72 $Y=1.53
+ $X2=6.695 $Y2=1.53
r135 37 66 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=6.215 $Y=1.53
+ $X2=6.235 $Y2=1.53
r136 36 62 4.59089 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=5.585 $Y=1.53
+ $X2=5.8 $Y2=1.53
r137 36 92 2.39067 $w=4.05e-07 $l=9.66954e-08 $layer=LI1_cond $X=5.585 $Y=1.53
+ $X2=5.56 $Y2=1.615
r138 36 94 11.8728 $w=8.5e-08 $l=2.55e-07 $layer=LI1_cond $X=5.707 $Y=1.615
+ $X2=5.707 $Y2=1.87
r139 36 37 25.9658 $w=1.68e-07 $l=3.98e-07 $layer=LI1_cond $X=5.817 $Y=1.53
+ $X2=6.215 $Y2=1.53
r140 36 62 1.10909 $w=1.68e-07 $l=1.7e-08 $layer=LI1_cond $X=5.817 $Y=1.53
+ $X2=5.8 $Y2=1.53
r141 33 36 13.3078 $w=5.63e-07 $l=5.95e-07 $layer=LI1_cond $X=5.585 $Y=0.85
+ $X2=5.585 $Y2=1.445
r142 33 35 2.62515 $w=4.3e-07 $l=1.08e-07 $layer=LI1_cond $X=5.585 $Y=0.85
+ $X2=5.585 $Y2=0.742
r143 29 31 50.3859 $w=2.13e-07 $l=9.4e-07 $layer=LI1_cond $X=7.465 $Y=0.742
+ $X2=8.405 $Y2=0.742
r144 27 29 50.3859 $w=2.13e-07 $l=9.4e-07 $layer=LI1_cond $X=6.525 $Y=0.742
+ $X2=7.465 $Y2=0.742
r145 25 35 5.226 $w=2.15e-07 $l=2.15e-07 $layer=LI1_cond $X=5.8 $Y=0.742
+ $X2=5.585 $Y2=0.742
r146 25 27 38.8615 $w=2.13e-07 $l=7.25e-07 $layer=LI1_cond $X=5.8 $Y=0.742
+ $X2=6.525 $Y2=0.742
r147 8 43 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=8.26
+ $Y=1.485 $X2=8.405 $Y2=1.61
r148 7 40 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=7.32
+ $Y=1.485 $X2=7.465 $Y2=1.61
r149 6 38 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=6.38
+ $Y=1.485 $X2=6.525 $Y2=1.61
r150 5 36 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=5.44
+ $Y=1.485 $X2=5.585 $Y2=1.61
r151 4 31 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=8.22
+ $Y=0.235 $X2=8.405 $Y2=0.76
r152 3 29 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=7.28
+ $Y=0.235 $X2=7.465 $Y2=0.76
r153 2 27 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=6.34
+ $Y=0.235 $X2=6.525 $Y2=0.76
r154 1 35 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=5.4
+ $Y=0.235 $X2=5.585 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_8%VGND 1 2 3 4 5 18 22 26 30 32 36 38 40 45
+ 50 55 65 66 69 72 75 78 81
r130 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r131 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r132 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r133 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r134 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r135 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r136 65 66 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r137 63 66 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=4.83 $Y=0 $X2=8.97
+ $Y2=0
r138 63 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=4.37
+ $Y2=0
r139 62 65 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=4.83 $Y=0 $X2=8.97
+ $Y2=0
r140 62 63 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r141 60 81 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.685 $Y=0 $X2=4.49
+ $Y2=0
r142 60 62 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.685 $Y=0
+ $X2=4.83 $Y2=0
r143 59 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r144 59 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r145 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r146 56 75 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.605
+ $Y2=0
r147 56 58 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.795 $Y=0
+ $X2=2.99 $Y2=0
r148 55 78 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.355 $Y=0 $X2=3.545
+ $Y2=0
r149 55 58 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.355 $Y=0
+ $X2=2.99 $Y2=0
r150 54 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r151 54 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r152 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r153 51 72 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.665
+ $Y2=0
r154 51 53 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.855 $Y=0
+ $X2=2.07 $Y2=0
r155 50 75 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=2.605
+ $Y2=0
r156 50 53 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=2.07
+ $Y2=0
r157 49 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r158 49 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r159 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r160 46 69 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r161 46 48 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r162 45 72 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.665
+ $Y2=0
r163 45 48 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.475 $Y=0
+ $X2=1.15 $Y2=0
r164 40 69 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r165 40 42 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r166 38 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r167 38 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r168 34 81 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=0.085
+ $X2=4.49 $Y2=0
r169 34 36 8.1262 $w=3.88e-07 $l=2.75e-07 $layer=LI1_cond $X=4.49 $Y=0.085
+ $X2=4.49 $Y2=0.36
r170 33 78 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.735 $Y=0 $X2=3.545
+ $Y2=0
r171 32 81 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.295 $Y=0 $X2=4.49
+ $Y2=0
r172 32 33 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.295 $Y=0
+ $X2=3.735 $Y2=0
r173 28 78 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.545 $Y=0.085
+ $X2=3.545 $Y2=0
r174 28 30 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=3.545 $Y=0.085
+ $X2=3.545 $Y2=0.36
r175 24 75 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=0.085
+ $X2=2.605 $Y2=0
r176 24 26 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=2.605 $Y=0.085
+ $X2=2.605 $Y2=0.36
r177 20 72 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=0.085
+ $X2=1.665 $Y2=0
r178 20 22 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=1.665 $Y=0.085
+ $X2=1.665 $Y2=0.36
r179 16 69 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r180 16 18 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.36
r181 5 36 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.375
+ $Y=0.235 $X2=4.51 $Y2=0.36
r182 4 30 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=3.385
+ $Y=0.235 $X2=3.57 $Y2=0.36
r183 3 26 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=2.445
+ $Y=0.235 $X2=2.63 $Y2=0.36
r184 2 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.235 $X2=1.69 $Y2=0.36
r185 1 18 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_8%A_213_47# 1 2 3 4 5 6 7 8 9 30 32 33 36 38
+ 42 44 48 50 55 56 64 66 67 68
c105 67 0 9.78995e-20 $X=3.1 $Y=0.74
c106 66 0 9.78995e-20 $X=2.16 $Y=0.74
c107 50 0 3.37278e-19 $X=4.855 $Y=0.74
c108 44 0 5.75845e-19 $X=3.955 $Y=0.74
c109 38 0 5.75845e-19 $X=3.015 $Y=0.74
c110 32 0 5.33433e-19 $X=2.075 $Y=0.74
r111 62 64 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=7.935 $Y=0.36
+ $X2=8.875 $Y2=0.36
r112 60 62 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=6.995 $Y=0.36
+ $X2=7.935 $Y2=0.36
r113 58 60 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=6.055 $Y=0.36
+ $X2=6.995 $Y2=0.36
r114 56 58 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=5.2 $Y=0.36
+ $X2=6.055 $Y2=0.36
r115 53 55 4.0085 $w=3.43e-07 $l=1.2e-07 $layer=LI1_cond $X=5.027 $Y=0.655
+ $X2=5.027 $Y2=0.535
r116 52 56 7.35458 $w=2.1e-07 $l=2.19303e-07 $layer=LI1_cond $X=5.027 $Y=0.465
+ $X2=5.2 $Y2=0.36
r117 52 55 2.33829 $w=3.43e-07 $l=7e-08 $layer=LI1_cond $X=5.027 $Y=0.465
+ $X2=5.027 $Y2=0.535
r118 51 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.125 $Y=0.74
+ $X2=4.04 $Y2=0.74
r119 50 53 7.89393 $w=1.7e-07 $l=2.10247e-07 $layer=LI1_cond $X=4.855 $Y=0.74
+ $X2=5.027 $Y2=0.655
r120 50 51 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.855 $Y=0.74
+ $X2=4.125 $Y2=0.74
r121 46 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=0.655
+ $X2=4.04 $Y2=0.74
r122 46 48 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.04 $Y=0.655
+ $X2=4.04 $Y2=0.535
r123 45 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=0.74
+ $X2=3.1 $Y2=0.74
r124 44 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.955 $Y=0.74
+ $X2=4.04 $Y2=0.74
r125 44 45 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.955 $Y=0.74
+ $X2=3.185 $Y2=0.74
r126 40 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=0.655 $X2=3.1
+ $Y2=0.74
r127 40 42 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.1 $Y=0.655
+ $X2=3.1 $Y2=0.535
r128 39 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0.74
+ $X2=2.16 $Y2=0.74
r129 38 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0.74
+ $X2=3.1 $Y2=0.74
r130 38 39 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.015 $Y=0.74
+ $X2=2.245 $Y2=0.74
r131 34 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.655
+ $X2=2.16 $Y2=0.74
r132 34 36 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.16 $Y=0.655
+ $X2=2.16 $Y2=0.535
r133 32 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0.74
+ $X2=2.16 $Y2=0.74
r134 32 33 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.075 $Y=0.74
+ $X2=1.305 $Y2=0.74
r135 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.22 $Y=0.655
+ $X2=1.305 $Y2=0.74
r136 28 30 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.22 $Y=0.655
+ $X2=1.22 $Y2=0.535
r137 9 64 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=8.69
+ $Y=0.235 $X2=8.875 $Y2=0.36
r138 8 62 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=7.75
+ $Y=0.235 $X2=7.935 $Y2=0.36
r139 7 60 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=6.81
+ $Y=0.235 $X2=6.995 $Y2=0.36
r140 6 58 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=5.87
+ $Y=0.235 $X2=6.055 $Y2=0.36
r141 5 55 182 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_NDIFF $count=1 $X=4.99
+ $Y=0.235 $X2=5.115 $Y2=0.535
r142 4 48 182 $w=1.7e-07 $l=3.81445e-07 $layer=licon1_NDIFF $count=1 $X=3.855
+ $Y=0.235 $X2=4.04 $Y2=0.535
r143 3 42 182 $w=1.7e-07 $l=3.81445e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.235 $X2=3.1 $Y2=0.535
r144 2 36 182 $w=1.7e-07 $l=3.81445e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.16 $Y2=0.535
r145 1 30 182 $w=1.7e-07 $l=3.69459e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.22 $Y2=0.535
.ends

