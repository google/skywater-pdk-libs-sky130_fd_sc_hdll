# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__clkinv_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkinv_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.332000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.065000 2.910000 1.290000 ;
    END
  END A
  PIN VGND
    ANTENNADIFFAREA  0.485100 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.270000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  1.177200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.725000 3.570000 0.895000 ;
        RECT 0.105000 0.895000 0.275000 1.460000 ;
        RECT 0.105000 1.460000 3.570000 1.630000 ;
        RECT 0.655000 1.630000 0.910000 2.435000 ;
        RECT 1.130000 0.280000 1.390000 0.725000 ;
        RECT 1.615000 1.630000 1.870000 2.435000 ;
        RECT 2.090000 0.280000 2.345000 0.725000 ;
        RECT 2.570000 1.630000 2.830000 2.435000 ;
        RECT 3.270000 0.895000 3.570000 1.460000 ;
    END
  END Y
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  1.800000 0.430000 2.635000 ;
      RECT 0.565000  0.085000 0.910000 0.555000 ;
      RECT 1.130000  1.800000 1.390000 2.635000 ;
      RECT 1.610000  0.085000 1.870000 0.555000 ;
      RECT 2.090000  1.800000 2.350000 2.635000 ;
      RECT 2.565000  0.085000 2.865000 0.555000 ;
      RECT 3.050000  1.800000 3.435000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinv_4
END LIBRARY
