* File: sky130_fd_sc_hdll__xnor2_4.pxi.spice
* Created: Thu Aug 27 19:29:15 2020
* 
x_PM_SKY130_FD_SC_HDLL__XNOR2_4%B N_B_c_153_n N_B_M1007_g N_B_c_164_n
+ N_B_M1005_g N_B_c_154_n N_B_M1021_g N_B_c_165_n N_B_M1012_g N_B_c_155_n
+ N_B_M1037_g N_B_c_166_n N_B_M1016_g N_B_c_167_n N_B_M1034_g N_B_c_156_n
+ N_B_M1038_g N_B_c_157_n N_B_M1002_g N_B_c_168_n N_B_M1006_g N_B_c_158_n
+ N_B_M1011_g N_B_c_169_n N_B_M1020_g N_B_c_159_n N_B_M1023_g N_B_c_170_n
+ N_B_M1028_g N_B_c_171_n N_B_M1036_g N_B_c_160_n N_B_M1039_g N_B_c_172_n
+ N_B_c_173_n N_B_c_174_n N_B_c_175_n N_B_c_197_p N_B_c_161_n N_B_c_194_p B
+ N_B_c_162_n N_B_c_163_n B PM_SKY130_FD_SC_HDLL__XNOR2_4%B
x_PM_SKY130_FD_SC_HDLL__XNOR2_4%A N_A_c_356_n N_A_M1009_g N_A_c_367_n
+ N_A_M1015_g N_A_c_357_n N_A_M1030_g N_A_c_368_n N_A_M1019_g N_A_c_358_n
+ N_A_M1031_g N_A_c_369_n N_A_M1027_g N_A_c_370_n N_A_M1035_g N_A_c_359_n
+ N_A_M1032_g N_A_c_360_n N_A_M1004_g N_A_c_371_n N_A_M1000_g N_A_c_361_n
+ N_A_M1022_g N_A_c_372_n N_A_M1013_g N_A_c_362_n N_A_M1025_g N_A_c_373_n
+ N_A_M1018_g N_A_c_374_n N_A_M1026_g N_A_c_363_n N_A_M1033_g A N_A_c_364_n
+ N_A_c_365_n N_A_c_366_n A PM_SKY130_FD_SC_HDLL__XNOR2_4%A
x_PM_SKY130_FD_SC_HDLL__XNOR2_4%A_38_297# N_A_38_297#_M1007_d
+ N_A_38_297#_M1037_d N_A_38_297#_M1005_d N_A_38_297#_M1012_d
+ N_A_38_297#_M1034_d N_A_38_297#_M1019_d N_A_38_297#_M1035_d
+ N_A_38_297#_c_508_n N_A_38_297#_M1003_g N_A_38_297#_c_519_n
+ N_A_38_297#_M1001_g N_A_38_297#_c_509_n N_A_38_297#_M1010_g
+ N_A_38_297#_c_520_n N_A_38_297#_M1008_g N_A_38_297#_c_510_n
+ N_A_38_297#_M1014_g N_A_38_297#_c_521_n N_A_38_297#_M1017_g
+ N_A_38_297#_c_522_n N_A_38_297#_M1029_g N_A_38_297#_c_511_n
+ N_A_38_297#_M1024_g N_A_38_297#_c_512_n N_A_38_297#_c_524_n
+ N_A_38_297#_c_513_n N_A_38_297#_c_514_n N_A_38_297#_c_525_n
+ N_A_38_297#_c_526_n N_A_38_297#_c_555_n N_A_38_297#_c_561_n
+ N_A_38_297#_c_562_n N_A_38_297#_c_515_n N_A_38_297#_c_516_n
+ N_A_38_297#_c_517_n N_A_38_297#_c_528_n N_A_38_297#_c_618_p
+ N_A_38_297#_c_567_n N_A_38_297#_c_568_n N_A_38_297#_c_529_n
+ N_A_38_297#_c_530_n N_A_38_297#_c_531_n N_A_38_297#_c_532_n
+ N_A_38_297#_c_533_n N_A_38_297#_c_518_n
+ PM_SKY130_FD_SC_HDLL__XNOR2_4%A_38_297#
x_PM_SKY130_FD_SC_HDLL__XNOR2_4%VPWR N_VPWR_M1005_s N_VPWR_M1016_s
+ N_VPWR_M1015_s N_VPWR_M1027_s N_VPWR_M1000_d N_VPWR_M1018_d N_VPWR_M1001_s
+ N_VPWR_M1017_s N_VPWR_c_732_n N_VPWR_c_733_n N_VPWR_c_734_n N_VPWR_c_735_n
+ N_VPWR_c_736_n N_VPWR_c_737_n N_VPWR_c_738_n N_VPWR_c_739_n N_VPWR_c_740_n
+ N_VPWR_c_741_n N_VPWR_c_742_n N_VPWR_c_743_n N_VPWR_c_744_n N_VPWR_c_745_n
+ N_VPWR_c_746_n N_VPWR_c_747_n N_VPWR_c_748_n N_VPWR_c_749_n N_VPWR_c_750_n
+ N_VPWR_c_751_n N_VPWR_c_752_n N_VPWR_c_753_n VPWR N_VPWR_c_754_n
+ N_VPWR_c_731_n N_VPWR_c_756_n PM_SKY130_FD_SC_HDLL__XNOR2_4%VPWR
x_PM_SKY130_FD_SC_HDLL__XNOR2_4%A_898_297# N_A_898_297#_M1000_s
+ N_A_898_297#_M1013_s N_A_898_297#_M1026_s N_A_898_297#_M1020_s
+ N_A_898_297#_M1036_s N_A_898_297#_c_894_n N_A_898_297#_c_895_n
+ N_A_898_297#_c_897_n N_A_898_297#_c_938_n N_A_898_297#_c_890_n
+ N_A_898_297#_c_891_n N_A_898_297#_c_903_n
+ PM_SKY130_FD_SC_HDLL__XNOR2_4%A_898_297#
x_PM_SKY130_FD_SC_HDLL__XNOR2_4%Y N_Y_M1003_s N_Y_M1014_s N_Y_M1006_d
+ N_Y_M1028_d N_Y_M1001_d N_Y_M1008_d N_Y_M1029_d N_Y_c_956_n N_Y_c_957_n
+ N_Y_c_958_n N_Y_c_954_n N_Y_c_1016_n N_Y_c_959_n N_Y_c_960_n N_Y_c_961_n
+ N_Y_c_962_n N_Y_c_963_n Y Y PM_SKY130_FD_SC_HDLL__XNOR2_4%Y
x_PM_SKY130_FD_SC_HDLL__XNOR2_4%A_38_47# N_A_38_47#_M1007_s N_A_38_47#_M1021_s
+ N_A_38_47#_M1038_s N_A_38_47#_M1030_d N_A_38_47#_M1032_d N_A_38_47#_c_1038_n
+ N_A_38_47#_c_1050_n N_A_38_47#_c_1039_n N_A_38_47#_c_1040_n
+ N_A_38_47#_c_1058_n N_A_38_47#_c_1041_n N_A_38_47#_c_1042_n
+ N_A_38_47#_c_1043_n PM_SKY130_FD_SC_HDLL__XNOR2_4%A_38_47#
x_PM_SKY130_FD_SC_HDLL__XNOR2_4%VGND N_VGND_M1009_s N_VGND_M1031_s
+ N_VGND_M1004_d N_VGND_M1022_d N_VGND_M1033_d N_VGND_M1011_d N_VGND_M1039_d
+ N_VGND_c_1110_n N_VGND_c_1111_n N_VGND_c_1112_n N_VGND_c_1113_n
+ N_VGND_c_1114_n N_VGND_c_1115_n N_VGND_c_1116_n N_VGND_c_1117_n
+ N_VGND_c_1118_n N_VGND_c_1119_n N_VGND_c_1120_n N_VGND_c_1121_n
+ N_VGND_c_1122_n N_VGND_c_1123_n N_VGND_c_1124_n N_VGND_c_1125_n
+ N_VGND_c_1126_n N_VGND_c_1127_n N_VGND_c_1128_n N_VGND_c_1129_n
+ N_VGND_c_1130_n VGND N_VGND_c_1131_n N_VGND_c_1132_n
+ PM_SKY130_FD_SC_HDLL__XNOR2_4%VGND
x_PM_SKY130_FD_SC_HDLL__XNOR2_4%A_980_47# N_A_980_47#_M1004_s
+ N_A_980_47#_M1025_s N_A_980_47#_M1002_s N_A_980_47#_M1023_s
+ N_A_980_47#_M1003_d N_A_980_47#_M1010_d N_A_980_47#_M1024_d
+ N_A_980_47#_c_1304_n N_A_980_47#_c_1269_n N_A_980_47#_c_1270_n
+ N_A_980_47#_c_1315_n N_A_980_47#_c_1271_n N_A_980_47#_c_1283_n
+ N_A_980_47#_c_1272_n N_A_980_47#_c_1290_n N_A_980_47#_c_1273_n
+ N_A_980_47#_c_1274_n N_A_980_47#_c_1275_n N_A_980_47#_c_1276_n
+ N_A_980_47#_c_1277_n N_A_980_47#_c_1278_n N_A_980_47#_c_1279_n
+ PM_SKY130_FD_SC_HDLL__XNOR2_4%A_980_47#
cc_1 VNB N_B_c_153_n 0.0197003f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_2 VNB N_B_c_154_n 0.016746f $X=-0.19 $Y=-0.24 $X2=1.015 $Y2=0.995
cc_3 VNB N_B_c_155_n 0.017207f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=0.995
cc_4 VNB N_B_c_156_n 0.0171597f $X=-0.19 $Y=-0.24 $X2=2.005 $Y2=0.995
cc_5 VNB N_B_c_157_n 0.0164943f $X=-0.19 $Y=-0.24 $X2=6.705 $Y2=0.995
cc_6 VNB N_B_c_158_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=7.175 $Y2=0.995
cc_7 VNB N_B_c_159_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=7.645 $Y2=0.995
cc_8 VNB N_B_c_160_n 0.0224106f $X=-0.19 $Y=-0.24 $X2=8.165 $Y2=0.995
cc_9 VNB N_B_c_161_n 0.00499013f $X=-0.19 $Y=-0.24 $X2=8 $Y2=1.16
cc_10 VNB N_B_c_162_n 0.0780001f $X=-0.19 $Y=-0.24 $X2=1.98 $Y2=1.202
cc_11 VNB N_B_c_163_n 0.0790137f $X=-0.19 $Y=-0.24 $X2=8.14 $Y2=1.202
cc_12 VNB N_A_c_356_n 0.0164797f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_13 VNB N_A_c_357_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=1.015 $Y2=0.995
cc_14 VNB N_A_c_358_n 0.0172028f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=0.995
cc_15 VNB N_A_c_359_n 0.0223965f $X=-0.19 $Y=-0.24 $X2=2.005 $Y2=0.995
cc_16 VNB N_A_c_360_n 0.0218461f $X=-0.19 $Y=-0.24 $X2=6.705 $Y2=0.995
cc_17 VNB N_A_c_361_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=7.175 $Y2=0.995
cc_18 VNB N_A_c_362_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=7.645 $Y2=0.995
cc_19 VNB N_A_c_363_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=8.165 $Y2=0.995
cc_20 VNB N_A_c_364_n 0.0818185f $X=-0.19 $Y=-0.24 $X2=1.835 $Y2=1.175
cc_21 VNB N_A_c_365_n 0.0220999f $X=-0.19 $Y=-0.24 $X2=1.51 $Y2=1.202
cc_22 VNB N_A_c_366_n 0.0805043f $X=-0.19 $Y=-0.24 $X2=1.825 $Y2=1.16
cc_23 VNB N_A_38_297#_c_508_n 0.0218502f $X=-0.19 $Y=-0.24 $X2=2.005 $Y2=0.995
cc_24 VNB N_A_38_297#_c_509_n 0.0167673f $X=-0.19 $Y=-0.24 $X2=6.73 $Y2=1.41
cc_25 VNB N_A_38_297#_c_510_n 0.0171817f $X=-0.19 $Y=-0.24 $X2=7.2 $Y2=1.41
cc_26 VNB N_A_38_297#_c_511_n 0.020075f $X=-0.19 $Y=-0.24 $X2=8.14 $Y2=1.41
cc_27 VNB N_A_38_297#_c_512_n 0.0205891f $X=-0.19 $Y=-0.24 $X2=8.165 $Y2=0.56
cc_28 VNB N_A_38_297#_c_513_n 0.0129845f $X=-0.19 $Y=-0.24 $X2=6.185 $Y2=1.445
cc_29 VNB N_A_38_297#_c_514_n 0.00940401f $X=-0.19 $Y=-0.24 $X2=6.83 $Y2=1.16
cc_30 VNB N_A_38_297#_c_515_n 7.96611e-19 $X=-0.19 $Y=-0.24 $X2=6.73 $Y2=1.202
cc_31 VNB N_A_38_297#_c_516_n 0.0041373f $X=-0.19 $Y=-0.24 $X2=6.83 $Y2=1.202
cc_32 VNB N_A_38_297#_c_517_n 0.0120004f $X=-0.19 $Y=-0.24 $X2=8 $Y2=1.202
cc_33 VNB N_A_38_297#_c_518_n 0.0827747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_731_n 0.459507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_Y_c_954_n 0.0195576f $X=-0.19 $Y=-0.24 $X2=7.2 $Y2=1.41
cc_36 VNB Y 0.0197952f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_37 VNB N_A_38_47#_c_1038_n 0.00936711f $X=-0.19 $Y=-0.24 $X2=1.51 $Y2=1.41
cc_38 VNB N_A_38_47#_c_1039_n 0.00321738f $X=-0.19 $Y=-0.24 $X2=2.005 $Y2=0.56
cc_39 VNB N_A_38_47#_c_1040_n 0.0023309f $X=-0.19 $Y=-0.24 $X2=2.005 $Y2=0.56
cc_40 VNB N_A_38_47#_c_1041_n 0.00688745f $X=-0.19 $Y=-0.24 $X2=6.73 $Y2=1.985
cc_41 VNB N_A_38_47#_c_1042_n 0.00435124f $X=-0.19 $Y=-0.24 $X2=7.2 $Y2=1.41
cc_42 VNB N_A_38_47#_c_1043_n 0.0023781f $X=-0.19 $Y=-0.24 $X2=7.67 $Y2=1.41
cc_43 VNB N_VGND_c_1110_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=2.005 $Y2=0.56
cc_44 VNB N_VGND_c_1111_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=6.73 $Y2=1.41
cc_45 VNB N_VGND_c_1112_n 0.0141878f $X=-0.19 $Y=-0.24 $X2=7.175 $Y2=0.56
cc_46 VNB N_VGND_c_1113_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=7.2 $Y2=1.985
cc_47 VNB N_VGND_c_1114_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=7.67 $Y2=1.41
cc_48 VNB N_VGND_c_1115_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=8.14 $Y2=1.985
cc_49 VNB N_VGND_c_1116_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=8.165 $Y2=0.56
cc_50 VNB N_VGND_c_1117_n 0.0622586f $X=-0.19 $Y=-0.24 $X2=6.1 $Y2=1.53
cc_51 VNB N_VGND_c_1118_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=2.005 $Y2=1.53
cc_52 VNB N_VGND_c_1119_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=6.185 $Y2=1.445
cc_53 VNB N_VGND_c_1120_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=6.27 $Y2=1.175
cc_54 VNB N_VGND_c_1121_n 0.0185093f $X=-0.19 $Y=-0.24 $X2=6.83 $Y2=1.16
cc_55 VNB N_VGND_c_1122_n 0.00519006f $X=-0.19 $Y=-0.24 $X2=6.83 $Y2=1.16
cc_56 VNB N_VGND_c_1123_n 0.0198149f $X=-0.19 $Y=-0.24 $X2=8 $Y2=1.16
cc_57 VNB N_VGND_c_1124_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=8 $Y2=1.16
cc_58 VNB N_VGND_c_1125_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=1.835 $Y2=1.175
cc_59 VNB N_VGND_c_1126_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_60 VNB N_VGND_c_1127_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.202
cc_61 VNB N_VGND_c_1128_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0.57 $Y2=1.202
cc_62 VNB N_VGND_c_1129_n 0.0192991f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_63 VNB N_VGND_c_1130_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_64 VNB N_VGND_c_1131_n 0.0644428f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1132_n 0.516244f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_980_47#_c_1269_n 0.0023309f $X=-0.19 $Y=-0.24 $X2=6.705 $Y2=0.56
cc_67 VNB N_A_980_47#_c_1270_n 0.0023781f $X=-0.19 $Y=-0.24 $X2=6.705 $Y2=0.56
cc_68 VNB N_A_980_47#_c_1271_n 0.00250477f $X=-0.19 $Y=-0.24 $X2=7.175 $Y2=0.56
cc_69 VNB N_A_980_47#_c_1272_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=7.645 $Y2=0.56
cc_70 VNB N_A_980_47#_c_1273_n 0.0129582f $X=-0.19 $Y=-0.24 $X2=8.14 $Y2=1.985
cc_71 VNB N_A_980_47#_c_1274_n 0.0020206f $X=-0.19 $Y=-0.24 $X2=8.165 $Y2=0.995
cc_72 VNB N_A_980_47#_c_1275_n 0.00295808f $X=-0.19 $Y=-0.24 $X2=1.92 $Y2=1.275
cc_73 VNB N_A_980_47#_c_1276_n 0.00777546f $X=-0.19 $Y=-0.24 $X2=6.185 $Y2=1.445
cc_74 VNB N_A_980_47#_c_1277_n 0.00291575f $X=-0.19 $Y=-0.24 $X2=6.83 $Y2=1.175
cc_75 VNB N_A_980_47#_c_1278_n 0.00241121f $X=-0.19 $Y=-0.24 $X2=6.83 $Y2=1.16
cc_76 VNB N_A_980_47#_c_1279_n 0.00280763f $X=-0.19 $Y=-0.24 $X2=6.83 $Y2=1.16
cc_77 VPB N_B_c_164_n 0.0191265f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=1.41
cc_78 VPB N_B_c_165_n 0.0156758f $X=-0.19 $Y=1.305 $X2=1.04 $Y2=1.41
cc_79 VPB N_B_c_166_n 0.0159744f $X=-0.19 $Y=1.305 $X2=1.51 $Y2=1.41
cc_80 VPB N_B_c_167_n 0.015791f $X=-0.19 $Y=1.305 $X2=1.98 $Y2=1.41
cc_81 VPB N_B_c_168_n 0.0157854f $X=-0.19 $Y=1.305 $X2=6.73 $Y2=1.41
cc_82 VPB N_B_c_169_n 0.0158194f $X=-0.19 $Y=1.305 $X2=7.2 $Y2=1.41
cc_83 VPB N_B_c_170_n 0.0158011f $X=-0.19 $Y=1.305 $X2=7.67 $Y2=1.41
cc_84 VPB N_B_c_171_n 0.0191981f $X=-0.19 $Y=1.305 $X2=8.14 $Y2=1.41
cc_85 VPB N_B_c_172_n 0.00102646f $X=-0.19 $Y=1.305 $X2=1.92 $Y2=1.445
cc_86 VPB N_B_c_173_n 0.0324742f $X=-0.19 $Y=1.305 $X2=6.1 $Y2=1.53
cc_87 VPB N_B_c_174_n 2.91493e-19 $X=-0.19 $Y=1.305 $X2=2.005 $Y2=1.53
cc_88 VPB N_B_c_175_n 0.00117844f $X=-0.19 $Y=1.305 $X2=6.185 $Y2=1.445
cc_89 VPB N_B_c_162_n 0.0468004f $X=-0.19 $Y=1.305 $X2=1.98 $Y2=1.202
cc_90 VPB N_B_c_163_n 0.0455105f $X=-0.19 $Y=1.305 $X2=8.14 $Y2=1.202
cc_91 VPB N_A_c_367_n 0.015982f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=1.41
cc_92 VPB N_A_c_368_n 0.0158911f $X=-0.19 $Y=1.305 $X2=1.04 $Y2=1.41
cc_93 VPB N_A_c_369_n 0.0158911f $X=-0.19 $Y=1.305 $X2=1.51 $Y2=1.41
cc_94 VPB N_A_c_370_n 0.0201091f $X=-0.19 $Y=1.305 $X2=1.98 $Y2=1.41
cc_95 VPB N_A_c_371_n 0.0201091f $X=-0.19 $Y=1.305 $X2=6.73 $Y2=1.41
cc_96 VPB N_A_c_372_n 0.0158729f $X=-0.19 $Y=1.305 $X2=7.2 $Y2=1.41
cc_97 VPB N_A_c_373_n 0.0158659f $X=-0.19 $Y=1.305 $X2=7.67 $Y2=1.41
cc_98 VPB N_A_c_374_n 0.0158788f $X=-0.19 $Y=1.305 $X2=8.14 $Y2=1.41
cc_99 VPB N_A_c_364_n 0.0482897f $X=-0.19 $Y=1.305 $X2=1.835 $Y2=1.175
cc_100 VPB N_A_c_366_n 0.0482108f $X=-0.19 $Y=1.305 $X2=1.825 $Y2=1.16
cc_101 VPB N_A_38_297#_c_519_n 0.0194229f $X=-0.19 $Y=1.305 $X2=6.705 $Y2=0.995
cc_102 VPB N_A_38_297#_c_520_n 0.0158911f $X=-0.19 $Y=1.305 $X2=7.175 $Y2=0.995
cc_103 VPB N_A_38_297#_c_521_n 0.0158722f $X=-0.19 $Y=1.305 $X2=7.645 $Y2=0.995
cc_104 VPB N_A_38_297#_c_522_n 0.0191994f $X=-0.19 $Y=1.305 $X2=7.67 $Y2=1.41
cc_105 VPB N_A_38_297#_c_512_n 0.00744189f $X=-0.19 $Y=1.305 $X2=8.165 $Y2=0.56
cc_106 VPB N_A_38_297#_c_524_n 0.0361631f $X=-0.19 $Y=1.305 $X2=1.92 $Y2=1.445
cc_107 VPB N_A_38_297#_c_525_n 0.00196613f $X=-0.19 $Y=1.305 $X2=8 $Y2=1.16
cc_108 VPB N_A_38_297#_c_526_n 0.00126656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_38_297#_c_515_n 0.00382418f $X=-0.19 $Y=1.305 $X2=6.73 $Y2=1.202
cc_110 VPB N_A_38_297#_c_528_n 0.00959806f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.175
cc_111 VPB N_A_38_297#_c_529_n 0.00172606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_38_297#_c_530_n 0.0108211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_38_297#_c_531_n 0.00276658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_38_297#_c_532_n 0.00216367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_38_297#_c_533_n 0.00176105f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_38_297#_c_518_n 0.0465016f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_732_n 0.00516582f $X=-0.19 $Y=1.305 $X2=6.73 $Y2=1.985
cc_118 VPB N_VPWR_c_733_n 0.00516582f $X=-0.19 $Y=1.305 $X2=7.175 $Y2=0.56
cc_119 VPB N_VPWR_c_734_n 0.00516582f $X=-0.19 $Y=1.305 $X2=7.645 $Y2=0.995
cc_120 VPB N_VPWR_c_735_n 0.00516582f $X=-0.19 $Y=1.305 $X2=7.67 $Y2=1.985
cc_121 VPB N_VPWR_c_736_n 0.00516582f $X=-0.19 $Y=1.305 $X2=8.14 $Y2=1.985
cc_122 VPB N_VPWR_c_737_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.92 $Y2=1.275
cc_123 VPB N_VPWR_c_738_n 0.00516582f $X=-0.19 $Y=1.305 $X2=6.185 $Y2=1.275
cc_124 VPB N_VPWR_c_739_n 0.00516582f $X=-0.19 $Y=1.305 $X2=6.83 $Y2=1.16
cc_125 VPB N_VPWR_c_740_n 0.0187181f $X=-0.19 $Y=1.305 $X2=8 $Y2=1.16
cc_126 VPB N_VPWR_c_741_n 0.00478085f $X=-0.19 $Y=1.305 $X2=8 $Y2=1.16
cc_127 VPB N_VPWR_c_742_n 0.0178757f $X=-0.19 $Y=1.305 $X2=1.835 $Y2=1.175
cc_128 VPB N_VPWR_c_743_n 0.00478085f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_129 VPB N_VPWR_c_744_n 0.0178757f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.202
cc_130 VPB N_VPWR_c_745_n 0.00478085f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=1.202
cc_131 VPB N_VPWR_c_746_n 0.0314785f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_132 VPB N_VPWR_c_747_n 0.00478085f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_133 VPB N_VPWR_c_748_n 0.0178757f $X=-0.19 $Y=1.305 $X2=1.04 $Y2=1.202
cc_134 VPB N_VPWR_c_749_n 0.00478085f $X=-0.19 $Y=1.305 $X2=1.485 $Y2=1.202
cc_135 VPB N_VPWR_c_750_n 0.0724778f $X=-0.19 $Y=1.305 $X2=1.825 $Y2=1.202
cc_136 VPB N_VPWR_c_751_n 0.0047828f $X=-0.19 $Y=1.305 $X2=1.825 $Y2=1.16
cc_137 VPB N_VPWR_c_752_n 0.0195604f $X=-0.19 $Y=1.305 $X2=1.98 $Y2=1.202
cc_138 VPB N_VPWR_c_753_n 0.0047828f $X=-0.19 $Y=1.305 $X2=2.005 $Y2=1.202
cc_139 VPB N_VPWR_c_754_n 0.0183432f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_731_n 0.0582357f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_756_n 0.025056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_898_297#_c_890_n 0.00290477f $X=-0.19 $Y=1.305 $X2=6.73 $Y2=1.985
cc_143 VPB N_A_898_297#_c_891_n 0.00772957f $X=-0.19 $Y=1.305 $X2=7.175 $Y2=0.56
cc_144 VPB N_Y_c_956_n 0.0087186f $X=-0.19 $Y=1.305 $X2=2.005 $Y2=0.995
cc_145 VPB N_Y_c_957_n 0.00511278f $X=-0.19 $Y=1.305 $X2=6.73 $Y2=1.985
cc_146 VPB N_Y_c_958_n 0.00182418f $X=-0.19 $Y=1.305 $X2=7.175 $Y2=0.56
cc_147 VPB N_Y_c_959_n 0.00182418f $X=-0.19 $Y=1.305 $X2=8.14 $Y2=1.985
cc_148 VPB N_Y_c_960_n 0.0312141f $X=-0.19 $Y=1.305 $X2=8.165 $Y2=0.56
cc_149 VPB N_Y_c_961_n 0.00804849f $X=-0.19 $Y=1.305 $X2=1.92 $Y2=1.445
cc_150 VPB N_Y_c_962_n 0.00150464f $X=-0.19 $Y=1.305 $X2=6.83 $Y2=1.175
cc_151 VPB N_Y_c_963_n 0.0103549f $X=-0.19 $Y=1.305 $X2=8 $Y2=1.175
cc_152 VPB Y 0.00695062f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_153 N_B_c_156_n N_A_c_356_n 0.0175558f $X=2.005 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_154 N_B_c_167_n N_A_c_367_n 0.0227832f $X=1.98 $Y=1.41 $X2=0 $Y2=0
cc_155 N_B_c_173_n N_A_c_367_n 0.0120485f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_156 N_B_c_173_n N_A_c_368_n 0.01191f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_157 N_B_c_173_n N_A_c_369_n 0.01191f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_158 N_B_c_173_n N_A_c_370_n 0.0139099f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_159 N_B_c_173_n N_A_c_371_n 0.0139099f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_160 N_B_c_173_n N_A_c_372_n 0.01191f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_161 N_B_c_173_n N_A_c_373_n 0.01191f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_162 N_B_c_175_n N_A_c_373_n 6.69584e-19 $X=6.185 $Y=1.445 $X2=0 $Y2=0
cc_163 N_B_c_168_n N_A_c_374_n 0.0229184f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_164 N_B_c_173_n N_A_c_374_n 0.00588725f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_165 N_B_c_175_n N_A_c_374_n 6.69704e-19 $X=6.185 $Y=1.445 $X2=0 $Y2=0
cc_166 N_B_c_157_n N_A_c_363_n 0.024015f $X=6.705 $Y=0.995 $X2=0 $Y2=0
cc_167 N_B_c_172_n N_A_c_364_n 7.95752e-19 $X=1.92 $Y=1.445 $X2=0 $Y2=0
cc_168 N_B_c_173_n N_A_c_364_n 0.0231984f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_169 N_B_c_194_p N_A_c_364_n 8.04129e-19 $X=1.835 $Y=1.175 $X2=0 $Y2=0
cc_170 N_B_c_162_n N_A_c_364_n 0.0175558f $X=1.98 $Y=1.202 $X2=0 $Y2=0
cc_171 N_B_c_173_n N_A_c_365_n 0.232463f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_172 N_B_c_197_p N_A_c_365_n 0.0167609f $X=6.27 $Y=1.175 $X2=0 $Y2=0
cc_173 N_B_c_194_p N_A_c_365_n 0.00892702f $X=1.835 $Y=1.175 $X2=0 $Y2=0
cc_174 N_B_c_162_n N_A_c_365_n 8.75854e-19 $X=1.98 $Y=1.202 $X2=0 $Y2=0
cc_175 N_B_c_173_n N_A_c_366_n 0.0216414f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_176 N_B_c_175_n N_A_c_366_n 0.00915008f $X=6.185 $Y=1.445 $X2=0 $Y2=0
cc_177 N_B_c_197_p N_A_c_366_n 0.00835678f $X=6.27 $Y=1.175 $X2=0 $Y2=0
cc_178 N_B_c_161_n N_A_c_366_n 0.0071501f $X=8 $Y=1.16 $X2=0 $Y2=0
cc_179 N_B_c_163_n N_A_c_366_n 0.024015f $X=8.14 $Y=1.202 $X2=0 $Y2=0
cc_180 N_B_c_173_n N_A_38_297#_M1034_d 0.00187091f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_181 N_B_c_173_n N_A_38_297#_M1019_d 0.00187091f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_182 N_B_c_173_n N_A_38_297#_M1035_d 0.00290685f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_183 N_B_c_153_n N_A_38_297#_c_512_n 0.01758f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_184 N_B_c_164_n N_A_38_297#_c_512_n 0.00124753f $X=0.57 $Y=1.41 $X2=0 $Y2=0
cc_185 N_B_c_194_p N_A_38_297#_c_512_n 0.0162001f $X=1.835 $Y=1.175 $X2=0 $Y2=0
cc_186 N_B_c_153_n N_A_38_297#_c_514_n 0.0137135f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_187 N_B_c_154_n N_A_38_297#_c_514_n 0.0114466f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_188 N_B_c_155_n N_A_38_297#_c_514_n 0.0114367f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_189 N_B_c_156_n N_A_38_297#_c_514_n 2.03781e-19 $X=2.005 $Y=0.995 $X2=0 $Y2=0
cc_190 N_B_c_194_p N_A_38_297#_c_514_n 0.102985f $X=1.835 $Y=1.175 $X2=0 $Y2=0
cc_191 N_B_c_162_n N_A_38_297#_c_514_n 0.0117089f $X=1.98 $Y=1.202 $X2=0 $Y2=0
cc_192 N_B_c_164_n N_A_38_297#_c_525_n 0.0162122f $X=0.57 $Y=1.41 $X2=0 $Y2=0
cc_193 N_B_c_165_n N_A_38_297#_c_525_n 0.0137157f $X=1.04 $Y=1.41 $X2=0 $Y2=0
cc_194 N_B_c_194_p N_A_38_297#_c_525_n 0.0456097f $X=1.835 $Y=1.175 $X2=0 $Y2=0
cc_195 N_B_c_162_n N_A_38_297#_c_525_n 0.00851578f $X=1.98 $Y=1.202 $X2=0 $Y2=0
cc_196 N_B_c_166_n N_A_38_297#_c_526_n 8.97035e-19 $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_197 N_B_c_174_n N_A_38_297#_c_526_n 0.00288939f $X=2.005 $Y=1.53 $X2=0 $Y2=0
cc_198 N_B_c_194_p N_A_38_297#_c_526_n 0.0163163f $X=1.835 $Y=1.175 $X2=0 $Y2=0
cc_199 N_B_c_162_n N_A_38_297#_c_526_n 0.00639652f $X=1.98 $Y=1.202 $X2=0 $Y2=0
cc_200 N_B_c_166_n N_A_38_297#_c_555_n 0.014974f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_201 N_B_c_167_n N_A_38_297#_c_555_n 0.0132187f $X=1.98 $Y=1.41 $X2=0 $Y2=0
cc_202 N_B_c_173_n N_A_38_297#_c_555_n 0.00401135f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_203 N_B_c_174_n N_A_38_297#_c_555_n 0.00797024f $X=2.005 $Y=1.53 $X2=0 $Y2=0
cc_204 N_B_c_194_p N_A_38_297#_c_555_n 0.00506447f $X=1.835 $Y=1.175 $X2=0 $Y2=0
cc_205 N_B_c_162_n N_A_38_297#_c_555_n 0.00412753f $X=1.98 $Y=1.202 $X2=0 $Y2=0
cc_206 N_B_c_173_n N_A_38_297#_c_561_n 0.0343218f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_207 N_B_c_173_n N_A_38_297#_c_562_n 0.0343218f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_208 N_B_c_171_n N_A_38_297#_c_515_n 0.00120137f $X=8.14 $Y=1.41 $X2=0 $Y2=0
cc_209 N_B_c_163_n N_A_38_297#_c_515_n 0.00517635f $X=8.14 $Y=1.202 $X2=0 $Y2=0
cc_210 N_B_c_161_n N_A_38_297#_c_516_n 0.0145269f $X=8 $Y=1.16 $X2=0 $Y2=0
cc_211 N_B_c_163_n N_A_38_297#_c_516_n 0.00578652f $X=8.14 $Y=1.202 $X2=0 $Y2=0
cc_212 N_B_c_173_n N_A_38_297#_c_567_n 0.0128801f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_213 N_B_c_173_n N_A_38_297#_c_568_n 0.0128801f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_214 N_B_c_173_n N_A_38_297#_c_529_n 0.0155879f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_215 N_B_c_168_n N_A_38_297#_c_530_n 0.010423f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_216 N_B_c_169_n N_A_38_297#_c_530_n 0.011867f $X=7.2 $Y=1.41 $X2=0 $Y2=0
cc_217 N_B_c_170_n N_A_38_297#_c_530_n 0.01191f $X=7.67 $Y=1.41 $X2=0 $Y2=0
cc_218 N_B_c_171_n N_A_38_297#_c_530_n 0.0140267f $X=8.14 $Y=1.41 $X2=0 $Y2=0
cc_219 N_B_c_173_n N_A_38_297#_c_530_n 0.00921168f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_220 N_B_c_161_n N_A_38_297#_c_530_n 0.11541f $X=8 $Y=1.16 $X2=0 $Y2=0
cc_221 N_B_c_163_n N_A_38_297#_c_530_n 0.0231155f $X=8.14 $Y=1.202 $X2=0 $Y2=0
cc_222 N_B_c_166_n N_A_38_297#_c_531_n 0.00493162f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_223 N_B_c_173_n N_A_38_297#_c_531_n 0.17462f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_224 N_B_c_174_n N_A_38_297#_c_531_n 0.0133283f $X=2.005 $Y=1.53 $X2=0 $Y2=0
cc_225 N_B_c_161_n N_A_38_297#_c_531_n 0.00734938f $X=8 $Y=1.16 $X2=0 $Y2=0
cc_226 N_B_c_194_p N_A_38_297#_c_531_n 0.0117308f $X=1.835 $Y=1.175 $X2=0 $Y2=0
cc_227 N_B_c_162_n N_A_38_297#_c_531_n 0.00659266f $X=1.98 $Y=1.202 $X2=0 $Y2=0
cc_228 N_B_c_164_n N_A_38_297#_c_532_n 2.9548e-19 $X=0.57 $Y=1.41 $X2=0 $Y2=0
cc_229 N_B_c_165_n N_A_38_297#_c_532_n 0.00492291f $X=1.04 $Y=1.41 $X2=0 $Y2=0
cc_230 N_B_c_166_n N_A_38_297#_c_532_n 5.37077e-19 $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_231 N_B_c_172_n N_A_38_297#_c_532_n 0.00112885f $X=1.92 $Y=1.445 $X2=0 $Y2=0
cc_232 N_B_c_174_n N_A_38_297#_c_532_n 2.37459e-19 $X=2.005 $Y=1.53 $X2=0 $Y2=0
cc_233 N_B_c_194_p N_A_38_297#_c_532_n 0.00923763f $X=1.835 $Y=1.175 $X2=0 $Y2=0
cc_234 N_B_c_162_n N_A_38_297#_c_532_n 0.0076923f $X=1.98 $Y=1.202 $X2=0 $Y2=0
cc_235 N_B_c_168_n N_A_38_297#_c_533_n 0.00454953f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_236 N_B_c_169_n N_A_38_297#_c_533_n 0.00105392f $X=7.2 $Y=1.41 $X2=0 $Y2=0
cc_237 N_B_c_175_n N_A_38_297#_c_533_n 9.7358e-19 $X=6.185 $Y=1.445 $X2=0 $Y2=0
cc_238 N_B_c_161_n N_A_38_297#_c_533_n 0.00917598f $X=8 $Y=1.16 $X2=0 $Y2=0
cc_239 N_B_c_163_n N_A_38_297#_c_533_n 0.00522958f $X=8.14 $Y=1.202 $X2=0 $Y2=0
cc_240 N_B_c_173_n N_VPWR_M1015_s 0.00187547f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_241 N_B_c_173_n N_VPWR_M1027_s 0.00187547f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_242 N_B_c_173_n N_VPWR_M1000_d 0.00187547f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_243 N_B_c_173_n N_VPWR_M1018_d 0.00186949f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_244 N_B_c_164_n N_VPWR_c_732_n 0.00300743f $X=0.57 $Y=1.41 $X2=0 $Y2=0
cc_245 N_B_c_165_n N_VPWR_c_732_n 0.00300743f $X=1.04 $Y=1.41 $X2=0 $Y2=0
cc_246 N_B_c_166_n N_VPWR_c_733_n 0.00300743f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_247 N_B_c_167_n N_VPWR_c_733_n 0.00300743f $X=1.98 $Y=1.41 $X2=0 $Y2=0
cc_248 N_B_c_165_n N_VPWR_c_740_n 0.00702461f $X=1.04 $Y=1.41 $X2=0 $Y2=0
cc_249 N_B_c_166_n N_VPWR_c_740_n 0.00523784f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_250 N_B_c_167_n N_VPWR_c_742_n 0.00523784f $X=1.98 $Y=1.41 $X2=0 $Y2=0
cc_251 N_B_c_168_n N_VPWR_c_750_n 0.00429453f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_252 N_B_c_169_n N_VPWR_c_750_n 0.00429453f $X=7.2 $Y=1.41 $X2=0 $Y2=0
cc_253 N_B_c_170_n N_VPWR_c_750_n 0.00429453f $X=7.67 $Y=1.41 $X2=0 $Y2=0
cc_254 N_B_c_171_n N_VPWR_c_750_n 0.00429453f $X=8.14 $Y=1.41 $X2=0 $Y2=0
cc_255 N_B_c_164_n N_VPWR_c_731_n 0.0133833f $X=0.57 $Y=1.41 $X2=0 $Y2=0
cc_256 N_B_c_165_n N_VPWR_c_731_n 0.0124092f $X=1.04 $Y=1.41 $X2=0 $Y2=0
cc_257 N_B_c_166_n N_VPWR_c_731_n 0.00678659f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_258 N_B_c_167_n N_VPWR_c_731_n 0.0068118f $X=1.98 $Y=1.41 $X2=0 $Y2=0
cc_259 N_B_c_168_n N_VPWR_c_731_n 0.00609021f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_260 N_B_c_169_n N_VPWR_c_731_n 0.00606499f $X=7.2 $Y=1.41 $X2=0 $Y2=0
cc_261 N_B_c_170_n N_VPWR_c_731_n 0.00606499f $X=7.67 $Y=1.41 $X2=0 $Y2=0
cc_262 N_B_c_171_n N_VPWR_c_731_n 0.00734734f $X=8.14 $Y=1.41 $X2=0 $Y2=0
cc_263 N_B_c_164_n N_VPWR_c_756_n 0.00702461f $X=0.57 $Y=1.41 $X2=0 $Y2=0
cc_264 N_B_c_173_n N_A_898_297#_M1000_s 0.00290685f $X=6.1 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_265 N_B_c_173_n N_A_898_297#_M1013_s 0.00187091f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_266 N_B_c_173_n N_A_898_297#_c_894_n 0.0343218f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_267 N_B_c_173_n N_A_898_297#_c_895_n 0.0300521f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_268 N_B_c_161_n N_A_898_297#_c_895_n 0.00111905f $X=8 $Y=1.16 $X2=0 $Y2=0
cc_269 N_B_c_161_n N_A_898_297#_c_897_n 0.00165733f $X=8 $Y=1.16 $X2=0 $Y2=0
cc_270 N_B_c_168_n N_A_898_297#_c_890_n 0.0127106f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_271 N_B_c_169_n N_A_898_297#_c_890_n 0.0112654f $X=7.2 $Y=1.41 $X2=0 $Y2=0
cc_272 N_B_c_170_n N_A_898_297#_c_890_n 0.0112654f $X=7.67 $Y=1.41 $X2=0 $Y2=0
cc_273 N_B_c_171_n N_A_898_297#_c_890_n 0.0112654f $X=8.14 $Y=1.41 $X2=0 $Y2=0
cc_274 N_B_c_173_n N_A_898_297#_c_891_n 0.0205254f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_275 N_B_c_173_n N_A_898_297#_c_903_n 0.0128801f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_276 N_B_c_168_n N_Y_c_956_n 0.00547764f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_277 N_B_c_169_n N_Y_c_956_n 0.0124936f $X=7.2 $Y=1.41 $X2=0 $Y2=0
cc_278 N_B_c_170_n N_Y_c_956_n 0.0124936f $X=7.67 $Y=1.41 $X2=0 $Y2=0
cc_279 N_B_c_171_n N_Y_c_956_n 0.0151292f $X=8.14 $Y=1.41 $X2=0 $Y2=0
cc_280 N_B_c_171_n N_Y_c_961_n 0.00901245f $X=8.14 $Y=1.41 $X2=0 $Y2=0
cc_281 N_B_c_153_n N_A_38_47#_c_1038_n 0.00931157f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_282 N_B_c_154_n N_A_38_47#_c_1038_n 0.00931157f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_283 N_B_c_155_n N_A_38_47#_c_1038_n 0.00964761f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_284 N_B_c_156_n N_A_38_47#_c_1038_n 0.013027f $X=2.005 $Y=0.995 $X2=0 $Y2=0
cc_285 N_B_c_194_p N_A_38_47#_c_1038_n 0.00229057f $X=1.835 $Y=1.175 $X2=0 $Y2=0
cc_286 N_B_c_173_n N_A_38_47#_c_1039_n 0.00704591f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_287 N_B_c_157_n N_VGND_c_1114_n 0.00268723f $X=6.705 $Y=0.995 $X2=0 $Y2=0
cc_288 N_B_c_158_n N_VGND_c_1115_n 0.00379224f $X=7.175 $Y=0.995 $X2=0 $Y2=0
cc_289 N_B_c_159_n N_VGND_c_1115_n 0.00276126f $X=7.645 $Y=0.995 $X2=0 $Y2=0
cc_290 N_B_c_160_n N_VGND_c_1116_n 0.00438629f $X=8.165 $Y=0.995 $X2=0 $Y2=0
cc_291 N_B_c_153_n N_VGND_c_1117_n 0.00357877f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_292 N_B_c_154_n N_VGND_c_1117_n 0.00357877f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_293 N_B_c_155_n N_VGND_c_1117_n 0.00357877f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_294 N_B_c_156_n N_VGND_c_1117_n 0.00357877f $X=2.005 $Y=0.995 $X2=0 $Y2=0
cc_295 N_B_c_157_n N_VGND_c_1127_n 0.00423334f $X=6.705 $Y=0.995 $X2=0 $Y2=0
cc_296 N_B_c_158_n N_VGND_c_1127_n 0.00423334f $X=7.175 $Y=0.995 $X2=0 $Y2=0
cc_297 N_B_c_159_n N_VGND_c_1129_n 0.00423334f $X=7.645 $Y=0.995 $X2=0 $Y2=0
cc_298 N_B_c_160_n N_VGND_c_1129_n 0.00438411f $X=8.165 $Y=0.995 $X2=0 $Y2=0
cc_299 N_B_c_153_n N_VGND_c_1132_n 0.0063758f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_300 N_B_c_154_n N_VGND_c_1132_n 0.00548399f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_301 N_B_c_155_n N_VGND_c_1132_n 0.00560377f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_302 N_B_c_156_n N_VGND_c_1132_n 0.005504f $X=2.005 $Y=0.995 $X2=0 $Y2=0
cc_303 N_B_c_157_n N_VGND_c_1132_n 0.00587047f $X=6.705 $Y=0.995 $X2=0 $Y2=0
cc_304 N_B_c_158_n N_VGND_c_1132_n 0.006093f $X=7.175 $Y=0.995 $X2=0 $Y2=0
cc_305 N_B_c_159_n N_VGND_c_1132_n 0.00608558f $X=7.645 $Y=0.995 $X2=0 $Y2=0
cc_306 N_B_c_160_n N_VGND_c_1132_n 0.00746524f $X=8.165 $Y=0.995 $X2=0 $Y2=0
cc_307 N_B_c_157_n N_A_980_47#_c_1271_n 0.00864883f $X=6.705 $Y=0.995 $X2=0
+ $Y2=0
cc_308 N_B_c_197_p N_A_980_47#_c_1271_n 0.0058811f $X=6.27 $Y=1.175 $X2=0 $Y2=0
cc_309 N_B_c_161_n N_A_980_47#_c_1271_n 0.0340427f $X=8 $Y=1.16 $X2=0 $Y2=0
cc_310 N_B_c_157_n N_A_980_47#_c_1283_n 0.00644736f $X=6.705 $Y=0.995 $X2=0
+ $Y2=0
cc_311 N_B_c_158_n N_A_980_47#_c_1283_n 0.00686626f $X=7.175 $Y=0.995 $X2=0
+ $Y2=0
cc_312 N_B_c_159_n N_A_980_47#_c_1283_n 5.45498e-19 $X=7.645 $Y=0.995 $X2=0
+ $Y2=0
cc_313 N_B_c_158_n N_A_980_47#_c_1272_n 0.00901745f $X=7.175 $Y=0.995 $X2=0
+ $Y2=0
cc_314 N_B_c_159_n N_A_980_47#_c_1272_n 0.00901745f $X=7.645 $Y=0.995 $X2=0
+ $Y2=0
cc_315 N_B_c_161_n N_A_980_47#_c_1272_n 0.0397461f $X=8 $Y=1.16 $X2=0 $Y2=0
cc_316 N_B_c_163_n N_A_980_47#_c_1272_n 0.00345541f $X=8.14 $Y=1.202 $X2=0 $Y2=0
cc_317 N_B_c_158_n N_A_980_47#_c_1290_n 5.24597e-19 $X=7.175 $Y=0.995 $X2=0
+ $Y2=0
cc_318 N_B_c_159_n N_A_980_47#_c_1290_n 0.00651696f $X=7.645 $Y=0.995 $X2=0
+ $Y2=0
cc_319 N_B_c_160_n N_A_980_47#_c_1273_n 0.00866308f $X=8.165 $Y=0.995 $X2=0
+ $Y2=0
cc_320 N_B_c_160_n N_A_980_47#_c_1275_n 0.00276108f $X=8.165 $Y=0.995 $X2=0
+ $Y2=0
cc_321 N_B_c_173_n N_A_980_47#_c_1277_n 0.00490376f $X=6.1 $Y=1.53 $X2=0 $Y2=0
cc_322 N_B_c_197_p N_A_980_47#_c_1277_n 0.00763057f $X=6.27 $Y=1.175 $X2=0 $Y2=0
cc_323 N_B_c_157_n N_A_980_47#_c_1278_n 0.00116416f $X=6.705 $Y=0.995 $X2=0
+ $Y2=0
cc_324 N_B_c_158_n N_A_980_47#_c_1278_n 0.00116636f $X=7.175 $Y=0.995 $X2=0
+ $Y2=0
cc_325 N_B_c_161_n N_A_980_47#_c_1278_n 0.0298141f $X=8 $Y=1.16 $X2=0 $Y2=0
cc_326 N_B_c_163_n N_A_980_47#_c_1278_n 0.00358305f $X=8.14 $Y=1.202 $X2=0 $Y2=0
cc_327 N_B_c_159_n N_A_980_47#_c_1279_n 0.00119564f $X=7.645 $Y=0.995 $X2=0
+ $Y2=0
cc_328 N_B_c_160_n N_A_980_47#_c_1279_n 0.0048839f $X=8.165 $Y=0.995 $X2=0 $Y2=0
cc_329 N_B_c_161_n N_A_980_47#_c_1279_n 0.0377434f $X=8 $Y=1.16 $X2=0 $Y2=0
cc_330 N_B_c_163_n N_A_980_47#_c_1279_n 0.00486271f $X=8.14 $Y=1.202 $X2=0 $Y2=0
cc_331 N_A_c_367_n N_A_38_297#_c_561_n 0.0132364f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_332 N_A_c_368_n N_A_38_297#_c_561_n 0.0132364f $X=2.92 $Y=1.41 $X2=0 $Y2=0
cc_333 N_A_c_369_n N_A_38_297#_c_562_n 0.0132364f $X=3.39 $Y=1.41 $X2=0 $Y2=0
cc_334 N_A_c_370_n N_A_38_297#_c_562_n 0.0132364f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_335 N_A_c_374_n N_A_38_297#_c_530_n 0.00104198f $X=6.26 $Y=1.41 $X2=0 $Y2=0
cc_336 N_A_c_374_n N_A_38_297#_c_531_n 0.00236547f $X=6.26 $Y=1.41 $X2=0 $Y2=0
cc_337 N_A_c_365_n N_A_38_297#_c_531_n 0.0256707f $X=5.715 $Y=1.16 $X2=0 $Y2=0
cc_338 N_A_c_366_n N_A_38_297#_c_531_n 2.99086e-19 $X=6.26 $Y=1.202 $X2=0 $Y2=0
cc_339 N_A_c_374_n N_A_38_297#_c_533_n 3.28186e-19 $X=6.26 $Y=1.41 $X2=0 $Y2=0
cc_340 N_A_c_367_n N_VPWR_c_734_n 0.00300743f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_341 N_A_c_368_n N_VPWR_c_734_n 0.00300743f $X=2.92 $Y=1.41 $X2=0 $Y2=0
cc_342 N_A_c_369_n N_VPWR_c_735_n 0.00300743f $X=3.39 $Y=1.41 $X2=0 $Y2=0
cc_343 N_A_c_370_n N_VPWR_c_735_n 0.00300743f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_344 N_A_c_371_n N_VPWR_c_736_n 0.00300743f $X=4.85 $Y=1.41 $X2=0 $Y2=0
cc_345 N_A_c_372_n N_VPWR_c_736_n 0.00300743f $X=5.32 $Y=1.41 $X2=0 $Y2=0
cc_346 N_A_c_373_n N_VPWR_c_737_n 0.00300743f $X=5.79 $Y=1.41 $X2=0 $Y2=0
cc_347 N_A_c_374_n N_VPWR_c_737_n 0.00300743f $X=6.26 $Y=1.41 $X2=0 $Y2=0
cc_348 N_A_c_367_n N_VPWR_c_742_n 0.00523784f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_349 N_A_c_368_n N_VPWR_c_744_n 0.00523784f $X=2.92 $Y=1.41 $X2=0 $Y2=0
cc_350 N_A_c_369_n N_VPWR_c_744_n 0.00523784f $X=3.39 $Y=1.41 $X2=0 $Y2=0
cc_351 N_A_c_370_n N_VPWR_c_746_n 0.00523784f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_352 N_A_c_371_n N_VPWR_c_746_n 0.00523784f $X=4.85 $Y=1.41 $X2=0 $Y2=0
cc_353 N_A_c_372_n N_VPWR_c_748_n 0.00523784f $X=5.32 $Y=1.41 $X2=0 $Y2=0
cc_354 N_A_c_373_n N_VPWR_c_748_n 0.00523784f $X=5.79 $Y=1.41 $X2=0 $Y2=0
cc_355 N_A_c_374_n N_VPWR_c_750_n 0.00523784f $X=6.26 $Y=1.41 $X2=0 $Y2=0
cc_356 N_A_c_367_n N_VPWR_c_731_n 0.0068118f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_357 N_A_c_368_n N_VPWR_c_731_n 0.00678659f $X=2.92 $Y=1.41 $X2=0 $Y2=0
cc_358 N_A_c_369_n N_VPWR_c_731_n 0.00678659f $X=3.39 $Y=1.41 $X2=0 $Y2=0
cc_359 N_A_c_370_n N_VPWR_c_731_n 0.00806894f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_360 N_A_c_371_n N_VPWR_c_731_n 0.00806894f $X=4.85 $Y=1.41 $X2=0 $Y2=0
cc_361 N_A_c_372_n N_VPWR_c_731_n 0.00678659f $X=5.32 $Y=1.41 $X2=0 $Y2=0
cc_362 N_A_c_373_n N_VPWR_c_731_n 0.00678659f $X=5.79 $Y=1.41 $X2=0 $Y2=0
cc_363 N_A_c_374_n N_VPWR_c_731_n 0.0068118f $X=6.26 $Y=1.41 $X2=0 $Y2=0
cc_364 N_A_c_371_n N_A_898_297#_c_894_n 0.0132364f $X=4.85 $Y=1.41 $X2=0 $Y2=0
cc_365 N_A_c_372_n N_A_898_297#_c_894_n 0.0132364f $X=5.32 $Y=1.41 $X2=0 $Y2=0
cc_366 N_A_c_373_n N_A_898_297#_c_895_n 0.0131805f $X=5.79 $Y=1.41 $X2=0 $Y2=0
cc_367 N_A_c_374_n N_A_898_297#_c_895_n 0.0139861f $X=6.26 $Y=1.41 $X2=0 $Y2=0
cc_368 N_A_c_366_n N_A_898_297#_c_895_n 3.96083e-19 $X=6.26 $Y=1.202 $X2=0 $Y2=0
cc_369 N_A_c_356_n N_A_38_47#_c_1050_n 0.00282739f $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_370 N_A_c_356_n N_A_38_47#_c_1039_n 0.00540206f $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_371 N_A_c_357_n N_A_38_47#_c_1039_n 4.74935e-19 $X=2.895 $Y=0.995 $X2=0 $Y2=0
cc_372 N_A_c_365_n N_A_38_47#_c_1039_n 3.71806e-19 $X=5.715 $Y=1.16 $X2=0 $Y2=0
cc_373 N_A_c_356_n N_A_38_47#_c_1040_n 0.00901129f $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_374 N_A_c_357_n N_A_38_47#_c_1040_n 0.00895282f $X=2.895 $Y=0.995 $X2=0 $Y2=0
cc_375 N_A_c_364_n N_A_38_47#_c_1040_n 0.00345541f $X=3.86 $Y=1.202 $X2=0 $Y2=0
cc_376 N_A_c_365_n N_A_38_47#_c_1040_n 0.0385731f $X=5.715 $Y=1.16 $X2=0 $Y2=0
cc_377 N_A_c_356_n N_A_38_47#_c_1058_n 5.24597e-19 $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_378 N_A_c_357_n N_A_38_47#_c_1058_n 0.00651696f $X=2.895 $Y=0.995 $X2=0 $Y2=0
cc_379 N_A_c_358_n N_A_38_47#_c_1058_n 0.00693563f $X=3.365 $Y=0.995 $X2=0 $Y2=0
cc_380 N_A_c_359_n N_A_38_47#_c_1058_n 5.34196e-19 $X=3.885 $Y=0.995 $X2=0 $Y2=0
cc_381 N_A_c_358_n N_A_38_47#_c_1041_n 0.00928566f $X=3.365 $Y=0.995 $X2=0 $Y2=0
cc_382 N_A_c_359_n N_A_38_47#_c_1041_n 0.00935869f $X=3.885 $Y=0.995 $X2=0 $Y2=0
cc_383 N_A_c_364_n N_A_38_47#_c_1041_n 0.00468948f $X=3.86 $Y=1.202 $X2=0 $Y2=0
cc_384 N_A_c_365_n N_A_38_47#_c_1041_n 0.0694337f $X=5.715 $Y=1.16 $X2=0 $Y2=0
cc_385 N_A_c_358_n N_A_38_47#_c_1042_n 5.69266e-19 $X=3.365 $Y=0.995 $X2=0 $Y2=0
cc_386 N_A_c_359_n N_A_38_47#_c_1042_n 0.00857123f $X=3.885 $Y=0.995 $X2=0 $Y2=0
cc_387 N_A_c_357_n N_A_38_47#_c_1043_n 0.00116477f $X=2.895 $Y=0.995 $X2=0 $Y2=0
cc_388 N_A_c_358_n N_A_38_47#_c_1043_n 0.00116477f $X=3.365 $Y=0.995 $X2=0 $Y2=0
cc_389 N_A_c_364_n N_A_38_47#_c_1043_n 0.00358305f $X=3.86 $Y=1.202 $X2=0 $Y2=0
cc_390 N_A_c_365_n N_A_38_47#_c_1043_n 0.0296122f $X=5.715 $Y=1.16 $X2=0 $Y2=0
cc_391 N_A_c_356_n N_VGND_c_1110_n 0.00378935f $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_392 N_A_c_357_n N_VGND_c_1110_n 0.00276126f $X=2.895 $Y=0.995 $X2=0 $Y2=0
cc_393 N_A_c_358_n N_VGND_c_1111_n 0.00385467f $X=3.365 $Y=0.995 $X2=0 $Y2=0
cc_394 N_A_c_359_n N_VGND_c_1111_n 0.00365402f $X=3.885 $Y=0.995 $X2=0 $Y2=0
cc_395 N_A_c_359_n N_VGND_c_1112_n 0.00334802f $X=3.885 $Y=0.995 $X2=0 $Y2=0
cc_396 N_A_c_360_n N_VGND_c_1112_n 0.00496201f $X=4.825 $Y=0.995 $X2=0 $Y2=0
cc_397 N_A_c_365_n N_VGND_c_1112_n 0.0221752f $X=5.715 $Y=1.16 $X2=0 $Y2=0
cc_398 N_A_c_361_n N_VGND_c_1113_n 0.00379224f $X=5.295 $Y=0.995 $X2=0 $Y2=0
cc_399 N_A_c_362_n N_VGND_c_1113_n 0.00276126f $X=5.765 $Y=0.995 $X2=0 $Y2=0
cc_400 N_A_c_363_n N_VGND_c_1114_n 0.00268723f $X=6.285 $Y=0.995 $X2=0 $Y2=0
cc_401 N_A_c_356_n N_VGND_c_1117_n 0.00421816f $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_402 N_A_c_357_n N_VGND_c_1119_n 0.00423334f $X=2.895 $Y=0.995 $X2=0 $Y2=0
cc_403 N_A_c_358_n N_VGND_c_1119_n 0.00423334f $X=3.365 $Y=0.995 $X2=0 $Y2=0
cc_404 N_A_c_359_n N_VGND_c_1121_n 0.00396605f $X=3.885 $Y=0.995 $X2=0 $Y2=0
cc_405 N_A_c_360_n N_VGND_c_1123_n 0.00541359f $X=4.825 $Y=0.995 $X2=0 $Y2=0
cc_406 N_A_c_361_n N_VGND_c_1123_n 0.00423334f $X=5.295 $Y=0.995 $X2=0 $Y2=0
cc_407 N_A_c_362_n N_VGND_c_1125_n 0.00423334f $X=5.765 $Y=0.995 $X2=0 $Y2=0
cc_408 N_A_c_363_n N_VGND_c_1125_n 0.00437852f $X=6.285 $Y=0.995 $X2=0 $Y2=0
cc_409 N_A_c_356_n N_VGND_c_1132_n 0.00600232f $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_410 N_A_c_357_n N_VGND_c_1132_n 0.00597024f $X=2.895 $Y=0.995 $X2=0 $Y2=0
cc_411 N_A_c_358_n N_VGND_c_1132_n 0.00620835f $X=3.365 $Y=0.995 $X2=0 $Y2=0
cc_412 N_A_c_359_n N_VGND_c_1132_n 0.00712929f $X=3.885 $Y=0.995 $X2=0 $Y2=0
cc_413 N_A_c_360_n N_VGND_c_1132_n 0.0109546f $X=4.825 $Y=0.995 $X2=0 $Y2=0
cc_414 N_A_c_361_n N_VGND_c_1132_n 0.006093f $X=5.295 $Y=0.995 $X2=0 $Y2=0
cc_415 N_A_c_362_n N_VGND_c_1132_n 0.00608558f $X=5.765 $Y=0.995 $X2=0 $Y2=0
cc_416 N_A_c_363_n N_VGND_c_1132_n 0.00615622f $X=6.285 $Y=0.995 $X2=0 $Y2=0
cc_417 N_A_c_360_n N_A_980_47#_c_1304_n 0.00539651f $X=4.825 $Y=0.995 $X2=0
+ $Y2=0
cc_418 N_A_c_361_n N_A_980_47#_c_1304_n 0.00686626f $X=5.295 $Y=0.995 $X2=0
+ $Y2=0
cc_419 N_A_c_362_n N_A_980_47#_c_1304_n 5.45498e-19 $X=5.765 $Y=0.995 $X2=0
+ $Y2=0
cc_420 N_A_c_361_n N_A_980_47#_c_1269_n 0.00901129f $X=5.295 $Y=0.995 $X2=0
+ $Y2=0
cc_421 N_A_c_362_n N_A_980_47#_c_1269_n 0.00901129f $X=5.765 $Y=0.995 $X2=0
+ $Y2=0
cc_422 N_A_c_365_n N_A_980_47#_c_1269_n 0.0385731f $X=5.715 $Y=1.16 $X2=0 $Y2=0
cc_423 N_A_c_366_n N_A_980_47#_c_1269_n 0.00345541f $X=6.26 $Y=1.202 $X2=0 $Y2=0
cc_424 N_A_c_360_n N_A_980_47#_c_1270_n 0.00265998f $X=4.825 $Y=0.995 $X2=0
+ $Y2=0
cc_425 N_A_c_361_n N_A_980_47#_c_1270_n 0.00116477f $X=5.295 $Y=0.995 $X2=0
+ $Y2=0
cc_426 N_A_c_365_n N_A_980_47#_c_1270_n 0.0296122f $X=5.715 $Y=1.16 $X2=0 $Y2=0
cc_427 N_A_c_366_n N_A_980_47#_c_1270_n 0.00358305f $X=6.26 $Y=1.202 $X2=0 $Y2=0
cc_428 N_A_c_361_n N_A_980_47#_c_1315_n 5.24597e-19 $X=5.295 $Y=0.995 $X2=0
+ $Y2=0
cc_429 N_A_c_362_n N_A_980_47#_c_1315_n 0.00651696f $X=5.765 $Y=0.995 $X2=0
+ $Y2=0
cc_430 N_A_c_363_n N_A_980_47#_c_1271_n 0.0106048f $X=6.285 $Y=0.995 $X2=0 $Y2=0
cc_431 N_A_c_363_n N_A_980_47#_c_1283_n 5.32212e-19 $X=6.285 $Y=0.995 $X2=0
+ $Y2=0
cc_432 N_A_c_362_n N_A_980_47#_c_1277_n 0.00119406f $X=5.765 $Y=0.995 $X2=0
+ $Y2=0
cc_433 N_A_c_365_n N_A_980_47#_c_1277_n 0.00930562f $X=5.715 $Y=1.16 $X2=0 $Y2=0
cc_434 N_A_c_366_n N_A_980_47#_c_1277_n 0.00588858f $X=6.26 $Y=1.202 $X2=0 $Y2=0
cc_435 N_A_38_297#_c_525_n N_VPWR_M1005_s 0.00209407f $X=1.15 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_436 N_A_38_297#_c_555_n N_VPWR_M1016_s 0.00412184f $X=2.09 $Y=1.895 $X2=0
+ $Y2=0
cc_437 N_A_38_297#_c_531_n N_VPWR_M1016_s 0.00187762f $X=6.655 $Y=1.53 $X2=0
+ $Y2=0
cc_438 N_A_38_297#_c_561_n N_VPWR_M1015_s 0.00334944f $X=3.03 $Y=1.895 $X2=0
+ $Y2=0
cc_439 N_A_38_297#_c_562_n N_VPWR_M1027_s 0.00334944f $X=3.97 $Y=1.895 $X2=0
+ $Y2=0
cc_440 N_A_38_297#_c_525_n N_VPWR_c_732_n 0.0118222f $X=1.15 $Y=1.53 $X2=0 $Y2=0
cc_441 N_A_38_297#_c_555_n N_VPWR_c_733_n 0.0135607f $X=2.09 $Y=1.895 $X2=0
+ $Y2=0
cc_442 N_A_38_297#_c_561_n N_VPWR_c_734_n 0.0135607f $X=3.03 $Y=1.895 $X2=0
+ $Y2=0
cc_443 N_A_38_297#_c_562_n N_VPWR_c_735_n 0.0135607f $X=3.97 $Y=1.895 $X2=0
+ $Y2=0
cc_444 N_A_38_297#_c_519_n N_VPWR_c_738_n 0.00300743f $X=9.13 $Y=1.41 $X2=0
+ $Y2=0
cc_445 N_A_38_297#_c_520_n N_VPWR_c_738_n 0.00300743f $X=9.6 $Y=1.41 $X2=0 $Y2=0
cc_446 N_A_38_297#_c_521_n N_VPWR_c_739_n 0.00300743f $X=10.07 $Y=1.41 $X2=0
+ $Y2=0
cc_447 N_A_38_297#_c_522_n N_VPWR_c_739_n 0.00300743f $X=10.54 $Y=1.41 $X2=0
+ $Y2=0
cc_448 N_A_38_297#_c_555_n N_VPWR_c_740_n 0.0028084f $X=2.09 $Y=1.895 $X2=0
+ $Y2=0
cc_449 N_A_38_297#_c_618_p N_VPWR_c_740_n 0.0149311f $X=1.275 $Y=1.96 $X2=0
+ $Y2=0
cc_450 N_A_38_297#_c_555_n N_VPWR_c_742_n 0.0028084f $X=2.09 $Y=1.895 $X2=0
+ $Y2=0
cc_451 N_A_38_297#_c_561_n N_VPWR_c_742_n 0.0028084f $X=3.03 $Y=1.895 $X2=0
+ $Y2=0
cc_452 N_A_38_297#_c_567_n N_VPWR_c_742_n 0.0149311f $X=2.215 $Y=1.96 $X2=0
+ $Y2=0
cc_453 N_A_38_297#_c_561_n N_VPWR_c_744_n 0.0028084f $X=3.03 $Y=1.895 $X2=0
+ $Y2=0
cc_454 N_A_38_297#_c_562_n N_VPWR_c_744_n 0.0028084f $X=3.97 $Y=1.895 $X2=0
+ $Y2=0
cc_455 N_A_38_297#_c_568_n N_VPWR_c_744_n 0.0149311f $X=3.155 $Y=1.96 $X2=0
+ $Y2=0
cc_456 N_A_38_297#_c_562_n N_VPWR_c_746_n 0.0028084f $X=3.97 $Y=1.895 $X2=0
+ $Y2=0
cc_457 N_A_38_297#_c_529_n N_VPWR_c_746_n 0.0161853f $X=4.095 $Y=1.96 $X2=0
+ $Y2=0
cc_458 N_A_38_297#_c_519_n N_VPWR_c_750_n 0.00673617f $X=9.13 $Y=1.41 $X2=0
+ $Y2=0
cc_459 N_A_38_297#_c_520_n N_VPWR_c_752_n 0.00702461f $X=9.6 $Y=1.41 $X2=0 $Y2=0
cc_460 N_A_38_297#_c_521_n N_VPWR_c_752_n 0.00702461f $X=10.07 $Y=1.41 $X2=0
+ $Y2=0
cc_461 N_A_38_297#_c_522_n N_VPWR_c_754_n 0.00673617f $X=10.54 $Y=1.41 $X2=0
+ $Y2=0
cc_462 N_A_38_297#_M1005_d N_VPWR_c_731_n 0.00303344f $X=0.19 $Y=1.485 $X2=0
+ $Y2=0
cc_463 N_A_38_297#_M1012_d N_VPWR_c_731_n 0.00309052f $X=1.13 $Y=1.485 $X2=0
+ $Y2=0
cc_464 N_A_38_297#_M1034_d N_VPWR_c_731_n 0.0024798f $X=2.07 $Y=1.485 $X2=0
+ $Y2=0
cc_465 N_A_38_297#_M1019_d N_VPWR_c_731_n 0.0024798f $X=3.01 $Y=1.485 $X2=0
+ $Y2=0
cc_466 N_A_38_297#_M1035_d N_VPWR_c_731_n 0.00225074f $X=3.95 $Y=1.485 $X2=0
+ $Y2=0
cc_467 N_A_38_297#_c_519_n N_VPWR_c_731_n 0.0130258f $X=9.13 $Y=1.41 $X2=0 $Y2=0
cc_468 N_A_38_297#_c_520_n N_VPWR_c_731_n 0.0124092f $X=9.6 $Y=1.41 $X2=0 $Y2=0
cc_469 N_A_38_297#_c_521_n N_VPWR_c_731_n 0.0124092f $X=10.07 $Y=1.41 $X2=0
+ $Y2=0
cc_470 N_A_38_297#_c_522_n N_VPWR_c_731_n 0.0126595f $X=10.54 $Y=1.41 $X2=0
+ $Y2=0
cc_471 N_A_38_297#_c_524_n N_VPWR_c_731_n 0.0143649f $X=0.335 $Y=1.62 $X2=0
+ $Y2=0
cc_472 N_A_38_297#_c_555_n N_VPWR_c_731_n 0.0108264f $X=2.09 $Y=1.895 $X2=0
+ $Y2=0
cc_473 N_A_38_297#_c_561_n N_VPWR_c_731_n 0.0108264f $X=3.03 $Y=1.895 $X2=0
+ $Y2=0
cc_474 N_A_38_297#_c_562_n N_VPWR_c_731_n 0.0108264f $X=3.97 $Y=1.895 $X2=0
+ $Y2=0
cc_475 N_A_38_297#_c_618_p N_VPWR_c_731_n 0.00955092f $X=1.275 $Y=1.96 $X2=0
+ $Y2=0
cc_476 N_A_38_297#_c_567_n N_VPWR_c_731_n 0.00955092f $X=2.215 $Y=1.96 $X2=0
+ $Y2=0
cc_477 N_A_38_297#_c_568_n N_VPWR_c_731_n 0.00955092f $X=3.155 $Y=1.96 $X2=0
+ $Y2=0
cc_478 N_A_38_297#_c_529_n N_VPWR_c_731_n 0.00955092f $X=4.095 $Y=1.96 $X2=0
+ $Y2=0
cc_479 N_A_38_297#_c_524_n N_VPWR_c_756_n 0.0251183f $X=0.335 $Y=1.62 $X2=0
+ $Y2=0
cc_480 N_A_38_297#_c_530_n N_A_898_297#_M1026_s 0.00178541f $X=8.39 $Y=1.53
+ $X2=0 $Y2=0
cc_481 N_A_38_297#_c_531_n N_A_898_297#_M1026_s 0.00119963f $X=6.655 $Y=1.53
+ $X2=0 $Y2=0
cc_482 N_A_38_297#_c_530_n N_A_898_297#_M1020_s 0.00187547f $X=8.39 $Y=1.53
+ $X2=0 $Y2=0
cc_483 N_A_38_297#_c_530_n N_A_898_297#_M1036_s 0.00294625f $X=8.39 $Y=1.53
+ $X2=0 $Y2=0
cc_484 N_A_38_297#_c_531_n N_A_898_297#_c_894_n 0.00508579f $X=6.655 $Y=1.53
+ $X2=0 $Y2=0
cc_485 N_A_38_297#_c_531_n N_A_898_297#_c_895_n 0.00692627f $X=6.655 $Y=1.53
+ $X2=0 $Y2=0
cc_486 N_A_38_297#_c_530_n N_A_898_297#_c_897_n 0.00658644f $X=8.39 $Y=1.53
+ $X2=0 $Y2=0
cc_487 N_A_38_297#_c_531_n N_A_898_297#_c_897_n 0.00456848f $X=6.655 $Y=1.53
+ $X2=0 $Y2=0
cc_488 N_A_38_297#_c_530_n N_A_898_297#_c_890_n 0.00151294f $X=8.39 $Y=1.53
+ $X2=0 $Y2=0
cc_489 N_A_38_297#_c_531_n N_A_898_297#_c_890_n 4.5081e-19 $X=6.655 $Y=1.53
+ $X2=0 $Y2=0
cc_490 N_A_38_297#_c_533_n N_A_898_297#_c_890_n 0.0020154f $X=6.81 $Y=1.53 $X2=0
+ $Y2=0
cc_491 N_A_38_297#_c_529_n N_A_898_297#_c_891_n 0.0496599f $X=4.095 $Y=1.96
+ $X2=0 $Y2=0
cc_492 N_A_38_297#_c_531_n N_A_898_297#_c_891_n 0.00264177f $X=6.655 $Y=1.53
+ $X2=0 $Y2=0
cc_493 N_A_38_297#_c_531_n N_A_898_297#_c_903_n 0.00209664f $X=6.655 $Y=1.53
+ $X2=0 $Y2=0
cc_494 N_A_38_297#_c_530_n N_Y_M1006_d 0.00111833f $X=8.39 $Y=1.53 $X2=0 $Y2=0
cc_495 N_A_38_297#_c_533_n N_Y_M1006_d 0.00201962f $X=6.81 $Y=1.53 $X2=0 $Y2=0
cc_496 N_A_38_297#_c_530_n N_Y_M1028_d 0.00187547f $X=8.39 $Y=1.53 $X2=0 $Y2=0
cc_497 N_A_38_297#_c_517_n N_Y_c_956_n 0.00624078f $X=10.37 $Y=1.16 $X2=0 $Y2=0
cc_498 N_A_38_297#_c_530_n N_Y_c_956_n 0.103198f $X=8.39 $Y=1.53 $X2=0 $Y2=0
cc_499 N_A_38_297#_c_533_n N_Y_c_956_n 0.00700584f $X=6.81 $Y=1.53 $X2=0 $Y2=0
cc_500 N_A_38_297#_c_519_n N_Y_c_957_n 0.00465871f $X=9.13 $Y=1.41 $X2=0 $Y2=0
cc_501 N_A_38_297#_c_519_n N_Y_c_958_n 0.0161605f $X=9.13 $Y=1.41 $X2=0 $Y2=0
cc_502 N_A_38_297#_c_520_n N_Y_c_958_n 0.0174772f $X=9.6 $Y=1.41 $X2=0 $Y2=0
cc_503 N_A_38_297#_c_517_n N_Y_c_958_n 0.0466668f $X=10.37 $Y=1.16 $X2=0 $Y2=0
cc_504 N_A_38_297#_c_518_n N_Y_c_958_n 0.00821262f $X=10.54 $Y=1.202 $X2=0 $Y2=0
cc_505 N_A_38_297#_c_508_n N_Y_c_954_n 0.00380374f $X=9.105 $Y=0.995 $X2=0 $Y2=0
cc_506 N_A_38_297#_c_509_n N_Y_c_954_n 0.0112301f $X=9.575 $Y=0.995 $X2=0 $Y2=0
cc_507 N_A_38_297#_c_510_n N_Y_c_954_n 0.0112578f $X=10.045 $Y=0.995 $X2=0 $Y2=0
cc_508 N_A_38_297#_c_511_n N_Y_c_954_n 0.0140989f $X=10.565 $Y=0.995 $X2=0 $Y2=0
cc_509 N_A_38_297#_c_517_n N_Y_c_954_n 0.101919f $X=10.37 $Y=1.16 $X2=0 $Y2=0
cc_510 N_A_38_297#_c_518_n N_Y_c_954_n 0.0116969f $X=10.54 $Y=1.202 $X2=0 $Y2=0
cc_511 N_A_38_297#_c_521_n N_Y_c_959_n 0.0174772f $X=10.07 $Y=1.41 $X2=0 $Y2=0
cc_512 N_A_38_297#_c_522_n N_Y_c_959_n 0.0162261f $X=10.54 $Y=1.41 $X2=0 $Y2=0
cc_513 N_A_38_297#_c_517_n N_Y_c_959_n 0.0414161f $X=10.37 $Y=1.16 $X2=0 $Y2=0
cc_514 N_A_38_297#_c_518_n N_Y_c_959_n 0.00800464f $X=10.54 $Y=1.202 $X2=0 $Y2=0
cc_515 N_A_38_297#_c_521_n N_Y_c_960_n 6.07675e-19 $X=10.07 $Y=1.41 $X2=0 $Y2=0
cc_516 N_A_38_297#_c_522_n N_Y_c_960_n 0.0102674f $X=10.54 $Y=1.41 $X2=0 $Y2=0
cc_517 N_A_38_297#_c_519_n N_Y_c_961_n 0.00772277f $X=9.13 $Y=1.41 $X2=0 $Y2=0
cc_518 N_A_38_297#_c_520_n N_Y_c_961_n 7.03686e-19 $X=9.6 $Y=1.41 $X2=0 $Y2=0
cc_519 N_A_38_297#_c_517_n N_Y_c_961_n 0.0278154f $X=10.37 $Y=1.16 $X2=0 $Y2=0
cc_520 N_A_38_297#_c_530_n N_Y_c_961_n 0.0150382f $X=8.39 $Y=1.53 $X2=0 $Y2=0
cc_521 N_A_38_297#_c_518_n N_Y_c_961_n 3.20658e-19 $X=10.54 $Y=1.202 $X2=0 $Y2=0
cc_522 N_A_38_297#_c_517_n N_Y_c_962_n 0.020385f $X=10.37 $Y=1.16 $X2=0 $Y2=0
cc_523 N_A_38_297#_c_518_n N_Y_c_962_n 0.00664519f $X=10.54 $Y=1.202 $X2=0 $Y2=0
cc_524 N_A_38_297#_c_522_n N_Y_c_963_n 0.00168966f $X=10.54 $Y=1.41 $X2=0 $Y2=0
cc_525 N_A_38_297#_c_518_n N_Y_c_963_n 3.89106e-19 $X=10.54 $Y=1.202 $X2=0 $Y2=0
cc_526 N_A_38_297#_c_522_n Y 0.00136862f $X=10.54 $Y=1.41 $X2=0 $Y2=0
cc_527 N_A_38_297#_c_511_n Y 0.0193348f $X=10.565 $Y=0.995 $X2=0 $Y2=0
cc_528 N_A_38_297#_c_517_n Y 0.0161986f $X=10.37 $Y=1.16 $X2=0 $Y2=0
cc_529 N_A_38_297#_c_513_n N_A_38_47#_M1007_s 0.00271814f $X=0.32 $Y=0.775
+ $X2=-0.19 $Y2=-0.24
cc_530 N_A_38_297#_c_514_n N_A_38_47#_M1007_s 9.57256e-19 $X=1.745 $Y=0.73
+ $X2=-0.19 $Y2=-0.24
cc_531 N_A_38_297#_c_514_n N_A_38_47#_M1021_s 0.00214342f $X=1.745 $Y=0.73 $X2=0
+ $Y2=0
cc_532 N_A_38_297#_M1007_d N_A_38_47#_c_1038_n 0.00400389f $X=0.62 $Y=0.235
+ $X2=0 $Y2=0
cc_533 N_A_38_297#_M1037_d N_A_38_47#_c_1038_n 0.00507817f $X=1.56 $Y=0.235
+ $X2=0 $Y2=0
cc_534 N_A_38_297#_c_513_n N_A_38_47#_c_1038_n 0.011822f $X=0.32 $Y=0.775 $X2=0
+ $Y2=0
cc_535 N_A_38_297#_c_514_n N_A_38_47#_c_1038_n 0.085575f $X=1.745 $Y=0.73 $X2=0
+ $Y2=0
cc_536 N_A_38_297#_c_514_n N_A_38_47#_c_1039_n 0.00140356f $X=1.745 $Y=0.73
+ $X2=0 $Y2=0
cc_537 N_A_38_297#_c_531_n N_A_38_47#_c_1039_n 0.00185567f $X=6.655 $Y=1.53
+ $X2=0 $Y2=0
cc_538 N_A_38_297#_c_508_n N_VGND_c_1116_n 0.00251964f $X=9.105 $Y=0.995 $X2=0
+ $Y2=0
cc_539 N_A_38_297#_c_513_n N_VGND_c_1117_n 0.00169073f $X=0.32 $Y=0.775 $X2=0
+ $Y2=0
cc_540 N_A_38_297#_c_508_n N_VGND_c_1131_n 0.00368123f $X=9.105 $Y=0.995 $X2=0
+ $Y2=0
cc_541 N_A_38_297#_c_509_n N_VGND_c_1131_n 0.00368123f $X=9.575 $Y=0.995 $X2=0
+ $Y2=0
cc_542 N_A_38_297#_c_510_n N_VGND_c_1131_n 0.00368123f $X=10.045 $Y=0.995 $X2=0
+ $Y2=0
cc_543 N_A_38_297#_c_511_n N_VGND_c_1131_n 0.00368123f $X=10.565 $Y=0.995 $X2=0
+ $Y2=0
cc_544 N_A_38_297#_M1007_d N_VGND_c_1132_n 0.00256987f $X=0.62 $Y=0.235 $X2=0
+ $Y2=0
cc_545 N_A_38_297#_M1037_d N_VGND_c_1132_n 0.00297142f $X=1.56 $Y=0.235 $X2=0
+ $Y2=0
cc_546 N_A_38_297#_c_508_n N_VGND_c_1132_n 0.00670426f $X=9.105 $Y=0.995 $X2=0
+ $Y2=0
cc_547 N_A_38_297#_c_509_n N_VGND_c_1132_n 0.00550516f $X=9.575 $Y=0.995 $X2=0
+ $Y2=0
cc_548 N_A_38_297#_c_510_n N_VGND_c_1132_n 0.00562494f $X=10.045 $Y=0.995 $X2=0
+ $Y2=0
cc_549 N_A_38_297#_c_511_n N_VGND_c_1132_n 0.00645695f $X=10.565 $Y=0.995 $X2=0
+ $Y2=0
cc_550 N_A_38_297#_c_513_n N_VGND_c_1132_n 0.00291453f $X=0.32 $Y=0.775 $X2=0
+ $Y2=0
cc_551 N_A_38_297#_c_531_n N_A_980_47#_c_1271_n 2.6706e-19 $X=6.655 $Y=1.53
+ $X2=0 $Y2=0
cc_552 N_A_38_297#_c_508_n N_A_980_47#_c_1273_n 4.83058e-19 $X=9.105 $Y=0.995
+ $X2=0 $Y2=0
cc_553 N_A_38_297#_c_516_n N_A_980_47#_c_1273_n 0.0140881f $X=8.56 $Y=1.175
+ $X2=0 $Y2=0
cc_554 N_A_38_297#_c_517_n N_A_980_47#_c_1273_n 0.0340191f $X=10.37 $Y=1.16
+ $X2=0 $Y2=0
cc_555 N_A_38_297#_c_530_n N_A_980_47#_c_1273_n 0.00691542f $X=8.39 $Y=1.53
+ $X2=0 $Y2=0
cc_556 N_A_38_297#_c_508_n N_A_980_47#_c_1276_n 0.00988409f $X=9.105 $Y=0.995
+ $X2=0 $Y2=0
cc_557 N_A_38_297#_c_509_n N_A_980_47#_c_1276_n 0.0083138f $X=9.575 $Y=0.995
+ $X2=0 $Y2=0
cc_558 N_A_38_297#_c_510_n N_A_980_47#_c_1276_n 0.00857276f $X=10.045 $Y=0.995
+ $X2=0 $Y2=0
cc_559 N_A_38_297#_c_511_n N_A_980_47#_c_1276_n 0.00857276f $X=10.565 $Y=0.995
+ $X2=0 $Y2=0
cc_560 N_A_38_297#_c_517_n N_A_980_47#_c_1276_n 0.00369351f $X=10.37 $Y=1.16
+ $X2=0 $Y2=0
cc_561 N_A_38_297#_c_531_n N_A_980_47#_c_1277_n 0.00188301f $X=6.655 $Y=1.53
+ $X2=0 $Y2=0
cc_562 N_VPWR_c_731_n N_A_898_297#_M1000_s 0.00225877f $X=10.81 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_563 N_VPWR_c_731_n N_A_898_297#_M1013_s 0.0024798f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_564 N_VPWR_c_731_n N_A_898_297#_M1026_s 0.00240429f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_565 N_VPWR_c_731_n N_A_898_297#_M1020_s 0.00231289f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_566 N_VPWR_c_731_n N_A_898_297#_M1036_s 0.00217543f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_567 N_VPWR_M1000_d N_A_898_297#_c_894_n 0.00334944f $X=4.94 $Y=1.485 $X2=0
+ $Y2=0
cc_568 N_VPWR_c_736_n N_A_898_297#_c_894_n 0.0135607f $X=5.085 $Y=2.34 $X2=0
+ $Y2=0
cc_569 N_VPWR_c_746_n N_A_898_297#_c_894_n 0.0028084f $X=4.96 $Y=2.72 $X2=0
+ $Y2=0
cc_570 N_VPWR_c_748_n N_A_898_297#_c_894_n 0.0028084f $X=5.9 $Y=2.72 $X2=0 $Y2=0
cc_571 N_VPWR_c_731_n N_A_898_297#_c_894_n 0.0108264f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_572 N_VPWR_M1018_d N_A_898_297#_c_895_n 0.00334064f $X=5.88 $Y=1.485 $X2=0
+ $Y2=0
cc_573 N_VPWR_c_737_n N_A_898_297#_c_895_n 0.0135607f $X=6.025 $Y=2.34 $X2=0
+ $Y2=0
cc_574 N_VPWR_c_748_n N_A_898_297#_c_895_n 0.0028084f $X=5.9 $Y=2.72 $X2=0 $Y2=0
cc_575 N_VPWR_c_750_n N_A_898_297#_c_895_n 0.0028084f $X=9.24 $Y=2.72 $X2=0
+ $Y2=0
cc_576 N_VPWR_c_731_n N_A_898_297#_c_895_n 0.0108264f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_577 N_VPWR_c_750_n N_A_898_297#_c_938_n 0.0134783f $X=9.24 $Y=2.72 $X2=0
+ $Y2=0
cc_578 N_VPWR_c_731_n N_A_898_297#_c_938_n 0.00808747f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_579 N_VPWR_c_750_n N_A_898_297#_c_890_n 0.112383f $X=9.24 $Y=2.72 $X2=0 $Y2=0
cc_580 N_VPWR_c_731_n N_A_898_297#_c_890_n 0.07004f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_581 N_VPWR_c_746_n N_A_898_297#_c_891_n 0.0208441f $X=4.96 $Y=2.72 $X2=0
+ $Y2=0
cc_582 N_VPWR_c_731_n N_A_898_297#_c_891_n 0.0120542f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_583 N_VPWR_c_748_n N_A_898_297#_c_903_n 0.0149311f $X=5.9 $Y=2.72 $X2=0 $Y2=0
cc_584 N_VPWR_c_731_n N_A_898_297#_c_903_n 0.00955092f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_585 N_VPWR_c_731_n N_Y_M1006_d 0.00232895f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_586 N_VPWR_c_731_n N_Y_M1028_d 0.00232895f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_587 N_VPWR_c_731_n N_Y_M1001_d 0.00217517f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_588 N_VPWR_c_731_n N_Y_M1008_d 0.00370124f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_589 N_VPWR_c_731_n N_Y_M1029_d 0.00217517f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_590 N_VPWR_c_750_n N_Y_c_956_n 0.00329726f $X=9.24 $Y=2.72 $X2=0 $Y2=0
cc_591 N_VPWR_c_731_n N_Y_c_956_n 0.00861215f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_592 N_VPWR_c_750_n N_Y_c_957_n 0.0210596f $X=9.24 $Y=2.72 $X2=0 $Y2=0
cc_593 N_VPWR_c_731_n N_Y_c_957_n 0.0124725f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_594 N_VPWR_M1001_s N_Y_c_958_n 0.00188585f $X=9.22 $Y=1.485 $X2=0 $Y2=0
cc_595 N_VPWR_c_738_n N_Y_c_958_n 0.014572f $X=9.365 $Y=2 $X2=0 $Y2=0
cc_596 N_VPWR_c_752_n N_Y_c_1016_n 0.0149311f $X=10.18 $Y=2.72 $X2=0 $Y2=0
cc_597 N_VPWR_c_731_n N_Y_c_1016_n 0.00955092f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_598 N_VPWR_M1017_s N_Y_c_959_n 0.00188585f $X=10.16 $Y=1.485 $X2=0 $Y2=0
cc_599 N_VPWR_c_739_n N_Y_c_959_n 0.014572f $X=10.305 $Y=2 $X2=0 $Y2=0
cc_600 N_VPWR_c_754_n N_Y_c_960_n 0.0210596f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_601 N_VPWR_c_731_n N_Y_c_960_n 0.0124725f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_602 N_A_898_297#_c_890_n N_Y_M1006_d 0.00354918f $X=8.375 $Y=2.3 $X2=0 $Y2=0
cc_603 N_A_898_297#_c_890_n N_Y_M1028_d 0.00357068f $X=8.375 $Y=2.3 $X2=0 $Y2=0
cc_604 N_A_898_297#_M1020_s N_Y_c_956_n 0.00350737f $X=7.29 $Y=1.485 $X2=0 $Y2=0
cc_605 N_A_898_297#_M1036_s N_Y_c_956_n 0.0058096f $X=8.23 $Y=1.485 $X2=0 $Y2=0
cc_606 N_A_898_297#_c_897_n N_Y_c_956_n 0.0191412f $X=6.475 $Y=2.005 $X2=0 $Y2=0
cc_607 N_A_898_297#_c_938_n N_Y_c_956_n 0.00307345f $X=6.475 $Y=2.215 $X2=0
+ $Y2=0
cc_608 N_A_898_297#_c_890_n N_Y_c_956_n 0.0990854f $X=8.375 $Y=2.3 $X2=0 $Y2=0
cc_609 N_A_898_297#_c_890_n N_Y_c_957_n 0.0202777f $X=8.375 $Y=2.3 $X2=0 $Y2=0
cc_610 N_Y_M1003_s N_VGND_c_1132_n 0.00261035f $X=9.18 $Y=0.235 $X2=0 $Y2=0
cc_611 N_Y_M1014_s N_VGND_c_1132_n 0.00301822f $X=10.12 $Y=0.235 $X2=0 $Y2=0
cc_612 N_Y_c_954_n N_A_980_47#_M1010_d 0.00219446f $X=10.705 $Y=0.78 $X2=0 $Y2=0
cc_613 N_Y_c_954_n N_A_980_47#_M1024_d 0.00323022f $X=10.705 $Y=0.78 $X2=0 $Y2=0
cc_614 N_Y_c_954_n N_A_980_47#_c_1273_n 0.00799569f $X=10.705 $Y=0.78 $X2=0
+ $Y2=0
cc_615 N_Y_M1003_s N_A_980_47#_c_1276_n 0.00423532f $X=9.18 $Y=0.235 $X2=0 $Y2=0
cc_616 N_Y_M1014_s N_A_980_47#_c_1276_n 0.00533758f $X=10.12 $Y=0.235 $X2=0
+ $Y2=0
cc_617 N_Y_c_954_n N_A_980_47#_c_1276_n 0.0930856f $X=10.705 $Y=0.78 $X2=0 $Y2=0
cc_618 N_A_38_47#_c_1040_n N_VGND_M1009_s 0.00251047f $X=2.94 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_619 N_A_38_47#_c_1041_n N_VGND_M1031_s 0.00348805f $X=3.88 $Y=0.815 $X2=0
+ $Y2=0
cc_620 N_A_38_47#_c_1050_n N_VGND_c_1110_n 0.0141571f $X=2.255 $Y=0.475 $X2=0
+ $Y2=0
cc_621 N_A_38_47#_c_1039_n N_VGND_c_1110_n 0.00471242f $X=2.255 $Y=0.725 $X2=0
+ $Y2=0
cc_622 N_A_38_47#_c_1040_n N_VGND_c_1110_n 0.0127273f $X=2.94 $Y=0.815 $X2=0
+ $Y2=0
cc_623 N_A_38_47#_c_1058_n N_VGND_c_1111_n 0.0183628f $X=3.155 $Y=0.39 $X2=0
+ $Y2=0
cc_624 N_A_38_47#_c_1041_n N_VGND_c_1111_n 0.0131987f $X=3.88 $Y=0.815 $X2=0
+ $Y2=0
cc_625 N_A_38_47#_c_1042_n N_VGND_c_1111_n 0.0223967f $X=4.095 $Y=0.39 $X2=0
+ $Y2=0
cc_626 N_A_38_47#_c_1041_n N_VGND_c_1112_n 0.0156976f $X=3.88 $Y=0.815 $X2=0
+ $Y2=0
cc_627 N_A_38_47#_c_1042_n N_VGND_c_1112_n 0.03893f $X=4.095 $Y=0.39 $X2=0 $Y2=0
cc_628 N_A_38_47#_c_1038_n N_VGND_c_1117_n 0.112055f $X=2.13 $Y=0.365 $X2=0
+ $Y2=0
cc_629 N_A_38_47#_c_1050_n N_VGND_c_1117_n 0.0152108f $X=2.255 $Y=0.475 $X2=0
+ $Y2=0
cc_630 N_A_38_47#_c_1040_n N_VGND_c_1117_n 0.00266636f $X=2.94 $Y=0.815 $X2=0
+ $Y2=0
cc_631 N_A_38_47#_c_1040_n N_VGND_c_1119_n 0.00198695f $X=2.94 $Y=0.815 $X2=0
+ $Y2=0
cc_632 N_A_38_47#_c_1058_n N_VGND_c_1119_n 0.0223596f $X=3.155 $Y=0.39 $X2=0
+ $Y2=0
cc_633 N_A_38_47#_c_1041_n N_VGND_c_1119_n 0.00266636f $X=3.88 $Y=0.815 $X2=0
+ $Y2=0
cc_634 N_A_38_47#_c_1041_n N_VGND_c_1121_n 0.00199443f $X=3.88 $Y=0.815 $X2=0
+ $Y2=0
cc_635 N_A_38_47#_c_1042_n N_VGND_c_1121_n 0.024373f $X=4.095 $Y=0.39 $X2=0
+ $Y2=0
cc_636 N_A_38_47#_M1007_s N_VGND_c_1132_n 0.00225742f $X=0.19 $Y=0.235 $X2=0
+ $Y2=0
cc_637 N_A_38_47#_M1021_s N_VGND_c_1132_n 0.00255381f $X=1.09 $Y=0.235 $X2=0
+ $Y2=0
cc_638 N_A_38_47#_M1038_s N_VGND_c_1132_n 0.00215206f $X=2.08 $Y=0.235 $X2=0
+ $Y2=0
cc_639 N_A_38_47#_M1030_d N_VGND_c_1132_n 0.0025535f $X=2.97 $Y=0.235 $X2=0
+ $Y2=0
cc_640 N_A_38_47#_M1032_d N_VGND_c_1132_n 0.00209319f $X=3.96 $Y=0.235 $X2=0
+ $Y2=0
cc_641 N_A_38_47#_c_1038_n N_VGND_c_1132_n 0.0703895f $X=2.13 $Y=0.365 $X2=0
+ $Y2=0
cc_642 N_A_38_47#_c_1050_n N_VGND_c_1132_n 0.00940698f $X=2.255 $Y=0.475 $X2=0
+ $Y2=0
cc_643 N_A_38_47#_c_1040_n N_VGND_c_1132_n 0.00972452f $X=2.94 $Y=0.815 $X2=0
+ $Y2=0
cc_644 N_A_38_47#_c_1058_n N_VGND_c_1132_n 0.0141302f $X=3.155 $Y=0.39 $X2=0
+ $Y2=0
cc_645 N_A_38_47#_c_1041_n N_VGND_c_1132_n 0.0100158f $X=3.88 $Y=0.815 $X2=0
+ $Y2=0
cc_646 N_A_38_47#_c_1042_n N_VGND_c_1132_n 0.0141066f $X=4.095 $Y=0.39 $X2=0
+ $Y2=0
cc_647 N_VGND_c_1132_n N_A_980_47#_M1004_s 0.0025535f $X=10.81 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_648 N_VGND_c_1132_n N_A_980_47#_M1025_s 0.00304143f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_649 N_VGND_c_1132_n N_A_980_47#_M1002_s 0.0025535f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_650 N_VGND_c_1132_n N_A_980_47#_M1023_s 0.00304114f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_651 N_VGND_c_1132_n N_A_980_47#_M1003_d 0.00212536f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_652 N_VGND_c_1132_n N_A_980_47#_M1010_d 0.00259403f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_653 N_VGND_c_1132_n N_A_980_47#_M1024_d 0.0021262f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_654 N_VGND_c_1113_n N_A_980_47#_c_1304_n 0.0183628f $X=5.555 $Y=0.39 $X2=0
+ $Y2=0
cc_655 N_VGND_c_1123_n N_A_980_47#_c_1304_n 0.0223596f $X=5.47 $Y=0 $X2=0 $Y2=0
cc_656 N_VGND_c_1132_n N_A_980_47#_c_1304_n 0.0141302f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_657 N_VGND_M1022_d N_A_980_47#_c_1269_n 0.00251047f $X=5.37 $Y=0.235 $X2=0
+ $Y2=0
cc_658 N_VGND_c_1113_n N_A_980_47#_c_1269_n 0.0127273f $X=5.555 $Y=0.39 $X2=0
+ $Y2=0
cc_659 N_VGND_c_1123_n N_A_980_47#_c_1269_n 0.00266636f $X=5.47 $Y=0 $X2=0 $Y2=0
cc_660 N_VGND_c_1125_n N_A_980_47#_c_1269_n 0.00198695f $X=6.41 $Y=0 $X2=0 $Y2=0
cc_661 N_VGND_c_1132_n N_A_980_47#_c_1269_n 0.00972452f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_662 N_VGND_c_1112_n N_A_980_47#_c_1270_n 0.00835241f $X=4.615 $Y=0.39 $X2=0
+ $Y2=0
cc_663 N_VGND_c_1125_n N_A_980_47#_c_1315_n 0.0231806f $X=6.41 $Y=0 $X2=0 $Y2=0
cc_664 N_VGND_c_1132_n N_A_980_47#_c_1315_n 0.0143352f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_665 N_VGND_M1033_d N_A_980_47#_c_1271_n 0.00162089f $X=6.36 $Y=0.235 $X2=0
+ $Y2=0
cc_666 N_VGND_c_1114_n N_A_980_47#_c_1271_n 0.0122559f $X=6.495 $Y=0.39 $X2=0
+ $Y2=0
cc_667 N_VGND_c_1125_n N_A_980_47#_c_1271_n 0.00254521f $X=6.41 $Y=0 $X2=0 $Y2=0
cc_668 N_VGND_c_1127_n N_A_980_47#_c_1271_n 0.00198695f $X=7.35 $Y=0 $X2=0 $Y2=0
cc_669 N_VGND_c_1132_n N_A_980_47#_c_1271_n 0.0094839f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_670 N_VGND_c_1115_n N_A_980_47#_c_1283_n 0.0183628f $X=7.435 $Y=0.39 $X2=0
+ $Y2=0
cc_671 N_VGND_c_1127_n N_A_980_47#_c_1283_n 0.0223596f $X=7.35 $Y=0 $X2=0 $Y2=0
cc_672 N_VGND_c_1132_n N_A_980_47#_c_1283_n 0.0141302f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_673 N_VGND_M1011_d N_A_980_47#_c_1272_n 0.00251047f $X=7.25 $Y=0.235 $X2=0
+ $Y2=0
cc_674 N_VGND_c_1115_n N_A_980_47#_c_1272_n 0.0127273f $X=7.435 $Y=0.39 $X2=0
+ $Y2=0
cc_675 N_VGND_c_1127_n N_A_980_47#_c_1272_n 0.00266636f $X=7.35 $Y=0 $X2=0 $Y2=0
cc_676 N_VGND_c_1129_n N_A_980_47#_c_1272_n 0.00198695f $X=8.29 $Y=0 $X2=0 $Y2=0
cc_677 N_VGND_c_1132_n N_A_980_47#_c_1272_n 0.00972452f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_678 N_VGND_c_1129_n N_A_980_47#_c_1290_n 0.0231806f $X=8.29 $Y=0 $X2=0 $Y2=0
cc_679 N_VGND_c_1132_n N_A_980_47#_c_1290_n 0.0143352f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_680 N_VGND_M1039_d N_A_980_47#_c_1273_n 0.00315719f $X=8.24 $Y=0.235 $X2=0
+ $Y2=0
cc_681 N_VGND_c_1116_n N_A_980_47#_c_1273_n 0.012101f $X=8.375 $Y=0.39 $X2=0
+ $Y2=0
cc_682 N_VGND_c_1129_n N_A_980_47#_c_1273_n 0.00128233f $X=8.29 $Y=0 $X2=0 $Y2=0
cc_683 N_VGND_c_1131_n N_A_980_47#_c_1273_n 0.00399176f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_684 N_VGND_c_1132_n N_A_980_47#_c_1273_n 0.0105081f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_685 N_VGND_c_1116_n N_A_980_47#_c_1274_n 0.0101441f $X=8.375 $Y=0.39 $X2=0
+ $Y2=0
cc_686 N_VGND_c_1131_n N_A_980_47#_c_1274_n 0.0130441f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_687 N_VGND_c_1132_n N_A_980_47#_c_1274_n 0.00935125f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_688 N_VGND_c_1116_n N_A_980_47#_c_1275_n 0.00435313f $X=8.375 $Y=0.39 $X2=0
+ $Y2=0
cc_689 N_VGND_c_1131_n N_A_980_47#_c_1276_n 0.0839473f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_690 N_VGND_c_1132_n N_A_980_47#_c_1276_n 0.0676908f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_691 N_VGND_c_1129_n N_A_980_47#_c_1279_n 0.00122796f $X=8.29 $Y=0 $X2=0 $Y2=0
cc_692 N_VGND_c_1132_n N_A_980_47#_c_1279_n 0.00220472f $X=10.81 $Y=0 $X2=0
+ $Y2=0
