* File: sky130_fd_sc_hdll__a21o_4.spice
* Created: Thu Aug 27 18:52:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a21o_4.pex.spice"
.subckt sky130_fd_sc_hdll__a21o_4  VNB VPB B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1002 N_X_M1002_d N_A_84_21#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.18525 PD=0.98 PS=1.87 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75005 A=0.0975 P=1.6 MULT=1
MM1005 N_X_M1002_d N_A_84_21#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75000.7
+ SB=75004.6 A=0.0975 P=1.6 MULT=1
MM1008 N_X_M1008_d N_A_84_21#_M1008_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1016 N_X_M1008_d N_A_84_21#_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.281125 PD=0.98 PS=1.515 NRD=0 NRS=29.532 M=1 R=4.33333
+ SA=75001.6 SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1016_s N_B1_M1000_g N_A_84_21#_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.281125 AS=0.12025 PD=1.515 PS=1.02 NRD=2.76 NRS=8.304 M=1 R=4.33333
+ SA=75002.7 SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_B1_M1006_g N_A_84_21#_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10075 AS=0.12025 PD=0.96 PS=1.02 NRD=6.456 NRS=8.304 M=1 R=4.33333
+ SA=75003.2 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1006_d N_A2_M1007_g A_801_47# VNB NSHORT L=0.15 W=0.65 AD=0.10075
+ AS=0.091 PD=0.96 PS=0.93 NRD=0 NRS=15.684 M=1 R=4.33333 SA=75003.6 SB=75001.6
+ A=0.0975 P=1.6 MULT=1
MM1017 A_801_47# N_A1_M1017_g N_A_84_21#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.12025 PD=0.93 PS=1.02 NRD=15.684 NRS=8.304 M=1 R=4.33333
+ SA=75004.1 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1009 A_991_47# N_A1_M1009_g N_A_84_21#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=14.76 NRS=8.304 M=1 R=4.33333
+ SA=75004.6 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1010_d N_A2_M1010_g A_991_47# VNB NSHORT L=0.15 W=0.65 AD=0.2015
+ AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=14.76 M=1 R=4.33333 SA=75005
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_84_21#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_A_84_21#_M1012_g N_X_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1012_d N_A_84_21#_M1018_g N_X_M1018_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.2
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1019 N_VPWR_M1019_d N_A_84_21#_M1019_g N_X_M1018_s VPB PHIGHVT L=0.18 W=1
+ AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1011 N_A_523_297#_M1011_d N_B1_M1011_g N_A_84_21#_M1011_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.7 A=0.18 P=2.36 MULT=1
MM1014 N_A_523_297#_M1014_d N_B1_M1014_g N_A_84_21#_M1011_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A2_M1004_g N_A_523_297#_M1014_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1001 N_A_523_297#_M1001_d N_A1_M1001_g N_VPWR_M1004_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1015 N_A_523_297#_M1001_d N_A1_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1015_s N_A2_M1013_g N_A_523_297#_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.405 PD=1.29 PS=2.81 NRD=0.9653 NRS=27.5603 M=1 R=5.55556
+ SA=90002.5 SB=90000.3 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.2078 P=15.93
pX21_noxref noxref_13 B1 B1 PROBETYPE=1
pX22_noxref noxref_14 A1 A1 PROBETYPE=1
pX23_noxref noxref_15 A2 A2 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__a21o_4.pxi.spice"
*
.ends
*
*
