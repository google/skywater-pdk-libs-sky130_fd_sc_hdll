* File: sky130_fd_sc_hdll__isobufsrc_2.spice
* Created: Thu Aug 27 19:09:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__isobufsrc_2.pex.spice"
.subckt sky130_fd_sc_hdll__isobufsrc_2  VNB VPB SLEEP A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* SLEEP	SLEEP
* VPB	VPB
* VNB	VNB
MM1004 N_X_M1004_d N_SLEEP_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.17875 PD=1.02 PS=1.85 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1004_d N_SLEEP_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1009_s N_A_271_21#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A_271_21#_M1008_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g N_A_271_21#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.1092 PD=1.46 PS=1.36 NRD=12.852 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_SLEEP_M1000_g N_A_27_297#_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1000_d N_SLEEP_M1007_g N_A_27_297#_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1002 N_A_27_297#_M1007_s N_A_271_21#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1003 N_A_27_297#_M1003_d N_A_271_21#_M1003_g N_X_M1002_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_271_21#_M1006_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.1134 AS=0.1134 PD=1.38 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
pX11_noxref noxref_10 A A PROBETYPE=1
*
.include "sky130_fd_sc_hdll__isobufsrc_2.pxi.spice"
*
.ends
*
*
