* File: sky130_fd_sc_hdll__and3b_2.pxi.spice
* Created: Thu Aug 27 18:58:25 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND3B_2%A_N N_A_N_c_67_n N_A_N_M1002_g N_A_N_M1000_g A_N
+ A_N PM_SKY130_FD_SC_HDLL__AND3B_2%A_N
x_PM_SKY130_FD_SC_HDLL__AND3B_2%A_117_311# N_A_117_311#_M1000_d
+ N_A_117_311#_M1002_d N_A_117_311#_c_91_n N_A_117_311#_M1007_g
+ N_A_117_311#_M1001_g N_A_117_311#_c_93_n N_A_117_311#_c_94_n
+ N_A_117_311#_c_95_n N_A_117_311#_c_96_n
+ PM_SKY130_FD_SC_HDLL__AND3B_2%A_117_311#
x_PM_SKY130_FD_SC_HDLL__AND3B_2%B N_B_c_132_n N_B_c_135_n N_B_M1003_g
+ N_B_M1009_g B B PM_SKY130_FD_SC_HDLL__AND3B_2%B
x_PM_SKY130_FD_SC_HDLL__AND3B_2%C N_C_M1010_g N_C_c_173_n N_C_M1004_g C C
+ N_C_c_175_n C PM_SKY130_FD_SC_HDLL__AND3B_2%C
x_PM_SKY130_FD_SC_HDLL__AND3B_2%A_225_311# N_A_225_311#_M1001_s
+ N_A_225_311#_M1007_s N_A_225_311#_M1003_d N_A_225_311#_c_223_n
+ N_A_225_311#_M1008_g N_A_225_311#_c_217_n N_A_225_311#_M1005_g
+ N_A_225_311#_c_224_n N_A_225_311#_M1011_g N_A_225_311#_c_218_n
+ N_A_225_311#_M1006_g N_A_225_311#_c_225_n N_A_225_311#_c_219_n
+ N_A_225_311#_c_226_n N_A_225_311#_c_227_n N_A_225_311#_c_220_n
+ N_A_225_311#_c_229_n N_A_225_311#_c_255_n N_A_225_311#_c_230_n
+ N_A_225_311#_c_221_n N_A_225_311#_c_274_p N_A_225_311#_c_232_n
+ N_A_225_311#_c_222_n PM_SKY130_FD_SC_HDLL__AND3B_2%A_225_311#
x_PM_SKY130_FD_SC_HDLL__AND3B_2%VPWR N_VPWR_M1002_s N_VPWR_M1007_d
+ N_VPWR_M1004_d N_VPWR_M1011_d N_VPWR_c_324_n N_VPWR_c_325_n N_VPWR_c_326_n
+ N_VPWR_c_327_n N_VPWR_c_328_n N_VPWR_c_329_n N_VPWR_c_340_n N_VPWR_c_330_n
+ N_VPWR_c_331_n VPWR N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_323_n
+ PM_SKY130_FD_SC_HDLL__AND3B_2%VPWR
x_PM_SKY130_FD_SC_HDLL__AND3B_2%X N_X_M1005_s N_X_M1008_s N_X_c_381_n X X X
+ N_X_c_399_n N_X_c_384_n X PM_SKY130_FD_SC_HDLL__AND3B_2%X
x_PM_SKY130_FD_SC_HDLL__AND3B_2%VGND N_VGND_M1000_s N_VGND_M1010_d
+ N_VGND_M1006_d N_VGND_c_414_n N_VGND_c_415_n N_VGND_c_416_n N_VGND_c_417_n
+ N_VGND_c_418_n N_VGND_c_419_n N_VGND_c_420_n VGND N_VGND_c_421_n
+ N_VGND_c_422_n PM_SKY130_FD_SC_HDLL__AND3B_2%VGND
cc_1 VNB N_A_N_c_67_n 0.0523483f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.48
cc_2 VNB N_A_N_M1000_g 0.035555f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_3 VNB A_N 0.0139484f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_4 VNB N_A_117_311#_c_91_n 0.0368975f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_117_311#_M1001_g 0.0340798f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_6 VNB N_A_117_311#_c_93_n 0.0144077f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_117_311#_c_94_n 0.00159635f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_117_311#_c_95_n 0.0151677f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_117_311#_c_96_n 0.00381195f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B_c_132_n 0.00835004f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.48
cc_11 VNB N_B_M1009_g 0.0346456f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_C_M1010_g 0.0268755f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.765
cc_13 VNB N_C_c_173_n 0.0223159f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_14 VNB C 5.99582e-19 $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_15 VNB N_C_c_175_n 0.00940708f $X=-0.19 $Y=-0.24 $X2=0.277 $Y2=0.85
cc_16 VNB N_A_225_311#_c_217_n 0.0190894f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_17 VNB N_A_225_311#_c_218_n 0.0207083f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_225_311#_c_219_n 0.00325624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_225_311#_c_220_n 0.0117236f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_225_311#_c_221_n 0.0052046f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_225_311#_c_222_n 0.0465687f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_323_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_X_c_381_n 8.34527e-19 $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_24 VNB X 0.0305864f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_25 VNB N_VGND_c_414_n 0.010079f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_415_n 0.0199242f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_27 VNB N_VGND_c_416_n 0.00598549f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_417_n 0.0109665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_418_n 0.0250577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_419_n 0.0598603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_420_n 0.00632082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_421_n 0.0220747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_422_n 0.244012f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VPB N_A_N_c_67_n 0.0509738f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.48
cc_35 VPB A_N 0.0026867f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_36 VPB N_A_117_311#_c_91_n 0.0398758f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_117_311#_c_94_n 0.0115999f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_B_c_132_n 0.0103921f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.48
cc_39 VPB N_B_c_135_n 0.0497316f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.765
cc_40 VPB N_B_M1003_g 0.0119497f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_41 VPB B 0.0111977f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_C_c_173_n 0.0272848f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.475
cc_43 VPB N_A_225_311#_c_223_n 0.0186516f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_225_311#_c_224_n 0.0192434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_225_311#_c_225_n 0.00361906f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_225_311#_c_226_n 0.00231847f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_225_311#_c_227_n 0.00337993f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_225_311#_c_220_n 0.00215932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_225_311#_c_229_n 0.00231379f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_225_311#_c_230_n 0.00647018f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_225_311#_c_221_n 0.00122146f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_225_311#_c_232_n 0.0014971f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_225_311#_c_222_n 0.025354f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_324_n 0.0109454f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_55 VPB N_VPWR_c_325_n 0.0616023f $X=-0.19 $Y=1.305 $X2=0.277 $Y2=0.85
cc_56 VPB N_VPWR_c_326_n 0.069176f $X=-0.19 $Y=1.305 $X2=0.277 $Y2=1.16
cc_57 VPB N_VPWR_c_327_n 0.00498362f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_328_n 0.0109406f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_329_n 0.03839f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_330_n 0.023503f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_331_n 0.00410958f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_332_n 0.0235637f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_333_n 0.00146642f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_323_n 0.0682922f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB X 0.0182412f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_66 VPB N_X_c_384_n 0.00203471f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 N_A_N_c_67_n N_A_117_311#_c_91_n 0.00524795f $X=0.495 $Y=1.48 $X2=0 $Y2=0
cc_68 N_A_N_M1000_g N_A_117_311#_c_93_n 0.00906231f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_69 A_N N_A_117_311#_c_93_n 0.0180715f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_70 N_A_N_c_67_n N_A_117_311#_c_94_n 0.0109697f $X=0.495 $Y=1.48 $X2=0 $Y2=0
cc_71 A_N N_A_117_311#_c_94_n 0.00502998f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_72 N_A_N_c_67_n N_A_117_311#_c_96_n 0.00345699f $X=0.495 $Y=1.48 $X2=0 $Y2=0
cc_73 A_N N_A_117_311#_c_96_n 0.0157538f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_74 N_A_N_c_67_n N_A_225_311#_c_225_n 0.00146303f $X=0.495 $Y=1.48 $X2=0 $Y2=0
cc_75 N_A_N_c_67_n N_VPWR_c_325_n 0.0108822f $X=0.495 $Y=1.48 $X2=0 $Y2=0
cc_76 A_N N_VPWR_c_325_n 0.0144894f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_77 N_A_N_c_67_n N_VPWR_c_326_n 0.00439574f $X=0.495 $Y=1.48 $X2=0 $Y2=0
cc_78 N_A_N_c_67_n N_VPWR_c_323_n 0.0052805f $X=0.495 $Y=1.48 $X2=0 $Y2=0
cc_79 N_A_N_c_67_n N_VGND_c_415_n 0.00226039f $X=0.495 $Y=1.48 $X2=0 $Y2=0
cc_80 N_A_N_M1000_g N_VGND_c_415_n 0.00639818f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_81 A_N N_VGND_c_415_n 0.0182064f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_82 N_A_N_M1000_g N_VGND_c_419_n 0.00555245f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_83 A_N N_VGND_c_419_n 8.67223e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_84 N_A_N_M1000_g N_VGND_c_422_n 0.0123489f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_85 A_N N_VGND_c_422_n 0.00238484f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_86 N_A_117_311#_c_91_n N_B_c_132_n 0.0115669f $X=1.485 $Y=1.48 $X2=-0.19
+ $Y2=-0.24
cc_87 N_A_117_311#_c_91_n N_B_c_135_n 8.20678e-19 $X=1.485 $Y=1.48 $X2=0 $Y2=0
cc_88 N_A_117_311#_c_91_n N_B_M1003_g 0.0125142f $X=1.485 $Y=1.48 $X2=0 $Y2=0
cc_89 N_A_117_311#_M1001_g N_B_M1009_g 0.0350576f $X=1.51 $Y=0.475 $X2=0 $Y2=0
cc_90 N_A_117_311#_M1001_g C 2.69787e-19 $X=1.51 $Y=0.475 $X2=0 $Y2=0
cc_91 N_A_117_311#_c_91_n N_A_225_311#_c_225_n 0.00426984f $X=1.485 $Y=1.48
+ $X2=0 $Y2=0
cc_92 N_A_117_311#_c_94_n N_A_225_311#_c_225_n 0.0224985f $X=0.73 $Y=1.74 $X2=0
+ $Y2=0
cc_93 N_A_117_311#_c_91_n N_A_225_311#_c_219_n 0.0056444f $X=1.485 $Y=1.48 $X2=0
+ $Y2=0
cc_94 N_A_117_311#_M1001_g N_A_225_311#_c_219_n 0.0141373f $X=1.51 $Y=0.475
+ $X2=0 $Y2=0
cc_95 N_A_117_311#_c_93_n N_A_225_311#_c_219_n 0.0205471f $X=0.75 $Y=0.47 $X2=0
+ $Y2=0
cc_96 N_A_117_311#_c_95_n N_A_225_311#_c_219_n 0.0117396f $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_97 N_A_117_311#_c_91_n N_A_225_311#_c_226_n 0.0191676f $X=1.485 $Y=1.48 $X2=0
+ $Y2=0
cc_98 N_A_117_311#_c_95_n N_A_225_311#_c_226_n 0.00876907f $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_99 N_A_117_311#_c_91_n N_A_225_311#_c_227_n 0.00506215f $X=1.485 $Y=1.48
+ $X2=0 $Y2=0
cc_100 N_A_117_311#_c_94_n N_A_225_311#_c_227_n 0.0134727f $X=0.73 $Y=1.74 $X2=0
+ $Y2=0
cc_101 N_A_117_311#_c_95_n N_A_225_311#_c_227_n 0.0182953f $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_102 N_A_117_311#_M1001_g N_A_225_311#_c_220_n 0.0171712f $X=1.51 $Y=0.475
+ $X2=0 $Y2=0
cc_103 N_A_117_311#_c_95_n N_A_225_311#_c_220_n 0.0174428f $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_104 N_A_117_311#_c_91_n N_VPWR_c_326_n 0.00448433f $X=1.485 $Y=1.48 $X2=0
+ $Y2=0
cc_105 N_A_117_311#_c_91_n N_VPWR_c_340_n 0.00389701f $X=1.485 $Y=1.48 $X2=0
+ $Y2=0
cc_106 N_A_117_311#_c_91_n N_VPWR_c_333_n 0.0107103f $X=1.485 $Y=1.48 $X2=0
+ $Y2=0
cc_107 N_A_117_311#_c_94_n N_VPWR_c_323_n 0.0109339f $X=0.73 $Y=1.74 $X2=0 $Y2=0
cc_108 N_A_117_311#_M1001_g N_VGND_c_419_n 0.00347765f $X=1.51 $Y=0.475 $X2=0
+ $Y2=0
cc_109 N_A_117_311#_c_93_n N_VGND_c_419_n 0.0140092f $X=0.75 $Y=0.47 $X2=0 $Y2=0
cc_110 N_A_117_311#_M1001_g N_VGND_c_422_n 0.0061559f $X=1.51 $Y=0.475 $X2=0
+ $Y2=0
cc_111 N_A_117_311#_c_93_n N_VGND_c_422_n 0.0102507f $X=0.75 $Y=0.47 $X2=0 $Y2=0
cc_112 N_B_M1009_g N_C_M1010_g 0.0386393f $X=1.98 $Y=0.475 $X2=0 $Y2=0
cc_113 N_B_c_132_n N_C_c_173_n 0.0447609f $X=1.955 $Y=1.48 $X2=0 $Y2=0
cc_114 N_B_M1003_g N_C_c_173_n 0.0115463f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_115 B N_C_c_173_n 0.00344582f $X=2.095 $Y=2.21 $X2=0 $Y2=0
cc_116 N_B_M1009_g C 0.0111354f $X=1.98 $Y=0.475 $X2=0 $Y2=0
cc_117 N_B_c_132_n N_C_c_175_n 0.00207038f $X=1.955 $Y=1.48 $X2=0 $Y2=0
cc_118 N_B_M1009_g N_C_c_175_n 0.0100724f $X=1.98 $Y=0.475 $X2=0 $Y2=0
cc_119 N_B_M1009_g N_A_225_311#_c_219_n 0.0021168f $X=1.98 $Y=0.475 $X2=0 $Y2=0
cc_120 N_B_c_132_n N_A_225_311#_c_220_n 0.00473301f $X=1.955 $Y=1.48 $X2=0 $Y2=0
cc_121 N_B_M1009_g N_A_225_311#_c_220_n 0.00440437f $X=1.98 $Y=0.475 $X2=0 $Y2=0
cc_122 N_B_c_132_n N_A_225_311#_c_229_n 0.00908193f $X=1.955 $Y=1.48 $X2=0 $Y2=0
cc_123 N_B_c_135_n N_A_225_311#_c_229_n 4.0052e-19 $X=1.955 $Y=2.105 $X2=0 $Y2=0
cc_124 N_B_M1003_g N_A_225_311#_c_229_n 0.00976113f $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_125 B N_A_225_311#_c_229_n 0.00670429f $X=2.095 $Y=2.21 $X2=0 $Y2=0
cc_126 N_B_M1003_g N_A_225_311#_c_255_n 0.00506553f $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_127 B N_A_225_311#_c_255_n 0.0113744f $X=2.095 $Y=2.21 $X2=0 $Y2=0
cc_128 B N_A_225_311#_c_230_n 0.00396479f $X=2.095 $Y=2.21 $X2=0 $Y2=0
cc_129 N_B_c_135_n N_VPWR_c_327_n 0.00251159f $X=1.955 $Y=2.105 $X2=0 $Y2=0
cc_130 N_B_M1003_g N_VPWR_c_327_n 0.0018517f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_131 B N_VPWR_c_327_n 0.0281462f $X=2.095 $Y=2.21 $X2=0 $Y2=0
cc_132 N_B_M1003_g N_VPWR_c_340_n 0.00357227f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_133 N_B_c_135_n N_VPWR_c_330_n 0.00690464f $X=1.955 $Y=2.105 $X2=0 $Y2=0
cc_134 B N_VPWR_c_330_n 0.0380394f $X=2.095 $Y=2.21 $X2=0 $Y2=0
cc_135 N_B_c_135_n N_VPWR_c_333_n 0.0103689f $X=1.955 $Y=2.105 $X2=0 $Y2=0
cc_136 N_B_M1003_g N_VPWR_c_333_n 0.0034845f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_137 B N_VPWR_c_333_n 0.0295124f $X=2.095 $Y=2.21 $X2=0 $Y2=0
cc_138 N_B_c_135_n N_VPWR_c_323_n 0.00959127f $X=1.955 $Y=2.105 $X2=0 $Y2=0
cc_139 B N_VPWR_c_323_n 0.020518f $X=2.095 $Y=2.21 $X2=0 $Y2=0
cc_140 N_B_M1009_g N_VGND_c_419_n 0.00459719f $X=1.98 $Y=0.475 $X2=0 $Y2=0
cc_141 N_B_M1009_g N_VGND_c_422_n 0.007918f $X=1.98 $Y=0.475 $X2=0 $Y2=0
cc_142 N_C_c_173_n N_A_225_311#_c_223_n 0.0152215f $X=2.48 $Y=1.41 $X2=0 $Y2=0
cc_143 N_C_M1010_g N_A_225_311#_c_217_n 0.0115903f $X=2.34 $Y=0.475 $X2=0 $Y2=0
cc_144 C N_A_225_311#_c_217_n 6.39831e-19 $X=2.04 $Y=0.425 $X2=0 $Y2=0
cc_145 N_C_c_175_n N_A_225_311#_c_217_n 0.00252666f $X=2.4 $Y=1.16 $X2=0 $Y2=0
cc_146 C N_A_225_311#_c_219_n 0.0221978f $X=2.04 $Y=0.425 $X2=0 $Y2=0
cc_147 C N_A_225_311#_c_220_n 0.0146415f $X=2.04 $Y=0.425 $X2=0 $Y2=0
cc_148 N_C_c_175_n N_A_225_311#_c_220_n 0.0379456f $X=2.4 $Y=1.16 $X2=0 $Y2=0
cc_149 N_C_c_175_n N_A_225_311#_c_229_n 0.0131276f $X=2.4 $Y=1.16 $X2=0 $Y2=0
cc_150 N_C_c_173_n N_A_225_311#_c_230_n 0.0161089f $X=2.48 $Y=1.41 $X2=0 $Y2=0
cc_151 N_C_c_175_n N_A_225_311#_c_230_n 0.0194667f $X=2.4 $Y=1.16 $X2=0 $Y2=0
cc_152 N_C_c_173_n N_A_225_311#_c_221_n 0.00452661f $X=2.48 $Y=1.41 $X2=0 $Y2=0
cc_153 N_C_c_175_n N_A_225_311#_c_221_n 0.0213462f $X=2.4 $Y=1.16 $X2=0 $Y2=0
cc_154 N_C_c_173_n N_A_225_311#_c_232_n 0.00250416f $X=2.48 $Y=1.41 $X2=0 $Y2=0
cc_155 N_C_c_175_n N_A_225_311#_c_232_n 0.0157434f $X=2.4 $Y=1.16 $X2=0 $Y2=0
cc_156 N_C_c_173_n N_A_225_311#_c_222_n 0.0228975f $X=2.48 $Y=1.41 $X2=0 $Y2=0
cc_157 N_C_c_175_n N_A_225_311#_c_222_n 9.04518e-19 $X=2.4 $Y=1.16 $X2=0 $Y2=0
cc_158 N_C_c_173_n N_VPWR_c_327_n 0.00459229f $X=2.48 $Y=1.41 $X2=0 $Y2=0
cc_159 N_C_c_173_n N_VPWR_c_340_n 2.9905e-19 $X=2.48 $Y=1.41 $X2=0 $Y2=0
cc_160 N_C_c_173_n N_VPWR_c_330_n 0.00180705f $X=2.48 $Y=1.41 $X2=0 $Y2=0
cc_161 N_C_c_173_n N_VPWR_c_323_n 0.00222661f $X=2.48 $Y=1.41 $X2=0 $Y2=0
cc_162 N_C_c_175_n N_X_c_381_n 0.0052023f $X=2.4 $Y=1.16 $X2=0 $Y2=0
cc_163 N_C_c_175_n X 0.00256979f $X=2.4 $Y=1.16 $X2=0 $Y2=0
cc_164 N_C_c_175_n N_VGND_M1010_d 0.0019417f $X=2.4 $Y=1.16 $X2=0 $Y2=0
cc_165 N_C_M1010_g N_VGND_c_416_n 0.00607497f $X=2.34 $Y=0.475 $X2=0 $Y2=0
cc_166 C N_VGND_c_416_n 0.0165713f $X=2.04 $Y=0.425 $X2=0 $Y2=0
cc_167 N_C_c_175_n N_VGND_c_416_n 7.23219e-19 $X=2.4 $Y=1.16 $X2=0 $Y2=0
cc_168 N_C_M1010_g N_VGND_c_419_n 0.00411264f $X=2.34 $Y=0.475 $X2=0 $Y2=0
cc_169 C N_VGND_c_419_n 0.0167205f $X=2.04 $Y=0.425 $X2=0 $Y2=0
cc_170 N_C_M1010_g N_VGND_c_422_n 0.00560252f $X=2.34 $Y=0.475 $X2=0 $Y2=0
cc_171 C N_VGND_c_422_n 0.0134002f $X=2.04 $Y=0.425 $X2=0 $Y2=0
cc_172 N_C_c_175_n N_VGND_c_422_n 0.00949801f $X=2.4 $Y=1.16 $X2=0 $Y2=0
cc_173 C A_411_53# 0.00103198f $X=2.04 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_174 N_A_225_311#_c_274_p N_VPWR_M1007_d 0.00180824f $X=1.73 $Y=1.51 $X2=0
+ $Y2=0
cc_175 N_A_225_311#_c_230_n N_VPWR_M1004_d 0.00364051f $X=2.79 $Y=1.51 $X2=0
+ $Y2=0
cc_176 N_A_225_311#_c_225_n N_VPWR_c_326_n 0.0204298f $X=1.25 $Y=1.76 $X2=0
+ $Y2=0
cc_177 N_A_225_311#_c_226_n N_VPWR_c_326_n 0.00498695f $X=1.645 $Y=1.51 $X2=0
+ $Y2=0
cc_178 N_A_225_311#_c_223_n N_VPWR_c_327_n 0.00450113f $X=3.015 $Y=1.41 $X2=0
+ $Y2=0
cc_179 N_A_225_311#_c_230_n N_VPWR_c_327_n 0.0157284f $X=2.79 $Y=1.51 $X2=0
+ $Y2=0
cc_180 N_A_225_311#_c_222_n N_VPWR_c_327_n 3.1527e-19 $X=3.485 $Y=1.202 $X2=0
+ $Y2=0
cc_181 N_A_225_311#_c_224_n N_VPWR_c_329_n 0.0101916f $X=3.485 $Y=1.41 $X2=0
+ $Y2=0
cc_182 N_A_225_311#_c_225_n N_VPWR_c_340_n 0.0144461f $X=1.25 $Y=1.76 $X2=0
+ $Y2=0
cc_183 N_A_225_311#_c_226_n N_VPWR_c_340_n 0.00566696f $X=1.645 $Y=1.51 $X2=0
+ $Y2=0
cc_184 N_A_225_311#_c_229_n N_VPWR_c_340_n 0.00133283f $X=2.16 $Y=1.51 $X2=0
+ $Y2=0
cc_185 N_A_225_311#_c_255_n N_VPWR_c_340_n 0.00647068f $X=2.245 $Y=1.725 $X2=0
+ $Y2=0
cc_186 N_A_225_311#_c_274_p N_VPWR_c_340_n 0.0133615f $X=1.73 $Y=1.51 $X2=0
+ $Y2=0
cc_187 N_A_225_311#_c_223_n N_VPWR_c_332_n 0.00702461f $X=3.015 $Y=1.41 $X2=0
+ $Y2=0
cc_188 N_A_225_311#_c_224_n N_VPWR_c_332_n 0.00429201f $X=3.485 $Y=1.41 $X2=0
+ $Y2=0
cc_189 N_A_225_311#_c_225_n N_VPWR_c_333_n 3.69269e-19 $X=1.25 $Y=1.76 $X2=0
+ $Y2=0
cc_190 N_A_225_311#_c_223_n N_VPWR_c_323_n 0.0137668f $X=3.015 $Y=1.41 $X2=0
+ $Y2=0
cc_191 N_A_225_311#_c_224_n N_VPWR_c_323_n 0.00713422f $X=3.485 $Y=1.41 $X2=0
+ $Y2=0
cc_192 N_A_225_311#_c_225_n N_VPWR_c_323_n 9.29713e-19 $X=1.25 $Y=1.76 $X2=0
+ $Y2=0
cc_193 N_A_225_311#_c_217_n N_X_c_381_n 0.0032307f $X=3.04 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_225_311#_c_218_n N_X_c_381_n 0.0122286f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_225_311#_c_222_n N_X_c_381_n 8.19151e-19 $X=3.485 $Y=1.202 $X2=0
+ $Y2=0
cc_196 N_A_225_311#_c_218_n X 0.0104443f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_225_311#_c_222_n X 0.00130953f $X=3.485 $Y=1.202 $X2=0 $Y2=0
cc_198 N_A_225_311#_c_223_n X 2.67766e-19 $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A_225_311#_c_217_n X 9.8064e-19 $X=3.04 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_225_311#_c_224_n X 0.00211583f $X=3.485 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A_225_311#_c_218_n X 0.0043268f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_225_311#_c_230_n X 0.00139394f $X=2.79 $Y=1.51 $X2=0 $Y2=0
cc_203 N_A_225_311#_c_221_n X 0.0275961f $X=2.935 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A_225_311#_c_222_n X 0.0324014f $X=3.485 $Y=1.202 $X2=0 $Y2=0
cc_205 N_A_225_311#_c_224_n N_X_c_399_n 0.0222707f $X=3.485 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A_225_311#_c_222_n N_X_c_399_n 0.00326491f $X=3.485 $Y=1.202 $X2=0
+ $Y2=0
cc_207 N_A_225_311#_c_223_n N_X_c_384_n 0.0059254f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A_225_311#_c_224_n N_X_c_384_n 0.0138798f $X=3.485 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A_225_311#_c_230_n N_X_c_384_n 0.0102321f $X=2.79 $Y=1.51 $X2=0 $Y2=0
cc_210 N_A_225_311#_c_222_n N_X_c_384_n 0.00106938f $X=3.485 $Y=1.202 $X2=0
+ $Y2=0
cc_211 N_A_225_311#_c_217_n N_VGND_c_416_n 0.00423828f $X=3.04 $Y=0.995 $X2=0
+ $Y2=0
cc_212 N_A_225_311#_c_221_n N_VGND_c_416_n 0.00572573f $X=2.935 $Y=1.16 $X2=0
+ $Y2=0
cc_213 N_A_225_311#_c_222_n N_VGND_c_416_n 8.28801e-19 $X=3.485 $Y=1.202 $X2=0
+ $Y2=0
cc_214 N_A_225_311#_c_218_n N_VGND_c_418_n 0.0138095f $X=3.51 $Y=0.995 $X2=0
+ $Y2=0
cc_215 N_A_225_311#_c_219_n N_VGND_c_419_n 0.0329523f $X=1.645 $Y=0.437 $X2=0
+ $Y2=0
cc_216 N_A_225_311#_c_217_n N_VGND_c_421_n 0.00585385f $X=3.04 $Y=0.995 $X2=0
+ $Y2=0
cc_217 N_A_225_311#_c_218_n N_VGND_c_421_n 0.00381957f $X=3.51 $Y=0.995 $X2=0
+ $Y2=0
cc_218 N_A_225_311#_c_217_n N_VGND_c_422_n 0.0115241f $X=3.04 $Y=0.995 $X2=0
+ $Y2=0
cc_219 N_A_225_311#_c_218_n N_VGND_c_422_n 0.00710512f $X=3.51 $Y=0.995 $X2=0
+ $Y2=0
cc_220 N_A_225_311#_c_219_n N_VGND_c_422_n 0.0253769f $X=1.645 $Y=0.437 $X2=0
+ $Y2=0
cc_221 N_A_225_311#_c_219_n A_317_53# 0.0046953f $X=1.645 $Y=0.437 $X2=-0.19
+ $Y2=-0.24
cc_222 N_A_225_311#_c_220_n A_317_53# 0.00244034f $X=1.73 $Y=1.425 $X2=-0.19
+ $Y2=-0.24
cc_223 N_VPWR_c_323_n N_X_M1008_s 0.00300692f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_224 N_VPWR_c_329_n X 0.0227078f $X=3.85 $Y=1.96 $X2=0 $Y2=0
cc_225 N_VPWR_c_332_n N_X_c_399_n 0.0284067f $X=3.76 $Y=2.72 $X2=0 $Y2=0
cc_226 N_VPWR_c_323_n N_X_c_399_n 0.0169336f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_227 X N_VGND_c_418_n 0.0347971f $X=3.36 $Y=0.425 $X2=0 $Y2=0
cc_228 X N_VGND_c_418_n 0.0227078f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_229 X N_VGND_c_421_n 0.0257037f $X=3.36 $Y=0.425 $X2=0 $Y2=0
cc_230 N_X_M1005_s N_VGND_c_422_n 0.00434007f $X=3.115 $Y=0.235 $X2=0 $Y2=0
cc_231 X N_VGND_c_422_n 0.0148742f $X=3.36 $Y=0.425 $X2=0 $Y2=0
