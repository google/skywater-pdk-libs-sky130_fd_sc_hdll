* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_521_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_409_297# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 Y a_119_47# a_409_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 VPWR A1_N a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 VGND a_119_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND A1_N a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_119_47# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y B2 a_521_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR B1 a_409_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 a_117_297# A2_N a_119_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
