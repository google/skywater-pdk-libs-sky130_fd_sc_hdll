* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_27_297# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VGND B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_109_47# B2 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_1259_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 Y a_831_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 VPWR A1_N a_1259_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_27_297# a_831_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 VPWR A1_N a_1259_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 Y B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Y a_831_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_831_21# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 Y B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 a_831_21# A2_N a_1259_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_1259_297# A2_N a_831_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 a_27_297# a_831_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 a_831_21# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_1259_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 VGND a_831_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_831_21# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_109_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_27_297# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 VGND a_831_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_831_21# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_109_47# B2 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VGND A1_N a_831_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X30 a_831_21# A2_N a_1259_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X31 VGND B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 Y a_831_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 Y a_831_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X34 a_1259_297# A2_N a_831_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X35 VGND A2_N a_831_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 VGND A1_N a_831_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 VPWR B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X38 a_109_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 VGND A2_N a_831_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
