* File: sky130_fd_sc_hdll__dlrtn_4.pxi.spice
* Created: Thu Aug 27 19:05:46 2020
* 
x_PM_SKY130_FD_SC_HDLL__DLRTN_4%GATE_N N_GATE_N_c_153_n N_GATE_N_c_154_n
+ N_GATE_N_M1003_g N_GATE_N_c_148_n N_GATE_N_M1018_g N_GATE_N_c_149_n GATE_N
+ N_GATE_N_c_151_n N_GATE_N_c_152_n PM_SKY130_FD_SC_HDLL__DLRTN_4%GATE_N
x_PM_SKY130_FD_SC_HDLL__DLRTN_4%A_27_363# N_A_27_363#_M1018_s
+ N_A_27_363#_M1003_s N_A_27_363#_M1005_g N_A_27_363#_c_198_n
+ N_A_27_363#_M1020_g N_A_27_363#_M1015_g N_A_27_363#_c_199_n
+ N_A_27_363#_M1019_g N_A_27_363#_c_200_n N_A_27_363#_c_335_p
+ N_A_27_363#_c_189_n N_A_27_363#_c_190_n N_A_27_363#_c_201_n
+ N_A_27_363#_c_191_n N_A_27_363#_c_264_p N_A_27_363#_c_192_n
+ N_A_27_363#_c_193_n N_A_27_363#_c_204_n N_A_27_363#_c_194_n
+ N_A_27_363#_c_195_n N_A_27_363#_c_196_n N_A_27_363#_c_205_n
+ N_A_27_363#_c_206_n N_A_27_363#_c_292_p N_A_27_363#_c_207_n
+ N_A_27_363#_c_197_n PM_SKY130_FD_SC_HDLL__DLRTN_4%A_27_363#
x_PM_SKY130_FD_SC_HDLL__DLRTN_4%D N_D_c_352_n N_D_c_353_n N_D_M1013_g
+ N_D_M1012_g N_D_c_349_n N_D_c_350_n D PM_SKY130_FD_SC_HDLL__DLRTN_4%D
x_PM_SKY130_FD_SC_HDLL__DLRTN_4%A_319_369# N_A_319_369#_M1012_s
+ N_A_319_369#_M1013_s N_A_319_369#_c_393_n N_A_319_369#_c_399_n
+ N_A_319_369#_M1008_g N_A_319_369#_M1023_g N_A_319_369#_c_400_n
+ N_A_319_369#_c_394_n N_A_319_369#_c_402_n N_A_319_369#_c_395_n
+ N_A_319_369#_c_396_n N_A_319_369#_c_397_n
+ PM_SKY130_FD_SC_HDLL__DLRTN_4%A_319_369#
x_PM_SKY130_FD_SC_HDLL__DLRTN_4%A_203_47# N_A_203_47#_M1005_d
+ N_A_203_47#_M1020_d N_A_203_47#_c_476_n N_A_203_47#_c_477_n
+ N_A_203_47#_M1021_g N_A_203_47#_c_471_n N_A_203_47#_M1009_g
+ N_A_203_47#_c_473_n N_A_203_47#_c_480_n N_A_203_47#_c_481_n
+ N_A_203_47#_c_482_n N_A_203_47#_c_483_n N_A_203_47#_c_515_n
+ N_A_203_47#_c_474_n N_A_203_47#_c_475_n
+ PM_SKY130_FD_SC_HDLL__DLRTN_4%A_203_47#
x_PM_SKY130_FD_SC_HDLL__DLRTN_4%A_750_21# N_A_750_21#_M1017_s
+ N_A_750_21#_M1024_d N_A_750_21#_M1001_g N_A_750_21#_c_586_n
+ N_A_750_21#_M1006_g N_A_750_21#_c_597_n N_A_750_21#_M1002_g
+ N_A_750_21#_c_587_n N_A_750_21#_M1000_g N_A_750_21#_c_588_n
+ N_A_750_21#_M1007_g N_A_750_21#_c_598_n N_A_750_21#_M1004_g
+ N_A_750_21#_c_599_n N_A_750_21#_M1011_g N_A_750_21#_c_589_n
+ N_A_750_21#_M1010_g N_A_750_21#_c_590_n N_A_750_21#_M1025_g
+ N_A_750_21#_c_600_n N_A_750_21#_M1022_g N_A_750_21#_c_601_n
+ N_A_750_21#_c_591_n N_A_750_21#_c_592_n N_A_750_21#_c_641_p
+ N_A_750_21#_c_603_n N_A_750_21#_c_593_n N_A_750_21#_c_685_p
+ N_A_750_21#_c_594_n N_A_750_21#_c_616_p N_A_750_21#_c_613_p
+ N_A_750_21#_c_595_n PM_SKY130_FD_SC_HDLL__DLRTN_4%A_750_21#
x_PM_SKY130_FD_SC_HDLL__DLRTN_4%A_604_47# N_A_604_47#_M1015_d
+ N_A_604_47#_M1021_d N_A_604_47#_c_742_n N_A_604_47#_c_750_n
+ N_A_604_47#_M1024_g N_A_604_47#_M1017_g N_A_604_47#_c_744_n
+ N_A_604_47#_c_755_n N_A_604_47#_c_759_n N_A_604_47#_c_745_n
+ N_A_604_47#_c_752_n N_A_604_47#_c_746_n N_A_604_47#_c_747_n
+ N_A_604_47#_c_748_n PM_SKY130_FD_SC_HDLL__DLRTN_4%A_604_47#
x_PM_SKY130_FD_SC_HDLL__DLRTN_4%RESET_B N_RESET_B_c_833_n N_RESET_B_M1014_g
+ N_RESET_B_c_834_n N_RESET_B_M1016_g RESET_B
+ PM_SKY130_FD_SC_HDLL__DLRTN_4%RESET_B
x_PM_SKY130_FD_SC_HDLL__DLRTN_4%VPWR N_VPWR_M1003_d N_VPWR_M1013_d
+ N_VPWR_M1006_d N_VPWR_M1016_d N_VPWR_M1004_s N_VPWR_M1022_s N_VPWR_c_868_n
+ N_VPWR_c_869_n N_VPWR_c_870_n N_VPWR_c_871_n N_VPWR_c_872_n N_VPWR_c_938_n
+ N_VPWR_c_873_n N_VPWR_c_874_n N_VPWR_c_875_n N_VPWR_c_876_n N_VPWR_c_877_n
+ N_VPWR_c_878_n VPWR N_VPWR_c_879_n N_VPWR_c_880_n N_VPWR_c_881_n
+ N_VPWR_c_867_n N_VPWR_c_883_n N_VPWR_c_884_n N_VPWR_c_885_n N_VPWR_c_886_n
+ PM_SKY130_FD_SC_HDLL__DLRTN_4%VPWR
x_PM_SKY130_FD_SC_HDLL__DLRTN_4%Q N_Q_M1000_d N_Q_M1010_d N_Q_M1002_d
+ N_Q_M1011_d N_Q_c_990_n N_Q_c_993_n N_Q_c_998_n N_Q_c_986_n N_Q_c_987_n
+ N_Q_c_1008_n N_Q_c_988_n N_Q_c_1019_n N_Q_c_1022_n N_Q_c_1024_n N_Q_c_1025_n
+ N_Q_c_1028_n Q PM_SKY130_FD_SC_HDLL__DLRTN_4%Q
x_PM_SKY130_FD_SC_HDLL__DLRTN_4%VGND N_VGND_M1018_d N_VGND_M1012_d
+ N_VGND_M1001_d N_VGND_M1014_d N_VGND_M1007_s N_VGND_M1025_s N_VGND_c_1058_n
+ N_VGND_c_1059_n N_VGND_c_1060_n N_VGND_c_1061_n N_VGND_c_1062_n
+ N_VGND_c_1063_n N_VGND_c_1064_n N_VGND_c_1065_n N_VGND_c_1066_n
+ N_VGND_c_1067_n N_VGND_c_1068_n N_VGND_c_1069_n VGND N_VGND_c_1070_n
+ N_VGND_c_1071_n N_VGND_c_1072_n N_VGND_c_1073_n N_VGND_c_1074_n
+ N_VGND_c_1075_n N_VGND_c_1076_n N_VGND_c_1077_n
+ PM_SKY130_FD_SC_HDLL__DLRTN_4%VGND
cc_1 VNB N_GATE_N_c_148_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_2 VNB N_GATE_N_c_149_n 0.0254388f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_3 VNB GATE_N 0.0196984f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_GATE_N_c_151_n 0.0178105f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.235
cc_5 VNB N_GATE_N_c_152_n 0.0157299f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.07
cc_6 VNB N_A_27_363#_M1005_g 0.0390164f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_7 VNB N_A_27_363#_M1015_g 0.0200544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_363#_c_189_n 0.00137507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_363#_c_190_n 0.00595335f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_363#_c_191_n 0.00235696f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_363#_c_192_n 5.38712e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_363#_c_193_n 0.00362448f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_363#_c_194_n 0.00401327f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_363#_c_195_n 0.0267668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_363#_c_196_n 0.00955011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_363#_c_197_n 0.0214946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_D_M1012_g 0.0323122f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_18 VNB N_D_c_349_n 0.0294753f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_19 VNB N_D_c_350_n 0.0116306f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=0.805
cc_20 VNB D 0.0124776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_319_369#_c_393_n 0.0137191f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_22 VNB N_A_319_369#_c_394_n 0.00197693f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_319_369#_c_395_n 0.0140494f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_319_369#_c_396_n 0.0231274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_319_369#_c_397_n 0.0172162f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_203_47#_c_471_n 0.0132521f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_203_47#_M1009_g 0.0385424f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_203_47#_c_473_n 0.0144111f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_203_47#_c_474_n 0.00964173f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_203_47#_c_475_n 0.00774225f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_750_21#_M1001_g 0.0440056f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_32 VNB N_A_750_21#_c_586_n 0.00267512f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=0.805
cc_33 VNB N_A_750_21#_c_587_n 0.0171447f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.665
cc_34 VNB N_A_750_21#_c_588_n 0.0167021f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_750_21#_c_589_n 0.0159577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_750_21#_c_590_n 0.0215085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_750_21#_c_591_n 0.00461115f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_750_21#_c_592_n 0.00473847f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_750_21#_c_593_n 0.00183578f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_750_21#_c_594_n 0.00314085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_750_21#_c_595_n 0.0852254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_604_47#_c_742_n 0.0116996f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_43 VNB N_A_604_47#_M1017_g 0.0273327f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_604_47#_c_744_n 0.00540275f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_604_47#_c_745_n 0.00311441f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_604_47#_c_746_n 0.0089303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_604_47#_c_747_n 0.00336267f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_604_47#_c_748_n 0.0289378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_RESET_B_c_833_n 0.0173376f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=0.88
cc_50 VNB N_RESET_B_c_834_n 0.0195736f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.59
cc_51 VNB RESET_B 0.0101451f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_52 VNB N_VPWR_c_867_n 0.326667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_Q_c_986_n 0.00165998f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.235
cc_54 VNB N_Q_c_987_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.07
cc_55 VNB N_Q_c_988_n 0.0107224f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1058_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.235
cc_57 VNB N_VGND_c_1059_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_58 VNB N_VGND_c_1060_n 0.00703343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1061_n 0.00557184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1062_n 0.00438892f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1063_n 0.00767379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1064_n 0.0321518f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1065_n 0.00634414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1066_n 0.0187037f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1067_n 0.00400911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1068_n 0.0173199f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1069_n 0.00403597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1070_n 0.0167943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1071_n 0.0299753f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1072_n 0.03956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1073_n 0.0134401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1074_n 0.411501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1075_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1076_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1077_n 0.00507956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VPB N_GATE_N_c_153_n 0.0130368f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.59
cc_77 VPB N_GATE_N_c_154_n 0.0457232f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.74
cc_78 VPB GATE_N 0.015162f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_79 VPB N_GATE_N_c_151_n 0.00836931f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.235
cc_80 VPB N_A_27_363#_c_198_n 0.0306782f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.805
cc_81 VPB N_A_27_363#_c_199_n 0.0478596f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_27_363#_c_200_n 0.0121265f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.235
cc_83 VPB N_A_27_363#_c_201_n 2.95372e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_27_363#_c_192_n 0.00385656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_27_363#_c_193_n 0.00298141f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_27_363#_c_204_n 0.0311606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_27_363#_c_205_n 0.0100987f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_27_363#_c_206_n 5.53836e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_27_363#_c_207_n 0.00859475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_27_363#_c_197_n 0.01105f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_D_c_352_n 0.0219473f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.07
cc_92 VPB N_D_c_353_n 0.0271128f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.4
cc_93 VPB N_D_c_349_n 0.0117743f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_94 VPB N_D_c_350_n 6.82386e-19 $X=-0.19 $Y=1.305 $X2=0.33 $Y2=0.805
cc_95 VPB N_A_319_369#_c_393_n 0.0175584f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_96 VPB N_A_319_369#_c_399_n 0.0233198f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_97 VPB N_A_319_369#_c_400_n 0.00828672f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.665
cc_98 VPB N_A_319_369#_c_394_n 0.00137236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_319_369#_c_402_n 0.00583579f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.235
cc_100 VPB N_A_203_47#_c_476_n 0.0136262f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_101 VPB N_A_203_47#_c_477_n 0.0232482f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_102 VPB N_A_203_47#_c_471_n 0.0170551f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_203_47#_c_473_n 0.00341069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_203_47#_c_480_n 0.0120963f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.07
cc_105 VPB N_A_203_47#_c_481_n 0.0116997f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_203_47#_c_482_n 0.00635095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_203_47#_c_483_n 0.00407738f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_203_47#_c_474_n 0.0231911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_203_47#_c_475_n 0.00381159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_750_21#_c_586_n 0.0878706f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=0.805
cc_111 VPB N_A_750_21#_c_597_n 0.0159868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_750_21#_c_598_n 0.0162464f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.235
cc_113 VPB N_A_750_21#_c_599_n 0.0155986f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_750_21#_c_600_n 0.0207627f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_750_21#_c_601_n 0.00310849f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_750_21#_c_592_n 0.00223949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_750_21#_c_603_n 0.00154179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_750_21#_c_595_n 0.0507666f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_604_47#_c_742_n 0.00770302f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_120 VPB N_A_604_47#_c_750_n 0.0198076f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_121 VPB N_A_604_47#_c_744_n 0.00700495f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_604_47#_c_752_n 0.0052925f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_604_47#_c_747_n 0.00167692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_604_47#_c_748_n 0.00663603f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_RESET_B_c_834_n 0.0245821f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.59
cc_126 VPB RESET_B 0.00222063f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_127 VPB N_VPWR_c_868_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.235
cc_128 VPB N_VPWR_c_869_n 0.0083008f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.4
cc_129 VPB N_VPWR_c_870_n 0.002048f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_871_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_872_n 0.00463848f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_873_n 0.0166118f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_874_n 0.00455763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_875_n 0.0178055f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_876_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_877_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_878_n 0.00487564f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_879_n 0.0157593f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_880_n 0.0302711f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_881_n 0.0120081f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_867_n 0.0596268f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_883_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_884_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_885_n 0.0472077f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_886_n 0.0201546f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_Q_c_988_n 0.00221657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 N_GATE_N_c_148_n N_A_27_363#_M1005_g 0.0188581f $X=0.52 $Y=0.73 $X2=0
+ $Y2=0
cc_148 N_GATE_N_c_152_n N_A_27_363#_M1005_g 0.00457196f $X=0.3 $Y=1.07 $X2=0
+ $Y2=0
cc_149 N_GATE_N_c_154_n N_A_27_363#_c_198_n 0.0262869f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_150 N_GATE_N_c_151_n N_A_27_363#_c_200_n 0.00540333f $X=0.3 $Y=1.235 $X2=0
+ $Y2=0
cc_151 N_GATE_N_c_148_n N_A_27_363#_c_189_n 0.00683119f $X=0.52 $Y=0.73 $X2=0
+ $Y2=0
cc_152 N_GATE_N_c_149_n N_A_27_363#_c_189_n 0.00930357f $X=0.52 $Y=0.805 $X2=0
+ $Y2=0
cc_153 GATE_N N_A_27_363#_c_189_n 0.00284891f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_154 N_GATE_N_c_149_n N_A_27_363#_c_190_n 0.0084621f $X=0.52 $Y=0.805 $X2=0
+ $Y2=0
cc_155 GATE_N N_A_27_363#_c_190_n 0.0133499f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_156 N_GATE_N_c_154_n N_A_27_363#_c_201_n 0.0162839f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_157 GATE_N N_A_27_363#_c_201_n 0.00301613f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_158 N_GATE_N_c_151_n N_A_27_363#_c_191_n 7.09938e-19 $X=0.3 $Y=1.235 $X2=0
+ $Y2=0
cc_159 N_GATE_N_c_153_n N_A_27_363#_c_192_n 7.09938e-19 $X=0.33 $Y=1.59 $X2=0
+ $Y2=0
cc_160 N_GATE_N_c_154_n N_A_27_363#_c_192_n 0.00497597f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_161 N_GATE_N_c_154_n N_A_27_363#_c_204_n 0.0055495f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_162 GATE_N N_A_27_363#_c_204_n 0.0279857f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_163 N_GATE_N_c_151_n N_A_27_363#_c_204_n 2.84016e-19 $X=0.3 $Y=1.235 $X2=0
+ $Y2=0
cc_164 N_GATE_N_c_149_n N_A_27_363#_c_194_n 0.00194152f $X=0.52 $Y=0.805 $X2=0
+ $Y2=0
cc_165 GATE_N N_A_27_363#_c_194_n 0.0495956f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_166 N_GATE_N_c_152_n N_A_27_363#_c_194_n 0.00309763f $X=0.3 $Y=1.07 $X2=0
+ $Y2=0
cc_167 N_GATE_N_c_154_n N_A_27_363#_c_206_n 0.00264502f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_168 GATE_N N_A_27_363#_c_197_n 3.13467e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_169 N_GATE_N_c_151_n N_A_27_363#_c_197_n 0.0175101f $X=0.3 $Y=1.235 $X2=0
+ $Y2=0
cc_170 N_GATE_N_c_154_n N_VPWR_c_868_n 0.00923212f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_171 N_GATE_N_c_154_n N_VPWR_c_879_n 0.0044329f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_172 N_GATE_N_c_154_n N_VPWR_c_867_n 0.00608656f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_173 N_GATE_N_c_148_n N_VGND_c_1058_n 0.00913236f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_174 N_GATE_N_c_148_n N_VGND_c_1070_n 0.00339367f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_175 N_GATE_N_c_149_n N_VGND_c_1070_n 5.87962e-19 $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_176 N_GATE_N_c_148_n N_VGND_c_1074_n 0.00502432f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_177 N_A_27_363#_c_205_n N_D_c_353_n 0.00409389f $X=3.22 $Y=1.87 $X2=0 $Y2=0
cc_178 N_A_27_363#_M1005_g N_D_c_349_n 0.0069171f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_179 N_A_27_363#_c_193_n N_A_319_369#_c_393_n 0.00350056f $X=3.21 $Y=1.575
+ $X2=0 $Y2=0
cc_180 N_A_27_363#_c_205_n N_A_319_369#_c_399_n 0.00677393f $X=3.22 $Y=1.87
+ $X2=0 $Y2=0
cc_181 N_A_27_363#_c_207_n N_A_319_369#_c_399_n 3.59161e-19 $X=3.365 $Y=1.87
+ $X2=0 $Y2=0
cc_182 N_A_27_363#_c_205_n N_A_319_369#_c_400_n 0.0211788f $X=3.22 $Y=1.87 $X2=0
+ $Y2=0
cc_183 N_A_27_363#_c_205_n N_A_319_369#_c_402_n 0.00465602f $X=3.22 $Y=1.87
+ $X2=0 $Y2=0
cc_184 N_A_27_363#_c_195_n N_A_319_369#_c_395_n 3.43721e-19 $X=2.945 $Y=0.9
+ $X2=0 $Y2=0
cc_185 N_A_27_363#_c_196_n N_A_319_369#_c_395_n 0.0212212f $X=3.21 $Y=0.915
+ $X2=0 $Y2=0
cc_186 N_A_27_363#_c_195_n N_A_319_369#_c_396_n 0.0144623f $X=2.945 $Y=0.9 $X2=0
+ $Y2=0
cc_187 N_A_27_363#_c_196_n N_A_319_369#_c_396_n 7.77092e-19 $X=3.21 $Y=0.915
+ $X2=0 $Y2=0
cc_188 N_A_27_363#_M1015_g N_A_319_369#_c_397_n 0.0220789f $X=2.945 $Y=0.415
+ $X2=0 $Y2=0
cc_189 N_A_27_363#_c_195_n N_A_319_369#_c_397_n 0.00124411f $X=2.945 $Y=0.9
+ $X2=0 $Y2=0
cc_190 N_A_27_363#_c_199_n N_A_203_47#_c_476_n 0.0053733f $X=3.42 $Y=1.99 $X2=0
+ $Y2=0
cc_191 N_A_27_363#_c_205_n N_A_203_47#_c_476_n 0.005923f $X=3.22 $Y=1.87 $X2=0
+ $Y2=0
cc_192 N_A_27_363#_c_199_n N_A_203_47#_c_477_n 0.0112656f $X=3.42 $Y=1.99 $X2=0
+ $Y2=0
cc_193 N_A_27_363#_c_205_n N_A_203_47#_c_477_n 0.00405726f $X=3.22 $Y=1.87 $X2=0
+ $Y2=0
cc_194 N_A_27_363#_c_199_n N_A_203_47#_c_471_n 0.018099f $X=3.42 $Y=1.99 $X2=0
+ $Y2=0
cc_195 N_A_27_363#_c_193_n N_A_203_47#_c_471_n 0.012296f $X=3.21 $Y=1.575 $X2=0
+ $Y2=0
cc_196 N_A_27_363#_c_196_n N_A_203_47#_c_471_n 8.98998e-19 $X=3.21 $Y=0.915
+ $X2=0 $Y2=0
cc_197 N_A_27_363#_c_205_n N_A_203_47#_c_471_n 0.00138393f $X=3.22 $Y=1.87 $X2=0
+ $Y2=0
cc_198 N_A_27_363#_c_207_n N_A_203_47#_c_471_n 0.00558349f $X=3.365 $Y=1.87
+ $X2=0 $Y2=0
cc_199 N_A_27_363#_M1015_g N_A_203_47#_M1009_g 0.00922459f $X=2.945 $Y=0.415
+ $X2=0 $Y2=0
cc_200 N_A_27_363#_c_193_n N_A_203_47#_M1009_g 0.00335377f $X=3.21 $Y=1.575
+ $X2=0 $Y2=0
cc_201 N_A_27_363#_c_195_n N_A_203_47#_M1009_g 0.0121069f $X=2.945 $Y=0.9 $X2=0
+ $Y2=0
cc_202 N_A_27_363#_c_196_n N_A_203_47#_M1009_g 0.00357812f $X=3.21 $Y=0.915
+ $X2=0 $Y2=0
cc_203 N_A_27_363#_M1005_g N_A_203_47#_c_473_n 0.00593261f $X=0.94 $Y=0.445
+ $X2=0 $Y2=0
cc_204 N_A_27_363#_c_189_n N_A_203_47#_c_473_n 0.00911803f $X=0.605 $Y=0.72
+ $X2=0 $Y2=0
cc_205 N_A_27_363#_c_191_n N_A_203_47#_c_473_n 0.025829f $X=0.75 $Y=1.215 $X2=0
+ $Y2=0
cc_206 N_A_27_363#_c_194_n N_A_203_47#_c_473_n 0.0136901f $X=0.75 $Y=1.07 $X2=0
+ $Y2=0
cc_207 N_A_27_363#_c_198_n N_A_203_47#_c_480_n 0.0057644f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_208 N_A_27_363#_c_200_n N_A_203_47#_c_480_n 0.00593261f $X=0.965 $Y=1.59
+ $X2=0 $Y2=0
cc_209 N_A_27_363#_c_264_p N_A_203_47#_c_480_n 0.00882838f $X=0.75 $Y=1.795
+ $X2=0 $Y2=0
cc_210 N_A_27_363#_c_205_n N_A_203_47#_c_480_n 0.0186521f $X=3.22 $Y=1.87 $X2=0
+ $Y2=0
cc_211 N_A_27_363#_c_206_n N_A_203_47#_c_480_n 0.00117183f $X=0.865 $Y=1.87
+ $X2=0 $Y2=0
cc_212 N_A_27_363#_c_205_n N_A_203_47#_c_481_n 0.105774f $X=3.22 $Y=1.87 $X2=0
+ $Y2=0
cc_213 N_A_27_363#_c_198_n N_A_203_47#_c_482_n 0.00170862f $X=0.965 $Y=1.74
+ $X2=0 $Y2=0
cc_214 N_A_27_363#_c_200_n N_A_203_47#_c_482_n 0.00515031f $X=0.965 $Y=1.59
+ $X2=0 $Y2=0
cc_215 N_A_27_363#_c_192_n N_A_203_47#_c_482_n 0.00721717f $X=0.81 $Y=1.235
+ $X2=0 $Y2=0
cc_216 N_A_27_363#_c_205_n N_A_203_47#_c_482_n 0.0251562f $X=3.22 $Y=1.87 $X2=0
+ $Y2=0
cc_217 N_A_27_363#_c_192_n N_A_203_47#_c_483_n 0.025829f $X=0.81 $Y=1.235 $X2=0
+ $Y2=0
cc_218 N_A_27_363#_c_197_n N_A_203_47#_c_483_n 0.00593261f $X=0.94 $Y=1.235
+ $X2=0 $Y2=0
cc_219 N_A_27_363#_c_193_n N_A_203_47#_c_515_n 0.00446852f $X=3.21 $Y=1.575
+ $X2=0 $Y2=0
cc_220 N_A_27_363#_c_196_n N_A_203_47#_c_515_n 9.8074e-19 $X=3.21 $Y=0.915 $X2=0
+ $Y2=0
cc_221 N_A_27_363#_c_205_n N_A_203_47#_c_515_n 0.0261499f $X=3.22 $Y=1.87 $X2=0
+ $Y2=0
cc_222 N_A_27_363#_c_207_n N_A_203_47#_c_515_n 0.00182791f $X=3.365 $Y=1.87
+ $X2=0 $Y2=0
cc_223 N_A_27_363#_c_199_n N_A_203_47#_c_474_n 0.016719f $X=3.42 $Y=1.99 $X2=0
+ $Y2=0
cc_224 N_A_27_363#_c_193_n N_A_203_47#_c_474_n 0.00411158f $X=3.21 $Y=1.575
+ $X2=0 $Y2=0
cc_225 N_A_27_363#_c_195_n N_A_203_47#_c_474_n 0.0211774f $X=2.945 $Y=0.9 $X2=0
+ $Y2=0
cc_226 N_A_27_363#_c_196_n N_A_203_47#_c_474_n 0.00551002f $X=3.21 $Y=0.915
+ $X2=0 $Y2=0
cc_227 N_A_27_363#_c_207_n N_A_203_47#_c_474_n 0.00863156f $X=3.365 $Y=1.87
+ $X2=0 $Y2=0
cc_228 N_A_27_363#_c_193_n N_A_203_47#_c_475_n 0.0212936f $X=3.21 $Y=1.575 $X2=0
+ $Y2=0
cc_229 N_A_27_363#_c_196_n N_A_203_47#_c_475_n 0.0132372f $X=3.21 $Y=0.915 $X2=0
+ $Y2=0
cc_230 N_A_27_363#_c_205_n N_A_203_47#_c_475_n 0.0156538f $X=3.22 $Y=1.87 $X2=0
+ $Y2=0
cc_231 N_A_27_363#_c_207_n N_A_203_47#_c_475_n 0.00800041f $X=3.365 $Y=1.87
+ $X2=0 $Y2=0
cc_232 N_A_27_363#_c_199_n N_A_750_21#_c_586_n 0.0476737f $X=3.42 $Y=1.99 $X2=0
+ $Y2=0
cc_233 N_A_27_363#_c_193_n N_A_750_21#_c_586_n 8.26114e-19 $X=3.21 $Y=1.575
+ $X2=0 $Y2=0
cc_234 N_A_27_363#_c_207_n N_A_750_21#_c_586_n 6.27988e-19 $X=3.365 $Y=1.87
+ $X2=0 $Y2=0
cc_235 N_A_27_363#_c_199_n N_A_604_47#_c_755_n 0.0127286f $X=3.42 $Y=1.99 $X2=0
+ $Y2=0
cc_236 N_A_27_363#_c_205_n N_A_604_47#_c_755_n 0.00338792f $X=3.22 $Y=1.87 $X2=0
+ $Y2=0
cc_237 N_A_27_363#_c_292_p N_A_604_47#_c_755_n 0.00120815f $X=3.365 $Y=1.87
+ $X2=0 $Y2=0
cc_238 N_A_27_363#_c_207_n N_A_604_47#_c_755_n 0.02443f $X=3.365 $Y=1.87 $X2=0
+ $Y2=0
cc_239 N_A_27_363#_c_195_n N_A_604_47#_c_759_n 0.00146696f $X=2.945 $Y=0.9 $X2=0
+ $Y2=0
cc_240 N_A_27_363#_c_196_n N_A_604_47#_c_759_n 0.0182656f $X=3.21 $Y=0.915 $X2=0
+ $Y2=0
cc_241 N_A_27_363#_M1015_g N_A_604_47#_c_745_n 7.58363e-19 $X=2.945 $Y=0.415
+ $X2=0 $Y2=0
cc_242 N_A_27_363#_c_195_n N_A_604_47#_c_745_n 2.13323e-19 $X=2.945 $Y=0.9 $X2=0
+ $Y2=0
cc_243 N_A_27_363#_c_196_n N_A_604_47#_c_745_n 0.0183748f $X=3.21 $Y=0.915 $X2=0
+ $Y2=0
cc_244 N_A_27_363#_c_199_n N_A_604_47#_c_752_n 0.0059256f $X=3.42 $Y=1.99 $X2=0
+ $Y2=0
cc_245 N_A_27_363#_c_193_n N_A_604_47#_c_752_n 0.0104035f $X=3.21 $Y=1.575 $X2=0
+ $Y2=0
cc_246 N_A_27_363#_c_292_p N_A_604_47#_c_752_n 0.0017055f $X=3.365 $Y=1.87 $X2=0
+ $Y2=0
cc_247 N_A_27_363#_c_207_n N_A_604_47#_c_752_n 0.0290753f $X=3.365 $Y=1.87 $X2=0
+ $Y2=0
cc_248 N_A_27_363#_c_199_n N_A_604_47#_c_746_n 0.00178452f $X=3.42 $Y=1.99 $X2=0
+ $Y2=0
cc_249 N_A_27_363#_c_193_n N_A_604_47#_c_746_n 0.012389f $X=3.21 $Y=1.575 $X2=0
+ $Y2=0
cc_250 N_A_27_363#_c_196_n N_A_604_47#_c_746_n 0.00778088f $X=3.21 $Y=0.915
+ $X2=0 $Y2=0
cc_251 N_A_27_363#_c_207_n N_A_604_47#_c_746_n 7.63243e-19 $X=3.365 $Y=1.87
+ $X2=0 $Y2=0
cc_252 N_A_27_363#_c_264_p N_VPWR_M1003_d 8.27335e-19 $X=0.75 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_253 N_A_27_363#_c_206_n N_VPWR_M1003_d 0.00205104f $X=0.865 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_254 N_A_27_363#_c_205_n N_VPWR_M1013_d 2.27104e-19 $X=3.22 $Y=1.87 $X2=0
+ $Y2=0
cc_255 N_A_27_363#_c_198_n N_VPWR_c_868_n 0.00922772f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_256 N_A_27_363#_c_201_n N_VPWR_c_868_n 0.0016327f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_257 N_A_27_363#_c_264_p N_VPWR_c_868_n 0.0156074f $X=0.75 $Y=1.795 $X2=0
+ $Y2=0
cc_258 N_A_27_363#_c_204_n N_VPWR_c_868_n 0.0127533f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_259 N_A_27_363#_c_206_n N_VPWR_c_868_n 0.00350507f $X=0.865 $Y=1.87 $X2=0
+ $Y2=0
cc_260 N_A_27_363#_c_205_n N_VPWR_c_869_n 0.0196711f $X=3.22 $Y=1.87 $X2=0 $Y2=0
cc_261 N_A_27_363#_c_201_n N_VPWR_c_879_n 0.00206959f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_262 N_A_27_363#_c_204_n N_VPWR_c_879_n 0.0220573f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_263 N_A_27_363#_c_198_n N_VPWR_c_880_n 0.00590576f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_264 N_A_27_363#_c_198_n N_VPWR_c_867_n 0.00667006f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_265 N_A_27_363#_c_199_n N_VPWR_c_867_n 0.00609959f $X=3.42 $Y=1.99 $X2=0
+ $Y2=0
cc_266 N_A_27_363#_c_201_n N_VPWR_c_867_n 0.00366495f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_267 N_A_27_363#_c_264_p N_VPWR_c_867_n 2.5417e-19 $X=0.75 $Y=1.795 $X2=0
+ $Y2=0
cc_268 N_A_27_363#_c_204_n N_VPWR_c_867_n 0.011857f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_269 N_A_27_363#_c_205_n N_VPWR_c_867_n 0.112853f $X=3.22 $Y=1.87 $X2=0 $Y2=0
cc_270 N_A_27_363#_c_206_n N_VPWR_c_867_n 0.0144885f $X=0.865 $Y=1.87 $X2=0
+ $Y2=0
cc_271 N_A_27_363#_c_292_p N_VPWR_c_867_n 0.0144105f $X=3.365 $Y=1.87 $X2=0
+ $Y2=0
cc_272 N_A_27_363#_c_199_n N_VPWR_c_885_n 0.00448856f $X=3.42 $Y=1.99 $X2=0
+ $Y2=0
cc_273 N_A_27_363#_c_205_n A_503_369# 0.00369043f $X=3.22 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_274 N_A_27_363#_c_189_n N_VGND_M1018_d 0.00151978f $X=0.605 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_275 N_A_27_363#_M1005_g N_VGND_c_1058_n 0.00953934f $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_276 N_A_27_363#_c_189_n N_VGND_c_1058_n 0.0123958f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_277 N_A_27_363#_c_191_n N_VGND_c_1058_n 0.00311311f $X=0.75 $Y=1.215 $X2=0
+ $Y2=0
cc_278 N_A_27_363#_c_197_n N_VGND_c_1058_n 6.85506e-19 $X=0.94 $Y=1.235 $X2=0
+ $Y2=0
cc_279 N_A_27_363#_M1015_g N_VGND_c_1059_n 0.00181512f $X=2.945 $Y=0.415 $X2=0
+ $Y2=0
cc_280 N_A_27_363#_c_335_p N_VGND_c_1070_n 0.00981821f $X=0.31 $Y=0.445 $X2=0
+ $Y2=0
cc_281 N_A_27_363#_c_189_n N_VGND_c_1070_n 0.00243651f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_282 N_A_27_363#_M1005_g N_VGND_c_1071_n 0.0046653f $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_283 N_A_27_363#_M1015_g N_VGND_c_1072_n 0.00439206f $X=2.945 $Y=0.415 $X2=0
+ $Y2=0
cc_284 N_A_27_363#_c_195_n N_VGND_c_1072_n 0.00155706f $X=2.945 $Y=0.9 $X2=0
+ $Y2=0
cc_285 N_A_27_363#_c_196_n N_VGND_c_1072_n 0.00358349f $X=3.21 $Y=0.915 $X2=0
+ $Y2=0
cc_286 N_A_27_363#_M1018_s N_VGND_c_1074_n 0.00366338f $X=0.185 $Y=0.235 $X2=0
+ $Y2=0
cc_287 N_A_27_363#_M1005_g N_VGND_c_1074_n 0.00934473f $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_288 N_A_27_363#_M1015_g N_VGND_c_1074_n 0.00664952f $X=2.945 $Y=0.415 $X2=0
+ $Y2=0
cc_289 N_A_27_363#_c_335_p N_VGND_c_1074_n 0.00634536f $X=0.31 $Y=0.445 $X2=0
+ $Y2=0
cc_290 N_A_27_363#_c_189_n N_VGND_c_1074_n 0.00525284f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_291 N_A_27_363#_c_195_n N_VGND_c_1074_n 0.00259944f $X=2.945 $Y=0.9 $X2=0
+ $Y2=0
cc_292 N_A_27_363#_c_196_n N_VGND_c_1074_n 0.00661169f $X=3.21 $Y=0.915 $X2=0
+ $Y2=0
cc_293 N_D_c_350_n N_A_319_369#_c_393_n 0.0154881f $X=1.955 $Y=1.16 $X2=0 $Y2=0
cc_294 N_D_c_352_n N_A_319_369#_c_399_n 0.0154881f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_295 N_D_c_353_n N_A_319_369#_c_399_n 0.009841f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_296 N_D_c_353_n N_A_319_369#_c_400_n 0.0134542f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_297 N_D_c_352_n N_A_319_369#_c_394_n 0.00766398f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_298 N_D_c_350_n N_A_319_369#_c_394_n 0.00732682f $X=1.955 $Y=1.16 $X2=0 $Y2=0
cc_299 D N_A_319_369#_c_394_n 0.0139513f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_300 N_D_c_352_n N_A_319_369#_c_402_n 0.0121171f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_301 N_D_c_349_n N_A_319_369#_c_402_n 0.00769683f $X=1.855 $Y=1.16 $X2=0 $Y2=0
cc_302 D N_A_319_369#_c_402_n 0.0118971f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_303 N_D_M1012_g N_A_319_369#_c_395_n 0.0222419f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_304 N_D_c_349_n N_A_319_369#_c_395_n 0.00632987f $X=1.855 $Y=1.16 $X2=0 $Y2=0
cc_305 N_D_c_350_n N_A_319_369#_c_395_n 0.00343492f $X=1.955 $Y=1.16 $X2=0 $Y2=0
cc_306 D N_A_319_369#_c_395_n 0.0196389f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_307 N_D_M1012_g N_A_319_369#_c_396_n 0.0213174f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_308 N_D_M1012_g N_A_319_369#_c_397_n 0.0138443f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_309 N_D_c_352_n N_A_203_47#_c_473_n 0.00250533f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_310 N_D_M1012_g N_A_203_47#_c_473_n 0.00569292f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_311 N_D_c_349_n N_A_203_47#_c_473_n 0.0015971f $X=1.855 $Y=1.16 $X2=0 $Y2=0
cc_312 D N_A_203_47#_c_473_n 0.0243991f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_313 N_D_c_352_n N_A_203_47#_c_480_n 4.03124e-19 $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_314 N_D_c_353_n N_A_203_47#_c_480_n 0.00118287f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_315 N_D_c_352_n N_A_203_47#_c_481_n 0.0041274f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_316 N_D_c_349_n N_A_203_47#_c_481_n 0.00959604f $X=1.855 $Y=1.16 $X2=0 $Y2=0
cc_317 D N_A_203_47#_c_481_n 0.0109338f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_318 N_D_c_352_n N_A_203_47#_c_482_n 6.03063e-19 $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_319 N_D_c_352_n N_A_203_47#_c_483_n 0.00118508f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_320 N_D_c_352_n N_A_203_47#_c_475_n 3.09224e-19 $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_321 N_D_c_350_n N_A_203_47#_c_475_n 2.52874e-19 $X=1.955 $Y=1.16 $X2=0 $Y2=0
cc_322 N_D_c_353_n N_VPWR_c_869_n 0.00329547f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_323 N_D_c_353_n N_VPWR_c_880_n 0.00673617f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_324 N_D_c_353_n N_VPWR_c_867_n 0.00835409f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_325 N_D_M1012_g N_VGND_c_1059_n 0.0111499f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_326 N_D_M1012_g N_VGND_c_1071_n 0.00336882f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_327 N_D_M1012_g N_VGND_c_1074_n 0.00532348f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_328 N_A_319_369#_c_393_n N_A_203_47#_c_476_n 0.00540817f $X=2.425 $Y=1.67
+ $X2=0 $Y2=0
cc_329 N_A_319_369#_c_399_n N_A_203_47#_c_476_n 0.00877513f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_330 N_A_319_369#_c_399_n N_A_203_47#_c_477_n 0.0230867f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_331 N_A_319_369#_c_395_n N_A_203_47#_c_473_n 0.0173676f $X=2.03 $Y=0.72 $X2=0
+ $Y2=0
cc_332 N_A_319_369#_c_400_n N_A_203_47#_c_480_n 0.0530041f $X=1.72 $Y=1.99 $X2=0
+ $Y2=0
cc_333 N_A_319_369#_c_393_n N_A_203_47#_c_481_n 0.00352657f $X=2.425 $Y=1.67
+ $X2=0 $Y2=0
cc_334 N_A_319_369#_c_400_n N_A_203_47#_c_481_n 4.87587e-19 $X=1.72 $Y=1.99
+ $X2=0 $Y2=0
cc_335 N_A_319_369#_c_394_n N_A_203_47#_c_481_n 0.0110072f $X=2.03 $Y=1.495
+ $X2=0 $Y2=0
cc_336 N_A_319_369#_c_402_n N_A_203_47#_c_481_n 0.01758f $X=2.03 $Y=1.58 $X2=0
+ $Y2=0
cc_337 N_A_319_369#_c_395_n N_A_203_47#_c_481_n 0.0126321f $X=2.03 $Y=0.72 $X2=0
+ $Y2=0
cc_338 N_A_319_369#_c_402_n N_A_203_47#_c_482_n 3.60176e-19 $X=2.03 $Y=1.58
+ $X2=0 $Y2=0
cc_339 N_A_319_369#_c_394_n N_A_203_47#_c_483_n 9.03084e-19 $X=2.03 $Y=1.495
+ $X2=0 $Y2=0
cc_340 N_A_319_369#_c_402_n N_A_203_47#_c_483_n 0.0100074f $X=2.03 $Y=1.58 $X2=0
+ $Y2=0
cc_341 N_A_319_369#_c_394_n N_A_203_47#_c_515_n 2.15582e-19 $X=2.03 $Y=1.495
+ $X2=0 $Y2=0
cc_342 N_A_319_369#_c_402_n N_A_203_47#_c_515_n 2.48695e-19 $X=2.03 $Y=1.58
+ $X2=0 $Y2=0
cc_343 N_A_319_369#_c_393_n N_A_203_47#_c_474_n 0.0253968f $X=2.425 $Y=1.67
+ $X2=0 $Y2=0
cc_344 N_A_319_369#_c_393_n N_A_203_47#_c_475_n 0.0118476f $X=2.425 $Y=1.67
+ $X2=0 $Y2=0
cc_345 N_A_319_369#_c_399_n N_A_203_47#_c_475_n 0.0018263f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_346 N_A_319_369#_c_400_n N_A_203_47#_c_475_n 5.53168e-19 $X=1.72 $Y=1.99
+ $X2=0 $Y2=0
cc_347 N_A_319_369#_c_394_n N_A_203_47#_c_475_n 0.0101463f $X=2.03 $Y=1.495
+ $X2=0 $Y2=0
cc_348 N_A_319_369#_c_402_n N_A_203_47#_c_475_n 0.0065905f $X=2.03 $Y=1.58 $X2=0
+ $Y2=0
cc_349 N_A_319_369#_c_395_n N_A_203_47#_c_475_n 0.00654622f $X=2.03 $Y=0.72
+ $X2=0 $Y2=0
cc_350 N_A_319_369#_c_399_n N_A_604_47#_c_755_n 9.84369e-19 $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_351 N_A_319_369#_c_399_n N_VPWR_c_869_n 0.00422565f $X=2.425 $Y=1.77 $X2=0
+ $Y2=0
cc_352 N_A_319_369#_c_400_n N_VPWR_c_869_n 0.025165f $X=1.72 $Y=1.99 $X2=0 $Y2=0
cc_353 N_A_319_369#_c_402_n N_VPWR_c_869_n 0.00394172f $X=2.03 $Y=1.58 $X2=0
+ $Y2=0
cc_354 N_A_319_369#_c_400_n N_VPWR_c_880_n 0.0210596f $X=1.72 $Y=1.99 $X2=0
+ $Y2=0
cc_355 N_A_319_369#_M1013_s N_VPWR_c_867_n 0.00179197f $X=1.595 $Y=1.845 $X2=0
+ $Y2=0
cc_356 N_A_319_369#_c_399_n N_VPWR_c_867_n 0.0074238f $X=2.425 $Y=1.77 $X2=0
+ $Y2=0
cc_357 N_A_319_369#_c_400_n N_VPWR_c_867_n 0.00594162f $X=1.72 $Y=1.99 $X2=0
+ $Y2=0
cc_358 N_A_319_369#_c_399_n N_VPWR_c_885_n 0.00702461f $X=2.425 $Y=1.77 $X2=0
+ $Y2=0
cc_359 N_A_319_369#_c_395_n N_VGND_M1012_d 5.4803e-19 $X=2.03 $Y=0.72 $X2=0
+ $Y2=0
cc_360 N_A_319_369#_c_395_n N_VGND_c_1059_n 0.0120795f $X=2.03 $Y=0.72 $X2=0
+ $Y2=0
cc_361 N_A_319_369#_c_396_n N_VGND_c_1059_n 3.80743e-19 $X=2.4 $Y=0.93 $X2=0
+ $Y2=0
cc_362 N_A_319_369#_c_397_n N_VGND_c_1059_n 0.00798806f $X=2.4 $Y=0.765 $X2=0
+ $Y2=0
cc_363 N_A_319_369#_c_395_n N_VGND_c_1071_n 0.0109521f $X=2.03 $Y=0.72 $X2=0
+ $Y2=0
cc_364 N_A_319_369#_c_396_n N_VGND_c_1072_n 2.5317e-19 $X=2.4 $Y=0.93 $X2=0
+ $Y2=0
cc_365 N_A_319_369#_c_397_n N_VGND_c_1072_n 0.00564095f $X=2.4 $Y=0.765 $X2=0
+ $Y2=0
cc_366 N_A_319_369#_M1012_s N_VGND_c_1074_n 0.00285324f $X=1.645 $Y=0.235 $X2=0
+ $Y2=0
cc_367 N_A_319_369#_c_395_n N_VGND_c_1074_n 0.0189897f $X=2.03 $Y=0.72 $X2=0
+ $Y2=0
cc_368 N_A_319_369#_c_397_n N_VGND_c_1074_n 0.00527362f $X=2.4 $Y=0.765 $X2=0
+ $Y2=0
cc_369 N_A_203_47#_M1009_g N_A_750_21#_M1001_g 0.0394664f $X=3.465 $Y=0.445
+ $X2=0 $Y2=0
cc_370 N_A_203_47#_c_471_n N_A_750_21#_c_586_n 0.0394664f $X=3.39 $Y=1.32 $X2=0
+ $Y2=0
cc_371 N_A_203_47#_c_474_n N_A_750_21#_c_586_n 2.81272e-19 $X=2.892 $Y=1.32
+ $X2=0 $Y2=0
cc_372 N_A_203_47#_c_477_n N_A_604_47#_c_755_n 0.00515668f $X=2.95 $Y=1.99 $X2=0
+ $Y2=0
cc_373 N_A_203_47#_c_471_n N_A_604_47#_c_759_n 0.00138963f $X=3.39 $Y=1.32 $X2=0
+ $Y2=0
cc_374 N_A_203_47#_M1009_g N_A_604_47#_c_759_n 0.0113891f $X=3.465 $Y=0.445
+ $X2=0 $Y2=0
cc_375 N_A_203_47#_M1009_g N_A_604_47#_c_745_n 0.00872448f $X=3.465 $Y=0.445
+ $X2=0 $Y2=0
cc_376 N_A_203_47#_c_471_n N_A_604_47#_c_752_n 6.06088e-19 $X=3.39 $Y=1.32 $X2=0
+ $Y2=0
cc_377 N_A_203_47#_c_474_n N_A_604_47#_c_752_n 4.18131e-19 $X=2.892 $Y=1.32
+ $X2=0 $Y2=0
cc_378 N_A_203_47#_M1009_g N_A_604_47#_c_746_n 0.0061787f $X=3.465 $Y=0.445
+ $X2=0 $Y2=0
cc_379 N_A_203_47#_c_480_n N_VPWR_c_868_n 0.0127456f $X=1.2 $Y=1.96 $X2=0 $Y2=0
cc_380 N_A_203_47#_c_481_n N_VPWR_c_869_n 0.00140184f $X=2.665 $Y=1.53 $X2=0
+ $Y2=0
cc_381 N_A_203_47#_c_480_n N_VPWR_c_880_n 0.0192143f $X=1.2 $Y=1.96 $X2=0 $Y2=0
cc_382 N_A_203_47#_c_477_n N_VPWR_c_867_n 0.00771671f $X=2.95 $Y=1.99 $X2=0
+ $Y2=0
cc_383 N_A_203_47#_c_480_n N_VPWR_c_867_n 0.00491647f $X=1.2 $Y=1.96 $X2=0 $Y2=0
cc_384 N_A_203_47#_c_477_n N_VPWR_c_885_n 0.00694986f $X=2.95 $Y=1.99 $X2=0
+ $Y2=0
cc_385 N_A_203_47#_M1009_g N_VGND_c_1060_n 0.0016369f $X=3.465 $Y=0.445 $X2=0
+ $Y2=0
cc_386 N_A_203_47#_c_473_n N_VGND_c_1071_n 0.00999887f $X=1.15 $Y=0.445 $X2=0
+ $Y2=0
cc_387 N_A_203_47#_M1009_g N_VGND_c_1072_n 0.00362991f $X=3.465 $Y=0.445 $X2=0
+ $Y2=0
cc_388 N_A_203_47#_M1005_d N_VGND_c_1074_n 0.00530224f $X=1.015 $Y=0.235 $X2=0
+ $Y2=0
cc_389 N_A_203_47#_M1009_g N_VGND_c_1074_n 0.00539993f $X=3.465 $Y=0.445 $X2=0
+ $Y2=0
cc_390 N_A_203_47#_c_473_n N_VGND_c_1074_n 0.00639171f $X=1.15 $Y=0.445 $X2=0
+ $Y2=0
cc_391 N_A_750_21#_c_592_n N_A_604_47#_c_742_n 0.010664f $X=4.635 $Y=1.535 $X2=0
+ $Y2=0
cc_392 N_A_750_21#_c_594_n N_A_604_47#_c_742_n 0.00309332f $X=4.62 $Y=0.825
+ $X2=0 $Y2=0
cc_393 N_A_750_21#_c_613_p N_A_604_47#_c_742_n 6.70661e-19 $X=5.175 $Y=1.7 $X2=0
+ $Y2=0
cc_394 N_A_750_21#_c_586_n N_A_604_47#_c_750_n 0.01028f $X=3.9 $Y=1.99 $X2=0
+ $Y2=0
cc_395 N_A_750_21#_c_592_n N_A_604_47#_c_750_n 0.00421619f $X=4.635 $Y=1.535
+ $X2=0 $Y2=0
cc_396 N_A_750_21#_c_616_p N_A_604_47#_c_750_n 0.0164274f $X=5.025 $Y=1.7 $X2=0
+ $Y2=0
cc_397 N_A_750_21#_c_613_p N_A_604_47#_c_750_n 0.0235927f $X=5.175 $Y=1.7 $X2=0
+ $Y2=0
cc_398 N_A_750_21#_c_591_n N_A_604_47#_M1017_g 0.00737376f $X=4.62 $Y=0.38 $X2=0
+ $Y2=0
cc_399 N_A_750_21#_c_592_n N_A_604_47#_M1017_g 0.00577472f $X=4.635 $Y=1.535
+ $X2=0 $Y2=0
cc_400 N_A_750_21#_c_594_n N_A_604_47#_M1017_g 0.00433812f $X=4.62 $Y=0.825
+ $X2=0 $Y2=0
cc_401 N_A_750_21#_c_592_n N_A_604_47#_c_744_n 0.00545235f $X=4.635 $Y=1.535
+ $X2=0 $Y2=0
cc_402 N_A_750_21#_c_586_n N_A_604_47#_c_755_n 0.00595901f $X=3.9 $Y=1.99 $X2=0
+ $Y2=0
cc_403 N_A_750_21#_M1001_g N_A_604_47#_c_759_n 0.00206262f $X=3.825 $Y=0.445
+ $X2=0 $Y2=0
cc_404 N_A_750_21#_M1001_g N_A_604_47#_c_745_n 0.00870159f $X=3.825 $Y=0.445
+ $X2=0 $Y2=0
cc_405 N_A_750_21#_c_586_n N_A_604_47#_c_752_n 0.0355361f $X=3.9 $Y=1.99 $X2=0
+ $Y2=0
cc_406 N_A_750_21#_c_601_n N_A_604_47#_c_752_n 0.0246758f $X=4.55 $Y=1.7 $X2=0
+ $Y2=0
cc_407 N_A_750_21#_M1001_g N_A_604_47#_c_746_n 0.00970956f $X=3.825 $Y=0.445
+ $X2=0 $Y2=0
cc_408 N_A_750_21#_c_586_n N_A_604_47#_c_746_n 6.43776e-19 $X=3.9 $Y=1.99 $X2=0
+ $Y2=0
cc_409 N_A_750_21#_M1001_g N_A_604_47#_c_747_n 0.00591896f $X=3.825 $Y=0.445
+ $X2=0 $Y2=0
cc_410 N_A_750_21#_c_586_n N_A_604_47#_c_747_n 0.0129533f $X=3.9 $Y=1.99 $X2=0
+ $Y2=0
cc_411 N_A_750_21#_c_601_n N_A_604_47#_c_747_n 0.0239061f $X=4.55 $Y=1.7 $X2=0
+ $Y2=0
cc_412 N_A_750_21#_c_592_n N_A_604_47#_c_747_n 0.0256838f $X=4.635 $Y=1.535
+ $X2=0 $Y2=0
cc_413 N_A_750_21#_M1001_g N_A_604_47#_c_748_n 0.0138805f $X=3.825 $Y=0.445
+ $X2=0 $Y2=0
cc_414 N_A_750_21#_c_586_n N_A_604_47#_c_748_n 0.00935438f $X=3.9 $Y=1.99 $X2=0
+ $Y2=0
cc_415 N_A_750_21#_c_601_n N_A_604_47#_c_748_n 0.00919786f $X=4.55 $Y=1.7 $X2=0
+ $Y2=0
cc_416 N_A_750_21#_c_592_n N_A_604_47#_c_748_n 0.00131564f $X=4.635 $Y=1.535
+ $X2=0 $Y2=0
cc_417 N_A_750_21#_c_587_n N_RESET_B_c_833_n 0.0161933f $X=5.77 $Y=0.995
+ $X2=-0.19 $Y2=-0.24
cc_418 N_A_750_21#_c_591_n N_RESET_B_c_833_n 0.00167505f $X=4.62 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_419 N_A_750_21#_c_597_n N_RESET_B_c_834_n 0.0210961f $X=5.745 $Y=1.41 $X2=0
+ $Y2=0
cc_420 N_A_750_21#_c_592_n N_RESET_B_c_834_n 0.00104943f $X=4.635 $Y=1.535 $X2=0
+ $Y2=0
cc_421 N_A_750_21#_c_641_p N_RESET_B_c_834_n 0.0152362f $X=5.555 $Y=1.62 $X2=0
+ $Y2=0
cc_422 N_A_750_21#_c_603_n N_RESET_B_c_834_n 0.00426133f $X=5.64 $Y=1.535 $X2=0
+ $Y2=0
cc_423 N_A_750_21#_c_593_n N_RESET_B_c_834_n 9.31102e-19 $X=5.725 $Y=1.2 $X2=0
+ $Y2=0
cc_424 N_A_750_21#_c_613_p N_RESET_B_c_834_n 0.00125633f $X=5.175 $Y=1.7 $X2=0
+ $Y2=0
cc_425 N_A_750_21#_c_595_n N_RESET_B_c_834_n 0.0253249f $X=7.13 $Y=1.202 $X2=0
+ $Y2=0
cc_426 N_A_750_21#_c_592_n RESET_B 0.0249612f $X=4.635 $Y=1.535 $X2=0 $Y2=0
cc_427 N_A_750_21#_c_593_n RESET_B 0.0217023f $X=5.725 $Y=1.2 $X2=0 $Y2=0
cc_428 N_A_750_21#_c_613_p RESET_B 0.0279176f $X=5.175 $Y=1.7 $X2=0 $Y2=0
cc_429 N_A_750_21#_c_595_n RESET_B 8.88102e-19 $X=7.13 $Y=1.202 $X2=0 $Y2=0
cc_430 N_A_750_21#_c_601_n N_VPWR_M1006_d 0.00480268f $X=4.55 $Y=1.7 $X2=0 $Y2=0
cc_431 N_A_750_21#_c_592_n N_VPWR_M1006_d 0.00115467f $X=4.635 $Y=1.535 $X2=0
+ $Y2=0
cc_432 N_A_750_21#_c_613_p N_VPWR_M1006_d 0.001673f $X=5.175 $Y=1.7 $X2=0 $Y2=0
cc_433 N_A_750_21#_c_641_p N_VPWR_M1016_d 0.00690342f $X=5.555 $Y=1.62 $X2=0
+ $Y2=0
cc_434 N_A_750_21#_c_603_n N_VPWR_M1016_d 5.76203e-19 $X=5.64 $Y=1.535 $X2=0
+ $Y2=0
cc_435 N_A_750_21#_c_597_n N_VPWR_c_870_n 0.0017544f $X=5.745 $Y=1.41 $X2=0
+ $Y2=0
cc_436 N_A_750_21#_c_598_n N_VPWR_c_871_n 0.00173895f $X=6.215 $Y=1.41 $X2=0
+ $Y2=0
cc_437 N_A_750_21#_c_599_n N_VPWR_c_871_n 0.00173895f $X=6.685 $Y=1.41 $X2=0
+ $Y2=0
cc_438 N_A_750_21#_c_595_n N_VPWR_c_871_n 6.152e-19 $X=7.13 $Y=1.202 $X2=0 $Y2=0
cc_439 N_A_750_21#_c_600_n N_VPWR_c_872_n 0.00354036f $X=7.155 $Y=1.41 $X2=0
+ $Y2=0
cc_440 N_A_750_21#_c_597_n N_VPWR_c_938_n 0.00351799f $X=5.745 $Y=1.41 $X2=0
+ $Y2=0
cc_441 N_A_750_21#_c_641_p N_VPWR_c_938_n 0.0174587f $X=5.555 $Y=1.62 $X2=0
+ $Y2=0
cc_442 N_A_750_21#_c_616_p N_VPWR_c_873_n 0.0143928f $X=5.025 $Y=1.7 $X2=0 $Y2=0
cc_443 N_A_750_21#_c_597_n N_VPWR_c_875_n 0.00652041f $X=5.745 $Y=1.41 $X2=0
+ $Y2=0
cc_444 N_A_750_21#_c_598_n N_VPWR_c_875_n 0.00673617f $X=6.215 $Y=1.41 $X2=0
+ $Y2=0
cc_445 N_A_750_21#_c_599_n N_VPWR_c_877_n 0.00673617f $X=6.685 $Y=1.41 $X2=0
+ $Y2=0
cc_446 N_A_750_21#_c_600_n N_VPWR_c_877_n 0.00673617f $X=7.155 $Y=1.41 $X2=0
+ $Y2=0
cc_447 N_A_750_21#_M1024_d N_VPWR_c_867_n 0.00268338f $X=4.895 $Y=1.485 $X2=0
+ $Y2=0
cc_448 N_A_750_21#_c_586_n N_VPWR_c_867_n 0.01305f $X=3.9 $Y=1.99 $X2=0 $Y2=0
cc_449 N_A_750_21#_c_597_n N_VPWR_c_867_n 0.0111327f $X=5.745 $Y=1.41 $X2=0
+ $Y2=0
cc_450 N_A_750_21#_c_598_n N_VPWR_c_867_n 0.0117184f $X=6.215 $Y=1.41 $X2=0
+ $Y2=0
cc_451 N_A_750_21#_c_599_n N_VPWR_c_867_n 0.0117184f $X=6.685 $Y=1.41 $X2=0
+ $Y2=0
cc_452 N_A_750_21#_c_600_n N_VPWR_c_867_n 0.0127538f $X=7.155 $Y=1.41 $X2=0
+ $Y2=0
cc_453 N_A_750_21#_c_601_n N_VPWR_c_867_n 0.00272145f $X=4.55 $Y=1.7 $X2=0 $Y2=0
cc_454 N_A_750_21#_c_616_p N_VPWR_c_867_n 0.0111526f $X=5.025 $Y=1.7 $X2=0 $Y2=0
cc_455 N_A_750_21#_c_613_p N_VPWR_c_867_n 0.00495438f $X=5.175 $Y=1.7 $X2=0
+ $Y2=0
cc_456 N_A_750_21#_c_586_n N_VPWR_c_885_n 0.00667791f $X=3.9 $Y=1.99 $X2=0 $Y2=0
cc_457 N_A_750_21#_c_586_n N_VPWR_c_886_n 0.0102041f $X=3.9 $Y=1.99 $X2=0 $Y2=0
cc_458 N_A_750_21#_c_601_n N_VPWR_c_886_n 0.03463f $X=4.55 $Y=1.7 $X2=0 $Y2=0
cc_459 N_A_750_21#_c_587_n N_Q_c_990_n 0.00532189f $X=5.77 $Y=0.995 $X2=0 $Y2=0
cc_460 N_A_750_21#_c_588_n N_Q_c_990_n 0.00878305f $X=6.19 $Y=0.995 $X2=0 $Y2=0
cc_461 N_A_750_21#_c_589_n N_Q_c_990_n 6.28488e-19 $X=6.71 $Y=0.995 $X2=0 $Y2=0
cc_462 N_A_750_21#_c_598_n N_Q_c_993_n 5.79575e-19 $X=6.215 $Y=1.41 $X2=0 $Y2=0
cc_463 N_A_750_21#_c_641_p N_Q_c_993_n 0.0113624f $X=5.555 $Y=1.62 $X2=0 $Y2=0
cc_464 N_A_750_21#_c_603_n N_Q_c_993_n 0.00312313f $X=5.64 $Y=1.535 $X2=0 $Y2=0
cc_465 N_A_750_21#_c_685_p N_Q_c_993_n 0.0175972f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_466 N_A_750_21#_c_595_n N_Q_c_993_n 0.00549457f $X=7.13 $Y=1.202 $X2=0 $Y2=0
cc_467 N_A_750_21#_c_598_n N_Q_c_998_n 0.0146847f $X=6.215 $Y=1.41 $X2=0 $Y2=0
cc_468 N_A_750_21#_c_685_p N_Q_c_998_n 0.00625258f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_469 N_A_750_21#_c_595_n N_Q_c_998_n 0.00224909f $X=7.13 $Y=1.202 $X2=0 $Y2=0
cc_470 N_A_750_21#_c_588_n N_Q_c_986_n 0.00668441f $X=6.19 $Y=0.995 $X2=0 $Y2=0
cc_471 N_A_750_21#_c_685_p N_Q_c_986_n 0.00276009f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_472 N_A_750_21#_c_595_n N_Q_c_986_n 0.00147082f $X=7.13 $Y=1.202 $X2=0 $Y2=0
cc_473 N_A_750_21#_c_587_n N_Q_c_987_n 0.00334627f $X=5.77 $Y=0.995 $X2=0 $Y2=0
cc_474 N_A_750_21#_c_588_n N_Q_c_987_n 0.00262934f $X=6.19 $Y=0.995 $X2=0 $Y2=0
cc_475 N_A_750_21#_c_685_p N_Q_c_987_n 0.0308404f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_476 N_A_750_21#_c_595_n N_Q_c_987_n 0.00230339f $X=7.13 $Y=1.202 $X2=0 $Y2=0
cc_477 N_A_750_21#_c_588_n N_Q_c_1008_n 5.66668e-19 $X=6.19 $Y=0.995 $X2=0 $Y2=0
cc_478 N_A_750_21#_c_589_n N_Q_c_1008_n 0.00668676f $X=6.71 $Y=0.995 $X2=0 $Y2=0
cc_479 N_A_750_21#_c_590_n N_Q_c_1008_n 0.00550646f $X=7.13 $Y=0.995 $X2=0 $Y2=0
cc_480 N_A_750_21#_c_588_n N_Q_c_988_n 0.0011926f $X=6.19 $Y=0.995 $X2=0 $Y2=0
cc_481 N_A_750_21#_c_598_n N_Q_c_988_n 0.00107237f $X=6.215 $Y=1.41 $X2=0 $Y2=0
cc_482 N_A_750_21#_c_599_n N_Q_c_988_n 0.0164448f $X=6.685 $Y=1.41 $X2=0 $Y2=0
cc_483 N_A_750_21#_c_589_n N_Q_c_988_n 0.0116647f $X=6.71 $Y=0.995 $X2=0 $Y2=0
cc_484 N_A_750_21#_c_590_n N_Q_c_988_n 0.00808017f $X=7.13 $Y=0.995 $X2=0 $Y2=0
cc_485 N_A_750_21#_c_600_n N_Q_c_988_n 0.00673489f $X=7.155 $Y=1.41 $X2=0 $Y2=0
cc_486 N_A_750_21#_c_685_p N_Q_c_988_n 0.0209934f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_487 N_A_750_21#_c_595_n N_Q_c_988_n 0.0821528f $X=7.13 $Y=1.202 $X2=0 $Y2=0
cc_488 N_A_750_21#_c_598_n N_Q_c_1019_n 5.91934e-19 $X=6.215 $Y=1.41 $X2=0 $Y2=0
cc_489 N_A_750_21#_c_599_n N_Q_c_1019_n 0.0100233f $X=6.685 $Y=1.41 $X2=0 $Y2=0
cc_490 N_A_750_21#_c_600_n N_Q_c_1019_n 0.00897418f $X=7.155 $Y=1.41 $X2=0 $Y2=0
cc_491 N_A_750_21#_c_597_n N_Q_c_1022_n 0.00317976f $X=5.745 $Y=1.41 $X2=0 $Y2=0
cc_492 N_A_750_21#_c_598_n N_Q_c_1022_n 0.00236301f $X=6.215 $Y=1.41 $X2=0 $Y2=0
cc_493 N_A_750_21#_c_598_n N_Q_c_1024_n 0.00239814f $X=6.215 $Y=1.41 $X2=0 $Y2=0
cc_494 N_A_750_21#_c_598_n N_Q_c_1025_n 0.00157772f $X=6.215 $Y=1.41 $X2=0 $Y2=0
cc_495 N_A_750_21#_c_685_p N_Q_c_1025_n 7.2795e-19 $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_496 N_A_750_21#_c_595_n N_Q_c_1025_n 8.10024e-19 $X=7.13 $Y=1.202 $X2=0 $Y2=0
cc_497 N_A_750_21#_c_598_n N_Q_c_1028_n 0.00365284f $X=6.215 $Y=1.41 $X2=0 $Y2=0
cc_498 N_A_750_21#_c_599_n N_Q_c_1028_n 5.92409e-19 $X=6.685 $Y=1.41 $X2=0 $Y2=0
cc_499 N_A_750_21#_c_641_p N_Q_c_1028_n 0.00319203f $X=5.555 $Y=1.62 $X2=0 $Y2=0
cc_500 N_A_750_21#_M1001_g N_VGND_c_1060_n 0.0114443f $X=3.825 $Y=0.445 $X2=0
+ $Y2=0
cc_501 N_A_750_21#_c_591_n N_VGND_c_1060_n 0.0222896f $X=4.62 $Y=0.38 $X2=0
+ $Y2=0
cc_502 N_A_750_21#_c_587_n N_VGND_c_1061_n 0.00633937f $X=5.77 $Y=0.995 $X2=0
+ $Y2=0
cc_503 N_A_750_21#_c_593_n N_VGND_c_1061_n 0.00572123f $X=5.725 $Y=1.2 $X2=0
+ $Y2=0
cc_504 N_A_750_21#_c_595_n N_VGND_c_1061_n 0.00117803f $X=7.13 $Y=1.202 $X2=0
+ $Y2=0
cc_505 N_A_750_21#_c_588_n N_VGND_c_1062_n 0.00376004f $X=6.19 $Y=0.995 $X2=0
+ $Y2=0
cc_506 N_A_750_21#_c_589_n N_VGND_c_1062_n 0.00163598f $X=6.71 $Y=0.995 $X2=0
+ $Y2=0
cc_507 N_A_750_21#_c_595_n N_VGND_c_1062_n 6.17468e-19 $X=7.13 $Y=1.202 $X2=0
+ $Y2=0
cc_508 N_A_750_21#_c_590_n N_VGND_c_1063_n 0.0031902f $X=7.13 $Y=0.995 $X2=0
+ $Y2=0
cc_509 N_A_750_21#_c_591_n N_VGND_c_1064_n 0.0209274f $X=4.62 $Y=0.38 $X2=0
+ $Y2=0
cc_510 N_A_750_21#_c_587_n N_VGND_c_1066_n 0.00541359f $X=5.77 $Y=0.995 $X2=0
+ $Y2=0
cc_511 N_A_750_21#_c_588_n N_VGND_c_1066_n 0.00397237f $X=6.19 $Y=0.995 $X2=0
+ $Y2=0
cc_512 N_A_750_21#_c_589_n N_VGND_c_1068_n 0.00424308f $X=6.71 $Y=0.995 $X2=0
+ $Y2=0
cc_513 N_A_750_21#_c_590_n N_VGND_c_1068_n 0.00541359f $X=7.13 $Y=0.995 $X2=0
+ $Y2=0
cc_514 N_A_750_21#_M1001_g N_VGND_c_1072_n 0.0046653f $X=3.825 $Y=0.445 $X2=0
+ $Y2=0
cc_515 N_A_750_21#_M1017_s N_VGND_c_1074_n 0.00209319f $X=4.495 $Y=0.235 $X2=0
+ $Y2=0
cc_516 N_A_750_21#_M1001_g N_VGND_c_1074_n 0.00783311f $X=3.825 $Y=0.445 $X2=0
+ $Y2=0
cc_517 N_A_750_21#_c_587_n N_VGND_c_1074_n 0.00987199f $X=5.77 $Y=0.995 $X2=0
+ $Y2=0
cc_518 N_A_750_21#_c_588_n N_VGND_c_1074_n 0.00581468f $X=6.19 $Y=0.995 $X2=0
+ $Y2=0
cc_519 N_A_750_21#_c_589_n N_VGND_c_1074_n 0.0059764f $X=6.71 $Y=0.995 $X2=0
+ $Y2=0
cc_520 N_A_750_21#_c_590_n N_VGND_c_1074_n 0.0106102f $X=7.13 $Y=0.995 $X2=0
+ $Y2=0
cc_521 N_A_750_21#_c_591_n N_VGND_c_1074_n 0.0123993f $X=4.62 $Y=0.38 $X2=0
+ $Y2=0
cc_522 N_A_604_47#_M1017_g N_RESET_B_c_833_n 0.0427647f $X=4.83 $Y=0.56
+ $X2=-0.19 $Y2=-0.24
cc_523 N_A_604_47#_c_750_n N_RESET_B_c_834_n 0.0183539f $X=4.805 $Y=1.41 $X2=0
+ $Y2=0
cc_524 N_A_604_47#_M1017_g N_RESET_B_c_834_n 0.0213675f $X=4.83 $Y=0.56 $X2=0
+ $Y2=0
cc_525 N_A_604_47#_c_744_n N_RESET_B_c_834_n 0.00398928f $X=4.805 $Y=1.25 $X2=0
+ $Y2=0
cc_526 N_A_604_47#_M1017_g RESET_B 0.00402529f $X=4.83 $Y=0.56 $X2=0 $Y2=0
cc_527 N_A_604_47#_c_744_n RESET_B 0.00387184f $X=4.805 $Y=1.25 $X2=0 $Y2=0
cc_528 N_A_604_47#_c_750_n N_VPWR_c_870_n 5.07375e-19 $X=4.805 $Y=1.41 $X2=0
+ $Y2=0
cc_529 N_A_604_47#_c_750_n N_VPWR_c_873_n 0.00674404f $X=4.805 $Y=1.41 $X2=0
+ $Y2=0
cc_530 N_A_604_47#_M1021_d N_VPWR_c_867_n 0.00194144f $X=3.04 $Y=2.065 $X2=0
+ $Y2=0
cc_531 N_A_604_47#_c_750_n N_VPWR_c_867_n 0.00838474f $X=4.805 $Y=1.41 $X2=0
+ $Y2=0
cc_532 N_A_604_47#_c_755_n N_VPWR_c_867_n 0.0194526f $X=3.68 $Y=2.275 $X2=0
+ $Y2=0
cc_533 N_A_604_47#_c_755_n N_VPWR_c_885_n 0.0311316f $X=3.68 $Y=2.275 $X2=0
+ $Y2=0
cc_534 N_A_604_47#_c_750_n N_VPWR_c_886_n 0.00365563f $X=4.805 $Y=1.41 $X2=0
+ $Y2=0
cc_535 N_A_604_47#_c_755_n A_702_413# 0.00588737f $X=3.68 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_536 N_A_604_47#_c_752_n A_702_413# 0.00114824f $X=3.765 $Y=2.165 $X2=-0.19
+ $Y2=-0.24
cc_537 N_A_604_47#_M1017_g N_VGND_c_1060_n 0.00210532f $X=4.83 $Y=0.56 $X2=0
+ $Y2=0
cc_538 N_A_604_47#_c_759_n N_VGND_c_1060_n 0.0198459f $X=3.49 $Y=0.422 $X2=0
+ $Y2=0
cc_539 N_A_604_47#_c_745_n N_VGND_c_1060_n 0.00279232f $X=3.575 $Y=0.995 $X2=0
+ $Y2=0
cc_540 N_A_604_47#_c_747_n N_VGND_c_1060_n 0.0141331f $X=4.295 $Y=1.16 $X2=0
+ $Y2=0
cc_541 N_A_604_47#_c_748_n N_VGND_c_1060_n 7.94156e-19 $X=4.295 $Y=1.16 $X2=0
+ $Y2=0
cc_542 N_A_604_47#_M1017_g N_VGND_c_1064_n 0.00541359f $X=4.83 $Y=0.56 $X2=0
+ $Y2=0
cc_543 N_A_604_47#_c_759_n N_VGND_c_1072_n 0.0313331f $X=3.49 $Y=0.422 $X2=0
+ $Y2=0
cc_544 N_A_604_47#_M1015_d N_VGND_c_1074_n 0.0030893f $X=3.02 $Y=0.235 $X2=0
+ $Y2=0
cc_545 N_A_604_47#_M1017_g N_VGND_c_1074_n 0.0110154f $X=4.83 $Y=0.56 $X2=0
+ $Y2=0
cc_546 N_A_604_47#_c_759_n N_VGND_c_1074_n 0.0224738f $X=3.49 $Y=0.422 $X2=0
+ $Y2=0
cc_547 N_A_604_47#_c_759_n A_708_47# 0.0032618f $X=3.49 $Y=0.422 $X2=-0.19
+ $Y2=-0.24
cc_548 N_A_604_47#_c_745_n A_708_47# 8.90683e-19 $X=3.575 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_549 N_RESET_B_c_834_n N_VPWR_c_870_n 0.00755919f $X=5.275 $Y=1.41 $X2=0 $Y2=0
cc_550 N_RESET_B_c_834_n N_VPWR_c_938_n 0.00315342f $X=5.275 $Y=1.41 $X2=0 $Y2=0
cc_551 N_RESET_B_c_834_n N_VPWR_c_873_n 0.00622633f $X=5.275 $Y=1.41 $X2=0 $Y2=0
cc_552 N_RESET_B_c_834_n N_VPWR_c_867_n 0.0105052f $X=5.275 $Y=1.41 $X2=0 $Y2=0
cc_553 N_RESET_B_c_833_n N_Q_c_987_n 2.45402e-19 $X=5.235 $Y=0.995 $X2=0 $Y2=0
cc_554 N_RESET_B_c_833_n N_VGND_c_1061_n 0.00332414f $X=5.235 $Y=0.995 $X2=0
+ $Y2=0
cc_555 N_RESET_B_c_834_n N_VGND_c_1061_n 0.00165613f $X=5.275 $Y=1.41 $X2=0
+ $Y2=0
cc_556 RESET_B N_VGND_c_1061_n 0.00340918f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_557 N_RESET_B_c_833_n N_VGND_c_1064_n 0.00585385f $X=5.235 $Y=0.995 $X2=0
+ $Y2=0
cc_558 N_RESET_B_c_833_n N_VGND_c_1074_n 0.0107732f $X=5.235 $Y=0.995 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_867_n A_503_369# 0.00493898f $X=7.59 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_560 N_VPWR_c_867_n A_702_413# 0.00249044f $X=7.59 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_561 N_VPWR_c_867_n N_Q_M1002_d 0.00231261f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_562 N_VPWR_c_867_n N_Q_M1011_d 0.00231261f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_563 N_VPWR_M1004_s N_Q_c_998_n 0.00100055f $X=6.305 $Y=1.485 $X2=0 $Y2=0
cc_564 N_VPWR_c_871_n N_Q_c_998_n 0.00346194f $X=6.45 $Y=2 $X2=0 $Y2=0
cc_565 N_VPWR_M1004_s N_Q_c_988_n 0.00147181f $X=6.305 $Y=1.485 $X2=0 $Y2=0
cc_566 N_VPWR_c_871_n N_Q_c_988_n 0.0119915f $X=6.45 $Y=2 $X2=0 $Y2=0
cc_567 N_VPWR_c_877_n N_Q_c_1019_n 0.0189467f $X=7.255 $Y=2.72 $X2=0 $Y2=0
cc_568 N_VPWR_c_867_n N_Q_c_1019_n 0.0123132f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_569 N_VPWR_c_875_n N_Q_c_1022_n 0.0188482f $X=6.315 $Y=2.72 $X2=0 $Y2=0
cc_570 N_VPWR_c_867_n N_Q_c_1022_n 0.0122778f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_571 N_VPWR_c_872_n N_VGND_c_1063_n 0.00621752f $X=7.39 $Y=1.66 $X2=0 $Y2=0
cc_572 N_Q_c_986_n N_VGND_M1007_s 0.00131825f $X=6.405 $Y=0.82 $X2=0 $Y2=0
cc_573 N_Q_c_988_n N_VGND_M1007_s 0.00191449f $X=6.92 $Y=1.665 $X2=0 $Y2=0
cc_574 N_Q_c_990_n N_VGND_c_1062_n 0.0224895f $X=5.98 $Y=0.38 $X2=0 $Y2=0
cc_575 N_Q_c_986_n N_VGND_c_1062_n 0.00224175f $X=6.405 $Y=0.82 $X2=0 $Y2=0
cc_576 N_Q_c_988_n N_VGND_c_1062_n 0.014999f $X=6.92 $Y=1.665 $X2=0 $Y2=0
cc_577 N_Q_c_988_n N_VGND_c_1063_n 5.02209e-19 $X=6.92 $Y=1.665 $X2=0 $Y2=0
cc_578 N_Q_c_990_n N_VGND_c_1066_n 0.0222529f $X=5.98 $Y=0.38 $X2=0 $Y2=0
cc_579 N_Q_c_986_n N_VGND_c_1066_n 0.00208744f $X=6.405 $Y=0.82 $X2=0 $Y2=0
cc_580 N_Q_c_1008_n N_VGND_c_1068_n 0.0189039f $X=6.92 $Y=0.38 $X2=0 $Y2=0
cc_581 N_Q_c_988_n N_VGND_c_1068_n 0.00210549f $X=6.92 $Y=1.665 $X2=0 $Y2=0
cc_582 N_Q_M1000_d N_VGND_c_1074_n 0.00215201f $X=5.845 $Y=0.235 $X2=0 $Y2=0
cc_583 N_Q_M1010_d N_VGND_c_1074_n 0.00215201f $X=6.785 $Y=0.235 $X2=0 $Y2=0
cc_584 N_Q_c_990_n N_VGND_c_1074_n 0.0139016f $X=5.98 $Y=0.38 $X2=0 $Y2=0
cc_585 N_Q_c_986_n N_VGND_c_1074_n 0.00447392f $X=6.405 $Y=0.82 $X2=0 $Y2=0
cc_586 N_Q_c_1008_n N_VGND_c_1074_n 0.0122217f $X=6.92 $Y=0.38 $X2=0 $Y2=0
cc_587 N_Q_c_988_n N_VGND_c_1074_n 0.00485861f $X=6.92 $Y=1.665 $X2=0 $Y2=0
cc_588 N_VGND_c_1074_n A_500_47# 0.0121316f $X=7.59 $Y=0 $X2=-0.19 $Y2=-0.24
cc_589 N_VGND_c_1074_n A_708_47# 0.00481582f $X=7.59 $Y=0 $X2=-0.19 $Y2=-0.24
cc_590 N_VGND_c_1074_n A_981_47# 0.0109001f $X=7.59 $Y=0 $X2=-0.19 $Y2=-0.24
