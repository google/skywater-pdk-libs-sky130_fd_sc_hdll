# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a31o_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.995000 2.275000 1.655000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 0.995000 1.815000 1.655000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 0.995000 1.340000 1.325000 ;
        RECT 1.075000 1.325000 1.340000 1.655000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 0.995000 2.745000 1.655000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.447300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.300000 0.425000 0.810000 ;
        RECT 0.095000 0.810000 0.285000 1.575000 ;
        RECT 0.095000 1.575000 0.425000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.455000  0.995000 0.815000 1.325000 ;
      RECT 0.605000  0.085000 0.935000 0.485000 ;
      RECT 0.645000  0.655000 3.085000 0.825000 ;
      RECT 0.645000  0.825000 0.815000 0.995000 ;
      RECT 0.645000  1.495000 0.895000 2.635000 ;
      RECT 1.085000  1.825000 2.525000 1.995000 ;
      RECT 1.085000  1.995000 1.385000 2.415000 ;
      RECT 1.665000  2.165000 1.995000 2.635000 ;
      RECT 2.125000  0.315000 2.505000 0.655000 ;
      RECT 2.275000  1.995000 2.525000 2.415000 ;
      RECT 2.725000  0.085000 3.055000 0.485000 ;
      RECT 2.755000  1.825000 3.085000 2.425000 ;
      RECT 2.915000  0.825000 3.085000 1.825000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a31o_1
END LIBRARY
