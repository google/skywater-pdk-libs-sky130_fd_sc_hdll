* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nor4_8 A B C D VGND VNB VPB VPWR Y
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_1635_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_869_297# C a_1635_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_869_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VGND D Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_27_297# B a_869_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 Y D a_1635_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_1635_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 a_1635_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 a_869_297# C a_1635_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 a_1635_297# C a_869_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 a_1635_297# C a_869_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X30 a_27_297# B a_869_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X31 Y D a_1635_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X32 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 a_869_297# C a_1635_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X34 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 Y D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X38 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X40 Y D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X41 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X42 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X43 Y D a_1635_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X44 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X45 a_869_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X46 VGND D Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X47 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X48 a_27_297# B a_869_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X49 a_869_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X50 a_869_297# C a_1635_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X51 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X52 a_869_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X53 a_27_297# B a_869_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X54 a_1635_297# C a_869_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X55 Y D a_1635_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X56 a_1635_297# C a_869_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X57 VGND D Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X58 a_1635_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X59 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X60 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X61 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X62 VGND D Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X63 Y D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
