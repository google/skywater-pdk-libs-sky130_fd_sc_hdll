* File: sky130_fd_sc_hdll__o31ai_2.spice
* Created: Wed Sep  2 08:46:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o31ai_2.pex.spice"
.subckt sky130_fd_sc_hdll__o31ai_2  VNB VPB A1 A2 A3 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A1_M1004_g N_A_27_47#_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.2145 PD=0.97 PS=1.96 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.3
+ SB=75004.2 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1004_d N_A1_M1015_g N_A_27_47#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1011 N_A_27_47#_M1015_s N_A2_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.247 PD=0.92 PS=1.41 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.1
+ SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1014 N_A_27_47#_M1014_d N_A2_M1014_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.247 PD=1.02 PS=1.41 NRD=6.456 NRS=17.532 M=1 R=4.33333
+ SA=75002.1 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1002 N_A_27_47#_M1014_d N_A3_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.15275 PD=1.02 PS=1.12 NRD=10.152 NRS=11.988 M=1 R=4.33333
+ SA=75002.6 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1003 N_A_27_47#_M1003_d N_A3_M1003_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.15275 PD=0.92 PS=1.12 NRD=0 NRS=23.076 M=1 R=4.33333
+ SA=75003.2 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1007 N_Y_M1007_d N_B1_M1007_g N_A_27_47#_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.143 AS=0.08775 PD=1.09 PS=0.92 NRD=23.076 NRS=0 M=1 R=4.33333 SA=75003.6
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1008 N_Y_M1007_d N_B1_M1008_g N_A_27_47#_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.143 AS=0.20475 PD=1.09 PS=1.93 NRD=6.456 NRS=9.228 M=1 R=4.33333
+ SA=75004.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g N_A_27_297#_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1000_d N_A1_M1013_g N_A_27_297#_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1006 N_A_27_297#_M1013_s N_A2_M1006_g N_A_309_297#_M1006_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1009 N_A_27_297#_M1009_d N_A2_M1009_g N_A_309_297#_M1006_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1005 N_Y_M1005_d N_A3_M1005_g N_A_309_297#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.29 AS=0.145 PD=2.58 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1012 N_Y_M1012_d N_A3_M1012_g N_A_309_297#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_B1_M1001_g N_Y_M1012_d VPB PHIGHVT L=0.18 W=1 AD=0.205
+ AS=0.145 PD=1.41 PS=1.29 NRD=16.7253 NRS=0.9653 M=1 R=5.55556 SA=90001.1
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1001_d N_B1_M1010_g N_Y_M1010_s VPB PHIGHVT L=0.18 W=1 AD=0.205
+ AS=0.27 PD=1.41 PS=2.54 NRD=8.8453 NRS=0.9653 M=1 R=5.55556 SA=90001.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.7312 P=14.09
*
.include "sky130_fd_sc_hdll__o31ai_2.pxi.spice"
*
.ends
*
*
