* NGSPICE file created from sky130_fd_sc_hdll__a21boi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 a_228_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.2e+12p pd=1.04e+07u as=7.055e+11p ps=6.57e+06u
M1001 VPWR A2 a_228_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_228_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_228_297# a_61_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1004 Y A1 a_529_47# VNB nshort w=650000u l=150000u
+  ad=4.225e+11p pd=3.9e+06u as=1.365e+11p ps=1.72e+06u
M1005 Y a_61_47# a_228_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_61_47# Y VNB nshort w=650000u l=150000u
+  ad=8.845e+11p pd=6.71e+06u as=0p ps=0u
M1007 a_61_47# B1_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.155e+11p pd=1.39e+06u as=0p ps=0u
M1008 VPWR A1 a_228_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_529_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B1_N a_61_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1011 a_697_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=0p ps=0u
M1012 Y a_61_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A2 a_697_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

