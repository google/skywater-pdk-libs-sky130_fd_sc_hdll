* File: sky130_fd_sc_hdll__o2bb2ai_1.pex.spice
* Created: Wed Sep  2 08:46:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_1%A1_N 1 3 4 6 7 12
c23 7 0 1.85093e-19 $X=0.23 $Y=1.19
r24 12 13 3.31956 $w=3.63e-07 $l=2.5e-08 $layer=POLY_cond $X=0.51 $Y=1.202
+ $X2=0.535 $Y2=1.202
r25 10 12 31.8678 $w=3.63e-07 $l=2.4e-07 $layer=POLY_cond $X=0.27 $Y=1.202
+ $X2=0.51 $Y2=1.202
r26 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r27 4 13 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.535 $Y=0.995
+ $X2=0.535 $Y2=1.202
r28 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.535 $Y=0.995
+ $X2=0.535 $Y2=0.56
r29 1 12 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.41
+ $X2=0.51 $Y2=1.202
r30 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.51 $Y=1.41 $X2=0.51
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_1%A2_N 1 3 4 6 9 13 17
c36 4 0 2.65272e-19 $X=0.98 $Y=1.41
r37 13 17 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.015 $Y=1.16
+ $X2=0.715 $Y2=1.16
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.015
+ $Y=1.16 $X2=1.015 $Y2=1.16
r39 9 17 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.69 $Y=1.16
+ $X2=0.715 $Y2=1.16
r40 4 12 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=1.015 $Y2=1.16
r41 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.98 $Y=1.41 $X2=0.98
+ $Y2=1.985
r42 1 12 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=1.015 $Y2=1.16
r43 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_1%A_120_297# 1 2 7 9 10 12 13 14 17 19 20
+ 24 26 30 32
c64 26 0 2.15831e-19 $X=1.165 $Y=0.39
c65 13 0 1.06764e-19 $X=1.78 $Y=1.16
c66 7 0 1.69324e-19 $X=1.88 $Y=1.41
r67 30 33 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=1.16
+ $X2=1.425 $Y2=1.325
r68 30 32 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=1.16
+ $X2=1.425 $Y2=0.995
r69 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.495
+ $Y=1.16 $X2=1.495 $Y2=1.16
r70 28 32 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.355 $Y=0.825
+ $X2=1.355 $Y2=0.995
r71 26 28 15.9071 $w=4.38e-07 $l=4.35e-07 $layer=LI1_cond $X=1.22 $Y=0.39
+ $X2=1.22 $Y2=0.825
r72 24 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.355 $Y=1.495
+ $X2=1.355 $Y2=1.325
r73 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.27 $Y=1.58
+ $X2=1.355 $Y2=1.495
r74 19 20 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.27 $Y=1.58 $X2=0.87
+ $Y2=1.58
r75 15 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.745 $Y=1.665
+ $X2=0.87 $Y2=1.58
r76 15 17 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.745 $Y=1.665
+ $X2=0.745 $Y2=1.96
r77 13 31 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=1.78 $Y=1.16
+ $X2=1.495 $Y2=1.16
r78 13 14 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.78 $Y=1.16
+ $X2=1.88 $Y2=1.202
r79 10 14 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=1.905 $Y=0.995
+ $X2=1.88 $Y2=1.202
r80 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.905 $Y=0.995
+ $X2=1.905 $Y2=0.56
r81 7 14 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=1.88 $Y=1.41
+ $X2=1.88 $Y2=1.202
r82 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.88 $Y=1.41 $X2=1.88
+ $Y2=1.985
r83 2 17 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.6
+ $Y=1.485 $X2=0.745 $Y2=1.96
r84 1 26 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.03
+ $Y=0.235 $X2=1.165 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_1%B2 1 3 4 6 7 13
c42 13 0 1.69324e-19 $X=2.53 $Y=1.53
c43 1 0 1.80417e-19 $X=2.37 $Y=1.41
r44 12 13 18.3 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.53 $Y=1.275 $X2=2.53
+ $Y2=1.53
r45 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.335
+ $Y=1.16 $X2=2.335 $Y2=1.16
r46 7 12 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.445 $Y=1.175
+ $X2=2.53 $Y2=1.275
r47 7 9 6.1 $w=1.98e-07 $l=1.1e-07 $layer=LI1_cond $X=2.445 $Y=1.175 $X2=2.335
+ $Y2=1.175
r48 4 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.395 $Y=0.995
+ $X2=2.335 $Y2=1.16
r49 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.395 $Y=0.995
+ $X2=2.395 $Y2=0.56
r50 1 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.37 $Y=1.41
+ $X2=2.335 $Y2=1.16
r51 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.37 $Y=1.41 $X2=2.37
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_1%B1 1 3 4 6 7 10 13
c26 13 0 1.80417e-19 $X=3.08 $Y=1.16
r27 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.08
+ $Y=1.16 $X2=3.08 $Y2=1.16
r28 10 12 31.8678 $w=3.63e-07 $l=2.4e-07 $layer=POLY_cond $X=2.84 $Y=1.202
+ $X2=3.08 $Y2=1.202
r29 9 10 3.31956 $w=3.63e-07 $l=2.5e-08 $layer=POLY_cond $X=2.815 $Y=1.202
+ $X2=2.84 $Y2=1.202
r30 7 13 4.75325 $w=2.08e-07 $l=9e-08 $layer=LI1_cond $X=2.99 $Y=1.18 $X2=3.08
+ $Y2=1.18
r31 4 10 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.84 $Y=1.41
+ $X2=2.84 $Y2=1.202
r32 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.84 $Y=1.41 $X2=2.84
+ $Y2=1.985
r33 1 9 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.815 $Y=0.995
+ $X2=2.815 $Y2=1.202
r34 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.815 $Y=0.995
+ $X2=2.815 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_1%VPWR 1 2 3 10 12 16 20 24 28 30 37 38 44
+ 49
r44 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 45 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r46 44 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r47 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r48 38 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r49 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r50 35 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.2 $Y=2.72
+ $X2=3.075 $Y2=2.72
r51 35 37 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.2 $Y=2.72 $X2=3.45
+ $Y2=2.72
r52 34 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 34 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r54 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r55 31 44 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=1.78 $Y=2.72
+ $X2=1.435 $Y2=2.72
r56 31 33 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.78 $Y=2.72
+ $X2=2.07 $Y2=2.72
r57 30 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.95 $Y=2.72
+ $X2=3.075 $Y2=2.72
r58 30 33 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=2.95 $Y=2.72
+ $X2=2.07 $Y2=2.72
r59 28 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r60 28 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r61 24 27 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=3.075 $Y=1.63
+ $X2=3.075 $Y2=2.31
r62 22 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=2.635
+ $X2=3.075 $Y2=2.72
r63 22 27 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=3.075 $Y=2.635
+ $X2=3.075 $Y2=2.31
r64 18 44 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=2.635
+ $X2=1.435 $Y2=2.72
r65 18 20 11.7008 $w=6.88e-07 $l=6.75e-07 $layer=LI1_cond $X=1.435 $Y=2.635
+ $X2=1.435 $Y2=1.96
r66 17 41 3.96842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=2.72 $X2=0.2
+ $Y2=2.72
r67 16 44 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=1.09 $Y=2.72
+ $X2=1.435 $Y2=2.72
r68 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.09 $Y=2.72 $X2=0.4
+ $Y2=2.72
r69 12 15 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.275 $Y=1.63
+ $X2=0.275 $Y2=2.31
r70 10 41 3.17474 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=0.275 $Y=2.635
+ $X2=0.2 $Y2=2.72
r71 10 15 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=0.275 $Y=2.635
+ $X2=0.275 $Y2=2.31
r72 3 27 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.485 $X2=3.075 $Y2=2.31
r73 3 24 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.485 $X2=3.075 $Y2=1.63
r74 2 20 150 $w=1.7e-07 $l=7.35085e-07 $layer=licon1_PDIFF $count=4 $X=1.07
+ $Y=1.485 $X2=1.605 $Y2=1.96
r75 1 15 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=2.31
r76 1 12 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_1%Y 1 2 8 12 17 20
c34 17 0 1.86943e-19 $X=2.112 $Y=1.665
r35 20 25 15.2477 $w=3.23e-07 $l=4.3e-07 $layer=LI1_cond $X=2.112 $Y=1.87
+ $X2=2.112 $Y2=2.3
r36 17 20 7.26926 $w=3.23e-07 $l=2.05e-07 $layer=LI1_cond $X=2.112 $Y=1.665
+ $X2=2.112 $Y2=1.87
r37 14 17 13.9865 $w=2.18e-07 $l=2.67e-07 $layer=LI1_cond $X=1.845 $Y=1.555
+ $X2=2.112 $Y2=1.555
r38 10 12 4.80185 $w=3.58e-07 $l=1.5e-07 $layer=LI1_cond $X=1.695 $Y=0.61
+ $X2=1.845 $Y2=0.61
r39 8 14 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.845 $Y=1.445
+ $X2=1.845 $Y2=1.555
r40 7 12 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.845 $Y=0.79
+ $X2=1.845 $Y2=0.61
r41 7 8 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.845 $Y=0.79
+ $X2=1.845 $Y2=1.445
r42 2 25 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.97
+ $Y=1.485 $X2=2.115 $Y2=2.3
r43 2 17 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.97
+ $Y=1.485 $X2=2.115 $Y2=1.62
r44 1 10 182 $w=1.7e-07 $l=4.32262e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.235 $X2=1.695 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_1%VGND 1 2 7 9 13 15 17 24 25 31
r42 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r43 25 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r44 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r45 22 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.605
+ $Y2=0
r46 22 24 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=3.45
+ $Y2=0
r47 21 32 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r48 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r49 18 28 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r50 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r51 17 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=0 $X2=2.605
+ $Y2=0
r52 17 20 119.39 $w=1.68e-07 $l=1.83e-06 $layer=LI1_cond $X=2.52 $Y=0 $X2=0.69
+ $Y2=0
r53 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r54 15 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r55 11 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=0.085
+ $X2=2.605 $Y2=0
r56 11 13 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.605 $Y=0.085
+ $X2=2.605 $Y2=0.39
r57 7 28 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.212 $Y2=0
r58 7 9 10.4924 $w=3.33e-07 $l=3.05e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.39
r59 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.47
+ $Y=0.235 $X2=2.605 $Y2=0.39
r60 1 9 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_1%A_396_47# 1 2 9 11 12 15
c32 12 0 3.28448e-20 $X=2.35 $Y=0.815
c33 9 0 1.82987e-19 $X=2.185 $Y=0.605
r34 13 15 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.05 $Y=0.725
+ $X2=3.05 $Y2=0.39
r35 11 13 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=2.86 $Y=0.815
+ $X2=3.05 $Y2=0.725
r36 11 12 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.86 $Y=0.815
+ $X2=2.35 $Y2=0.815
r37 7 12 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=2.225 $Y=0.725
+ $X2=2.35 $Y2=0.815
r38 7 9 5.53173 $w=2.48e-07 $l=1.2e-07 $layer=LI1_cond $X=2.225 $Y=0.725
+ $X2=2.225 $Y2=0.605
r39 2 15 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=2.89
+ $Y=0.235 $X2=3.075 $Y2=0.39
r40 1 9 182 $w=1.7e-07 $l=4.61248e-07 $layer=licon1_NDIFF $count=1 $X=1.98
+ $Y=0.235 $X2=2.185 $Y2=0.605
.ends

