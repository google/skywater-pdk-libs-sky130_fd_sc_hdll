* File: sky130_fd_sc_hdll__clkinv_12.pxi.spice
* Created: Wed Sep  2 08:26:01 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKINV_12%A N_A_c_142_n N_A_M1000_g N_A_c_143_n
+ N_A_M1001_g N_A_c_144_n N_A_M1003_g N_A_c_145_n N_A_M1004_g N_A_M1002_g
+ N_A_M1006_g N_A_c_146_n N_A_M1005_g N_A_c_147_n N_A_M1007_g N_A_M1009_g
+ N_A_M1010_g N_A_c_148_n N_A_M1008_g N_A_c_149_n N_A_M1011_g N_A_M1013_g
+ N_A_M1014_g N_A_c_150_n N_A_M1012_g N_A_c_151_n N_A_M1015_g N_A_M1017_g
+ N_A_M1020_g N_A_c_152_n N_A_M1016_g N_A_c_153_n N_A_M1018_g N_A_M1024_g
+ N_A_M1026_g N_A_c_154_n N_A_M1019_g N_A_c_155_n N_A_M1021_g N_A_M1027_g
+ N_A_M1028_g N_A_c_156_n N_A_M1022_g N_A_c_157_n N_A_M1023_g N_A_c_158_n
+ N_A_M1025_g N_A_c_159_n N_A_M1029_g A N_A_c_234_p N_A_c_141_n
+ PM_SKY130_FD_SC_HDLL__CLKINV_12%A
x_PM_SKY130_FD_SC_HDLL__CLKINV_12%VPWR N_VPWR_M1000_d N_VPWR_M1001_d
+ N_VPWR_M1004_d N_VPWR_M1007_d N_VPWR_M1011_d N_VPWR_M1015_d N_VPWR_M1018_d
+ N_VPWR_M1021_d N_VPWR_M1023_d N_VPWR_M1029_d N_VPWR_c_393_n N_VPWR_c_394_n
+ N_VPWR_c_395_n N_VPWR_c_396_n N_VPWR_c_397_n N_VPWR_c_398_n N_VPWR_c_399_n
+ N_VPWR_c_400_n N_VPWR_c_401_n N_VPWR_c_402_n N_VPWR_c_403_n N_VPWR_c_404_n
+ N_VPWR_c_405_n N_VPWR_c_406_n N_VPWR_c_407_n N_VPWR_c_408_n N_VPWR_c_409_n
+ N_VPWR_c_410_n N_VPWR_c_411_n N_VPWR_c_412_n N_VPWR_c_413_n VPWR
+ N_VPWR_c_414_n N_VPWR_c_415_n N_VPWR_c_416_n N_VPWR_c_392_n N_VPWR_c_418_n
+ N_VPWR_c_419_n N_VPWR_c_420_n N_VPWR_c_421_n N_VPWR_c_422_n N_VPWR_c_423_n
+ PM_SKY130_FD_SC_HDLL__CLKINV_12%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKINV_12%Y N_Y_M1002_d N_Y_M1009_d N_Y_M1013_d
+ N_Y_M1017_d N_Y_M1024_d N_Y_M1027_d N_Y_M1000_s N_Y_M1003_s N_Y_M1005_s
+ N_Y_M1008_s N_Y_M1012_s N_Y_M1016_s N_Y_M1019_s N_Y_M1022_s N_Y_M1025_s
+ N_Y_c_545_n N_Y_c_546_n N_Y_c_547_n N_Y_c_568_n N_Y_c_569_n N_Y_c_724_n
+ N_Y_c_570_n N_Y_c_728_n N_Y_c_571_n N_Y_c_548_n N_Y_c_549_n N_Y_c_732_n
+ N_Y_c_572_n N_Y_c_550_n N_Y_c_551_n N_Y_c_736_n N_Y_c_573_n N_Y_c_552_n
+ N_Y_c_553_n N_Y_c_740_n N_Y_c_574_n N_Y_c_554_n N_Y_c_555_n N_Y_c_744_n
+ N_Y_c_575_n N_Y_c_556_n N_Y_c_557_n N_Y_c_748_n N_Y_c_576_n N_Y_c_558_n
+ N_Y_c_559_n N_Y_c_752_n N_Y_c_577_n N_Y_c_756_n N_Y_c_578_n N_Y_c_579_n
+ N_Y_c_560_n N_Y_c_580_n N_Y_c_561_n N_Y_c_581_n N_Y_c_562_n N_Y_c_582_n
+ N_Y_c_563_n N_Y_c_583_n N_Y_c_564_n N_Y_c_584_n N_Y_c_565_n N_Y_c_585_n
+ N_Y_c_586_n Y PM_SKY130_FD_SC_HDLL__CLKINV_12%Y
x_PM_SKY130_FD_SC_HDLL__CLKINV_12%VGND N_VGND_M1002_s N_VGND_M1006_s
+ N_VGND_M1010_s N_VGND_M1014_s N_VGND_M1020_s N_VGND_M1026_s N_VGND_M1028_s
+ N_VGND_c_808_n N_VGND_c_809_n N_VGND_c_810_n N_VGND_c_811_n N_VGND_c_812_n
+ N_VGND_c_813_n N_VGND_c_814_n N_VGND_c_815_n N_VGND_c_816_n VGND
+ N_VGND_c_817_n N_VGND_c_818_n N_VGND_c_819_n N_VGND_c_820_n N_VGND_c_821_n
+ N_VGND_c_822_n N_VGND_c_823_n N_VGND_c_824_n N_VGND_c_825_n N_VGND_c_826_n
+ N_VGND_c_827_n N_VGND_c_828_n PM_SKY130_FD_SC_HDLL__CLKINV_12%VGND
cc_1 VNB N_A_M1002_g 0.0365543f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.445
cc_2 VNB N_A_M1006_g 0.0278467f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=0.445
cc_3 VNB N_A_M1009_g 0.0278467f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=0.445
cc_4 VNB N_A_M1010_g 0.0278467f $X=-0.19 $Y=-0.24 $X2=3.29 $Y2=0.445
cc_5 VNB N_A_M1013_g 0.0278467f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.445
cc_6 VNB N_A_M1014_g 0.0278467f $X=-0.19 $Y=-0.24 $X2=4.23 $Y2=0.445
cc_7 VNB N_A_M1017_g 0.0278467f $X=-0.19 $Y=-0.24 $X2=4.75 $Y2=0.445
cc_8 VNB N_A_M1020_g 0.0278467f $X=-0.19 $Y=-0.24 $X2=5.17 $Y2=0.445
cc_9 VNB N_A_M1024_g 0.0278467f $X=-0.19 $Y=-0.24 $X2=5.69 $Y2=0.445
cc_10 VNB N_A_M1026_g 0.0278467f $X=-0.19 $Y=-0.24 $X2=6.11 $Y2=0.445
cc_11 VNB N_A_M1027_g 0.0278467f $X=-0.19 $Y=-0.24 $X2=6.63 $Y2=0.445
cc_12 VNB N_A_M1028_g 0.0365543f $X=-0.19 $Y=-0.24 $X2=7.05 $Y2=0.445
cc_13 VNB N_A_c_141_n 0.394759f $X=-0.19 $Y=-0.24 $X2=8.015 $Y2=1.202
cc_14 VNB N_VPWR_c_392_n 0.383598f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.202
cc_15 VNB N_Y_c_545_n 0.0240607f $X=-0.19 $Y=-0.24 $X2=4.23 $Y2=0.445
cc_16 VNB N_Y_c_546_n 0.0366113f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_Y_c_547_n 0.0104149f $X=-0.19 $Y=-0.24 $X2=4.255 $Y2=1.41
cc_18 VNB N_Y_c_548_n 6.87798e-19 $X=-0.19 $Y=-0.24 $X2=5.665 $Y2=1.41
cc_19 VNB N_Y_c_549_n 0.00614847f $X=-0.19 $Y=-0.24 $X2=5.665 $Y2=1.985
cc_20 VNB N_Y_c_550_n 6.50236e-19 $X=-0.19 $Y=-0.24 $X2=6.135 $Y2=1.985
cc_21 VNB N_Y_c_551_n 0.00614847f $X=-0.19 $Y=-0.24 $X2=6.605 $Y2=1.41
cc_22 VNB N_Y_c_552_n 6.50236e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_Y_c_553_n 0.00614847f $X=-0.19 $Y=-0.24 $X2=7.075 $Y2=1.985
cc_24 VNB N_Y_c_554_n 6.50236e-19 $X=-0.19 $Y=-0.24 $X2=8.485 $Y2=1.985
cc_25 VNB N_Y_c_555_n 0.00614847f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_Y_c_556_n 6.50236e-19 $X=-0.19 $Y=-0.24 $X2=2.375 $Y2=1.202
cc_27 VNB N_Y_c_557_n 0.00614847f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=1.202
cc_28 VNB N_Y_c_558_n 6.87798e-19 $X=-0.19 $Y=-0.24 $X2=5.195 $Y2=1.202
cc_29 VNB N_Y_c_559_n 0.0377569f $X=-0.19 $Y=-0.24 $X2=5.69 $Y2=1.202
cc_30 VNB N_Y_c_560_n 0.002211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_Y_c_561_n 0.002211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_562_n 0.002211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_Y_c_563_n 0.002211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_Y_c_564_n 0.002211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_Y_c_565_n 0.002211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB Y 0.0225583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_808_n 0.00441949f $X=-0.19 $Y=-0.24 $X2=2.845 $Y2=1.41
cc_38 VNB N_VGND_c_809_n 0.0154684f $X=-0.19 $Y=-0.24 $X2=2.845 $Y2=1.985
cc_39 VNB N_VGND_c_810_n 0.00442069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_811_n 0.0154684f $X=-0.19 $Y=-0.24 $X2=3.29 $Y2=0.445
cc_41 VNB N_VGND_c_812_n 0.00442069f $X=-0.19 $Y=-0.24 $X2=3.315 $Y2=1.985
cc_42 VNB N_VGND_c_813_n 0.0154684f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.41
cc_43 VNB N_VGND_c_814_n 0.00442069f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.445
cc_44 VNB N_VGND_c_815_n 0.0154684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_816_n 0.00441949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_817_n 0.0154684f $X=-0.19 $Y=-0.24 $X2=5.17 $Y2=0.445
cc_47 VNB N_VGND_c_818_n 0.0429047f $X=-0.19 $Y=-0.24 $X2=6.11 $Y2=0.445
cc_48 VNB N_VGND_c_819_n 0.470351f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_820_n 0.035079f $X=-0.19 $Y=-0.24 $X2=6.605 $Y2=1.985
cc_50 VNB N_VGND_c_821_n 0.0321546f $X=-0.19 $Y=-0.24 $X2=6.63 $Y2=0.445
cc_51 VNB N_VGND_c_822_n 0.00631792f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_823_n 0.00631792f $X=-0.19 $Y=-0.24 $X2=7.05 $Y2=0.445
cc_53 VNB N_VGND_c_824_n 0.00631792f $X=-0.19 $Y=-0.24 $X2=7.075 $Y2=1.985
cc_54 VNB N_VGND_c_825_n 0.00631792f $X=-0.19 $Y=-0.24 $X2=7.545 $Y2=1.985
cc_55 VNB N_VGND_c_826_n 0.00631792f $X=-0.19 $Y=-0.24 $X2=8.015 $Y2=1.985
cc_56 VNB N_VGND_c_827_n 0.0154684f $X=-0.19 $Y=-0.24 $X2=4.285 $Y2=1.105
cc_57 VNB N_VGND_c_828_n 0.0321546f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.202
cc_58 VPB N_A_c_142_n 0.0183051f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_59 VPB N_A_c_143_n 0.0158261f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_60 VPB N_A_c_144_n 0.0158451f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_61 VPB N_A_c_145_n 0.0158451f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_62 VPB N_A_c_146_n 0.0158451f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_63 VPB N_A_c_147_n 0.0158451f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_64 VPB N_A_c_148_n 0.0158451f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.41
cc_65 VPB N_A_c_149_n 0.0158451f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_66 VPB N_A_c_150_n 0.0158451f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.41
cc_67 VPB N_A_c_151_n 0.0158451f $X=-0.19 $Y=1.305 $X2=4.725 $Y2=1.41
cc_68 VPB N_A_c_152_n 0.0158451f $X=-0.19 $Y=1.305 $X2=5.195 $Y2=1.41
cc_69 VPB N_A_c_153_n 0.0158451f $X=-0.19 $Y=1.305 $X2=5.665 $Y2=1.41
cc_70 VPB N_A_c_154_n 0.0158451f $X=-0.19 $Y=1.305 $X2=6.135 $Y2=1.41
cc_71 VPB N_A_c_155_n 0.0158451f $X=-0.19 $Y=1.305 $X2=6.605 $Y2=1.41
cc_72 VPB N_A_c_156_n 0.0158451f $X=-0.19 $Y=1.305 $X2=7.075 $Y2=1.41
cc_73 VPB N_A_c_157_n 0.0158245f $X=-0.19 $Y=1.305 $X2=7.545 $Y2=1.41
cc_74 VPB N_A_c_158_n 0.0156225f $X=-0.19 $Y=1.305 $X2=8.015 $Y2=1.41
cc_75 VPB N_A_c_159_n 0.0184001f $X=-0.19 $Y=1.305 $X2=8.485 $Y2=1.41
cc_76 VPB N_A_c_141_n 0.225867f $X=-0.19 $Y=1.305 $X2=8.015 $Y2=1.202
cc_77 VPB N_VPWR_c_393_n 0.0103693f $X=-0.19 $Y=1.305 $X2=3.29 $Y2=0.995
cc_78 VPB N_VPWR_c_394_n 0.0301438f $X=-0.19 $Y=1.305 $X2=3.29 $Y2=0.445
cc_79 VPB N_VPWR_c_395_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.985
cc_80 VPB N_VPWR_c_396_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=3.81 $Y2=0.995
cc_81 VPB N_VPWR_c_397_n 0.0147329f $X=-0.19 $Y=1.305 $X2=3.81 $Y2=0.445
cc_82 VPB N_VPWR_c_398_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=4.23 $Y2=0.445
cc_83 VPB N_VPWR_c_399_n 0.0147329f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.41
cc_84 VPB N_VPWR_c_400_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=4.725 $Y2=1.985
cc_85 VPB N_VPWR_c_401_n 0.0147329f $X=-0.19 $Y=1.305 $X2=4.75 $Y2=0.995
cc_86 VPB N_VPWR_c_402_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=5.17 $Y2=0.995
cc_87 VPB N_VPWR_c_403_n 0.0147329f $X=-0.19 $Y=1.305 $X2=5.17 $Y2=0.445
cc_88 VPB N_VPWR_c_404_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=5.195 $Y2=1.985
cc_89 VPB N_VPWR_c_405_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=5.69 $Y2=0.995
cc_90 VPB N_VPWR_c_406_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=6.11 $Y2=0.995
cc_91 VPB N_VPWR_c_407_n 0.0307803f $X=-0.19 $Y=1.305 $X2=6.135 $Y2=1.41
cc_92 VPB N_VPWR_c_408_n 0.0147329f $X=-0.19 $Y=1.305 $X2=6.605 $Y2=1.41
cc_93 VPB N_VPWR_c_409_n 0.00436868f $X=-0.19 $Y=1.305 $X2=6.605 $Y2=1.985
cc_94 VPB N_VPWR_c_410_n 0.0147329f $X=-0.19 $Y=1.305 $X2=6.63 $Y2=0.995
cc_95 VPB N_VPWR_c_411_n 0.00436868f $X=-0.19 $Y=1.305 $X2=6.63 $Y2=0.445
cc_96 VPB N_VPWR_c_412_n 0.0147329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_413_n 0.00513801f $X=-0.19 $Y=1.305 $X2=7.05 $Y2=0.995
cc_98 VPB N_VPWR_c_414_n 0.0147329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_415_n 0.0147329f $X=-0.19 $Y=1.305 $X2=7.545 $Y2=1.985
cc_100 VPB N_VPWR_c_416_n 0.0121672f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_101 VPB N_VPWR_c_392_n 0.0529516f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=1.202
cc_102 VPB N_VPWR_c_418_n 0.00436868f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.202
cc_103 VPB N_VPWR_c_419_n 0.00436868f $X=-0.19 $Y=1.305 $X2=4.23 $Y2=1.202
cc_104 VPB N_VPWR_c_420_n 0.00436868f $X=-0.19 $Y=1.305 $X2=4.75 $Y2=1.202
cc_105 VPB N_VPWR_c_421_n 0.00436868f $X=-0.19 $Y=1.305 $X2=5.665 $Y2=1.202
cc_106 VPB N_VPWR_c_422_n 0.00436868f $X=-0.19 $Y=1.305 $X2=6.135 $Y2=1.202
cc_107 VPB N_VPWR_c_423_n 0.00436868f $X=-0.19 $Y=1.305 $X2=7.05 $Y2=1.202
cc_108 VPB N_Y_c_545_n 0.00734091f $X=-0.19 $Y=1.305 $X2=4.23 $Y2=0.445
cc_109 VPB N_Y_c_568_n 0.00166909f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.985
cc_110 VPB N_Y_c_569_n 0.00731071f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.985
cc_111 VPB N_Y_c_570_n 0.00181842f $X=-0.19 $Y=1.305 $X2=4.75 $Y2=0.445
cc_112 VPB N_Y_c_571_n 0.00181842f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_Y_c_572_n 0.00181842f $X=-0.19 $Y=1.305 $X2=6.11 $Y2=0.445
cc_114 VPB N_Y_c_573_n 0.00181842f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_Y_c_574_n 0.00181842f $X=-0.19 $Y=1.305 $X2=8.015 $Y2=1.985
cc_116 VPB N_Y_c_575_n 0.00181842f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.202
cc_117 VPB N_Y_c_576_n 0.00181842f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.202
cc_118 VPB N_Y_c_577_n 0.00176637f $X=-0.19 $Y=1.305 $X2=7.075 $Y2=1.202
cc_119 VPB N_Y_c_578_n 0.00163387f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.162
cc_120 VPB N_Y_c_579_n 0.00163387f $X=-0.19 $Y=1.305 $X2=4.37 $Y2=1.162
cc_121 VPB N_Y_c_580_n 0.00163387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_Y_c_581_n 0.00163387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_Y_c_582_n 0.00163387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_Y_c_583_n 0.00163387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_Y_c_584_n 0.00163387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_Y_c_585_n 0.00163387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_Y_c_586_n 0.00101819f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB Y 0.00611616f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 N_A_c_142_n N_VPWR_c_394_n 0.0129769f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_c_143_n N_VPWR_c_394_n 6.03055e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A_c_142_n N_VPWR_c_395_n 6.03055e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A_c_143_n N_VPWR_c_395_n 0.0119993f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A_c_144_n N_VPWR_c_395_n 0.0119993f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_c_145_n N_VPWR_c_395_n 6.03055e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_c_144_n N_VPWR_c_396_n 6.03055e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A_c_145_n N_VPWR_c_396_n 0.0119993f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A_c_146_n N_VPWR_c_396_n 0.0119993f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_c_147_n N_VPWR_c_396_n 6.03055e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_c_146_n N_VPWR_c_397_n 0.00622633f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_c_147_n N_VPWR_c_397_n 0.00622633f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_c_146_n N_VPWR_c_398_n 6.03055e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_c_147_n N_VPWR_c_398_n 0.0119993f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_c_148_n N_VPWR_c_398_n 0.0119993f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_149_n N_VPWR_c_398_n 6.03055e-19 $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_c_148_n N_VPWR_c_399_n 0.00622633f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_c_149_n N_VPWR_c_399_n 0.00622633f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_c_148_n N_VPWR_c_400_n 6.03055e-19 $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_c_149_n N_VPWR_c_400_n 0.0119993f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_c_150_n N_VPWR_c_400_n 0.0119993f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_c_151_n N_VPWR_c_400_n 6.03055e-19 $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_c_150_n N_VPWR_c_401_n 0.00622633f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_c_151_n N_VPWR_c_401_n 0.00622633f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_c_150_n N_VPWR_c_402_n 6.03055e-19 $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_c_151_n N_VPWR_c_402_n 0.0119993f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_c_152_n N_VPWR_c_402_n 0.0119993f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_c_153_n N_VPWR_c_402_n 6.03055e-19 $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_c_152_n N_VPWR_c_403_n 0.00622633f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_c_153_n N_VPWR_c_403_n 0.00622633f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_c_152_n N_VPWR_c_404_n 6.03055e-19 $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A_c_153_n N_VPWR_c_404_n 0.0119993f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A_c_154_n N_VPWR_c_404_n 0.0119993f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_c_155_n N_VPWR_c_404_n 6.03055e-19 $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A_c_154_n N_VPWR_c_405_n 6.03055e-19 $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_c_155_n N_VPWR_c_405_n 0.0119993f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A_c_156_n N_VPWR_c_405_n 0.0119993f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_c_157_n N_VPWR_c_405_n 6.03055e-19 $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_c_156_n N_VPWR_c_406_n 6.03055e-19 $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A_c_157_n N_VPWR_c_406_n 0.0119993f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_c_158_n N_VPWR_c_406_n 0.0119993f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_c_159_n N_VPWR_c_406_n 6.03055e-19 $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_c_158_n N_VPWR_c_407_n 6.03055e-19 $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A_c_159_n N_VPWR_c_407_n 0.0129761f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_c_154_n N_VPWR_c_408_n 0.00622633f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_c_155_n N_VPWR_c_408_n 0.00622633f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_c_156_n N_VPWR_c_410_n 0.00622633f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A_c_157_n N_VPWR_c_410_n 0.00622633f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A_c_158_n N_VPWR_c_412_n 0.00622633f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A_c_159_n N_VPWR_c_412_n 0.00622633f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_c_142_n N_VPWR_c_414_n 0.00622633f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_c_143_n N_VPWR_c_414_n 0.00622633f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_c_144_n N_VPWR_c_415_n 0.00622633f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A_c_145_n N_VPWR_c_415_n 0.00622633f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A_c_142_n N_VPWR_c_392_n 0.0104011f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A_c_143_n N_VPWR_c_392_n 0.0104011f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A_c_144_n N_VPWR_c_392_n 0.0104011f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_186 N_A_c_145_n N_VPWR_c_392_n 0.0104011f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_187 N_A_c_146_n N_VPWR_c_392_n 0.0104011f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A_c_147_n N_VPWR_c_392_n 0.0104011f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A_c_148_n N_VPWR_c_392_n 0.0104011f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_190 N_A_c_149_n N_VPWR_c_392_n 0.0104011f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_191 N_A_c_150_n N_VPWR_c_392_n 0.0104011f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_192 N_A_c_151_n N_VPWR_c_392_n 0.0104011f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A_c_152_n N_VPWR_c_392_n 0.0104011f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A_c_153_n N_VPWR_c_392_n 0.0104011f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A_c_154_n N_VPWR_c_392_n 0.0104011f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A_c_155_n N_VPWR_c_392_n 0.0104011f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A_c_156_n N_VPWR_c_392_n 0.0104011f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_c_157_n N_VPWR_c_392_n 0.0104011f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A_c_158_n N_VPWR_c_392_n 0.0104011f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_200 N_A_c_159_n N_VPWR_c_392_n 0.0104011f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A_c_142_n N_Y_c_545_n 0.00180824f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A_c_234_p N_Y_c_545_n 0.0202172f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A_c_141_n N_Y_c_545_n 0.0137702f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_204 N_A_M1002_g N_Y_c_546_n 0.0121037f $X=1.93 $Y=0.445 $X2=0 $Y2=0
cc_205 N_A_c_234_p N_Y_c_546_n 0.113639f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A_c_141_n N_Y_c_546_n 0.0370545f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_207 N_A_c_142_n N_Y_c_568_n 0.0167971f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A_c_234_p N_Y_c_568_n 0.00979398f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A_c_141_n N_Y_c_568_n 5.92681e-19 $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_210 N_A_c_143_n N_Y_c_570_n 0.0149843f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A_c_144_n N_Y_c_570_n 0.0149843f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A_c_234_p N_Y_c_570_n 0.0479566f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A_c_141_n N_Y_c_570_n 0.00738631f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_214 N_A_c_145_n N_Y_c_571_n 0.0149843f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A_c_146_n N_Y_c_571_n 0.0149843f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A_c_234_p N_Y_c_571_n 0.0479566f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A_c_141_n N_Y_c_571_n 0.00822052f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_218 N_A_M1002_g N_Y_c_548_n 0.00113469f $X=1.93 $Y=0.445 $X2=0 $Y2=0
cc_219 N_A_M1006_g N_Y_c_548_n 6.66199e-19 $X=2.35 $Y=0.445 $X2=0 $Y2=0
cc_220 N_A_M1006_g N_Y_c_549_n 0.0105559f $X=2.35 $Y=0.445 $X2=0 $Y2=0
cc_221 N_A_M1009_g N_Y_c_549_n 0.0105559f $X=2.87 $Y=0.445 $X2=0 $Y2=0
cc_222 N_A_c_234_p N_Y_c_549_n 0.0481922f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A_c_141_n N_Y_c_549_n 0.00446519f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_224 N_A_c_147_n N_Y_c_572_n 0.0149843f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A_c_148_n N_Y_c_572_n 0.0149843f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_226 N_A_c_234_p N_Y_c_572_n 0.0479566f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A_c_141_n N_Y_c_572_n 0.00825306f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_228 N_A_M1009_g N_Y_c_550_n 6.66199e-19 $X=2.87 $Y=0.445 $X2=0 $Y2=0
cc_229 N_A_M1010_g N_Y_c_550_n 6.66199e-19 $X=3.29 $Y=0.445 $X2=0 $Y2=0
cc_230 N_A_M1010_g N_Y_c_551_n 0.0105559f $X=3.29 $Y=0.445 $X2=0 $Y2=0
cc_231 N_A_M1013_g N_Y_c_551_n 0.0105559f $X=3.81 $Y=0.445 $X2=0 $Y2=0
cc_232 N_A_c_234_p N_Y_c_551_n 0.0481922f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_233 N_A_c_141_n N_Y_c_551_n 0.00446519f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_234 N_A_c_149_n N_Y_c_573_n 0.0149843f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A_c_150_n N_Y_c_573_n 0.0149843f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A_c_234_p N_Y_c_573_n 0.0479566f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A_c_141_n N_Y_c_573_n 0.00825306f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_238 N_A_M1013_g N_Y_c_552_n 6.66199e-19 $X=3.81 $Y=0.445 $X2=0 $Y2=0
cc_239 N_A_M1014_g N_Y_c_552_n 6.66199e-19 $X=4.23 $Y=0.445 $X2=0 $Y2=0
cc_240 N_A_M1014_g N_Y_c_553_n 0.0105559f $X=4.23 $Y=0.445 $X2=0 $Y2=0
cc_241 N_A_M1017_g N_Y_c_553_n 0.0105559f $X=4.75 $Y=0.445 $X2=0 $Y2=0
cc_242 N_A_c_234_p N_Y_c_553_n 0.0481922f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_243 N_A_c_141_n N_Y_c_553_n 0.00446519f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_244 N_A_c_151_n N_Y_c_574_n 0.0149843f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_245 N_A_c_152_n N_Y_c_574_n 0.0149843f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_246 N_A_c_234_p N_Y_c_574_n 0.0479566f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_247 N_A_c_141_n N_Y_c_574_n 0.00825306f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_248 N_A_M1017_g N_Y_c_554_n 6.66199e-19 $X=4.75 $Y=0.445 $X2=0 $Y2=0
cc_249 N_A_M1020_g N_Y_c_554_n 6.66199e-19 $X=5.17 $Y=0.445 $X2=0 $Y2=0
cc_250 N_A_M1020_g N_Y_c_555_n 0.0105559f $X=5.17 $Y=0.445 $X2=0 $Y2=0
cc_251 N_A_M1024_g N_Y_c_555_n 0.0105559f $X=5.69 $Y=0.445 $X2=0 $Y2=0
cc_252 N_A_c_234_p N_Y_c_555_n 0.0481922f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_253 N_A_c_141_n N_Y_c_555_n 0.00446519f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_254 N_A_c_153_n N_Y_c_575_n 0.0149843f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_255 N_A_c_154_n N_Y_c_575_n 0.0149843f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_256 N_A_c_234_p N_Y_c_575_n 0.0479566f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_257 N_A_c_141_n N_Y_c_575_n 0.00825306f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_258 N_A_M1024_g N_Y_c_556_n 6.66199e-19 $X=5.69 $Y=0.445 $X2=0 $Y2=0
cc_259 N_A_M1026_g N_Y_c_556_n 6.66199e-19 $X=6.11 $Y=0.445 $X2=0 $Y2=0
cc_260 N_A_M1026_g N_Y_c_557_n 0.0105559f $X=6.11 $Y=0.445 $X2=0 $Y2=0
cc_261 N_A_M1027_g N_Y_c_557_n 0.0105559f $X=6.63 $Y=0.445 $X2=0 $Y2=0
cc_262 N_A_c_234_p N_Y_c_557_n 0.0481922f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_263 N_A_c_141_n N_Y_c_557_n 0.00446519f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_264 N_A_c_155_n N_Y_c_576_n 0.0149843f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A_c_156_n N_Y_c_576_n 0.0149843f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A_c_234_p N_Y_c_576_n 0.0479566f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_267 N_A_c_141_n N_Y_c_576_n 0.00822052f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_268 N_A_M1027_g N_Y_c_558_n 6.66199e-19 $X=6.63 $Y=0.445 $X2=0 $Y2=0
cc_269 N_A_M1028_g N_Y_c_558_n 0.00113469f $X=7.05 $Y=0.445 $X2=0 $Y2=0
cc_270 N_A_M1028_g N_Y_c_559_n 0.0121037f $X=7.05 $Y=0.445 $X2=0 $Y2=0
cc_271 N_A_c_234_p N_Y_c_559_n 0.0694192f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_272 N_A_c_141_n N_Y_c_559_n 0.0253858f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_273 N_A_c_157_n N_Y_c_577_n 0.0149843f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_274 N_A_c_158_n N_Y_c_577_n 0.0161446f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_275 N_A_c_234_p N_Y_c_577_n 0.0346647f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_276 N_A_c_141_n N_Y_c_577_n 0.0071181f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_277 N_A_c_234_p N_Y_c_578_n 0.0223745f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_278 N_A_c_141_n N_Y_c_578_n 0.00656124f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_279 N_A_c_234_p N_Y_c_579_n 0.0223745f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_280 N_A_c_141_n N_Y_c_579_n 0.00656124f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_281 N_A_M1002_g N_Y_c_560_n 0.00196728f $X=1.93 $Y=0.445 $X2=0 $Y2=0
cc_282 N_A_M1006_g N_Y_c_560_n 0.00196728f $X=2.35 $Y=0.445 $X2=0 $Y2=0
cc_283 N_A_c_234_p N_Y_c_560_n 0.0221763f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_284 N_A_c_141_n N_Y_c_560_n 0.00218937f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_285 N_A_c_234_p N_Y_c_580_n 0.0223745f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_286 N_A_c_141_n N_Y_c_580_n 0.00688898f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_287 N_A_M1009_g N_Y_c_561_n 0.00196728f $X=2.87 $Y=0.445 $X2=0 $Y2=0
cc_288 N_A_M1010_g N_Y_c_561_n 0.00196728f $X=3.29 $Y=0.445 $X2=0 $Y2=0
cc_289 N_A_c_234_p N_Y_c_561_n 0.0221763f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_290 N_A_c_141_n N_Y_c_561_n 0.00218937f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_291 N_A_c_234_p N_Y_c_581_n 0.0223745f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_292 N_A_c_141_n N_Y_c_581_n 0.00688898f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_293 N_A_M1013_g N_Y_c_562_n 0.00196728f $X=3.81 $Y=0.445 $X2=0 $Y2=0
cc_294 N_A_M1014_g N_Y_c_562_n 0.00196728f $X=4.23 $Y=0.445 $X2=0 $Y2=0
cc_295 N_A_c_234_p N_Y_c_562_n 0.0221763f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_296 N_A_c_141_n N_Y_c_562_n 0.00218937f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_297 N_A_c_234_p N_Y_c_582_n 0.0223745f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_298 N_A_c_141_n N_Y_c_582_n 0.00688898f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_299 N_A_M1017_g N_Y_c_563_n 0.00196728f $X=4.75 $Y=0.445 $X2=0 $Y2=0
cc_300 N_A_M1020_g N_Y_c_563_n 0.00196728f $X=5.17 $Y=0.445 $X2=0 $Y2=0
cc_301 N_A_c_234_p N_Y_c_563_n 0.0221763f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_302 N_A_c_141_n N_Y_c_563_n 0.00218937f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_303 N_A_c_234_p N_Y_c_583_n 0.0223745f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_304 N_A_c_141_n N_Y_c_583_n 0.00688898f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_305 N_A_M1024_g N_Y_c_564_n 0.00196728f $X=5.69 $Y=0.445 $X2=0 $Y2=0
cc_306 N_A_M1026_g N_Y_c_564_n 0.00196728f $X=6.11 $Y=0.445 $X2=0 $Y2=0
cc_307 N_A_c_234_p N_Y_c_564_n 0.0221763f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_308 N_A_c_141_n N_Y_c_564_n 0.00218937f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_309 N_A_c_234_p N_Y_c_584_n 0.0223745f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_310 N_A_c_141_n N_Y_c_584_n 0.00688898f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_311 N_A_M1027_g N_Y_c_565_n 0.00196728f $X=6.63 $Y=0.445 $X2=0 $Y2=0
cc_312 N_A_M1028_g N_Y_c_565_n 0.00196728f $X=7.05 $Y=0.445 $X2=0 $Y2=0
cc_313 N_A_c_234_p N_Y_c_565_n 0.0221763f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_314 N_A_c_141_n N_Y_c_565_n 0.00218937f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_315 N_A_c_234_p N_Y_c_585_n 0.0223745f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_316 N_A_c_141_n N_Y_c_585_n 0.00656124f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_317 N_A_c_158_n N_Y_c_586_n 3.55576e-19 $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_318 N_A_c_159_n N_Y_c_586_n 0.0144247f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_319 N_A_c_157_n Y 2.17606e-19 $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_320 N_A_c_158_n Y 0.00145782f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_321 N_A_c_159_n Y 0.00215997f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_322 N_A_c_234_p Y 0.0204994f $X=7.76 $Y=1.16 $X2=0 $Y2=0
cc_323 N_A_c_141_n Y 0.0515261f $X=8.015 $Y=1.202 $X2=0 $Y2=0
cc_324 N_A_M1006_g N_VGND_c_808_n 0.00175491f $X=2.35 $Y=0.445 $X2=0 $Y2=0
cc_325 N_A_M1009_g N_VGND_c_808_n 0.00175624f $X=2.87 $Y=0.445 $X2=0 $Y2=0
cc_326 N_A_M1009_g N_VGND_c_809_n 0.00433717f $X=2.87 $Y=0.445 $X2=0 $Y2=0
cc_327 N_A_M1010_g N_VGND_c_809_n 0.00433717f $X=3.29 $Y=0.445 $X2=0 $Y2=0
cc_328 N_A_M1010_g N_VGND_c_810_n 0.00175624f $X=3.29 $Y=0.445 $X2=0 $Y2=0
cc_329 N_A_M1013_g N_VGND_c_810_n 0.00175624f $X=3.81 $Y=0.445 $X2=0 $Y2=0
cc_330 N_A_M1013_g N_VGND_c_811_n 0.00433717f $X=3.81 $Y=0.445 $X2=0 $Y2=0
cc_331 N_A_M1014_g N_VGND_c_811_n 0.00433717f $X=4.23 $Y=0.445 $X2=0 $Y2=0
cc_332 N_A_M1014_g N_VGND_c_812_n 0.00175624f $X=4.23 $Y=0.445 $X2=0 $Y2=0
cc_333 N_A_M1017_g N_VGND_c_812_n 0.00175624f $X=4.75 $Y=0.445 $X2=0 $Y2=0
cc_334 N_A_M1017_g N_VGND_c_813_n 0.00433717f $X=4.75 $Y=0.445 $X2=0 $Y2=0
cc_335 N_A_M1020_g N_VGND_c_813_n 0.00433717f $X=5.17 $Y=0.445 $X2=0 $Y2=0
cc_336 N_A_M1020_g N_VGND_c_814_n 0.00175624f $X=5.17 $Y=0.445 $X2=0 $Y2=0
cc_337 N_A_M1024_g N_VGND_c_814_n 0.00175624f $X=5.69 $Y=0.445 $X2=0 $Y2=0
cc_338 N_A_M1024_g N_VGND_c_815_n 0.00433717f $X=5.69 $Y=0.445 $X2=0 $Y2=0
cc_339 N_A_M1026_g N_VGND_c_815_n 0.00433717f $X=6.11 $Y=0.445 $X2=0 $Y2=0
cc_340 N_A_M1026_g N_VGND_c_816_n 0.00175624f $X=6.11 $Y=0.445 $X2=0 $Y2=0
cc_341 N_A_M1027_g N_VGND_c_816_n 0.00175491f $X=6.63 $Y=0.445 $X2=0 $Y2=0
cc_342 N_A_M1002_g N_VGND_c_817_n 0.00433717f $X=1.93 $Y=0.445 $X2=0 $Y2=0
cc_343 N_A_M1006_g N_VGND_c_817_n 0.00433717f $X=2.35 $Y=0.445 $X2=0 $Y2=0
cc_344 N_A_M1002_g N_VGND_c_819_n 0.00710548f $X=1.93 $Y=0.445 $X2=0 $Y2=0
cc_345 N_A_M1006_g N_VGND_c_819_n 0.00602419f $X=2.35 $Y=0.445 $X2=0 $Y2=0
cc_346 N_A_M1009_g N_VGND_c_819_n 0.00602419f $X=2.87 $Y=0.445 $X2=0 $Y2=0
cc_347 N_A_M1010_g N_VGND_c_819_n 0.00602419f $X=3.29 $Y=0.445 $X2=0 $Y2=0
cc_348 N_A_M1013_g N_VGND_c_819_n 0.00602419f $X=3.81 $Y=0.445 $X2=0 $Y2=0
cc_349 N_A_M1014_g N_VGND_c_819_n 0.00602419f $X=4.23 $Y=0.445 $X2=0 $Y2=0
cc_350 N_A_M1017_g N_VGND_c_819_n 0.00602419f $X=4.75 $Y=0.445 $X2=0 $Y2=0
cc_351 N_A_M1020_g N_VGND_c_819_n 0.00602419f $X=5.17 $Y=0.445 $X2=0 $Y2=0
cc_352 N_A_M1024_g N_VGND_c_819_n 0.00602419f $X=5.69 $Y=0.445 $X2=0 $Y2=0
cc_353 N_A_M1026_g N_VGND_c_819_n 0.00602419f $X=6.11 $Y=0.445 $X2=0 $Y2=0
cc_354 N_A_M1027_g N_VGND_c_819_n 0.00602419f $X=6.63 $Y=0.445 $X2=0 $Y2=0
cc_355 N_A_M1028_g N_VGND_c_819_n 0.00710548f $X=7.05 $Y=0.445 $X2=0 $Y2=0
cc_356 N_A_M1002_g N_VGND_c_821_n 0.00348282f $X=1.93 $Y=0.445 $X2=0 $Y2=0
cc_357 N_A_M1027_g N_VGND_c_827_n 0.00433717f $X=6.63 $Y=0.445 $X2=0 $Y2=0
cc_358 N_A_M1028_g N_VGND_c_827_n 0.00433717f $X=7.05 $Y=0.445 $X2=0 $Y2=0
cc_359 N_A_M1028_g N_VGND_c_828_n 0.00348282f $X=7.05 $Y=0.445 $X2=0 $Y2=0
cc_360 N_VPWR_c_392_n N_Y_M1000_s 0.00300692f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_361 N_VPWR_c_392_n N_Y_M1003_s 0.00300692f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_362 N_VPWR_c_392_n N_Y_M1005_s 0.00300692f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_363 N_VPWR_c_392_n N_Y_M1008_s 0.00300692f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_364 N_VPWR_c_392_n N_Y_M1012_s 0.00300692f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_365 N_VPWR_c_392_n N_Y_M1016_s 0.00300692f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_366 N_VPWR_c_392_n N_Y_M1019_s 0.00300692f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_367 N_VPWR_c_392_n N_Y_M1022_s 0.00300692f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_368 N_VPWR_c_392_n N_Y_M1025_s 0.00300692f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_369 N_VPWR_M1000_d N_Y_c_568_n 6.59072e-19 $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_370 N_VPWR_c_394_n N_Y_c_568_n 0.00649432f $X=0.26 $Y=1.925 $X2=0 $Y2=0
cc_371 N_VPWR_M1000_d N_Y_c_569_n 0.00238226f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_372 N_VPWR_c_394_n N_Y_c_569_n 0.0153514f $X=0.26 $Y=1.925 $X2=0 $Y2=0
cc_373 N_VPWR_c_414_n N_Y_c_724_n 0.0156407f $X=1.035 $Y=2.72 $X2=0 $Y2=0
cc_374 N_VPWR_c_392_n N_Y_c_724_n 0.0103212f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_375 N_VPWR_M1001_d N_Y_c_570_n 0.00187091f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_376 N_VPWR_c_395_n N_Y_c_570_n 0.0171295f $X=1.2 $Y=1.925 $X2=0 $Y2=0
cc_377 N_VPWR_c_415_n N_Y_c_728_n 0.0156407f $X=1.975 $Y=2.72 $X2=0 $Y2=0
cc_378 N_VPWR_c_392_n N_Y_c_728_n 0.0103212f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_379 N_VPWR_M1004_d N_Y_c_571_n 0.00187091f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_380 N_VPWR_c_396_n N_Y_c_571_n 0.0171295f $X=2.14 $Y=1.925 $X2=0 $Y2=0
cc_381 N_VPWR_c_397_n N_Y_c_732_n 0.0156407f $X=2.915 $Y=2.72 $X2=0 $Y2=0
cc_382 N_VPWR_c_392_n N_Y_c_732_n 0.0103212f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_383 N_VPWR_M1007_d N_Y_c_572_n 0.00187091f $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_384 N_VPWR_c_398_n N_Y_c_572_n 0.0171295f $X=3.08 $Y=1.925 $X2=0 $Y2=0
cc_385 N_VPWR_c_399_n N_Y_c_736_n 0.0156407f $X=3.855 $Y=2.72 $X2=0 $Y2=0
cc_386 N_VPWR_c_392_n N_Y_c_736_n 0.0103212f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_387 N_VPWR_M1011_d N_Y_c_573_n 0.00187091f $X=3.875 $Y=1.485 $X2=0 $Y2=0
cc_388 N_VPWR_c_400_n N_Y_c_573_n 0.0171295f $X=4.02 $Y=1.925 $X2=0 $Y2=0
cc_389 N_VPWR_c_401_n N_Y_c_740_n 0.0156407f $X=4.795 $Y=2.72 $X2=0 $Y2=0
cc_390 N_VPWR_c_392_n N_Y_c_740_n 0.0103212f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_391 N_VPWR_M1015_d N_Y_c_574_n 0.00187091f $X=4.815 $Y=1.485 $X2=0 $Y2=0
cc_392 N_VPWR_c_402_n N_Y_c_574_n 0.0171295f $X=4.96 $Y=1.925 $X2=0 $Y2=0
cc_393 N_VPWR_c_403_n N_Y_c_744_n 0.0156407f $X=5.735 $Y=2.72 $X2=0 $Y2=0
cc_394 N_VPWR_c_392_n N_Y_c_744_n 0.0103212f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_395 N_VPWR_M1018_d N_Y_c_575_n 0.00187091f $X=5.755 $Y=1.485 $X2=0 $Y2=0
cc_396 N_VPWR_c_404_n N_Y_c_575_n 0.0171295f $X=5.9 $Y=1.925 $X2=0 $Y2=0
cc_397 N_VPWR_c_408_n N_Y_c_748_n 0.0156407f $X=6.675 $Y=2.72 $X2=0 $Y2=0
cc_398 N_VPWR_c_392_n N_Y_c_748_n 0.0103212f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_399 N_VPWR_M1021_d N_Y_c_576_n 0.00187091f $X=6.695 $Y=1.485 $X2=0 $Y2=0
cc_400 N_VPWR_c_405_n N_Y_c_576_n 0.0171295f $X=6.84 $Y=1.925 $X2=0 $Y2=0
cc_401 N_VPWR_c_410_n N_Y_c_752_n 0.0156407f $X=7.615 $Y=2.72 $X2=0 $Y2=0
cc_402 N_VPWR_c_392_n N_Y_c_752_n 0.0103212f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_403 N_VPWR_M1023_d N_Y_c_577_n 0.00187091f $X=7.635 $Y=1.485 $X2=0 $Y2=0
cc_404 N_VPWR_c_406_n N_Y_c_577_n 0.0171295f $X=7.78 $Y=1.925 $X2=0 $Y2=0
cc_405 N_VPWR_c_412_n N_Y_c_756_n 0.0156407f $X=8.555 $Y=2.72 $X2=0 $Y2=0
cc_406 N_VPWR_c_392_n N_Y_c_756_n 0.0103212f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_407 N_VPWR_M1029_d N_Y_c_586_n 0.00679555f $X=8.575 $Y=1.485 $X2=0 $Y2=0
cc_408 N_VPWR_c_407_n N_Y_c_586_n 0.00363976f $X=8.72 $Y=1.925 $X2=0 $Y2=0
cc_409 N_Y_c_549_n N_VGND_c_808_n 0.0226915f $X=2.945 $Y=0.78 $X2=0 $Y2=0
cc_410 N_Y_c_549_n N_VGND_c_809_n 0.00245234f $X=2.945 $Y=0.78 $X2=0 $Y2=0
cc_411 N_Y_c_550_n N_VGND_c_809_n 0.0148571f $X=3.08 $Y=0.445 $X2=0 $Y2=0
cc_412 N_Y_c_551_n N_VGND_c_809_n 0.00245234f $X=3.885 $Y=0.78 $X2=0 $Y2=0
cc_413 N_Y_c_551_n N_VGND_c_810_n 0.0226915f $X=3.885 $Y=0.78 $X2=0 $Y2=0
cc_414 N_Y_c_551_n N_VGND_c_811_n 0.00245234f $X=3.885 $Y=0.78 $X2=0 $Y2=0
cc_415 N_Y_c_552_n N_VGND_c_811_n 0.0148571f $X=4.02 $Y=0.445 $X2=0 $Y2=0
cc_416 N_Y_c_553_n N_VGND_c_811_n 0.00245234f $X=4.825 $Y=0.78 $X2=0 $Y2=0
cc_417 N_Y_c_553_n N_VGND_c_812_n 0.0226915f $X=4.825 $Y=0.78 $X2=0 $Y2=0
cc_418 N_Y_c_553_n N_VGND_c_813_n 0.00245234f $X=4.825 $Y=0.78 $X2=0 $Y2=0
cc_419 N_Y_c_554_n N_VGND_c_813_n 0.0148571f $X=4.96 $Y=0.445 $X2=0 $Y2=0
cc_420 N_Y_c_555_n N_VGND_c_813_n 0.00245234f $X=5.765 $Y=0.78 $X2=0 $Y2=0
cc_421 N_Y_c_555_n N_VGND_c_814_n 0.0226915f $X=5.765 $Y=0.78 $X2=0 $Y2=0
cc_422 N_Y_c_555_n N_VGND_c_815_n 0.00245234f $X=5.765 $Y=0.78 $X2=0 $Y2=0
cc_423 N_Y_c_556_n N_VGND_c_815_n 0.0148571f $X=5.9 $Y=0.445 $X2=0 $Y2=0
cc_424 N_Y_c_557_n N_VGND_c_815_n 0.00245234f $X=6.705 $Y=0.78 $X2=0 $Y2=0
cc_425 N_Y_c_557_n N_VGND_c_816_n 0.0226915f $X=6.705 $Y=0.78 $X2=0 $Y2=0
cc_426 N_Y_c_546_n N_VGND_c_817_n 0.00245234f $X=2.005 $Y=0.78 $X2=0 $Y2=0
cc_427 N_Y_c_548_n N_VGND_c_817_n 0.0148571f $X=2.14 $Y=0.445 $X2=0 $Y2=0
cc_428 N_Y_c_549_n N_VGND_c_817_n 0.00245234f $X=2.945 $Y=0.78 $X2=0 $Y2=0
cc_429 N_Y_c_559_n N_VGND_c_818_n 0.0145882f $X=8.1 $Y=0.78 $X2=0 $Y2=0
cc_430 N_Y_M1002_d N_VGND_c_819_n 0.00215201f $X=2.005 $Y=0.235 $X2=0 $Y2=0
cc_431 N_Y_M1009_d N_VGND_c_819_n 0.00215201f $X=2.945 $Y=0.235 $X2=0 $Y2=0
cc_432 N_Y_M1013_d N_VGND_c_819_n 0.00215201f $X=3.885 $Y=0.235 $X2=0 $Y2=0
cc_433 N_Y_M1017_d N_VGND_c_819_n 0.00215201f $X=4.825 $Y=0.235 $X2=0 $Y2=0
cc_434 N_Y_M1024_d N_VGND_c_819_n 0.00215201f $X=5.765 $Y=0.235 $X2=0 $Y2=0
cc_435 N_Y_M1027_d N_VGND_c_819_n 0.00215201f $X=6.705 $Y=0.235 $X2=0 $Y2=0
cc_436 N_Y_c_546_n N_VGND_c_819_n 0.0302627f $X=2.005 $Y=0.78 $X2=0 $Y2=0
cc_437 N_Y_c_547_n N_VGND_c_819_n 0.00489372f $X=0.285 $Y=0.78 $X2=0 $Y2=0
cc_438 N_Y_c_548_n N_VGND_c_819_n 0.0102919f $X=2.14 $Y=0.445 $X2=0 $Y2=0
cc_439 N_Y_c_549_n N_VGND_c_819_n 0.00891516f $X=2.945 $Y=0.78 $X2=0 $Y2=0
cc_440 N_Y_c_550_n N_VGND_c_819_n 0.0102919f $X=3.08 $Y=0.445 $X2=0 $Y2=0
cc_441 N_Y_c_551_n N_VGND_c_819_n 0.00891516f $X=3.885 $Y=0.78 $X2=0 $Y2=0
cc_442 N_Y_c_552_n N_VGND_c_819_n 0.0102919f $X=4.02 $Y=0.445 $X2=0 $Y2=0
cc_443 N_Y_c_553_n N_VGND_c_819_n 0.00891516f $X=4.825 $Y=0.78 $X2=0 $Y2=0
cc_444 N_Y_c_554_n N_VGND_c_819_n 0.0102919f $X=4.96 $Y=0.445 $X2=0 $Y2=0
cc_445 N_Y_c_555_n N_VGND_c_819_n 0.00891516f $X=5.765 $Y=0.78 $X2=0 $Y2=0
cc_446 N_Y_c_556_n N_VGND_c_819_n 0.0102919f $X=5.9 $Y=0.445 $X2=0 $Y2=0
cc_447 N_Y_c_557_n N_VGND_c_819_n 0.00891516f $X=6.705 $Y=0.78 $X2=0 $Y2=0
cc_448 N_Y_c_558_n N_VGND_c_819_n 0.0102919f $X=6.84 $Y=0.445 $X2=0 $Y2=0
cc_449 N_Y_c_559_n N_VGND_c_819_n 0.030148f $X=8.1 $Y=0.78 $X2=0 $Y2=0
cc_450 N_Y_c_546_n N_VGND_c_820_n 0.0142044f $X=2.005 $Y=0.78 $X2=0 $Y2=0
cc_451 N_Y_c_547_n N_VGND_c_820_n 0.0030627f $X=0.285 $Y=0.78 $X2=0 $Y2=0
cc_452 N_Y_c_546_n N_VGND_c_821_n 0.051019f $X=2.005 $Y=0.78 $X2=0 $Y2=0
cc_453 N_Y_c_557_n N_VGND_c_827_n 0.00245234f $X=6.705 $Y=0.78 $X2=0 $Y2=0
cc_454 N_Y_c_558_n N_VGND_c_827_n 0.0148571f $X=6.84 $Y=0.445 $X2=0 $Y2=0
cc_455 N_Y_c_559_n N_VGND_c_827_n 0.00245234f $X=8.1 $Y=0.78 $X2=0 $Y2=0
cc_456 N_Y_c_559_n N_VGND_c_828_n 0.051019f $X=8.1 $Y=0.78 $X2=0 $Y2=0
