* File: sky130_fd_sc_hdll__and4_4.spice
* Created: Thu Aug 27 18:58:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and4_4.pex.spice"
.subckt sky130_fd_sc_hdll__and4_4  VNB VPB A B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1012 A_119_47# N_A_M1012_g N_A_27_47#_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.079625 AS=0.2015 PD=0.895 PS=1.92 NRD=12.456 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1001 A_198_47# N_B_M1001_g A_119_47# VNB NSHORT L=0.15 W=0.65 AD=0.1235
+ AS=0.079625 PD=1.03 PS=0.895 NRD=24.912 NRS=12.456 M=1 R=4.33333 SA=75000.6
+ SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1015 A_304_47# N_C_M1015_g A_198_47# VNB NSHORT L=0.15 W=0.65 AD=0.157625
+ AS=0.1235 PD=1.135 PS=1.03 NRD=34.608 NRS=24.912 M=1 R=4.33333 SA=75001.2
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_D_M1005_g A_304_47# VNB NSHORT L=0.15 W=0.65 AD=0.1235
+ AS=0.157625 PD=1.03 PS=1.135 NRD=17.532 NRS=34.608 M=1 R=4.33333 SA=75001.8
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1005_d N_A_27_47#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.104 PD=1.03 PS=0.97 NRD=0.912 NRS=8.304 M=1 R=4.33333
+ SA=75002.3 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A_27_47#_M1008_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.8
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1008_d N_A_27_47#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.3
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_A_27_47#_M1013_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_A_27_47#_M1006_d N_A_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.7 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_B_M1002_g N_A_27_47#_M1006_d VPB PHIGHVT L=0.18 W=1
+ AD=0.165 AS=0.145 PD=1.33 PS=1.29 NRD=4.9053 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003.3 A=0.18 P=2.36 MULT=1
MM1003 N_A_27_47#_M1003_d N_C_M1003_g N_VPWR_M1002_d VPB PHIGHVT L=0.18 W=1
+ AD=0.225 AS=0.165 PD=1.45 PS=1.33 NRD=0.9653 NRS=4.9053 M=1 R=5.55556
+ SA=90001.2 SB=90002.7 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_D_M1000_g N_A_27_47#_M1003_d VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.225 PD=1.35 PS=1.45 NRD=10.8153 NRS=32.4853 M=1 R=5.55556
+ SA=90001.8 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1000_d N_A_27_47#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.145 PD=1.35 PS=1.29 NRD=2.9353 NRS=0.9653 M=1 R=5.55556
+ SA=90002.3 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1010_d N_A_27_47#_M1010_g N_X_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.8 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1010_d N_A_27_47#_M1011_g N_X_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.3 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1014 N_VPWR_M1014_d N_A_27_47#_M1014_g N_X_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.7 SB=90000.2 A=0.18 P=2.36 MULT=1
DX16_noxref VNB VPB NWDIODE A=7.9929 P=13.17
*
.include "sky130_fd_sc_hdll__and4_4.pxi.spice"
*
.ends
*
*
