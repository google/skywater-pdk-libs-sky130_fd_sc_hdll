* File: sky130_fd_sc_hdll__ebufn_8.pex.spice
* Created: Thu Aug 27 19:07:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__EBUFN_8%A 1 3 4 6 7 9 12 14 15 23
c44 23 0 1.55488e-19 $X=1 $Y=1.202
c45 12 0 1.13485e-20 $X=1.025 $Y=0.56
c46 7 0 1.41448e-19 $X=1 $Y=1.41
r47 23 24 3.52339 $w=3.42e-07 $l=2.5e-08 $layer=POLY_cond $X=1 $Y=1.202
+ $X2=1.025 $Y2=1.202
r48 22 23 62.7164 $w=3.42e-07 $l=4.45e-07 $layer=POLY_cond $X=0.555 $Y=1.202
+ $X2=1 $Y2=1.202
r49 21 22 3.52339 $w=3.42e-07 $l=2.5e-08 $layer=POLY_cond $X=0.53 $Y=1.202
+ $X2=0.555 $Y2=1.202
r50 19 21 33.1199 $w=3.42e-07 $l=2.35e-07 $layer=POLY_cond $X=0.295 $Y=1.202
+ $X2=0.53 $Y2=1.202
r51 14 15 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.257 $Y=1.16
+ $X2=0.257 $Y2=1.53
r52 14 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.295
+ $Y=1.16 $X2=0.295 $Y2=1.16
r53 10 24 22.0749 $w=1.5e-07 $l=1.77e-07 $layer=POLY_cond $X=1.025 $Y=1.025
+ $X2=1.025 $Y2=1.202
r54 10 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.025 $Y=1.025
+ $X2=1.025 $Y2=0.56
r55 7 23 17.7656 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1 $Y=1.41 $X2=1
+ $Y2=1.202
r56 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1 $Y=1.41 $X2=1
+ $Y2=1.985
r57 4 22 22.0749 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.555 $Y=0.995
+ $X2=0.555 $Y2=1.202
r58 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.555 $Y=0.995
+ $X2=0.555 $Y2=0.56
r59 1 21 17.7656 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.53 $Y=1.41
+ $X2=0.53 $Y2=1.202
r60 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.53 $Y=1.41 $X2=0.53
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_8%TE_B 1 3 4 6 8 9 11 13 14 16 18 19 21 23
+ 24 26 28 29 31 33 34 36 38 39 41 43 44 46 48 49 50 51 52 53 54 55 56 57 58 59
c174 39 0 7.91225e-20 $X=5.575 $Y=1.395
c175 29 0 7.91225e-20 $X=4.535 $Y=1.395
c176 19 0 7.91225e-20 $X=3.495 $Y=1.395
r177 65 66 3.17942 $w=3.79e-07 $l=2.5e-08 $layer=POLY_cond $X=1.53 $Y=1.202
+ $X2=1.555 $Y2=1.202
r178 63 65 10.81 $w=3.79e-07 $l=8.5e-08 $layer=POLY_cond $X=1.445 $Y=1.202
+ $X2=1.53 $Y2=1.202
r179 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.445
+ $Y=1.16 $X2=1.445 $Y2=1.16
r180 59 64 10.6714 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.275 $Y=1.53
+ $X2=1.275 $Y2=1.16
r181 58 64 8.9409 $w=4.23e-07 $l=3.1e-07 $layer=LI1_cond $X=1.275 $Y=0.85
+ $X2=1.275 $Y2=1.16
r182 49 50 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.07 $Y=1.232
+ $X2=2.22 $Y2=1.232
r183 46 48 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=6.185 $Y=1.47
+ $X2=6.185 $Y2=2.015
r184 45 57 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.755 $Y=1.395
+ $X2=5.665 $Y2=1.395
r185 44 46 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.095 $Y=1.395
+ $X2=6.185 $Y2=1.47
r186 44 45 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=6.095 $Y=1.395
+ $X2=5.755 $Y2=1.395
r187 41 57 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.665 $Y=1.47
+ $X2=5.665 $Y2=1.395
r188 41 43 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=5.665 $Y=1.47
+ $X2=5.665 $Y2=2.015
r189 40 56 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.235 $Y=1.395
+ $X2=5.145 $Y2=1.395
r190 39 57 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.575 $Y=1.395
+ $X2=5.665 $Y2=1.395
r191 39 40 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=5.575 $Y=1.395
+ $X2=5.235 $Y2=1.395
r192 36 56 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.145 $Y=1.47
+ $X2=5.145 $Y2=1.395
r193 36 38 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=5.145 $Y=1.47
+ $X2=5.145 $Y2=2.015
r194 35 55 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.715 $Y=1.395
+ $X2=4.625 $Y2=1.395
r195 34 56 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.055 $Y=1.395
+ $X2=5.145 $Y2=1.395
r196 34 35 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=5.055 $Y=1.395
+ $X2=4.715 $Y2=1.395
r197 31 55 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.625 $Y=1.47
+ $X2=4.625 $Y2=1.395
r198 31 33 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=4.625 $Y=1.47
+ $X2=4.625 $Y2=2.015
r199 30 54 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.195 $Y=1.395
+ $X2=4.105 $Y2=1.395
r200 29 55 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.535 $Y=1.395
+ $X2=4.625 $Y2=1.395
r201 29 30 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=4.535 $Y=1.395
+ $X2=4.195 $Y2=1.395
r202 26 54 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.105 $Y=1.47
+ $X2=4.105 $Y2=1.395
r203 26 28 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=4.105 $Y=1.47
+ $X2=4.105 $Y2=2.015
r204 25 53 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.675 $Y=1.395
+ $X2=3.585 $Y2=1.395
r205 24 54 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.015 $Y=1.395
+ $X2=4.105 $Y2=1.395
r206 24 25 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=4.015 $Y=1.395
+ $X2=3.675 $Y2=1.395
r207 21 53 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.585 $Y=1.47
+ $X2=3.585 $Y2=1.395
r208 21 23 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=3.585 $Y=1.47
+ $X2=3.585 $Y2=2.015
r209 20 52 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.155 $Y=1.395
+ $X2=3.065 $Y2=1.395
r210 19 53 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.495 $Y=1.395
+ $X2=3.585 $Y2=1.395
r211 19 20 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.495 $Y=1.395
+ $X2=3.155 $Y2=1.395
r212 16 52 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.065 $Y=1.47
+ $X2=3.065 $Y2=1.395
r213 16 18 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=3.065 $Y=1.47
+ $X2=3.065 $Y2=2.015
r214 15 51 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.635 $Y=1.395
+ $X2=2.545 $Y2=1.395
r215 14 52 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.975 $Y=1.395
+ $X2=3.065 $Y2=1.395
r216 14 15 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.975 $Y=1.395
+ $X2=2.635 $Y2=1.395
r217 11 51 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.545 $Y=1.47
+ $X2=2.545 $Y2=1.395
r218 11 13 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.545 $Y=1.47
+ $X2=2.545 $Y2=2.015
r219 9 51 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.455 $Y=1.395
+ $X2=2.545 $Y2=1.395
r220 9 50 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=2.455 $Y=1.395
+ $X2=2.22 $Y2=1.395
r221 8 66 13.6516 $w=3.79e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.655 $Y=1.16
+ $X2=1.555 $Y2=1.202
r222 8 49 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=1.655 $Y=1.16
+ $X2=2.07 $Y2=1.16
r223 4 66 20.1817 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.555 $Y=1.41
+ $X2=1.555 $Y2=1.202
r224 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.555 $Y=1.41
+ $X2=1.555 $Y2=1.985
r225 1 65 24.5487 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.53 $Y=0.995
+ $X2=1.53 $Y2=1.202
r226 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.53 $Y=0.995
+ $X2=1.53 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_8%A_321_47# 1 2 7 9 10 11 12 14 15 17 19 20
+ 22 24 25 27 29 30 32 34 35 37 39 40 42 44 45 46 47 48 49 50 52 55 58 63 64 67
+ 71 72 73
c157 73 0 1.36178e-19 $X=1.942 $Y=1.15
c158 72 0 1.93101e-20 $X=1.775 $Y=1.495
c159 71 0 1.41448e-19 $X=1.79 $Y=1.63
c160 58 0 1.13485e-20 $X=1.942 $Y=1.025
r161 71 72 6.07748 $w=3.98e-07 $l=1.35e-07 $layer=LI1_cond $X=1.775 $Y=1.63
+ $X2=1.775 $Y2=1.495
r162 67 69 6.83773 $w=5.58e-07 $l=2.65e-07 $layer=LI1_cond $X=1.855 $Y=0.56
+ $X2=1.855 $Y2=0.825
r163 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.71
+ $Y=1.16 $X2=6.71 $Y2=1.16
r164 61 73 2.06747 $w=2.5e-07 $l=1.93e-07 $layer=LI1_cond $X=2.135 $Y=1.15
+ $X2=1.942 $Y2=1.15
r165 61 63 210.897 $w=2.48e-07 $l=4.575e-06 $layer=LI1_cond $X=2.135 $Y=1.15
+ $X2=6.71 $Y2=1.15
r166 59 73 4.36486 $w=3.05e-07 $l=1.60078e-07 $layer=LI1_cond $X=1.862 $Y=1.275
+ $X2=1.942 $Y2=1.15
r167 59 72 11.2683 $w=2.23e-07 $l=2.2e-07 $layer=LI1_cond $X=1.862 $Y=1.275
+ $X2=1.862 $Y2=1.495
r168 58 73 4.36486 $w=3.05e-07 $l=1.25e-07 $layer=LI1_cond $X=1.942 $Y=1.025
+ $X2=1.942 $Y2=1.15
r169 58 69 5.98672 $w=3.83e-07 $l=2e-07 $layer=LI1_cond $X=1.942 $Y=1.025
+ $X2=1.942 $Y2=0.825
r170 53 71 1.87272 $w=3.98e-07 $l=6.5e-08 $layer=LI1_cond $X=1.775 $Y=1.695
+ $X2=1.775 $Y2=1.63
r171 53 55 17.7188 $w=3.98e-07 $l=6.15e-07 $layer=LI1_cond $X=1.775 $Y=1.695
+ $X2=1.775 $Y2=2.31
r172 51 64 31.8665 $w=3.35e-07 $l=1.85e-07 $layer=POLY_cond $X=6.525 $Y=1.127
+ $X2=6.71 $Y2=1.127
r173 51 52 13.4622 $w=2.42e-07 $l=2.30085e-07 $layer=POLY_cond $X=6.525 $Y=1.127
+ $X2=6.375 $Y2=0.96
r174 42 52 12.3158 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.45 $Y=0.96
+ $X2=6.375 $Y2=0.96
r175 42 44 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=6.45 $Y=0.96 $X2=6.45
+ $Y2=0.56
r176 41 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.005 $Y=1.035
+ $X2=5.93 $Y2=1.035
r177 40 52 13.4622 $w=2.42e-07 $l=7.5e-08 $layer=POLY_cond $X=6.375 $Y=1.035
+ $X2=6.375 $Y2=0.96
r178 40 41 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.375 $Y=1.035
+ $X2=6.005 $Y2=1.035
r179 37 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.93 $Y=0.96
+ $X2=5.93 $Y2=1.035
r180 37 39 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.93 $Y=0.96 $X2=5.93
+ $Y2=0.56
r181 36 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.485 $Y=1.035
+ $X2=5.41 $Y2=1.035
r182 35 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.855 $Y=1.035
+ $X2=5.93 $Y2=1.035
r183 35 36 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.855 $Y=1.035
+ $X2=5.485 $Y2=1.035
r184 32 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.41 $Y=0.96
+ $X2=5.41 $Y2=1.035
r185 32 34 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.41 $Y=0.96 $X2=5.41
+ $Y2=0.56
r186 31 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.965 $Y=1.035
+ $X2=4.89 $Y2=1.035
r187 30 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.335 $Y=1.035
+ $X2=5.41 $Y2=1.035
r188 30 31 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.335 $Y=1.035
+ $X2=4.965 $Y2=1.035
r189 27 48 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.89 $Y=0.96
+ $X2=4.89 $Y2=1.035
r190 27 29 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.89 $Y=0.96 $X2=4.89
+ $Y2=0.56
r191 26 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.445 $Y=1.035
+ $X2=4.37 $Y2=1.035
r192 25 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.815 $Y=1.035
+ $X2=4.89 $Y2=1.035
r193 25 26 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.815 $Y=1.035
+ $X2=4.445 $Y2=1.035
r194 22 47 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.37 $Y=0.96
+ $X2=4.37 $Y2=1.035
r195 22 24 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.37 $Y=0.96 $X2=4.37
+ $Y2=0.56
r196 21 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.925 $Y=1.035
+ $X2=3.85 $Y2=1.035
r197 20 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.295 $Y=1.035
+ $X2=4.37 $Y2=1.035
r198 20 21 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.295 $Y=1.035
+ $X2=3.925 $Y2=1.035
r199 17 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.85 $Y=0.96
+ $X2=3.85 $Y2=1.035
r200 17 19 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.85 $Y=0.96 $X2=3.85
+ $Y2=0.56
r201 16 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.405 $Y=1.035
+ $X2=3.33 $Y2=1.035
r202 15 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.775 $Y=1.035
+ $X2=3.85 $Y2=1.035
r203 15 16 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.775 $Y=1.035
+ $X2=3.405 $Y2=1.035
r204 12 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.33 $Y=0.96
+ $X2=3.33 $Y2=1.035
r205 12 14 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.33 $Y=0.96 $X2=3.33
+ $Y2=0.56
r206 10 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.255 $Y=1.035
+ $X2=3.33 $Y2=1.035
r207 10 11 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.255 $Y=1.035
+ $X2=2.885 $Y2=1.035
r208 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.81 $Y=0.96
+ $X2=2.885 $Y2=1.035
r209 7 9 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.81 $Y=0.96 $X2=2.81
+ $Y2=0.56
r210 2 71 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.645
+ $Y=1.485 $X2=1.79 $Y2=1.63
r211 2 55 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=1.645
+ $Y=1.485 $X2=1.79 $Y2=2.31
r212 1 67 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.605
+ $Y=0.235 $X2=1.79 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_8%A_124_297# 1 2 9 11 13 16 18 20 23 25 27
+ 30 32 34 37 39 41 44 46 48 51 53 55 56 58 61 65 75 77 79 98 101 104
r138 101 102 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=10.495 $Y=1.217
+ $X2=10.52 $Y2=1.217
r139 100 101 70.354 $w=3.22e-07 $l=4.7e-07 $layer=POLY_cond $X=10.025 $Y=1.217
+ $X2=10.495 $Y2=1.217
r140 99 100 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=10 $Y=1.217
+ $X2=10.025 $Y2=1.217
r141 97 99 1.49689 $w=3.22e-07 $l=1e-08 $layer=POLY_cond $X=9.99 $Y=1.217 $X2=10
+ $Y2=1.217
r142 97 98 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=9.99
+ $Y=1.16 $X2=9.99 $Y2=1.16
r143 95 97 65.1149 $w=3.22e-07 $l=4.35e-07 $layer=POLY_cond $X=9.555 $Y=1.217
+ $X2=9.99 $Y2=1.217
r144 94 95 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=9.53 $Y=1.217
+ $X2=9.555 $Y2=1.217
r145 93 94 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=9.085 $Y=1.217
+ $X2=9.53 $Y2=1.217
r146 92 93 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=9.06 $Y=1.217
+ $X2=9.085 $Y2=1.217
r147 91 92 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=8.615 $Y=1.217
+ $X2=9.06 $Y2=1.217
r148 90 91 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=8.59 $Y=1.217
+ $X2=8.615 $Y2=1.217
r149 89 90 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=8.145 $Y=1.217
+ $X2=8.59 $Y2=1.217
r150 88 89 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=8.12 $Y=1.217
+ $X2=8.145 $Y2=1.217
r151 87 88 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=7.675 $Y=1.217
+ $X2=8.12 $Y2=1.217
r152 86 87 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=7.65 $Y=1.217
+ $X2=7.675 $Y2=1.217
r153 84 86 50.8944 $w=3.22e-07 $l=3.4e-07 $layer=POLY_cond $X=7.31 $Y=1.217
+ $X2=7.65 $Y2=1.217
r154 84 85 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=7.31
+ $Y=1.16 $X2=7.31 $Y2=1.16
r155 82 84 15.7174 $w=3.22e-07 $l=1.05e-07 $layer=POLY_cond $X=7.205 $Y=1.217
+ $X2=7.31 $Y2=1.217
r156 81 82 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=7.18 $Y=1.217
+ $X2=7.205 $Y2=1.217
r157 78 98 104.872 $w=2.48e-07 $l=2.275e-06 $layer=LI1_cond $X=7.715 $Y=1.15
+ $X2=9.99 $Y2=1.15
r158 78 85 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=7.715 $Y=1.15
+ $X2=7.31 $Y2=1.15
r159 77 79 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=7.715 $Y=1.145
+ $X2=7.52 $Y2=1.145
r160 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.715 $Y=1.145
+ $X2=7.715 $Y2=1.145
r161 75 79 8.21162 $w=1.4e-07 $l=6.635e-06 $layer=MET1_cond $X=0.885 $Y=1.19
+ $X2=7.52 $Y2=1.19
r162 73 104 38.8182 $w=1.98e-07 $l=7e-07 $layer=LI1_cond $X=0.75 $Y=1.145
+ $X2=0.75 $Y2=0.445
r163 72 75 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.74 $Y=1.145
+ $X2=0.885 $Y2=1.145
r164 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.74 $Y=1.145
+ $X2=0.74 $Y2=1.145
r165 67 73 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.75 $Y=1.515
+ $X2=0.75 $Y2=1.145
r166 67 68 5.62585 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=0.75 $Y=1.515
+ $X2=0.75 $Y2=1.615
r167 65 68 36.2703 $w=1.83e-07 $l=6.05e-07 $layer=LI1_cond $X=0.757 $Y=2.22
+ $X2=0.757 $Y2=1.615
r168 59 102 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=10.52 $Y=1.025
+ $X2=10.52 $Y2=1.217
r169 59 61 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=10.52 $Y=1.025
+ $X2=10.52 $Y2=0.56
r170 56 101 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=10.495 $Y=1.41
+ $X2=10.495 $Y2=1.217
r171 56 58 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.495 $Y=1.41
+ $X2=10.495 $Y2=1.985
r172 53 100 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=10.025 $Y=1.41
+ $X2=10.025 $Y2=1.217
r173 53 55 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.025 $Y=1.41
+ $X2=10.025 $Y2=1.985
r174 49 99 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=10 $Y=1.025 $X2=10
+ $Y2=1.217
r175 49 51 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=10 $Y=1.025 $X2=10
+ $Y2=0.56
r176 46 95 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=9.555 $Y=1.41
+ $X2=9.555 $Y2=1.217
r177 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.555 $Y=1.41
+ $X2=9.555 $Y2=1.985
r178 42 94 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=9.53 $Y=1.025
+ $X2=9.53 $Y2=1.217
r179 42 44 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.53 $Y=1.025
+ $X2=9.53 $Y2=0.56
r180 39 93 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=9.085 $Y=1.41
+ $X2=9.085 $Y2=1.217
r181 39 41 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.085 $Y=1.41
+ $X2=9.085 $Y2=1.985
r182 35 92 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=9.06 $Y=1.025
+ $X2=9.06 $Y2=1.217
r183 35 37 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.06 $Y=1.025
+ $X2=9.06 $Y2=0.56
r184 32 91 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=8.615 $Y=1.41
+ $X2=8.615 $Y2=1.217
r185 32 34 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.615 $Y=1.41
+ $X2=8.615 $Y2=1.985
r186 28 90 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=8.59 $Y=1.025
+ $X2=8.59 $Y2=1.217
r187 28 30 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.59 $Y=1.025
+ $X2=8.59 $Y2=0.56
r188 25 89 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=8.145 $Y=1.41
+ $X2=8.145 $Y2=1.217
r189 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.145 $Y=1.41
+ $X2=8.145 $Y2=1.985
r190 21 88 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=8.12 $Y=1.025
+ $X2=8.12 $Y2=1.217
r191 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.12 $Y=1.025
+ $X2=8.12 $Y2=0.56
r192 18 87 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.675 $Y=1.41
+ $X2=7.675 $Y2=1.217
r193 18 20 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.675 $Y=1.41
+ $X2=7.675 $Y2=1.985
r194 14 86 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.65 $Y=1.025
+ $X2=7.65 $Y2=1.217
r195 14 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.65 $Y=1.025
+ $X2=7.65 $Y2=0.56
r196 11 82 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.205 $Y=1.41
+ $X2=7.205 $Y2=1.217
r197 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.205 $Y=1.41
+ $X2=7.205 $Y2=1.985
r198 7 81 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.18 $Y=1.025
+ $X2=7.18 $Y2=1.217
r199 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.18 $Y=1.025
+ $X2=7.18 $Y2=0.56
r200 2 65 600 $w=1.7e-07 $l=8.04239e-07 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.485 $X2=0.765 $Y2=2.22
r201 1 104 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.63
+ $Y=0.235 $X2=0.765 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_8%VPWR 1 2 3 4 5 6 19 21 25 27 30 33 36 38
+ 50 54 64 65 71 74 81 88
r143 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r144 88 91 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=5.9 $Y=2.36 $X2=5.9
+ $Y2=2.72
r145 85 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r146 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r147 81 84 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=4.86 $Y=2.36
+ $X2=4.86 $Y2=2.72
r148 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r149 74 77 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.82 $Y=2.36
+ $X2=3.82 $Y2=2.72
r150 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r151 64 65 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r152 62 65 1.30889 $w=4.8e-07 $l=4.6e-06 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=10.81 $Y2=2.72
r153 62 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r154 61 64 300.107 $w=1.68e-07 $l=4.6e-06 $layer=LI1_cond $X=6.21 $Y=2.72
+ $X2=10.81 $Y2=2.72
r155 61 62 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r156 59 91 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=6.115 $Y=2.72
+ $X2=5.9 $Y2=2.72
r157 59 61 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=6.115 $Y=2.72
+ $X2=6.21 $Y2=2.72
r158 58 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r159 58 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r160 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r161 55 77 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=4.035 $Y=2.72
+ $X2=3.82 $Y2=2.72
r162 55 57 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.035 $Y=2.72
+ $X2=4.37 $Y2=2.72
r163 54 84 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=4.645 $Y=2.72
+ $X2=4.86 $Y2=2.72
r164 54 57 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.645 $Y=2.72
+ $X2=4.37 $Y2=2.72
r165 53 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r166 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r167 50 77 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=3.605 $Y=2.72
+ $X2=3.82 $Y2=2.72
r168 50 52 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.605 $Y=2.72
+ $X2=3.45 $Y2=2.72
r169 49 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r170 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r171 46 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r172 46 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r173 45 48 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r174 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r175 43 71 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.405 $Y=2.72
+ $X2=1.212 $Y2=2.72
r176 43 45 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.405 $Y=2.72
+ $X2=1.61 $Y2=2.72
r177 42 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r178 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r179 39 68 5.0973 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=2.72
+ $X2=0.222 $Y2=2.72
r180 39 41 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.445 $Y=2.72
+ $X2=0.69 $Y2=2.72
r181 38 71 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=1.02 $Y=2.72
+ $X2=1.212 $Y2=2.72
r182 38 41 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.02 $Y=2.72
+ $X2=0.69 $Y2=2.72
r183 36 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r184 36 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r185 34 52 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.995 $Y=2.72
+ $X2=3.45 $Y2=2.72
r186 33 48 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.565 $Y=2.72
+ $X2=2.53 $Y2=2.72
r187 32 34 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.78 $Y=2.72
+ $X2=2.995 $Y2=2.72
r188 32 33 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.78 $Y=2.72
+ $X2=2.565 $Y2=2.72
r189 30 32 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.78 $Y=2.36
+ $X2=2.78 $Y2=2.72
r190 28 84 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=5.075 $Y=2.72
+ $X2=4.86 $Y2=2.72
r191 27 91 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=5.685 $Y=2.72
+ $X2=5.9 $Y2=2.72
r192 27 28 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.685 $Y=2.72
+ $X2=5.075 $Y2=2.72
r193 23 71 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.212 $Y=2.635
+ $X2=1.212 $Y2=2.72
r194 23 25 18.4092 $w=3.83e-07 $l=6.15e-07 $layer=LI1_cond $X=1.212 $Y=2.635
+ $X2=1.212 $Y2=2.02
r195 19 68 2.92581 $w=3.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.222 $Y2=2.72
r196 19 21 19.6876 $w=3.58e-07 $l=6.15e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.265 $Y2=2.02
r197 6 88 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.755
+ $Y=1.545 $X2=5.9 $Y2=2.36
r198 5 81 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.715
+ $Y=1.545 $X2=4.86 $Y2=2.36
r199 4 74 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.675
+ $Y=1.545 $X2=3.82 $Y2=2.36
r200 3 30 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=1.545 $X2=2.78 $Y2=2.36
r201 2 25 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=1.09
+ $Y=1.485 $X2=1.235 $Y2=2.02
r202 1 21 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_8%A_437_309# 1 2 3 4 5 6 7 8 9 30 32 33 36
+ 38 42 44 48 52 60 62 63 64 67
c107 67 0 7.91225e-20 $X=6.335 $Y=2.18
c108 44 0 7.91225e-20 $X=5.295 $Y=1.98
c109 38 0 7.91225e-20 $X=4.255 $Y=1.98
r110 66 67 18.2496 $w=5.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.895 $Y=2.18
+ $X2=6.335 $Y2=2.18
r111 58 60 19.7248 $w=5.68e-07 $l=9.4e-07 $layer=LI1_cond $X=9.79 $Y=2.18
+ $X2=10.73 $Y2=2.18
r112 56 58 19.7248 $w=5.68e-07 $l=9.4e-07 $layer=LI1_cond $X=8.85 $Y=2.18
+ $X2=9.79 $Y2=2.18
r113 54 56 19.7248 $w=5.68e-07 $l=9.4e-07 $layer=LI1_cond $X=7.91 $Y=2.18
+ $X2=8.85 $Y2=2.18
r114 52 66 0.209838 $w=5.68e-07 $l=1e-08 $layer=LI1_cond $X=6.905 $Y=2.18
+ $X2=6.895 $Y2=2.18
r115 52 54 21.0888 $w=5.68e-07 $l=1.005e-06 $layer=LI1_cond $X=6.905 $Y=2.18
+ $X2=7.91 $Y2=2.18
r116 51 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.465 $Y=1.98
+ $X2=5.38 $Y2=1.98
r117 51 67 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=5.465 $Y=1.98
+ $X2=6.335 $Y2=1.98
r118 46 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.38 $Y=2.065
+ $X2=5.38 $Y2=1.98
r119 46 48 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.38 $Y=2.065
+ $X2=5.38 $Y2=2.3
r120 45 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.425 $Y=1.98
+ $X2=4.34 $Y2=1.98
r121 44 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.295 $Y=1.98
+ $X2=5.38 $Y2=1.98
r122 44 45 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=5.295 $Y=1.98
+ $X2=4.425 $Y2=1.98
r123 40 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=2.065
+ $X2=4.34 $Y2=1.98
r124 40 42 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.34 $Y=2.065
+ $X2=4.34 $Y2=2.3
r125 39 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.385 $Y=1.98
+ $X2=3.3 $Y2=1.98
r126 38 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.255 $Y=1.98
+ $X2=4.34 $Y2=1.98
r127 38 39 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=4.255 $Y=1.98
+ $X2=3.385 $Y2=1.98
r128 34 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=2.065 $X2=3.3
+ $Y2=1.98
r129 34 36 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.3 $Y=2.065
+ $X2=3.3 $Y2=2.3
r130 32 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=1.98
+ $X2=3.3 $Y2=1.98
r131 32 33 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=3.215 $Y=1.98
+ $X2=2.395 $Y2=1.98
r132 28 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.27 $Y=2.065
+ $X2=2.395 $Y2=1.98
r133 28 30 10.833 $w=2.48e-07 $l=2.35e-07 $layer=LI1_cond $X=2.27 $Y=2.065
+ $X2=2.27 $Y2=2.3
r134 9 60 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=10.585
+ $Y=1.485 $X2=10.73 $Y2=2.02
r135 8 58 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=9.645
+ $Y=1.485 $X2=9.79 $Y2=2.02
r136 7 56 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=8.705
+ $Y=1.485 $X2=8.85 $Y2=2.02
r137 6 54 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=7.765
+ $Y=1.485 $X2=7.91 $Y2=2.02
r138 5 66 300 $w=1.7e-07 $l=1.01888e-06 $layer=licon1_PDIFF $count=2 $X=6.275
+ $Y=1.545 $X2=6.895 $Y2=2.3
r139 4 48 600 $w=1.7e-07 $l=8.24318e-07 $layer=licon1_PDIFF $count=1 $X=5.235
+ $Y=1.545 $X2=5.38 $Y2=2.3
r140 3 42 600 $w=1.7e-07 $l=8.24318e-07 $layer=licon1_PDIFF $count=1 $X=4.195
+ $Y=1.545 $X2=4.34 $Y2=2.3
r141 2 36 600 $w=1.7e-07 $l=8.24318e-07 $layer=licon1_PDIFF $count=1 $X=3.155
+ $Y=1.545 $X2=3.3 $Y2=2.3
r142 1 30 600 $w=1.7e-07 $l=8.15107e-07 $layer=licon1_PDIFF $count=1 $X=2.185
+ $Y=1.545 $X2=2.31 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_8%Z 1 2 3 4 5 6 7 8 25 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 71 75 77 81 88 90 93 96 101 106 109 115 120 121
r108 115 117 20.5793 $w=2.78e-07 $l=5e-07 $layer=LI1_cond $X=9.76 $Y=1.585
+ $X2=10.26 $Y2=1.585
r109 104 106 11.7302 $w=2.78e-07 $l=2.85e-07 $layer=LI1_cond $X=8.38 $Y=1.585
+ $X2=8.665 $Y2=1.585
r110 99 101 30.2516 $w=2.78e-07 $l=7.35e-07 $layer=LI1_cond $X=7.44 $Y=1.585
+ $X2=8.175 $Y2=1.585
r111 88 90 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=5.49 $Y=1.585
+ $X2=6.125 $Y2=1.585
r112 75 77 21.8141 $w=2.78e-07 $l=5.3e-07 $layer=LI1_cond $X=2.755 $Y=1.585
+ $X2=3.285 $Y2=1.585
r113 71 120 16.4635 $w=2.78e-07 $l=4e-07 $layer=LI1_cond $X=10.675 $Y=1.585
+ $X2=10.275 $Y2=1.585
r114 51 71 3.22874 $w=2.8e-07 $l=1.25e-07 $layer=LI1_cond $X=10.8 $Y=1.585
+ $X2=10.675 $Y2=1.585
r115 50 51 8.86994 $w=4.18e-07 $l=2.55e-07 $layer=LI1_cond $X=10.8 $Y=1.19
+ $X2=10.8 $Y2=1.445
r116 49 121 3.3405 $w=2.5e-07 $l=1.2e-07 $layer=LI1_cond $X=10.8 $Y=0.735
+ $X2=10.8 $Y2=0.855
r117 49 50 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=10.8 $Y=0.895
+ $X2=10.8 $Y2=1.19
r118 49 121 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=10.8 $Y=0.895
+ $X2=10.8 $Y2=0.855
r119 48 120 0.411587 $w=2.78e-07 $l=1e-08 $layer=LI1_cond $X=10.265 $Y=1.585
+ $X2=10.275 $Y2=1.585
r120 48 117 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=10.265 $Y=1.585
+ $X2=10.26 $Y2=1.585
r121 47 115 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=9.755 $Y=1.585
+ $X2=9.76 $Y2=1.585
r122 47 112 17.904 $w=2.78e-07 $l=4.35e-07 $layer=LI1_cond $X=9.755 $Y=1.585
+ $X2=9.32 $Y2=1.585
r123 46 112 4.73325 $w=2.78e-07 $l=1.15e-07 $layer=LI1_cond $X=9.205 $Y=1.585
+ $X2=9.32 $Y2=1.585
r124 46 109 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=9.205 $Y=1.585
+ $X2=9.2 $Y2=1.585
r125 45 109 21.8141 $w=2.78e-07 $l=5.3e-07 $layer=LI1_cond $X=8.67 $Y=1.585
+ $X2=9.2 $Y2=1.585
r126 45 106 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=8.67 $Y=1.585
+ $X2=8.665 $Y2=1.585
r127 44 104 8.02594 $w=2.78e-07 $l=1.95e-07 $layer=LI1_cond $X=8.185 $Y=1.585
+ $X2=8.38 $Y2=1.585
r128 44 101 0.411587 $w=2.78e-07 $l=1e-08 $layer=LI1_cond $X=8.185 $Y=1.585
+ $X2=8.175 $Y2=1.585
r129 43 99 11.7302 $w=2.78e-07 $l=2.85e-07 $layer=LI1_cond $X=7.155 $Y=1.585
+ $X2=7.44 $Y2=1.585
r130 43 96 1.23476 $w=2.78e-07 $l=3e-08 $layer=LI1_cond $X=7.155 $Y=1.585
+ $X2=7.125 $Y2=1.585
r131 42 96 17.4924 $w=2.78e-07 $l=4.25e-07 $layer=LI1_cond $X=6.7 $Y=1.585
+ $X2=7.125 $Y2=1.585
r132 42 93 0.823174 $w=2.78e-07 $l=2e-08 $layer=LI1_cond $X=6.7 $Y=1.585
+ $X2=6.68 $Y2=1.585
r133 41 93 22.2257 $w=2.78e-07 $l=5.4e-07 $layer=LI1_cond $X=6.14 $Y=1.585
+ $X2=6.68 $Y2=1.585
r134 41 90 0.61738 $w=2.78e-07 $l=1.5e-08 $layer=LI1_cond $X=6.14 $Y=1.585
+ $X2=6.125 $Y2=1.585
r135 40 88 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=5.485 $Y=1.585
+ $X2=5.49 $Y2=1.585
r136 39 40 22.8431 $w=2.78e-07 $l=5.55e-07 $layer=LI1_cond $X=4.93 $Y=1.585
+ $X2=5.485 $Y2=1.585
r137 38 39 23.0489 $w=2.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.37 $Y=1.585
+ $X2=4.93 $Y2=1.585
r138 38 81 18.933 $w=2.78e-07 $l=4.6e-07 $layer=LI1_cond $X=4.37 $Y=1.585
+ $X2=3.91 $Y2=1.585
r139 37 81 3.0869 $w=2.78e-07 $l=7.5e-08 $layer=LI1_cond $X=3.835 $Y=1.585
+ $X2=3.91 $Y2=1.585
r140 36 37 22.4315 $w=2.78e-07 $l=5.45e-07 $layer=LI1_cond $X=3.29 $Y=1.585
+ $X2=3.835 $Y2=1.585
r141 36 77 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=3.29 $Y=1.585
+ $X2=3.285 $Y2=1.585
r142 35 75 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=2.73 $Y=1.585
+ $X2=2.755 $Y2=1.585
r143 32 34 45.1374 $w=2.38e-07 $l=9.4e-07 $layer=LI1_cond $X=9.32 $Y=0.735
+ $X2=10.26 $Y2=0.735
r144 30 32 45.1374 $w=2.38e-07 $l=9.4e-07 $layer=LI1_cond $X=8.38 $Y=0.735
+ $X2=9.32 $Y2=0.735
r145 27 30 45.1374 $w=2.38e-07 $l=9.4e-07 $layer=LI1_cond $X=7.44 $Y=0.735
+ $X2=8.38 $Y2=0.735
r146 25 49 3.47969 $w=2.4e-07 $l=1.25e-07 $layer=LI1_cond $X=10.675 $Y=0.735
+ $X2=10.8 $Y2=0.735
r147 25 34 19.9277 $w=2.38e-07 $l=4.15e-07 $layer=LI1_cond $X=10.675 $Y=0.735
+ $X2=10.26 $Y2=0.735
r148 8 117 600 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=10.115
+ $Y=1.485 $X2=10.26 $Y2=1.64
r149 7 112 600 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=9.175
+ $Y=1.485 $X2=9.32 $Y2=1.64
r150 6 104 600 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=8.235
+ $Y=1.485 $X2=8.38 $Y2=1.64
r151 5 99 600 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=7.295
+ $Y=1.485 $X2=7.44 $Y2=1.64
r152 4 34 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=10.075
+ $Y=0.235 $X2=10.26 $Y2=0.76
r153 3 32 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=9.135
+ $Y=0.235 $X2=9.32 $Y2=0.76
r154 2 30 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=8.195
+ $Y=0.235 $X2=8.38 $Y2=0.76
r155 1 27 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=7.255
+ $Y=0.235 $X2=7.44 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_8%VGND 1 2 3 4 5 6 19 21 23 25 26 32 34 39
+ 51 60 61 75 82 89
r128 89 92 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=6.19 $Y=0 $X2=6.19
+ $Y2=0.36
r129 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r130 82 85 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=4.11 $Y=0 $X2=4.11
+ $Y2=0.36
r131 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r132 76 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r133 75 78 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.07 $Y=0 $X2=3.07
+ $Y2=0.36
r134 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r135 60 61 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r136 58 61 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=6.67 $Y=0 $X2=10.81
+ $Y2=0
r137 58 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r138 57 60 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=6.67 $Y=0
+ $X2=10.81 $Y2=0
r139 57 58 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r140 55 89 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=6.405 $Y=0 $X2=6.19
+ $Y2=0
r141 55 57 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.405 $Y=0
+ $X2=6.67 $Y2=0
r142 54 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r143 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r144 51 89 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=5.975 $Y=0 $X2=6.19
+ $Y2=0
r145 51 53 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.975 $Y=0
+ $X2=5.75 $Y2=0
r146 50 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r147 50 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=3.91
+ $Y2=0
r148 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r149 47 82 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=4.325 $Y=0 $X2=4.11
+ $Y2=0
r150 47 49 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.325 $Y=0
+ $X2=4.83 $Y2=0
r151 46 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r152 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r153 43 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r154 43 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r155 42 45 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r156 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r157 40 42 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.405 $Y=0
+ $X2=1.61 $Y2=0
r158 39 75 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.855 $Y=0 $X2=3.07
+ $Y2=0
r159 39 45 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.855 $Y=0
+ $X2=2.53 $Y2=0
r160 38 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r161 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r162 35 64 5.0973 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r163 35 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.69
+ $Y2=0
r164 34 71 10.7761 $w=3.83e-07 $l=3.6e-07 $layer=LI1_cond $X=1.212 $Y=0
+ $X2=1.212 $Y2=0.36
r165 34 40 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.212 $Y=0
+ $X2=1.405 $Y2=0
r166 34 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r167 34 37 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=0.69
+ $Y2=0
r168 32 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r169 32 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r170 28 53 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.365 $Y=0
+ $X2=5.75 $Y2=0
r171 26 49 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.935 $Y=0
+ $X2=4.83 $Y2=0
r172 25 30 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=5.15 $Y=0 $X2=5.15
+ $Y2=0.36
r173 25 28 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=5.15 $Y=0 $X2=5.365
+ $Y2=0
r174 25 26 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=5.15 $Y=0 $X2=4.935
+ $Y2=0
r175 24 75 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=3.285 $Y=0 $X2=3.07
+ $Y2=0
r176 23 82 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=3.895 $Y=0 $X2=4.11
+ $Y2=0
r177 23 24 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.895 $Y=0
+ $X2=3.285 $Y2=0
r178 19 64 2.92581 $w=3.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.222 $Y2=0
r179 19 21 8.80338 $w=3.58e-07 $l=2.75e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.265 $Y2=0.36
r180 6 92 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=6.005
+ $Y=0.235 $X2=6.19 $Y2=0.36
r181 5 30 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=4.965
+ $Y=0.235 $X2=5.15 $Y2=0.36
r182 4 85 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=3.925
+ $Y=0.235 $X2=4.11 $Y2=0.36
r183 3 78 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=2.885
+ $Y=0.235 $X2=3.07 $Y2=0.36
r184 2 71 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.235 $X2=1.235 $Y2=0.36
r185 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_8%A_485_47# 1 2 3 4 5 6 7 8 9 28 31 32 33 36
+ 38 41 43 46 56 58 59 60 61
r115 64 65 5.22619 $w=4.28e-07 $l=1.95e-07 $layer=LI1_cond $X=6.84 $Y=0.56
+ $X2=6.84 $Y2=0.755
r116 61 64 5.62821 $w=4.28e-07 $l=2.1e-07 $layer=LI1_cond $X=6.84 $Y=0.35
+ $X2=6.84 $Y2=0.56
r117 54 56 54.8708 $w=1.88e-07 $l=9.4e-07 $layer=LI1_cond $X=9.79 $Y=0.35
+ $X2=10.73 $Y2=0.35
r118 52 54 54.8708 $w=1.88e-07 $l=9.4e-07 $layer=LI1_cond $X=8.85 $Y=0.35
+ $X2=9.79 $Y2=0.35
r119 50 52 54.8708 $w=1.88e-07 $l=9.4e-07 $layer=LI1_cond $X=7.91 $Y=0.35
+ $X2=8.85 $Y2=0.35
r120 48 61 5.54258 $w=1.9e-07 $l=2.15e-07 $layer=LI1_cond $X=7.055 $Y=0.35
+ $X2=6.84 $Y2=0.35
r121 48 50 49.9091 $w=1.88e-07 $l=8.55e-07 $layer=LI1_cond $X=7.055 $Y=0.35
+ $X2=7.91 $Y2=0.35
r122 47 60 5.58832 $w=2e-07 $l=1.1e-07 $layer=LI1_cond $X=5.805 $Y=0.755
+ $X2=5.695 $Y2=0.755
r123 46 65 5.23352 $w=2e-07 $l=2.15e-07 $layer=LI1_cond $X=6.625 $Y=0.755
+ $X2=6.84 $Y2=0.755
r124 46 47 45.4727 $w=1.98e-07 $l=8.2e-07 $layer=LI1_cond $X=6.625 $Y=0.755
+ $X2=5.805 $Y2=0.755
r125 43 60 1.0017 $w=2.2e-07 $l=1e-07 $layer=LI1_cond $X=5.695 $Y=0.655
+ $X2=5.695 $Y2=0.755
r126 43 45 5.26818 $w=2.2e-07 $l=9.5e-08 $layer=LI1_cond $X=5.695 $Y=0.655
+ $X2=5.695 $Y2=0.56
r127 42 59 5.58832 $w=2e-07 $l=1.1e-07 $layer=LI1_cond $X=4.765 $Y=0.755
+ $X2=4.655 $Y2=0.755
r128 41 60 5.58832 $w=2e-07 $l=1.1e-07 $layer=LI1_cond $X=5.585 $Y=0.755
+ $X2=5.695 $Y2=0.755
r129 41 42 45.4727 $w=1.98e-07 $l=8.2e-07 $layer=LI1_cond $X=5.585 $Y=0.755
+ $X2=4.765 $Y2=0.755
r130 38 59 1.0017 $w=2.2e-07 $l=1e-07 $layer=LI1_cond $X=4.655 $Y=0.655
+ $X2=4.655 $Y2=0.755
r131 38 40 5.26818 $w=2.2e-07 $l=9.5e-08 $layer=LI1_cond $X=4.655 $Y=0.655
+ $X2=4.655 $Y2=0.56
r132 37 58 5.58832 $w=2e-07 $l=1.1e-07 $layer=LI1_cond $X=3.725 $Y=0.755
+ $X2=3.615 $Y2=0.755
r133 36 59 5.58832 $w=2e-07 $l=1.1e-07 $layer=LI1_cond $X=4.545 $Y=0.755
+ $X2=4.655 $Y2=0.755
r134 36 37 45.4727 $w=1.98e-07 $l=8.2e-07 $layer=LI1_cond $X=4.545 $Y=0.755
+ $X2=3.725 $Y2=0.755
r135 33 58 1.0017 $w=2.2e-07 $l=1e-07 $layer=LI1_cond $X=3.615 $Y=0.655
+ $X2=3.615 $Y2=0.755
r136 33 35 5.26818 $w=2.2e-07 $l=9.5e-08 $layer=LI1_cond $X=3.615 $Y=0.655
+ $X2=3.615 $Y2=0.56
r137 31 58 5.58832 $w=2e-07 $l=1.1e-07 $layer=LI1_cond $X=3.505 $Y=0.755
+ $X2=3.615 $Y2=0.755
r138 31 32 45.4727 $w=1.98e-07 $l=8.2e-07 $layer=LI1_cond $X=3.505 $Y=0.755
+ $X2=2.685 $Y2=0.755
r139 28 32 7.70722 $w=2e-07 $l=2.34734e-07 $layer=LI1_cond $X=2.495 $Y=0.655
+ $X2=2.685 $Y2=0.755
r140 28 30 3.05 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.495 $Y=0.655
+ $X2=2.495 $Y2=0.56
r141 9 56 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=10.595
+ $Y=0.235 $X2=10.73 $Y2=0.36
r142 8 54 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=9.605
+ $Y=0.235 $X2=9.79 $Y2=0.36
r143 7 52 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=8.665
+ $Y=0.235 $X2=8.85 $Y2=0.36
r144 6 50 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=7.725
+ $Y=0.235 $X2=7.91 $Y2=0.36
r145 5 64 182 $w=1.7e-07 $l=4.57848e-07 $layer=licon1_NDIFF $count=1 $X=6.525
+ $Y=0.235 $X2=6.845 $Y2=0.56
r146 4 45 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=5.485
+ $Y=0.235 $X2=5.67 $Y2=0.56
r147 3 40 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=4.445
+ $Y=0.235 $X2=4.63 $Y2=0.56
r148 2 35 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=3.405
+ $Y=0.235 $X2=3.59 $Y2=0.56
r149 1 30 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.55 $Y2=0.56
.ends

