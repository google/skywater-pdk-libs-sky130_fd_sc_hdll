* NGSPICE file created from sky130_fd_sc_hdll__nand4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__nand4_4 A B C D VGND VNB VPB VPWR Y
M1000 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=3.15e+12p pd=2.43e+07u as=2.32e+12p ps=2.064e+07u
M1001 VPWR D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_27_47# D VGND VNB nshort w=650000u l=150000u
+  ad=9.62e+11p pd=9.46e+06u as=4.16e+11p ps=3.88e+06u
M1003 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_883_47# B a_485_47# VNB nshort w=650000u l=150000u
+  ad=1.0335e+12p pd=9.68e+06u as=8.645e+11p ps=7.86e+06u
M1006 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_485_47# B a_883_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_883_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1009 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y A a_883_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_47# C a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_883_47# B a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_485_47# C a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_485_47# B a_883_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND D a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_47# D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_883_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_27_47# C a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y A a_883_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_485_47# C a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND D a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

