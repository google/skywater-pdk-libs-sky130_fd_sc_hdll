* File: sky130_fd_sc_hdll__a2bb2o_1.spice
* Created: Thu Aug 27 18:54:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a2bb2o_1.pex.spice"
.subckt sky130_fd_sc_hdll__a2bb2o_1  VNB VPB A1_N A2_N B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_79_21#_M1011_g N_X_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.174589 AS=0.169 PD=1.4215 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1008 N_A_243_47#_M1008_d N_A1_N_M1008_g N_VGND_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.112811 PD=0.69 PS=0.918505 NRD=0 NRS=55.704 M=1 R=2.8
+ SA=75000.9 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A2_N_M1006_g N_A_243_47#_M1008_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1785 AS=0.0567 PD=1.27 PS=0.69 NRD=17.136 NRS=0 M=1 R=2.8
+ SA=75001.3 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1002 N_A_79_21#_M1002_d N_A_243_47#_M1002_g N_VGND_M1006_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1785 PD=0.69 PS=1.27 NRD=0 NRS=34.284 M=1 R=2.8
+ SA=75002.3 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 A_611_47# N_B2_M1001_g N_A_79_21#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0567 PD=0.75 PS=0.69 NRD=31.428 NRS=0 M=1 R=2.8 SA=75002.7
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_B1_M1007_g A_611_47# VNB NSHORT L=0.15 W=0.42 AD=0.1302
+ AS=0.0693 PD=1.46 PS=0.75 NRD=12.852 NRS=31.428 M=1 R=2.8 SA=75003.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_79_21#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.240423 AS=0.27 PD=2.02817 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1004 A_241_297# N_A1_N_M1004_g N_VPWR_M1003_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.05145 AS=0.100977 PD=0.665 PS=0.851831 NRD=31.6579 NRS=86.9558 M=1
+ R=2.33333 SA=90000.8 SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1009 N_A_243_47#_M1009_d N_A2_N_M1009_g A_241_297# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.1155 AS=0.05145 PD=1.39 PS=0.665 NRD=2.3443 NRS=31.6579 M=1 R=2.33333
+ SA=90001.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1000 N_A_525_413#_M1000_d N_A_243_47#_M1000_g N_A_79_21#_M1000_s VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.0609 AS=0.1134 PD=0.71 PS=1.38 NRD=2.3443 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_B2_M1010_g N_A_525_413#_M1000_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.063 AS=0.0609 PD=0.72 PS=0.71 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.6 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1005 N_A_525_413#_M1005_d N_B1_M1005_g N_VPWR_M1010_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.063 PD=1.38 PS=0.72 NRD=2.3443 NRS=7.0329 M=1 R=2.33333
+ SA=90001.1 SB=90000.2 A=0.0756 P=1.2 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hdll__a2bb2o_1.pxi.spice"
*
.ends
*
*
