* File: sky130_fd_sc_hdll__a31oi_2.pxi.spice
* Created: Wed Sep  2 08:20:20 2020
* 
x_PM_SKY130_FD_SC_HDLL__A31OI_2%A3 N_A3_c_67_n N_A3_M1001_g N_A3_c_64_n
+ N_A3_M1002_g N_A3_c_68_n N_A3_M1006_g N_A3_c_65_n N_A3_M1012_g A3 A3
+ N_A3_c_66_n A3 PM_SKY130_FD_SC_HDLL__A31OI_2%A3
x_PM_SKY130_FD_SC_HDLL__A31OI_2%A2 N_A2_c_104_n N_A2_M1005_g N_A2_c_108_n
+ N_A2_M1011_g N_A2_c_109_n N_A2_M1015_g N_A2_c_105_n N_A2_M1013_g A2 A2
+ N_A2_c_106_n A2 A2 A2 PM_SKY130_FD_SC_HDLL__A31OI_2%A2
x_PM_SKY130_FD_SC_HDLL__A31OI_2%A1 N_A1_c_155_n N_A1_M1007_g N_A1_c_150_n
+ N_A1_c_151_n N_A1_c_152_n N_A1_M1000_g N_A1_c_158_n N_A1_M1009_g N_A1_c_153_n
+ N_A1_M1004_g A1 A1 N_A1_c_154_n A1 A1 A1 A1 PM_SKY130_FD_SC_HDLL__A31OI_2%A1
x_PM_SKY130_FD_SC_HDLL__A31OI_2%B1 N_B1_c_208_n N_B1_M1003_g N_B1_c_214_n
+ N_B1_M1008_g N_B1_c_209_n N_B1_c_210_n N_B1_M1014_g N_B1_c_216_n N_B1_M1010_g
+ N_B1_c_211_n B1 B1 B1 N_B1_c_213_n N_B1_c_228_p B1
+ PM_SKY130_FD_SC_HDLL__A31OI_2%B1
x_PM_SKY130_FD_SC_HDLL__A31OI_2%A_27_297# N_A_27_297#_M1001_d
+ N_A_27_297#_M1006_d N_A_27_297#_M1015_d N_A_27_297#_M1009_d
+ N_A_27_297#_M1010_s N_A_27_297#_c_263_n N_A_27_297#_c_270_n
+ N_A_27_297#_c_275_n N_A_27_297#_c_322_p N_A_27_297#_c_280_n
+ N_A_27_297#_c_283_n N_A_27_297#_c_281_n N_A_27_297#_c_285_n
+ N_A_27_297#_c_267_n N_A_27_297#_c_274_n N_A_27_297#_c_296_p
+ PM_SKY130_FD_SC_HDLL__A31OI_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A31OI_2%VPWR N_VPWR_M1001_s N_VPWR_M1011_s
+ N_VPWR_M1007_s N_VPWR_c_330_n N_VPWR_c_331_n VPWR N_VPWR_c_332_n
+ N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_329_n N_VPWR_c_336_n N_VPWR_c_337_n
+ N_VPWR_c_338_n N_VPWR_c_339_n PM_SKY130_FD_SC_HDLL__A31OI_2%VPWR
x_PM_SKY130_FD_SC_HDLL__A31OI_2%Y N_Y_M1000_d N_Y_M1004_d N_Y_M1014_s
+ N_Y_M1008_d N_Y_c_400_n N_Y_c_419_n N_Y_c_403_n N_Y_c_427_n N_Y_c_431_n
+ N_Y_c_401_n Y Y Y Y PM_SKY130_FD_SC_HDLL__A31OI_2%Y
x_PM_SKY130_FD_SC_HDLL__A31OI_2%A_27_47# N_A_27_47#_M1002_d N_A_27_47#_M1012_d
+ N_A_27_47#_M1013_s N_A_27_47#_c_475_n PM_SKY130_FD_SC_HDLL__A31OI_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__A31OI_2%VGND N_VGND_M1002_s N_VGND_M1003_d
+ N_VGND_c_497_n N_VGND_c_498_n VGND N_VGND_c_499_n N_VGND_c_500_n
+ N_VGND_c_501_n N_VGND_c_502_n PM_SKY130_FD_SC_HDLL__A31OI_2%VGND
x_PM_SKY130_FD_SC_HDLL__A31OI_2%A_297_47# N_A_297_47#_M1005_d
+ N_A_297_47#_M1000_s N_A_297_47#_c_551_n
+ PM_SKY130_FD_SC_HDLL__A31OI_2%A_297_47#
cc_1 VNB N_A3_c_64_n 0.0219558f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB N_A3_c_65_n 0.0167331f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB N_A3_c_66_n 0.0660896f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_4 VNB N_A2_c_104_n 0.0171772f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_A2_c_105_n 0.0229091f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_6 VNB N_A2_c_106_n 0.0366368f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_7 VNB A2 0.00396393f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A1_c_150_n 0.0243424f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_9 VNB N_A1_c_151_n 0.0191259f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_10 VNB N_A1_c_152_n 0.0227091f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_11 VNB N_A1_c_153_n 0.0166589f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_12 VNB N_A1_c_154_n 0.030534f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.202
cc_13 VNB N_B1_c_208_n 0.0179375f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_14 VNB N_B1_c_209_n 0.0167081f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_15 VNB N_B1_c_210_n 0.023158f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_16 VNB N_B1_c_211_n 0.0136431f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_17 VNB B1 0.00812034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B1_c_213_n 0.0358329f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.16
cc_19 VNB N_VPWR_c_329_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_400_n 0.00222757f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_21 VNB N_Y_c_401_n 0.0226742f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB Y 0.00568277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_475_n 0.0110136f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_497_n 0.00913142f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_25 VNB N_VGND_c_498_n 0.07583f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_26 VNB N_VGND_c_499_n 0.0157127f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_500_n 0.0189906f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_501_n 0.261129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_502_n 0.0085923f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_30 VNB N_A_297_47#_c_551_n 0.00778212f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_31 VPB N_A3_c_67_n 0.0188351f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_32 VPB N_A3_c_68_n 0.0162218f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_33 VPB A3 0.00703028f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_34 VPB N_A3_c_66_n 0.0311433f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_35 VPB N_A2_c_108_n 0.0152026f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_36 VPB N_A2_c_109_n 0.0159312f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_37 VPB N_A2_c_106_n 0.0194368f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_38 VPB A2 0.00129908f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A1_c_155_n 0.0197872f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_40 VPB N_A1_c_150_n 0.0128374f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_41 VPB N_A1_c_151_n 0.00722592f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_42 VPB N_A1_c_158_n 0.019949f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_43 VPB N_A1_c_154_n 0.0212068f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.202
cc_44 VPB A1 0.00115016f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_B1_c_214_n 0.0172362f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_46 VPB N_B1_c_209_n 0.00918527f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_47 VPB N_B1_c_216_n 0.0195761f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_48 VPB N_B1_c_211_n 0.0067642f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_49 VPB B1 0.0131071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_B1_c_213_n 0.0175721f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.16
cc_51 VPB N_VPWR_c_330_n 4.04661e-19 $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_52 VPB N_VPWR_c_331_n 4.04661e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_332_n 0.0159043f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_333_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.16
cc_55 VPB N_VPWR_c_334_n 0.047288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_329_n 0.0475109f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_336_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_337_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_338_n 0.02038f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_339_n 0.0217026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_Y_c_403_n 0.00626458f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_62 VPB Y 4.15115e-19 $X=-0.19 $Y=1.305 $X2=0.745 $Y2=1.305
cc_63 VPB Y 0.00279783f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 N_A3_c_65_n N_A2_c_104_n 0.0230895f $X=0.99 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_65 N_A3_c_68_n N_A2_c_108_n 0.0213366f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_66 A3 N_A2_c_106_n 3.06355e-19 $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_67 N_A3_c_66_n N_A2_c_106_n 0.0230895f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_68 N_A3_c_68_n A2 0.00198172f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_69 A3 A2 0.0342759f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_70 N_A3_c_66_n A2 0.00450289f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_71 A3 N_A_27_297#_M1001_d 0.00947317f $X=0.66 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_72 N_A3_c_67_n N_A_27_297#_c_263_n 0.0106972f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_73 N_A3_c_68_n N_A_27_297#_c_263_n 0.0165376f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_74 A3 N_A_27_297#_c_263_n 0.0277816f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_75 N_A3_c_66_n N_A_27_297#_c_263_n 8.79699e-19 $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_76 A3 N_A_27_297#_c_267_n 0.0151524f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_77 N_A3_c_66_n N_A_27_297#_c_267_n 7.14729e-19 $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_78 A3 N_VPWR_M1001_s 0.00199847f $X=0.66 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_79 N_A3_c_67_n N_VPWR_c_330_n 0.0139279f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A3_c_68_n N_VPWR_c_330_n 0.00931793f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A3_c_68_n N_VPWR_c_331_n 5.73683e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A3_c_67_n N_VPWR_c_332_n 0.00427505f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A3_c_68_n N_VPWR_c_333_n 0.00622633f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A3_c_67_n N_VPWR_c_329_n 0.00485802f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A3_c_68_n N_VPWR_c_329_n 0.00550537f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A3_c_64_n N_A_27_47#_c_475_n 0.00938548f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_87 N_A3_c_65_n N_A_27_47#_c_475_n 0.0146664f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_88 A3 N_A_27_47#_c_475_n 0.0513119f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_89 N_A3_c_66_n N_A_27_47#_c_475_n 0.0112233f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_90 N_A3_c_65_n N_VGND_c_498_n 0.00428022f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A3_c_64_n N_VGND_c_499_n 0.00199743f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_92 N_A3_c_64_n N_VGND_c_501_n 0.00369362f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A3_c_65_n N_VGND_c_501_n 0.00583944f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_94 N_A3_c_64_n N_VGND_c_502_n 0.0184487f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A3_c_65_n N_VGND_c_502_n 0.00317372f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A3_c_65_n N_A_297_47#_c_551_n 5.01868e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A2_c_109_n N_A1_c_155_n 0.0213245f $X=1.905 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_98 A2 N_A1_c_155_n 6.32254e-19 $X=1.775 $Y=1.22 $X2=-0.19 $Y2=-0.24
cc_99 N_A2_c_106_n N_A1_c_151_n 0.020839f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_100 A2 N_A1_c_151_n 0.00153975f $X=1.775 $Y=1.22 $X2=0 $Y2=0
cc_101 N_A2_c_109_n A1 6.92457e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A2_c_106_n A1 0.00166684f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_103 A2 A1 0.0247718f $X=1.775 $Y=1.22 $X2=0 $Y2=0
cc_104 A2 N_A_27_297#_M1006_d 0.00288073f $X=1.775 $Y=1.22 $X2=0 $Y2=0
cc_105 N_A2_c_108_n N_A_27_297#_c_270_n 0.0106972f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_106 N_A2_c_109_n N_A_27_297#_c_270_n 0.0138319f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_107 N_A2_c_106_n N_A_27_297#_c_270_n 8.82066e-19 $X=1.905 $Y=1.202 $X2=0
+ $Y2=0
cc_108 A2 N_A_27_297#_c_270_n 0.0345505f $X=1.775 $Y=1.22 $X2=0 $Y2=0
cc_109 A2 N_A_27_297#_c_274_n 0.0120328f $X=1.775 $Y=1.22 $X2=0 $Y2=0
cc_110 A2 N_VPWR_M1011_s 0.00195154f $X=1.775 $Y=1.22 $X2=0 $Y2=0
cc_111 N_A2_c_108_n N_VPWR_c_330_n 5.29587e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A2_c_108_n N_VPWR_c_331_n 0.0122621f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A2_c_109_n N_VPWR_c_331_n 0.010376f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A2_c_108_n N_VPWR_c_333_n 0.00427505f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A2_c_108_n N_VPWR_c_329_n 0.0039718f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A2_c_109_n N_VPWR_c_329_n 0.00550537f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A2_c_109_n N_VPWR_c_338_n 0.00622633f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A2_c_104_n N_A_27_47#_c_475_n 0.0101179f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A2_c_105_n N_A_27_47#_c_475_n 0.0120394f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A2_c_106_n N_A_27_47#_c_475_n 0.0042599f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_121 A2 N_A_27_47#_c_475_n 0.0527138f $X=1.775 $Y=1.22 $X2=0 $Y2=0
cc_122 N_A2_c_104_n N_VGND_c_498_n 0.00415639f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A2_c_105_n N_VGND_c_498_n 0.00366111f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A2_c_104_n N_VGND_c_501_n 0.0060278f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A2_c_105_n N_VGND_c_501_n 0.00685947f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A2_c_104_n N_A_297_47#_c_551_n 0.00379151f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A2_c_105_n N_A_297_47#_c_551_n 0.0101156f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A1_c_153_n N_B1_c_208_n 0.0152532f $X=3.47 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_129 N_A1_c_158_n N_B1_c_214_n 0.0250036f $X=3.445 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A1_c_154_n N_B1_c_211_n 0.0152532f $X=3.445 $Y=1.202 $X2=0 $Y2=0
cc_131 N_A1_c_155_n N_A_27_297#_c_275_n 0.0146157f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A1_c_150_n N_A_27_297#_c_275_n 0.00221727f $X=2.895 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A1_c_158_n N_A_27_297#_c_275_n 0.0154731f $X=3.445 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A1_c_154_n N_A_27_297#_c_275_n 0.00645621f $X=3.445 $Y=1.202 $X2=0
+ $Y2=0
cc_135 A1 N_A_27_297#_c_275_n 0.0558049f $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_136 N_A1_c_158_n N_A_27_297#_c_280_n 0.00544766f $X=3.445 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A1_c_158_n N_A_27_297#_c_281_n 0.00197231f $X=3.445 $Y=1.41 $X2=0 $Y2=0
cc_138 A1 N_VPWR_M1007_s 0.0102719f $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_139 N_A1_c_155_n N_VPWR_c_331_n 0.00111357f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A1_c_158_n N_VPWR_c_334_n 0.00702461f $X=3.445 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A1_c_155_n N_VPWR_c_329_n 0.00852407f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A1_c_158_n N_VPWR_c_329_n 0.00872812f $X=3.445 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A1_c_155_n N_VPWR_c_338_n 0.00702461f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A1_c_155_n N_VPWR_c_339_n 0.0140185f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A1_c_158_n N_VPWR_c_339_n 0.0148324f $X=3.445 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A1_c_150_n N_Y_c_400_n 0.00770192f $X=2.895 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A1_c_152_n N_Y_c_400_n 0.0089331f $X=2.97 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A1_c_154_n N_Y_c_400_n 0.00638627f $X=3.445 $Y=1.202 $X2=0 $Y2=0
cc_149 A1 N_Y_c_400_n 0.0382206f $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_150 N_A1_c_152_n Y 4.93458e-19 $X=2.97 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A1_c_153_n Y 0.00871709f $X=3.47 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A1_c_158_n Y 0.0104403f $X=3.445 $Y=1.41 $X2=0 $Y2=0
cc_153 A1 Y 0.0073984f $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_154 N_A1_c_152_n Y 0.00312095f $X=2.97 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A1_c_158_n Y 0.00131249f $X=3.445 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A1_c_153_n Y 0.00389735f $X=3.47 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A1_c_154_n Y 0.0188789f $X=3.445 $Y=1.202 $X2=0 $Y2=0
cc_158 A1 Y 0.0281152f $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_159 N_A1_c_151_n N_A_27_47#_c_475_n 0.00121664f $X=2.475 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A1_c_153_n N_VGND_c_497_n 0.001051f $X=3.47 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A1_c_152_n N_VGND_c_498_n 0.00366111f $X=2.97 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A1_c_153_n N_VGND_c_498_n 0.00427876f $X=3.47 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A1_c_152_n N_VGND_c_501_n 0.00681466f $X=2.97 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A1_c_153_n N_VGND_c_501_n 0.00626657f $X=3.47 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A1_c_151_n N_A_297_47#_c_551_n 0.00514306f $X=2.475 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A1_c_152_n N_A_297_47#_c_551_n 0.0101156f $X=2.97 $Y=0.995 $X2=0 $Y2=0
cc_167 A1 N_A_297_47#_c_551_n 0.00716467f $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_168 B1 N_A_27_297#_M1010_s 0.0061467f $X=4.73 $Y=1.445 $X2=0 $Y2=0
cc_169 N_B1_c_214_n N_A_27_297#_c_283_n 0.0147897f $X=4.005 $Y=1.41 $X2=0 $Y2=0
cc_170 N_B1_c_216_n N_A_27_297#_c_283_n 0.0142164f $X=4.555 $Y=1.41 $X2=0 $Y2=0
cc_171 B1 N_A_27_297#_c_285_n 0.0140093f $X=4.73 $Y=1.445 $X2=0 $Y2=0
cc_172 N_B1_c_213_n N_A_27_297#_c_285_n 8.57558e-19 $X=4.555 $Y=1.202 $X2=0
+ $Y2=0
cc_173 N_B1_c_228_p N_A_27_297#_c_285_n 2.86897e-19 $X=4.715 $Y=1.175 $X2=0
+ $Y2=0
cc_174 N_B1_c_214_n N_VPWR_c_334_n 0.00429453f $X=4.005 $Y=1.41 $X2=0 $Y2=0
cc_175 N_B1_c_216_n N_VPWR_c_334_n 0.00429453f $X=4.555 $Y=1.41 $X2=0 $Y2=0
cc_176 N_B1_c_214_n N_VPWR_c_329_n 0.00648608f $X=4.005 $Y=1.41 $X2=0 $Y2=0
cc_177 N_B1_c_216_n N_VPWR_c_329_n 0.00718299f $X=4.555 $Y=1.41 $X2=0 $Y2=0
cc_178 N_B1_c_208_n N_Y_c_419_n 0.00593249f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_179 N_B1_c_214_n N_Y_c_403_n 0.020604f $X=4.005 $Y=1.41 $X2=0 $Y2=0
cc_180 N_B1_c_209_n N_Y_c_403_n 0.00974235f $X=4.455 $Y=1.16 $X2=0 $Y2=0
cc_181 N_B1_c_216_n N_Y_c_403_n 0.00300916f $X=4.555 $Y=1.41 $X2=0 $Y2=0
cc_182 N_B1_c_211_n N_Y_c_403_n 7.29089e-19 $X=4.005 $Y=1.202 $X2=0 $Y2=0
cc_183 B1 N_Y_c_403_n 0.0108421f $X=4.73 $Y=1.445 $X2=0 $Y2=0
cc_184 N_B1_c_213_n N_Y_c_403_n 3.20002e-19 $X=4.555 $Y=1.202 $X2=0 $Y2=0
cc_185 N_B1_c_228_p N_Y_c_403_n 0.0214558f $X=4.715 $Y=1.175 $X2=0 $Y2=0
cc_186 N_B1_c_208_n N_Y_c_427_n 0.015503f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_187 N_B1_c_209_n N_Y_c_427_n 0.0055165f $X=4.455 $Y=1.16 $X2=0 $Y2=0
cc_188 N_B1_c_210_n N_Y_c_427_n 0.0104224f $X=4.53 $Y=0.995 $X2=0 $Y2=0
cc_189 N_B1_c_228_p N_Y_c_427_n 0.0181676f $X=4.715 $Y=1.175 $X2=0 $Y2=0
cc_190 N_B1_c_214_n N_Y_c_431_n 0.00836442f $X=4.005 $Y=1.41 $X2=0 $Y2=0
cc_191 N_B1_c_216_n N_Y_c_431_n 0.0118164f $X=4.555 $Y=1.41 $X2=0 $Y2=0
cc_192 B1 N_Y_c_431_n 5.68138e-19 $X=4.73 $Y=1.445 $X2=0 $Y2=0
cc_193 N_B1_c_208_n N_Y_c_401_n 7.05755e-19 $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_194 N_B1_c_210_n N_Y_c_401_n 0.00760167f $X=4.53 $Y=0.995 $X2=0 $Y2=0
cc_195 B1 N_Y_c_401_n 0.0151122f $X=4.73 $Y=1.105 $X2=0 $Y2=0
cc_196 N_B1_c_213_n N_Y_c_401_n 0.00819476f $X=4.555 $Y=1.202 $X2=0 $Y2=0
cc_197 N_B1_c_228_p N_Y_c_401_n 0.00651646f $X=4.715 $Y=1.175 $X2=0 $Y2=0
cc_198 N_B1_c_208_n Y 0.0103672f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_199 N_B1_c_214_n Y 7.38675e-19 $X=4.005 $Y=1.41 $X2=0 $Y2=0
cc_200 N_B1_c_228_p Y 0.00656374f $X=4.715 $Y=1.175 $X2=0 $Y2=0
cc_201 N_B1_c_208_n N_VGND_c_497_n 0.00858015f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_202 N_B1_c_210_n N_VGND_c_497_n 0.00443041f $X=4.53 $Y=0.995 $X2=0 $Y2=0
cc_203 N_B1_c_208_n N_VGND_c_498_n 0.00342417f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_204 N_B1_c_210_n N_VGND_c_500_n 0.00417062f $X=4.53 $Y=0.995 $X2=0 $Y2=0
cc_205 N_B1_c_208_n N_VGND_c_501_n 0.00426775f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_206 N_B1_c_210_n N_VGND_c_501_n 0.00695019f $X=4.53 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A_27_297#_c_263_n N_VPWR_M1001_s 0.00347905f $X=1.115 $Y=1.87 $X2=0.495
+ $Y2=1.41
cc_208 N_A_27_297#_c_270_n N_VPWR_M1011_s 0.00347905f $X=2.055 $Y=1.87 $X2=0.495
+ $Y2=1.985
cc_209 N_A_27_297#_c_275_n N_VPWR_M1007_s 0.021908f $X=3.685 $Y=1.87 $X2=0.495
+ $Y2=1.985
cc_210 N_A_27_297#_c_263_n N_VPWR_c_330_n 0.0203395f $X=1.115 $Y=1.87 $X2=0.99
+ $Y2=0.56
cc_211 N_A_27_297#_c_267_n N_VPWR_c_330_n 0.0253827f $X=0.26 $Y=1.95 $X2=0.99
+ $Y2=0.56
cc_212 N_A_27_297#_c_274_n N_VPWR_c_330_n 0.0208108f $X=1.2 $Y=1.95 $X2=0.99
+ $Y2=0.56
cc_213 N_A_27_297#_c_270_n N_VPWR_c_331_n 0.0203395f $X=2.055 $Y=1.87 $X2=0
+ $Y2=0
cc_214 N_A_27_297#_c_274_n N_VPWR_c_331_n 0.0253827f $X=1.2 $Y=1.95 $X2=0 $Y2=0
cc_215 N_A_27_297#_c_296_p N_VPWR_c_331_n 0.0208108f $X=2.14 $Y=1.95 $X2=0 $Y2=0
cc_216 N_A_27_297#_c_267_n N_VPWR_c_332_n 0.0118139f $X=0.26 $Y=1.95 $X2=0 $Y2=0
cc_217 N_A_27_297#_c_274_n N_VPWR_c_333_n 0.0118139f $X=1.2 $Y=1.95 $X2=0.605
+ $Y2=1.16
cc_218 N_A_27_297#_c_283_n N_VPWR_c_334_n 0.0585163f $X=4.705 $Y=2.38 $X2=0
+ $Y2=0
cc_219 N_A_27_297#_c_281_n N_VPWR_c_334_n 0.0119545f $X=3.855 $Y=2.38 $X2=0
+ $Y2=0
cc_220 N_A_27_297#_M1001_d N_VPWR_c_329_n 0.00391905f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_221 N_A_27_297#_M1006_d N_VPWR_c_329_n 0.00295369f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_222 N_A_27_297#_M1015_d N_VPWR_c_329_n 0.00295369f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_223 N_A_27_297#_M1009_d N_VPWR_c_329_n 0.00387873f $X=3.535 $Y=1.485 $X2=0
+ $Y2=0
cc_224 N_A_27_297#_M1010_s N_VPWR_c_329_n 0.00356385f $X=4.645 $Y=1.485 $X2=0
+ $Y2=0
cc_225 N_A_27_297#_c_263_n N_VPWR_c_329_n 0.0134894f $X=1.115 $Y=1.87 $X2=0
+ $Y2=0
cc_226 N_A_27_297#_c_270_n N_VPWR_c_329_n 0.0134894f $X=2.055 $Y=1.87 $X2=0
+ $Y2=0
cc_227 N_A_27_297#_c_275_n N_VPWR_c_329_n 0.0269697f $X=3.685 $Y=1.87 $X2=0
+ $Y2=0
cc_228 N_A_27_297#_c_283_n N_VPWR_c_329_n 0.0364022f $X=4.705 $Y=2.38 $X2=0
+ $Y2=0
cc_229 N_A_27_297#_c_281_n N_VPWR_c_329_n 0.006547f $X=3.855 $Y=2.38 $X2=0 $Y2=0
cc_230 N_A_27_297#_c_267_n N_VPWR_c_329_n 0.00646998f $X=0.26 $Y=1.95 $X2=0
+ $Y2=0
cc_231 N_A_27_297#_c_274_n N_VPWR_c_329_n 0.00646998f $X=1.2 $Y=1.95 $X2=0 $Y2=0
cc_232 N_A_27_297#_c_296_p N_VPWR_c_329_n 0.00646998f $X=2.14 $Y=1.95 $X2=0
+ $Y2=0
cc_233 N_A_27_297#_c_296_p N_VPWR_c_338_n 0.0118139f $X=2.14 $Y=1.95 $X2=0 $Y2=0
cc_234 N_A_27_297#_c_275_n N_VPWR_c_339_n 0.0566177f $X=3.685 $Y=1.87 $X2=0
+ $Y2=0
cc_235 N_A_27_297#_c_280_n N_VPWR_c_339_n 0.00723947f $X=3.77 $Y=2.295 $X2=0
+ $Y2=0
cc_236 N_A_27_297#_c_281_n N_VPWR_c_339_n 0.00806765f $X=3.855 $Y=2.38 $X2=0
+ $Y2=0
cc_237 N_A_27_297#_c_296_p N_VPWR_c_339_n 0.0167779f $X=2.14 $Y=1.95 $X2=0 $Y2=0
cc_238 N_A_27_297#_c_283_n N_Y_M1008_d 0.00524122f $X=4.705 $Y=2.38 $X2=0.52
+ $Y2=0.995
cc_239 N_A_27_297#_M1009_d N_Y_c_403_n 0.00230741f $X=3.535 $Y=1.485 $X2=0.495
+ $Y2=1.202
cc_240 N_A_27_297#_c_275_n N_Y_c_403_n 0.0028327f $X=3.685 $Y=1.87 $X2=0.495
+ $Y2=1.202
cc_241 N_A_27_297#_c_322_p N_Y_c_403_n 0.013831f $X=3.77 $Y=1.955 $X2=0.495
+ $Y2=1.202
cc_242 N_A_27_297#_c_322_p N_Y_c_431_n 0.0095104f $X=3.77 $Y=1.955 $X2=0.99
+ $Y2=1.202
cc_243 N_A_27_297#_c_280_n N_Y_c_431_n 0.00802388f $X=3.77 $Y=2.295 $X2=0.99
+ $Y2=1.202
cc_244 N_A_27_297#_c_283_n N_Y_c_431_n 0.0195098f $X=4.705 $Y=2.38 $X2=0.99
+ $Y2=1.202
cc_245 N_A_27_297#_c_285_n N_Y_c_431_n 0.0193734f $X=4.79 $Y=1.96 $X2=0.99
+ $Y2=1.202
cc_246 N_A_27_297#_M1009_d Y 5.87954e-19 $X=3.535 $Y=1.485 $X2=0.745 $Y2=1.305
cc_247 N_A_27_297#_c_275_n Y 0.0180236f $X=3.685 $Y=1.87 $X2=0.745 $Y2=1.305
cc_248 N_VPWR_c_329_n N_Y_M1008_d 0.00297142f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_249 N_Y_c_400_n N_A_27_47#_c_475_n 0.0123435f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_250 N_Y_c_427_n N_VGND_M1003_d 0.00687004f $X=4.575 $Y=0.75 $X2=0 $Y2=0
cc_251 N_Y_c_419_n N_VGND_c_497_n 0.0116547f $X=3.69 $Y=0.42 $X2=0 $Y2=0
cc_252 N_Y_c_427_n N_VGND_c_497_n 0.0218854f $X=4.575 $Y=0.75 $X2=0 $Y2=0
cc_253 N_Y_c_419_n N_VGND_c_498_n 0.0117202f $X=3.69 $Y=0.42 $X2=0 $Y2=0
cc_254 N_Y_c_427_n N_VGND_c_498_n 0.00364243f $X=4.575 $Y=0.75 $X2=0 $Y2=0
cc_255 Y N_VGND_c_498_n 0.00333995f $X=3.435 $Y=0.765 $X2=0 $Y2=0
cc_256 N_Y_c_427_n N_VGND_c_500_n 0.00235272f $X=4.575 $Y=0.75 $X2=0 $Y2=0
cc_257 N_Y_c_401_n N_VGND_c_500_n 0.0192822f $X=4.79 $Y=0.38 $X2=0 $Y2=0
cc_258 N_Y_M1000_d N_VGND_c_501_n 0.00253905f $X=2.585 $Y=0.235 $X2=0 $Y2=0
cc_259 N_Y_M1004_d N_VGND_c_501_n 0.00361011f $X=3.545 $Y=0.235 $X2=0 $Y2=0
cc_260 N_Y_M1014_s N_VGND_c_501_n 0.00252987f $X=4.605 $Y=0.235 $X2=0 $Y2=0
cc_261 N_Y_c_419_n N_VGND_c_501_n 0.00645161f $X=3.69 $Y=0.42 $X2=0 $Y2=0
cc_262 N_Y_c_427_n N_VGND_c_501_n 0.0122934f $X=4.575 $Y=0.75 $X2=0 $Y2=0
cc_263 N_Y_c_401_n N_VGND_c_501_n 0.0139745f $X=4.79 $Y=0.38 $X2=0 $Y2=0
cc_264 Y N_VGND_c_501_n 0.00607689f $X=3.435 $Y=0.765 $X2=0 $Y2=0
cc_265 N_Y_c_400_n N_A_297_47#_M1000_s 0.0065896f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_266 Y N_A_297_47#_M1000_s 3.89508e-19 $X=3.435 $Y=0.765 $X2=0 $Y2=0
cc_267 Y N_A_297_47#_M1000_s 5.33276e-19 $X=3.515 $Y=0.85 $X2=0 $Y2=0
cc_268 N_Y_M1000_d N_A_297_47#_c_551_n 0.00632442f $X=2.585 $Y=0.235 $X2=0 $Y2=0
cc_269 N_Y_c_400_n N_A_297_47#_c_551_n 0.0414707f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_270 Y N_A_297_47#_c_551_n 5.59064e-19 $X=3.435 $Y=0.765 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_475_n N_VGND_M1002_s 0.00408716f $X=2.14 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_272 N_A_27_47#_c_475_n N_VGND_c_498_n 0.00806484f $X=2.14 $Y=0.74 $X2=0 $Y2=0
cc_273 N_A_27_47#_c_475_n N_VGND_c_499_n 0.00655693f $X=2.14 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A_27_47#_M1002_d N_VGND_c_501_n 0.00375731f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_M1012_d N_VGND_c_501_n 0.00323135f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_M1013_s N_VGND_c_501_n 0.00212464f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_475_n N_VGND_c_501_n 0.0289625f $X=2.14 $Y=0.74 $X2=0 $Y2=0
cc_278 N_A_27_47#_c_475_n N_VGND_c_502_n 0.0193991f $X=2.14 $Y=0.74 $X2=0 $Y2=0
cc_279 N_A_27_47#_c_475_n N_A_297_47#_M1005_d 0.00513712f $X=2.14 $Y=0.74
+ $X2=-0.19 $Y2=-0.24
cc_280 N_A_27_47#_M1013_s N_A_297_47#_c_551_n 0.00508809f $X=2.005 $Y=0.235
+ $X2=0 $Y2=0
cc_281 N_A_27_47#_c_475_n N_A_297_47#_c_551_n 0.0418342f $X=2.14 $Y=0.74 $X2=0
+ $Y2=0
cc_282 N_VGND_c_501_n N_A_297_47#_M1005_d 0.00298815f $X=4.83 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_283 N_VGND_c_501_n N_A_297_47#_M1000_s 0.00289859f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_284 N_VGND_c_498_n N_A_297_47#_c_551_n 0.0897105f $X=4.025 $Y=0 $X2=0 $Y2=0
cc_285 N_VGND_c_501_n N_A_297_47#_c_551_n 0.0680333f $X=4.83 $Y=0 $X2=0 $Y2=0
