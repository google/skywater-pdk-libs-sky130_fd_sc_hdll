* File: sky130_fd_sc_hdll__o31ai_1.spice
* Created: Thu Aug 27 19:22:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o31ai_1.pex.spice"
.subckt sky130_fd_sc_hdll__o31ai_1  VNB VPB A1 A2 A3 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1005 N_A_119_47#_M1005_d N_A1_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.2015 PD=0.98 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g N_A_119_47#_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.10725 PD=0.92 PS=0.98 NRD=0 NRS=10.152 M=1 R=4.33333
+ SA=75000.7 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1004 N_A_119_47#_M1004_d N_A3_M1004_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.15925 AS=0.08775 PD=1.14 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_B1_M1002_g N_A_119_47#_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2535 AS=0.15925 PD=2.08 PS=1.14 NRD=10.152 NRS=39.684 M=1 R=4.33333
+ SA=75001.8 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1000 A_117_297# N_A1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.27 PD=1.3 PS=2.54 NRD=18.6953 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90001.9 A=0.18 P=2.36 MULT=1
MM1006 A_213_297# N_A2_M1006_g A_117_297# VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.15 PD=1.29 PS=1.3 NRD=17.7103 NRS=18.6953 M=1 R=5.55556 SA=90000.7
+ SB=90001.4 A=0.18 P=2.36 MULT=1
MM1003 N_Y_M1003_d N_A3_M1003_g A_213_297# VPB PHIGHVT L=0.18 W=1 AD=0.29
+ AS=0.145 PD=1.58 PS=1.29 NRD=58.0953 NRS=17.7103 M=1 R=5.55556 SA=90001.1
+ SB=90000.9 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_B1_M1007_g N_Y_M1003_d VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.29 PD=2.54 PS=1.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.9
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hdll__o31ai_1.pxi.spice"
*
.ends
*
*
