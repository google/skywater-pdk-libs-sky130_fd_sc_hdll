* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__and3b_4 A_N B C VGND VNB VPB VPWR X
X0 VPWR B a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 X a_56_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 X a_56_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_56_297# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 VGND a_56_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR a_56_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 X a_56_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_56_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 a_56_297# a_98_199# a_162_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_162_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND a_56_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR a_56_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 VPWR A_N a_98_199# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X14 a_56_297# a_98_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 VGND A_N a_98_199# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
