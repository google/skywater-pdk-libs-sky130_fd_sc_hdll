* File: sky130_fd_sc_hdll__a221oi_2.pex.spice
* Created: Wed Sep  2 08:18:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A221OI_2%C1 1 3 4 6 7 9 10 12 13 14 22
r40 22 23 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.975 $Y=1.202
+ $X2=1 $Y2=1.202
r41 21 22 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=0.53 $Y=1.202
+ $X2=0.975 $Y2=1.202
r42 20 21 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.505 $Y=1.202
+ $X2=0.53 $Y2=1.202
r43 18 20 33.0137 $w=3.65e-07 $l=2.5e-07 $layer=POLY_cond $X=0.255 $Y=1.202
+ $X2=0.505 $Y2=1.202
r44 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.16
+ $X2=0.255 $Y2=1.53
r45 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.255
+ $Y=1.16 $X2=0.255 $Y2=1.16
r46 10 23 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1 $Y=0.995 $X2=1
+ $Y2=1.202
r47 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1 $Y=0.995 $X2=1
+ $Y2=0.56
r48 7 22 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.975 $Y=1.41
+ $X2=0.975 $Y2=1.202
r49 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.975 $Y=1.41
+ $X2=0.975 $Y2=1.985
r50 4 21 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.53 $Y=0.995
+ $X2=0.53 $Y2=1.202
r51 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.53 $Y=0.995 $X2=0.53
+ $Y2=0.56
r52 1 20 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.41
+ $X2=0.505 $Y2=1.202
r53 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.41
+ $X2=0.505 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_2%B2 1 3 4 6 7 9 10 12 13 16 21 22
c77 7 0 1.81434e-19 $X=3.375 $Y=1.41
c78 1 0 1.39491e-19 $X=1.965 $Y=1.41
r79 21 22 9.62063 $w=4.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.96 $Y=1.16
+ $X2=1.96 $Y2=1.53
r80 21 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.94
+ $Y=1.16 $X2=1.94 $Y2=1.16
r81 16 19 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.375 $Y=1.16
+ $X2=3.375 $Y2=1.53
r82 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.35
+ $Y=1.16 $X2=3.35 $Y2=1.16
r83 14 22 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.19 $Y=1.53 $X2=1.96
+ $Y2=1.53
r84 13 19 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.185 $Y=1.53
+ $X2=3.375 $Y2=1.53
r85 13 14 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=3.185 $Y=1.53
+ $X2=2.19 $Y2=1.53
r86 10 17 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=3.4 $Y=0.995
+ $X2=3.375 $Y2=1.16
r87 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.4 $Y=0.995 $X2=3.4
+ $Y2=0.56
r88 7 17 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=3.375 $Y=1.41
+ $X2=3.375 $Y2=1.16
r89 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.375 $Y=1.41
+ $X2=3.375 $Y2=1.985
r90 4 26 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.99 $Y=0.995
+ $X2=1.965 $Y2=1.16
r91 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.99 $Y=0.995 $X2=1.99
+ $Y2=0.56
r92 1 26 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=1.965 $Y=1.41
+ $X2=1.965 $Y2=1.16
r93 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.965 $Y=1.41
+ $X2=1.965 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_2%B1 1 3 4 6 7 9 10 12 13 20 23
r44 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=2.905 $Y=1.202
+ $X2=2.93 $Y2=1.202
r45 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=2.67 $Y=1.202
+ $X2=2.905 $Y2=1.202
r46 16 18 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=2.435 $Y=1.202
+ $X2=2.67 $Y2=1.202
r47 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=2.41 $Y=1.202
+ $X2=2.435 $Y2=1.202
r48 13 23 6.37727 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=2.67 $Y=1.175
+ $X2=2.555 $Y2=1.175
r49 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.16 $X2=2.67 $Y2=1.16
r50 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.93 $Y=0.995
+ $X2=2.93 $Y2=1.202
r51 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.93 $Y=0.995
+ $X2=2.93 $Y2=0.56
r52 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.905 $Y=1.41
+ $X2=2.905 $Y2=1.202
r53 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.905 $Y=1.41
+ $X2=2.905 $Y2=1.985
r54 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.435 $Y=1.41
+ $X2=2.435 $Y2=1.202
r55 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.435 $Y=1.41
+ $X2=2.435 $Y2=1.985
r56 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.41 $Y=0.995
+ $X2=2.41 $Y2=1.202
r57 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.41 $Y=0.995 $X2=2.41
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_2%A2 1 3 4 6 7 9 10 12 15 18 19 21 22 23 30
c77 10 0 1.80188e-19 $X=5.36 $Y=0.995
c78 7 0 1.96071e-19 $X=5.335 $Y=1.41
c79 1 0 4.1943e-20 $X=3.925 $Y=1.41
r80 27 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.31
+ $Y=1.16 $X2=5.31 $Y2=1.16
r81 23 30 24.1227 $w=1.98e-07 $l=4.35e-07 $layer=LI1_cond $X=5.725 $Y=1.175
+ $X2=5.29 $Y2=1.175
r82 22 30 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=5.27 $Y=1.175 $X2=5.29
+ $Y2=1.175
r83 20 22 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.185 $Y=1.275
+ $X2=5.27 $Y2=1.175
r84 20 21 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.185 $Y=1.275
+ $X2=5.185 $Y2=1.445
r85 18 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.1 $Y=1.53
+ $X2=5.185 $Y2=1.445
r86 18 19 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=5.1 $Y=1.53
+ $X2=4.065 $Y2=1.53
r87 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.9
+ $Y=1.16 $X2=3.9 $Y2=1.16
r88 13 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.9 $Y=1.445
+ $X2=4.065 $Y2=1.53
r89 13 15 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.9 $Y=1.445
+ $X2=3.9 $Y2=1.16
r90 10 27 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=5.36 $Y=0.995
+ $X2=5.335 $Y2=1.16
r91 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.36 $Y=0.995
+ $X2=5.36 $Y2=0.56
r92 7 27 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=5.335 $Y=1.41
+ $X2=5.335 $Y2=1.16
r93 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.335 $Y=1.41
+ $X2=5.335 $Y2=1.985
r94 4 16 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=3.95 $Y=0.995
+ $X2=3.925 $Y2=1.16
r95 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.95 $Y=0.995 $X2=3.95
+ $Y2=0.56
r96 1 16 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=3.925 $Y=1.41
+ $X2=3.925 $Y2=1.16
r97 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.925 $Y=1.41
+ $X2=3.925 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_2%A1 1 3 4 6 7 9 10 12 13 20 24
c45 13 0 1.96071e-19 $X=4.725 $Y=1.105
c46 10 0 1.86655e-19 $X=4.89 $Y=0.995
r47 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.865 $Y=1.202
+ $X2=4.89 $Y2=1.202
r48 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=4.63 $Y=1.202
+ $X2=4.865 $Y2=1.202
r49 18 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.63
+ $Y=1.16 $X2=4.63 $Y2=1.16
r50 16 18 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=4.395 $Y=1.202
+ $X2=4.63 $Y2=1.202
r51 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.37 $Y=1.202
+ $X2=4.395 $Y2=1.202
r52 13 24 9.98182 $w=1.98e-07 $l=1.8e-07 $layer=LI1_cond $X=4.81 $Y=1.175
+ $X2=4.63 $Y2=1.175
r53 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.89 $Y=0.995
+ $X2=4.89 $Y2=1.202
r54 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.89 $Y=0.995
+ $X2=4.89 $Y2=0.56
r55 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.865 $Y=1.41
+ $X2=4.865 $Y2=1.202
r56 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.865 $Y=1.41
+ $X2=4.865 $Y2=1.985
r57 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.395 $Y=1.41
+ $X2=4.395 $Y2=1.202
r58 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.395 $Y=1.41
+ $X2=4.395 $Y2=1.985
r59 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.37 $Y=0.995
+ $X2=4.37 $Y2=1.202
r60 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.37 $Y=0.995 $X2=4.37
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_2%A_27_297# 1 2 3 4 15 17 18 21 24 25 27 29
+ 30 35
c62 35 0 1.39491e-19 $X=3.14 $Y=1.87
c63 30 0 1.39491e-19 $X=2.2 $Y=1.87
r64 35 38 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=3.14 $Y=1.87 $X2=3.14
+ $Y2=1.96
r65 30 33 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.2 $Y=1.87 $X2=2.2
+ $Y2=1.96
r66 28 30 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.325 $Y=1.87
+ $X2=2.2 $Y2=1.87
r67 27 35 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.015 $Y=1.87
+ $X2=3.14 $Y2=1.87
r68 27 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.015 $Y=1.87
+ $X2=2.325 $Y2=1.87
r69 26 29 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.375 $Y=1.87
+ $X2=1.25 $Y2=1.87
r70 25 30 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.075 $Y=1.87
+ $X2=2.2 $Y2=1.87
r71 25 26 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.075 $Y=1.87
+ $X2=1.375 $Y2=1.87
r72 23 29 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=1.955
+ $X2=1.25 $Y2=1.87
r73 23 24 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=1.25 $Y=1.955
+ $X2=1.25 $Y2=2.295
r74 19 29 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=1.785
+ $X2=1.25 $Y2=1.87
r75 19 21 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.25 $Y=1.785
+ $X2=1.25 $Y2=1.66
r76 17 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.125 $Y=2.38
+ $X2=1.25 $Y2=2.295
r77 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.125 $Y=2.38
+ $X2=0.435 $Y2=2.38
r78 13 18 7.89393 $w=1.7e-07 $l=2.11268e-07 $layer=LI1_cond $X=0.262 $Y=2.295
+ $X2=0.435 $Y2=2.38
r79 13 15 13.8627 $w=3.43e-07 $l=4.15e-07 $layer=LI1_cond $X=0.262 $Y=2.295
+ $X2=0.262 $Y2=1.88
r80 4 38 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=2.995
+ $Y=1.485 $X2=3.14 $Y2=1.96
r81 3 33 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=2.055
+ $Y=1.485 $X2=2.2 $Y2=1.96
r82 2 21 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=1.065
+ $Y=1.485 $X2=1.21 $Y2=1.66
r83 1 15 300 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.27 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_2%Y 1 2 3 4 15 16 21 22 24 25 27 28 29 30
+ 31 40
r74 31 49 9.60369 $w=2.98e-07 $l=2.5e-07 $layer=LI1_cond $X=0.755 $Y=1.87
+ $X2=0.755 $Y2=1.62
r75 30 49 3.45733 $w=2.98e-07 $l=9e-08 $layer=LI1_cond $X=0.755 $Y=1.53
+ $X2=0.755 $Y2=1.62
r76 29 30 13.061 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.755 $Y=1.19
+ $X2=0.755 $Y2=1.53
r77 28 38 2.9604 $w=3.4e-07 $l=1.9e-07 $layer=LI1_cond $X=0.525 $Y=0.725
+ $X2=0.715 $Y2=0.725
r78 28 43 2.9604 $w=3.4e-07 $l=3.07083e-07 $layer=LI1_cond $X=0.525 $Y=0.725
+ $X2=0.755 $Y2=0.905
r79 28 29 10.372 $w=2.98e-07 $l=2.7e-07 $layer=LI1_cond $X=0.755 $Y=0.92
+ $X2=0.755 $Y2=1.19
r80 28 43 0.576222 $w=2.98e-07 $l=1.5e-08 $layer=LI1_cond $X=0.755 $Y=0.92
+ $X2=0.755 $Y2=0.905
r81 27 38 6.5204 $w=3.78e-07 $l=2.15e-07 $layer=LI1_cond $X=0.715 $Y=0.51
+ $X2=0.715 $Y2=0.725
r82 27 40 3.63929 $w=3.78e-07 $l=1.2e-07 $layer=LI1_cond $X=0.715 $Y=0.51
+ $X2=0.715 $Y2=0.39
r83 24 25 10.6316 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=4.63 $Y=0.775
+ $X2=4.415 $Y2=0.775
r84 22 25 97.3535 $w=1.78e-07 $l=1.58e-06 $layer=LI1_cond $X=2.835 $Y=0.815
+ $X2=4.415 $Y2=0.815
r85 16 21 6.86404 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=2.565 $Y=0.775
+ $X2=2.435 $Y2=0.775
r86 16 18 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=2.565 $Y=0.775
+ $X2=2.67 $Y2=0.775
r87 15 22 6.86404 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=2.705 $Y=0.775
+ $X2=2.835 $Y2=0.775
r88 15 18 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=2.705 $Y=0.775
+ $X2=2.67 $Y2=0.775
r89 14 28 3.70584 $w=1.8e-07 $l=4.22611e-07 $layer=LI1_cond $X=0.905 $Y=0.815
+ $X2=0.525 $Y2=0.725
r90 14 21 94.2727 $w=1.78e-07 $l=1.53e-06 $layer=LI1_cond $X=0.905 $Y=0.815
+ $X2=2.435 $Y2=0.815
r91 4 49 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.485 $X2=0.74 $Y2=1.62
r92 3 24 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=4.445
+ $Y=0.235 $X2=4.63 $Y2=0.73
r93 2 18 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.235 $X2=2.67 $Y2=0.73
r94 1 40 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.605
+ $Y=0.235 $X2=0.74 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_2%A_321_297# 1 2 3 4 5 16 18 20 22 26 28 32
+ 36 39 44 50
c60 20 0 8.3886e-20 $X=3.65 $Y=1.955
r61 44 46 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.67 $Y=2.3 $X2=2.67
+ $Y2=2.38
r62 39 41 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=1.73 $Y=2.3 $X2=1.73
+ $Y2=2.38
r63 34 51 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.592 $Y=1.955
+ $X2=5.592 $Y2=1.87
r64 34 36 0.27051 $w=2.03e-07 $l=5e-09 $layer=LI1_cond $X=5.592 $Y=1.955
+ $X2=5.592 $Y2=1.96
r65 30 51 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.592 $Y=1.785
+ $X2=5.592 $Y2=1.87
r66 30 32 8.92683 $w=2.03e-07 $l=1.65e-07 $layer=LI1_cond $X=5.592 $Y=1.785
+ $X2=5.592 $Y2=1.62
r67 29 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.755 $Y=1.87
+ $X2=4.63 $Y2=1.87
r68 28 51 2.0246 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=5.49 $Y=1.87
+ $X2=5.592 $Y2=1.87
r69 28 29 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=5.49 $Y=1.87
+ $X2=4.755 $Y2=1.87
r70 24 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.63 $Y=1.955
+ $X2=4.63 $Y2=1.87
r71 24 26 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=4.63 $Y=1.955
+ $X2=4.63 $Y2=1.96
r72 23 49 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.775 $Y=1.87
+ $X2=3.65 $Y2=1.87
r73 22 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.505 $Y=1.87
+ $X2=4.63 $Y2=1.87
r74 22 23 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.505 $Y=1.87
+ $X2=3.775 $Y2=1.87
r75 20 49 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.65 $Y=1.955
+ $X2=3.65 $Y2=1.87
r76 20 21 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=3.65 $Y=1.955
+ $X2=3.65 $Y2=2.295
r77 19 46 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.795 $Y=2.38
+ $X2=2.67 $Y2=2.38
r78 18 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.525 $Y=2.38
+ $X2=3.65 $Y2=2.295
r79 18 19 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.525 $Y=2.38
+ $X2=2.795 $Y2=2.38
r80 17 41 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.855 $Y=2.38
+ $X2=1.73 $Y2=2.38
r81 16 46 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.545 $Y=2.38
+ $X2=2.67 $Y2=2.38
r82 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.545 $Y=2.38
+ $X2=1.855 $Y2=2.38
r83 5 36 300 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=2 $X=5.425
+ $Y=1.485 $X2=5.575 $Y2=1.96
r84 5 32 600 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=1 $X=5.425
+ $Y=1.485 $X2=5.575 $Y2=1.62
r85 4 26 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.485
+ $Y=1.485 $X2=4.63 $Y2=1.96
r86 3 49 300 $w=1.7e-07 $l=5.49773e-07 $layer=licon1_PDIFF $count=2 $X=3.465
+ $Y=1.485 $X2=3.65 $Y2=1.95
r87 2 44 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=1.485 $X2=2.67 $Y2=2.3
r88 1 39 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=1.605
+ $Y=1.485 $X2=1.73 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_2%VPWR 1 2 9 13 16 17 19 20 21 34 35
r69 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r70 32 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r71 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r72 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r73 28 29 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r74 24 28 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=3.91 $Y2=2.72
r75 21 29 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=3.91 $Y2=2.72
r76 21 24 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r77 19 31 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.975 $Y=2.72
+ $X2=4.83 $Y2=2.72
r78 19 20 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.975 $Y=2.72
+ $X2=5.1 $Y2=2.72
r79 18 34 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=5.225 $Y=2.72
+ $X2=5.75 $Y2=2.72
r80 18 20 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.225 $Y=2.72
+ $X2=5.1 $Y2=2.72
r81 16 28 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.035 $Y=2.72
+ $X2=3.91 $Y2=2.72
r82 16 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.035 $Y=2.72
+ $X2=4.16 $Y2=2.72
r83 15 31 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=4.285 $Y=2.72
+ $X2=4.83 $Y2=2.72
r84 15 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.285 $Y=2.72
+ $X2=4.16 $Y2=2.72
r85 11 20 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.1 $Y=2.635
+ $X2=5.1 $Y2=2.72
r86 11 13 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.1 $Y=2.635
+ $X2=5.1 $Y2=2.3
r87 7 17 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.16 $Y=2.635
+ $X2=4.16 $Y2=2.72
r88 7 9 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.16 $Y=2.635
+ $X2=4.16 $Y2=2.3
r89 2 13 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.955
+ $Y=1.485 $X2=5.1 $Y2=2.3
r90 1 9 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.015
+ $Y=1.485 $X2=4.16 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_2%VGND 1 2 3 4 13 15 21 25 28 29 31 32 33
+ 49 50 58 64
r72 63 64 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=0.235
+ $X2=1.815 $Y2=0.235
r73 60 63 2.24265 $w=6.38e-07 $l=1.2e-07 $layer=LI1_cond $X=1.61 $Y=0.235
+ $X2=1.73 $Y2=0.235
r74 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r75 57 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r76 56 60 8.59681 $w=6.38e-07 $l=4.6e-07 $layer=LI1_cond $X=1.15 $Y=0.235
+ $X2=1.61 $Y2=0.235
r77 56 58 7.80044 $w=6.38e-07 $l=2.5e-08 $layer=LI1_cond $X=1.15 $Y=0.235
+ $X2=1.125 $Y2=0.235
r78 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r79 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r80 47 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r81 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r82 44 47 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=0 $X2=5.29
+ $Y2=0
r83 43 46 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=5.29
+ $Y2=0
r84 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r85 41 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r86 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r87 38 41 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r88 38 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r89 37 40 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r90 37 64 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.815
+ $Y2=0
r91 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r92 33 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r93 33 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r94 31 46 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.485 $Y=0 $X2=5.29
+ $Y2=0
r95 31 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.485 $Y=0 $X2=5.57
+ $Y2=0
r96 30 49 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=5.655 $Y=0 $X2=5.75
+ $Y2=0
r97 30 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.655 $Y=0 $X2=5.57
+ $Y2=0
r98 28 40 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.45
+ $Y2=0
r99 28 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.655
+ $Y2=0
r100 27 43 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.91
+ $Y2=0
r101 27 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.655
+ $Y2=0
r102 23 32 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=0.085
+ $X2=5.57 $Y2=0
r103 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.57 $Y=0.085
+ $X2=5.57 $Y2=0.39
r104 19 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=0.085
+ $X2=3.655 $Y2=0
r105 19 21 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.655 $Y=0.085
+ $X2=3.655 $Y2=0.39
r106 18 53 4.02368 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=0
+ $X2=0.177 $Y2=0
r107 18 58 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.355 $Y=0
+ $X2=1.125 $Y2=0
r108 13 53 3.11948 $w=2.5e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.23 $Y=0.085
+ $X2=0.177 $Y2=0
r109 13 15 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.23 $Y=0.085
+ $X2=0.23 $Y2=0.39
r110 4 25 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.435
+ $Y=0.235 $X2=5.57 $Y2=0.39
r111 3 21 182 $w=1.7e-07 $l=2.45561e-07 $layer=licon1_NDIFF $count=1 $X=3.475
+ $Y=0.235 $X2=3.655 $Y2=0.39
r112 2 63 91 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_NDIFF $count=2 $X=1.075
+ $Y=0.235 $X2=1.73 $Y2=0.39
r113 1 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.27 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_2%A_413_47# 1 2 11
r14 8 11 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=2.2 $Y=0.365 $X2=3.14
+ $Y2=0.365
r15 2 11 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.005
+ $Y=0.235 $X2=3.14 $Y2=0.39
r16 1 8 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.065
+ $Y=0.235 $X2=2.2 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_2%A_805_47# 1 2 7 11 13
c21 13 0 3.66843e-19 $X=5.1 $Y=0.73
r22 11 16 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=5.14 $Y=0.475
+ $X2=5.14 $Y2=0.365
r23 11 13 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=5.14 $Y=0.475
+ $X2=5.14 $Y2=0.73
r24 7 16 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=5.015 $Y=0.365
+ $X2=5.14 $Y2=0.365
r25 7 9 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=5.015 $Y=0.365
+ $X2=4.16 $Y2=0.365
r26 2 16 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.965
+ $Y=0.235 $X2=5.1 $Y2=0.39
r27 2 13 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.965
+ $Y=0.235 $X2=5.1 $Y2=0.73
r28 1 9 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.025
+ $Y=0.235 $X2=4.16 $Y2=0.39
.ends

