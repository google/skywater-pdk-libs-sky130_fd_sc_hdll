* File: sky130_fd_sc_hdll__muxb4to1_1.pxi.spice
* Created: Thu Aug 27 19:11:45 2020
* 
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%D[0] N_D[0]_c_140_n N_D[0]_M1021_g
+ N_D[0]_c_141_n N_D[0]_M1007_g N_D[0]_c_142_n N_D[0]_c_143_n D[0]
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%D[0]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%A_184_265# N_A_184_265#_M1017_s
+ N_A_184_265#_M1013_s N_A_184_265#_M1009_g N_A_184_265#_c_168_n
+ N_A_184_265#_c_169_n N_A_184_265#_c_173_n N_A_184_265#_c_170_n
+ N_A_184_265#_c_171_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%A_184_265#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%S[0] N_S[0]_c_224_n N_S[0]_M1023_g
+ N_S[0]_c_225_n N_S[0]_c_226_n N_S[0]_c_227_n N_S[0]_M1013_g N_S[0]_c_228_n
+ N_S[0]_M1017_g S[0] N_S[0]_c_229_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%S[0]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%S[1] N_S[1]_c_270_n N_S[1]_M1010_g
+ N_S[1]_c_271_n N_S[1]_M1016_g N_S[1]_c_272_n N_S[1]_c_273_n N_S[1]_M1006_g
+ S[1] N_S[1]_c_274_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%S[1]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%A_533_47# N_A_533_47#_M1016_d
+ N_A_533_47#_M1010_d N_A_533_47#_M1003_g N_A_533_47#_c_319_n
+ N_A_533_47#_c_314_n N_A_533_47#_c_315_n N_A_533_47#_c_316_n
+ N_A_533_47#_c_317_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%A_533_47#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%D[1] N_D[1]_c_369_n N_D[1]_M1019_g
+ N_D[1]_c_370_n N_D[1]_M1018_g N_D[1]_c_371_n N_D[1]_c_372_n D[1]
+ N_D[1]_c_401_p PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%D[1]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%D[2] N_D[2]_c_406_n N_D[2]_M1000_g
+ N_D[2]_c_407_n N_D[2]_M1011_g N_D[2]_c_408_n N_D[2]_c_409_n D[2]
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%D[2]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%A_1012_265# N_A_1012_265#_M1022_s
+ N_A_1012_265#_M1014_s N_A_1012_265#_M1012_g N_A_1012_265#_c_443_n
+ N_A_1012_265#_c_444_n N_A_1012_265#_c_448_n N_A_1012_265#_c_445_n
+ N_A_1012_265#_c_446_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%A_1012_265#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%S[2] N_S[2]_c_499_n N_S[2]_M1004_g
+ N_S[2]_c_500_n N_S[2]_c_501_n N_S[2]_c_502_n N_S[2]_M1014_g N_S[2]_c_503_n
+ N_S[2]_M1022_g S[2] N_S[2]_c_504_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%S[2]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%S[3] N_S[3]_c_546_n N_S[3]_M1001_g
+ N_S[3]_c_547_n N_S[3]_M1015_g N_S[3]_c_548_n N_S[3]_c_549_n N_S[3]_M1002_g
+ S[3] N_S[3]_c_550_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%S[3]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%A_1361_47# N_A_1361_47#_M1015_d
+ N_A_1361_47#_M1001_d N_A_1361_47#_M1005_g N_A_1361_47#_c_594_n
+ N_A_1361_47#_c_589_n N_A_1361_47#_c_590_n N_A_1361_47#_c_591_n
+ N_A_1361_47#_c_592_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%A_1361_47#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%D[3] N_D[3]_c_644_n N_D[3]_M1008_g
+ N_D[3]_c_645_n N_D[3]_M1020_g N_D[3]_c_646_n N_D[3]_c_647_n D[3]
+ N_D[3]_c_667_p PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%D[3]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%VPWR N_VPWR_M1007_s N_VPWR_M1013_d
+ N_VPWR_M1019_d N_VPWR_M1014_d N_VPWR_M1008_d N_VPWR_c_673_n N_VPWR_c_674_n
+ N_VPWR_c_675_n N_VPWR_c_676_n N_VPWR_c_677_n N_VPWR_c_678_n N_VPWR_c_679_n
+ N_VPWR_c_680_n N_VPWR_c_681_n N_VPWR_c_682_n N_VPWR_c_683_n VPWR
+ N_VPWR_c_684_n N_VPWR_c_685_n N_VPWR_c_686_n N_VPWR_c_672_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%VPWR
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%Z N_Z_M1023_d N_Z_M1006_s N_Z_M1004_d
+ N_Z_M1002_s N_Z_M1009_d N_Z_M1003_s N_Z_M1012_d N_Z_M1005_s N_Z_c_804_n
+ N_Z_c_805_n N_Z_c_806_n N_Z_c_817_n N_Z_c_818_n N_Z_c_807_n N_Z_c_808_n
+ N_Z_c_809_n N_Z_c_810_n N_Z_c_811_n N_Z_c_821_n N_Z_c_822_n N_Z_c_812_n
+ N_Z_c_813_n N_Z_c_814_n N_Z_c_815_n N_Z_c_824_n N_Z_c_850_n N_Z_c_897_n
+ N_Z_c_884_n N_Z_c_825_n N_Z_c_923_n N_Z_c_826_n N_Z_c_827_n N_Z_c_957_n
+ N_Z_c_828_n Z N_Z_c_829_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%Z
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%VGND N_VGND_M1021_s N_VGND_M1017_d
+ N_VGND_M1018_d N_VGND_M1022_d N_VGND_M1020_d N_VGND_c_1039_n N_VGND_c_1040_n
+ N_VGND_c_1041_n N_VGND_c_1042_n N_VGND_c_1043_n N_VGND_c_1044_n
+ N_VGND_c_1045_n N_VGND_c_1046_n N_VGND_c_1047_n N_VGND_c_1048_n
+ N_VGND_c_1049_n VGND N_VGND_c_1050_n N_VGND_c_1051_n N_VGND_c_1052_n
+ N_VGND_c_1053_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%VGND
cc_1 VNB N_D[0]_c_140_n 0.0226847f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_D[0]_c_141_n 0.0309471f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_3 VNB N_D[0]_c_142_n 0.00249376f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_4 VNB N_D[0]_c_143_n 0.012124f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.19
cc_5 VNB N_A_184_265#_c_168_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_6 VNB N_A_184_265#_c_169_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_184_265#_c_170_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_184_265#_c_171_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_S[0]_c_224_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_10 VNB N_S[0]_c_225_n 0.0502713f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_11 VNB N_S[0]_c_226_n 0.00937382f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_12 VNB N_S[0]_c_227_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_13 VNB N_S[0]_c_228_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_14 VNB N_S[0]_c_229_n 0.0083332f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_15 VNB N_S[1]_c_270_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_16 VNB N_S[1]_c_271_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_17 VNB N_S[1]_c_272_n 0.0596452f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.625
cc_18 VNB N_S[1]_c_273_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_19 VNB N_S[1]_c_274_n 0.00817678f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_20 VNB N_A_533_47#_c_314_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_533_47#_c_315_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_533_47#_c_316_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_533_47#_c_317_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_D[1]_c_369_n 0.0251359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_25 VNB N_D[1]_c_370_n 0.0174886f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_26 VNB N_D[1]_c_371_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_27 VNB N_D[1]_c_372_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_D[2]_c_406_n 0.0174886f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_29 VNB N_D[2]_c_407_n 0.0251359f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_30 VNB N_D[2]_c_408_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_31 VNB N_D[2]_c_409_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.19
cc_32 VNB N_A_1012_265#_c_443_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_33 VNB N_A_1012_265#_c_444_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_1012_265#_c_445_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_1012_265#_c_446_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_S[2]_c_499_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_37 VNB N_S[2]_c_500_n 0.0502713f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_38 VNB N_S[2]_c_501_n 0.00937382f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_39 VNB N_S[2]_c_502_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_40 VNB N_S[2]_c_503_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_41 VNB N_S[2]_c_504_n 0.00817678f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_42 VNB N_S[3]_c_546_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_43 VNB N_S[3]_c_547_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_44 VNB N_S[3]_c_548_n 0.0596452f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.625
cc_45 VNB N_S[3]_c_549_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_46 VNB N_S[3]_c_550_n 0.0083332f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_47 VNB N_A_1361_47#_c_589_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_1361_47#_c_590_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_1361_47#_c_591_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_1361_47#_c_592_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_D[3]_c_644_n 0.0309471f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_52 VNB N_D[3]_c_645_n 0.0226847f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_53 VNB N_D[3]_c_646_n 0.00249376f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_54 VNB N_D[3]_c_647_n 0.012124f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VPWR_c_672_n 0.364621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_Z_c_804_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_Z_c_805_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_Z_c_806_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_Z_c_807_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_Z_c_808_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_Z_c_809_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_Z_c_810_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_Z_c_811_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_Z_c_812_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_Z_c_813_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_Z_c_814_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_Z_c_815_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1039_n 0.0113488f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1040_n 0.0320435f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.51
cc_70 VNB N_VGND_c_1041_n 0.00561737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1042_n 0.00902444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1043_n 0.00561737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1044_n 0.0113488f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1045_n 0.0320435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1046_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1047_n 0.00634747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1048_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1049_n 0.00634747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1050_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1051_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1052_n 0.00615512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1053_n 0.434155f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VPB N_D[0]_c_141_n 0.0335483f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_84 VPB N_D[0]_c_143_n 0.00458905f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_85 VPB N_A_184_265#_M1009_g 0.0269712f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_86 VPB N_A_184_265#_c_173_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.425
cc_87 VPB N_A_184_265#_c_170_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_184_265#_c_171_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_S[0]_c_227_n 0.0280252f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_90 VPB N_S[1]_c_270_n 0.0280248f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_91 VPB N_A_533_47#_M1003_g 0.0269712f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_92 VPB N_A_533_47#_c_319_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_93 VPB N_A_533_47#_c_315_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_533_47#_c_316_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_D[1]_c_369_n 0.0267097f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_96 VPB N_D[1]_c_372_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_D[2]_c_407_n 0.0267097f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_98 VPB N_D[2]_c_409_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_99 VPB N_A_1012_265#_M1012_g 0.0269712f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_100 VPB N_A_1012_265#_c_448_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.605
+ $Y2=0.425
cc_101 VPB N_A_1012_265#_c_445_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_1012_265#_c_446_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_S[2]_c_502_n 0.0280248f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_104 VPB N_S[3]_c_546_n 0.0280252f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_105 VPB N_A_1361_47#_M1005_g 0.0269712f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_106 VPB N_A_1361_47#_c_594_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_107 VPB N_A_1361_47#_c_590_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_1361_47#_c_591_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_D[3]_c_644_n 0.0335483f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_110 VPB N_D[3]_c_647_n 0.00458905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_673_n 0.0103693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_674_n 0.0425009f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=0.51
cc_113 VPB N_VPWR_c_675_n 0.017394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_676_n 4.89801e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_677_n 0.017394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_678_n 0.0103693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_679_n 0.0425009f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_680_n 0.0471219f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_681_n 0.00574453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_682_n 0.0461673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_683_n 0.00574453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_684_n 0.0461673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_685_n 0.0471219f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_686_n 0.0051677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_672_n 0.0575211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_Z_c_804_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_Z_c_817_n 0.00457032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_Z_c_818_n 0.00457032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_Z_c_808_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_Z_c_809_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_Z_c_821_n 0.00457032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_Z_c_822_n 0.00457032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_Z_c_813_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_Z_c_824_n 0.00809084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_Z_c_825_n 0.00809084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_Z_c_826_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_Z_c_827_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_Z_c_828_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_Z_c_829_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 N_D[0]_c_141_n N_A_184_265#_M1009_g 0.0381613f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_141 N_D[0]_c_141_n N_A_184_265#_c_171_n 0.00712672f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_142 N_D[0]_c_140_n N_S[0]_c_224_n 0.0286599f $X=0.47 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_143 N_D[0]_c_142_n N_S[0]_c_224_n 0.00289497f $X=0.645 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_144 N_D[0]_c_141_n N_VPWR_c_674_n 0.0245615f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_145 N_D[0]_c_143_n N_VPWR_c_674_n 0.00471543f $X=0.645 $Y=1.19 $X2=0 $Y2=0
cc_146 N_D[0]_c_141_n N_VPWR_c_680_n 0.00622633f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_147 N_D[0]_c_141_n N_VPWR_c_672_n 0.0106352f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_148 N_D[0]_c_141_n N_Z_c_804_n 0.00605747f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_149 N_D[0]_c_142_n N_Z_c_804_n 0.00376465f $X=0.645 $Y=1.055 $X2=0 $Y2=0
cc_150 N_D[0]_c_143_n N_Z_c_804_n 0.0216525f $X=0.645 $Y=1.19 $X2=0 $Y2=0
cc_151 N_D[0]_c_142_n N_Z_c_805_n 0.0128881f $X=0.645 $Y=1.055 $X2=0 $Y2=0
cc_152 N_D[0]_c_142_n N_Z_c_806_n 0.00686805f $X=0.645 $Y=1.055 $X2=0 $Y2=0
cc_153 N_D[0]_c_141_n N_Z_c_817_n 0.00145364f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_154 N_D[0]_c_140_n N_VGND_c_1040_n 0.00487865f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_155 N_D[0]_c_143_n N_VGND_c_1040_n 0.00222881f $X=0.645 $Y=1.19 $X2=0 $Y2=0
cc_156 N_D[0]_c_140_n N_VGND_c_1046_n 0.00585385f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_157 D[0] N_VGND_c_1046_n 0.00842546f $X=0.605 $Y=0.425 $X2=0 $Y2=0
cc_158 N_D[0]_c_140_n N_VGND_c_1053_n 0.011617f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_159 D[0] N_VGND_c_1053_n 0.00942277f $X=0.605 $Y=0.425 $X2=0 $Y2=0
cc_160 N_D[0]_c_142_n A_109_47# 0.00426617f $X=0.645 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_161 D[0] A_109_47# 0.00894235f $X=0.605 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_162 N_A_184_265#_c_168_n N_S[0]_c_225_n 0.00827389f $X=1.545 $Y=0.755 $X2=0
+ $Y2=0
cc_163 N_A_184_265#_c_169_n N_S[0]_c_225_n 0.0164662f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_164 N_A_184_265#_c_170_n N_S[0]_c_225_n 0.00928634f $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_165 N_A_184_265#_c_171_n N_S[0]_c_225_n 0.0184911f $X=1.02 $Y=1.34 $X2=0
+ $Y2=0
cc_166 N_A_184_265#_c_171_n N_S[0]_c_226_n 0.00820745f $X=1.02 $Y=1.34 $X2=0
+ $Y2=0
cc_167 N_A_184_265#_c_169_n N_S[0]_c_227_n 0.0012443f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_168 N_A_184_265#_c_173_n N_S[0]_c_227_n 0.00960233f $X=1.775 $Y=2.31 $X2=0
+ $Y2=0
cc_169 N_A_184_265#_c_170_n N_S[0]_c_227_n 0.00779252f $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_170 N_A_184_265#_c_171_n N_S[0]_c_227_n 0.00659591f $X=1.02 $Y=1.34 $X2=0
+ $Y2=0
cc_171 N_A_184_265#_c_169_n N_S[0]_c_228_n 0.00219336f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_172 N_A_184_265#_c_168_n N_S[0]_c_229_n 0.00603567f $X=1.545 $Y=0.755 $X2=0
+ $Y2=0
cc_173 N_A_184_265#_c_169_n N_S[0]_c_229_n 0.0176329f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_174 N_A_184_265#_c_170_n N_S[0]_c_229_n 0.0213691f $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_175 N_A_184_265#_c_171_n N_S[0]_c_229_n 2.54352e-19 $X=1.02 $Y=1.34 $X2=0
+ $Y2=0
cc_176 N_A_184_265#_M1009_g N_VPWR_c_674_n 0.00298082f $X=1.02 $Y=2.075 $X2=0
+ $Y2=0
cc_177 N_A_184_265#_c_173_n N_VPWR_c_675_n 0.0498301f $X=1.775 $Y=2.31 $X2=0
+ $Y2=0
cc_178 N_A_184_265#_c_170_n N_VPWR_c_675_n 0.0110094f $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_179 N_A_184_265#_M1009_g N_VPWR_c_680_n 0.00522699f $X=1.02 $Y=2.075 $X2=0
+ $Y2=0
cc_180 N_A_184_265#_c_173_n N_VPWR_c_680_n 0.0210596f $X=1.775 $Y=2.31 $X2=0
+ $Y2=0
cc_181 N_A_184_265#_M1013_s N_VPWR_c_672_n 0.00179197f $X=1.65 $Y=1.485 $X2=0
+ $Y2=0
cc_182 N_A_184_265#_M1009_g N_VPWR_c_672_n 0.00828927f $X=1.02 $Y=2.075 $X2=0
+ $Y2=0
cc_183 N_A_184_265#_c_173_n N_VPWR_c_672_n 0.00594162f $X=1.775 $Y=2.31 $X2=0
+ $Y2=0
cc_184 N_A_184_265#_M1009_g N_Z_c_804_n 0.00862328f $X=1.02 $Y=2.075 $X2=0 $Y2=0
cc_185 N_A_184_265#_c_169_n N_Z_c_804_n 0.00719188f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_186 N_A_184_265#_c_173_n N_Z_c_804_n 0.00378484f $X=1.775 $Y=2.31 $X2=0 $Y2=0
cc_187 N_A_184_265#_c_170_n N_Z_c_804_n 0.0304368f $X=1.775 $Y=1.63 $X2=0 $Y2=0
cc_188 N_A_184_265#_c_171_n N_Z_c_804_n 0.00814206f $X=1.02 $Y=1.34 $X2=0 $Y2=0
cc_189 N_A_184_265#_c_169_n N_Z_c_805_n 0.0124144f $X=1.545 $Y=1.175 $X2=0 $Y2=0
cc_190 N_A_184_265#_c_170_n N_Z_c_805_n 0.00398133f $X=1.775 $Y=1.63 $X2=0 $Y2=0
cc_191 N_A_184_265#_c_171_n N_Z_c_805_n 0.00349316f $X=1.02 $Y=1.34 $X2=0 $Y2=0
cc_192 N_A_184_265#_c_168_n N_Z_c_806_n 0.0259454f $X=1.545 $Y=0.755 $X2=0 $Y2=0
cc_193 N_A_184_265#_c_169_n N_Z_c_806_n 0.00611965f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_194 N_A_184_265#_M1009_g N_Z_c_817_n 0.00988241f $X=1.02 $Y=2.075 $X2=0 $Y2=0
cc_195 N_A_184_265#_c_173_n N_Z_c_817_n 0.0369227f $X=1.775 $Y=2.31 $X2=0 $Y2=0
cc_196 N_A_184_265#_c_173_n N_Z_c_824_n 0.0293762f $X=1.775 $Y=2.31 $X2=0 $Y2=0
cc_197 N_A_184_265#_c_170_n N_Z_c_824_n 0.0126642f $X=1.775 $Y=1.63 $X2=0 $Y2=0
cc_198 N_A_184_265#_M1009_g N_Z_c_850_n 0.00289142f $X=1.02 $Y=2.075 $X2=0 $Y2=0
cc_199 N_A_184_265#_c_173_n N_Z_c_850_n 6.03258e-19 $X=1.775 $Y=2.31 $X2=0 $Y2=0
cc_200 N_A_184_265#_c_170_n N_Z_c_850_n 4.25753e-19 $X=1.775 $Y=1.63 $X2=0 $Y2=0
cc_201 N_A_184_265#_M1009_g N_Z_c_829_n 0.0105217f $X=1.02 $Y=2.075 $X2=0 $Y2=0
cc_202 N_A_184_265#_c_173_n N_Z_c_829_n 0.0139746f $X=1.775 $Y=2.31 $X2=0 $Y2=0
cc_203 N_A_184_265#_c_170_n N_Z_c_829_n 0.00749676f $X=1.775 $Y=1.63 $X2=0 $Y2=0
cc_204 N_A_184_265#_c_171_n N_Z_c_829_n 0.00449162f $X=1.02 $Y=1.34 $X2=0 $Y2=0
cc_205 N_A_184_265#_c_168_n N_VGND_c_1046_n 0.015238f $X=1.545 $Y=0.755 $X2=0
+ $Y2=0
cc_206 N_A_184_265#_M1017_s N_VGND_c_1053_n 0.00358139f $X=1.65 $Y=0.235 $X2=0
+ $Y2=0
cc_207 N_A_184_265#_c_168_n N_VGND_c_1053_n 0.0150148f $X=1.545 $Y=0.755 $X2=0
+ $Y2=0
cc_208 N_S[0]_c_227_n N_S[1]_c_270_n 0.057922f $X=2.01 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_209 N_S[0]_c_229_n N_S[1]_c_270_n 0.00132881f $X=1.975 $Y=1.03 $X2=-0.19
+ $Y2=-0.24
cc_210 N_S[0]_c_228_n N_S[1]_c_271_n 0.0091402f $X=2.01 $Y=0.83 $X2=0 $Y2=0
cc_211 N_S[0]_c_227_n N_S[1]_c_274_n 0.00132881f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_212 N_S[0]_c_229_n N_S[1]_c_274_n 0.0202885f $X=1.975 $Y=1.03 $X2=0 $Y2=0
cc_213 N_S[0]_c_227_n N_VPWR_c_675_n 0.013047f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_214 N_S[0]_c_227_n N_VPWR_c_680_n 0.00673617f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_215 N_S[0]_c_227_n N_VPWR_c_672_n 0.00878911f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_216 N_S[0]_c_226_n N_Z_c_804_n 7.46972e-19 $X=1.02 $Y=0.905 $X2=0 $Y2=0
cc_217 N_S[0]_c_225_n N_Z_c_805_n 0.00806549f $X=1.84 $Y=0.905 $X2=0 $Y2=0
cc_218 N_S[0]_c_226_n N_Z_c_805_n 0.00605736f $X=1.02 $Y=0.905 $X2=0 $Y2=0
cc_219 N_S[0]_c_224_n N_Z_c_806_n 0.00316445f $X=0.945 $Y=0.83 $X2=0 $Y2=0
cc_220 N_S[0]_c_225_n N_Z_c_806_n 0.00501353f $X=1.84 $Y=0.905 $X2=0 $Y2=0
cc_221 N_S[0]_c_227_n N_Z_c_824_n 0.00637646f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_222 N_S[0]_c_229_n N_Z_c_824_n 0.00698535f $X=1.975 $Y=1.03 $X2=0 $Y2=0
cc_223 N_S[0]_c_228_n N_VGND_c_1041_n 0.00570474f $X=2.01 $Y=0.83 $X2=0 $Y2=0
cc_224 N_S[0]_c_229_n N_VGND_c_1041_n 8.9983e-19 $X=1.975 $Y=1.03 $X2=0 $Y2=0
cc_225 N_S[0]_c_224_n N_VGND_c_1046_n 0.00585385f $X=0.945 $Y=0.83 $X2=0 $Y2=0
cc_226 N_S[0]_c_228_n N_VGND_c_1046_n 0.00585385f $X=2.01 $Y=0.83 $X2=0 $Y2=0
cc_227 N_S[0]_c_224_n N_VGND_c_1053_n 0.00880034f $X=0.945 $Y=0.83 $X2=0 $Y2=0
cc_228 N_S[0]_c_225_n N_VGND_c_1053_n 0.00349917f $X=1.84 $Y=0.905 $X2=0 $Y2=0
cc_229 N_S[0]_c_227_n N_VGND_c_1053_n 6.15795e-19 $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_230 N_S[0]_c_228_n N_VGND_c_1053_n 0.0124506f $X=2.01 $Y=0.83 $X2=0 $Y2=0
cc_231 N_S[1]_c_270_n N_A_533_47#_c_319_n 0.00903826f $X=2.59 $Y=1.41 $X2=0
+ $Y2=0
cc_232 N_S[1]_c_270_n N_A_533_47#_c_314_n 0.0012443f $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_233 N_S[1]_c_271_n N_A_533_47#_c_314_n 0.00219336f $X=2.59 $Y=0.83 $X2=0
+ $Y2=0
cc_234 N_S[1]_c_272_n N_A_533_47#_c_314_n 0.0164662f $X=3.58 $Y=0.905 $X2=0
+ $Y2=0
cc_235 N_S[1]_c_274_n N_A_533_47#_c_314_n 0.0176329f $X=2.625 $Y=1.03 $X2=0
+ $Y2=0
cc_236 N_S[1]_c_270_n N_A_533_47#_c_315_n 0.00767015f $X=2.59 $Y=1.41 $X2=0
+ $Y2=0
cc_237 N_S[1]_c_272_n N_A_533_47#_c_315_n 0.00928634f $X=3.58 $Y=0.905 $X2=0
+ $Y2=0
cc_238 N_S[1]_c_274_n N_A_533_47#_c_315_n 0.0213691f $X=2.625 $Y=1.03 $X2=0
+ $Y2=0
cc_239 N_S[1]_c_270_n N_A_533_47#_c_316_n 0.00659591f $X=2.59 $Y=1.41 $X2=0
+ $Y2=0
cc_240 N_S[1]_c_272_n N_A_533_47#_c_316_n 0.0266986f $X=3.58 $Y=0.905 $X2=0
+ $Y2=0
cc_241 N_S[1]_c_274_n N_A_533_47#_c_316_n 2.54352e-19 $X=2.625 $Y=1.03 $X2=0
+ $Y2=0
cc_242 N_S[1]_c_270_n N_A_533_47#_c_317_n 0.00827389f $X=2.59 $Y=1.41 $X2=0
+ $Y2=0
cc_243 N_S[1]_c_274_n N_A_533_47#_c_317_n 0.00603567f $X=2.625 $Y=1.03 $X2=0
+ $Y2=0
cc_244 N_S[1]_c_273_n N_D[1]_c_370_n 0.0286599f $X=3.655 $Y=0.83 $X2=0 $Y2=0
cc_245 N_S[1]_c_273_n N_D[1]_c_371_n 0.00289497f $X=3.655 $Y=0.83 $X2=0 $Y2=0
cc_246 N_S[1]_c_270_n N_VPWR_c_675_n 0.00962409f $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_247 N_S[1]_c_274_n N_VPWR_c_675_n 0.00155482f $X=2.625 $Y=1.03 $X2=0 $Y2=0
cc_248 N_S[1]_c_270_n N_VPWR_c_684_n 0.00673617f $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_249 N_S[1]_c_270_n N_VPWR_c_672_n 0.00871384f $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_250 N_S[1]_c_272_n N_Z_c_807_n 0.00501353f $X=3.58 $Y=0.905 $X2=0 $Y2=0
cc_251 N_S[1]_c_273_n N_Z_c_807_n 0.00316445f $X=3.655 $Y=0.83 $X2=0 $Y2=0
cc_252 N_S[1]_c_272_n N_Z_c_808_n 7.46972e-19 $X=3.58 $Y=0.905 $X2=0 $Y2=0
cc_253 N_S[1]_c_272_n N_Z_c_814_n 0.0141229f $X=3.58 $Y=0.905 $X2=0 $Y2=0
cc_254 N_S[1]_c_270_n N_Z_c_824_n 0.0062071f $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_255 N_S[1]_c_274_n N_Z_c_824_n 0.00638667f $X=2.625 $Y=1.03 $X2=0 $Y2=0
cc_256 N_S[1]_c_271_n N_VGND_c_1041_n 0.00570474f $X=2.59 $Y=0.83 $X2=0 $Y2=0
cc_257 N_S[1]_c_274_n N_VGND_c_1041_n 8.9983e-19 $X=2.625 $Y=1.03 $X2=0 $Y2=0
cc_258 N_S[1]_c_271_n N_VGND_c_1050_n 0.00585385f $X=2.59 $Y=0.83 $X2=0 $Y2=0
cc_259 N_S[1]_c_273_n N_VGND_c_1050_n 0.00585385f $X=3.655 $Y=0.83 $X2=0 $Y2=0
cc_260 N_S[1]_c_270_n N_VGND_c_1053_n 6.15795e-19 $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_261 N_S[1]_c_271_n N_VGND_c_1053_n 0.0124506f $X=2.59 $Y=0.83 $X2=0 $Y2=0
cc_262 N_S[1]_c_272_n N_VGND_c_1053_n 0.00349917f $X=3.58 $Y=0.905 $X2=0 $Y2=0
cc_263 N_S[1]_c_273_n N_VGND_c_1053_n 0.00880034f $X=3.655 $Y=0.83 $X2=0 $Y2=0
cc_264 N_A_533_47#_M1003_g N_D[1]_c_369_n 0.0388862f $X=3.58 $Y=2.075 $X2=-0.19
+ $Y2=-0.24
cc_265 N_A_533_47#_c_316_n N_D[1]_c_369_n 0.00712672f $X=3.275 $Y=1.34 $X2=-0.19
+ $Y2=-0.24
cc_266 N_A_533_47#_c_319_n N_VPWR_c_675_n 0.02928f $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_267 N_A_533_47#_c_315_n N_VPWR_c_675_n 0.00687548f $X=3.055 $Y=1.405 $X2=0
+ $Y2=0
cc_268 N_A_533_47#_M1003_g N_VPWR_c_676_n 0.0030953f $X=3.58 $Y=2.075 $X2=0
+ $Y2=0
cc_269 N_A_533_47#_M1003_g N_VPWR_c_684_n 0.00522699f $X=3.58 $Y=2.075 $X2=0
+ $Y2=0
cc_270 N_A_533_47#_c_319_n N_VPWR_c_684_n 0.0210596f $X=2.825 $Y=2.31 $X2=0
+ $Y2=0
cc_271 N_A_533_47#_M1010_d N_VPWR_c_672_n 0.00179197f $X=2.68 $Y=1.485 $X2=0
+ $Y2=0
cc_272 N_A_533_47#_M1003_g N_VPWR_c_672_n 0.00809563f $X=3.58 $Y=2.075 $X2=0
+ $Y2=0
cc_273 N_A_533_47#_c_319_n N_VPWR_c_672_n 0.00594162f $X=2.825 $Y=2.31 $X2=0
+ $Y2=0
cc_274 N_A_533_47#_M1003_g N_Z_c_818_n 0.00988241f $X=3.58 $Y=2.075 $X2=0 $Y2=0
cc_275 N_A_533_47#_c_319_n N_Z_c_818_n 0.0369227f $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_276 N_A_533_47#_c_314_n N_Z_c_807_n 0.00611965f $X=3.055 $Y=1.175 $X2=0 $Y2=0
cc_277 N_A_533_47#_c_317_n N_Z_c_807_n 0.0259454f $X=2.825 $Y=0.495 $X2=0 $Y2=0
cc_278 N_A_533_47#_M1003_g N_Z_c_808_n 0.00862328f $X=3.58 $Y=2.075 $X2=0 $Y2=0
cc_279 N_A_533_47#_c_319_n N_Z_c_808_n 0.00378484f $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_280 N_A_533_47#_c_314_n N_Z_c_808_n 0.00719188f $X=3.055 $Y=1.175 $X2=0 $Y2=0
cc_281 N_A_533_47#_c_315_n N_Z_c_808_n 0.0304368f $X=3.055 $Y=1.405 $X2=0 $Y2=0
cc_282 N_A_533_47#_c_316_n N_Z_c_808_n 0.00814206f $X=3.275 $Y=1.34 $X2=0 $Y2=0
cc_283 N_A_533_47#_c_314_n N_Z_c_814_n 0.0124144f $X=3.055 $Y=1.175 $X2=0 $Y2=0
cc_284 N_A_533_47#_c_315_n N_Z_c_814_n 0.00398133f $X=3.055 $Y=1.405 $X2=0 $Y2=0
cc_285 N_A_533_47#_c_316_n N_Z_c_814_n 0.00349316f $X=3.275 $Y=1.34 $X2=0 $Y2=0
cc_286 N_A_533_47#_c_319_n N_Z_c_824_n 0.0291787f $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_287 N_A_533_47#_c_315_n N_Z_c_824_n 0.0126642f $X=3.055 $Y=1.405 $X2=0 $Y2=0
cc_288 N_A_533_47#_M1003_g N_Z_c_884_n 0.00289142f $X=3.58 $Y=2.075 $X2=0 $Y2=0
cc_289 N_A_533_47#_c_319_n N_Z_c_884_n 6.03258e-19 $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_290 N_A_533_47#_c_315_n N_Z_c_884_n 4.25753e-19 $X=3.055 $Y=1.405 $X2=0 $Y2=0
cc_291 N_A_533_47#_M1003_g N_Z_c_826_n 0.0105217f $X=3.58 $Y=2.075 $X2=0 $Y2=0
cc_292 N_A_533_47#_c_319_n N_Z_c_826_n 0.0139746f $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_293 N_A_533_47#_c_315_n N_Z_c_826_n 0.00749676f $X=3.055 $Y=1.405 $X2=0 $Y2=0
cc_294 N_A_533_47#_c_316_n N_Z_c_826_n 0.00449162f $X=3.275 $Y=1.34 $X2=0 $Y2=0
cc_295 N_A_533_47#_c_317_n N_VGND_c_1050_n 0.015238f $X=2.825 $Y=0.495 $X2=0
+ $Y2=0
cc_296 N_A_533_47#_M1016_d N_VGND_c_1053_n 0.00358139f $X=2.665 $Y=0.235 $X2=0
+ $Y2=0
cc_297 N_A_533_47#_c_317_n N_VGND_c_1053_n 0.0150148f $X=2.825 $Y=0.495 $X2=0
+ $Y2=0
cc_298 N_D[1]_c_370_n N_D[2]_c_406_n 0.00915308f $X=4.13 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_299 N_D[1]_c_369_n N_D[2]_c_407_n 0.0270908f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_300 N_D[1]_c_372_n N_D[2]_c_407_n 9.4377e-19 $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_301 N_D[1]_c_371_n N_D[2]_c_408_n 0.00442615f $X=3.955 $Y=1.055 $X2=0 $Y2=0
cc_302 N_D[1]_c_369_n N_D[2]_c_409_n 9.4377e-19 $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_303 N_D[1]_c_372_n N_D[2]_c_409_n 0.0199139f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_304 N_D[1]_c_369_n N_VPWR_c_676_n 0.0231278f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_305 N_D[1]_c_372_n N_VPWR_c_676_n 0.0044581f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_306 N_D[1]_c_369_n N_VPWR_c_684_n 0.00622633f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_307 N_D[1]_c_369_n N_VPWR_c_672_n 0.00594051f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_308 N_D[1]_c_369_n N_Z_c_818_n 0.00145364f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_309 N_D[1]_c_371_n N_Z_c_807_n 0.00686805f $X=3.955 $Y=1.055 $X2=0 $Y2=0
cc_310 N_D[1]_c_369_n N_Z_c_808_n 0.00605747f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_311 N_D[1]_c_371_n N_Z_c_808_n 0.00376465f $X=3.955 $Y=1.055 $X2=0 $Y2=0
cc_312 N_D[1]_c_372_n N_Z_c_808_n 0.0216525f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_313 N_D[1]_c_371_n N_Z_c_814_n 0.0128881f $X=3.955 $Y=1.055 $X2=0 $Y2=0
cc_314 N_D[1]_c_369_n N_Z_c_897_n 0.00719456f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_315 N_D[1]_c_372_n N_Z_c_897_n 0.00989895f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_316 N_D[1]_c_369_n N_Z_c_826_n 8.42164e-19 $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_317 N_D[1]_c_370_n N_VGND_c_1042_n 0.00322791f $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_318 N_D[1]_c_372_n N_VGND_c_1042_n 0.00222881f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_319 N_D[1]_c_370_n N_VGND_c_1050_n 0.00585385f $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_320 N_D[1]_c_401_p N_VGND_c_1050_n 0.00842546f $X=3.955 $Y=0.51 $X2=0 $Y2=0
cc_321 N_D[1]_c_370_n N_VGND_c_1053_n 0.0108306f $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_322 N_D[1]_c_401_p N_VGND_c_1053_n 0.00942277f $X=3.955 $Y=0.51 $X2=0 $Y2=0
cc_323 N_D[1]_c_371_n A_746_47# 0.00426617f $X=3.955 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_324 N_D[1]_c_401_p A_746_47# 0.00894235f $X=3.955 $Y=0.51 $X2=-0.19 $Y2=-0.24
cc_325 N_D[2]_c_407_n N_A_1012_265#_M1012_g 0.0388862f $X=4.635 $Y=1.41 $X2=0
+ $Y2=0
cc_326 N_D[2]_c_407_n N_A_1012_265#_c_446_n 0.00712672f $X=4.635 $Y=1.41 $X2=0
+ $Y2=0
cc_327 N_D[2]_c_406_n N_S[2]_c_499_n 0.0286599f $X=4.61 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_328 N_D[2]_c_408_n N_S[2]_c_499_n 0.00289497f $X=4.785 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_329 N_D[2]_c_407_n N_VPWR_c_676_n 0.0231278f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_330 N_D[2]_c_409_n N_VPWR_c_676_n 0.0044581f $X=4.785 $Y=1.19 $X2=0 $Y2=0
cc_331 N_D[2]_c_407_n N_VPWR_c_682_n 0.00622633f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_332 N_D[2]_c_407_n N_VPWR_c_672_n 0.00594051f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_333 N_D[2]_c_407_n N_Z_c_809_n 0.00605747f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_334 N_D[2]_c_408_n N_Z_c_809_n 0.00376465f $X=4.785 $Y=1.055 $X2=0 $Y2=0
cc_335 N_D[2]_c_409_n N_Z_c_809_n 0.0216525f $X=4.785 $Y=1.19 $X2=0 $Y2=0
cc_336 N_D[2]_c_408_n N_Z_c_810_n 0.0128881f $X=4.785 $Y=1.055 $X2=0 $Y2=0
cc_337 N_D[2]_c_408_n N_Z_c_811_n 0.00686805f $X=4.785 $Y=1.055 $X2=0 $Y2=0
cc_338 N_D[2]_c_407_n N_Z_c_821_n 0.00145364f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_339 N_D[2]_c_407_n N_Z_c_897_n 0.00719456f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_340 N_D[2]_c_409_n N_Z_c_897_n 0.00989895f $X=4.785 $Y=1.19 $X2=0 $Y2=0
cc_341 N_D[2]_c_407_n N_Z_c_827_n 8.42164e-19 $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_342 N_D[2]_c_406_n N_VGND_c_1042_n 0.00322791f $X=4.61 $Y=0.995 $X2=0 $Y2=0
cc_343 N_D[2]_c_409_n N_VGND_c_1042_n 0.00222881f $X=4.785 $Y=1.19 $X2=0 $Y2=0
cc_344 N_D[2]_c_406_n N_VGND_c_1048_n 0.00585385f $X=4.61 $Y=0.995 $X2=0 $Y2=0
cc_345 D[2] N_VGND_c_1048_n 0.00842546f $X=4.745 $Y=0.425 $X2=0 $Y2=0
cc_346 N_D[2]_c_406_n N_VGND_c_1053_n 0.0108306f $X=4.61 $Y=0.995 $X2=0 $Y2=0
cc_347 D[2] N_VGND_c_1053_n 0.00942277f $X=4.745 $Y=0.425 $X2=0 $Y2=0
cc_348 N_D[2]_c_408_n A_937_47# 0.00426617f $X=4.785 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_349 D[2] A_937_47# 0.00894235f $X=4.745 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_350 N_A_1012_265#_c_443_n N_S[2]_c_500_n 0.00827389f $X=5.685 $Y=0.755 $X2=0
+ $Y2=0
cc_351 N_A_1012_265#_c_444_n N_S[2]_c_500_n 0.0164662f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_352 N_A_1012_265#_c_445_n N_S[2]_c_500_n 0.00928634f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_353 N_A_1012_265#_c_446_n N_S[2]_c_500_n 0.0184911f $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_354 N_A_1012_265#_c_446_n N_S[2]_c_501_n 0.00820745f $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_355 N_A_1012_265#_c_444_n N_S[2]_c_502_n 0.0012443f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_356 N_A_1012_265#_c_448_n N_S[2]_c_502_n 0.00903826f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_357 N_A_1012_265#_c_445_n N_S[2]_c_502_n 0.00767015f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_358 N_A_1012_265#_c_446_n N_S[2]_c_502_n 0.00659591f $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_359 N_A_1012_265#_c_444_n N_S[2]_c_503_n 0.00219336f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_360 N_A_1012_265#_c_443_n N_S[2]_c_504_n 0.00603567f $X=5.685 $Y=0.755 $X2=0
+ $Y2=0
cc_361 N_A_1012_265#_c_444_n N_S[2]_c_504_n 0.0176329f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_362 N_A_1012_265#_c_445_n N_S[2]_c_504_n 0.0213691f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_363 N_A_1012_265#_c_446_n N_S[2]_c_504_n 2.54352e-19 $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_364 N_A_1012_265#_M1012_g N_VPWR_c_676_n 0.0030953f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_365 N_A_1012_265#_c_448_n N_VPWR_c_677_n 0.02928f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_366 N_A_1012_265#_c_445_n N_VPWR_c_677_n 0.00687548f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_367 N_A_1012_265#_M1012_g N_VPWR_c_682_n 0.00522699f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_368 N_A_1012_265#_c_448_n N_VPWR_c_682_n 0.0210596f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_369 N_A_1012_265#_M1014_s N_VPWR_c_672_n 0.00179197f $X=5.79 $Y=1.485 $X2=0
+ $Y2=0
cc_370 N_A_1012_265#_M1012_g N_VPWR_c_672_n 0.00809563f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_371 N_A_1012_265#_c_448_n N_VPWR_c_672_n 0.00594162f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_372 N_A_1012_265#_M1012_g N_Z_c_809_n 0.00862328f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_373 N_A_1012_265#_c_444_n N_Z_c_809_n 0.00719188f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_374 N_A_1012_265#_c_448_n N_Z_c_809_n 0.00378484f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_375 N_A_1012_265#_c_445_n N_Z_c_809_n 0.0304368f $X=5.915 $Y=1.63 $X2=0 $Y2=0
cc_376 N_A_1012_265#_c_446_n N_Z_c_809_n 0.00814206f $X=5.16 $Y=1.34 $X2=0 $Y2=0
cc_377 N_A_1012_265#_c_444_n N_Z_c_810_n 0.0124144f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_378 N_A_1012_265#_c_445_n N_Z_c_810_n 0.00398133f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_379 N_A_1012_265#_c_446_n N_Z_c_810_n 0.00349316f $X=5.16 $Y=1.34 $X2=0 $Y2=0
cc_380 N_A_1012_265#_c_443_n N_Z_c_811_n 0.0259454f $X=5.685 $Y=0.755 $X2=0
+ $Y2=0
cc_381 N_A_1012_265#_c_444_n N_Z_c_811_n 0.00611965f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_382 N_A_1012_265#_M1012_g N_Z_c_821_n 0.00988241f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_383 N_A_1012_265#_c_448_n N_Z_c_821_n 0.0369227f $X=5.915 $Y=2.31 $X2=0 $Y2=0
cc_384 N_A_1012_265#_c_448_n N_Z_c_825_n 0.0291787f $X=5.915 $Y=2.31 $X2=0 $Y2=0
cc_385 N_A_1012_265#_c_445_n N_Z_c_825_n 0.0126642f $X=5.915 $Y=1.63 $X2=0 $Y2=0
cc_386 N_A_1012_265#_M1012_g N_Z_c_923_n 0.00289142f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_387 N_A_1012_265#_c_448_n N_Z_c_923_n 6.03258e-19 $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_388 N_A_1012_265#_c_445_n N_Z_c_923_n 4.25753e-19 $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_389 N_A_1012_265#_M1012_g N_Z_c_827_n 0.0105217f $X=5.16 $Y=2.075 $X2=0 $Y2=0
cc_390 N_A_1012_265#_c_448_n N_Z_c_827_n 0.0139746f $X=5.915 $Y=2.31 $X2=0 $Y2=0
cc_391 N_A_1012_265#_c_445_n N_Z_c_827_n 0.00749676f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_392 N_A_1012_265#_c_446_n N_Z_c_827_n 0.00449162f $X=5.16 $Y=1.34 $X2=0 $Y2=0
cc_393 N_A_1012_265#_c_443_n N_VGND_c_1048_n 0.015238f $X=5.685 $Y=0.755 $X2=0
+ $Y2=0
cc_394 N_A_1012_265#_M1022_s N_VGND_c_1053_n 0.00358139f $X=5.79 $Y=0.235 $X2=0
+ $Y2=0
cc_395 N_A_1012_265#_c_443_n N_VGND_c_1053_n 0.0150148f $X=5.685 $Y=0.755 $X2=0
+ $Y2=0
cc_396 N_S[2]_c_502_n N_S[3]_c_546_n 0.057922f $X=6.15 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_397 N_S[2]_c_504_n N_S[3]_c_546_n 0.00132881f $X=6.115 $Y=1.03 $X2=-0.19
+ $Y2=-0.24
cc_398 N_S[2]_c_503_n N_S[3]_c_547_n 0.0091402f $X=6.15 $Y=0.83 $X2=0 $Y2=0
cc_399 N_S[2]_c_502_n N_S[3]_c_550_n 0.00132881f $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_400 N_S[2]_c_504_n N_S[3]_c_550_n 0.0202885f $X=6.115 $Y=1.03 $X2=0 $Y2=0
cc_401 N_S[2]_c_502_n N_VPWR_c_677_n 0.00962409f $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_402 N_S[2]_c_504_n N_VPWR_c_677_n 0.00155482f $X=6.115 $Y=1.03 $X2=0 $Y2=0
cc_403 N_S[2]_c_502_n N_VPWR_c_682_n 0.00673617f $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_404 N_S[2]_c_502_n N_VPWR_c_672_n 0.00871384f $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_405 N_S[2]_c_501_n N_Z_c_809_n 7.46972e-19 $X=5.16 $Y=0.905 $X2=0 $Y2=0
cc_406 N_S[2]_c_500_n N_Z_c_810_n 0.00806549f $X=5.98 $Y=0.905 $X2=0 $Y2=0
cc_407 N_S[2]_c_501_n N_Z_c_810_n 0.00605736f $X=5.16 $Y=0.905 $X2=0 $Y2=0
cc_408 N_S[2]_c_499_n N_Z_c_811_n 0.00316445f $X=5.085 $Y=0.83 $X2=0 $Y2=0
cc_409 N_S[2]_c_500_n N_Z_c_811_n 0.00501353f $X=5.98 $Y=0.905 $X2=0 $Y2=0
cc_410 N_S[2]_c_502_n N_Z_c_825_n 0.0062071f $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_411 N_S[2]_c_504_n N_Z_c_825_n 0.00638667f $X=6.115 $Y=1.03 $X2=0 $Y2=0
cc_412 N_S[2]_c_503_n N_VGND_c_1043_n 0.00570474f $X=6.15 $Y=0.83 $X2=0 $Y2=0
cc_413 N_S[2]_c_504_n N_VGND_c_1043_n 8.9983e-19 $X=6.115 $Y=1.03 $X2=0 $Y2=0
cc_414 N_S[2]_c_499_n N_VGND_c_1048_n 0.00585385f $X=5.085 $Y=0.83 $X2=0 $Y2=0
cc_415 N_S[2]_c_503_n N_VGND_c_1048_n 0.00585385f $X=6.15 $Y=0.83 $X2=0 $Y2=0
cc_416 N_S[2]_c_499_n N_VGND_c_1053_n 0.00880034f $X=5.085 $Y=0.83 $X2=0 $Y2=0
cc_417 N_S[2]_c_500_n N_VGND_c_1053_n 0.00349917f $X=5.98 $Y=0.905 $X2=0 $Y2=0
cc_418 N_S[2]_c_502_n N_VGND_c_1053_n 6.15795e-19 $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_419 N_S[2]_c_503_n N_VGND_c_1053_n 0.0124506f $X=6.15 $Y=0.83 $X2=0 $Y2=0
cc_420 N_S[3]_c_546_n N_A_1361_47#_c_594_n 0.00960233f $X=6.73 $Y=1.41 $X2=0
+ $Y2=0
cc_421 N_S[3]_c_546_n N_A_1361_47#_c_589_n 0.0012443f $X=6.73 $Y=1.41 $X2=0
+ $Y2=0
cc_422 N_S[3]_c_547_n N_A_1361_47#_c_589_n 0.00219336f $X=6.73 $Y=0.83 $X2=0
+ $Y2=0
cc_423 N_S[3]_c_548_n N_A_1361_47#_c_589_n 0.0164662f $X=7.72 $Y=0.905 $X2=0
+ $Y2=0
cc_424 N_S[3]_c_550_n N_A_1361_47#_c_589_n 0.0176329f $X=6.765 $Y=1.03 $X2=0
+ $Y2=0
cc_425 N_S[3]_c_546_n N_A_1361_47#_c_590_n 0.00779252f $X=6.73 $Y=1.41 $X2=0
+ $Y2=0
cc_426 N_S[3]_c_548_n N_A_1361_47#_c_590_n 0.00928634f $X=7.72 $Y=0.905 $X2=0
+ $Y2=0
cc_427 N_S[3]_c_550_n N_A_1361_47#_c_590_n 0.0213691f $X=6.765 $Y=1.03 $X2=0
+ $Y2=0
cc_428 N_S[3]_c_546_n N_A_1361_47#_c_591_n 0.00659591f $X=6.73 $Y=1.41 $X2=0
+ $Y2=0
cc_429 N_S[3]_c_548_n N_A_1361_47#_c_591_n 0.0266986f $X=7.72 $Y=0.905 $X2=0
+ $Y2=0
cc_430 N_S[3]_c_550_n N_A_1361_47#_c_591_n 2.54352e-19 $X=6.765 $Y=1.03 $X2=0
+ $Y2=0
cc_431 N_S[3]_c_546_n N_A_1361_47#_c_592_n 0.00827389f $X=6.73 $Y=1.41 $X2=0
+ $Y2=0
cc_432 N_S[3]_c_550_n N_A_1361_47#_c_592_n 0.00603567f $X=6.765 $Y=1.03 $X2=0
+ $Y2=0
cc_433 N_S[3]_c_549_n N_D[3]_c_645_n 0.0286599f $X=7.795 $Y=0.83 $X2=0 $Y2=0
cc_434 N_S[3]_c_549_n N_D[3]_c_646_n 0.00289497f $X=7.795 $Y=0.83 $X2=0 $Y2=0
cc_435 N_S[3]_c_546_n N_VPWR_c_677_n 0.013047f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_436 N_S[3]_c_546_n N_VPWR_c_685_n 0.00673617f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_437 N_S[3]_c_546_n N_VPWR_c_672_n 0.00878911f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_438 N_S[3]_c_548_n N_Z_c_812_n 0.00501353f $X=7.72 $Y=0.905 $X2=0 $Y2=0
cc_439 N_S[3]_c_549_n N_Z_c_812_n 0.00316445f $X=7.795 $Y=0.83 $X2=0 $Y2=0
cc_440 N_S[3]_c_548_n N_Z_c_813_n 7.46972e-19 $X=7.72 $Y=0.905 $X2=0 $Y2=0
cc_441 N_S[3]_c_548_n N_Z_c_815_n 0.0141229f $X=7.72 $Y=0.905 $X2=0 $Y2=0
cc_442 N_S[3]_c_546_n N_Z_c_825_n 0.00637646f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_443 N_S[3]_c_550_n N_Z_c_825_n 0.00698535f $X=6.765 $Y=1.03 $X2=0 $Y2=0
cc_444 N_S[3]_c_547_n N_VGND_c_1043_n 0.00570474f $X=6.73 $Y=0.83 $X2=0 $Y2=0
cc_445 N_S[3]_c_550_n N_VGND_c_1043_n 8.9983e-19 $X=6.765 $Y=1.03 $X2=0 $Y2=0
cc_446 N_S[3]_c_547_n N_VGND_c_1051_n 0.00585385f $X=6.73 $Y=0.83 $X2=0 $Y2=0
cc_447 N_S[3]_c_549_n N_VGND_c_1051_n 0.00585385f $X=7.795 $Y=0.83 $X2=0 $Y2=0
cc_448 N_S[3]_c_546_n N_VGND_c_1053_n 6.15795e-19 $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_449 N_S[3]_c_547_n N_VGND_c_1053_n 0.0124506f $X=6.73 $Y=0.83 $X2=0 $Y2=0
cc_450 N_S[3]_c_548_n N_VGND_c_1053_n 0.00349917f $X=7.72 $Y=0.905 $X2=0 $Y2=0
cc_451 N_S[3]_c_549_n N_VGND_c_1053_n 0.00880034f $X=7.795 $Y=0.83 $X2=0 $Y2=0
cc_452 N_A_1361_47#_M1005_g N_D[3]_c_644_n 0.0381613f $X=7.72 $Y=2.075 $X2=-0.19
+ $Y2=-0.24
cc_453 N_A_1361_47#_c_591_n N_D[3]_c_644_n 0.00712672f $X=7.415 $Y=1.34
+ $X2=-0.19 $Y2=-0.24
cc_454 N_A_1361_47#_c_594_n N_VPWR_c_677_n 0.0498301f $X=6.965 $Y=2.31 $X2=0
+ $Y2=0
cc_455 N_A_1361_47#_c_590_n N_VPWR_c_677_n 0.0110094f $X=7.195 $Y=1.405 $X2=0
+ $Y2=0
cc_456 N_A_1361_47#_M1005_g N_VPWR_c_679_n 0.00298082f $X=7.72 $Y=2.075 $X2=0
+ $Y2=0
cc_457 N_A_1361_47#_M1005_g N_VPWR_c_685_n 0.00522699f $X=7.72 $Y=2.075 $X2=0
+ $Y2=0
cc_458 N_A_1361_47#_c_594_n N_VPWR_c_685_n 0.0210596f $X=6.965 $Y=2.31 $X2=0
+ $Y2=0
cc_459 N_A_1361_47#_M1001_d N_VPWR_c_672_n 0.00179197f $X=6.82 $Y=1.485 $X2=0
+ $Y2=0
cc_460 N_A_1361_47#_M1005_g N_VPWR_c_672_n 0.00828927f $X=7.72 $Y=2.075 $X2=0
+ $Y2=0
cc_461 N_A_1361_47#_c_594_n N_VPWR_c_672_n 0.00594162f $X=6.965 $Y=2.31 $X2=0
+ $Y2=0
cc_462 N_A_1361_47#_M1005_g N_Z_c_822_n 0.00988241f $X=7.72 $Y=2.075 $X2=0 $Y2=0
cc_463 N_A_1361_47#_c_594_n N_Z_c_822_n 0.0369227f $X=6.965 $Y=2.31 $X2=0 $Y2=0
cc_464 N_A_1361_47#_c_589_n N_Z_c_812_n 0.00611965f $X=7.195 $Y=1.175 $X2=0
+ $Y2=0
cc_465 N_A_1361_47#_c_592_n N_Z_c_812_n 0.0259454f $X=6.965 $Y=0.495 $X2=0 $Y2=0
cc_466 N_A_1361_47#_M1005_g N_Z_c_813_n 0.00862328f $X=7.72 $Y=2.075 $X2=0 $Y2=0
cc_467 N_A_1361_47#_c_594_n N_Z_c_813_n 0.00378484f $X=6.965 $Y=2.31 $X2=0 $Y2=0
cc_468 N_A_1361_47#_c_589_n N_Z_c_813_n 0.00719188f $X=7.195 $Y=1.175 $X2=0
+ $Y2=0
cc_469 N_A_1361_47#_c_590_n N_Z_c_813_n 0.0304368f $X=7.195 $Y=1.405 $X2=0 $Y2=0
cc_470 N_A_1361_47#_c_591_n N_Z_c_813_n 0.00814206f $X=7.415 $Y=1.34 $X2=0 $Y2=0
cc_471 N_A_1361_47#_c_589_n N_Z_c_815_n 0.0124144f $X=7.195 $Y=1.175 $X2=0 $Y2=0
cc_472 N_A_1361_47#_c_590_n N_Z_c_815_n 0.00398133f $X=7.195 $Y=1.405 $X2=0
+ $Y2=0
cc_473 N_A_1361_47#_c_591_n N_Z_c_815_n 0.00349316f $X=7.415 $Y=1.34 $X2=0 $Y2=0
cc_474 N_A_1361_47#_c_594_n N_Z_c_825_n 0.0293762f $X=6.965 $Y=2.31 $X2=0 $Y2=0
cc_475 N_A_1361_47#_c_590_n N_Z_c_825_n 0.0126642f $X=7.195 $Y=1.405 $X2=0 $Y2=0
cc_476 N_A_1361_47#_M1005_g N_Z_c_957_n 0.00289142f $X=7.72 $Y=2.075 $X2=0 $Y2=0
cc_477 N_A_1361_47#_c_594_n N_Z_c_957_n 6.03258e-19 $X=6.965 $Y=2.31 $X2=0 $Y2=0
cc_478 N_A_1361_47#_c_590_n N_Z_c_957_n 4.25753e-19 $X=7.195 $Y=1.405 $X2=0
+ $Y2=0
cc_479 N_A_1361_47#_M1005_g N_Z_c_828_n 0.0105217f $X=7.72 $Y=2.075 $X2=0 $Y2=0
cc_480 N_A_1361_47#_c_594_n N_Z_c_828_n 0.0139746f $X=6.965 $Y=2.31 $X2=0 $Y2=0
cc_481 N_A_1361_47#_c_590_n N_Z_c_828_n 0.00749676f $X=7.195 $Y=1.405 $X2=0
+ $Y2=0
cc_482 N_A_1361_47#_c_591_n N_Z_c_828_n 0.00449162f $X=7.415 $Y=1.34 $X2=0 $Y2=0
cc_483 N_A_1361_47#_c_592_n N_VGND_c_1051_n 0.015238f $X=6.965 $Y=0.495 $X2=0
+ $Y2=0
cc_484 N_A_1361_47#_M1015_d N_VGND_c_1053_n 0.00358139f $X=6.805 $Y=0.235 $X2=0
+ $Y2=0
cc_485 N_A_1361_47#_c_592_n N_VGND_c_1053_n 0.0150148f $X=6.965 $Y=0.495 $X2=0
+ $Y2=0
cc_486 N_D[3]_c_644_n N_VPWR_c_679_n 0.0245615f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_487 N_D[3]_c_647_n N_VPWR_c_679_n 0.00471543f $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_488 N_D[3]_c_644_n N_VPWR_c_685_n 0.00622633f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_489 N_D[3]_c_644_n N_VPWR_c_672_n 0.0106352f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_490 N_D[3]_c_644_n N_Z_c_822_n 0.00145364f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_491 N_D[3]_c_646_n N_Z_c_812_n 0.00686805f $X=8.095 $Y=1.055 $X2=0 $Y2=0
cc_492 N_D[3]_c_644_n N_Z_c_813_n 0.00605747f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_493 N_D[3]_c_646_n N_Z_c_813_n 0.00376465f $X=8.095 $Y=1.055 $X2=0 $Y2=0
cc_494 N_D[3]_c_647_n N_Z_c_813_n 0.0216525f $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_495 N_D[3]_c_646_n N_Z_c_815_n 0.0128881f $X=8.095 $Y=1.055 $X2=0 $Y2=0
cc_496 N_D[3]_c_645_n N_VGND_c_1045_n 0.00487865f $X=8.27 $Y=0.995 $X2=0 $Y2=0
cc_497 N_D[3]_c_647_n N_VGND_c_1045_n 0.00222881f $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_498 N_D[3]_c_645_n N_VGND_c_1051_n 0.00585385f $X=8.27 $Y=0.995 $X2=0 $Y2=0
cc_499 N_D[3]_c_667_p N_VGND_c_1051_n 0.00842546f $X=8.095 $Y=0.51 $X2=0 $Y2=0
cc_500 N_D[3]_c_645_n N_VGND_c_1053_n 0.011617f $X=8.27 $Y=0.995 $X2=0 $Y2=0
cc_501 N_D[3]_c_667_p N_VGND_c_1053_n 0.00942277f $X=8.095 $Y=0.51 $X2=0 $Y2=0
cc_502 N_D[3]_c_646_n A_1574_47# 0.00426617f $X=8.095 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_503 N_D[3]_c_667_p A_1574_47# 0.00894235f $X=8.095 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_504 N_VPWR_c_672_n A_117_297# 0.0138589f $X=8.51 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_505 N_VPWR_c_672_n N_Z_M1009_d 0.00174926f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_506 N_VPWR_c_672_n N_Z_M1003_s 0.00174926f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_507 N_VPWR_c_672_n N_Z_M1012_d 0.00174926f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_508 N_VPWR_c_672_n N_Z_M1005_s 0.00174926f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_509 N_VPWR_c_674_n N_Z_c_804_n 0.00734981f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_510 N_VPWR_c_674_n N_Z_c_817_n 0.0115091f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_511 N_VPWR_c_680_n N_Z_c_817_n 0.0210727f $X=2.165 $Y=2.72 $X2=0 $Y2=0
cc_512 N_VPWR_c_672_n N_Z_c_817_n 0.00577491f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_513 N_VPWR_c_676_n N_Z_c_818_n 0.0116583f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_514 N_VPWR_c_684_n N_Z_c_818_n 0.0210727f $X=4.175 $Y=2.72 $X2=0 $Y2=0
cc_515 N_VPWR_c_672_n N_Z_c_818_n 0.00577491f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_516 N_VPWR_c_676_n N_Z_c_808_n 0.0074594f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_517 N_VPWR_c_676_n N_Z_c_809_n 0.0074594f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_518 N_VPWR_c_676_n N_Z_c_821_n 0.0116583f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_519 N_VPWR_c_682_n N_Z_c_821_n 0.0210727f $X=6.275 $Y=2.72 $X2=0 $Y2=0
cc_520 N_VPWR_c_672_n N_Z_c_821_n 0.00577491f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_521 N_VPWR_c_679_n N_Z_c_822_n 0.0115091f $X=8.48 $Y=1.66 $X2=0 $Y2=0
cc_522 N_VPWR_c_685_n N_Z_c_822_n 0.0210727f $X=8.315 $Y=2.72 $X2=0 $Y2=0
cc_523 N_VPWR_c_672_n N_Z_c_822_n 0.00577491f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_524 N_VPWR_c_679_n N_Z_c_813_n 0.00734981f $X=8.48 $Y=1.66 $X2=0 $Y2=0
cc_525 N_VPWR_M1013_d N_Z_c_824_n 0.00291605f $X=2.1 $Y=1.485 $X2=0 $Y2=0
cc_526 N_VPWR_c_675_n N_Z_c_824_n 0.0300023f $X=2.3 $Y=1.63 $X2=0 $Y2=0
cc_527 N_VPWR_c_672_n N_Z_c_824_n 0.0951133f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_528 N_VPWR_c_674_n N_Z_c_850_n 0.00119119f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_529 N_VPWR_c_672_n N_Z_c_850_n 0.0144722f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_530 N_VPWR_c_676_n N_Z_c_897_n 0.0355595f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_531 N_VPWR_c_672_n N_Z_c_897_n 0.0739714f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_532 N_VPWR_c_676_n N_Z_c_884_n 4.83404e-19 $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_533 N_VPWR_c_672_n N_Z_c_884_n 0.0144722f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_534 N_VPWR_M1014_d N_Z_c_825_n 0.00291605f $X=6.24 $Y=1.485 $X2=0 $Y2=0
cc_535 N_VPWR_c_677_n N_Z_c_825_n 0.0300023f $X=6.44 $Y=1.63 $X2=0 $Y2=0
cc_536 N_VPWR_c_672_n N_Z_c_825_n 0.0951133f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_537 N_VPWR_c_676_n N_Z_c_923_n 4.83404e-19 $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_538 N_VPWR_c_672_n N_Z_c_923_n 0.0144722f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_539 N_VPWR_c_676_n N_Z_c_826_n 0.00305596f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_540 N_VPWR_c_684_n N_Z_c_826_n 0.00233997f $X=4.175 $Y=2.72 $X2=0 $Y2=0
cc_541 N_VPWR_c_672_n N_Z_c_826_n 0.00180522f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_542 N_VPWR_c_676_n N_Z_c_827_n 0.00305596f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_543 N_VPWR_c_682_n N_Z_c_827_n 0.00233997f $X=6.275 $Y=2.72 $X2=0 $Y2=0
cc_544 N_VPWR_c_672_n N_Z_c_827_n 0.00180522f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_545 N_VPWR_c_679_n N_Z_c_957_n 0.00119119f $X=8.48 $Y=1.66 $X2=0 $Y2=0
cc_546 N_VPWR_c_672_n N_Z_c_957_n 0.0144722f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_547 N_VPWR_c_685_n N_Z_c_828_n 0.00233997f $X=8.315 $Y=2.72 $X2=0 $Y2=0
cc_548 N_VPWR_c_672_n N_Z_c_828_n 0.00317613f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_549 N_VPWR_c_680_n N_Z_c_829_n 0.00233997f $X=2.165 $Y=2.72 $X2=0 $Y2=0
cc_550 N_VPWR_c_672_n N_Z_c_829_n 0.00317613f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_551 N_VPWR_c_672_n A_734_333# 0.00481681f $X=8.51 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_552 N_VPWR_c_672_n A_945_297# 0.00481681f $X=8.51 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_553 N_VPWR_c_672_n A_1562_333# 0.0138589f $X=8.51 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_554 N_VPWR_c_674_n N_VGND_c_1040_n 0.00704239f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_555 N_VPWR_c_676_n N_VGND_c_1042_n 0.00723368f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_556 N_VPWR_c_679_n N_VGND_c_1045_n 0.00704239f $X=8.48 $Y=1.66 $X2=0 $Y2=0
cc_557 N_Z_c_897_n A_734_333# 0.0127078f $X=5.145 $Y=1.87 $X2=-0.19 $Y2=-0.24
cc_558 N_Z_c_897_n A_945_297# 0.0127078f $X=5.145 $Y=1.87 $X2=-0.19 $Y2=-0.24
cc_559 N_Z_c_806_n N_VGND_c_1046_n 0.0106022f $X=1.155 $Y=0.495 $X2=0 $Y2=0
cc_560 N_Z_c_811_n N_VGND_c_1048_n 0.0106022f $X=5.295 $Y=0.495 $X2=0 $Y2=0
cc_561 N_Z_c_807_n N_VGND_c_1050_n 0.0106022f $X=3.445 $Y=0.495 $X2=0 $Y2=0
cc_562 N_Z_c_812_n N_VGND_c_1051_n 0.0106022f $X=7.585 $Y=0.495 $X2=0 $Y2=0
cc_563 N_Z_M1023_d N_VGND_c_1053_n 0.00232956f $X=1.02 $Y=0.235 $X2=0 $Y2=0
cc_564 N_Z_M1006_s N_VGND_c_1053_n 0.00232956f $X=3.32 $Y=0.235 $X2=0 $Y2=0
cc_565 N_Z_M1004_d N_VGND_c_1053_n 0.00232956f $X=5.16 $Y=0.235 $X2=0 $Y2=0
cc_566 N_Z_M1002_s N_VGND_c_1053_n 0.00232956f $X=7.46 $Y=0.235 $X2=0 $Y2=0
cc_567 N_Z_c_805_n N_VGND_c_1053_n 0.00409585f $X=1.167 $Y=0.835 $X2=0 $Y2=0
cc_568 N_Z_c_806_n N_VGND_c_1053_n 0.00891193f $X=1.155 $Y=0.495 $X2=0 $Y2=0
cc_569 N_Z_c_807_n N_VGND_c_1053_n 0.00891193f $X=3.445 $Y=0.495 $X2=0 $Y2=0
cc_570 N_Z_c_810_n N_VGND_c_1053_n 0.00409585f $X=5.307 $Y=0.835 $X2=0 $Y2=0
cc_571 N_Z_c_811_n N_VGND_c_1053_n 0.00891193f $X=5.295 $Y=0.495 $X2=0 $Y2=0
cc_572 N_Z_c_812_n N_VGND_c_1053_n 0.00891193f $X=7.585 $Y=0.495 $X2=0 $Y2=0
cc_573 N_Z_c_814_n N_VGND_c_1053_n 0.00409585f $X=3.615 $Y=0.92 $X2=0 $Y2=0
cc_574 N_Z_c_815_n N_VGND_c_1053_n 0.00409585f $X=7.755 $Y=0.92 $X2=0 $Y2=0
cc_575 N_VGND_c_1053_n A_109_47# 0.00453173f $X=8.51 $Y=0 $X2=-0.19 $Y2=-0.24
cc_576 N_VGND_c_1053_n A_746_47# 0.00453173f $X=8.51 $Y=0 $X2=-0.19 $Y2=-0.24
cc_577 N_VGND_c_1053_n A_937_47# 0.00453173f $X=8.51 $Y=0 $X2=-0.19 $Y2=-0.24
cc_578 N_VGND_c_1053_n A_1574_47# 0.00453173f $X=8.51 $Y=0 $X2=-0.19 $Y2=-0.24
