* NGSPICE file created from sky130_fd_sc_hdll__dlygate4sd2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__dlygate4sd2_1 A VGND VNB VPB VPWR X
M1000 a_213_47# a_27_47# VGND VNB nshort w=420000u l=180000u
+  ad=1.092e+11p pd=1.36e+06u as=4.913e+11p ps=3.91e+06u
M1001 X a_319_93# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1002 VPWR a_213_47# a_319_93# VPB phighvt w=420000u l=180000u
+  ad=6.233e+11p pd=4.51e+06u as=1.176e+11p ps=1.4e+06u
M1003 X a_319_93# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1004 a_213_47# a_27_47# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1005 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1006 VGND a_213_47# a_319_93# VNB nshort w=420000u l=180000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1007 VPWR A a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
.ends

