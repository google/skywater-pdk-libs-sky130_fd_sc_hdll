* File: sky130_fd_sc_hdll__and2_4.spice
* Created: Thu Aug 27 18:56:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and2_4.pex.spice"
.subckt sky130_fd_sc_hdll__and2_4  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 A_120_47# N_A_M1002_g N_A_27_47#_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.20475 PD=0.86 PS=1.93 NRD=9.228 NRS=9.228 M=1 R=4.33333
+ SA=75000.2 SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_B_M1009_g A_120_47# VNB NSHORT L=0.15 W=0.65 AD=0.154375
+ AS=0.06825 PD=1.125 PS=0.86 NRD=22.152 NRS=9.228 M=1 R=4.33333 SA=75000.6
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1009_d N_A_27_47#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.154375 AS=0.10725 PD=1.125 PS=0.98 NRD=13.836 NRS=9.228 M=1 R=4.33333
+ SA=75001.2 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_A_27_47#_M1003_g N_X_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1003_d N_A_27_47#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.1235 PD=0.98 PS=1.03 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75002.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1010_d N_A_27_47#_M1010_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.18525 AS=0.1235 PD=1.87 PS=1.03 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75002.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_27_47#_M1004_d N_A_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90002.7 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_B_M1008_g N_A_27_47#_M1004_d VPB PHIGHVT L=0.18 W=1
+ AD=0.1875 AS=0.15 PD=1.375 PS=1.3 NRD=8.8453 NRS=1.9503 M=1 R=5.55556
+ SA=90000.7 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1000 N_X_M1000_d N_A_27_47#_M1000_g N_VPWR_M1008_d VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.1875 PD=1.3 PS=1.375 NRD=1.9503 NRS=9.8303 M=1 R=5.55556
+ SA=90001.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1005 N_X_M1000_d N_A_27_47#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.7
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1006 N_X_M1006_d N_A_27_47#_M1006_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.2
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1011 N_X_M1006_d N_A_27_47#_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hdll__and2_4.pxi.spice"
*
.ends
*
*
