# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__clkbuf_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.243000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.755000 0.825000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.898200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.345000 1.405000 0.735000 ;
        RECT 1.050000 0.735000 2.910000 0.905000 ;
        RECT 1.145000 1.835000 2.365000 2.005000 ;
        RECT 1.145000 2.005000 1.405000 2.465000 ;
        RECT 2.105000 0.345000 2.365000 0.735000 ;
        RECT 2.105000 1.415000 2.910000 1.650000 ;
        RECT 2.105000 1.650000 2.365000 1.835000 ;
        RECT 2.105000 2.005000 2.365000 2.465000 ;
        RECT 2.410000 0.905000 2.910000 1.415000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.255000 0.385000 0.585000 ;
      RECT 0.085000  0.585000 0.255000 1.495000 ;
      RECT 0.085000  1.495000 1.215000 1.665000 ;
      RECT 0.085000  1.665000 0.395000 2.465000 ;
      RECT 0.605000  0.085000 0.880000 0.565000 ;
      RECT 0.615000  1.835000 0.925000 2.635000 ;
      RECT 0.995000  1.075000 2.240000 1.245000 ;
      RECT 0.995000  1.245000 1.215000 1.495000 ;
      RECT 1.625000  0.085000 1.880000 0.565000 ;
      RECT 1.625000  2.175000 1.880000 2.635000 ;
      RECT 2.545000  1.845000 2.875000 2.635000 ;
      RECT 2.585000  0.085000 2.865000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkbuf_4
END LIBRARY
