* File: sky130_fd_sc_hdll__or3b_2.pex.spice
* Created: Wed Sep  2 08:48:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR3B_2%C_N 2 3 5 8 10 11 19
c32 19 0 1.20913e-19 $X=0.52 $Y=1.16
r33 18 19 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r34 15 18 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.495 $Y2=1.16
r35 10 11 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.16
+ $X2=0.255 $Y2=1.53
r36 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r37 6 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.16
r38 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r39 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.725
+ $X2=0.495 $Y2=2.01
r40 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.625 $X2=0.495
+ $Y2=1.725
r41 1 18 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r42 1 2 99.4732 $w=2e-07 $l=3e-07 $layer=POLY_cond $X=0.495 $Y=1.325 $X2=0.495
+ $Y2=1.625
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_2%A_186_21# 1 2 3 10 12 13 15 16 18 20 21 23
+ 24 27 30 31 34 36 40 43 44 45 49
c103 31 0 1.58571e-19 $X=1.655 $Y=0.82
c104 13 0 1.43265e-20 $X=1.03 $Y=1.41
r105 47 49 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.325 $Y=1.71
+ $X2=3.46 $Y2=1.71
r106 43 49 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=3.46 $Y=1.495
+ $X2=3.46 $Y2=1.71
r107 42 45 3.87901 $w=2.37e-07 $l=1.14039e-07 $layer=LI1_cond $X=3.46 $Y=0.825
+ $X2=3.392 $Y2=0.74
r108 42 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.46 $Y=0.825
+ $X2=3.46 $Y2=1.495
r109 38 45 3.87901 $w=2.37e-07 $l=8.5e-08 $layer=LI1_cond $X=3.392 $Y=0.655
+ $X2=3.392 $Y2=0.74
r110 38 40 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=3.392 $Y=0.655
+ $X2=3.392 $Y2=0.47
r111 37 44 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=2.535 $Y=0.74
+ $X2=2.45 $Y2=0.78
r112 36 45 2.57001 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.24 $Y=0.74
+ $X2=3.392 $Y2=0.74
r113 36 37 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=3.24 $Y=0.74
+ $X2=2.535 $Y2=0.74
r114 32 44 1.34256 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.45 $Y=0.655
+ $X2=2.45 $Y2=0.78
r115 32 34 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.45 $Y=0.655
+ $X2=2.45 $Y2=0.47
r116 30 44 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=2.365 $Y=0.82
+ $X2=2.45 $Y2=0.78
r117 30 31 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.365 $Y=0.82
+ $X2=1.655 $Y2=0.82
r118 25 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.57 $Y=0.905
+ $X2=1.655 $Y2=0.82
r119 25 27 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.57 $Y=0.905
+ $X2=1.57 $Y2=1.16
r120 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.68 $Y=0.995
+ $X2=1.68 $Y2=0.56
r121 18 20 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.61 $Y=1.41
+ $X2=1.61 $Y2=1.985
r122 17 24 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.13 $Y=1.16
+ $X2=1.03 $Y2=1.202
r123 16 18 54.0377 $w=2.35e-07 $l=2.60768e-07 $layer=POLY_cond $X=1.632 $Y=1.16
+ $X2=1.61 $Y2=1.41
r124 16 21 40.1263 $w=2.35e-07 $l=1.8747e-07 $layer=POLY_cond $X=1.632 $Y=1.16
+ $X2=1.68 $Y2=0.995
r125 16 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.57
+ $Y=1.16 $X2=1.57 $Y2=1.16
r126 16 17 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=1.51 $Y=1.16
+ $X2=1.13 $Y2=1.16
r127 13 24 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.03 $Y2=1.202
r128 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.03 $Y2=1.985
r129 10 24 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.03 $Y2=1.202
r130 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=0.56
r131 3 47 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=3.18
+ $Y=1.485 $X2=3.325 $Y2=1.685
r132 2 40 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=3.19
+ $Y=0.265 $X2=3.325 $Y2=0.47
r133 1 34 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=2.31
+ $Y=0.265 $X2=2.45 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_2%A 1 3 6 8 9
r36 8 9 7.56494 $w=5.83e-07 $l=3.7e-07 $layer=LI1_cond $X=2.247 $Y=1.16
+ $X2=2.247 $Y2=1.53
r37 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.125
+ $Y=1.16 $X2=2.125 $Y2=1.16
r38 4 13 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.235 $Y=0.995
+ $X2=2.15 $Y2=1.16
r39 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.235 $Y=0.995
+ $X2=2.235 $Y2=0.475
r40 1 13 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=2.15 $Y=1.41
+ $X2=2.15 $Y2=1.16
r41 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.15 $Y=1.41 $X2=2.15
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_2%B 1 2 4 7 10 11 20
r37 16 20 13.4452 $w=2.38e-07 $l=2.8e-07 $layer=LI1_cond $X=2.595 $Y=2.245
+ $X2=2.875 $Y2=2.245
r38 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.595
+ $Y=2.28 $X2=2.595 $Y2=2.28
r39 10 11 19.9277 $w=2.38e-07 $l=4.15e-07 $layer=LI1_cond $X=2.99 $Y=2.245
+ $X2=3.405 $Y2=2.245
r40 10 20 5.52212 $w=2.38e-07 $l=1.15e-07 $layer=LI1_cond $X=2.99 $Y=2.245
+ $X2=2.875 $Y2=2.245
r41 7 9 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.665 $Y=0.475
+ $X2=2.665 $Y2=1.11
r42 2 15 45.7813 $w=3.27e-07 $l=2.54804e-07 $layer=POLY_cond $X=2.64 $Y=2.035
+ $X2=2.62 $Y2=2.28
r43 2 4 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=2.64 $Y=2.035 $X2=2.64
+ $Y2=1.695
r44 1 9 118.763 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=2.64 $Y=1.41 $X2=2.64
+ $Y2=1.11
r45 1 4 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.64 $Y=1.41 $X2=2.64
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_2%A_27_47# 1 2 7 9 12 16 18 19 20 23 26 29 32
+ 34 35 36 40
c102 32 0 1.43265e-20 $X=0.26 $Y=1.975
c103 20 0 1.20913e-19 $X=0.645 $Y=1.925
r104 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.085
+ $Y=1.16 $X2=3.085 $Y2=1.16
r105 37 40 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.935 $Y=1.16
+ $X2=3.085 $Y2=1.16
r106 35 36 7.68295 $w=2.53e-07 $l=1.7e-07 $layer=LI1_cond $X=1.81 $Y=1.912
+ $X2=1.98 $Y2=1.912
r107 28 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.935 $Y=1.325
+ $X2=2.935 $Y2=1.16
r108 28 29 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.935 $Y=1.325
+ $X2=2.935 $Y2=1.785
r109 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.85 $Y=1.87
+ $X2=2.935 $Y2=1.785
r110 26 36 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=2.85 $Y=1.87
+ $X2=1.98 $Y2=1.87
r111 25 34 4.50329 $w=2e-07 $l=9.88686e-08 $layer=LI1_cond $X=0.815 $Y=1.955
+ $X2=0.73 $Y2=1.925
r112 25 35 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=0.815 $Y=1.955
+ $X2=1.81 $Y2=1.955
r113 23 34 1.93381 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.73 $Y=1.81
+ $X2=0.73 $Y2=1.925
r114 22 23 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=0.73 $Y=0.905
+ $X2=0.73 $Y2=1.81
r115 21 32 1.45362 $w=2.3e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.925
+ $X2=0.215 $Y2=1.925
r116 20 34 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.645 $Y=1.925
+ $X2=0.73 $Y2=1.925
r117 20 21 15.0319 $w=2.28e-07 $l=3e-07 $layer=LI1_cond $X=0.645 $Y=1.925
+ $X2=0.345 $Y2=1.925
r118 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.645 $Y=0.82
+ $X2=0.73 $Y2=0.905
r119 18 19 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.645 $Y=0.82
+ $X2=0.345 $Y2=0.82
r120 14 19 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.735
+ $X2=0.345 $Y2=0.82
r121 14 16 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=0.215 $Y=0.735
+ $X2=0.215 $Y2=0.455
r122 10 41 38.7444 $w=2.79e-07 $l=1.72337e-07 $layer=POLY_cond $X=3.115 $Y=0.995
+ $X2=3.1 $Y2=1.16
r123 10 12 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=3.115 $Y=0.995
+ $X2=3.115 $Y2=0.475
r124 7 41 49.2447 $w=2.79e-07 $l=2.54951e-07 $layer=POLY_cond $X=3.09 $Y=1.41
+ $X2=3.1 $Y2=1.16
r125 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.09 $Y=1.41
+ $X2=3.09 $Y2=1.695
r126 2 32 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.8 $X2=0.26 $Y2=1.975
r127 1 16 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_2%VPWR 1 2 9 13 16 17 18 20 33 34 37
r48 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r49 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r50 31 34 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r51 30 33 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r52 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r53 28 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r54 28 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r55 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r56 25 37 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.96 $Y=2.72 $X2=0.78
+ $Y2=2.72
r57 25 27 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=0.96 $Y=2.72
+ $X2=1.61 $Y2=2.72
r58 20 37 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.6 $Y=2.72 $X2=0.78
+ $Y2=2.72
r59 20 22 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.6 $Y=2.72 $X2=0.23
+ $Y2=2.72
r60 18 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r62 16 27 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=1.685 $Y=2.72
+ $X2=1.61 $Y2=2.72
r63 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=2.72
+ $X2=1.85 $Y2=2.72
r64 15 30 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.015 $Y=2.72
+ $X2=2.07 $Y2=2.72
r65 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=2.72
+ $X2=1.85 $Y2=2.72
r66 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.85 $Y=2.635
+ $X2=1.85 $Y2=2.72
r67 11 13 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.85 $Y=2.635
+ $X2=1.85 $Y2=2.295
r68 7 37 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=2.635 $X2=0.78
+ $Y2=2.72
r69 7 9 10.8842 $w=3.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.78 $Y=2.635 $X2=0.78
+ $Y2=2.295
r70 2 13 600 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=1.7
+ $Y=1.485 $X2=1.85 $Y2=2.295
r71 1 9 600 $w=1.7e-07 $l=5.90741e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.8 $X2=0.795 $Y2=2.295
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_2%X 1 2 8 11 13 21
r32 18 21 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=1.11 $Y=0.43
+ $X2=1.155 $Y2=0.43
r33 13 21 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.255 $Y=0.43
+ $X2=1.155 $Y2=0.43
r34 13 18 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=1.11 $Y=0.595
+ $X2=1.11 $Y2=0.43
r35 8 13 33.4503 $w=3.13e-07 $l=9e-07 $layer=LI1_cond $X=1.11 $Y=1.495 $X2=1.11
+ $Y2=0.595
r36 8 11 8.38581 $w=2.03e-07 $l=1.55e-07 $layer=LI1_cond $X=1.11 $Y=1.597
+ $X2=1.265 $Y2=1.597
r37 2 11 600 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.485 $X2=1.265 $Y2=1.615
r38 1 13 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.235 $X2=1.265 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_2%VGND 1 2 3 14 18 22 25 26 28 29 30 40 41 44
r56 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r57 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r58 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r59 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r60 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r61 35 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r62 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r63 32 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.73
+ $Y2=0
r64 32 34 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=1.61
+ $Y2=0
r65 30 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r66 28 37 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.74 $Y=0 $X2=2.53
+ $Y2=0
r67 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.74 $Y=0 $X2=2.905
+ $Y2=0
r68 27 40 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.07 $Y=0 $X2=3.45
+ $Y2=0
r69 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.07 $Y=0 $X2=2.905
+ $Y2=0
r70 25 34 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.61
+ $Y2=0
r71 25 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.95
+ $Y2=0
r72 24 37 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=2.53
+ $Y2=0
r73 24 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.035 $Y=0 $X2=1.95
+ $Y2=0
r74 20 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.905 $Y=0.085
+ $X2=2.905 $Y2=0
r75 20 22 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.905 $Y=0.085
+ $X2=2.905 $Y2=0.4
r76 16 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=0.085
+ $X2=1.95 $Y2=0
r77 16 18 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.95 $Y=0.085
+ $X2=1.95 $Y2=0.4
r78 12 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r79 12 14 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.4
r80 3 22 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.74
+ $Y=0.265 $X2=2.905 $Y2=0.4
r81 2 18 182 $w=1.7e-07 $l=2.64953e-07 $layer=licon1_NDIFF $count=1 $X=1.755
+ $Y=0.235 $X2=1.95 $Y2=0.4
r82 1 14 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.4
.ends

