* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__sedfxbp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 a_1787_159# a_1611_413# VPWR VPB phighvt w=750000u l=180000u
+  ad=2.025e+11p pd=2.04e+06u as=1.93535e+12p ps=1.705e+07u
M1001 Q a_2266_413# VGND VNB nshort w=650000u l=150000u
+  ad=1.9825e+11p pd=1.91e+06u as=1.4487e+12p ps=1.404e+07u
M1002 a_211_363# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1003 a_2165_413# a_1787_159# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.365e+11p pd=1.49e+06u as=0p ps=0u
M1004 a_2266_413# a_27_47# a_2165_413# VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
M1005 VPWR DE a_455_324# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1006 VPWR CLK a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1007 a_319_47# a_851_264# a_779_47# VNB nshort w=420000u l=150000u
+  ad=2.478e+11p pd=2.86e+06u as=1.932e+11p ps=1.76e+06u
M1008 a_2181_47# a_1787_159# VGND VNB nshort w=420000u l=150000u
+  ad=1.356e+11p pd=1.51e+06u as=0p ps=0u
M1009 Q a_2266_413# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.15e+11p pd=2.63e+06u as=0p ps=0u
M1010 a_2266_413# a_211_363# a_2181_47# VNB nshort w=360000u l=150000u
+  ad=1.494e+11p pd=1.55e+06u as=0p ps=0u
M1011 a_1611_413# a_27_47# a_985_47# VNB nshort w=360000u l=150000u
+  ad=1.404e+11p pd=1.5e+06u as=6.015e+11p ps=4.57e+06u
M1012 a_985_47# a_955_21# a_1376_369# VPB phighvt w=640000u l=180000u
+  ad=4.837e+11p pd=4.13e+06u as=2.24e+11p ps=1.98e+06u
M1013 VGND SCE a_955_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1014 VGND a_2266_413# a_851_264# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1015 a_985_47# a_955_21# a_319_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Q_N a_851_264# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1017 VPWR SCE a_955_21# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.76e+11p ps=1.83e+06u
M1018 a_409_369# D a_319_47# VPB phighvt w=640000u l=180000u
+  ad=1.472e+11p pd=1.74e+06u as=3.84e+11p ps=3.76e+06u
M1019 a_985_47# SCE a_1373_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1020 VGND a_851_264# a_2391_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.32e+11p ps=1.49e+06u
M1021 a_787_369# DE VPWR VPB phighvt w=640000u l=180000u
+  ad=2.432e+11p pd=2.04e+06u as=0p ps=0u
M1022 a_319_47# a_851_264# a_787_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1611_413# a_211_363# a_985_47# VPB phighvt w=420000u l=180000u
+  ad=1.365e+11p pd=1.49e+06u as=0p ps=0u
M1024 VPWR a_1787_159# a_1712_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.617e+11p ps=1.61e+06u
M1025 VPWR a_455_324# a_409_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_985_47# SCE a_319_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Q_N a_851_264# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1028 a_1712_413# a_27_47# a_1611_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_2266_413# a_851_264# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1030 VGND DE a_455_324# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1031 a_779_47# a_455_324# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1376_369# SCD VPWR VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1034 a_1373_119# SCD VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR a_851_264# a_2360_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=2.058e+11p ps=1.82e+06u
M1036 VGND a_1787_159# a_1738_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.518e+11p ps=1.6e+06u
M1037 a_211_363# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1038 a_1738_47# a_211_363# a_1611_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_2391_47# a_27_47# a_2266_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_413_47# D a_319_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1041 VGND DE a_413_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_2360_413# a_211_363# a_2266_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_1787_159# a_1611_413# VGND VNB nshort w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=0p ps=0u
.ends
