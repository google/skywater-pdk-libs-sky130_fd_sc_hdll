* File: sky130_fd_sc_hdll__o2bb2a_1.pex.spice
* Created: Thu Aug 27 19:21:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_1%A_76_199# 1 2 7 9 10 12 15 19 20 21 25 28
+ 31 34 35 36
c98 7 0 1.12461e-19 $X=0.495 $Y=1.41
r99 36 38 2.04089 $w=5.38e-07 $l=9e-08 $layer=LI1_cond $X=2.632 $Y=1.97
+ $X2=2.632 $Y2=2.06
r100 34 35 9.669 $w=1.93e-07 $l=1.7e-07 $layer=LI1_cond $X=2.402 $Y=1.075
+ $X2=2.402 $Y2=1.245
r101 33 34 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.39 $Y=0.69
+ $X2=2.39 $Y2=1.075
r102 31 33 10.6372 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=2.35 $Y=0.485
+ $X2=2.35 $Y2=0.69
r103 25 36 16.98 $w=5.38e-07 $l=5.73324e-07 $layer=LI1_cond $X=2.415 $Y=1.495
+ $X2=2.632 $Y2=1.97
r104 25 35 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.415 $Y=1.495
+ $X2=2.415 $Y2=1.245
r105 20 36 7.61904 $w=1.7e-07 $l=3.02e-07 $layer=LI1_cond $X=2.33 $Y=1.97
+ $X2=2.632 $Y2=1.97
r106 20 21 94.9251 $w=1.68e-07 $l=1.455e-06 $layer=LI1_cond $X=2.33 $Y=1.97
+ $X2=0.875 $Y2=1.97
r107 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.79 $Y=1.885
+ $X2=0.875 $Y2=1.97
r108 18 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=1.615
+ $X2=0.79 $Y2=1.53
r109 18 19 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.79 $Y=1.615
+ $X2=0.79 $Y2=1.885
r110 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.16 $X2=0.515 $Y2=1.16
r111 13 28 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.54 $Y=1.53
+ $X2=0.79 $Y2=1.53
r112 13 15 14.9294 $w=2.18e-07 $l=2.85e-07 $layer=LI1_cond $X=0.54 $Y=1.445
+ $X2=0.54 $Y2=1.16
r113 10 16 38.578 $w=2.95e-07 $l=1.74714e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.54 $Y2=1.16
r114 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=0.56
r115 7 16 48.1208 $w=2.95e-07 $l=2.7157e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.54 $Y2=1.16
r116 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r117 2 38 600 $w=1.7e-07 $l=2.82046e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=1.845 $X2=2.79 $Y2=2.06
r118 1 31 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=2.185
+ $Y=0.235 $X2=2.31 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_1%A1_N 2 3 5 8 10 13 21
c45 21 0 1.56868e-19 $X=1.155 $Y=1.19
c46 8 0 1.42981e-19 $X=1.05 $Y=0.445
r47 13 16 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.07 $Y=1.16
+ $X2=1.07 $Y2=1.325
r48 13 15 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.07 $Y=1.16
+ $X2=1.07 $Y2=0.995
r49 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.045
+ $Y=1.16 $X2=1.045 $Y2=1.16
r50 10 21 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=1.14 $Y=1.175
+ $X2=1.155 $Y2=1.175
r51 10 14 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=1.14 $Y=1.175
+ $X2=1.045 $Y2=1.175
r52 8 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.05 $Y=0.445
+ $X2=1.05 $Y2=0.995
r53 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.03 $Y=1.77 $X2=1.03
+ $Y2=2.055
r54 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.03 $Y=1.67 $X2=1.03
+ $Y2=1.77
r55 2 16 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=1.03 $Y=1.67 $X2=1.03
+ $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_1%A2_N 3 5 6 8 9 10 16 18 21
c53 16 0 1.56868e-19 $X=1.575 $Y=0.935
r54 16 22 37.7065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=0.935
+ $X2=1.61 $Y2=1.1
r55 16 21 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=0.935
+ $X2=1.61 $Y2=0.77
r56 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.575
+ $Y=0.935 $X2=1.575 $Y2=0.935
r57 11 18 9.09823 $w=2.83e-07 $l=2.25e-07 $layer=LI1_cond $X=1.157 $Y=0.735
+ $X2=1.157 $Y2=0.51
r58 10 11 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=1.3 $Y=0.82
+ $X2=1.157 $Y2=0.735
r59 9 15 5.89026 $w=2.23e-07 $l=1.15e-07 $layer=LI1_cond $X=1.602 $Y=0.82
+ $X2=1.602 $Y2=0.935
r60 9 10 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.49 $Y=0.82 $X2=1.3
+ $Y2=0.82
r61 6 8 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.63 $Y=1.77 $X2=1.63
+ $Y2=2.055
r62 5 6 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.63 $Y=1.67 $X2=1.63
+ $Y2=1.77
r63 5 22 188.999 $w=2e-07 $l=5.7e-07 $layer=POLY_cond $X=1.63 $Y=1.67 $X2=1.63
+ $Y2=1.1
r64 3 21 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=1.515 $Y=0.445
+ $X2=1.515 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_1%A_224_369# 1 2 7 9 12 14 15 16 20 27 29
c70 20 0 1.42981e-19 $X=1.885 $Y=0.48
c71 16 0 1.12461e-19 $X=1.885 $Y=1.605
r72 27 29 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=2.022 $Y=1.52
+ $X2=2.022 $Y2=1.355
r73 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.075
+ $Y=1.52 $X2=2.075 $Y2=1.52
r74 24 29 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.97 $Y=0.565
+ $X2=1.97 $Y2=1.355
r75 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.885 $Y=0.48
+ $X2=1.97 $Y2=0.565
r76 20 22 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.885 $Y=0.48
+ $X2=1.775 $Y2=0.48
r77 16 27 3.5621 $w=2.73e-07 $l=8.5e-08 $layer=LI1_cond $X=2.022 $Y=1.605
+ $X2=2.022 $Y2=1.52
r78 16 18 29.073 $w=2.18e-07 $l=5.55e-07 $layer=LI1_cond $X=1.885 $Y=1.605
+ $X2=1.33 $Y2=1.605
r79 14 28 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=2.445 $Y=1.52
+ $X2=2.075 $Y2=1.52
r80 14 15 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=2.445 $Y=1.52
+ $X2=2.545 $Y2=1.562
r81 10 15 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=2.57 $Y=1.355
+ $X2=2.545 $Y2=1.562
r82 10 12 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=2.57 $Y=1.355
+ $X2=2.57 $Y2=0.445
r83 7 15 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=2.545 $Y=1.77
+ $X2=2.545 $Y2=1.562
r84 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.545 $Y=1.77
+ $X2=2.545 $Y2=2.055
r85 2 18 600 $w=1.7e-07 $l=3.02283e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.845 $X2=1.33 $Y2=1.63
r86 1 22 182 $w=1.7e-07 $l=3.24577e-07 $layer=licon1_NDIFF $count=1 $X=1.59
+ $Y=0.235 $X2=1.775 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_1%B2 3 6 7 9 10 13 15 17 18
r48 17 18 12.505 $w=2e-07 $l=2.05e-07 $layer=LI1_cond $X=3.435 $Y=1.325
+ $X2=3.435 $Y2=1.53
r49 13 22 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.015 $Y=1.16
+ $X2=3.015 $Y2=1.325
r50 13 21 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.015 $Y=1.16
+ $X2=3.015 $Y2=0.995
r51 13 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=1.16 $X2=2.99 $Y2=1.16
r52 10 17 6.92652 $w=2.5e-07 $l=1.67705e-07 $layer=LI1_cond $X=3.335 $Y=1.2
+ $X2=3.435 $Y2=1.325
r53 10 15 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=3.335 $Y=1.2
+ $X2=2.99 $Y2=1.2
r54 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.075 $Y=1.77
+ $X2=3.075 $Y2=2.055
r55 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.075 $Y=1.67 $X2=3.075
+ $Y2=1.77
r56 6 22 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=3.075 $Y=1.67
+ $X2=3.075 $Y2=1.325
r57 3 21 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.04 $Y=0.445
+ $X2=3.04 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_1%B1 3 6 7 9 10 11 18
r29 16 18 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.645 $Y=1.16
+ $X2=3.875 $Y2=1.16
r30 14 16 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=3.62 $Y=1.16
+ $X2=3.645 $Y2=1.16
r31 10 11 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.88 $Y=1.16 $X2=3.88
+ $Y2=1.53
r32 10 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.875
+ $Y=1.16 $X2=3.875 $Y2=1.16
r33 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.645 $Y=1.77
+ $X2=3.645 $Y2=2.055
r34 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.645 $Y=1.67 $X2=3.645
+ $Y2=1.77
r35 5 16 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.645 $Y=1.325
+ $X2=3.645 $Y2=1.16
r36 5 6 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=3.645 $Y=1.325
+ $X2=3.645 $Y2=1.67
r37 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.62 $Y=0.995
+ $X2=3.62 $Y2=1.16
r38 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.62 $Y=0.995 $X2=3.62
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_1%X 1 2 9 13 14 15 16 19
r21 16 19 11.0812 $w=2.58e-07 $l=2.5e-07 $layer=LI1_cond $X=0.215 $Y=2.21
+ $X2=0.215 $Y2=1.96
r22 14 19 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=0.215 $Y=1.925
+ $X2=0.215 $Y2=1.96
r23 14 15 6.99888 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.215 $Y=1.925
+ $X2=0.215 $Y2=1.795
r24 13 15 61.4753 $w=1.73e-07 $l=9.7e-07 $layer=LI1_cond $X=0.172 $Y=0.825
+ $X2=0.172 $Y2=1.795
r25 7 13 8.46734 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.255 $Y=0.655
+ $X2=0.255 $Y2=0.825
r26 7 9 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=0.255 $Y=0.655
+ $X2=0.255 $Y2=0.38
r27 2 19 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
r28 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_1%VPWR 1 2 3 12 14 16 18 20 25 30 39 42 50
r53 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r54 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r55 42 45 11.5244 $w=3.98e-07 $l=4e-07 $layer=LI1_cond $X=2.065 $Y=2.32
+ $X2=2.065 $Y2=2.72
r56 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r57 37 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r58 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r59 34 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r60 34 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r61 33 36 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r62 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r63 31 45 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.265 $Y=2.72 $X2=2.065
+ $Y2=2.72
r64 31 33 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.265 $Y=2.72
+ $X2=2.53 $Y2=2.72
r65 30 49 5.00668 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=3.705 $Y=2.72
+ $X2=3.922 $Y2=2.72
r66 30 36 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.705 $Y=2.72
+ $X2=3.45 $Y2=2.72
r67 29 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r68 29 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r70 26 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r71 26 28 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r72 25 45 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=1.865 $Y=2.72 $X2=2.065
+ $Y2=2.72
r73 25 28 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.865 $Y=2.72
+ $X2=1.61 $Y2=2.72
r74 20 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r75 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r76 18 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r77 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r78 14 49 2.93018 $w=3.5e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.88 $Y=2.635
+ $X2=3.922 $Y2=2.72
r79 14 16 18.933 $w=3.48e-07 $l=5.75e-07 $layer=LI1_cond $X=3.88 $Y=2.635
+ $X2=3.88 $Y2=2.06
r80 10 39 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r81 10 12 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.32
r82 3 16 600 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=1 $X=3.735
+ $Y=1.845 $X2=3.88 $Y2=2.06
r83 2 42 600 $w=1.7e-07 $l=6.24099e-07 $layer=licon1_PDIFF $count=1 $X=1.72
+ $Y=1.845 $X2=2.065 $Y2=2.32
r84 1 12 600 $w=1.7e-07 $l=9.04599e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.32
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_1%VGND 1 2 11 15 18 19 20 30 31 34 37
r52 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r53 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r54 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r55 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r56 25 28 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r57 25 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r58 24 27 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r59 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r60 22 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.84 $Y=0 $X2=0.755
+ $Y2=0
r61 22 24 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.84 $Y=0 $X2=1.15
+ $Y2=0
r62 20 35 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r63 20 37 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r64 18 27 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.135 $Y=0 $X2=2.99
+ $Y2=0
r65 18 19 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.135 $Y=0 $X2=3.31
+ $Y2=0
r66 17 30 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.485 $Y=0 $X2=3.91
+ $Y2=0
r67 17 19 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.485 $Y=0 $X2=3.31
+ $Y2=0
r68 13 19 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=0.085
+ $X2=3.31 $Y2=0
r69 13 15 10.0427 $w=3.48e-07 $l=3.05e-07 $layer=LI1_cond $X=3.31 $Y=0.085
+ $X2=3.31 $Y2=0.39
r70 9 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0
r71 9 11 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0.525
r72 2 15 182 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.235 $X2=3.315 $Y2=0.39
r73 1 11 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.755 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_1%A_529_47# 1 2 9 11 12 15
r31 13 15 8.56945 $w=3.88e-07 $l=2.9e-07 $layer=LI1_cond $X=3.86 $Y=0.725
+ $X2=3.86 $Y2=0.435
r32 11 13 8.0953 $w=1.8e-07 $l=2.35743e-07 $layer=LI1_cond $X=3.665 $Y=0.815
+ $X2=3.86 $Y2=0.725
r33 11 12 44.3636 $w=1.78e-07 $l=7.2e-07 $layer=LI1_cond $X=3.665 $Y=0.815
+ $X2=2.945 $Y2=0.815
r34 7 12 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=2.82 $Y=0.725
+ $X2=2.945 $Y2=0.815
r35 7 9 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=2.82 $Y=0.725 $X2=2.82
+ $Y2=0.485
r36 2 15 182 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_NDIFF $count=1 $X=3.695
+ $Y=0.235 $X2=3.88 $Y2=0.435
r37 1 9 182 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.485
.ends

