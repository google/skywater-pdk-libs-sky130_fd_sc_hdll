* File: sky130_fd_sc_hdll__dlxtn_4.spice
* Created: Wed Sep  2 08:30:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__dlxtn_4.pex.spice"
.subckt sky130_fd_sc_hdll__dlxtn_4  VNB VPB GATE_N D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* GATE_N	GATE_N
* VPB	VPB
* VNB	VNB
MM1016 N_VGND_M1016_d N_GATE_N_M1016_g N_A_27_47#_M1016_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_A_211_363#_M1001_d N_A_27_47#_M1001_g N_VGND_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0672 PD=1.36 PS=0.74 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_D_M1010_g N_A_319_47#_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1007 A_505_47# N_A_319_47#_M1007_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0933692 AS=0.0672 PD=0.926154 PS=0.74 NRD=47.796 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1008 N_A_609_413#_M1008_d N_A_27_47#_M1008_g A_505_47# VNB NSHORT L=0.15
+ W=0.36 AD=0.0504 AS=0.0800308 PD=0.64 PS=0.793846 NRD=0 NRS=55.764 M=1 R=2.4
+ SA=75001.3 SB=75001.1 A=0.054 P=1.02 MULT=1
MM1000 A_709_47# N_A_211_363#_M1000_g N_A_609_413#_M1008_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0609231 AS=0.0504 PD=0.687692 PS=0.64 NRD=38.076 NRS=0 M=1 R=2.4
+ SA=75001.7 SB=75000.7 A=0.054 P=1.02 MULT=1
MM1009 N_VGND_M1009_d N_A_774_21#_M1009_g A_709_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0710769 PD=1.46 PS=0.802308 NRD=12.852 NRS=32.628 M=1 R=2.8
+ SA=75001.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_609_413#_M1014_g N_A_774_21#_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.108875 AS=0.2015 PD=0.985 PS=1.92 NRD=1.836 NRS=2.76 M=1 R=4.33333
+ SA=75000.2 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1003 N_Q_M1003_d N_A_774_21#_M1003_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.108875 PD=0.97 PS=0.985 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1005 N_Q_M1003_d N_A_774_21#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1012 N_Q_M1012_d N_A_774_21#_M1012_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.7
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1021 N_Q_M1012_d N_A_774_21#_M1021_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.169 PD=0.97 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_GATE_N_M1004_g N_A_27_47#_M1004_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1019 N_A_211_363#_M1019_d N_A_27_47#_M1019_g N_VPWR_M1004_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1011 N_VPWR_M1011_d N_D_M1011_g N_A_319_47#_M1011_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90001.7 A=0.1152 P=1.64 MULT=1
MM1006 A_503_369# N_A_319_47#_M1006_g N_VPWR_M1011_d VPB PHIGHVT L=0.18 W=0.64
+ AD=0.123291 AS=0.0928 PD=1.19547 PS=0.93 NRD=42.355 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90001.2 A=0.1152 P=1.64 MULT=1
MM1018 N_A_609_413#_M1018_d N_A_211_363#_M1018_g A_503_369# VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0609 AS=0.0809094 PD=0.71 PS=0.784528 NRD=2.3443 NRS=64.5569 M=1
+ R=2.33333 SA=90001.2 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1015 A_703_413# N_A_27_47#_M1015_g N_A_609_413#_M1018_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.07665 AS=0.0609 PD=0.785 PS=0.71 NRD=59.7895 NRS=2.3443 M=1
+ R=2.33333 SA=90001.6 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1022 N_VPWR_M1022_d N_A_774_21#_M1022_g A_703_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.1134 AS=0.07665 PD=1.38 PS=0.785 NRD=2.3443 NRS=59.7895 M=1 R=2.33333
+ SA=90002.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1017 N_VPWR_M1017_d N_A_609_413#_M1017_g N_A_774_21#_M1017_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.1525 AS=0.27 PD=1.305 PS=2.54 NRD=3.9203 NRS=0.9653 M=1
+ R=5.55556 SA=90000.2 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1002 N_Q_M1002_d N_A_774_21#_M1002_g N_VPWR_M1017_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.1525 PD=1.29 PS=1.305 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1013 N_Q_M1002_d N_A_774_21#_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1020 N_Q_M1020_d N_A_774_21#_M1020_g N_VPWR_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1023 N_Q_M1020_d N_A_774_21#_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90000.2 A=0.18 P=2.36 MULT=1
DX24_noxref VNB VPB NWDIODE A=12.4227 P=18.69
c_136 VPB 0 1.69345e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__dlxtn_4.pxi.spice"
*
.ends
*
*
