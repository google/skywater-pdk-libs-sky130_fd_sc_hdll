* File: sky130_fd_sc_hdll__a21o_6.pex.spice
* Created: Thu Aug 27 18:53:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A21O_6%A2 1 3 4 6 7 9 10 12 14 15 16 18 19 23 26
c88 18 0 1.53044e-19 $X=1.79 $Y=1.46
c89 14 0 1.34369e-19 $X=0.61 $Y=1.46
c90 10 0 1.86168e-19 $X=1.905 $Y=1.41
r91 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.49
+ $Y=1.16 $X2=0.49 $Y2=1.16
r92 26 30 12.7504 $w=2.33e-07 $l=2.6e-07 $layer=LI1_cond $X=0.23 $Y=1.172
+ $X2=0.49 $Y2=1.172
r93 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.16 $X2=1.88 $Y2=1.16
r94 20 23 4.41361 $w=2.33e-07 $l=9e-08 $layer=LI1_cond $X=1.79 $Y=1.172 $X2=1.88
+ $Y2=1.172
r95 19 30 1.7164 $w=2.33e-07 $l=3.5e-08 $layer=LI1_cond $X=0.525 $Y=1.172
+ $X2=0.49 $Y2=1.172
r96 17 20 2.6346 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=1.79 $Y=1.29 $X2=1.79
+ $Y2=1.172
r97 17 18 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.79 $Y=1.29
+ $X2=1.79 $Y2=1.46
r98 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.705 $Y=1.545
+ $X2=1.79 $Y2=1.46
r99 15 16 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=1.705 $Y=1.545
+ $X2=0.695 $Y2=1.545
r100 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.46
+ $X2=0.695 $Y2=1.545
r101 13 19 7.04737 $w=2.35e-07 $l=1.54771e-07 $layer=LI1_cond $X=0.61 $Y=1.29
+ $X2=0.525 $Y2=1.172
r102 13 14 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.61 $Y=1.29
+ $X2=0.61 $Y2=1.46
r103 10 24 51.486 $w=2.55e-07 $l=2.62202e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.88 $Y2=1.16
r104 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r105 7 24 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.82 $Y=0.995
+ $X2=1.88 $Y2=1.16
r106 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.82 $Y=0.995
+ $X2=1.82 $Y2=0.56
r107 4 29 38.5416 $w=3.03e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.58 $Y=0.995
+ $X2=0.49 $Y2=1.16
r108 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.58 $Y=0.995
+ $X2=0.58 $Y2=0.56
r109 1 29 47.6478 $w=3.03e-07 $l=2.52488e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.49 $Y2=1.16
r110 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_6%A1 1 3 4 6 7 9 10 12 13 19 20
r52 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.202
+ $X2=1.435 $Y2=1.202
r53 18 20 5.07368 $w=3.8e-07 $l=4e-08 $layer=POLY_cond $X=1.37 $Y=1.202 $X2=1.41
+ $Y2=1.202
r54 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.37
+ $Y=1.16 $X2=1.37 $Y2=1.16
r55 16 18 48.2 $w=3.8e-07 $l=3.8e-07 $layer=POLY_cond $X=0.99 $Y=1.202 $X2=1.37
+ $Y2=1.202
r56 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r57 13 19 10.7888 $w=2.33e-07 $l=2.2e-07 $layer=LI1_cond $X=1.15 $Y=1.172
+ $X2=1.37 $Y2=1.172
r58 10 21 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r59 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r60 7 20 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.202
r61 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995 $X2=1.41
+ $Y2=0.56
r62 4 16 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r63 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995 $X2=0.99
+ $Y2=0.56
r64 1 15 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r65 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_6%B1 1 3 4 6 7 9 10 12 13 18
c54 1 0 1.53044e-19 $X=2.375 $Y=1.41
r55 18 20 24.3634 $w=3.66e-07 $l=1.85e-07 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=3.03 $Y2=1.202
r56 17 18 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.845 $Y2=1.202
r57 16 17 55.3115 $w=3.66e-07 $l=4.2e-07 $layer=POLY_cond $X=2.4 $Y=1.202
+ $X2=2.82 $Y2=1.202
r58 15 16 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.4 $Y2=1.202
r59 13 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.03
+ $Y=1.16 $X2=3.03 $Y2=1.16
r60 10 18 19.3576 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r61 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r62 7 17 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=1.202
r63 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.82 $Y=0.995 $X2=2.82
+ $Y2=0.56
r64 4 16 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.4 $Y=0.995 $X2=2.4
+ $Y2=1.202
r65 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.4 $Y=0.995 $X2=2.4
+ $Y2=0.56
r66 1 15 19.3576 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r67 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_6%A_213_47# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 39 40 42 43 45 48 50 51 54 59 60 63 64 69 72 74
+ 89
r180 89 90 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=6.16 $Y=1.202
+ $X2=6.185 $Y2=1.202
r181 88 89 54.8618 $w=3.69e-07 $l=4.2e-07 $layer=POLY_cond $X=5.74 $Y=1.202
+ $X2=6.16 $Y2=1.202
r182 87 88 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=5.715 $Y=1.202
+ $X2=5.74 $Y2=1.202
r183 84 85 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=5.22 $Y=1.202
+ $X2=5.245 $Y2=1.202
r184 83 84 54.8618 $w=3.69e-07 $l=4.2e-07 $layer=POLY_cond $X=4.8 $Y=1.202
+ $X2=5.22 $Y2=1.202
r185 82 83 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=4.775 $Y=1.202
+ $X2=4.8 $Y2=1.202
r186 81 82 61.393 $w=3.69e-07 $l=4.7e-07 $layer=POLY_cond $X=4.305 $Y=1.202
+ $X2=4.775 $Y2=1.202
r187 80 81 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=4.28 $Y=1.202
+ $X2=4.305 $Y2=1.202
r188 77 78 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=3.835 $Y=1.202
+ $X2=3.86 $Y2=1.202
r189 74 75 6.88461 $w=2.98e-07 $l=1.7e-07 $layer=LI1_cond $X=2.595 $Y=1.96
+ $X2=2.595 $Y2=1.79
r190 70 87 55.5149 $w=3.69e-07 $l=4.25e-07 $layer=POLY_cond $X=5.29 $Y=1.202
+ $X2=5.715 $Y2=1.202
r191 70 85 5.87805 $w=3.69e-07 $l=4.5e-08 $layer=POLY_cond $X=5.29 $Y=1.202
+ $X2=5.245 $Y2=1.202
r192 69 70 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.29
+ $Y=1.16 $X2=5.29 $Y2=1.16
r193 67 80 45.7182 $w=3.69e-07 $l=3.5e-07 $layer=POLY_cond $X=3.93 $Y=1.202
+ $X2=4.28 $Y2=1.202
r194 67 78 9.14363 $w=3.69e-07 $l=7e-08 $layer=POLY_cond $X=3.93 $Y=1.202
+ $X2=3.86 $Y2=1.202
r195 66 69 65.3051 $w=2.38e-07 $l=1.36e-06 $layer=LI1_cond $X=3.93 $Y=1.155
+ $X2=5.29 $Y2=1.155
r196 66 67 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.93
+ $Y=1.16 $X2=3.93 $Y2=1.16
r197 64 66 9.3636 $w=2.38e-07 $l=1.95e-07 $layer=LI1_cond $X=3.735 $Y=1.155
+ $X2=3.93 $Y2=1.155
r198 63 64 7.07814 $w=2.4e-07 $l=1.56844e-07 $layer=LI1_cond $X=3.65 $Y=1.035
+ $X2=3.735 $Y2=1.155
r199 62 63 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.65 $Y=0.885
+ $X2=3.65 $Y2=1.035
r200 61 72 3.9099 $w=2.1e-07 $l=1.5e-07 $layer=LI1_cond $X=2.745 $Y=0.78
+ $X2=2.595 $Y2=0.78
r201 60 62 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.565 $Y=0.78
+ $X2=3.65 $Y2=0.885
r202 60 61 43.3074 $w=2.08e-07 $l=8.2e-07 $layer=LI1_cond $X=3.565 $Y=0.78
+ $X2=2.745 $Y2=0.78
r203 59 75 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=2.57 $Y=1.62
+ $X2=2.57 $Y2=1.79
r204 56 72 2.27033 $w=2.5e-07 $l=1.16833e-07 $layer=LI1_cond $X=2.57 $Y=0.885
+ $X2=2.595 $Y2=0.78
r205 56 59 33.8818 $w=2.48e-07 $l=7.35e-07 $layer=LI1_cond $X=2.57 $Y=0.885
+ $X2=2.57 $Y2=1.62
r206 52 72 2.27033 $w=3e-07 $l=1.05e-07 $layer=LI1_cond $X=2.595 $Y=0.675
+ $X2=2.595 $Y2=0.78
r207 52 54 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=2.595 $Y=0.675
+ $X2=2.595 $Y2=0.42
r208 50 72 3.9099 $w=2.1e-07 $l=1.5e-07 $layer=LI1_cond $X=2.445 $Y=0.78
+ $X2=2.595 $Y2=0.78
r209 50 51 57.039 $w=2.08e-07 $l=1.08e-06 $layer=LI1_cond $X=2.445 $Y=0.78
+ $X2=1.365 $Y2=0.78
r210 46 51 7.26367 $w=2.1e-07 $l=2.11069e-07 $layer=LI1_cond $X=1.2 $Y=0.675
+ $X2=1.365 $Y2=0.78
r211 46 48 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=0.675
+ $X2=1.2 $Y2=0.38
r212 43 90 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.202
r213 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.985
r214 40 89 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=1.202
r215 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=0.56
r216 37 88 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.74 $Y=0.995
+ $X2=5.74 $Y2=1.202
r217 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.74 $Y=0.995
+ $X2=5.74 $Y2=0.56
r218 34 87 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.202
r219 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.985
r220 31 85 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.202
r221 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.985
r222 28 84 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.22 $Y=0.995
+ $X2=5.22 $Y2=1.202
r223 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.22 $Y=0.995
+ $X2=5.22 $Y2=0.56
r224 25 83 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.8 $Y=0.995
+ $X2=4.8 $Y2=1.202
r225 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.8 $Y=0.995
+ $X2=4.8 $Y2=0.56
r226 22 82 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.202
r227 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
r228 19 81 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.202
r229 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.985
r230 16 80 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.28 $Y=0.995
+ $X2=4.28 $Y2=1.202
r231 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.28 $Y=0.995
+ $X2=4.28 $Y2=0.56
r232 13 78 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.86 $Y=0.995
+ $X2=3.86 $Y2=1.202
r233 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.86 $Y=0.995
+ $X2=3.86 $Y2=0.56
r234 10 77 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.202
r235 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.985
r236 3 74 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.96
r237 3 59 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.62
r238 2 54 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=2.475
+ $Y=0.235 $X2=2.61 $Y2=0.42
r239 1 48 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_6%A_27_297# 1 2 3 4 15 19 21 25 28 33 35 36
+ 39 41 43 44
c71 33 0 1.86168e-19 $X=2.14 $Y=1.63
r72 37 39 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=3.08 $Y=2.295
+ $X2=3.08 $Y2=1.87
r73 35 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.915 $Y=2.38
+ $X2=3.08 $Y2=2.295
r74 35 36 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.915 $Y=2.38
+ $X2=2.275 $Y2=2.38
r75 31 44 3.52026 $w=2.65e-07 $l=1.00995e-07 $layer=LI1_cond $X=2.16 $Y=1.8
+ $X2=2.125 $Y2=1.885
r76 31 33 8.51806 $w=2.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.16 $Y=1.8 $X2=2.16
+ $Y2=1.63
r77 30 44 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=1.97
+ $X2=2.125 $Y2=1.885
r78 28 36 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.125 $Y=2.295
+ $X2=2.275 $Y2=2.38
r79 28 30 12.4848 $w=2.98e-07 $l=3.25e-07 $layer=LI1_cond $X=2.125 $Y=2.295
+ $X2=2.125 $Y2=1.97
r80 26 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=1.885
+ $X2=1.2 $Y2=1.885
r81 25 44 2.98021 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.975 $Y=1.885
+ $X2=2.125 $Y2=1.885
r82 25 26 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.975 $Y=1.885
+ $X2=1.365 $Y2=1.885
r83 22 41 3.3845 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=1.885
+ $X2=0.26 $Y2=1.885
r84 21 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=1.885
+ $X2=1.2 $Y2=1.885
r85 21 22 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.035 $Y=1.885
+ $X2=0.425 $Y2=1.885
r86 17 41 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.97
+ $X2=0.26 $Y2=1.885
r87 17 19 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=0.26 $Y=1.97 $X2=0.26
+ $Y2=2
r88 13 41 3.19717 $w=2.95e-07 $l=1.00995e-07 $layer=LI1_cond $X=0.225 $Y=1.8
+ $X2=0.26 $Y2=1.885
r89 13 15 6.20546 $w=2.58e-07 $l=1.4e-07 $layer=LI1_cond $X=0.225 $Y=1.8
+ $X2=0.225 $Y2=1.66
r90 4 39 300 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=1.87
r91 3 33 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.63
r92 3 30 300 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.97
r93 2 43 300 $w=1.7e-07 $l=4.66905e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.885
r94 1 19 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
r95 1 15 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_6%VPWR 1 2 3 4 5 6 21 23 27 31 37 41 45 50 51
+ 53 54 56 57 59 60 61 63 85 86 89 92
r108 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r109 90 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r110 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r111 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r112 83 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r113 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r114 80 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r115 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r116 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r117 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r118 74 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r119 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r120 71 74 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r121 71 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r122 70 73 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r123 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r124 68 92 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=1.67 $Y2=2.72
r125 68 70 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=2.07 $Y2=2.72
r126 63 89 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.73 $Y2=2.72
r127 63 65 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r128 61 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r129 61 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r130 59 82 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=6.265 $Y=2.72
+ $X2=6.21 $Y2=2.72
r131 59 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.265 $Y=2.72
+ $X2=6.43 $Y2=2.72
r132 58 85 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.595 $Y=2.72
+ $X2=6.67 $Y2=2.72
r133 58 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.595 $Y=2.72
+ $X2=6.43 $Y2=2.72
r134 56 79 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.315 $Y=2.72
+ $X2=5.29 $Y2=2.72
r135 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.315 $Y=2.72
+ $X2=5.48 $Y2=2.72
r136 55 82 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.645 $Y=2.72
+ $X2=6.21 $Y2=2.72
r137 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.645 $Y=2.72
+ $X2=5.48 $Y2=2.72
r138 53 76 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.375 $Y=2.72
+ $X2=4.37 $Y2=2.72
r139 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.375 $Y=2.72
+ $X2=4.54 $Y2=2.72
r140 52 79 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.705 $Y=2.72
+ $X2=5.29 $Y2=2.72
r141 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=2.72
+ $X2=4.54 $Y2=2.72
r142 50 73 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.485 $Y=2.72
+ $X2=3.45 $Y2=2.72
r143 50 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.485 $Y=2.72
+ $X2=3.61 $Y2=2.72
r144 49 76 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.735 $Y=2.72
+ $X2=4.37 $Y2=2.72
r145 49 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.735 $Y=2.72
+ $X2=3.61 $Y2=2.72
r146 45 48 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.43 $Y=1.63
+ $X2=6.43 $Y2=2.31
r147 43 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.43 $Y=2.635
+ $X2=6.43 $Y2=2.72
r148 43 48 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6.43 $Y=2.635
+ $X2=6.43 $Y2=2.31
r149 39 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2.72
r150 39 41 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=1.87
r151 35 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=2.635
+ $X2=4.54 $Y2=2.72
r152 35 37 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=4.54 $Y=2.635
+ $X2=4.54 $Y2=1.87
r153 31 34 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=3.61 $Y=1.66
+ $X2=3.61 $Y2=2.34
r154 29 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.61 $Y=2.635
+ $X2=3.61 $Y2=2.72
r155 29 34 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.61 $Y=2.635
+ $X2=3.61 $Y2=2.34
r156 25 92 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.72
r157 25 27 14.0854 $w=2.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.305
r158 24 89 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.865 $Y=2.72
+ $X2=0.73 $Y2=2.72
r159 23 92 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.535 $Y=2.72
+ $X2=1.67 $Y2=2.72
r160 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.535 $Y=2.72
+ $X2=0.865 $Y2=2.72
r161 19 89 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.72
r162 19 21 14.0854 $w=2.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.305
r163 6 48 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=6.275
+ $Y=1.485 $X2=6.42 $Y2=2.31
r164 6 45 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.275
+ $Y=1.485 $X2=6.42 $Y2=1.63
r165 5 41 300 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_PDIFF $count=2 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=1.87
r166 4 37 300 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_PDIFF $count=2 $X=4.395
+ $Y=1.485 $X2=4.54 $Y2=1.87
r167 3 34 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=3.475
+ $Y=1.485 $X2=3.6 $Y2=2.34
r168 3 31 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=3.475
+ $Y=1.485 $X2=3.6 $Y2=1.66
r169 2 27 600 $w=1.7e-07 $l=8.8955e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.305
r170 1 21 600 $w=1.7e-07 $l=8.8955e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.305
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_6%X 1 2 3 4 5 6 21 25 29 30 31 32 35 39 43 45
+ 49 51 53 57 58 60 65
r93 62 65 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=5.75 $Y=1.445
+ $X2=5.75 $Y2=1.19
r94 59 65 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=5.75 $Y=0.865
+ $X2=5.75 $Y2=1.19
r95 59 60 3.24686 $w=2.9e-07 $l=1.56844e-07 $layer=LI1_cond $X=5.75 $Y=0.865
+ $X2=5.87 $Y2=0.78
r96 53 55 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.95 $Y=1.62
+ $X2=5.95 $Y2=2.3
r97 51 62 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=5.95 $Y=1.53 $X2=5.75
+ $Y2=1.53
r98 51 53 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=5.95 $Y=1.615
+ $X2=5.95 $Y2=1.62
r99 47 60 3.24686 $w=2.9e-07 $l=1.18427e-07 $layer=LI1_cond $X=5.95 $Y=0.695
+ $X2=5.87 $Y2=0.78
r100 47 49 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.95 $Y=0.695
+ $X2=5.95 $Y2=0.36
r101 46 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.175 $Y=0.78
+ $X2=5.01 $Y2=0.78
r102 45 60 3.3199 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=5.625 $Y=0.78
+ $X2=5.87 $Y2=0.78
r103 45 46 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.625 $Y=0.78
+ $X2=5.175 $Y2=0.78
r104 44 58 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.145 $Y=1.53
+ $X2=5.01 $Y2=1.53
r105 43 62 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.625 $Y=1.53
+ $X2=5.75 $Y2=1.53
r106 43 44 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=5.625 $Y=1.53
+ $X2=5.145 $Y2=1.53
r107 39 41 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.01 $Y=1.62
+ $X2=5.01 $Y2=2.3
r108 37 58 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.01 $Y=1.615
+ $X2=5.01 $Y2=1.53
r109 37 39 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=5.01 $Y=1.615
+ $X2=5.01 $Y2=1.62
r110 33 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.01 $Y=0.695
+ $X2=5.01 $Y2=0.78
r111 33 35 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.01 $Y=0.695
+ $X2=5.01 $Y2=0.36
r112 31 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.845 $Y=0.78
+ $X2=5.01 $Y2=0.78
r113 31 32 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.845 $Y=0.78
+ $X2=4.235 $Y2=0.78
r114 29 58 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.875 $Y=1.53
+ $X2=5.01 $Y2=1.53
r115 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.875 $Y=1.53
+ $X2=4.205 $Y2=1.53
r116 25 27 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.07 $Y=1.62
+ $X2=4.07 $Y2=2.3
r117 23 30 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.07 $Y=1.615
+ $X2=4.205 $Y2=1.53
r118 23 25 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=4.07 $Y=1.615
+ $X2=4.07 $Y2=1.62
r119 19 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.07 $Y=0.695
+ $X2=4.235 $Y2=0.78
r120 19 21 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.07 $Y=0.695
+ $X2=4.07 $Y2=0.36
r121 6 55 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=2.3
r122 6 53 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=1.62
r123 5 41 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=2.3
r124 5 39 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=1.62
r125 4 27 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=2.3
r126 4 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=1.62
r127 3 49 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=5.815
+ $Y=0.235 $X2=5.95 $Y2=0.36
r128 2 35 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=4.875
+ $Y=0.235 $X2=5.01 $Y2=0.36
r129 1 21 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=3.935
+ $Y=0.235 $X2=4.07 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_6%VGND 1 2 3 4 5 6 19 21 25 31 35 39 42 43 45
+ 46 48 49 50 52 71 72 78 83 89
r97 88 89 10.0909 $w=5.88e-07 $l=1.65e-07 $layer=LI1_cond $X=3.57 $Y=0.21
+ $X2=3.735 $Y2=0.21
r98 85 88 2.4327 $w=5.88e-07 $l=1.2e-07 $layer=LI1_cond $X=3.45 $Y=0.21 $X2=3.57
+ $Y2=0.21
r99 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r100 82 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r101 81 85 9.32536 $w=5.88e-07 $l=4.6e-07 $layer=LI1_cond $X=2.99 $Y=0.21
+ $X2=3.45 $Y2=0.21
r102 81 83 8.2664 $w=5.88e-07 $l=7.5e-08 $layer=LI1_cond $X=2.99 $Y=0.21
+ $X2=2.915 $Y2=0.21
r103 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r104 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r105 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r106 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r107 69 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r108 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r109 66 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r110 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r111 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r112 63 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.45
+ $Y2=0
r113 62 89 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.37 $Y=0
+ $X2=3.735 $Y2=0
r114 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r115 59 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r116 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r117 56 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r118 55 58 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r119 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r120 53 75 4.56433 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=0.535 $Y=0
+ $X2=0.267 $Y2=0
r121 53 55 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.535 $Y=0
+ $X2=0.69 $Y2=0
r122 52 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=2.11
+ $Y2=0
r123 52 58 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.945 $Y=0
+ $X2=1.61 $Y2=0
r124 50 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r125 50 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r126 48 68 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.285 $Y=0 $X2=6.21
+ $Y2=0
r127 48 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.285 $Y=0 $X2=6.41
+ $Y2=0
r128 47 71 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.535 $Y=0
+ $X2=6.67 $Y2=0
r129 47 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.535 $Y=0 $X2=6.41
+ $Y2=0
r130 45 65 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=5.345 $Y=0 $X2=5.29
+ $Y2=0
r131 45 46 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.345 $Y=0 $X2=5.48
+ $Y2=0
r132 44 68 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.615 $Y=0
+ $X2=6.21 $Y2=0
r133 44 46 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.615 $Y=0 $X2=5.48
+ $Y2=0
r134 42 62 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.405 $Y=0 $X2=4.37
+ $Y2=0
r135 42 43 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.405 $Y=0 $X2=4.54
+ $Y2=0
r136 41 65 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.675 $Y=0 $X2=5.29
+ $Y2=0
r137 41 43 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.675 $Y=0 $X2=4.54
+ $Y2=0
r138 37 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.41 $Y=0.085
+ $X2=6.41 $Y2=0
r139 37 39 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=6.41 $Y=0.085
+ $X2=6.41 $Y2=0.36
r140 33 46 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0
r141 33 35 11.7378 $w=2.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.36
r142 29 43 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0
r143 29 31 11.7378 $w=2.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0.36
r144 28 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.11
+ $Y2=0
r145 28 83 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.915
+ $Y2=0
r146 23 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.11 $Y2=0
r147 23 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.11 $Y2=0.38
r148 19 75 3.20184 $w=3.3e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.37 $Y=0.085
+ $X2=0.267 $Y2=0
r149 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.37 $Y=0.085
+ $X2=0.37 $Y2=0.38
r150 6 39 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=6.235
+ $Y=0.235 $X2=6.37 $Y2=0.36
r151 5 35 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=5.295
+ $Y=0.235 $X2=5.48 $Y2=0.36
r152 4 31 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=4.355
+ $Y=0.235 $X2=4.54 $Y2=0.36
r153 3 88 91 $w=1.7e-07 $l=7.43976e-07 $layer=licon1_NDIFF $count=2 $X=2.895
+ $Y=0.235 $X2=3.57 $Y2=0.38
r154 2 25 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.235 $X2=2.11 $Y2=0.38
r155 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.245
+ $Y=0.235 $X2=0.37 $Y2=0.38
.ends

