* File: sky130_fd_sc_hdll__and4_4.pxi.spice
* Created: Thu Aug 27 18:58:53 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND4_4%A N_A_c_71_n N_A_M1006_g N_A_c_68_n N_A_M1012_g A
+ A N_A_c_70_n PM_SKY130_FD_SC_HDLL__AND4_4%A
x_PM_SKY130_FD_SC_HDLL__AND4_4%B N_B_c_97_n N_B_M1001_g N_B_c_98_n N_B_M1002_g B
+ B B PM_SKY130_FD_SC_HDLL__AND4_4%B
x_PM_SKY130_FD_SC_HDLL__AND4_4%C N_C_c_128_n N_C_M1015_g N_C_c_129_n N_C_M1003_g
+ C C C PM_SKY130_FD_SC_HDLL__AND4_4%C
x_PM_SKY130_FD_SC_HDLL__AND4_4%D N_D_c_159_n N_D_M1005_g N_D_c_160_n N_D_M1000_g
+ D PM_SKY130_FD_SC_HDLL__AND4_4%D
x_PM_SKY130_FD_SC_HDLL__AND4_4%A_27_47# N_A_27_47#_M1012_s N_A_27_47#_M1006_d
+ N_A_27_47#_M1003_d N_A_27_47#_c_196_n N_A_27_47#_M1004_g N_A_27_47#_c_203_n
+ N_A_27_47#_M1007_g N_A_27_47#_c_197_n N_A_27_47#_M1008_g N_A_27_47#_c_204_n
+ N_A_27_47#_M1010_g N_A_27_47#_c_198_n N_A_27_47#_M1009_g N_A_27_47#_c_205_n
+ N_A_27_47#_M1011_g N_A_27_47#_c_206_n N_A_27_47#_M1014_g N_A_27_47#_c_199_n
+ N_A_27_47#_M1013_g N_A_27_47#_c_200_n N_A_27_47#_c_223_n N_A_27_47#_c_224_n
+ N_A_27_47#_c_236_n N_A_27_47#_c_237_n N_A_27_47#_c_208_n N_A_27_47#_c_201_n
+ N_A_27_47#_c_278_p N_A_27_47#_c_215_n N_A_27_47#_c_218_n N_A_27_47#_c_230_n
+ N_A_27_47#_c_202_n PM_SKY130_FD_SC_HDLL__AND4_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__AND4_4%VPWR N_VPWR_M1006_s N_VPWR_M1002_d N_VPWR_M1000_d
+ N_VPWR_M1010_d N_VPWR_M1014_d N_VPWR_c_331_n N_VPWR_c_332_n N_VPWR_c_333_n
+ N_VPWR_c_334_n N_VPWR_c_335_n N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n
+ N_VPWR_c_339_n N_VPWR_c_340_n N_VPWR_c_341_n VPWR N_VPWR_c_342_n
+ N_VPWR_c_343_n N_VPWR_c_344_n N_VPWR_c_330_n PM_SKY130_FD_SC_HDLL__AND4_4%VPWR
x_PM_SKY130_FD_SC_HDLL__AND4_4%X N_X_M1004_s N_X_M1009_s N_X_M1007_s N_X_M1011_s
+ N_X_c_410_n N_X_c_411_n N_X_c_415_n N_X_c_409_n N_X_c_422_n N_X_c_405_n
+ N_X_c_432_n N_X_c_434_n N_X_c_436_n N_X_c_439_n N_X_c_440_n N_X_c_406_n X X X
+ N_X_c_403_n N_X_c_407_n X PM_SKY130_FD_SC_HDLL__AND4_4%X
x_PM_SKY130_FD_SC_HDLL__AND4_4%VGND N_VGND_M1005_d N_VGND_M1008_d N_VGND_M1013_d
+ N_VGND_c_493_n N_VGND_c_494_n N_VGND_c_495_n N_VGND_c_496_n N_VGND_c_497_n
+ N_VGND_c_498_n N_VGND_c_499_n N_VGND_c_500_n VGND N_VGND_c_501_n
+ N_VGND_c_502_n PM_SKY130_FD_SC_HDLL__AND4_4%VGND
cc_1 VNB N_A_c_68_n 0.0185442f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB A 0.00892312f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_A_c_70_n 0.0461216f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_B_c_97_n 0.0165235f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_B_c_98_n 0.0241017f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB B 0.0024573f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_7 VNB N_C_c_128_n 0.0184065f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_8 VNB N_C_c_129_n 0.0318223f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_9 VNB C 7.25139e-19 $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_10 VNB N_D_c_159_n 0.0162318f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_11 VNB N_D_c_160_n 0.0259683f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_12 VNB D 0.00372234f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_13 VNB N_A_27_47#_c_196_n 0.0174554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_197_n 0.0167427f $X=-0.19 $Y=-0.24 $X2=0.227 $Y2=0.85
cc_15 VNB N_A_27_47#_c_198_n 0.0171812f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_199_n 0.0189221f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_200_n 0.00248426f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_201_n 0.00273989f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_202_n 0.076126f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_330_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_X_c_403_n 0.00770055f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB X 0.0247728f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_493_n 0.00489575f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_24 VNB N_VGND_c_494_n 3.24573e-19 $X=-0.19 $Y=-0.24 $X2=0.227 $Y2=0.85
cc_25 VNB N_VGND_c_495_n 0.0128379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_496_n 0.0122245f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_497_n 0.0619174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_498_n 0.00593471f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_499_n 0.0153278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_500_n 0.00502664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_501_n 0.0123502f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_502_n 0.24128f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VPB N_A_c_71_n 0.0188726f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_34 VPB A 0.0126686f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_35 VPB N_A_c_70_n 0.0164787f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_36 VPB N_B_c_98_n 0.0270758f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_37 VPB B 0.00273724f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_38 VPB N_C_c_129_n 0.0317805f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_39 VPB C 0.00191243f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_40 VPB N_D_c_160_n 0.0287616f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_41 VPB D 9.54851e-19 $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_42 VPB N_A_27_47#_c_203_n 0.0162781f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_43 VPB N_A_27_47#_c_204_n 0.0162026f $X=-0.19 $Y=1.305 $X2=0.227 $Y2=1.16
cc_44 VPB N_A_27_47#_c_205_n 0.0160348f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_47#_c_206_n 0.0179643f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_27_47#_c_200_n 0.00168395f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_27_47#_c_208_n 0.00173767f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_27_47#_c_202_n 0.0470977f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_331_n 0.0109102f $X=-0.19 $Y=1.305 $X2=0.227 $Y2=0.85
cc_50 VPB N_VPWR_c_332_n 0.0294551f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_333_n 0.00508424f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_334_n 0.00291475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_335_n 0.00234357f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_336_n 0.0129491f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_337_n 0.0254666f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_338_n 0.0248982f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_339_n 0.00519718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_340_n 0.018706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_341_n 0.00359922f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_342_n 0.0193003f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_343_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_344_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_330_n 0.0462084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_X_c_405_n 0.00105739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_X_c_406_n 0.00105739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_X_c_407_n 0.0118427f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB X 0.00909869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 N_A_c_68_n N_B_c_97_n 0.0299922f $X=0.52 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_69 N_A_c_71_n N_B_c_98_n 0.0203669f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_70 N_A_c_70_n N_B_c_98_n 0.0345682f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_71 N_A_c_68_n B 8.43474e-19 $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_72 A N_A_27_47#_M1012_s 0.00411512f $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_73 N_A_c_71_n N_A_27_47#_c_200_n 0.00189679f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_74 N_A_c_68_n N_A_27_47#_c_200_n 0.0150149f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_75 A N_A_27_47#_c_200_n 0.0524527f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_76 N_A_c_70_n N_A_27_47#_c_200_n 0.0116298f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_77 N_A_c_68_n N_A_27_47#_c_215_n 0.0107557f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_78 A N_A_27_47#_c_215_n 0.0120742f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_79 N_A_c_70_n N_A_27_47#_c_215_n 0.00355245f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_80 N_A_c_71_n N_A_27_47#_c_218_n 0.00943614f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_81 A N_A_27_47#_c_218_n 0.0127418f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_82 A N_VPWR_M1006_s 0.00511992f $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_83 N_A_c_71_n N_VPWR_c_332_n 0.0034823f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_84 A N_VPWR_c_332_n 0.0175645f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_85 N_A_c_70_n N_VPWR_c_332_n 0.00240218f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_86 N_A_c_71_n N_VPWR_c_342_n 0.00702461f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_c_71_n N_VPWR_c_330_n 0.0133458f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A_c_68_n N_VGND_c_497_n 0.00357877f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_89 N_A_c_68_n N_VGND_c_502_n 0.00618659f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_90 A N_VGND_c_502_n 0.00238628f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_91 N_B_c_97_n N_C_c_128_n 0.0259777f $X=0.915 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_92 B N_C_c_128_n 0.00641522f $X=1.065 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_93 N_B_c_98_n N_C_c_129_n 0.0454118f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_94 N_B_c_97_n C 3.71388e-19 $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_95 N_B_c_98_n C 2.37481e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_96 B C 0.0517906f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_97 N_B_c_97_n N_A_27_47#_c_200_n 0.00439784f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_98 N_B_c_98_n N_A_27_47#_c_200_n 0.00392522f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_99 B N_A_27_47#_c_200_n 0.0576674f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_100 N_B_c_98_n N_A_27_47#_c_223_n 0.00805815f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_101 N_B_c_98_n N_A_27_47#_c_224_n 0.0185904f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_102 B N_A_27_47#_c_224_n 0.0333788f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_103 N_B_c_97_n N_A_27_47#_c_215_n 0.00552502f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_104 B N_A_27_47#_c_215_n 0.0136168f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_105 N_B_c_98_n N_VPWR_c_333_n 0.00186534f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_106 N_B_c_98_n N_VPWR_c_342_n 0.00700684f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_107 N_B_c_98_n N_VPWR_c_330_n 0.0124944f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_108 B A_198_47# 0.00670646f $X=1.065 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_109 N_B_c_97_n N_VGND_c_497_n 0.00456292f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_110 B N_VGND_c_497_n 0.0137432f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_111 N_B_c_97_n N_VGND_c_502_n 0.00750031f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_112 B N_VGND_c_502_n 0.0153723f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_113 N_C_c_128_n N_D_c_159_n 0.0201458f $X=1.445 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_114 C N_D_c_159_n 0.00639764f $X=1.525 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_115 N_C_c_129_n N_D_c_160_n 0.0421471f $X=1.475 $Y=1.41 $X2=0 $Y2=0
cc_116 C N_D_c_160_n 4.00479e-19 $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_117 N_C_c_128_n D 3.53395e-19 $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_118 N_C_c_129_n D 0.00197007f $X=1.475 $Y=1.41 $X2=0 $Y2=0
cc_119 C D 0.0351393f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_120 N_C_c_129_n N_A_27_47#_c_224_n 0.0222976f $X=1.475 $Y=1.41 $X2=0 $Y2=0
cc_121 C N_A_27_47#_c_224_n 0.00541755f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_122 N_C_c_129_n N_A_27_47#_c_230_n 0.00159229f $X=1.475 $Y=1.41 $X2=0 $Y2=0
cc_123 C N_A_27_47#_c_230_n 0.014442f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_124 N_C_c_129_n N_VPWR_c_333_n 0.00324396f $X=1.475 $Y=1.41 $X2=0 $Y2=0
cc_125 N_C_c_129_n N_VPWR_c_338_n 0.00700684f $X=1.475 $Y=1.41 $X2=0 $Y2=0
cc_126 N_C_c_129_n N_VPWR_c_330_n 0.0128264f $X=1.475 $Y=1.41 $X2=0 $Y2=0
cc_127 C A_304_47# 0.00980595f $X=1.525 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_128 C N_VGND_c_493_n 0.00481639f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_129 N_C_c_128_n N_VGND_c_497_n 0.00580193f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_130 C N_VGND_c_497_n 0.0078455f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_131 N_C_c_128_n N_VGND_c_502_n 0.0113971f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_132 C N_VGND_c_502_n 0.0091588f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_133 N_D_c_159_n N_A_27_47#_c_196_n 0.0201098f $X=2.08 $Y=0.965 $X2=0 $Y2=0
cc_134 N_D_c_160_n N_A_27_47#_c_196_n 0.0232139f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_135 D N_A_27_47#_c_196_n 0.00478837f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_136 N_D_c_160_n N_A_27_47#_c_203_n 0.0191714f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_137 N_D_c_160_n N_A_27_47#_c_236_n 0.00985619f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_138 N_D_c_160_n N_A_27_47#_c_237_n 0.0207127f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_139 D N_A_27_47#_c_237_n 0.0189039f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_140 N_D_c_160_n N_A_27_47#_c_208_n 0.0034303f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_141 D N_A_27_47#_c_208_n 0.0014507f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_142 N_D_c_160_n N_A_27_47#_c_201_n 0.00155435f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_143 D N_A_27_47#_c_201_n 0.0192253f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_144 N_D_c_160_n N_A_27_47#_c_202_n 0.00286121f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_145 D N_A_27_47#_c_202_n 2.40851e-19 $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_146 N_D_c_160_n N_VPWR_c_334_n 0.00312764f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_147 N_D_c_160_n N_VPWR_c_338_n 0.00702461f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_148 N_D_c_160_n N_VPWR_c_330_n 0.0130442f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_149 D N_X_c_409_n 0.00297167f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_150 D N_VGND_M1005_d 0.00290666f $X=1.985 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_151 N_D_c_159_n N_VGND_c_493_n 0.00962767f $X=2.08 $Y=0.965 $X2=0 $Y2=0
cc_152 N_D_c_160_n N_VGND_c_493_n 0.00196019f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_153 D N_VGND_c_493_n 0.0039159f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_154 N_D_c_159_n N_VGND_c_497_n 0.00438395f $X=2.08 $Y=0.965 $X2=0 $Y2=0
cc_155 D N_VGND_c_497_n 0.0029498f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_156 N_D_c_159_n N_VGND_c_502_n 0.00680522f $X=2.08 $Y=0.965 $X2=0 $Y2=0
cc_157 D N_VGND_c_502_n 0.00614246f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_158 N_A_27_47#_c_224_n N_VPWR_M1002_d 0.00501866f $X=1.605 $Y=1.58 $X2=0
+ $Y2=0
cc_159 N_A_27_47#_c_237_n N_VPWR_M1000_d 0.00794077f $X=2.445 $Y=1.58 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_223_n N_VPWR_c_333_n 0.032721f $X=0.73 $Y=1.96 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_224_n N_VPWR_c_333_n 0.0124807f $X=1.605 $Y=1.58 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_203_n N_VPWR_c_334_n 0.0117861f $X=2.635 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_204_n N_VPWR_c_334_n 9.76587e-19 $X=3.105 $Y=1.41 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_c_237_n N_VPWR_c_334_n 0.018556f $X=2.445 $Y=1.58 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_204_n N_VPWR_c_335_n 0.0055474f $X=3.105 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_205_n N_VPWR_c_335_n 0.011332f $X=3.575 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_206_n N_VPWR_c_335_n 6.15458e-19 $X=4.045 $Y=1.41 $X2=0
+ $Y2=0
cc_168 N_A_27_47#_c_205_n N_VPWR_c_337_n 6.33692e-19 $X=3.575 $Y=1.41 $X2=0
+ $Y2=0
cc_169 N_A_27_47#_c_206_n N_VPWR_c_337_n 0.0152179f $X=4.045 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_236_n N_VPWR_c_338_n 0.0126629f $X=1.71 $Y=1.96 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_203_n N_VPWR_c_340_n 0.00661659f $X=2.635 $Y=1.41 $X2=0
+ $Y2=0
cc_172 N_A_27_47#_c_204_n N_VPWR_c_340_n 0.00673617f $X=3.105 $Y=1.41 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_c_223_n N_VPWR_c_342_n 0.0133725f $X=0.73 $Y=1.96 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_205_n N_VPWR_c_343_n 0.00622633f $X=3.575 $Y=1.41 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_c_206_n N_VPWR_c_343_n 0.00427505f $X=4.045 $Y=1.41 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_M1006_d N_VPWR_c_330_n 0.00508986f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_M1003_d N_VPWR_c_330_n 0.0126813f $X=1.565 $Y=1.485 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_203_n N_VPWR_c_330_n 0.0110154f $X=2.635 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_204_n N_VPWR_c_330_n 0.0118438f $X=3.105 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_205_n N_VPWR_c_330_n 0.0104011f $X=3.575 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_27_47#_c_206_n N_VPWR_c_330_n 0.00732977f $X=4.045 $Y=1.41 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_223_n N_VPWR_c_330_n 0.00801045f $X=0.73 $Y=1.96 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_236_n N_VPWR_c_330_n 0.00724021f $X=1.71 $Y=1.96 $X2=0 $Y2=0
cc_184 N_A_27_47#_c_196_n N_X_c_410_n 0.00283085f $X=2.61 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_27_47#_c_203_n N_X_c_411_n 0.0069886f $X=2.635 $Y=1.41 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_204_n N_X_c_411_n 0.0117859f $X=3.105 $Y=1.41 $X2=0 $Y2=0
cc_187 N_A_27_47#_c_205_n N_X_c_411_n 7.71987e-19 $X=3.575 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_237_n N_X_c_411_n 7.69026e-19 $X=2.445 $Y=1.58 $X2=0 $Y2=0
cc_189 N_A_27_47#_c_197_n N_X_c_415_n 0.0120328f $X=3.08 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_27_47#_c_198_n N_X_c_415_n 0.0128176f $X=3.55 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_27_47#_c_278_p N_X_c_415_n 0.0327997f $X=3.77 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_27_47#_c_202_n N_X_c_415_n 0.00346052f $X=4.045 $Y=1.202 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_196_n N_X_c_409_n 0.00381713f $X=2.61 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_27_47#_c_278_p N_X_c_409_n 0.00935716f $X=3.77 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_202_n N_X_c_409_n 0.00313409f $X=4.045 $Y=1.202 $X2=0 $Y2=0
cc_196 N_A_27_47#_c_204_n N_X_c_422_n 0.0138566f $X=3.105 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_205_n N_X_c_422_n 0.0168647f $X=3.575 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_278_p N_X_c_422_n 0.0404986f $X=3.77 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A_27_47#_c_202_n N_X_c_422_n 0.00645354f $X=4.045 $Y=1.202 $X2=0 $Y2=0
cc_200 N_A_27_47#_c_203_n N_X_c_405_n 0.00140886f $X=2.635 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_204_n N_X_c_405_n 0.00221763f $X=3.105 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A_27_47#_c_237_n N_X_c_405_n 0.0139845f $X=2.445 $Y=1.58 $X2=0 $Y2=0
cc_203 N_A_27_47#_c_208_n N_X_c_405_n 7.55245e-19 $X=2.53 $Y=1.495 $X2=0 $Y2=0
cc_204 N_A_27_47#_c_278_p N_X_c_405_n 0.0167596f $X=3.77 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A_27_47#_c_202_n N_X_c_405_n 0.005429f $X=4.045 $Y=1.202 $X2=0 $Y2=0
cc_206 N_A_27_47#_c_198_n N_X_c_432_n 0.00397179f $X=3.55 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A_27_47#_c_199_n N_X_c_432_n 0.00382799f $X=4.07 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A_27_47#_c_205_n N_X_c_434_n 0.0040177f $X=3.575 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A_27_47#_c_206_n N_X_c_434_n 0.00490547f $X=4.045 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A_27_47#_c_199_n N_X_c_436_n 0.0152217f $X=4.07 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A_27_47#_c_278_p N_X_c_436_n 0.00201745f $X=3.77 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_27_47#_c_202_n N_X_c_436_n 2.27724e-19 $X=4.045 $Y=1.202 $X2=0 $Y2=0
cc_213 N_A_27_47#_c_206_n N_X_c_439_n 0.0238149f $X=4.045 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A_27_47#_c_278_p N_X_c_440_n 0.00957732f $X=3.77 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A_27_47#_c_202_n N_X_c_440_n 0.0040986f $X=4.045 $Y=1.202 $X2=0 $Y2=0
cc_216 N_A_27_47#_c_205_n N_X_c_406_n 0.0028587f $X=3.575 $Y=1.41 $X2=0 $Y2=0
cc_217 N_A_27_47#_c_278_p N_X_c_406_n 0.013101f $X=3.77 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A_27_47#_c_202_n N_X_c_406_n 0.00403689f $X=4.045 $Y=1.202 $X2=0 $Y2=0
cc_219 N_A_27_47#_c_206_n X 0.00304104f $X=4.045 $Y=1.41 $X2=0 $Y2=0
cc_220 N_A_27_47#_c_199_n X 0.021725f $X=4.07 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A_27_47#_c_278_p X 0.0134334f $X=3.77 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A_27_47#_c_200_n A_119_47# 0.00268512f $X=0.61 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_223 N_A_27_47#_c_215_n A_119_47# 0.00437339f $X=0.61 $Y=0.42 $X2=-0.19
+ $Y2=-0.24
cc_224 N_A_27_47#_c_196_n N_VGND_c_493_n 0.00181406f $X=2.61 $Y=0.995 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_201_n N_VGND_c_493_n 0.00249284f $X=2.615 $Y=1.19 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_196_n N_VGND_c_494_n 5.10718e-19 $X=2.61 $Y=0.995 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_197_n N_VGND_c_494_n 0.00713159f $X=3.08 $Y=0.995 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_c_198_n N_VGND_c_494_n 0.0073378f $X=3.55 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A_27_47#_c_199_n N_VGND_c_494_n 4.79843e-19 $X=4.07 $Y=0.995 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_198_n N_VGND_c_496_n 5.27041e-19 $X=3.55 $Y=0.995 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_199_n N_VGND_c_496_n 0.0108274f $X=4.07 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_27_47#_c_215_n N_VGND_c_497_n 0.0322786f $X=0.61 $Y=0.42 $X2=0 $Y2=0
cc_233 N_A_27_47#_c_196_n N_VGND_c_499_n 0.00583607f $X=2.61 $Y=0.995 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_197_n N_VGND_c_499_n 0.00339951f $X=3.08 $Y=0.995 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_198_n N_VGND_c_501_n 0.00339951f $X=3.55 $Y=0.995 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_199_n N_VGND_c_501_n 0.00198008f $X=4.07 $Y=0.995 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_M1012_s N_VGND_c_502_n 0.00272551f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_196_n N_VGND_c_502_n 0.0108044f $X=2.61 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A_27_47#_c_197_n N_VGND_c_502_n 0.00408071f $X=3.08 $Y=0.995 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_c_198_n N_VGND_c_502_n 0.00419605f $X=3.55 $Y=0.995 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_199_n N_VGND_c_502_n 0.00283856f $X=4.07 $Y=0.995 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_215_n N_VGND_c_502_n 0.0198456f $X=0.61 $Y=0.42 $X2=0 $Y2=0
cc_243 N_VPWR_c_330_n N_X_M1007_s 0.00439555f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_244 N_VPWR_c_330_n N_X_M1011_s 0.00647849f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_245 N_VPWR_c_334_n N_X_c_411_n 0.0367474f $X=2.39 $Y=2.02 $X2=0 $Y2=0
cc_246 N_VPWR_c_335_n N_X_c_411_n 0.0384644f $X=3.34 $Y=2 $X2=0 $Y2=0
cc_247 N_VPWR_c_340_n N_X_c_411_n 0.0153803f $X=3.255 $Y=2.72 $X2=0 $Y2=0
cc_248 N_VPWR_c_330_n N_X_c_411_n 0.00939158f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_249 N_VPWR_M1010_d N_X_c_422_n 0.00337289f $X=3.195 $Y=1.485 $X2=0 $Y2=0
cc_250 N_VPWR_c_335_n N_X_c_422_n 0.0147499f $X=3.34 $Y=2 $X2=0 $Y2=0
cc_251 N_VPWR_c_335_n N_X_c_434_n 0.0373402f $X=3.34 $Y=2 $X2=0 $Y2=0
cc_252 N_VPWR_c_337_n N_X_c_434_n 0.0410603f $X=4.28 $Y=2 $X2=0 $Y2=0
cc_253 N_VPWR_c_343_n N_X_c_434_n 0.0118139f $X=4.065 $Y=2.72 $X2=0 $Y2=0
cc_254 N_VPWR_c_330_n N_X_c_434_n 0.00646998f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_255 N_VPWR_M1014_d N_X_c_439_n 2.163e-19 $X=4.135 $Y=1.485 $X2=0 $Y2=0
cc_256 N_VPWR_c_337_n N_X_c_439_n 0.00600363f $X=4.28 $Y=2 $X2=0 $Y2=0
cc_257 N_VPWR_M1014_d N_X_c_407_n 0.00356378f $X=4.135 $Y=1.485 $X2=0 $Y2=0
cc_258 N_VPWR_c_337_n N_X_c_407_n 0.0221374f $X=4.28 $Y=2 $X2=0 $Y2=0
cc_259 N_X_c_415_n N_VGND_M1008_d 0.00437503f $X=3.725 $Y=0.725 $X2=0 $Y2=0
cc_260 N_X_c_403_n N_VGND_M1013_d 0.00291581f $X=4.327 $Y=0.81 $X2=0 $Y2=0
cc_261 X N_VGND_M1013_d 3.27674e-19 $X=4.355 $Y=0.85 $X2=0 $Y2=0
cc_262 N_X_c_410_n N_VGND_c_493_n 0.0173435f $X=2.87 $Y=0.42 $X2=0 $Y2=0
cc_263 N_X_c_415_n N_VGND_c_494_n 0.0198084f $X=3.725 $Y=0.725 $X2=0 $Y2=0
cc_264 N_X_c_432_n N_VGND_c_494_n 0.01316f $X=3.81 $Y=0.42 $X2=0 $Y2=0
cc_265 N_X_c_403_n N_VGND_c_495_n 2.01513e-19 $X=4.327 $Y=0.81 $X2=0 $Y2=0
cc_266 N_X_c_432_n N_VGND_c_496_n 0.0160509f $X=3.81 $Y=0.42 $X2=0 $Y2=0
cc_267 N_X_c_436_n N_VGND_c_496_n 0.00560946f $X=4.2 $Y=0.725 $X2=0 $Y2=0
cc_268 N_X_c_403_n N_VGND_c_496_n 0.0205549f $X=4.327 $Y=0.81 $X2=0 $Y2=0
cc_269 N_X_c_410_n N_VGND_c_499_n 0.0114373f $X=2.87 $Y=0.42 $X2=0 $Y2=0
cc_270 N_X_c_415_n N_VGND_c_499_n 0.0024142f $X=3.725 $Y=0.725 $X2=0 $Y2=0
cc_271 N_X_c_415_n N_VGND_c_501_n 0.00321855f $X=3.725 $Y=0.725 $X2=0 $Y2=0
cc_272 N_X_c_432_n N_VGND_c_501_n 0.0116402f $X=3.81 $Y=0.42 $X2=0 $Y2=0
cc_273 N_X_c_436_n N_VGND_c_501_n 0.0024098f $X=4.2 $Y=0.725 $X2=0 $Y2=0
cc_274 N_X_M1004_s N_VGND_c_502_n 0.00619934f $X=2.685 $Y=0.235 $X2=0 $Y2=0
cc_275 N_X_M1009_s N_VGND_c_502_n 0.00370264f $X=3.625 $Y=0.235 $X2=0 $Y2=0
cc_276 N_X_c_410_n N_VGND_c_502_n 0.00643596f $X=2.87 $Y=0.42 $X2=0 $Y2=0
cc_277 N_X_c_415_n N_VGND_c_502_n 0.0114234f $X=3.725 $Y=0.725 $X2=0 $Y2=0
cc_278 N_X_c_432_n N_VGND_c_502_n 0.00643596f $X=3.81 $Y=0.42 $X2=0 $Y2=0
cc_279 N_X_c_436_n N_VGND_c_502_n 0.00499324f $X=4.2 $Y=0.725 $X2=0 $Y2=0
cc_280 N_X_c_403_n N_VGND_c_502_n 0.00156067f $X=4.327 $Y=0.81 $X2=0 $Y2=0
cc_281 A_119_47# N_VGND_c_502_n 0.0061253f $X=0.595 $Y=0.235 $X2=2.445 $Y2=1.58
cc_282 A_198_47# N_VGND_c_502_n 0.00428291f $X=0.99 $Y=0.235 $X2=0 $Y2=0
cc_283 A_304_47# N_VGND_c_502_n 0.0114506f $X=1.52 $Y=0.235 $X2=0 $Y2=0
