* File: sky130_fd_sc_hdll__nand2b_4.pxi.spice
* Created: Wed Sep  2 08:37:26 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND2B_4%A_N N_A_N_c_89_n N_A_N_M1006_g N_A_N_M1013_g
+ A_N N_A_N_c_88_n PM_SKY130_FD_SC_HDLL__NAND2B_4%A_N
x_PM_SKY130_FD_SC_HDLL__NAND2B_4%A_27_47# N_A_27_47#_M1013_s N_A_27_47#_M1006_s
+ N_A_27_47#_c_130_n N_A_27_47#_M1003_g N_A_27_47#_M1004_g N_A_27_47#_c_131_n
+ N_A_27_47#_M1010_g N_A_27_47#_M1005_g N_A_27_47#_c_132_n N_A_27_47#_M1012_g
+ N_A_27_47#_M1009_g N_A_27_47#_c_133_n N_A_27_47#_M1017_g N_A_27_47#_M1014_g
+ N_A_27_47#_c_121_n N_A_27_47#_c_134_n N_A_27_47#_c_135_n N_A_27_47#_c_122_n
+ N_A_27_47#_c_123_n N_A_27_47#_c_136_n N_A_27_47#_c_124_n N_A_27_47#_c_125_n
+ N_A_27_47#_c_126_n N_A_27_47#_c_127_n N_A_27_47#_c_128_n N_A_27_47#_c_129_n
+ PM_SKY130_FD_SC_HDLL__NAND2B_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NAND2B_4%B N_B_M1000_g N_B_c_252_n N_B_M1002_g
+ N_B_M1001_g N_B_c_253_n N_B_M1008_g N_B_M1007_g N_B_c_254_n N_B_M1011_g
+ N_B_c_255_n N_B_M1016_g N_B_M1015_g B B B B N_B_c_250_n N_B_c_251_n B B
+ N_B_X23_noxref_CONDUCTOR B B PM_SKY130_FD_SC_HDLL__NAND2B_4%B
x_PM_SKY130_FD_SC_HDLL__NAND2B_4%VPWR N_VPWR_M1006_d N_VPWR_M1003_d
+ N_VPWR_M1010_d N_VPWR_M1017_d N_VPWR_M1008_d N_VPWR_M1016_d N_VPWR_c_332_n
+ N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_335_n N_VPWR_c_336_n N_VPWR_c_337_n
+ N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n
+ N_VPWR_c_343_n N_VPWR_c_344_n N_VPWR_c_345_n VPWR N_VPWR_c_346_n
+ N_VPWR_c_347_n N_VPWR_c_331_n PM_SKY130_FD_SC_HDLL__NAND2B_4%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND2B_4%Y N_Y_M1004_s N_Y_M1009_s N_Y_M1003_s
+ N_Y_M1012_s N_Y_M1002_s N_Y_M1011_s N_Y_c_418_n N_Y_c_420_n N_Y_c_437_n
+ N_Y_c_421_n N_Y_c_444_n N_Y_c_419_n N_Y_c_423_n N_Y_c_453_n N_Y_c_424_n
+ N_Y_c_425_n N_Y_c_475_n N_Y_c_426_n Y Y Y PM_SKY130_FD_SC_HDLL__NAND2B_4%Y
x_PM_SKY130_FD_SC_HDLL__NAND2B_4%VGND N_VGND_M1013_d N_VGND_M1000_d
+ N_VGND_M1007_d N_VGND_c_522_n N_VGND_c_523_n N_VGND_c_524_n N_VGND_c_525_n
+ N_VGND_c_526_n N_VGND_c_527_n N_VGND_c_528_n VGND N_VGND_c_529_n
+ N_VGND_c_530_n N_VGND_c_531_n VGND PM_SKY130_FD_SC_HDLL__NAND2B_4%VGND
x_PM_SKY130_FD_SC_HDLL__NAND2B_4%A_225_47# N_A_225_47#_M1004_d
+ N_A_225_47#_M1005_d N_A_225_47#_M1014_d N_A_225_47#_M1001_s
+ N_A_225_47#_M1015_s N_A_225_47#_c_596_n N_A_225_47#_c_597_n
+ N_A_225_47#_c_608_n N_A_225_47#_c_616_n N_A_225_47#_c_598_n
+ N_A_225_47#_c_599_n N_A_225_47#_c_623_n N_A_225_47#_c_600_n
+ N_A_225_47#_c_601_n N_A_225_47#_c_602_n
+ PM_SKY130_FD_SC_HDLL__NAND2B_4%A_225_47#
cc_1 VNB N_A_N_M1013_g 0.0265299f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_2 VNB A_N 0.00738464f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_N_c_88_n 0.0406188f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.212
cc_4 VNB N_A_27_47#_M1004_g 0.0223139f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_5 VNB N_A_27_47#_M1005_g 0.0183647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_M1009_g 0.0183209f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_M1014_g 0.0184382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_121_n 0.0182049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_122_n 0.00117716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_123_n 0.0102254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_124_n 0.00402801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_125_n 6.57408e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_126_n 0.0112315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_127_n 0.00245604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_128_n 0.0328703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_129_n 0.0869195f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_B_M1000_g 0.0182567f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_18 VNB N_B_M1001_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.212
cc_19 VNB N_B_M1007_g 0.0188821f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B_M1015_g 0.0249344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB B 0.0159396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_B_c_250_n 0.084785f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_B_c_251_n 0.0366487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_331_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_Y_c_418_n 0.00572335f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_Y_c_419_n 0.00236899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_522_n 0.00487042f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.212
cc_28 VNB N_VGND_c_523_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_524_n 0.00512401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_525_n 0.0631322f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_526_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_527_n 0.0191455f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_528_n 0.00458858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_529_n 0.0238395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_530_n 0.291301f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_531_n 0.0224167f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_225_47#_c_596_n 0.00232453f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_225_47#_c_597_n 0.00653732f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_225_47#_c_598_n 0.00356157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_225_47#_c_599_n 0.00248276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_225_47#_c_600_n 0.0134401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_225_47#_c_601_n 0.0175671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_225_47#_c_602_n 0.00253093f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VPB N_A_N_c_89_n 0.0233693f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_45 VPB N_A_N_c_88_n 0.0167949f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.212
cc_46 VPB N_A_27_47#_c_130_n 0.0192398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_27_47#_c_131_n 0.0158679f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.212
cc_48 VPB N_A_27_47#_c_132_n 0.0158755f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_27_47#_c_133_n 0.0159631f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_47#_c_134_n 0.0114656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_c_135_n 0.0314532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_47#_c_136_n 0.00133315f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_c_125_n 0.00347213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_47#_c_129_n 0.0267f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_B_c_252_n 0.0160961f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_56 VPB N_B_c_253_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_57 VPB N_B_c_254_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_B_c_255_n 0.0209048f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_B_c_250_n 0.0290861f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_332_n 0.0106419f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_333_n 0.00742108f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_334_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_335_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_336_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_337_n 0.0155402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_338_n 0.043309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_339_n 0.00605347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_340_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_341_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_342_n 0.0209721f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_343_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_344_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_345_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_346_n 0.0215955f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_347_n 0.0326527f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_331_n 0.0489345f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_Y_c_420_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_Y_c_421_n 0.00173134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_Y_c_419_n 0.00133237f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_Y_c_423_n 0.00581507f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_Y_c_424_n 0.00173134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_Y_c_425_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_Y_c_426_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB Y 4.72977e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 N_A_N_c_89_n N_A_27_47#_c_134_n 0.00148112f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_86 A_N N_A_27_47#_c_134_n 0.0255956f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_87 N_A_N_c_88_n N_A_27_47#_c_134_n 0.0069955f $X=0.495 $Y=1.212 $X2=0 $Y2=0
cc_88 N_A_N_c_89_n N_A_27_47#_c_135_n 0.0115092f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A_N_M1013_g N_A_27_47#_c_122_n 0.0140823f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_90 A_N N_A_27_47#_c_122_n 0.001057f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_91 N_A_N_c_88_n N_A_27_47#_c_122_n 5.86027e-19 $X=0.495 $Y=1.212 $X2=0 $Y2=0
cc_92 A_N N_A_27_47#_c_123_n 0.0255857f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_93 N_A_N_c_88_n N_A_27_47#_c_123_n 0.00778107f $X=0.495 $Y=1.212 $X2=0 $Y2=0
cc_94 N_A_N_c_89_n N_A_27_47#_c_136_n 0.0185198f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_95 A_N N_A_27_47#_c_136_n 0.00101487f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_96 N_A_N_c_88_n N_A_27_47#_c_136_n 3.62813e-19 $X=0.495 $Y=1.212 $X2=0 $Y2=0
cc_97 N_A_N_M1013_g N_A_27_47#_c_124_n 0.00598965f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_98 N_A_N_c_89_n N_A_27_47#_c_125_n 0.00131797f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A_N_c_88_n N_A_27_47#_c_125_n 0.00514132f $X=0.495 $Y=1.212 $X2=0 $Y2=0
cc_100 A_N N_A_27_47#_c_127_n 0.0138154f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_101 N_A_N_c_88_n N_A_27_47#_c_127_n 0.00264337f $X=0.495 $Y=1.212 $X2=0 $Y2=0
cc_102 N_A_N_c_88_n N_A_27_47#_c_128_n 0.00571372f $X=0.495 $Y=1.212 $X2=0 $Y2=0
cc_103 N_A_N_c_89_n N_VPWR_c_333_n 0.00361231f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_N_c_89_n N_VPWR_c_339_n 0.00824863f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A_N_c_89_n N_VPWR_c_347_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_106 N_A_N_c_89_n N_VPWR_c_331_n 0.0140376f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_107 N_A_N_M1013_g N_VGND_c_522_n 0.00442456f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_108 N_A_N_M1013_g N_VGND_c_530_n 0.00818709f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_109 N_A_N_M1013_g N_VGND_c_531_n 0.00436487f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_110 N_A_N_M1013_g N_A_225_47#_c_597_n 0.0034126f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_111 N_A_27_47#_M1014_g N_B_M1000_g 0.0160481f $X=2.92 $Y=0.56 $X2=0 $Y2=0
cc_112 N_A_27_47#_c_133_n N_B_c_252_n 0.0216251f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_27_47#_c_129_n B 7.75916e-19 $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_114 N_A_27_47#_c_129_n N_B_c_250_n 0.0160481f $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_115 N_A_27_47#_c_136_n N_VPWR_M1006_d 0.00455976f $X=0.66 $Y=1.555 $X2=-0.19
+ $Y2=-0.24
cc_116 N_A_27_47#_c_130_n N_VPWR_c_333_n 0.00964359f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_117 N_A_27_47#_c_135_n N_VPWR_c_333_n 0.00517368f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_118 N_A_27_47#_c_136_n N_VPWR_c_333_n 0.0176016f $X=0.66 $Y=1.555 $X2=0 $Y2=0
cc_119 N_A_27_47#_c_126_n N_VPWR_c_333_n 0.0256544f $X=2.19 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A_27_47#_c_128_n N_VPWR_c_333_n 0.0063996f $X=1.385 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_27_47#_c_131_n N_VPWR_c_334_n 0.0052072f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A_27_47#_c_132_n N_VPWR_c_334_n 0.004751f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A_27_47#_c_133_n N_VPWR_c_335_n 0.00507848f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_124 N_A_27_47#_c_135_n N_VPWR_c_339_n 0.0425456f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_125 N_A_27_47#_c_136_n N_VPWR_c_339_n 0.0164487f $X=0.66 $Y=1.555 $X2=0 $Y2=0
cc_126 N_A_27_47#_c_126_n N_VPWR_c_339_n 0.00701209f $X=2.19 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A_27_47#_c_130_n N_VPWR_c_340_n 0.00597712f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_128 N_A_27_47#_c_131_n N_VPWR_c_340_n 0.00673617f $X=1.955 $Y=1.41 $X2=0
+ $Y2=0
cc_129 N_A_27_47#_c_132_n N_VPWR_c_342_n 0.00597712f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_130 N_A_27_47#_c_133_n N_VPWR_c_342_n 0.00650846f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_131 N_A_27_47#_c_135_n N_VPWR_c_347_n 0.021418f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_132 N_A_27_47#_M1006_s N_VPWR_c_331_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_133 N_A_27_47#_c_130_n N_VPWR_c_331_n 0.0112769f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_27_47#_c_131_n N_VPWR_c_331_n 0.0118438f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_27_47#_c_132_n N_VPWR_c_331_n 0.00999457f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_136 N_A_27_47#_c_133_n N_VPWR_c_331_n 0.0113873f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A_27_47#_c_135_n N_VPWR_c_331_n 0.0126651f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_138 N_A_27_47#_M1004_g N_Y_c_418_n 0.00630077f $X=1.51 $Y=0.56 $X2=0 $Y2=0
cc_139 N_A_27_47#_M1005_g N_Y_c_418_n 0.0117281f $X=1.98 $Y=0.56 $X2=0 $Y2=0
cc_140 N_A_27_47#_M1009_g N_Y_c_418_n 0.0133472f $X=2.45 $Y=0.56 $X2=0 $Y2=0
cc_141 N_A_27_47#_c_126_n N_Y_c_418_n 0.0629398f $X=2.19 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_27_47#_c_129_n N_Y_c_418_n 0.00646758f $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_143 N_A_27_47#_c_130_n N_Y_c_420_n 0.0046976f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_27_47#_c_131_n N_Y_c_420_n 0.00116723f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_27_47#_c_126_n N_Y_c_420_n 0.0305808f $X=2.19 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A_27_47#_c_129_n N_Y_c_420_n 0.0074788f $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_147 N_A_27_47#_c_130_n N_Y_c_437_n 0.0121679f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_27_47#_c_131_n N_Y_c_437_n 0.0106251f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_27_47#_c_132_n N_Y_c_437_n 6.24674e-19 $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_27_47#_c_131_n N_Y_c_421_n 0.0153933f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_27_47#_c_132_n N_Y_c_421_n 0.0123979f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_27_47#_c_126_n N_Y_c_421_n 0.0339925f $X=2.19 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A_27_47#_c_129_n N_Y_c_421_n 0.00725062f $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_154 N_A_27_47#_M1014_g N_Y_c_444_n 2.07927e-19 $X=2.92 $Y=0.56 $X2=0 $Y2=0
cc_155 N_A_27_47#_c_132_n N_Y_c_419_n 8.88477e-19 $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_27_47#_M1009_g N_Y_c_419_n 0.00317383f $X=2.45 $Y=0.56 $X2=0 $Y2=0
cc_157 N_A_27_47#_c_133_n N_Y_c_419_n 9.57924e-19 $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_27_47#_M1014_g N_Y_c_419_n 0.00336253f $X=2.92 $Y=0.56 $X2=0 $Y2=0
cc_159 N_A_27_47#_c_126_n N_Y_c_419_n 0.0126464f $X=2.19 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_27_47#_c_129_n N_Y_c_419_n 0.0327055f $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_133_n N_Y_c_423_n 0.0188175f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_129_n N_Y_c_423_n 4.93319e-19 $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_133_n N_Y_c_453_n 6.42345e-19 $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_132_n Y 0.00366797f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_133_n Y 0.00118805f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_129_n Y 0.00206076f $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_131_n Y 6.48075e-19 $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_132_n Y 0.0130707f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_133_n Y 0.0116194f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_122_n N_VGND_M1013_d 0.00447436f $X=0.66 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_171 N_A_27_47#_M1004_g N_VGND_c_522_n 0.00188749f $X=1.51 $Y=0.56 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_122_n N_VGND_c_522_n 0.0152582f $X=0.66 $Y=0.81 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_126_n N_VGND_c_522_n 3.11831e-19 $X=2.19 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_27_47#_M1004_g N_VGND_c_525_n 0.00357877f $X=1.51 $Y=0.56 $X2=0 $Y2=0
cc_175 N_A_27_47#_M1005_g N_VGND_c_525_n 0.00357877f $X=1.98 $Y=0.56 $X2=0 $Y2=0
cc_176 N_A_27_47#_M1009_g N_VGND_c_525_n 0.00357877f $X=2.45 $Y=0.56 $X2=0 $Y2=0
cc_177 N_A_27_47#_M1014_g N_VGND_c_525_n 0.00357877f $X=2.92 $Y=0.56 $X2=0 $Y2=0
cc_178 N_A_27_47#_M1013_s N_VGND_c_530_n 0.00258669f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_M1004_g N_VGND_c_530_n 0.00668309f $X=1.51 $Y=0.56 $X2=0 $Y2=0
cc_180 N_A_27_47#_M1005_g N_VGND_c_530_n 0.00548399f $X=1.98 $Y=0.56 $X2=0 $Y2=0
cc_181 N_A_27_47#_M1009_g N_VGND_c_530_n 0.00548399f $X=2.45 $Y=0.56 $X2=0 $Y2=0
cc_182 N_A_27_47#_M1014_g N_VGND_c_530_n 0.00542082f $X=2.92 $Y=0.56 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_121_n N_VGND_c_530_n 0.0128092f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_184 N_A_27_47#_c_122_n N_VGND_c_530_n 0.0058392f $X=0.66 $Y=0.81 $X2=0 $Y2=0
cc_185 N_A_27_47#_c_121_n N_VGND_c_531_n 0.0221535f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_122_n N_VGND_c_531_n 0.00260993f $X=0.66 $Y=0.81 $X2=0 $Y2=0
cc_187 N_A_27_47#_M1004_g N_A_225_47#_c_597_n 0.00459803f $X=1.51 $Y=0.56 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_122_n N_A_225_47#_c_597_n 0.012088f $X=0.66 $Y=0.81 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_126_n N_A_225_47#_c_597_n 0.0201437f $X=2.19 $Y=1.16 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_128_n N_A_225_47#_c_597_n 0.00588114f $X=1.385 $Y=1.16 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_M1004_g N_A_225_47#_c_608_n 0.00999874f $X=1.51 $Y=0.56 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_M1005_g N_A_225_47#_c_608_n 0.00903374f $X=1.98 $Y=0.56 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_M1009_g N_A_225_47#_c_608_n 0.00903374f $X=2.45 $Y=0.56 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_M1014_g N_A_225_47#_c_608_n 0.0137288f $X=2.92 $Y=0.56 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_126_n N_A_225_47#_c_608_n 0.00348133f $X=2.19 $Y=1.16 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_128_n N_A_225_47#_c_608_n 0.00156368f $X=1.385 $Y=1.16 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_129_n N_A_225_47#_c_608_n 4.47034e-19 $X=2.895 $Y=1.217
+ $X2=0 $Y2=0
cc_198 N_A_27_47#_M1014_g N_A_225_47#_c_598_n 9.88618e-19 $X=2.92 $Y=0.56 $X2=0
+ $Y2=0
cc_199 N_B_c_252_n N_VPWR_c_335_n 0.00477308f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_200 N_B_c_253_n N_VPWR_c_336_n 0.0052072f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_201 N_B_c_254_n N_VPWR_c_336_n 0.004751f $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_202 N_B_c_255_n N_VPWR_c_338_n 0.0278322f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_203 B N_VPWR_c_338_n 0.0218086f $X=5.22 $Y=1.105 $X2=0 $Y2=0
cc_204 N_B_c_251_n N_VPWR_c_338_n 0.00557f $X=5.055 $Y=1.16 $X2=0 $Y2=0
cc_205 N_B_c_252_n N_VPWR_c_344_n 0.00597712f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_206 N_B_c_253_n N_VPWR_c_344_n 0.00673617f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_207 N_B_c_254_n N_VPWR_c_346_n 0.00597712f $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_208 N_B_c_255_n N_VPWR_c_346_n 0.00673617f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_209 N_B_c_252_n N_VPWR_c_331_n 0.0100552f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_210 N_B_c_253_n N_VPWR_c_331_n 0.0118438f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_211 N_B_c_254_n N_VPWR_c_331_n 0.00999457f $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_212 N_B_c_255_n N_VPWR_c_331_n 0.0131061f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_213 B N_Y_c_419_n 0.00577061f $X=5.22 $Y=1.105 $X2=0 $Y2=0
cc_214 N_B_c_250_n N_Y_c_419_n 0.00167906f $X=4.89 $Y=1.16 $X2=0 $Y2=0
cc_215 N_B_c_252_n N_Y_c_423_n 0.0127889f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_216 N_B_c_250_n N_Y_c_423_n 3.62694e-19 $X=4.89 $Y=1.16 $X2=0 $Y2=0
cc_217 N_B_c_252_n N_Y_c_453_n 0.0130996f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_218 N_B_c_253_n N_Y_c_453_n 0.0106251f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_219 N_B_c_254_n N_Y_c_453_n 6.24674e-19 $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_220 N_B_c_253_n N_Y_c_424_n 0.0153933f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_221 N_B_c_254_n N_Y_c_424_n 0.0113962f $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_222 B N_Y_c_424_n 0.040258f $X=5.22 $Y=1.105 $X2=0 $Y2=0
cc_223 N_B_c_250_n N_Y_c_424_n 0.00725062f $X=4.89 $Y=1.16 $X2=0 $Y2=0
cc_224 N_B_c_254_n N_Y_c_425_n 0.00292783f $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_225 N_B_c_255_n N_Y_c_425_n 0.0053659f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_226 B N_Y_c_425_n 0.0305808f $X=5.22 $Y=1.105 $X2=0 $Y2=0
cc_227 N_B_c_250_n N_Y_c_425_n 0.00723098f $X=4.89 $Y=1.16 $X2=0 $Y2=0
cc_228 N_B_c_253_n N_Y_c_475_n 6.48386e-19 $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_229 N_B_c_254_n N_Y_c_475_n 0.0130707f $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_230 N_B_c_255_n N_Y_c_475_n 0.0106395f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_231 N_B_c_252_n N_Y_c_426_n 0.00299279f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_232 N_B_c_253_n N_Y_c_426_n 0.00116723f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_233 B N_Y_c_426_n 0.0301956f $X=5.22 $Y=1.105 $X2=0 $Y2=0
cc_234 N_B_c_250_n N_Y_c_426_n 0.0074788f $X=4.89 $Y=1.16 $X2=0 $Y2=0
cc_235 N_B_c_252_n Y 6.38511e-19 $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_236 N_B_M1000_g N_VGND_c_523_n 0.00375751f $X=3.355 $Y=0.56 $X2=0 $Y2=0
cc_237 N_B_M1001_g N_VGND_c_523_n 0.00276126f $X=3.825 $Y=0.56 $X2=0 $Y2=0
cc_238 N_B_M1007_g N_VGND_c_524_n 0.00401373f $X=4.295 $Y=0.56 $X2=0 $Y2=0
cc_239 N_B_M1015_g N_VGND_c_524_n 0.00304644f $X=4.815 $Y=0.56 $X2=0 $Y2=0
cc_240 N_B_M1000_g N_VGND_c_525_n 0.00420723f $X=3.355 $Y=0.56 $X2=0 $Y2=0
cc_241 N_B_M1001_g N_VGND_c_527_n 0.00422241f $X=3.825 $Y=0.56 $X2=0 $Y2=0
cc_242 N_B_M1007_g N_VGND_c_527_n 0.00422241f $X=4.295 $Y=0.56 $X2=0 $Y2=0
cc_243 N_B_M1015_g N_VGND_c_529_n 0.00436487f $X=4.815 $Y=0.56 $X2=0 $Y2=0
cc_244 N_B_M1000_g N_VGND_c_530_n 0.00601917f $X=3.355 $Y=0.56 $X2=0 $Y2=0
cc_245 N_B_M1001_g N_VGND_c_530_n 0.0059505f $X=3.825 $Y=0.56 $X2=0 $Y2=0
cc_246 N_B_M1007_g N_VGND_c_530_n 0.00618861f $X=4.295 $Y=0.56 $X2=0 $Y2=0
cc_247 N_B_M1015_g N_VGND_c_530_n 0.0072574f $X=4.815 $Y=0.56 $X2=0 $Y2=0
cc_248 N_B_M1000_g N_A_225_47#_c_616_n 0.00271016f $X=3.355 $Y=0.56 $X2=0 $Y2=0
cc_249 N_B_M1000_g N_A_225_47#_c_598_n 0.00552237f $X=3.355 $Y=0.56 $X2=0 $Y2=0
cc_250 N_B_M1001_g N_A_225_47#_c_598_n 4.74935e-19 $X=3.825 $Y=0.56 $X2=0 $Y2=0
cc_251 N_B_M1000_g N_A_225_47#_c_599_n 0.0103821f $X=3.355 $Y=0.56 $X2=0 $Y2=0
cc_252 N_B_M1001_g N_A_225_47#_c_599_n 0.0091744f $X=3.825 $Y=0.56 $X2=0 $Y2=0
cc_253 B N_A_225_47#_c_599_n 0.033373f $X=5.22 $Y=1.105 $X2=0 $Y2=0
cc_254 N_B_c_250_n N_A_225_47#_c_599_n 0.00320443f $X=4.89 $Y=1.16 $X2=0 $Y2=0
cc_255 N_B_M1000_g N_A_225_47#_c_623_n 5.22028e-19 $X=3.355 $Y=0.56 $X2=0 $Y2=0
cc_256 N_B_M1001_g N_A_225_47#_c_623_n 0.00641183f $X=3.825 $Y=0.56 $X2=0 $Y2=0
cc_257 N_B_M1007_g N_A_225_47#_c_623_n 0.00707713f $X=4.295 $Y=0.56 $X2=0 $Y2=0
cc_258 N_B_M1015_g N_A_225_47#_c_623_n 8.10277e-19 $X=4.815 $Y=0.56 $X2=0 $Y2=0
cc_259 N_B_M1007_g N_A_225_47#_c_600_n 0.00952594f $X=4.295 $Y=0.56 $X2=0 $Y2=0
cc_260 N_B_M1015_g N_A_225_47#_c_600_n 0.0153414f $X=4.815 $Y=0.56 $X2=0 $Y2=0
cc_261 B N_A_225_47#_c_600_n 0.0785594f $X=5.22 $Y=1.105 $X2=0 $Y2=0
cc_262 N_B_c_250_n N_A_225_47#_c_600_n 0.00434886f $X=4.89 $Y=1.16 $X2=0 $Y2=0
cc_263 N_B_c_251_n N_A_225_47#_c_600_n 0.00773686f $X=5.055 $Y=1.16 $X2=0 $Y2=0
cc_264 N_B_M1015_g N_A_225_47#_c_601_n 0.013644f $X=4.815 $Y=0.56 $X2=0 $Y2=0
cc_265 N_B_M1001_g N_A_225_47#_c_602_n 0.00119366f $X=3.825 $Y=0.56 $X2=0 $Y2=0
cc_266 N_B_M1007_g N_A_225_47#_c_602_n 0.00119366f $X=4.295 $Y=0.56 $X2=0 $Y2=0
cc_267 B N_A_225_47#_c_602_n 0.030602f $X=5.22 $Y=1.105 $X2=0 $Y2=0
cc_268 N_B_c_250_n N_A_225_47#_c_602_n 0.00332f $X=4.89 $Y=1.16 $X2=0 $Y2=0
cc_269 N_VPWR_c_331_n N_Y_M1003_s 0.00231261f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_270 N_VPWR_c_331_n N_Y_M1012_s 0.00231261f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_271 N_VPWR_c_331_n N_Y_M1002_s 0.00231261f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_272 N_VPWR_c_331_n N_Y_M1011_s 0.00231261f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_273 N_VPWR_c_333_n N_Y_c_420_n 0.0181268f $X=1.25 $Y=1.66 $X2=0 $Y2=0
cc_274 N_VPWR_c_333_n N_Y_c_437_n 0.0655186f $X=1.25 $Y=1.66 $X2=0 $Y2=0
cc_275 N_VPWR_c_334_n N_Y_c_437_n 0.0385613f $X=2.19 $Y=2 $X2=0 $Y2=0
cc_276 N_VPWR_c_340_n N_Y_c_437_n 0.0223557f $X=2.105 $Y=2.72 $X2=0 $Y2=0
cc_277 N_VPWR_c_331_n N_Y_c_437_n 0.0140101f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_278 N_VPWR_M1010_d N_Y_c_421_n 0.00180012f $X=2.045 $Y=1.485 $X2=0 $Y2=0
cc_279 N_VPWR_c_334_n N_Y_c_421_n 0.0139097f $X=2.19 $Y=2 $X2=0 $Y2=0
cc_280 N_VPWR_M1017_d N_Y_c_423_n 0.00254806f $X=2.985 $Y=1.485 $X2=0 $Y2=0
cc_281 N_VPWR_c_335_n N_Y_c_423_n 0.0139097f $X=3.145 $Y=2 $X2=0 $Y2=0
cc_282 N_VPWR_c_335_n N_Y_c_453_n 0.0470327f $X=3.145 $Y=2 $X2=0 $Y2=0
cc_283 N_VPWR_c_336_n N_Y_c_453_n 0.0385613f $X=4.085 $Y=2 $X2=0 $Y2=0
cc_284 N_VPWR_c_344_n N_Y_c_453_n 0.0223557f $X=4 $Y=2.72 $X2=0 $Y2=0
cc_285 N_VPWR_c_331_n N_Y_c_453_n 0.0140101f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_286 N_VPWR_M1008_d N_Y_c_424_n 0.00180012f $X=3.94 $Y=1.485 $X2=0 $Y2=0
cc_287 N_VPWR_c_336_n N_Y_c_424_n 0.0139097f $X=4.085 $Y=2 $X2=0 $Y2=0
cc_288 N_VPWR_c_338_n N_Y_c_425_n 0.0103987f $X=5.135 $Y=1.66 $X2=0 $Y2=0
cc_289 N_VPWR_c_336_n N_Y_c_475_n 0.0470327f $X=4.085 $Y=2 $X2=0 $Y2=0
cc_290 N_VPWR_c_338_n N_Y_c_475_n 0.0466499f $X=5.135 $Y=1.66 $X2=0 $Y2=0
cc_291 N_VPWR_c_346_n N_Y_c_475_n 0.0223557f $X=4.97 $Y=2.72 $X2=0 $Y2=0
cc_292 N_VPWR_c_331_n N_Y_c_475_n 0.0140101f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_293 N_VPWR_c_334_n Y 0.0471762f $X=2.19 $Y=2 $X2=0 $Y2=0
cc_294 N_VPWR_c_335_n Y 0.0386782f $X=3.145 $Y=2 $X2=0 $Y2=0
cc_295 N_VPWR_c_342_n Y 0.0233784f $X=3.06 $Y=2.72 $X2=0 $Y2=0
cc_296 N_VPWR_c_331_n Y 0.0145192f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_297 N_Y_M1004_s N_VGND_c_530_n 0.00256987f $X=1.585 $Y=0.235 $X2=0 $Y2=0
cc_298 N_Y_M1009_s N_VGND_c_530_n 0.00256987f $X=2.525 $Y=0.235 $X2=0 $Y2=0
cc_299 N_Y_c_418_n N_A_225_47#_M1005_d 0.00214196f $X=2.575 $Y=0.77 $X2=0 $Y2=0
cc_300 N_Y_c_418_n N_A_225_47#_c_597_n 0.0216726f $X=2.575 $Y=0.77 $X2=0 $Y2=0
cc_301 N_Y_M1004_s N_A_225_47#_c_608_n 0.00401386f $X=1.585 $Y=0.235 $X2=0 $Y2=0
cc_302 N_Y_M1009_s N_A_225_47#_c_608_n 0.00400901f $X=2.525 $Y=0.235 $X2=0 $Y2=0
cc_303 N_Y_c_418_n N_A_225_47#_c_608_n 0.0553961f $X=2.575 $Y=0.77 $X2=0 $Y2=0
cc_304 N_Y_c_444_n N_A_225_47#_c_608_n 0.016068f $X=2.707 $Y=0.905 $X2=0 $Y2=0
cc_305 N_Y_c_444_n N_A_225_47#_c_598_n 0.00783997f $X=2.707 $Y=0.905 $X2=0 $Y2=0
cc_306 N_Y_c_423_n N_A_225_47#_c_598_n 0.00936811f $X=3.4 $Y=1.555 $X2=0 $Y2=0
cc_307 N_Y_c_423_n N_A_225_47#_c_599_n 0.00240615f $X=3.4 $Y=1.555 $X2=0 $Y2=0
cc_308 N_VGND_c_530_n N_A_225_47#_M1004_d 0.00250318f $X=5.29 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_309 N_VGND_c_530_n N_A_225_47#_M1005_d 0.00255381f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_310 N_VGND_c_530_n N_A_225_47#_M1014_d 0.00227252f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_311 N_VGND_c_530_n N_A_225_47#_M1001_s 0.0025535f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_312 N_VGND_c_530_n N_A_225_47#_M1015_s 0.00354473f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_313 N_VGND_c_522_n N_A_225_47#_c_596_n 0.0135471f $X=0.73 $Y=0.38 $X2=0 $Y2=0
cc_314 N_VGND_c_525_n N_A_225_47#_c_596_n 0.017577f $X=3.53 $Y=0 $X2=0 $Y2=0
cc_315 N_VGND_c_530_n N_A_225_47#_c_596_n 0.00961661f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_316 N_VGND_c_522_n N_A_225_47#_c_597_n 0.00470956f $X=0.73 $Y=0.38 $X2=0
+ $Y2=0
cc_317 N_VGND_c_525_n N_A_225_47#_c_608_n 0.0963611f $X=3.53 $Y=0 $X2=0 $Y2=0
cc_318 N_VGND_c_530_n N_A_225_47#_c_608_n 0.0615191f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_319 N_VGND_c_523_n N_A_225_47#_c_616_n 0.0135136f $X=3.615 $Y=0.38 $X2=0
+ $Y2=0
cc_320 N_VGND_c_525_n N_A_225_47#_c_616_n 0.015453f $X=3.53 $Y=0 $X2=0 $Y2=0
cc_321 N_VGND_c_530_n N_A_225_47#_c_616_n 0.00940698f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_322 N_VGND_c_523_n N_A_225_47#_c_598_n 0.00471242f $X=3.615 $Y=0.38 $X2=0
+ $Y2=0
cc_323 N_VGND_M1000_d N_A_225_47#_c_599_n 0.0025045f $X=3.43 $Y=0.235 $X2=0
+ $Y2=0
cc_324 N_VGND_c_523_n N_A_225_47#_c_599_n 0.0127393f $X=3.615 $Y=0.38 $X2=0
+ $Y2=0
cc_325 N_VGND_c_525_n N_A_225_47#_c_599_n 0.00273345f $X=3.53 $Y=0 $X2=0 $Y2=0
cc_326 N_VGND_c_527_n N_A_225_47#_c_599_n 0.00203746f $X=4.47 $Y=0 $X2=0 $Y2=0
cc_327 N_VGND_c_530_n N_A_225_47#_c_599_n 0.00983903f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_328 N_VGND_c_524_n N_A_225_47#_c_623_n 0.0182121f $X=4.555 $Y=0.38 $X2=0
+ $Y2=0
cc_329 N_VGND_c_527_n N_A_225_47#_c_623_n 0.0223596f $X=4.47 $Y=0 $X2=0 $Y2=0
cc_330 N_VGND_c_530_n N_A_225_47#_c_623_n 0.0141302f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_331 N_VGND_M1007_d N_A_225_47#_c_600_n 0.00311775f $X=4.37 $Y=0.235 $X2=0
+ $Y2=0
cc_332 N_VGND_c_524_n N_A_225_47#_c_600_n 0.0166712f $X=4.555 $Y=0.38 $X2=0
+ $Y2=0
cc_333 N_VGND_c_527_n N_A_225_47#_c_600_n 0.00273345f $X=4.47 $Y=0 $X2=0 $Y2=0
cc_334 N_VGND_c_529_n N_A_225_47#_c_600_n 0.00308655f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_335 N_VGND_c_530_n N_A_225_47#_c_600_n 0.0123689f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_336 N_VGND_c_529_n N_A_225_47#_c_601_n 0.0230148f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_337 N_VGND_c_530_n N_A_225_47#_c_601_n 0.0126169f $X=5.29 $Y=0 $X2=0 $Y2=0
