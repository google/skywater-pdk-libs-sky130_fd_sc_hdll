* File: sky130_fd_sc_hdll__inv_12.spice
* Created: Thu Aug 27 19:08:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__inv_12.pex.spice"
.subckt sky130_fd_sc_hdll__inv_12  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.169 PD=0.97 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75005.4
+ A=0.0975 P=1.6 MULT=1
MM1001 N_Y_M1000_d N_A_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7 SB=75004.9
+ A=0.0975 P=1.6 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.1 SB=75004.5
+ A=0.0975 P=1.6 MULT=1
MM1007 N_Y_M1005_d N_A_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.6 SB=75004
+ A=0.0975 P=1.6 MULT=1
MM1011 N_Y_M1011_d N_A_M1011_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.1 SB=75003.5
+ A=0.0975 P=1.6 MULT=1
MM1012 N_Y_M1011_d N_A_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.5 SB=75003.1
+ A=0.0975 P=1.6 MULT=1
MM1013 N_Y_M1013_d N_A_M1013_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003 SB=75002.6
+ A=0.0975 P=1.6 MULT=1
MM1014 N_Y_M1013_d N_A_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.5 SB=75002.1
+ A=0.0975 P=1.6 MULT=1
MM1016 N_Y_M1016_d N_A_M1016_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.9 SB=75001.7
+ A=0.0975 P=1.6 MULT=1
MM1020 N_Y_M1016_d N_A_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.4 SB=75001.2
+ A=0.0975 P=1.6 MULT=1
MM1022 N_Y_M1022_d N_A_M1022_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75004.9
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1023 N_Y_M1022_d N_A_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.1755 PD=1.02 PS=1.84 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75005.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90005.4 A=0.18 P=2.36 MULT=1
MM1003 N_Y_M1002_d N_A_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.6
+ SB=90004.9 A=0.18 P=2.36 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g N_VPWR_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.1
+ SB=90004.4 A=0.18 P=2.36 MULT=1
MM1006 N_Y_M1004_d N_A_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.6
+ SB=90003.9 A=0.18 P=2.36 MULT=1
MM1008 N_Y_M1008_d N_A_M1008_g N_VPWR_M1006_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.1
+ SB=90003.5 A=0.18 P=2.36 MULT=1
MM1009 N_Y_M1008_d N_A_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.5
+ SB=90003 A=0.18 P=2.36 MULT=1
MM1010 N_Y_M1010_d N_A_M1010_g N_VPWR_M1009_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90002.5 A=0.18 P=2.36 MULT=1
MM1015 N_Y_M1010_d N_A_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003.5
+ SB=90002.1 A=0.18 P=2.36 MULT=1
MM1017 N_Y_M1017_d N_A_M1017_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003.9
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1018 N_Y_M1017_d N_A_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90004.4
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1019 N_Y_M1019_d N_A_M1019_g N_VPWR_M1018_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90004.9
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1021 N_Y_M1019_d N_A_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.28 PD=1.29 PS=2.56 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90005.3
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX24_noxref VNB VPB NWDIODE A=10.9461 P=16.85
*
.include "sky130_fd_sc_hdll__inv_12.pxi.spice"
*
.ends
*
*
