* File: sky130_fd_sc_hdll__a2bb2o_1.pex.spice
* Created: Thu Aug 27 18:54:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_1%A_79_21# 1 2 7 9 10 12 15 18 19 21 22 23
+ 25 28 31 35
c91 31 0 1.66009e-19 $X=2.3 $Y=2.275
c92 25 0 6.17718e-20 $X=2.49 $Y=1.895
r93 31 32 0.382445 $w=3.19e-07 $l=1e-08 $layer=LI1_cond $X=2.365 $Y=2.275
+ $X2=2.365 $Y2=2.285
r94 26 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.77 $Y=0.7 $X2=2.77
+ $Y2=0.785
r95 26 28 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.77 $Y=0.7
+ $X2=2.77 $Y2=0.445
r96 25 31 15.7185 $w=3.19e-07 $l=4.38064e-07 $layer=LI1_cond $X=2.49 $Y=1.895
+ $X2=2.365 $Y2=2.275
r97 24 35 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.49 $Y=0.785
+ $X2=2.77 $Y2=0.785
r98 24 25 53.6934 $w=2.18e-07 $l=1.025e-06 $layer=LI1_cond $X=2.49 $Y=0.87
+ $X2=2.49 $Y2=1.895
r99 22 32 4.42298 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=2.13 $Y=2.285
+ $X2=2.365 $Y2=2.285
r100 22 23 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.13 $Y=2.285
+ $X2=1.375 $Y2=2.285
r101 21 23 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.265 $Y=2.2
+ $X2=1.375 $Y2=2.285
r102 20 21 11.7863 $w=2.18e-07 $l=2.25e-07 $layer=LI1_cond $X=1.265 $Y=1.975
+ $X2=1.265 $Y2=2.2
r103 18 20 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.155 $Y=1.89
+ $X2=1.265 $Y2=1.975
r104 18 19 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=1.155 $Y=1.89
+ $X2=0.685 $Y2=1.89
r105 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.16 $X2=0.6 $Y2=1.16
r106 13 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.6 $Y=1.805
+ $X2=0.685 $Y2=1.89
r107 13 15 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=0.6 $Y=1.805
+ $X2=0.6 $Y2=1.16
r108 10 16 47.2262 $w=3.11e-07 $l=2.82843e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.565 $Y2=1.16
r109 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r110 7 16 38.532 $w=3.11e-07 $l=2.07123e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.565 $Y2=1.16
r111 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r112 2 31 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=2.175
+ $Y=2.065 $X2=2.3 $Y2=2.275
r113 1 28 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=2.635
+ $Y=0.235 $X2=2.77 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_1%A1_N 1 3 6 8 9
r30 8 9 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.135 $Y=1.16
+ $X2=1.135 $Y2=1.53
r31 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.08
+ $Y=1.16 $X2=1.08 $Y2=1.16
r32 4 13 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.14 $Y=0.995
+ $X2=1.08 $Y2=1.16
r33 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.14 $Y=0.995 $X2=1.14
+ $Y2=0.445
r34 1 13 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.115 $Y=1.41
+ $X2=1.08 $Y2=1.16
r35 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.115 $Y=1.41
+ $X2=1.115 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_1%A2_N 1 3 6 8 16
c28 1 0 1.5683e-19 $X=1.54 $Y=1.41
r29 8 16 1.06146 $w=3.78e-07 $l=3.5e-08 $layer=LI1_cond $X=1.58 $Y=1.185
+ $X2=1.615 $Y2=1.185
r30 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.58
+ $Y=1.16 $X2=1.58 $Y2=1.16
r31 4 11 39.1718 $w=2.59e-07 $l=1.73292e-07 $layer=POLY_cond $X=1.56 $Y=0.995
+ $X2=1.577 $Y2=1.16
r32 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.56 $Y=0.995 $X2=1.56
+ $Y2=0.445
r33 1 11 51.0578 $w=2.59e-07 $l=2.67862e-07 $layer=POLY_cond $X=1.54 $Y=1.41
+ $X2=1.577 $Y2=1.16
r34 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.54 $Y=1.41 $X2=1.54
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_1%A_243_47# 1 2 8 9 11 14 16 17 20 22 23 24
+ 29 33
c67 33 0 1.5683e-19 $X=1.775 $Y=1.71
c68 29 0 2.83004e-20 $X=2.125 $Y=1.07
c69 9 0 1.62791e-19 $X=2.535 $Y=1.99
r70 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.125
+ $Y=1.07 $X2=2.125 $Y2=1.07
r71 27 29 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.125 $Y=1.545
+ $X2=2.125 $Y2=1.07
r72 26 29 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.125 $Y=0.825
+ $X2=2.125 $Y2=1.07
r73 25 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.86 $Y=1.63
+ $X2=1.775 $Y2=1.63
r74 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.04 $Y=1.63
+ $X2=2.125 $Y2=1.545
r75 24 25 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.04 $Y=1.63
+ $X2=1.86 $Y2=1.63
r76 22 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.04 $Y=0.74
+ $X2=2.125 $Y2=0.825
r77 22 23 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.04 $Y=0.74
+ $X2=1.435 $Y2=0.74
r78 18 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.35 $Y=0.655
+ $X2=1.435 $Y2=0.74
r79 18 20 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.35 $Y=0.655
+ $X2=1.35 $Y2=0.445
r80 16 30 43.1019 $w=4e-07 $l=3.1e-07 $layer=POLY_cond $X=2.435 $Y=1.065
+ $X2=2.125 $Y2=1.065
r81 16 17 5.47071 $w=4e-07 $l=1e-07 $layer=POLY_cond $X=2.435 $Y=1.065 $X2=2.535
+ $Y2=1.065
r82 12 17 38.0281 $w=1.75e-07 $l=2.12132e-07 $layer=POLY_cond $X=2.56 $Y=0.865
+ $X2=2.535 $Y2=1.065
r83 12 14 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.56 $Y=0.865
+ $X2=2.56 $Y2=0.445
r84 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.535 $Y=1.99
+ $X2=2.535 $Y2=2.275
r85 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.535 $Y=1.89 $X2=2.535
+ $Y2=1.99
r86 7 17 38.0281 $w=1.75e-07 $l=2e-07 $layer=POLY_cond $X=2.535 $Y=1.265
+ $X2=2.535 $Y2=1.065
r87 7 8 207.236 $w=2e-07 $l=6.25e-07 $layer=POLY_cond $X=2.535 $Y=1.265
+ $X2=2.535 $Y2=1.89
r88 2 33 600 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=1 $X=1.63
+ $Y=1.485 $X2=1.775 $Y2=1.71
r89 1 20 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.215
+ $Y=0.235 $X2=1.35 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_1%B2 3 6 7 9 10 13
c40 10 0 6.42894e-20 $X=2.985 $Y=1.53
c41 7 0 1.66009e-19 $X=3.005 $Y=1.99
c42 6 0 5.91615e-20 $X=3.005 $Y=1.89
c43 3 0 2.83004e-20 $X=2.98 $Y=0.445
r44 13 16 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.04 $Y=1.47
+ $X2=3.04 $Y2=1.635
r45 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.04 $Y=1.47
+ $X2=3.04 $Y2=1.305
r46 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.04
+ $Y=1.47 $X2=3.04 $Y2=1.47
r47 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.005 $Y=1.99
+ $X2=3.005 $Y2=2.275
r48 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.005 $Y=1.89 $X2=3.005
+ $Y2=1.99
r49 6 16 84.5522 $w=2e-07 $l=2.55e-07 $layer=POLY_cond $X=3.005 $Y=1.89
+ $X2=3.005 $Y2=1.635
r50 3 15 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.98 $Y=0.445
+ $X2=2.98 $Y2=1.305
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_1%B1 3 6 7 9 10 11 12 17
c31 10 0 5.91615e-20 $X=3.525 $Y=0.85
c32 6 0 6.42894e-20 $X=3.485 $Y=1.89
r33 17 20 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.52 $Y=1.16
+ $X2=3.52 $Y2=1.325
r34 17 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.52 $Y=1.16
+ $X2=3.52 $Y2=0.995
r35 11 12 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.495 $Y=1.16
+ $X2=3.495 $Y2=1.53
r36 11 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.52
+ $Y=1.16 $X2=3.52 $Y2=1.16
r37 10 11 13.7407 $w=2.58e-07 $l=3.1e-07 $layer=LI1_cond $X=3.495 $Y=0.85
+ $X2=3.495 $Y2=1.16
r38 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.485 $Y=1.99
+ $X2=3.485 $Y2=2.275
r39 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.485 $Y=1.89 $X2=3.485
+ $Y2=1.99
r40 6 20 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=3.485 $Y=1.89
+ $X2=3.485 $Y2=1.325
r41 3 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.46 $Y=0.445
+ $X2=3.46 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_1%X 1 2 7 8 9
r13 8 9 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.215 $Y=1.87
+ $X2=0.215 $Y2=2.21
r14 8 18 4.87572 $w=2.58e-07 $l=1.1e-07 $layer=LI1_cond $X=0.215 $Y=1.87
+ $X2=0.215 $Y2=1.76
r15 7 18 55.4059 $w=2.58e-07 $l=1.25e-06 $layer=LI1_cond $X=0.215 $Y=0.51
+ $X2=0.215 $Y2=1.76
r16 2 18 300 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.76
r17 1 7 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_1%VPWR 1 2 9 13 16 17 18 20 22 27 37 38 41
r56 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r57 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r58 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r59 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r60 32 35 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r61 32 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r62 31 34 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r63 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r64 29 41 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r65 29 31 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r66 22 41 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r67 20 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r68 20 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r69 18 22 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.235 $Y=2.72
+ $X2=0.515 $Y2=2.72
r70 18 27 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r71 16 34 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=2.72
+ $X2=2.99 $Y2=2.72
r72 16 17 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.155 $Y=2.72
+ $X2=3.285 $Y2=2.72
r73 15 37 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.415 $Y=2.72
+ $X2=3.91 $Y2=2.72
r74 15 17 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.415 $Y=2.72
+ $X2=3.285 $Y2=2.72
r75 11 17 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=2.635
+ $X2=3.285 $Y2=2.72
r76 11 13 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.285 $Y=2.635
+ $X2=3.285 $Y2=2.34
r77 7 41 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r78 7 9 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.32
r79 2 13 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=3.095
+ $Y=2.065 $X2=3.24 $Y2=2.34
r80 1 9 600 $w=1.7e-07 $l=9.04599e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.32
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_1%A_525_413# 1 2 8 9 10 13 18
c39 10 0 1.01019e-19 $X=2.945 $Y=1.92
r40 16 18 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.77 $Y=2.34 $X2=2.86
+ $Y2=2.34
r41 11 13 16.6364 $w=1.78e-07 $l=2.7e-07 $layer=LI1_cond $X=3.725 $Y=2.005
+ $X2=3.725 $Y2=2.275
r42 9 11 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.635 $Y=1.92
+ $X2=3.725 $Y2=2.005
r43 9 10 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.635 $Y=1.92
+ $X2=2.945 $Y2=1.92
r44 8 18 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=2.255
+ $X2=2.86 $Y2=2.34
r45 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.86 $Y=2.005
+ $X2=2.945 $Y2=1.92
r46 7 8 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.86 $Y=2.005 $X2=2.86
+ $Y2=2.255
r47 2 13 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=3.575
+ $Y=2.065 $X2=3.72 $Y2=2.275
r48 1 16 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=2.625
+ $Y=2.065 $X2=2.77 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_1%VGND 1 2 3 10 12 14 16 18 23 30 40 48 51
+ 54
r51 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r52 50 51 9.96101 $w=5.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=0.2
+ $X2=2.39 $Y2=0.2
r53 46 50 3.25249 $w=5.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.07 $Y=0.2
+ $X2=2.225 $Y2=0.2
r54 46 48 14.8922 $w=5.68e-07 $l=4e-07 $layer=LI1_cond $X=2.07 $Y=0.2 $X2=1.67
+ $Y2=0.2
r55 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r56 40 43 11.0886 $w=4.78e-07 $l=4.45e-07 $layer=LI1_cond $X=0.755 $Y=0
+ $X2=0.755 $Y2=0.445
r57 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r58 37 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r59 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r60 34 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r61 34 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r62 33 36 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r63 33 51 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=2.39
+ $Y2=0
r64 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r65 30 53 5.61088 $w=1.7e-07 $l=3.25e-07 $layer=LI1_cond $X=3.49 $Y=0 $X2=3.815
+ $Y2=0
r66 30 36 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=3.49 $Y=0 $X2=3.45
+ $Y2=0
r67 29 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r68 29 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r69 28 48 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.67
+ $Y2=0
r70 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r71 26 40 6.90116 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=0.755
+ $Y2=0
r72 26 28 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=1.61
+ $Y2=0
r73 18 40 6.90116 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.755
+ $Y2=0
r74 16 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r75 16 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r76 14 18 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.235 $Y=0 $X2=0.515
+ $Y2=0
r77 14 23 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r78 10 53 3.19389 $w=4.5e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.715 $Y=0.085
+ $X2=3.815 $Y2=0
r79 10 12 9.16993 $w=4.48e-07 $l=3.45e-07 $layer=LI1_cond $X=3.715 $Y=0.085
+ $X2=3.715 $Y2=0.43
r80 3 12 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=3.535
+ $Y=0.235 $X2=3.72 $Y2=0.43
r81 2 50 91 $w=1.7e-07 $l=6.6742e-07 $layer=licon1_NDIFF $count=2 $X=1.635
+ $Y=0.235 $X2=2.225 $Y2=0.4
r82 1 43 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.445
.ends

