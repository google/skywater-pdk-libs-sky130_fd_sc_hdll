* File: sky130_fd_sc_hdll__sdlclkp_4.pxi.spice
* Created: Thu Aug 27 19:28:25 2020
* 
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_4%SCE N_SCE_c_160_n N_SCE_c_161_n N_SCE_M1007_g
+ N_SCE_M1016_g SCE SCE N_SCE_c_159_n PM_SKY130_FD_SC_HDLL__SDLCLKP_4%SCE
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_4%GATE N_GATE_c_190_n N_GATE_c_191_n
+ N_GATE_M1002_g N_GATE_M1001_g GATE GATE N_GATE_c_188_n N_GATE_c_189_n
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_4%GATE
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_280_21# N_A_280_21#_M1006_d
+ N_A_280_21#_M1023_d N_A_280_21#_M1026_g N_A_280_21#_c_244_n
+ N_A_280_21#_M1005_g N_A_280_21#_c_234_n N_A_280_21#_M1013_g
+ N_A_280_21#_M1008_g N_A_280_21#_c_236_n N_A_280_21#_c_237_n
+ N_A_280_21#_c_238_n N_A_280_21#_c_247_n N_A_280_21#_c_239_n
+ N_A_280_21#_c_248_n N_A_280_21#_c_240_n N_A_280_21#_c_241_n
+ N_A_280_21#_c_242_n N_A_280_21#_c_243_n N_A_280_21#_c_249_n
+ N_A_280_21#_c_258_n N_A_280_21#_c_250_n N_A_280_21#_c_251_n
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_280_21#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_277_243# N_A_277_243#_M1008_s
+ N_A_277_243#_M1013_s N_A_277_243#_c_417_n N_A_277_243#_c_418_n
+ N_A_277_243#_M1012_g N_A_277_243#_c_405_n N_A_277_243#_c_406_n
+ N_A_277_243#_M1000_g N_A_277_243#_c_407_n N_A_277_243#_c_408_n
+ N_A_277_243#_c_409_n N_A_277_243#_c_422_n N_A_277_243#_c_410_n
+ N_A_277_243#_c_411_n N_A_277_243#_c_412_n N_A_277_243#_c_413_n
+ N_A_277_243#_c_414_n N_A_277_243#_c_415_n N_A_277_243#_c_416_n
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_277_243#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_505_315# N_A_505_315#_M1027_d
+ N_A_505_315#_M1019_d N_A_505_315#_c_534_n N_A_505_315#_M1010_g
+ N_A_505_315#_M1015_g N_A_505_315#_c_530_n N_A_505_315#_M1011_g
+ N_A_505_315#_c_531_n N_A_505_315#_M1018_g N_A_505_315#_c_537_n
+ N_A_505_315#_c_532_n N_A_505_315#_c_548_n N_A_505_315#_c_539_n
+ N_A_505_315#_c_533_n N_A_505_315#_c_558_n N_A_505_315#_c_559_n
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_505_315#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_310_47# N_A_310_47#_M1026_d
+ N_A_310_47#_M1012_d N_A_310_47#_c_651_n N_A_310_47#_M1019_g
+ N_A_310_47#_c_652_n N_A_310_47#_M1027_g N_A_310_47#_c_662_n
+ N_A_310_47#_c_660_n N_A_310_47#_c_657_n N_A_310_47#_c_653_n
+ N_A_310_47#_c_654_n N_A_310_47#_c_655_n
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_310_47#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_4%CLK N_CLK_c_744_n N_CLK_M1006_g N_CLK_c_745_n
+ N_CLK_M1023_g N_CLK_c_746_n N_CLK_M1021_g N_CLK_c_747_n N_CLK_M1009_g
+ N_CLK_c_748_n N_CLK_c_749_n N_CLK_c_750_n CLK N_CLK_c_756_n N_CLK_c_751_n CLK
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_4%CLK
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_1125_47# N_A_1125_47#_M1018_s
+ N_A_1125_47#_M1011_d N_A_1125_47#_M1004_g N_A_1125_47#_c_848_n
+ N_A_1125_47#_M1003_g N_A_1125_47#_M1014_g N_A_1125_47#_c_849_n
+ N_A_1125_47#_M1017_g N_A_1125_47#_M1022_g N_A_1125_47#_c_850_n
+ N_A_1125_47#_M1020_g N_A_1125_47#_c_841_n N_A_1125_47#_c_842_n
+ N_A_1125_47#_c_852_n N_A_1125_47#_M1025_g N_A_1125_47#_M1024_g
+ N_A_1125_47#_c_844_n N_A_1125_47#_c_858_n N_A_1125_47#_c_861_n
+ N_A_1125_47#_c_845_n N_A_1125_47#_c_854_n N_A_1125_47#_c_855_n
+ N_A_1125_47#_c_846_n N_A_1125_47#_c_865_n N_A_1125_47#_c_847_n
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_1125_47#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_4%VPWR N_VPWR_M1007_s N_VPWR_M1010_d
+ N_VPWR_M1013_d N_VPWR_M1011_s N_VPWR_M1009_d N_VPWR_M1017_s N_VPWR_M1025_s
+ N_VPWR_c_994_n N_VPWR_c_995_n N_VPWR_c_996_n N_VPWR_c_997_n N_VPWR_c_998_n
+ N_VPWR_c_999_n N_VPWR_c_1000_n N_VPWR_c_1001_n VPWR N_VPWR_c_1002_n
+ N_VPWR_c_1003_n N_VPWR_c_1004_n N_VPWR_c_1005_n N_VPWR_c_1006_n
+ N_VPWR_c_1007_n N_VPWR_c_1008_n N_VPWR_c_1009_n N_VPWR_c_1010_n N_VPWR_c_993_n
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_4%VPWR
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_27_47# N_A_27_47#_M1016_s N_A_27_47#_M1001_d
+ N_A_27_47#_M1002_d N_A_27_47#_c_1115_n N_A_27_47#_c_1116_n N_A_27_47#_c_1117_n
+ N_A_27_47#_c_1118_n N_A_27_47#_c_1128_n N_A_27_47#_c_1137_n
+ N_A_27_47#_c_1141_n PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_4%GCLK N_GCLK_M1004_d N_GCLK_M1022_d
+ N_GCLK_M1003_d N_GCLK_M1020_d N_GCLK_c_1179_n N_GCLK_c_1183_n N_GCLK_c_1187_n
+ N_GCLK_c_1170_n N_GCLK_c_1197_n N_GCLK_c_1174_n N_GCLK_c_1171_n
+ N_GCLK_c_1175_n N_GCLK_c_1212_n N_GCLK_c_1215_n GCLK GCLK GCLK GCLK GCLK GCLK
+ GCLK N_GCLK_c_1178_n N_GCLK_c_1173_n PM_SKY130_FD_SC_HDLL__SDLCLKP_4%GCLK
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_4%VGND N_VGND_M1016_d N_VGND_M1015_d
+ N_VGND_M1008_d N_VGND_M1021_d N_VGND_M1014_s N_VGND_M1024_s N_VGND_c_1259_n
+ N_VGND_c_1260_n N_VGND_c_1261_n N_VGND_c_1262_n N_VGND_c_1263_n
+ N_VGND_c_1264_n N_VGND_c_1265_n N_VGND_c_1266_n VGND N_VGND_c_1267_n
+ N_VGND_c_1268_n N_VGND_c_1269_n N_VGND_c_1270_n N_VGND_c_1271_n
+ N_VGND_c_1272_n N_VGND_c_1273_n N_VGND_c_1274_n
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_4%VGND
cc_1 VNB N_SCE_M1016_g 0.0359819f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB SCE 0.0153286f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_SCE_c_159_n 0.0372557f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_4 VNB N_GATE_M1001_g 0.0287519f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_5 VNB N_GATE_c_188_n 0.0304502f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_6 VNB N_GATE_c_189_n 0.0049723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_280_21#_M1026_g 0.0199677f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_280_21#_c_234_n 0.0264962f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_9 VNB N_A_280_21#_M1008_g 0.0394488f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_280_21#_c_236_n 0.0073558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_280_21#_c_237_n 0.029308f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_280_21#_c_238_n 0.001574f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_280_21#_c_239_n 0.00448089f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_280_21#_c_240_n 0.00288442f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_280_21#_c_241_n 0.00359034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_280_21#_c_242_n 0.00214704f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_280_21#_c_243_n 0.00111161f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_277_243#_c_405_n 0.0158179f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_277_243#_c_406_n 0.00659755f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_277_243#_c_407_n 0.0125358f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_21 VNB N_A_277_243#_c_408_n 0.00834345f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=1.16
cc_22 VNB N_A_277_243#_c_409_n 0.00748877f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=1.53
cc_23 VNB N_A_277_243#_c_410_n 0.00925015f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_277_243#_c_411_n 0.00127255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_277_243#_c_412_n 0.00298048f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_277_243#_c_413_n 0.00716656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_277_243#_c_414_n 0.0306656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_277_243#_c_415_n 0.00252522f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_277_243#_c_416_n 0.0199296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_505_315#_M1015_g 0.0466327f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_505_315#_c_530_n 0.030909f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_32 VNB N_A_505_315#_c_531_n 0.0191045f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_505_315#_c_532_n 0.00951002f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=1.53
cc_34 VNB N_A_505_315#_c_533_n 0.0051523f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_310_47#_c_651_n 0.0328946f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_36 VNB N_A_310_47#_c_652_n 0.0214259f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_37 VNB N_A_310_47#_c_653_n 0.00186374f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=1.53
cc_38 VNB N_A_310_47#_c_654_n 0.00657086f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_310_47#_c_655_n 0.00187427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_CLK_c_744_n 0.0179045f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_41 VNB N_CLK_c_745_n 0.0685883f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.165
cc_42 VNB N_CLK_c_746_n 0.0161966f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_43 VNB N_CLK_c_747_n 0.023896f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_44 VNB N_CLK_c_748_n 0.0114221f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_45 VNB N_CLK_c_749_n 7.01061e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_46 VNB N_CLK_c_750_n 9.64156e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_47 VNB N_CLK_c_751_n 0.00309142f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_1125_47#_M1004_g 0.0188583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_1125_47#_M1014_g 0.0184824f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_50 VNB N_A_1125_47#_M1022_g 0.019851f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_1125_47#_c_841_n 0.0354607f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_1125_47#_c_842_n 0.0596402f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_1125_47#_M1024_g 0.0258397f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1125_47#_c_844_n 0.014941f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_1125_47#_c_845_n 0.00151223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_1125_47#_c_846_n 0.0120421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1125_47#_c_847_n 0.00134722f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VPWR_c_993_n 0.383598f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_27_47#_c_1115_n 0.0141581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_27_47#_c_1116_n 0.00412536f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_61 VNB N_A_27_47#_c_1117_n 0.00642239f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_62 VNB N_A_27_47#_c_1118_n 0.0109465f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_GCLK_c_1170_n 0.00108392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_GCLK_c_1171_n 0.0022023f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=1.53
cc_65 VNB GCLK 0.0207825f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_GCLK_c_1173_n 9.63901e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1259_n 0.00572759f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=1.16
cc_68 VNB N_VGND_c_1260_n 0.00237268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1261_n 0.0126543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1262_n 0.0322355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1263_n 0.00859087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1264_n 0.029725f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1265_n 0.0194567f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1266_n 0.0035381f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1267_n 0.0142754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1268_n 0.0496938f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1269_n 0.0242007f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1270_n 0.00859087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1271_n 0.00663599f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1272_n 0.0299624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1273_n 0.0154142f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1274_n 0.442125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VPB N_SCE_c_160_n 0.0181951f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.67
cc_84 VPB N_SCE_c_161_n 0.0288642f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_85 VPB SCE 0.0189103f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_86 VPB N_SCE_c_159_n 0.0110967f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_87 VPB N_GATE_c_190_n 0.0186063f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.67
cc_88 VPB N_GATE_c_191_n 0.022443f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_89 VPB GATE 0.00673107f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_90 VPB N_GATE_c_188_n 0.00617752f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_91 VPB N_GATE_c_189_n 8.51712e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_280_21#_c_244_n 0.0527117f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_93 VPB N_A_280_21#_c_234_n 0.0150615f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_94 VPB N_A_280_21#_M1013_g 0.0430086f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_280_21#_c_247_n 0.00363029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_280_21#_c_248_n 0.00509907f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_280_21#_c_249_n 0.0181954f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_280_21#_c_250_n 0.00420831f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_280_21#_c_251_n 7.50236e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_277_243#_c_417_n 0.0319868f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_101 VPB N_A_277_243#_c_418_n 0.0245485f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_277_243#_c_405_n 0.0176049f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_277_243#_c_406_n 0.00253968f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_277_243#_c_409_n 0.00477958f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=1.53
cc_105 VPB N_A_277_243#_c_422_n 0.00295943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_505_315#_c_534_n 0.0586229f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_107 VPB N_A_505_315#_M1015_g 0.0172482f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_505_315#_c_530_n 0.0337699f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_109 VPB N_A_505_315#_c_537_n 0.00359991f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_505_315#_c_532_n 0.00409689f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=1.53
cc_111 VPB N_A_505_315#_c_539_n 0.0182773f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_505_315#_c_533_n 0.00735128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_310_47#_c_651_n 0.0357479f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_114 VPB N_A_310_47#_c_657_n 0.0140731f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_310_47#_c_654_n 0.00313868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_310_47#_c_655_n 0.0039199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_CLK_c_745_n 0.0183302f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.165
cc_118 VPB N_CLK_M1023_g 0.0444237f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_119 VPB N_CLK_c_747_n 0.0269316f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_120 VPB N_CLK_c_750_n 0.00130257f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.16
cc_121 VPB N_CLK_c_756_n 0.002495f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_CLK_c_751_n 0.00160768f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_1125_47#_c_848_n 0.0164062f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_124 VPB N_A_1125_47#_c_849_n 0.0161818f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.16
cc_125 VPB N_A_1125_47#_c_850_n 0.0170248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_1125_47#_c_842_n 0.0195582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_1125_47#_c_852_n 0.0217107f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_1125_47#_c_844_n 0.00982363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_1125_47#_c_854_n 0.00160457f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_1125_47#_c_855_n 0.00384171f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_994_n 0.0098838f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_995_n 0.0318655f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=1.53
cc_133 VPB N_VPWR_c_996_n 0.00505078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_997_n 0.00242779f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_998_n 0.0126284f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_999_n 0.0454674f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_1000_n 0.0200898f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_1001_n 0.00359922f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_1002_n 0.0349567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_1003_n 0.0132524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_1004_n 0.0165457f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_1005_n 0.0241871f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_1006_n 0.0531491f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_1007_n 0.0150015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_1008_n 0.0160577f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_1009_n 0.00468713f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_1010_n 0.00631443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_993_n 0.0485335f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_27_47#_c_1116_n 0.00314985f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_150 VPB N_GCLK_c_1174_n 0.00107206f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_GCLK_c_1175_n 0.00262324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB GCLK 0.00115012f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB GCLK 0.00878868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_GCLK_c_1178_n 0.00665993f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 N_SCE_c_160_n N_GATE_c_190_n 0.0156526f $X=0.495 $Y=1.67 $X2=0 $Y2=0
cc_156 N_SCE_c_161_n N_GATE_c_191_n 0.0632062f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_157 N_SCE_M1016_g N_GATE_M1001_g 0.0211542f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_158 N_SCE_c_160_n GATE 3.16667e-19 $X=0.495 $Y=1.67 $X2=0 $Y2=0
cc_159 N_SCE_c_159_n N_GATE_c_188_n 0.0156526f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_160 N_SCE_c_159_n N_GATE_c_189_n 3.16667e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_161 N_SCE_c_161_n N_VPWR_c_995_n 0.00695514f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_162 SCE N_VPWR_c_995_n 0.0242525f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_163 N_SCE_c_159_n N_VPWR_c_995_n 9.03791e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_164 N_SCE_c_161_n N_VPWR_c_1006_n 0.00596194f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_165 N_SCE_c_161_n N_VPWR_c_993_n 0.0107787f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_166 N_SCE_c_160_n N_A_27_47#_c_1116_n 0.0072321f $X=0.495 $Y=1.67 $X2=0 $Y2=0
cc_167 N_SCE_c_161_n N_A_27_47#_c_1116_n 0.014751f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_168 N_SCE_M1016_g N_A_27_47#_c_1116_n 0.0103107f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_169 SCE N_A_27_47#_c_1116_n 0.0521526f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_170 N_SCE_c_159_n N_A_27_47#_c_1116_n 0.00880008f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_171 N_SCE_M1016_g N_A_27_47#_c_1118_n 0.0138857f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_172 SCE N_A_27_47#_c_1118_n 0.0218663f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_173 N_SCE_c_159_n N_A_27_47#_c_1118_n 0.00529806f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_174 N_SCE_c_161_n N_A_27_47#_c_1128_n 0.0089029f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_175 N_SCE_M1016_g N_VGND_c_1267_n 0.00196986f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_176 N_SCE_M1016_g N_VGND_c_1270_n 0.010927f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_177 N_SCE_M1016_g N_VGND_c_1274_n 0.00356708f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_178 N_GATE_M1001_g N_A_280_21#_M1026_g 0.023537f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_179 N_GATE_M1001_g N_A_280_21#_c_236_n 0.00100038f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_180 N_GATE_c_188_n N_A_280_21#_c_236_n 0.0011781f $X=0.99 $Y=1.16 $X2=0 $Y2=0
cc_181 N_GATE_c_189_n N_A_280_21#_c_236_n 0.0311277f $X=0.99 $Y=1.16 $X2=0 $Y2=0
cc_182 N_GATE_c_188_n N_A_280_21#_c_237_n 5.71837e-19 $X=0.99 $Y=1.16 $X2=0
+ $Y2=0
cc_183 N_GATE_c_189_n N_A_280_21#_c_237_n 4.0759e-19 $X=0.99 $Y=1.16 $X2=0 $Y2=0
cc_184 GATE N_A_280_21#_c_258_n 0.00121224f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_185 N_GATE_c_190_n N_A_280_21#_c_250_n 3.08624e-19 $X=0.905 $Y=1.67 $X2=0
+ $Y2=0
cc_186 GATE N_A_280_21#_c_250_n 0.0412461f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_187 N_GATE_c_189_n N_A_280_21#_c_250_n 0.00801744f $X=0.99 $Y=1.16 $X2=0
+ $Y2=0
cc_188 N_GATE_c_191_n N_A_277_243#_c_417_n 0.0118466f $X=0.905 $Y=1.77 $X2=0
+ $Y2=0
cc_189 GATE N_A_277_243#_c_417_n 0.00485806f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_190 N_GATE_c_191_n N_A_277_243#_c_418_n 0.0179326f $X=0.905 $Y=1.77 $X2=0
+ $Y2=0
cc_191 N_GATE_c_190_n N_A_277_243#_c_406_n 0.00594096f $X=0.905 $Y=1.67 $X2=0
+ $Y2=0
cc_192 N_GATE_c_188_n N_A_277_243#_c_406_n 0.00721875f $X=0.99 $Y=1.16 $X2=0
+ $Y2=0
cc_193 N_GATE_c_189_n N_A_277_243#_c_406_n 0.00200251f $X=0.99 $Y=1.16 $X2=0
+ $Y2=0
cc_194 N_GATE_c_191_n N_A_310_47#_c_660_n 2.19657e-19 $X=0.905 $Y=1.77 $X2=0
+ $Y2=0
cc_195 N_GATE_c_191_n N_VPWR_c_1006_n 0.00429453f $X=0.905 $Y=1.77 $X2=0 $Y2=0
cc_196 N_GATE_c_191_n N_VPWR_c_993_n 0.00624845f $X=0.905 $Y=1.77 $X2=0 $Y2=0
cc_197 GATE N_A_27_47#_M1002_d 0.00356778f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_198 N_GATE_c_191_n N_A_27_47#_c_1116_n 0.00518472f $X=0.905 $Y=1.77 $X2=0
+ $Y2=0
cc_199 N_GATE_M1001_g N_A_27_47#_c_1116_n 0.00385412f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_200 N_GATE_c_188_n N_A_27_47#_c_1116_n 0.00498289f $X=0.99 $Y=1.16 $X2=0
+ $Y2=0
cc_201 N_GATE_c_189_n N_A_27_47#_c_1116_n 0.0778137f $X=0.99 $Y=1.16 $X2=0 $Y2=0
cc_202 N_GATE_M1001_g N_A_27_47#_c_1117_n 0.0116943f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_203 N_GATE_c_188_n N_A_27_47#_c_1117_n 0.00479945f $X=0.99 $Y=1.16 $X2=0
+ $Y2=0
cc_204 N_GATE_c_189_n N_A_27_47#_c_1117_n 0.0328353f $X=0.99 $Y=1.16 $X2=0 $Y2=0
cc_205 N_GATE_c_191_n N_A_27_47#_c_1137_n 0.0208897f $X=0.905 $Y=1.77 $X2=0
+ $Y2=0
cc_206 GATE N_A_27_47#_c_1137_n 0.0304797f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_207 N_GATE_M1001_g N_VGND_c_1268_n 0.00422112f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_208 N_GATE_M1001_g N_VGND_c_1270_n 0.00317372f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_209 N_GATE_M1001_g N_VGND_c_1274_n 0.00586994f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_210 N_A_280_21#_c_244_n N_A_277_243#_c_417_n 0.0213218f $X=2.015 $Y=1.99
+ $X2=0 $Y2=0
cc_211 N_A_280_21#_c_250_n N_A_277_243#_c_417_n 0.0153505f $X=1.765 $Y=1.53
+ $X2=0 $Y2=0
cc_212 N_A_280_21#_c_244_n N_A_277_243#_c_418_n 0.0134129f $X=2.015 $Y=1.99
+ $X2=0 $Y2=0
cc_213 N_A_280_21#_c_250_n N_A_277_243#_c_418_n 0.00297656f $X=1.765 $Y=1.53
+ $X2=0 $Y2=0
cc_214 N_A_280_21#_c_244_n N_A_277_243#_c_405_n 0.0218656f $X=2.015 $Y=1.99
+ $X2=0 $Y2=0
cc_215 N_A_280_21#_c_242_n N_A_277_243#_c_405_n 0.010838f $X=1.74 $Y=1.325 $X2=0
+ $Y2=0
cc_216 N_A_280_21#_c_249_n N_A_277_243#_c_405_n 0.0028057f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_217 N_A_280_21#_c_250_n N_A_277_243#_c_405_n 0.00878186f $X=1.765 $Y=1.53
+ $X2=0 $Y2=0
cc_218 N_A_280_21#_c_237_n N_A_277_243#_c_406_n 0.0248786f $X=1.565 $Y=0.87
+ $X2=0 $Y2=0
cc_219 N_A_280_21#_c_242_n N_A_277_243#_c_406_n 0.00531293f $X=1.74 $Y=1.325
+ $X2=0 $Y2=0
cc_220 N_A_280_21#_c_250_n N_A_277_243#_c_406_n 6.29157e-19 $X=1.765 $Y=1.53
+ $X2=0 $Y2=0
cc_221 N_A_280_21#_c_242_n N_A_277_243#_c_407_n 0.00153026f $X=1.74 $Y=1.325
+ $X2=0 $Y2=0
cc_222 N_A_280_21#_M1008_g N_A_277_243#_c_408_n 0.00719655f $X=4.4 $Y=0.445
+ $X2=0 $Y2=0
cc_223 N_A_280_21#_c_240_n N_A_277_243#_c_408_n 0.00782756f $X=5.12 $Y=0.615
+ $X2=0 $Y2=0
cc_224 N_A_280_21#_c_234_n N_A_277_243#_c_409_n 0.00643314f $X=4.375 $Y=1.44
+ $X2=0 $Y2=0
cc_225 N_A_280_21#_M1013_g N_A_277_243#_c_409_n 0.00152654f $X=4.375 $Y=1.835
+ $X2=0 $Y2=0
cc_226 N_A_280_21#_M1008_g N_A_277_243#_c_409_n 0.00225643f $X=4.4 $Y=0.445
+ $X2=0 $Y2=0
cc_227 N_A_280_21#_c_238_n N_A_277_243#_c_409_n 0.0132835f $X=4.525 $Y=1.19
+ $X2=0 $Y2=0
cc_228 N_A_280_21#_c_247_n N_A_277_243#_c_409_n 0.00949266f $X=4.677 $Y=1.495
+ $X2=0 $Y2=0
cc_229 N_A_280_21#_c_239_n N_A_277_243#_c_409_n 0.00563849f $X=4.685 $Y=1.105
+ $X2=0 $Y2=0
cc_230 N_A_280_21#_c_249_n N_A_277_243#_c_409_n 0.0105724f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_231 N_A_280_21#_c_251_n N_A_277_243#_c_409_n 2.64595e-19 $X=4.745 $Y=1.53
+ $X2=0 $Y2=0
cc_232 N_A_280_21#_c_234_n N_A_277_243#_c_422_n 9.91151e-19 $X=4.375 $Y=1.44
+ $X2=0 $Y2=0
cc_233 N_A_280_21#_M1013_g N_A_277_243#_c_422_n 0.00240904f $X=4.375 $Y=1.835
+ $X2=0 $Y2=0
cc_234 N_A_280_21#_c_238_n N_A_277_243#_c_422_n 0.00178751f $X=4.525 $Y=1.19
+ $X2=0 $Y2=0
cc_235 N_A_280_21#_c_247_n N_A_277_243#_c_422_n 0.0108783f $X=4.677 $Y=1.495
+ $X2=0 $Y2=0
cc_236 N_A_280_21#_c_249_n N_A_277_243#_c_422_n 0.00992705f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_237 N_A_280_21#_c_251_n N_A_277_243#_c_422_n 2.76111e-19 $X=4.745 $Y=1.53
+ $X2=0 $Y2=0
cc_238 N_A_280_21#_c_249_n N_A_277_243#_c_410_n 0.0741886f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_239 N_A_280_21#_c_236_n N_A_277_243#_c_411_n 0.00139598f $X=1.565 $Y=0.87
+ $X2=0 $Y2=0
cc_240 N_A_280_21#_c_249_n N_A_277_243#_c_411_n 0.0132091f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_241 N_A_280_21#_c_234_n N_A_277_243#_c_412_n 0.00181472f $X=4.375 $Y=1.44
+ $X2=0 $Y2=0
cc_242 N_A_280_21#_M1008_g N_A_277_243#_c_412_n 0.00655519f $X=4.4 $Y=0.445
+ $X2=0 $Y2=0
cc_243 N_A_280_21#_c_238_n N_A_277_243#_c_412_n 0.00258532f $X=4.525 $Y=1.19
+ $X2=0 $Y2=0
cc_244 N_A_280_21#_c_239_n N_A_277_243#_c_412_n 0.00545288f $X=4.685 $Y=1.105
+ $X2=0 $Y2=0
cc_245 N_A_280_21#_c_240_n N_A_277_243#_c_412_n 0.00140104f $X=5.12 $Y=0.615
+ $X2=0 $Y2=0
cc_246 N_A_280_21#_c_249_n N_A_277_243#_c_412_n 0.0151503f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_247 N_A_280_21#_c_234_n N_A_277_243#_c_413_n 0.00207242f $X=4.375 $Y=1.44
+ $X2=0 $Y2=0
cc_248 N_A_280_21#_M1008_g N_A_277_243#_c_413_n 0.00372865f $X=4.4 $Y=0.445
+ $X2=0 $Y2=0
cc_249 N_A_280_21#_c_238_n N_A_277_243#_c_413_n 0.00527536f $X=4.525 $Y=1.19
+ $X2=0 $Y2=0
cc_250 N_A_280_21#_c_239_n N_A_277_243#_c_413_n 0.00790702f $X=4.685 $Y=1.105
+ $X2=0 $Y2=0
cc_251 N_A_280_21#_c_240_n N_A_277_243#_c_413_n 0.00107367f $X=5.12 $Y=0.615
+ $X2=0 $Y2=0
cc_252 N_A_280_21#_c_249_n N_A_277_243#_c_413_n 9.62924e-19 $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_253 N_A_280_21#_c_236_n N_A_277_243#_c_414_n 0.00753732f $X=1.565 $Y=0.87
+ $X2=0 $Y2=0
cc_254 N_A_280_21#_c_237_n N_A_277_243#_c_414_n 0.0167373f $X=1.565 $Y=0.87
+ $X2=0 $Y2=0
cc_255 N_A_280_21#_c_249_n N_A_277_243#_c_414_n 8.52878e-19 $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_256 N_A_280_21#_c_244_n N_A_277_243#_c_415_n 2.78293e-19 $X=2.015 $Y=1.99
+ $X2=0 $Y2=0
cc_257 N_A_280_21#_c_236_n N_A_277_243#_c_415_n 0.0250263f $X=1.565 $Y=0.87
+ $X2=0 $Y2=0
cc_258 N_A_280_21#_c_237_n N_A_277_243#_c_415_n 2.60115e-19 $X=1.565 $Y=0.87
+ $X2=0 $Y2=0
cc_259 N_A_280_21#_c_249_n N_A_277_243#_c_415_n 0.00617415f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_260 N_A_280_21#_M1026_g N_A_277_243#_c_416_n 0.0135285f $X=1.475 $Y=0.415
+ $X2=0 $Y2=0
cc_261 N_A_280_21#_c_249_n N_A_505_315#_M1019_d 4.4047e-19 $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_262 N_A_280_21#_c_244_n N_A_505_315#_c_534_n 0.0241503f $X=2.015 $Y=1.99
+ $X2=0 $Y2=0
cc_263 N_A_280_21#_c_249_n N_A_505_315#_c_534_n 0.00434872f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_264 N_A_280_21#_c_249_n N_A_505_315#_M1015_g 0.00429637f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_265 N_A_280_21#_c_248_n N_A_505_315#_c_530_n 9.95993e-19 $X=5.21 $Y=1.66
+ $X2=0 $Y2=0
cc_266 N_A_280_21#_c_249_n N_A_505_315#_c_537_n 0.0253368f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_267 N_A_280_21#_c_249_n N_A_505_315#_c_532_n 0.027531f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_268 N_A_280_21#_M1013_g N_A_505_315#_c_548_n 0.00469303f $X=4.375 $Y=1.835
+ $X2=0 $Y2=0
cc_269 N_A_280_21#_M1023_d N_A_505_315#_c_539_n 0.00506445f $X=5.065 $Y=1.515
+ $X2=0 $Y2=0
cc_270 N_A_280_21#_c_234_n N_A_505_315#_c_539_n 9.14009e-19 $X=4.375 $Y=1.44
+ $X2=0 $Y2=0
cc_271 N_A_280_21#_M1013_g N_A_505_315#_c_539_n 0.0164643f $X=4.375 $Y=1.835
+ $X2=0 $Y2=0
cc_272 N_A_280_21#_c_238_n N_A_505_315#_c_539_n 0.0016708f $X=4.525 $Y=1.19
+ $X2=0 $Y2=0
cc_273 N_A_280_21#_c_247_n N_A_505_315#_c_539_n 0.0230625f $X=4.677 $Y=1.495
+ $X2=0 $Y2=0
cc_274 N_A_280_21#_c_248_n N_A_505_315#_c_539_n 0.0311518f $X=5.21 $Y=1.66 $X2=0
+ $Y2=0
cc_275 N_A_280_21#_c_249_n N_A_505_315#_c_539_n 0.0151471f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_276 N_A_280_21#_c_251_n N_A_505_315#_c_539_n 0.00170291f $X=4.745 $Y=1.53
+ $X2=0 $Y2=0
cc_277 N_A_280_21#_c_248_n N_A_505_315#_c_533_n 0.0203634f $X=5.21 $Y=1.66 $X2=0
+ $Y2=0
cc_278 N_A_280_21#_c_249_n N_A_505_315#_c_558_n 0.00655646f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_279 N_A_280_21#_M1013_g N_A_505_315#_c_559_n 0.00335363f $X=4.375 $Y=1.835
+ $X2=0 $Y2=0
cc_280 N_A_280_21#_c_249_n N_A_310_47#_c_651_n 0.00920654f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_281 N_A_280_21#_M1026_g N_A_310_47#_c_662_n 0.0102897f $X=1.475 $Y=0.415
+ $X2=0 $Y2=0
cc_282 N_A_280_21#_c_236_n N_A_310_47#_c_662_n 0.0290877f $X=1.565 $Y=0.87 $X2=0
+ $Y2=0
cc_283 N_A_280_21#_c_237_n N_A_310_47#_c_662_n 0.00131912f $X=1.565 $Y=0.87
+ $X2=0 $Y2=0
cc_284 N_A_280_21#_c_242_n N_A_310_47#_c_662_n 0.00398233f $X=1.74 $Y=1.325
+ $X2=0 $Y2=0
cc_285 N_A_280_21#_c_244_n N_A_310_47#_c_660_n 0.015797f $X=2.015 $Y=1.99 $X2=0
+ $Y2=0
cc_286 N_A_280_21#_c_249_n N_A_310_47#_c_660_n 0.00736596f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_287 N_A_280_21#_c_258_n N_A_310_47#_c_660_n 0.00121651f $X=1.91 $Y=1.53 $X2=0
+ $Y2=0
cc_288 N_A_280_21#_c_250_n N_A_310_47#_c_660_n 0.0341068f $X=1.765 $Y=1.53 $X2=0
+ $Y2=0
cc_289 N_A_280_21#_c_244_n N_A_310_47#_c_657_n 0.00739196f $X=2.015 $Y=1.99
+ $X2=0 $Y2=0
cc_290 N_A_280_21#_c_249_n N_A_310_47#_c_657_n 0.020911f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_291 N_A_280_21#_c_258_n N_A_310_47#_c_657_n 5.20903e-19 $X=1.91 $Y=1.53 $X2=0
+ $Y2=0
cc_292 N_A_280_21#_c_250_n N_A_310_47#_c_657_n 0.0356414f $X=1.765 $Y=1.53 $X2=0
+ $Y2=0
cc_293 N_A_280_21#_c_236_n N_A_310_47#_c_654_n 0.00573093f $X=1.565 $Y=0.87
+ $X2=0 $Y2=0
cc_294 N_A_280_21#_c_242_n N_A_310_47#_c_654_n 0.0121979f $X=1.74 $Y=1.325 $X2=0
+ $Y2=0
cc_295 N_A_280_21#_c_249_n N_A_310_47#_c_654_n 0.00793238f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_296 N_A_280_21#_c_249_n N_A_310_47#_c_655_n 0.00804876f $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_297 N_A_280_21#_M1008_g N_CLK_c_744_n 0.0163343f $X=4.4 $Y=0.445 $X2=-0.19
+ $Y2=-0.24
cc_298 N_A_280_21#_c_240_n N_CLK_c_744_n 0.00757408f $X=5.12 $Y=0.615 $X2=-0.19
+ $Y2=-0.24
cc_299 N_A_280_21#_c_234_n N_CLK_c_745_n 0.0155716f $X=4.375 $Y=1.44 $X2=0 $Y2=0
cc_300 N_A_280_21#_M1008_g N_CLK_c_745_n 0.00391642f $X=4.4 $Y=0.445 $X2=0 $Y2=0
cc_301 N_A_280_21#_c_247_n N_CLK_c_745_n 0.00366095f $X=4.677 $Y=1.495 $X2=0
+ $Y2=0
cc_302 N_A_280_21#_c_239_n N_CLK_c_745_n 0.0111099f $X=4.685 $Y=1.105 $X2=0
+ $Y2=0
cc_303 N_A_280_21#_c_248_n N_CLK_c_745_n 0.00358328f $X=5.21 $Y=1.66 $X2=0 $Y2=0
cc_304 N_A_280_21#_c_240_n N_CLK_c_745_n 0.0208647f $X=5.12 $Y=0.615 $X2=0 $Y2=0
cc_305 N_A_280_21#_c_241_n N_CLK_c_745_n 0.0014877f $X=5.08 $Y=0.465 $X2=0 $Y2=0
cc_306 N_A_280_21#_c_243_n N_CLK_c_745_n 0.00171819f $X=4.677 $Y=1.19 $X2=0
+ $Y2=0
cc_307 N_A_280_21#_c_251_n N_CLK_c_745_n 0.00292718f $X=4.745 $Y=1.53 $X2=0
+ $Y2=0
cc_308 N_A_280_21#_M1013_g N_CLK_M1023_g 0.0345002f $X=4.375 $Y=1.835 $X2=0
+ $Y2=0
cc_309 N_A_280_21#_c_247_n N_CLK_M1023_g 0.00125292f $X=4.677 $Y=1.495 $X2=0
+ $Y2=0
cc_310 N_A_280_21#_c_248_n N_CLK_M1023_g 0.0184633f $X=5.21 $Y=1.66 $X2=0 $Y2=0
cc_311 N_A_280_21#_c_251_n N_CLK_M1023_g 0.00256658f $X=4.745 $Y=1.53 $X2=0
+ $Y2=0
cc_312 N_A_280_21#_c_248_n N_CLK_c_748_n 0.00130707f $X=5.21 $Y=1.66 $X2=0 $Y2=0
cc_313 N_A_280_21#_c_247_n N_CLK_c_749_n 7.24764e-19 $X=4.677 $Y=1.495 $X2=0
+ $Y2=0
cc_314 N_A_280_21#_c_239_n N_CLK_c_749_n 7.23675e-19 $X=4.685 $Y=1.105 $X2=0
+ $Y2=0
cc_315 N_A_280_21#_c_248_n N_CLK_c_749_n 0.00213681f $X=5.21 $Y=1.66 $X2=0 $Y2=0
cc_316 N_A_280_21#_c_240_n N_CLK_c_749_n 0.00106475f $X=5.12 $Y=0.615 $X2=0
+ $Y2=0
cc_317 N_A_280_21#_c_243_n N_CLK_c_749_n 0.00480639f $X=4.677 $Y=1.19 $X2=0
+ $Y2=0
cc_318 N_A_280_21#_c_234_n N_CLK_c_756_n 2.94772e-19 $X=4.375 $Y=1.44 $X2=0
+ $Y2=0
cc_319 N_A_280_21#_c_247_n N_CLK_c_756_n 0.0027056f $X=4.677 $Y=1.495 $X2=0
+ $Y2=0
cc_320 N_A_280_21#_c_239_n N_CLK_c_756_n 0.0064702f $X=4.685 $Y=1.105 $X2=0
+ $Y2=0
cc_321 N_A_280_21#_c_248_n N_CLK_c_756_n 0.0203035f $X=5.21 $Y=1.66 $X2=0 $Y2=0
cc_322 N_A_280_21#_c_240_n N_CLK_c_756_n 0.0103459f $X=5.12 $Y=0.615 $X2=0 $Y2=0
cc_323 N_A_280_21#_c_243_n N_CLK_c_756_n 0.00881118f $X=4.677 $Y=1.19 $X2=0
+ $Y2=0
cc_324 N_A_280_21#_c_240_n N_A_1125_47#_c_846_n 0.0149176f $X=5.12 $Y=0.615
+ $X2=0 $Y2=0
cc_325 N_A_280_21#_c_241_n N_A_1125_47#_c_846_n 0.0299163f $X=5.08 $Y=0.465
+ $X2=0 $Y2=0
cc_326 N_A_280_21#_c_249_n N_VPWR_M1010_d 0.0021747f $X=4.6 $Y=1.53 $X2=0 $Y2=0
cc_327 N_A_280_21#_c_247_n N_VPWR_M1013_d 0.00773199f $X=4.677 $Y=1.495 $X2=0
+ $Y2=0
cc_328 N_A_280_21#_c_249_n N_VPWR_M1013_d 5.63848e-19 $X=4.6 $Y=1.53 $X2=0 $Y2=0
cc_329 N_A_280_21#_M1013_g N_VPWR_c_1002_n 0.0263319f $X=4.375 $Y=1.835 $X2=0
+ $Y2=0
cc_330 N_A_280_21#_c_244_n N_VPWR_c_1006_n 0.00429453f $X=2.015 $Y=1.99 $X2=0
+ $Y2=0
cc_331 N_A_280_21#_c_244_n N_VPWR_c_1007_n 0.00142567f $X=2.015 $Y=1.99 $X2=0
+ $Y2=0
cc_332 N_A_280_21#_c_249_n N_VPWR_c_1007_n 9.58092e-19 $X=4.6 $Y=1.53 $X2=0
+ $Y2=0
cc_333 N_A_280_21#_c_244_n N_VPWR_c_993_n 0.00655921f $X=2.015 $Y=1.99 $X2=0
+ $Y2=0
cc_334 N_A_280_21#_c_250_n N_VPWR_c_993_n 0.0015855f $X=1.765 $Y=1.53 $X2=0
+ $Y2=0
cc_335 N_A_280_21#_M1026_g N_A_27_47#_c_1117_n 0.00341791f $X=1.475 $Y=0.415
+ $X2=0 $Y2=0
cc_336 N_A_280_21#_c_236_n N_A_27_47#_c_1117_n 0.00678546f $X=1.565 $Y=0.87
+ $X2=0 $Y2=0
cc_337 N_A_280_21#_M1026_g N_A_27_47#_c_1141_n 0.00382934f $X=1.475 $Y=0.415
+ $X2=0 $Y2=0
cc_338 N_A_280_21#_c_240_n N_VGND_M1008_d 0.0025681f $X=5.12 $Y=0.615 $X2=0
+ $Y2=0
cc_339 N_A_280_21#_c_234_n N_VGND_c_1263_n 8.44957e-19 $X=4.375 $Y=1.44 $X2=0
+ $Y2=0
cc_340 N_A_280_21#_M1008_g N_VGND_c_1263_n 0.0121645f $X=4.4 $Y=0.445 $X2=0
+ $Y2=0
cc_341 N_A_280_21#_c_238_n N_VGND_c_1263_n 0.0024167f $X=4.525 $Y=1.19 $X2=0
+ $Y2=0
cc_342 N_A_280_21#_c_240_n N_VGND_c_1263_n 0.01501f $X=5.12 $Y=0.615 $X2=0 $Y2=0
cc_343 N_A_280_21#_c_243_n N_VGND_c_1263_n 3.25845e-19 $X=4.677 $Y=1.19 $X2=0
+ $Y2=0
cc_344 N_A_280_21#_M1008_g N_VGND_c_1264_n 0.00273179f $X=4.4 $Y=0.445 $X2=0
+ $Y2=0
cc_345 N_A_280_21#_M1026_g N_VGND_c_1268_n 0.00456464f $X=1.475 $Y=0.415 $X2=0
+ $Y2=0
cc_346 N_A_280_21#_c_240_n N_VGND_c_1272_n 0.00331726f $X=5.12 $Y=0.615 $X2=0
+ $Y2=0
cc_347 N_A_280_21#_c_241_n N_VGND_c_1272_n 0.0165187f $X=5.08 $Y=0.465 $X2=0
+ $Y2=0
cc_348 N_A_280_21#_M1006_d N_VGND_c_1274_n 0.00227267f $X=4.945 $Y=0.235 $X2=0
+ $Y2=0
cc_349 N_A_280_21#_M1026_g N_VGND_c_1274_n 0.00821985f $X=1.475 $Y=0.415 $X2=0
+ $Y2=0
cc_350 N_A_280_21#_M1008_g N_VGND_c_1274_n 0.00469827f $X=4.4 $Y=0.445 $X2=0
+ $Y2=0
cc_351 N_A_280_21#_c_240_n N_VGND_c_1274_n 0.00666319f $X=5.12 $Y=0.615 $X2=0
+ $Y2=0
cc_352 N_A_280_21#_c_241_n N_VGND_c_1274_n 0.00940011f $X=5.08 $Y=0.465 $X2=0
+ $Y2=0
cc_353 N_A_277_243#_c_410_n N_A_505_315#_M1027_d 5.81953e-19 $X=4.09 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_354 N_A_277_243#_c_407_n N_A_505_315#_M1015_g 0.00590251f $X=2.075 $Y=1.215
+ $X2=0 $Y2=0
cc_355 N_A_277_243#_c_410_n N_A_505_315#_M1015_g 0.0049111f $X=4.09 $Y=0.85
+ $X2=0 $Y2=0
cc_356 N_A_277_243#_c_414_n N_A_505_315#_M1015_g 0.00952673f $X=2.11 $Y=0.87
+ $X2=0 $Y2=0
cc_357 N_A_277_243#_c_415_n N_A_505_315#_M1015_g 7.27229e-19 $X=2.11 $Y=0.87
+ $X2=0 $Y2=0
cc_358 N_A_277_243#_c_416_n N_A_505_315#_M1015_g 0.0102362f $X=2.135 $Y=0.705
+ $X2=0 $Y2=0
cc_359 N_A_277_243#_c_408_n N_A_505_315#_c_532_n 0.0925201f $X=4.14 $Y=0.465
+ $X2=0 $Y2=0
cc_360 N_A_277_243#_c_422_n N_A_505_315#_c_532_n 0.00411251f $X=4.14 $Y=1.66
+ $X2=0 $Y2=0
cc_361 N_A_277_243#_c_410_n N_A_505_315#_c_532_n 0.02109f $X=4.09 $Y=0.85 $X2=0
+ $Y2=0
cc_362 N_A_277_243#_c_412_n N_A_505_315#_c_532_n 2.94771e-19 $X=4.235 $Y=0.85
+ $X2=0 $Y2=0
cc_363 N_A_277_243#_M1013_s N_A_505_315#_c_539_n 0.00516605f $X=4.015 $Y=1.515
+ $X2=0 $Y2=0
cc_364 N_A_277_243#_c_422_n N_A_505_315#_c_539_n 0.024093f $X=4.14 $Y=1.66 $X2=0
+ $Y2=0
cc_365 N_A_277_243#_c_422_n N_A_505_315#_c_559_n 0.00889198f $X=4.14 $Y=1.66
+ $X2=0 $Y2=0
cc_366 N_A_277_243#_c_422_n N_A_310_47#_c_651_n 5.9685e-19 $X=4.14 $Y=1.66 $X2=0
+ $Y2=0
cc_367 N_A_277_243#_c_410_n N_A_310_47#_c_651_n 0.00556045f $X=4.09 $Y=0.85
+ $X2=0 $Y2=0
cc_368 N_A_277_243#_c_410_n N_A_310_47#_c_652_n 0.00867797f $X=4.09 $Y=0.85
+ $X2=0 $Y2=0
cc_369 N_A_277_243#_c_406_n N_A_310_47#_c_662_n 7.42828e-19 $X=1.585 $Y=1.29
+ $X2=0 $Y2=0
cc_370 N_A_277_243#_c_410_n N_A_310_47#_c_662_n 0.00173863f $X=4.09 $Y=0.85
+ $X2=0 $Y2=0
cc_371 N_A_277_243#_c_411_n N_A_310_47#_c_662_n 0.0020552f $X=2.42 $Y=0.85 $X2=0
+ $Y2=0
cc_372 N_A_277_243#_c_414_n N_A_310_47#_c_662_n 0.00388987f $X=2.11 $Y=0.87
+ $X2=0 $Y2=0
cc_373 N_A_277_243#_c_415_n N_A_310_47#_c_662_n 0.021194f $X=2.11 $Y=0.87 $X2=0
+ $Y2=0
cc_374 N_A_277_243#_c_416_n N_A_310_47#_c_662_n 0.0134113f $X=2.135 $Y=0.705
+ $X2=0 $Y2=0
cc_375 N_A_277_243#_c_418_n N_A_310_47#_c_660_n 0.00520514f $X=1.485 $Y=1.99
+ $X2=0 $Y2=0
cc_376 N_A_277_243#_c_417_n N_A_310_47#_c_657_n 6.1349e-19 $X=1.485 $Y=1.89
+ $X2=0 $Y2=0
cc_377 N_A_277_243#_c_410_n N_A_310_47#_c_653_n 0.0163852f $X=4.09 $Y=0.85 $X2=0
+ $Y2=0
cc_378 N_A_277_243#_c_411_n N_A_310_47#_c_653_n 0.00275249f $X=2.42 $Y=0.85
+ $X2=0 $Y2=0
cc_379 N_A_277_243#_c_414_n N_A_310_47#_c_653_n 7.76087e-19 $X=2.11 $Y=0.87
+ $X2=0 $Y2=0
cc_380 N_A_277_243#_c_415_n N_A_310_47#_c_653_n 0.0206688f $X=2.11 $Y=0.87 $X2=0
+ $Y2=0
cc_381 N_A_277_243#_c_416_n N_A_310_47#_c_653_n 0.00295563f $X=2.135 $Y=0.705
+ $X2=0 $Y2=0
cc_382 N_A_277_243#_c_407_n N_A_310_47#_c_654_n 0.00427003f $X=2.075 $Y=1.215
+ $X2=0 $Y2=0
cc_383 N_A_277_243#_c_410_n N_A_310_47#_c_654_n 0.00154998f $X=4.09 $Y=0.85
+ $X2=0 $Y2=0
cc_384 N_A_277_243#_c_411_n N_A_310_47#_c_654_n 0.00160742f $X=2.42 $Y=0.85
+ $X2=0 $Y2=0
cc_385 N_A_277_243#_c_414_n N_A_310_47#_c_654_n 0.00154097f $X=2.11 $Y=0.87
+ $X2=0 $Y2=0
cc_386 N_A_277_243#_c_415_n N_A_310_47#_c_654_n 0.0128918f $X=2.11 $Y=0.87 $X2=0
+ $Y2=0
cc_387 N_A_277_243#_c_410_n N_A_310_47#_c_655_n 0.0123454f $X=4.09 $Y=0.85 $X2=0
+ $Y2=0
cc_388 N_A_277_243#_c_418_n N_VPWR_c_1006_n 0.00654912f $X=1.485 $Y=1.99 $X2=0
+ $Y2=0
cc_389 N_A_277_243#_c_418_n N_VPWR_c_993_n 0.0111791f $X=1.485 $Y=1.99 $X2=0
+ $Y2=0
cc_390 N_A_277_243#_c_410_n N_VGND_M1015_d 0.00116391f $X=4.09 $Y=0.85 $X2=0
+ $Y2=0
cc_391 N_A_277_243#_c_410_n N_VGND_c_1259_n 0.0142651f $X=4.09 $Y=0.85 $X2=0
+ $Y2=0
cc_392 N_A_277_243#_c_408_n N_VGND_c_1263_n 0.0149043f $X=4.14 $Y=0.465 $X2=0
+ $Y2=0
cc_393 N_A_277_243#_c_408_n N_VGND_c_1264_n 0.0232287f $X=4.14 $Y=0.465 $X2=0
+ $Y2=0
cc_394 N_A_277_243#_c_416_n N_VGND_c_1268_n 0.00357877f $X=2.135 $Y=0.705 $X2=0
+ $Y2=0
cc_395 N_A_277_243#_M1008_s N_VGND_c_1274_n 0.00235995f $X=4.015 $Y=0.235 $X2=0
+ $Y2=0
cc_396 N_A_277_243#_c_408_n N_VGND_c_1274_n 0.00590194f $X=4.14 $Y=0.465 $X2=0
+ $Y2=0
cc_397 N_A_277_243#_c_410_n N_VGND_c_1274_n 0.0787253f $X=4.09 $Y=0.85 $X2=0
+ $Y2=0
cc_398 N_A_277_243#_c_411_n N_VGND_c_1274_n 0.0148704f $X=2.42 $Y=0.85 $X2=0
+ $Y2=0
cc_399 N_A_277_243#_c_412_n N_VGND_c_1274_n 0.0154936f $X=4.235 $Y=0.85 $X2=0
+ $Y2=0
cc_400 N_A_277_243#_c_413_n N_VGND_c_1274_n 6.80412e-19 $X=4.235 $Y=0.85 $X2=0
+ $Y2=0
cc_401 N_A_277_243#_c_416_n N_VGND_c_1274_n 0.00619361f $X=2.135 $Y=0.705 $X2=0
+ $Y2=0
cc_402 N_A_505_315#_c_534_n N_A_310_47#_c_651_n 0.0122345f $X=2.625 $Y=1.99
+ $X2=0 $Y2=0
cc_403 N_A_505_315#_M1015_g N_A_310_47#_c_651_n 0.0356301f $X=2.76 $Y=0.445
+ $X2=0 $Y2=0
cc_404 N_A_505_315#_c_537_n N_A_310_47#_c_651_n 0.0225684f $X=3.485 $Y=1.77
+ $X2=0 $Y2=0
cc_405 N_A_505_315#_c_532_n N_A_310_47#_c_651_n 0.00694438f $X=3.62 $Y=0.42
+ $X2=0 $Y2=0
cc_406 N_A_505_315#_c_558_n N_A_310_47#_c_651_n 3.5205e-19 $X=2.795 $Y=1.74
+ $X2=0 $Y2=0
cc_407 N_A_505_315#_M1015_g N_A_310_47#_c_652_n 0.0162405f $X=2.76 $Y=0.445
+ $X2=0 $Y2=0
cc_408 N_A_505_315#_c_532_n N_A_310_47#_c_652_n 0.0232068f $X=3.62 $Y=0.42 $X2=0
+ $Y2=0
cc_409 N_A_505_315#_M1015_g N_A_310_47#_c_662_n 0.00845805f $X=2.76 $Y=0.445
+ $X2=0 $Y2=0
cc_410 N_A_505_315#_c_534_n N_A_310_47#_c_660_n 0.00297601f $X=2.625 $Y=1.99
+ $X2=0 $Y2=0
cc_411 N_A_505_315#_c_534_n N_A_310_47#_c_657_n 0.00719955f $X=2.625 $Y=1.99
+ $X2=0 $Y2=0
cc_412 N_A_505_315#_M1015_g N_A_310_47#_c_657_n 0.00512785f $X=2.76 $Y=0.445
+ $X2=0 $Y2=0
cc_413 N_A_505_315#_c_558_n N_A_310_47#_c_657_n 0.0256974f $X=2.795 $Y=1.74
+ $X2=0 $Y2=0
cc_414 N_A_505_315#_M1015_g N_A_310_47#_c_653_n 0.011367f $X=2.76 $Y=0.445 $X2=0
+ $Y2=0
cc_415 N_A_505_315#_c_534_n N_A_310_47#_c_654_n 0.00397597f $X=2.625 $Y=1.99
+ $X2=0 $Y2=0
cc_416 N_A_505_315#_M1015_g N_A_310_47#_c_654_n 0.00603625f $X=2.76 $Y=0.445
+ $X2=0 $Y2=0
cc_417 N_A_505_315#_c_558_n N_A_310_47#_c_654_n 0.00717065f $X=2.795 $Y=1.74
+ $X2=0 $Y2=0
cc_418 N_A_505_315#_M1015_g N_A_310_47#_c_655_n 0.012652f $X=2.76 $Y=0.445 $X2=0
+ $Y2=0
cc_419 N_A_505_315#_c_537_n N_A_310_47#_c_655_n 0.0173332f $X=3.485 $Y=1.77
+ $X2=0 $Y2=0
cc_420 N_A_505_315#_c_532_n N_A_310_47#_c_655_n 0.0255496f $X=3.62 $Y=0.42 $X2=0
+ $Y2=0
cc_421 N_A_505_315#_c_558_n N_A_310_47#_c_655_n 0.00489539f $X=2.795 $Y=1.74
+ $X2=0 $Y2=0
cc_422 N_A_505_315#_c_530_n N_CLK_c_745_n 0.0138439f $X=5.985 $Y=1.41 $X2=0
+ $Y2=0
cc_423 N_A_505_315#_c_531_n N_CLK_c_745_n 0.00666663f $X=6.01 $Y=0.995 $X2=0
+ $Y2=0
cc_424 N_A_505_315#_c_533_n N_CLK_c_745_n 0.00513169f $X=5.79 $Y=1.16 $X2=0
+ $Y2=0
cc_425 N_A_505_315#_c_539_n N_CLK_M1023_g 0.014475f $X=5.565 $Y=2 $X2=0 $Y2=0
cc_426 N_A_505_315#_c_533_n N_CLK_M1023_g 0.0051364f $X=5.79 $Y=1.16 $X2=0 $Y2=0
cc_427 N_A_505_315#_c_531_n N_CLK_c_746_n 0.0391676f $X=6.01 $Y=0.995 $X2=0
+ $Y2=0
cc_428 N_A_505_315#_c_530_n N_CLK_c_747_n 0.0756686f $X=5.985 $Y=1.41 $X2=0
+ $Y2=0
cc_429 N_A_505_315#_c_533_n N_CLK_c_747_n 0.00141065f $X=5.79 $Y=1.16 $X2=0
+ $Y2=0
cc_430 N_A_505_315#_c_530_n N_CLK_c_748_n 0.00963676f $X=5.985 $Y=1.41 $X2=0
+ $Y2=0
cc_431 N_A_505_315#_c_533_n N_CLK_c_748_n 0.0321395f $X=5.79 $Y=1.16 $X2=0 $Y2=0
cc_432 N_A_505_315#_c_533_n N_CLK_c_749_n 0.00220187f $X=5.79 $Y=1.16 $X2=0
+ $Y2=0
cc_433 N_A_505_315#_c_530_n N_CLK_c_750_n 0.00155353f $X=5.985 $Y=1.41 $X2=0
+ $Y2=0
cc_434 N_A_505_315#_c_533_n N_CLK_c_750_n 0.00259415f $X=5.79 $Y=1.16 $X2=0
+ $Y2=0
cc_435 N_A_505_315#_c_530_n N_CLK_c_756_n 4.9817e-19 $X=5.985 $Y=1.41 $X2=0
+ $Y2=0
cc_436 N_A_505_315#_c_533_n N_CLK_c_756_n 0.0184047f $X=5.79 $Y=1.16 $X2=0 $Y2=0
cc_437 N_A_505_315#_c_530_n N_CLK_c_751_n 0.00245047f $X=5.985 $Y=1.41 $X2=0
+ $Y2=0
cc_438 N_A_505_315#_c_533_n N_CLK_c_751_n 0.0185868f $X=5.79 $Y=1.16 $X2=0 $Y2=0
cc_439 N_A_505_315#_c_530_n N_A_1125_47#_c_858_n 4.42321e-19 $X=5.985 $Y=1.41
+ $X2=0 $Y2=0
cc_440 N_A_505_315#_c_531_n N_A_1125_47#_c_858_n 0.0111203f $X=6.01 $Y=0.995
+ $X2=0 $Y2=0
cc_441 N_A_505_315#_c_533_n N_A_1125_47#_c_858_n 0.00390405f $X=5.79 $Y=1.16
+ $X2=0 $Y2=0
cc_442 N_A_505_315#_c_530_n N_A_1125_47#_c_861_n 0.00471521f $X=5.985 $Y=1.41
+ $X2=0 $Y2=0
cc_443 N_A_505_315#_c_530_n N_A_1125_47#_c_846_n 0.00133868f $X=5.985 $Y=1.41
+ $X2=0 $Y2=0
cc_444 N_A_505_315#_c_531_n N_A_1125_47#_c_846_n 0.00537171f $X=6.01 $Y=0.995
+ $X2=0 $Y2=0
cc_445 N_A_505_315#_c_533_n N_A_1125_47#_c_846_n 0.0182023f $X=5.79 $Y=1.16
+ $X2=0 $Y2=0
cc_446 N_A_505_315#_c_530_n N_A_1125_47#_c_865_n 0.00478514f $X=5.985 $Y=1.41
+ $X2=0 $Y2=0
cc_447 N_A_505_315#_c_539_n N_A_1125_47#_c_865_n 0.0120899f $X=5.565 $Y=2 $X2=0
+ $Y2=0
cc_448 N_A_505_315#_c_533_n N_A_1125_47#_c_865_n 0.0284482f $X=5.79 $Y=1.16
+ $X2=0 $Y2=0
cc_449 N_A_505_315#_c_537_n N_VPWR_M1010_d 0.0052367f $X=3.485 $Y=1.77 $X2=0
+ $Y2=0
cc_450 N_A_505_315#_c_539_n N_VPWR_M1013_d 0.00659411f $X=5.565 $Y=2 $X2=0 $Y2=0
cc_451 N_A_505_315#_c_539_n N_VPWR_M1011_s 0.00352128f $X=5.565 $Y=2 $X2=0 $Y2=0
cc_452 N_A_505_315#_c_533_n N_VPWR_M1011_s 0.00244316f $X=5.79 $Y=1.16 $X2=0
+ $Y2=0
cc_453 N_A_505_315#_c_539_n N_VPWR_c_1002_n 0.0243816f $X=5.565 $Y=2 $X2=0 $Y2=0
cc_454 N_A_505_315#_c_548_n N_VPWR_c_1003_n 0.0163045f $X=3.62 $Y=2.205 $X2=0
+ $Y2=0
cc_455 N_A_505_315#_c_539_n N_VPWR_c_1003_n 0.119041f $X=5.565 $Y=2 $X2=0 $Y2=0
cc_456 N_A_505_315#_c_530_n N_VPWR_c_1004_n 0.00622633f $X=5.985 $Y=1.41 $X2=0
+ $Y2=0
cc_457 N_A_505_315#_c_534_n N_VPWR_c_1006_n 0.00173281f $X=2.625 $Y=1.99 $X2=0
+ $Y2=0
cc_458 N_A_505_315#_c_534_n N_VPWR_c_1007_n 0.0293133f $X=2.625 $Y=1.99 $X2=0
+ $Y2=0
cc_459 N_A_505_315#_c_558_n N_VPWR_c_1007_n 0.0489027f $X=2.795 $Y=1.74 $X2=0
+ $Y2=0
cc_460 N_A_505_315#_c_548_n N_VPWR_c_1008_n 0.0137273f $X=3.62 $Y=2.205 $X2=0
+ $Y2=0
cc_461 N_A_505_315#_c_539_n N_VPWR_c_1008_n 0.00252001f $X=5.565 $Y=2 $X2=0
+ $Y2=0
cc_462 N_A_505_315#_c_530_n N_VPWR_c_1009_n 0.00851749f $X=5.985 $Y=1.41 $X2=0
+ $Y2=0
cc_463 N_A_505_315#_M1019_d N_VPWR_c_993_n 0.00237624f $X=3.475 $Y=1.485 $X2=0
+ $Y2=0
cc_464 N_A_505_315#_c_534_n N_VPWR_c_993_n 0.00379144f $X=2.625 $Y=1.99 $X2=0
+ $Y2=0
cc_465 N_A_505_315#_c_530_n N_VPWR_c_993_n 0.0104567f $X=5.985 $Y=1.41 $X2=0
+ $Y2=0
cc_466 N_A_505_315#_c_537_n N_VPWR_c_993_n 0.00668636f $X=3.485 $Y=1.77 $X2=0
+ $Y2=0
cc_467 N_A_505_315#_c_548_n N_VPWR_c_993_n 0.00839556f $X=3.62 $Y=2.205 $X2=0
+ $Y2=0
cc_468 N_A_505_315#_c_539_n N_VPWR_c_993_n 0.0150759f $X=5.565 $Y=2 $X2=0 $Y2=0
cc_469 N_A_505_315#_c_558_n N_VPWR_c_993_n 0.00230693f $X=2.795 $Y=1.74 $X2=0
+ $Y2=0
cc_470 N_A_505_315#_M1015_g N_VGND_c_1259_n 0.00931121f $X=2.76 $Y=0.445 $X2=0
+ $Y2=0
cc_471 N_A_505_315#_c_532_n N_VGND_c_1259_n 0.0310922f $X=3.62 $Y=0.42 $X2=0
+ $Y2=0
cc_472 N_A_505_315#_c_532_n N_VGND_c_1264_n 0.0133789f $X=3.62 $Y=0.42 $X2=0
+ $Y2=0
cc_473 N_A_505_315#_M1015_g N_VGND_c_1268_n 0.00562613f $X=2.76 $Y=0.445 $X2=0
+ $Y2=0
cc_474 N_A_505_315#_c_531_n N_VGND_c_1272_n 0.00196297f $X=6.01 $Y=0.995 $X2=0
+ $Y2=0
cc_475 N_A_505_315#_c_531_n N_VGND_c_1273_n 0.0126251f $X=6.01 $Y=0.995 $X2=0
+ $Y2=0
cc_476 N_A_505_315#_M1027_d N_VGND_c_1274_n 0.00204319f $X=3.485 $Y=0.235 $X2=0
+ $Y2=0
cc_477 N_A_505_315#_M1015_g N_VGND_c_1274_n 0.00739808f $X=2.76 $Y=0.445 $X2=0
+ $Y2=0
cc_478 N_A_505_315#_c_531_n N_VGND_c_1274_n 0.00397487f $X=6.01 $Y=0.995 $X2=0
+ $Y2=0
cc_479 N_A_505_315#_c_532_n N_VGND_c_1274_n 0.00399922f $X=3.62 $Y=0.42 $X2=0
+ $Y2=0
cc_480 N_A_310_47#_c_651_n N_VPWR_c_1003_n 0.00240134f $X=3.385 $Y=1.41 $X2=0
+ $Y2=0
cc_481 N_A_310_47#_c_660_n N_VPWR_c_1006_n 0.0528678f $X=2.235 $Y=2.295 $X2=0
+ $Y2=0
cc_482 N_A_310_47#_c_651_n N_VPWR_c_1007_n 0.0055899f $X=3.385 $Y=1.41 $X2=0
+ $Y2=0
cc_483 N_A_310_47#_c_660_n N_VPWR_c_1007_n 0.0297493f $X=2.235 $Y=2.295 $X2=0
+ $Y2=0
cc_484 N_A_310_47#_c_657_n N_VPWR_c_1007_n 0.00381946f $X=2.32 $Y=2.125 $X2=0
+ $Y2=0
cc_485 N_A_310_47#_c_651_n N_VPWR_c_1008_n 0.0062441f $X=3.385 $Y=1.41 $X2=0
+ $Y2=0
cc_486 N_A_310_47#_M1012_d N_VPWR_c_993_n 0.00279474f $X=1.575 $Y=2.065 $X2=0
+ $Y2=0
cc_487 N_A_310_47#_c_651_n N_VPWR_c_993_n 0.00911855f $X=3.385 $Y=1.41 $X2=0
+ $Y2=0
cc_488 N_A_310_47#_c_660_n N_VPWR_c_993_n 0.0320307f $X=2.235 $Y=2.295 $X2=0
+ $Y2=0
cc_489 N_A_310_47#_c_662_n N_A_27_47#_c_1141_n 0.0219377f $X=2.53 $Y=0.395 $X2=0
+ $Y2=0
cc_490 N_A_310_47#_c_660_n A_421_413# 0.00880176f $X=2.235 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_491 N_A_310_47#_c_657_n A_421_413# 0.00154763f $X=2.32 $Y=2.125 $X2=-0.19
+ $Y2=-0.24
cc_492 N_A_310_47#_c_651_n N_VGND_c_1259_n 0.00488531f $X=3.385 $Y=1.41 $X2=0
+ $Y2=0
cc_493 N_A_310_47#_c_652_n N_VGND_c_1259_n 0.00959698f $X=3.41 $Y=0.995 $X2=0
+ $Y2=0
cc_494 N_A_310_47#_c_662_n N_VGND_c_1259_n 0.0189594f $X=2.53 $Y=0.395 $X2=0
+ $Y2=0
cc_495 N_A_310_47#_c_653_n N_VGND_c_1259_n 0.0170088f $X=2.615 $Y=0.995 $X2=0
+ $Y2=0
cc_496 N_A_310_47#_c_655_n N_VGND_c_1259_n 0.0229573f $X=3.18 $Y=1.16 $X2=0
+ $Y2=0
cc_497 N_A_310_47#_c_652_n N_VGND_c_1264_n 0.00585385f $X=3.41 $Y=0.995 $X2=0
+ $Y2=0
cc_498 N_A_310_47#_c_662_n N_VGND_c_1268_n 0.0740696f $X=2.53 $Y=0.395 $X2=0
+ $Y2=0
cc_499 N_A_310_47#_M1026_d N_VGND_c_1274_n 0.00341601f $X=1.55 $Y=0.235 $X2=0
+ $Y2=0
cc_500 N_A_310_47#_c_652_n N_VGND_c_1274_n 0.00815534f $X=3.41 $Y=0.995 $X2=0
+ $Y2=0
cc_501 N_A_310_47#_c_662_n N_VGND_c_1274_n 0.0337317f $X=2.53 $Y=0.395 $X2=0
+ $Y2=0
cc_502 N_A_310_47#_c_662_n A_425_47# 0.0116337f $X=2.53 $Y=0.395 $X2=-0.19
+ $Y2=-0.24
cc_503 N_A_310_47#_c_653_n A_425_47# 0.00168313f $X=2.615 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_504 N_CLK_c_746_n N_A_1125_47#_M1004_g 0.0218983f $X=6.37 $Y=0.995 $X2=0
+ $Y2=0
cc_505 N_CLK_c_747_n N_A_1125_47#_M1004_g 0.0151521f $X=6.455 $Y=1.41 $X2=0
+ $Y2=0
cc_506 N_CLK_c_751_n N_A_1125_47#_M1004_g 3.03821e-19 $X=6.43 $Y=1.16 $X2=0
+ $Y2=0
cc_507 N_CLK_c_747_n N_A_1125_47#_c_848_n 0.0307988f $X=6.455 $Y=1.41 $X2=0
+ $Y2=0
cc_508 N_CLK_c_747_n N_A_1125_47#_c_842_n 0.00288585f $X=6.455 $Y=1.41 $X2=0
+ $Y2=0
cc_509 N_CLK_c_746_n N_A_1125_47#_c_858_n 0.0108765f $X=6.37 $Y=0.995 $X2=0
+ $Y2=0
cc_510 N_CLK_c_747_n N_A_1125_47#_c_858_n 0.00466689f $X=6.455 $Y=1.41 $X2=0
+ $Y2=0
cc_511 N_CLK_c_748_n N_A_1125_47#_c_858_n 0.00646417f $X=6.1 $Y=1.19 $X2=0 $Y2=0
cc_512 N_CLK_c_750_n N_A_1125_47#_c_858_n 0.00300199f $X=6.245 $Y=1.19 $X2=0
+ $Y2=0
cc_513 N_CLK_c_751_n N_A_1125_47#_c_858_n 0.0223668f $X=6.43 $Y=1.16 $X2=0 $Y2=0
cc_514 N_CLK_c_747_n N_A_1125_47#_c_861_n 0.00479018f $X=6.455 $Y=1.41 $X2=0
+ $Y2=0
cc_515 N_CLK_c_746_n N_A_1125_47#_c_845_n 0.00398268f $X=6.37 $Y=0.995 $X2=0
+ $Y2=0
cc_516 N_CLK_c_747_n N_A_1125_47#_c_845_n 4.08409e-19 $X=6.455 $Y=1.41 $X2=0
+ $Y2=0
cc_517 N_CLK_c_751_n N_A_1125_47#_c_845_n 0.00441122f $X=6.43 $Y=1.16 $X2=0
+ $Y2=0
cc_518 N_CLK_c_747_n N_A_1125_47#_c_854_n 0.0036352f $X=6.455 $Y=1.41 $X2=0
+ $Y2=0
cc_519 N_CLK_c_751_n N_A_1125_47#_c_854_n 6.41528e-19 $X=6.43 $Y=1.16 $X2=0
+ $Y2=0
cc_520 N_CLK_c_744_n N_A_1125_47#_c_846_n 3.56754e-19 $X=4.87 $Y=0.73 $X2=0
+ $Y2=0
cc_521 N_CLK_c_745_n N_A_1125_47#_c_846_n 7.62216e-19 $X=4.975 $Y=1.44 $X2=0
+ $Y2=0
cc_522 N_CLK_c_748_n N_A_1125_47#_c_846_n 0.00824021f $X=6.1 $Y=1.19 $X2=0 $Y2=0
cc_523 N_CLK_c_747_n N_A_1125_47#_c_865_n 0.0318428f $X=6.455 $Y=1.41 $X2=0
+ $Y2=0
cc_524 N_CLK_c_750_n N_A_1125_47#_c_865_n 0.0020289f $X=6.245 $Y=1.19 $X2=0
+ $Y2=0
cc_525 N_CLK_c_751_n N_A_1125_47#_c_865_n 0.0301791f $X=6.43 $Y=1.16 $X2=0 $Y2=0
cc_526 N_CLK_c_747_n N_A_1125_47#_c_847_n 0.00195414f $X=6.455 $Y=1.41 $X2=0
+ $Y2=0
cc_527 N_CLK_c_750_n N_A_1125_47#_c_847_n 0.00127984f $X=6.245 $Y=1.19 $X2=0
+ $Y2=0
cc_528 N_CLK_c_751_n N_A_1125_47#_c_847_n 0.0206769f $X=6.43 $Y=1.16 $X2=0 $Y2=0
cc_529 N_CLK_c_747_n N_VPWR_c_996_n 0.00181837f $X=6.455 $Y=1.41 $X2=0 $Y2=0
cc_530 N_CLK_M1023_g N_VPWR_c_1002_n 0.0274117f $X=4.975 $Y=1.835 $X2=0 $Y2=0
cc_531 N_CLK_c_747_n N_VPWR_c_1004_n 0.00510113f $X=6.455 $Y=1.41 $X2=0 $Y2=0
cc_532 N_CLK_c_747_n N_VPWR_c_1009_n 5.70534e-19 $X=6.455 $Y=1.41 $X2=0 $Y2=0
cc_533 N_CLK_c_747_n N_VPWR_c_993_n 0.0067498f $X=6.455 $Y=1.41 $X2=0 $Y2=0
cc_534 N_CLK_c_744_n N_VGND_c_1263_n 0.00317372f $X=4.87 $Y=0.73 $X2=0 $Y2=0
cc_535 N_CLK_c_744_n N_VGND_c_1272_n 0.00422112f $X=4.87 $Y=0.73 $X2=0 $Y2=0
cc_536 N_CLK_c_745_n N_VGND_c_1272_n 0.00230382f $X=4.975 $Y=1.44 $X2=0 $Y2=0
cc_537 N_CLK_c_746_n N_VGND_c_1273_n 0.0176987f $X=6.37 $Y=0.995 $X2=0 $Y2=0
cc_538 N_CLK_c_744_n N_VGND_c_1274_n 0.00711082f $X=4.87 $Y=0.73 $X2=0 $Y2=0
cc_539 N_CLK_c_745_n N_VGND_c_1274_n 0.00262886f $X=4.975 $Y=1.44 $X2=0 $Y2=0
cc_540 N_A_1125_47#_c_854_n N_VPWR_M1009_d 3.90052e-19 $X=6.825 $Y=1.495 $X2=0
+ $Y2=0
cc_541 N_A_1125_47#_c_865_n N_VPWR_M1009_d 0.00848749f $X=6.825 $Y=1.79 $X2=0
+ $Y2=0
cc_542 N_A_1125_47#_c_848_n N_VPWR_c_996_n 0.00327647f $X=6.98 $Y=1.41 $X2=0
+ $Y2=0
cc_543 N_A_1125_47#_c_865_n N_VPWR_c_996_n 0.0191719f $X=6.825 $Y=1.79 $X2=0
+ $Y2=0
cc_544 N_A_1125_47#_c_849_n N_VPWR_c_997_n 0.00558536f $X=7.45 $Y=1.41 $X2=0
+ $Y2=0
cc_545 N_A_1125_47#_c_850_n N_VPWR_c_997_n 0.0148874f $X=7.92 $Y=1.41 $X2=0
+ $Y2=0
cc_546 N_A_1125_47#_c_842_n N_VPWR_c_997_n 5.58063e-19 $X=8.02 $Y=1.16 $X2=0
+ $Y2=0
cc_547 N_A_1125_47#_c_852_n N_VPWR_c_997_n 0.00113408f $X=8.525 $Y=1.41 $X2=0
+ $Y2=0
cc_548 N_A_1125_47#_c_852_n N_VPWR_c_999_n 0.0246404f $X=8.525 $Y=1.41 $X2=0
+ $Y2=0
cc_549 N_A_1125_47#_c_848_n N_VPWR_c_1000_n 0.00681089f $X=6.98 $Y=1.41 $X2=0
+ $Y2=0
cc_550 N_A_1125_47#_c_849_n N_VPWR_c_1000_n 0.00673617f $X=7.45 $Y=1.41 $X2=0
+ $Y2=0
cc_551 N_A_1125_47#_c_865_n N_VPWR_c_1000_n 3.86084e-19 $X=6.825 $Y=1.79 $X2=0
+ $Y2=0
cc_552 N_A_1125_47#_c_861_n N_VPWR_c_1004_n 0.0113299f $X=6.22 $Y=2.085 $X2=0
+ $Y2=0
cc_553 N_A_1125_47#_c_865_n N_VPWR_c_1004_n 0.00392738f $X=6.825 $Y=1.79 $X2=0
+ $Y2=0
cc_554 N_A_1125_47#_c_850_n N_VPWR_c_1005_n 0.00622633f $X=7.92 $Y=1.41 $X2=0
+ $Y2=0
cc_555 N_A_1125_47#_c_852_n N_VPWR_c_1005_n 0.00461082f $X=8.525 $Y=1.41 $X2=0
+ $Y2=0
cc_556 N_A_1125_47#_c_861_n N_VPWR_c_1009_n 0.013449f $X=6.22 $Y=2.085 $X2=0
+ $Y2=0
cc_557 N_A_1125_47#_M1011_d N_VPWR_c_993_n 0.00462612f $X=6.075 $Y=1.485 $X2=0
+ $Y2=0
cc_558 N_A_1125_47#_c_848_n N_VPWR_c_993_n 0.0119747f $X=6.98 $Y=1.41 $X2=0
+ $Y2=0
cc_559 N_A_1125_47#_c_849_n N_VPWR_c_993_n 0.0118847f $X=7.45 $Y=1.41 $X2=0
+ $Y2=0
cc_560 N_A_1125_47#_c_850_n N_VPWR_c_993_n 0.0107955f $X=7.92 $Y=1.41 $X2=0
+ $Y2=0
cc_561 N_A_1125_47#_c_852_n N_VPWR_c_993_n 0.00827986f $X=8.525 $Y=1.41 $X2=0
+ $Y2=0
cc_562 N_A_1125_47#_c_861_n N_VPWR_c_993_n 0.00637602f $X=6.22 $Y=2.085 $X2=0
+ $Y2=0
cc_563 N_A_1125_47#_c_865_n N_VPWR_c_993_n 0.00878273f $X=6.825 $Y=1.79 $X2=0
+ $Y2=0
cc_564 N_A_1125_47#_M1004_g N_GCLK_c_1179_n 0.00451142f $X=6.955 $Y=0.56 $X2=0
+ $Y2=0
cc_565 N_A_1125_47#_M1014_g N_GCLK_c_1179_n 0.0060766f $X=7.425 $Y=0.56 $X2=0
+ $Y2=0
cc_566 N_A_1125_47#_M1022_g N_GCLK_c_1179_n 7.5358e-19 $X=7.895 $Y=0.56 $X2=0
+ $Y2=0
cc_567 N_A_1125_47#_c_858_n N_GCLK_c_1179_n 0.00658218f $X=6.74 $Y=0.7 $X2=0
+ $Y2=0
cc_568 N_A_1125_47#_c_848_n N_GCLK_c_1183_n 0.00666419f $X=6.98 $Y=1.41 $X2=0
+ $Y2=0
cc_569 N_A_1125_47#_c_849_n N_GCLK_c_1183_n 0.0117872f $X=7.45 $Y=1.41 $X2=0
+ $Y2=0
cc_570 N_A_1125_47#_c_850_n N_GCLK_c_1183_n 7.46878e-19 $X=7.92 $Y=1.41 $X2=0
+ $Y2=0
cc_571 N_A_1125_47#_c_865_n N_GCLK_c_1183_n 0.0283421f $X=6.825 $Y=1.79 $X2=0
+ $Y2=0
cc_572 N_A_1125_47#_M1014_g N_GCLK_c_1187_n 0.00959347f $X=7.425 $Y=0.56 $X2=0
+ $Y2=0
cc_573 N_A_1125_47#_M1022_g N_GCLK_c_1187_n 0.0024022f $X=7.895 $Y=0.56 $X2=0
+ $Y2=0
cc_574 N_A_1125_47#_c_842_n N_GCLK_c_1187_n 0.00160552f $X=8.02 $Y=1.16 $X2=0
+ $Y2=0
cc_575 N_A_1125_47#_c_855_n N_GCLK_c_1187_n 0.00346944f $X=6.91 $Y=1.185 $X2=0
+ $Y2=0
cc_576 N_A_1125_47#_M1004_g N_GCLK_c_1170_n 0.00148274f $X=6.955 $Y=0.56 $X2=0
+ $Y2=0
cc_577 N_A_1125_47#_M1014_g N_GCLK_c_1170_n 0.00257181f $X=7.425 $Y=0.56 $X2=0
+ $Y2=0
cc_578 N_A_1125_47#_c_842_n N_GCLK_c_1170_n 0.00297398f $X=8.02 $Y=1.16 $X2=0
+ $Y2=0
cc_579 N_A_1125_47#_c_858_n N_GCLK_c_1170_n 0.00501335f $X=6.74 $Y=0.7 $X2=0
+ $Y2=0
cc_580 N_A_1125_47#_c_845_n N_GCLK_c_1170_n 0.00645302f $X=6.825 $Y=1.055 $X2=0
+ $Y2=0
cc_581 N_A_1125_47#_c_855_n N_GCLK_c_1170_n 0.0171333f $X=6.91 $Y=1.185 $X2=0
+ $Y2=0
cc_582 N_A_1125_47#_c_849_n N_GCLK_c_1197_n 0.0148879f $X=7.45 $Y=1.41 $X2=0
+ $Y2=0
cc_583 N_A_1125_47#_c_842_n N_GCLK_c_1197_n 0.00240839f $X=8.02 $Y=1.16 $X2=0
+ $Y2=0
cc_584 N_A_1125_47#_c_855_n N_GCLK_c_1197_n 0.00346944f $X=6.91 $Y=1.185 $X2=0
+ $Y2=0
cc_585 N_A_1125_47#_c_848_n N_GCLK_c_1174_n 0.00143834f $X=6.98 $Y=1.41 $X2=0
+ $Y2=0
cc_586 N_A_1125_47#_c_849_n N_GCLK_c_1174_n 0.00186704f $X=7.45 $Y=1.41 $X2=0
+ $Y2=0
cc_587 N_A_1125_47#_c_842_n N_GCLK_c_1174_n 0.00150749f $X=8.02 $Y=1.16 $X2=0
+ $Y2=0
cc_588 N_A_1125_47#_c_854_n N_GCLK_c_1174_n 6.48059e-19 $X=6.825 $Y=1.495 $X2=0
+ $Y2=0
cc_589 N_A_1125_47#_c_855_n N_GCLK_c_1174_n 0.0185691f $X=6.91 $Y=1.185 $X2=0
+ $Y2=0
cc_590 N_A_1125_47#_c_865_n N_GCLK_c_1174_n 0.0113873f $X=6.825 $Y=1.79 $X2=0
+ $Y2=0
cc_591 N_A_1125_47#_M1014_g N_GCLK_c_1171_n 0.00300631f $X=7.425 $Y=0.56 $X2=0
+ $Y2=0
cc_592 N_A_1125_47#_M1022_g N_GCLK_c_1171_n 0.00162504f $X=7.895 $Y=0.56 $X2=0
+ $Y2=0
cc_593 N_A_1125_47#_c_842_n N_GCLK_c_1171_n 0.00393239f $X=8.02 $Y=1.16 $X2=0
+ $Y2=0
cc_594 N_A_1125_47#_c_849_n N_GCLK_c_1175_n 0.00166886f $X=7.45 $Y=1.41 $X2=0
+ $Y2=0
cc_595 N_A_1125_47#_c_850_n N_GCLK_c_1175_n 8.30867e-19 $X=7.92 $Y=1.41 $X2=0
+ $Y2=0
cc_596 N_A_1125_47#_c_842_n N_GCLK_c_1175_n 0.00320044f $X=8.02 $Y=1.16 $X2=0
+ $Y2=0
cc_597 N_A_1125_47#_M1004_g N_GCLK_c_1212_n 0.00306258f $X=6.955 $Y=0.56 $X2=0
+ $Y2=0
cc_598 N_A_1125_47#_M1014_g N_GCLK_c_1212_n 0.00254186f $X=7.425 $Y=0.56 $X2=0
+ $Y2=0
cc_599 N_A_1125_47#_c_855_n N_GCLK_c_1212_n 0.00261564f $X=6.91 $Y=1.185 $X2=0
+ $Y2=0
cc_600 N_A_1125_47#_c_842_n N_GCLK_c_1215_n 0.0117085f $X=8.02 $Y=1.16 $X2=0
+ $Y2=0
cc_601 N_A_1125_47#_c_855_n N_GCLK_c_1215_n 0.0178399f $X=6.91 $Y=1.185 $X2=0
+ $Y2=0
cc_602 N_A_1125_47#_c_841_n GCLK 0.0103356f $X=8.425 $Y=1.16 $X2=0 $Y2=0
cc_603 N_A_1125_47#_c_844_n GCLK 0.00447884f $X=8.525 $Y=1.217 $X2=0 $Y2=0
cc_604 N_A_1125_47#_c_850_n GCLK 0.0129232f $X=7.92 $Y=1.41 $X2=0 $Y2=0
cc_605 N_A_1125_47#_c_842_n GCLK 9.57476e-19 $X=8.02 $Y=1.16 $X2=0 $Y2=0
cc_606 N_A_1125_47#_c_852_n GCLK 0.0293036f $X=8.525 $Y=1.41 $X2=0 $Y2=0
cc_607 N_A_1125_47#_c_844_n GCLK 0.00665286f $X=8.525 $Y=1.217 $X2=0 $Y2=0
cc_608 N_A_1125_47#_c_844_n GCLK 0.00896406f $X=8.525 $Y=1.217 $X2=0 $Y2=0
cc_609 N_A_1125_47#_c_841_n N_GCLK_c_1178_n 0.0141146f $X=8.425 $Y=1.16 $X2=0
+ $Y2=0
cc_610 N_A_1125_47#_c_842_n N_GCLK_c_1178_n 0.0222994f $X=8.02 $Y=1.16 $X2=0
+ $Y2=0
cc_611 N_A_1125_47#_M1022_g N_GCLK_c_1173_n 0.00992861f $X=7.895 $Y=0.56 $X2=0
+ $Y2=0
cc_612 N_A_1125_47#_c_841_n N_GCLK_c_1173_n 0.00556565f $X=8.425 $Y=1.16 $X2=0
+ $Y2=0
cc_613 N_A_1125_47#_M1024_g N_GCLK_c_1173_n 0.0246222f $X=8.55 $Y=0.56 $X2=0
+ $Y2=0
cc_614 N_A_1125_47#_c_844_n N_GCLK_c_1173_n 0.00164051f $X=8.525 $Y=1.217 $X2=0
+ $Y2=0
cc_615 N_A_1125_47#_c_858_n N_VGND_M1021_d 0.00990816f $X=6.74 $Y=0.7 $X2=0
+ $Y2=0
cc_616 N_A_1125_47#_c_845_n N_VGND_M1021_d 0.00126753f $X=6.825 $Y=1.055 $X2=0
+ $Y2=0
cc_617 N_A_1125_47#_M1014_g N_VGND_c_1260_n 0.00400589f $X=7.425 $Y=0.56 $X2=0
+ $Y2=0
cc_618 N_A_1125_47#_M1022_g N_VGND_c_1260_n 0.0102164f $X=7.895 $Y=0.56 $X2=0
+ $Y2=0
cc_619 N_A_1125_47#_c_842_n N_VGND_c_1260_n 4.15508e-19 $X=8.02 $Y=1.16 $X2=0
+ $Y2=0
cc_620 N_A_1125_47#_M1024_g N_VGND_c_1260_n 7.75959e-19 $X=8.55 $Y=0.56 $X2=0
+ $Y2=0
cc_621 N_A_1125_47#_M1024_g N_VGND_c_1262_n 0.0171624f $X=8.55 $Y=0.56 $X2=0
+ $Y2=0
cc_622 N_A_1125_47#_M1004_g N_VGND_c_1265_n 0.00507199f $X=6.955 $Y=0.56 $X2=0
+ $Y2=0
cc_623 N_A_1125_47#_M1014_g N_VGND_c_1265_n 0.00420765f $X=7.425 $Y=0.56 $X2=0
+ $Y2=0
cc_624 N_A_1125_47#_c_858_n N_VGND_c_1265_n 0.00107125f $X=6.74 $Y=0.7 $X2=0
+ $Y2=0
cc_625 N_A_1125_47#_M1022_g N_VGND_c_1269_n 0.0046653f $X=7.895 $Y=0.56 $X2=0
+ $Y2=0
cc_626 N_A_1125_47#_M1024_g N_VGND_c_1269_n 0.00404729f $X=8.55 $Y=0.56 $X2=0
+ $Y2=0
cc_627 N_A_1125_47#_c_858_n N_VGND_c_1272_n 0.00255844f $X=6.74 $Y=0.7 $X2=0
+ $Y2=0
cc_628 N_A_1125_47#_c_846_n N_VGND_c_1272_n 0.0291387f $X=5.75 $Y=0.46 $X2=0
+ $Y2=0
cc_629 N_A_1125_47#_M1004_g N_VGND_c_1273_n 0.00465365f $X=6.955 $Y=0.56 $X2=0
+ $Y2=0
cc_630 N_A_1125_47#_c_858_n N_VGND_c_1273_n 0.0482871f $X=6.74 $Y=0.7 $X2=0
+ $Y2=0
cc_631 N_A_1125_47#_c_846_n N_VGND_c_1273_n 0.015853f $X=5.75 $Y=0.46 $X2=0
+ $Y2=0
cc_632 N_A_1125_47#_M1018_s N_VGND_c_1274_n 0.00286449f $X=5.625 $Y=0.235 $X2=0
+ $Y2=0
cc_633 N_A_1125_47#_M1004_g N_VGND_c_1274_n 0.00906214f $X=6.955 $Y=0.56 $X2=0
+ $Y2=0
cc_634 N_A_1125_47#_M1014_g N_VGND_c_1274_n 0.00607329f $X=7.425 $Y=0.56 $X2=0
+ $Y2=0
cc_635 N_A_1125_47#_M1022_g N_VGND_c_1274_n 0.00849071f $X=7.895 $Y=0.56 $X2=0
+ $Y2=0
cc_636 N_A_1125_47#_M1024_g N_VGND_c_1274_n 0.00800476f $X=8.55 $Y=0.56 $X2=0
+ $Y2=0
cc_637 N_A_1125_47#_c_858_n N_VGND_c_1274_n 0.0105743f $X=6.74 $Y=0.7 $X2=0
+ $Y2=0
cc_638 N_A_1125_47#_c_846_n N_VGND_c_1274_n 0.0159946f $X=5.75 $Y=0.46 $X2=0
+ $Y2=0
cc_639 N_A_1125_47#_c_858_n A_1217_47# 0.00202671f $X=6.74 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_640 N_VPWR_c_993_n A_117_369# 0.00184695f $X=8.97 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_641 N_VPWR_c_993_n N_A_27_47#_M1002_d 0.0041952f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_642 N_VPWR_c_995_n N_A_27_47#_c_1116_n 0.0214275f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_643 N_VPWR_c_995_n N_A_27_47#_c_1128_n 0.027538f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_644 N_VPWR_c_1006_n N_A_27_47#_c_1128_n 0.0132673f $X=2.575 $Y=2.44 $X2=0
+ $Y2=0
cc_645 N_VPWR_c_993_n N_A_27_47#_c_1128_n 0.00814261f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_646 N_VPWR_c_1006_n N_A_27_47#_c_1137_n 0.0369062f $X=2.575 $Y=2.44 $X2=0
+ $Y2=0
cc_647 N_VPWR_c_993_n N_A_27_47#_c_1137_n 0.0228157f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_648 N_VPWR_c_993_n A_421_413# 0.0077658f $X=8.97 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_649 N_VPWR_c_993_n N_GCLK_M1003_d 0.00444633f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_650 N_VPWR_c_993_n N_GCLK_M1020_d 0.0102279f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_651 N_VPWR_c_997_n N_GCLK_c_1183_n 0.039075f $X=7.685 $Y=2 $X2=0 $Y2=0
cc_652 N_VPWR_c_1000_n N_GCLK_c_1183_n 0.015413f $X=7.6 $Y=2.72 $X2=0 $Y2=0
cc_653 N_VPWR_c_993_n N_GCLK_c_1183_n 0.00946403f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_654 N_VPWR_M1017_s N_GCLK_c_1197_n 0.00301189f $X=7.54 $Y=1.485 $X2=0 $Y2=0
cc_655 N_VPWR_c_997_n N_GCLK_c_1197_n 0.01504f $X=7.685 $Y=2 $X2=0 $Y2=0
cc_656 N_VPWR_c_997_n GCLK 0.0280512f $X=7.685 $Y=2 $X2=0 $Y2=0
cc_657 N_VPWR_c_999_n GCLK 0.0758651f $X=8.85 $Y=1.66 $X2=0 $Y2=0
cc_658 N_VPWR_c_1005_n GCLK 0.0249582f $X=8.765 $Y=2.72 $X2=0 $Y2=0
cc_659 N_VPWR_c_993_n GCLK 0.0142154f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_660 N_VPWR_c_999_n GCLK 0.022905f $X=8.85 $Y=1.66 $X2=0 $Y2=0
cc_661 N_VPWR_c_997_n N_GCLK_c_1178_n 7.2207e-19 $X=7.685 $Y=2 $X2=0 $Y2=0
cc_662 A_117_369# N_A_27_47#_c_1116_n 0.00283574f $X=0.585 $Y=1.845 $X2=0 $Y2=0
cc_663 A_117_369# N_A_27_47#_c_1128_n 8.99713e-19 $X=0.585 $Y=1.845 $X2=0 $Y2=0
cc_664 A_117_369# N_A_27_47#_c_1137_n 0.00112381f $X=0.585 $Y=1.845 $X2=0 $Y2=0
cc_665 N_A_27_47#_c_1117_n N_VGND_M1016_d 0.00124282f $X=1.115 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_666 N_A_27_47#_c_1118_n N_VGND_M1016_d 8.45526e-19 $X=0.735 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_667 N_A_27_47#_c_1115_n N_VGND_c_1267_n 0.0173928f $X=0.26 $Y=0.43 $X2=0
+ $Y2=0
cc_668 N_A_27_47#_c_1118_n N_VGND_c_1267_n 0.00260613f $X=0.735 $Y=0.7 $X2=0
+ $Y2=0
cc_669 N_A_27_47#_c_1117_n N_VGND_c_1268_n 0.0032947f $X=1.115 $Y=0.7 $X2=0
+ $Y2=0
cc_670 N_A_27_47#_c_1141_n N_VGND_c_1268_n 0.0120906f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_671 N_A_27_47#_c_1115_n N_VGND_c_1270_n 0.0146378f $X=0.26 $Y=0.43 $X2=0
+ $Y2=0
cc_672 N_A_27_47#_c_1118_n N_VGND_c_1270_n 0.0211481f $X=0.735 $Y=0.7 $X2=0
+ $Y2=0
cc_673 N_A_27_47#_M1016_s N_VGND_c_1274_n 0.00286466f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_674 N_A_27_47#_M1001_d N_VGND_c_1274_n 0.00651855f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_675 N_A_27_47#_c_1115_n N_VGND_c_1274_n 0.00977915f $X=0.26 $Y=0.43 $X2=0
+ $Y2=0
cc_676 N_A_27_47#_c_1117_n N_VGND_c_1274_n 0.00548642f $X=1.115 $Y=0.7 $X2=0
+ $Y2=0
cc_677 N_A_27_47#_c_1118_n N_VGND_c_1274_n 0.00629427f $X=0.735 $Y=0.7 $X2=0
+ $Y2=0
cc_678 N_A_27_47#_c_1141_n N_VGND_c_1274_n 0.00681108f $X=1.2 $Y=0.42 $X2=0
+ $Y2=0
cc_679 N_GCLK_c_1187_n N_VGND_M1014_s 0.00447771f $X=7.65 $Y=0.8 $X2=0 $Y2=0
cc_680 N_GCLK_c_1179_n N_VGND_c_1260_n 0.00610556f $X=7.255 $Y=0.715 $X2=0 $Y2=0
cc_681 N_GCLK_c_1187_n N_VGND_c_1260_n 0.0135386f $X=7.65 $Y=0.8 $X2=0 $Y2=0
cc_682 N_GCLK_c_1212_n N_VGND_c_1260_n 0.011889f $X=7.215 $Y=0.36 $X2=0 $Y2=0
cc_683 N_GCLK_c_1178_n N_VGND_c_1260_n 8.87795e-19 $X=8.205 $Y=1.185 $X2=0 $Y2=0
cc_684 N_GCLK_c_1173_n N_VGND_c_1260_n 0.012712f $X=8.29 $Y=0.42 $X2=0 $Y2=0
cc_685 GCLK N_VGND_c_1262_n 0.022905f $X=8.885 $Y=1.105 $X2=0 $Y2=0
cc_686 N_GCLK_c_1173_n N_VGND_c_1262_n 0.0487704f $X=8.29 $Y=0.42 $X2=0 $Y2=0
cc_687 N_GCLK_c_1187_n N_VGND_c_1265_n 0.00271675f $X=7.65 $Y=0.8 $X2=0 $Y2=0
cc_688 N_GCLK_c_1212_n N_VGND_c_1265_n 0.020842f $X=7.215 $Y=0.36 $X2=0 $Y2=0
cc_689 N_GCLK_c_1173_n N_VGND_c_1269_n 0.0250111f $X=8.29 $Y=0.42 $X2=0 $Y2=0
cc_690 N_GCLK_M1004_d N_VGND_c_1274_n 0.00255381f $X=7.03 $Y=0.235 $X2=0 $Y2=0
cc_691 N_GCLK_M1022_d N_VGND_c_1274_n 0.0122643f $X=7.97 $Y=0.235 $X2=0 $Y2=0
cc_692 N_GCLK_c_1187_n N_VGND_c_1274_n 0.00619043f $X=7.65 $Y=0.8 $X2=0 $Y2=0
cc_693 N_GCLK_c_1212_n N_VGND_c_1274_n 0.0137736f $X=7.215 $Y=0.36 $X2=0 $Y2=0
cc_694 N_GCLK_c_1173_n N_VGND_c_1274_n 0.0143259f $X=8.29 $Y=0.42 $X2=0 $Y2=0
cc_695 N_VGND_c_1274_n A_425_47# 0.00367269f $X=8.97 $Y=0 $X2=-0.19 $Y2=-0.24
cc_696 N_VGND_c_1273_n A_1217_47# 0.00105937f $X=6.83 $Y=0.18 $X2=-0.19
+ $Y2=-0.24
