* File: sky130_fd_sc_hdll__buf_4.pxi.spice
* Created: Thu Aug 27 19:00:26 2020
* 
x_PM_SKY130_FD_SC_HDLL__BUF_4%A N_A_c_54_n N_A_M1002_g N_A_M1006_g A
+ PM_SKY130_FD_SC_HDLL__BUF_4%A
x_PM_SKY130_FD_SC_HDLL__BUF_4%A_27_47# N_A_27_47#_M1006_s N_A_27_47#_M1002_s
+ N_A_27_47#_c_94_n N_A_27_47#_M1000_g N_A_27_47#_M1001_g N_A_27_47#_c_95_n
+ N_A_27_47#_M1003_g N_A_27_47#_M1004_g N_A_27_47#_c_96_n N_A_27_47#_M1005_g
+ N_A_27_47#_M1007_g N_A_27_47#_c_97_n N_A_27_47#_M1008_g N_A_27_47#_M1009_g
+ N_A_27_47#_c_98_n N_A_27_47#_c_99_n N_A_27_47#_c_107_n N_A_27_47#_c_88_n
+ N_A_27_47#_c_89_n N_A_27_47#_c_113_n N_A_27_47#_c_90_n N_A_27_47#_c_91_n
+ N_A_27_47#_c_126_p N_A_27_47#_c_92_n N_A_27_47#_c_93_n
+ PM_SKY130_FD_SC_HDLL__BUF_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__BUF_4%VPWR N_VPWR_M1002_d N_VPWR_M1003_s N_VPWR_M1008_s
+ N_VPWR_c_196_n N_VPWR_c_197_n N_VPWR_c_198_n VPWR VPWR N_VPWR_c_199_n
+ N_VPWR_c_200_n N_VPWR_c_201_n N_VPWR_c_195_n N_VPWR_c_203_n N_VPWR_c_204_n
+ N_VPWR_c_205_n N_VPWR_c_206_n PM_SKY130_FD_SC_HDLL__BUF_4%VPWR
x_PM_SKY130_FD_SC_HDLL__BUF_4%X N_X_M1001_d N_X_M1007_d N_X_M1000_d N_X_M1005_d
+ N_X_c_254_n N_X_c_255_n N_X_c_247_n N_X_c_248_n N_X_c_250_n N_X_c_251_n
+ N_X_c_271_n X X X N_X_c_280_n PM_SKY130_FD_SC_HDLL__BUF_4%X
x_PM_SKY130_FD_SC_HDLL__BUF_4%VGND N_VGND_M1006_d N_VGND_M1004_s N_VGND_M1009_s
+ N_VGND_c_311_n N_VGND_c_312_n N_VGND_c_313_n VGND VGND N_VGND_c_314_n
+ N_VGND_c_315_n N_VGND_c_316_n N_VGND_c_317_n N_VGND_c_318_n N_VGND_c_319_n
+ N_VGND_c_320_n N_VGND_c_321_n PM_SKY130_FD_SC_HDLL__BUF_4%VGND
cc_1 VNB N_A_c_54_n 0.0373727f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_A_M1006_g 0.0232772f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_3 VNB A 0.0104808f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_A_27_47#_M1001_g 0.0187886f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.16
cc_5 VNB N_A_27_47#_M1004_g 0.0178228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_M1007_g 0.0178704f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_M1009_g 0.0236446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_88_n 0.00204016f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_89_n 0.00185886f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_90_n 0.00306916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_91_n 9.05057e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_92_n 0.00108293f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_93_n 0.105347f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_VPWR_c_195_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_X_c_247_n 0.00474317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_X_c_248_n 0.00137901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB X 0.00149571f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_311_n 0.00181111f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.16
cc_19 VNB N_VGND_c_312_n 0.00207171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_313_n 0.0321553f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_314_n 0.0155583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_315_n 0.0168868f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_316_n 0.0143186f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_317_n 0.0163041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_318_n 0.196828f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_319_n 0.00407139f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_320_n 0.00574292f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_321_n 0.00577057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_A_c_54_n 0.0380348f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_30 VPB A 0.0032877f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_31 VPB N_A_27_47#_c_94_n 0.0162447f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_A_27_47#_c_95_n 0.015418f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A_27_47#_c_96_n 0.0155598f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_27_47#_c_97_n 0.0198847f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_27_47#_c_98_n 0.00886215f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_27_47#_c_99_n 0.0316012f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_27_47#_c_91_n 0.00334531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_27_47#_c_93_n 0.0289015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_196_n 0.00234463f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.16
cc_40 VPB N_VPWR_c_197_n 3.21306e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_198_n 0.0461502f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_199_n 0.0144008f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_200_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_201_n 0.0163041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_195_n 0.0580909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_203_n 0.0194569f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_204_n 0.00346606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_205_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_206_n 0.00580385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_X_c_250_n 0.00276239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_X_c_251_n 0.00150118f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB X 0.00135553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB X 4.42593e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 N_A_c_54_n N_A_27_47#_c_94_n 0.021252f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_55 N_A_M1006_g N_A_27_47#_M1001_g 0.0194936f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_56 N_A_c_54_n N_A_27_47#_c_98_n 0.00240898f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_57 A N_A_27_47#_c_98_n 0.0252552f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_58 N_A_c_54_n N_A_27_47#_c_99_n 0.0108491f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_59 N_A_M1006_g N_A_27_47#_c_107_n 0.0059937f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_60 N_A_c_54_n N_A_27_47#_c_88_n 0.00254997f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_61 N_A_M1006_g N_A_27_47#_c_88_n 0.0136545f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_62 A N_A_27_47#_c_88_n 0.00903933f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_63 N_A_c_54_n N_A_27_47#_c_89_n 0.00413894f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_64 A N_A_27_47#_c_89_n 0.0139772f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_65 N_A_c_54_n N_A_27_47#_c_113_n 0.0148788f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_66 A N_A_27_47#_c_113_n 0.00309924f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_67 N_A_M1006_g N_A_27_47#_c_90_n 0.00392971f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_68 N_A_c_54_n N_A_27_47#_c_91_n 0.00441126f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_69 A N_A_27_47#_c_91_n 0.00430437f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_70 N_A_c_54_n N_A_27_47#_c_92_n 0.00154783f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_71 A N_A_27_47#_c_92_n 0.0116998f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_72 N_A_c_54_n N_A_27_47#_c_93_n 0.017092f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_73 N_A_c_54_n N_VPWR_c_196_n 0.00551021f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_74 N_A_c_54_n N_VPWR_c_195_n 0.0127805f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_75 N_A_c_54_n N_VPWR_c_203_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_76 N_A_M1006_g N_VGND_c_311_n 0.0118905f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_77 N_A_M1006_g N_VGND_c_314_n 0.0023344f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_78 N_A_M1006_g N_VGND_c_318_n 0.00406386f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_79 N_A_27_47#_c_113_n N_VPWR_M1002_d 0.00327879f $X=0.69 $Y=1.57 $X2=-0.19
+ $Y2=-0.24
cc_80 N_A_27_47#_c_94_n N_VPWR_c_196_n 0.0107285f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_27_47#_c_95_n N_VPWR_c_196_n 6.4992e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A_27_47#_c_99_n N_VPWR_c_196_n 0.0391438f $X=0.26 $Y=2.31 $X2=0 $Y2=0
cc_83 N_A_27_47#_c_113_n N_VPWR_c_196_n 0.0144498f $X=0.69 $Y=1.57 $X2=0 $Y2=0
cc_84 N_A_27_47#_c_126_p N_VPWR_c_196_n 3.99599e-19 $X=1.025 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_27_47#_c_94_n N_VPWR_c_197_n 7.03572e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A_27_47#_c_95_n N_VPWR_c_197_n 0.0154767f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_27_47#_c_96_n N_VPWR_c_197_n 0.0117392f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A_27_47#_c_97_n N_VPWR_c_197_n 6.61031e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A_27_47#_c_96_n N_VPWR_c_198_n 8.34825e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_27_47#_c_97_n N_VPWR_c_198_n 0.022204f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_91 N_A_27_47#_c_94_n N_VPWR_c_199_n 0.00661659f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_95_n N_VPWR_c_199_n 0.00427505f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_93 N_A_27_47#_c_96_n N_VPWR_c_200_n 0.00622633f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_27_47#_c_97_n N_VPWR_c_200_n 0.00427505f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A_27_47#_M1002_s N_VPWR_c_195_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_96 N_A_27_47#_c_94_n N_VPWR_c_195_n 0.0110933f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A_27_47#_c_95_n N_VPWR_c_195_n 0.00740765f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A_27_47#_c_96_n N_VPWR_c_195_n 0.010479f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A_27_47#_c_97_n N_VPWR_c_195_n 0.00740765f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A_27_47#_c_99_n N_VPWR_c_195_n 0.0124725f $X=0.26 $Y=2.31 $X2=0 $Y2=0
cc_101 N_A_27_47#_c_99_n N_VPWR_c_203_n 0.0210596f $X=0.26 $Y=2.31 $X2=0 $Y2=0
cc_102 N_A_27_47#_M1004_g N_X_c_254_n 0.00442074f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_103 N_A_27_47#_c_94_n N_X_c_255_n 0.0065097f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_27_47#_c_95_n N_X_c_255_n 0.00657309f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A_27_47#_M1004_g N_X_c_247_n 0.0127539f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_106 N_A_27_47#_M1007_g N_X_c_247_n 0.00649735f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_107 N_A_27_47#_c_93_n N_X_c_247_n 0.00404505f $X=2.375 $Y=1.217 $X2=0 $Y2=0
cc_108 N_A_27_47#_M1001_g N_X_c_248_n 8.24763e-19 $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_109 N_A_27_47#_c_88_n N_X_c_248_n 0.00133678f $X=0.69 $Y=0.82 $X2=0 $Y2=0
cc_110 N_A_27_47#_c_126_p N_X_c_248_n 0.0100467f $X=1.025 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A_27_47#_c_93_n N_X_c_248_n 0.0033396f $X=2.375 $Y=1.217 $X2=0 $Y2=0
cc_112 N_A_27_47#_c_95_n N_X_c_250_n 0.0163916f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_27_47#_c_96_n N_X_c_250_n 0.0103364f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_27_47#_c_93_n N_X_c_250_n 0.0102269f $X=2.375 $Y=1.217 $X2=0 $Y2=0
cc_115 N_A_27_47#_c_94_n N_X_c_251_n 0.00145092f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A_27_47#_c_91_n N_X_c_251_n 0.00251068f $X=0.775 $Y=1.485 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_126_p N_X_c_251_n 0.00893013f $X=1.025 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_27_47#_c_93_n N_X_c_251_n 0.00441044f $X=2.375 $Y=1.217 $X2=0 $Y2=0
cc_119 N_A_27_47#_M1009_g N_X_c_271_n 0.00168609f $X=2.4 $Y=0.56 $X2=0 $Y2=0
cc_120 N_A_27_47#_M1004_g X 6.34671e-19 $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_121 N_A_27_47#_c_96_n X 0.00105816f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A_27_47#_M1007_g X 0.00888778f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_123 N_A_27_47#_c_97_n X 9.12643e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A_27_47#_M1009_g X 0.00475854f $X=2.4 $Y=0.56 $X2=0 $Y2=0
cc_125 N_A_27_47#_c_93_n X 0.0478308f $X=2.375 $Y=1.217 $X2=0 $Y2=0
cc_126 N_A_27_47#_c_96_n X 0.00605739f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A_27_47#_c_97_n X 0.00210361f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A_27_47#_c_96_n N_X_c_280_n 0.00702928f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_27_47#_c_97_n N_X_c_280_n 0.00289399f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_27_47#_c_88_n N_VGND_M1006_d 0.00328906f $X=0.69 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_131 N_A_27_47#_M1001_g N_VGND_c_311_n 0.00300899f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_132 N_A_27_47#_c_107_n N_VGND_c_311_n 0.021682f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_133 N_A_27_47#_c_88_n N_VGND_c_311_n 0.0187264f $X=0.69 $Y=0.82 $X2=0 $Y2=0
cc_134 N_A_27_47#_M1001_g N_VGND_c_312_n 6.7227e-19 $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_135 N_A_27_47#_M1004_g N_VGND_c_312_n 0.0111872f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_136 N_A_27_47#_M1007_g N_VGND_c_312_n 0.00162962f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_137 N_A_27_47#_M1007_g N_VGND_c_313_n 8.031e-19 $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_138 N_A_27_47#_M1009_g N_VGND_c_313_n 0.0176565f $X=2.4 $Y=0.56 $X2=0 $Y2=0
cc_139 N_A_27_47#_c_107_n N_VGND_c_314_n 0.0117748f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_140 N_A_27_47#_c_88_n N_VGND_c_314_n 0.00206995f $X=0.69 $Y=0.82 $X2=0 $Y2=0
cc_141 N_A_27_47#_M1001_g N_VGND_c_315_n 0.00585385f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_142 N_A_27_47#_M1004_g N_VGND_c_315_n 0.0020416f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_143 N_A_27_47#_c_88_n N_VGND_c_315_n 6.84867e-19 $X=0.69 $Y=0.82 $X2=0 $Y2=0
cc_144 N_A_27_47#_M1007_g N_VGND_c_316_n 0.00439129f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_145 N_A_27_47#_M1009_g N_VGND_c_316_n 0.00271402f $X=2.4 $Y=0.56 $X2=0 $Y2=0
cc_146 N_A_27_47#_M1006_s N_VGND_c_318_n 0.00446555f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_147 N_A_27_47#_M1001_g N_VGND_c_318_n 0.011013f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_148 N_A_27_47#_M1004_g N_VGND_c_318_n 0.00288181f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_149 N_A_27_47#_M1007_g N_VGND_c_318_n 0.00613805f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_150 N_A_27_47#_M1009_g N_VGND_c_318_n 0.00510095f $X=2.4 $Y=0.56 $X2=0 $Y2=0
cc_151 N_A_27_47#_c_107_n N_VGND_c_318_n 0.0064623f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_152 N_A_27_47#_c_88_n N_VGND_c_318_n 0.00673892f $X=0.69 $Y=0.82 $X2=0 $Y2=0
cc_153 N_VPWR_c_195_n N_X_M1000_d 0.00656398f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_154 N_VPWR_c_195_n N_X_M1005_d 0.00656398f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_155 N_VPWR_c_196_n N_X_c_255_n 0.0359797f $X=0.73 $Y=2 $X2=0 $Y2=0
cc_156 N_VPWR_c_197_n N_X_c_255_n 0.0470327f $X=1.67 $Y=2 $X2=0 $Y2=0
cc_157 N_VPWR_c_199_n N_X_c_255_n 0.0118139f $X=1.455 $Y=2.72 $X2=0 $Y2=0
cc_158 N_VPWR_c_195_n N_X_c_255_n 0.00646998f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_159 N_VPWR_M1003_s N_X_c_250_n 0.00209407f $X=1.525 $Y=1.485 $X2=0 $Y2=0
cc_160 N_VPWR_c_197_n N_X_c_250_n 0.0172025f $X=1.67 $Y=2 $X2=0 $Y2=0
cc_161 N_VPWR_c_198_n X 0.0108422f $X=2.61 $Y=1.66 $X2=0 $Y2=0
cc_162 N_VPWR_c_197_n N_X_c_280_n 0.0385613f $X=1.67 $Y=2 $X2=0 $Y2=0
cc_163 N_VPWR_c_198_n N_X_c_280_n 0.0634205f $X=2.61 $Y=1.66 $X2=0 $Y2=0
cc_164 N_VPWR_c_200_n N_X_c_280_n 0.0118139f $X=2.395 $Y=2.72 $X2=0 $Y2=0
cc_165 N_VPWR_c_195_n N_X_c_280_n 0.00646998f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_166 N_VPWR_c_198_n N_VGND_c_313_n 0.0109366f $X=2.61 $Y=1.66 $X2=0 $Y2=0
cc_167 N_X_c_247_n N_VGND_M1004_s 0.00213931f $X=1.92 $Y=0.82 $X2=0 $Y2=0
cc_168 N_X_c_254_n N_VGND_c_312_n 0.0231432f $X=1.2 $Y=0.56 $X2=0 $Y2=0
cc_169 N_X_c_247_n N_VGND_c_312_n 0.0219272f $X=1.92 $Y=0.82 $X2=0 $Y2=0
cc_170 N_X_c_271_n N_VGND_c_313_n 0.0357983f $X=2.14 $Y=0.56 $X2=0 $Y2=0
cc_171 X N_VGND_c_313_n 0.0125104f $X=1.975 $Y=0.765 $X2=0 $Y2=0
cc_172 N_X_c_254_n N_VGND_c_315_n 0.0115672f $X=1.2 $Y=0.56 $X2=0 $Y2=0
cc_173 N_X_c_247_n N_VGND_c_315_n 0.00193889f $X=1.92 $Y=0.82 $X2=0 $Y2=0
cc_174 N_X_c_247_n N_VGND_c_316_n 9.89991e-19 $X=1.92 $Y=0.82 $X2=0 $Y2=0
cc_175 N_X_c_271_n N_VGND_c_316_n 0.0116048f $X=2.14 $Y=0.56 $X2=0 $Y2=0
cc_176 X N_VGND_c_316_n 0.00160042f $X=1.975 $Y=0.765 $X2=0 $Y2=0
cc_177 N_X_M1001_d N_VGND_c_318_n 0.00486275f $X=1.065 $Y=0.235 $X2=0 $Y2=0
cc_178 N_X_M1007_d N_VGND_c_318_n 0.00634176f $X=2.005 $Y=0.235 $X2=0 $Y2=0
cc_179 N_X_c_254_n N_VGND_c_318_n 0.0064623f $X=1.2 $Y=0.56 $X2=0 $Y2=0
cc_180 N_X_c_247_n N_VGND_c_318_n 0.00737166f $X=1.92 $Y=0.82 $X2=0 $Y2=0
cc_181 N_X_c_271_n N_VGND_c_318_n 0.00646998f $X=2.14 $Y=0.56 $X2=0 $Y2=0
cc_182 X N_VGND_c_318_n 0.0033156f $X=1.975 $Y=0.765 $X2=0 $Y2=0
