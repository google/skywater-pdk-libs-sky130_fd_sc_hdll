* File: sky130_fd_sc_hdll__a2bb2oi_1.spice
* Created: Thu Aug 27 18:55:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a2bb2oi_1.pex.spice"
.subckt sky130_fd_sc_hdll__a2bb2oi_1  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1007 N_A_119_47#_M1007_d N_A1_N_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.10725 AS=0.2015 PD=0.98 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_A2_N_M1003_g N_A_119_47#_M1007_d VNB NSHORT L=0.15
+ W=0.65 AD=0.26975 AS=0.10725 PD=1.48 PS=0.98 NRD=0 NRS=10.152 M=1 R=4.33333
+ SA=75000.7 SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_A_119_47#_M1004_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.13 AS=0.26975 PD=1.05 PS=1.48 NRD=0 NRS=39.684 M=1 R=4.33333 SA=75001.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1000 A_521_47# N_B2_M1000_g N_Y_M1004_d VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.13 PD=0.93 PS=1.05 NRD=15.684 NRS=23.076 M=1 R=4.33333 SA=75002.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_B1_M1008_g A_521_47# VNB NSHORT L=0.15 W=0.65 AD=0.2015
+ AS=0.091 PD=1.92 PS=0.93 NRD=8.304 NRS=15.684 M=1 R=4.33333 SA=75002.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 A_117_297# N_A1_N_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18 W=1 AD=0.115
+ AS=0.27 PD=1.23 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1001 N_A_119_47#_M1001_d N_A2_N_M1001_g A_117_297# VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.115 PD=2.54 PS=1.23 NRD=0.9653 NRS=11.8003 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1006 N_A_409_297#_M1006_d N_A_119_47#_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.18
+ W=1 AD=0.185 AS=0.27 PD=1.37 PS=2.54 NRD=16.7253 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_B2_M1009_g N_A_409_297#_M1006_d VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.185 PD=1.3 PS=1.37 NRD=2.9353 NRS=0.9653 M=1 R=5.55556 SA=90000.7
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1005 N_A_409_297#_M1005_d N_B1_M1005_g N_VPWR_M1009_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.15 PD=2.54 PS=1.3 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
pX11_noxref noxref_14 A2_N A2_N PROBETYPE=1
pX12_noxref noxref_15 Y Y PROBETYPE=1
pX13_noxref noxref_16 Y Y PROBETYPE=1
pX14_noxref noxref_17 Y Y PROBETYPE=1
*
.include "sky130_fd_sc_hdll__a2bb2oi_1.pxi.spice"
*
.ends
*
*
