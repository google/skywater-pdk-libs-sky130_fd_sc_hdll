* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 Q a_1972_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VPWR RESET_B a_1324_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X2 VPWR a_1972_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 a_1972_21# a_1757_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X4 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 a_618_389# D a_700_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=180000u
X6 VGND a_1202_413# a_1380_303# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X7 a_870_389# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=180000u
X8 a_1322_47# a_1380_303# a_1428_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND a_27_47# a_213_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Q a_1972_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_700_389# a_331_66# a_870_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=180000u
X12 a_700_389# SCE a_899_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=500000u
X13 a_1202_413# a_213_47# a_1322_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X14 a_1757_47# a_27_47# a_1866_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X15 VPWR SCE a_618_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=180000u
X16 a_631_119# D a_700_389# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_331_66# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=180000u
X18 a_331_66# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_1866_47# a_1972_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR a_1202_413# a_1380_303# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X21 a_1428_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_1324_413# a_1380_303# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X24 a_1380_303# a_213_47# a_1757_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X25 a_1202_413# a_27_47# a_1324_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X26 a_1380_303# a_27_47# a_1757_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X27 a_2157_47# a_1757_47# a_1972_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VGND a_1972_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_1757_47# a_213_47# a_1951_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X30 a_700_389# a_213_47# a_1202_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X31 VGND RESET_B a_2157_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 VGND a_331_66# a_631_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_1951_413# a_1972_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X34 VPWR a_27_47# a_213_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X35 a_899_66# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=180000u
X36 VPWR RESET_B a_1972_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X37 a_700_389# a_27_47# a_1202_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
.ends
