* File: sky130_fd_sc_hdll__o32ai_2.spice
* Created: Wed Sep  2 08:47:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o32ai_2.pex.spice"
.subckt sky130_fd_sc_hdll__o32ai_2  VNB VPB B2 B1 A3 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* A3	A3
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1003 N_A_27_47#_M1003_d N_B2_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75005.6 A=0.0975 P=1.6 MULT=1
MM1019 N_A_27_47#_M1019_d N_B2_M1019_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75005.1 A=0.0975 P=1.6 MULT=1
MM1005 N_Y_M1005_d N_B1_M1005_g N_A_27_47#_M1019_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75004.7 A=0.0975 P=1.6 MULT=1
MM1013 N_Y_M1005_d N_B1_M1013_g N_A_27_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75004.2 A=0.0975 P=1.6 MULT=1
MM1014 N_A_27_47#_M1013_s N_A3_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.3055 PD=0.92 PS=1.59 NRD=0 NRS=86.76 M=1 R=4.33333 SA=75002.1
+ SB=75003.8 A=0.0975 P=1.6 MULT=1
MM1016 N_A_27_47#_M1016_d N_A3_M1016_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.3055 PD=0.92 PS=1.59 NRD=0 NRS=35.076 M=1 R=4.33333 SA=75003.2
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_27_47#_M1016_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.6
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1000_d N_A2_M1008_g N_A_27_47#_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.25675 PD=1.02 PS=1.44 NRD=8.304 NRS=13.836 M=1 R=4.33333
+ SA=75004.1 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A1_M1004_g N_A_27_47#_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.25675 PD=0.97 PS=1.44 NRD=8.304 NRS=17.532 M=1 R=4.33333
+ SA=75005 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1004_d N_A1_M1017_g N_A_27_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.26 PD=0.97 PS=2.1 NRD=0 NRS=24.912 M=1 R=4.33333 SA=75005.5
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1001 N_A_27_297#_M1001_d N_B2_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1007 N_A_27_297#_M1007_d N_B2_M1007_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1012 N_A_27_297#_M1007_d N_B1_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1018 N_A_27_297#_M1018_d N_B1_M1018_g N_VPWR_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1002 N_Y_M1002_d N_A3_M1002_g N_A_525_297#_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=4.9053 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1015 N_Y_M1002_d N_A3_M1015_g N_A_525_297#_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1009 N_A_525_297#_M1015_s N_A2_M1009_g N_A_807_297#_M1009_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1011 N_A_525_297#_M1011_d N_A2_M1011_g N_A_807_297#_M1009_s VPB PHIGHVT L=0.18
+ W=1 AD=0.29 AS=0.145 PD=2.58 PS=1.29 NRD=4.9053 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g N_A_807_297#_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1010_d N_A1_M1010_g N_A_807_297#_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.29 AS=0.145 PD=2.58 PS=1.29 NRD=4.9053 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.9461 P=16.85
c_46 VNB 0 6.17784e-20 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hdll__o32ai_2.pxi.spice"
*
.ends
*
*
