* File: sky130_fd_sc_hdll__a22oi_2.pex.spice
* Created: Thu Aug 27 18:54:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A22OI_2%B2 1 3 4 6 7 9 10 12 13 14 22 30
c42 30 0 1.14332e-19 $X=0.695 $Y=1.19
c43 10 0 8.29508e-20 $X=0.99 $Y=0.995
r44 22 23 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r45 21 22 57.504 $w=3.73e-07 $l=4.45e-07 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.965 $Y2=1.202
r46 20 21 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r47 18 20 10.9839 $w=3.73e-07 $l=8.5e-08 $layer=POLY_cond $X=0.41 $Y=1.202
+ $X2=0.495 $Y2=1.202
r48 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r49 14 30 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=0.69 $Y=1.175
+ $X2=0.695 $Y2=1.175
r50 14 19 15.5273 $w=1.98e-07 $l=2.8e-07 $layer=LI1_cond $X=0.69 $Y=1.175
+ $X2=0.41 $Y2=1.175
r51 13 19 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.41 $Y2=1.175
r52 10 23 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r53 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r54 7 22 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r55 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r56 4 21 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r57 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r58 1 20 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r59 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_2%B1 1 3 4 6 7 9 10 12 13 14 22 25 31
c51 22 0 1.14332e-19 $X=1.905 $Y=1.202
r52 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=1.93 $Y2=1.202
r53 20 22 51.3711 $w=3.8e-07 $l=4.05e-07 $layer=POLY_cond $X=1.5 $Y=1.202
+ $X2=1.905 $Y2=1.202
r54 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.5
+ $Y=1.16 $X2=1.5 $Y2=1.16
r55 18 20 8.24474 $w=3.8e-07 $l=6.5e-08 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.5 $Y2=1.202
r56 17 18 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.202
+ $X2=1.435 $Y2=1.202
r57 14 31 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=1.605 $Y=1.175
+ $X2=1.615 $Y2=1.175
r58 14 21 5.82273 $w=1.98e-07 $l=1.05e-07 $layer=LI1_cond $X=1.605 $Y=1.175
+ $X2=1.5 $Y2=1.175
r59 13 21 18.3 $w=1.98e-07 $l=3.3e-07 $layer=LI1_cond $X=1.17 $Y=1.175 $X2=1.5
+ $Y2=1.175
r60 13 25 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=1.17 $Y=1.175
+ $X2=1.155 $Y2=1.175
r61 10 23 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r62 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r63 7 22 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r64 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r65 4 18 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r66 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r67 1 17 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.202
r68 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995 $X2=1.41
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_2%A1 1 3 4 6 7 9 10 12 13 14 22 28 31
r52 22 23 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=3.365 $Y=1.202
+ $X2=3.39 $Y2=1.202
r53 21 22 57.504 $w=3.73e-07 $l=4.45e-07 $layer=POLY_cond $X=2.92 $Y=1.202
+ $X2=3.365 $Y2=1.202
r54 20 21 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=2.895 $Y=1.202
+ $X2=2.92 $Y2=1.202
r55 18 20 10.9839 $w=3.73e-07 $l=8.5e-08 $layer=POLY_cond $X=2.81 $Y=1.202
+ $X2=2.895 $Y2=1.202
r56 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.81
+ $Y=1.16 $X2=2.81 $Y2=1.16
r57 14 31 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=3.405 $Y=1.175
+ $X2=3.415 $Y2=1.175
r58 14 28 21.6273 $w=1.98e-07 $l=3.9e-07 $layer=LI1_cond $X=3.405 $Y=1.175
+ $X2=3.015 $Y2=1.175
r59 13 28 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=3.01 $Y=1.175
+ $X2=3.015 $Y2=1.175
r60 13 19 11.0909 $w=1.98e-07 $l=2e-07 $layer=LI1_cond $X=3.01 $Y=1.175 $X2=2.81
+ $Y2=1.175
r61 10 23 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.39 $Y=0.995
+ $X2=3.39 $Y2=1.202
r62 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.39 $Y=0.995
+ $X2=3.39 $Y2=0.56
r63 7 22 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.202
r64 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.985
r65 4 21 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.92 $Y=0.995
+ $X2=2.92 $Y2=1.202
r66 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.92 $Y=0.995 $X2=2.92
+ $Y2=0.56
r67 1 20 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.202
r68 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_2%A2 1 3 4 6 7 9 10 12 13 14 22 25
r40 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.405 $Y=1.202
+ $X2=4.43 $Y2=1.202
r41 20 22 51.3711 $w=3.8e-07 $l=4.05e-07 $layer=POLY_cond $X=4 $Y=1.202
+ $X2=4.405 $Y2=1.202
r42 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4 $Y=1.16
+ $X2=4 $Y2=1.16
r43 18 20 8.24474 $w=3.8e-07 $l=6.5e-08 $layer=POLY_cond $X=3.935 $Y=1.202 $X2=4
+ $Y2=1.202
r44 17 18 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.91 $Y=1.202
+ $X2=3.935 $Y2=1.202
r45 14 21 21.35 $w=1.98e-07 $l=3.85e-07 $layer=LI1_cond $X=4.385 $Y=1.175 $X2=4
+ $Y2=1.175
r46 13 21 6.93182 $w=1.98e-07 $l=1.25e-07 $layer=LI1_cond $X=3.875 $Y=1.175
+ $X2=4 $Y2=1.175
r47 13 25 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=3.875 $Y=1.175
+ $X2=3.86 $Y2=1.175
r48 10 23 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.43 $Y=0.995
+ $X2=4.43 $Y2=1.202
r49 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.43 $Y=0.995
+ $X2=4.43 $Y2=0.56
r50 7 22 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.405 $Y=1.41
+ $X2=4.405 $Y2=1.202
r51 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.405 $Y=1.41
+ $X2=4.405 $Y2=1.985
r52 4 18 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.935 $Y=1.41
+ $X2=3.935 $Y2=1.202
r53 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.935 $Y=1.41
+ $X2=3.935 $Y2=1.985
r54 1 17 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.91 $Y=0.995
+ $X2=3.91 $Y2=1.202
r55 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.91 $Y=0.995 $X2=3.91
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_2%Y 1 2 3 4 5 18 20 21 24 26 28 34 36 37 38
+ 39 40 50 57
c88 50 0 1.72693e-19 $X=2.075 $Y=0.85
c89 28 0 8.29508e-20 $X=1.93 $Y=0.76
r90 55 57 0.132465 $w=4.33e-07 $l=5e-09 $layer=LI1_cond $X=2.142 $Y=1.655
+ $X2=2.142 $Y2=1.66
r91 47 50 0.134005 $w=4.28e-07 $l=5e-09 $layer=LI1_cond $X=2.145 $Y=0.845
+ $X2=2.145 $Y2=0.85
r92 40 57 5.56352 $w=4.33e-07 $l=2.1e-07 $layer=LI1_cond $X=2.142 $Y=1.87
+ $X2=2.142 $Y2=1.66
r93 39 48 2.24864 $w=4.32e-07 $l=8.6487e-08 $layer=LI1_cond $X=2.142 $Y=1.57
+ $X2=2.145 $Y2=1.485
r94 39 55 2.24864 $w=4.32e-07 $l=8.5e-08 $layer=LI1_cond $X=2.142 $Y=1.57
+ $X2=2.142 $Y2=1.655
r95 39 48 0.53602 $w=4.28e-07 $l=2e-08 $layer=LI1_cond $X=2.145 $Y=1.465
+ $X2=2.145 $Y2=1.485
r96 38 39 7.37028 $w=4.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.145 $Y=1.19
+ $X2=2.145 $Y2=1.465
r97 37 47 1.67165 $w=4.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=0.76
+ $X2=2.145 $Y2=0.845
r98 37 38 8.0403 $w=4.28e-07 $l=3e-07 $layer=LI1_cond $X=2.145 $Y=0.89 $X2=2.145
+ $Y2=1.19
r99 37 50 1.07204 $w=4.28e-07 $l=4e-08 $layer=LI1_cond $X=2.145 $Y=0.89
+ $X2=2.145 $Y2=0.85
r100 32 37 10.2816 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.36 $Y=0.76
+ $X2=2.145 $Y2=0.76
r101 32 34 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.36 $Y=0.76
+ $X2=3.13 $Y2=0.76
r102 28 37 10.2816 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=1.93 $Y=0.76
+ $X2=2.145 $Y2=0.76
r103 28 30 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.93 $Y=0.76
+ $X2=1.67 $Y2=0.76
r104 27 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.365 $Y=1.57
+ $X2=1.175 $Y2=1.57
r105 26 39 4.84258 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=1.925 $Y=1.57
+ $X2=2.142 $Y2=1.57
r106 26 27 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.925 $Y=1.57
+ $X2=1.365 $Y2=1.57
r107 22 36 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=1.655
+ $X2=1.175 $Y2=1.57
r108 22 24 0.151637 $w=3.78e-07 $l=5e-09 $layer=LI1_cond $X=1.175 $Y=1.655
+ $X2=1.175 $Y2=1.66
r109 20 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.985 $Y=1.57
+ $X2=1.175 $Y2=1.57
r110 20 21 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.985 $Y=1.57
+ $X2=0.345 $Y2=1.57
r111 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.22 $Y=1.655
+ $X2=0.345 $Y2=1.57
r112 16 18 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=0.22 $Y=1.655
+ $X2=0.22 $Y2=1.8
r113 5 57 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.66
r114 4 24 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.66
r115 3 18 300 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.8
r116 2 34 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=2.995
+ $Y=0.235 $X2=3.13 $Y2=0.76
r117 1 30 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_2%A_117_297# 1 2 3 4 5 18 20 21 24 26 29 31
+ 32 33 36 40 44 48 51
r84 44 46 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=4.615 $Y=1.66
+ $X2=4.615 $Y2=2.34
r85 42 44 0.151637 $w=3.78e-07 $l=5e-09 $layer=LI1_cond $X=4.615 $Y=1.655
+ $X2=4.615 $Y2=1.66
r86 41 51 11.015 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=3.865 $Y=1.57
+ $X2=3.625 $Y2=1.57
r87 40 42 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=4.425 $Y=1.57
+ $X2=4.615 $Y2=1.655
r88 40 41 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.425 $Y=1.57
+ $X2=3.865 $Y2=1.57
r89 36 38 16.9444 $w=4.78e-07 $l=6.8e-07 $layer=LI1_cond $X=3.625 $Y=1.66
+ $X2=3.625 $Y2=2.34
r90 34 51 1.96841 $w=4.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=1.655
+ $X2=3.625 $Y2=1.57
r91 34 36 0.124591 $w=4.78e-07 $l=5e-09 $layer=LI1_cond $X=3.625 $Y=1.655
+ $X2=3.625 $Y2=1.66
r92 32 51 11.015 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=3.385 $Y=1.57
+ $X2=3.625 $Y2=1.57
r93 32 33 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.385 $Y=1.57
+ $X2=2.825 $Y2=1.57
r94 29 50 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.7 $Y=2.295 $X2=2.7
+ $Y2=2.38
r95 29 31 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=2.7 $Y=2.295
+ $X2=2.7 $Y2=1.66
r96 28 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.7 $Y=1.655
+ $X2=2.825 $Y2=1.57
r97 28 31 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=2.7 $Y=1.655 $X2=2.7
+ $Y2=1.66
r98 27 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=2.38
+ $X2=1.67 $Y2=2.38
r99 26 50 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.575 $Y=2.38
+ $X2=2.7 $Y2=2.38
r100 26 27 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=2.575 $Y=2.38
+ $X2=1.755 $Y2=2.38
r101 22 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=2.295
+ $X2=1.67 $Y2=2.38
r102 22 24 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.67 $Y=2.295
+ $X2=1.67 $Y2=2
r103 20 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=2.38
+ $X2=1.67 $Y2=2.38
r104 20 21 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.585 $Y=2.38
+ $X2=0.815 $Y2=2.38
r105 16 21 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=0.665 $Y=2.295
+ $X2=0.815 $Y2=2.38
r106 16 18 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.665 $Y=2.295
+ $X2=0.665 $Y2=2
r107 5 46 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.495
+ $Y=1.485 $X2=4.64 $Y2=2.34
r108 5 44 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.495
+ $Y=1.485 $X2=4.64 $Y2=1.66
r109 4 38 400 $w=1.7e-07 $l=9.69794e-07 $layer=licon1_PDIFF $count=1 $X=3.455
+ $Y=1.485 $X2=3.7 $Y2=2.34
r110 4 36 400 $w=1.7e-07 $l=3.2078e-07 $layer=licon1_PDIFF $count=1 $X=3.455
+ $Y=1.485 $X2=3.7 $Y2=1.66
r111 3 50 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.535
+ $Y=1.485 $X2=2.66 $Y2=2.34
r112 3 31 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=2.535
+ $Y=1.485 $X2=2.66 $Y2=1.66
r113 2 24 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2
r114 1 18 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_2%VPWR 1 2 9 13 16 17 19 20 21 23 30 39 40
r62 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r63 37 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r64 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r65 34 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r66 33 34 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r67 26 30 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.695 $Y2=2.72
r68 23 34 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.99 $Y2=2.72
r69 23 26 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r70 21 33 146.465 $w=1.68e-07 $l=2.245e-06 $layer=LI1_cond $X=0.745 $Y=2.72
+ $X2=2.99 $Y2=2.72
r71 21 30 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=0.745 $Y=2.72
+ $X2=0.695 $Y2=2.72
r72 19 36 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.085 $Y=2.72
+ $X2=3.91 $Y2=2.72
r73 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.085 $Y=2.72
+ $X2=4.17 $Y2=2.72
r74 18 39 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=4.255 $Y=2.72
+ $X2=4.83 $Y2=2.72
r75 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.255 $Y=2.72
+ $X2=4.17 $Y2=2.72
r76 16 33 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.045 $Y=2.72
+ $X2=2.99 $Y2=2.72
r77 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.045 $Y=2.72
+ $X2=3.13 $Y2=2.72
r78 15 36 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=3.91 $Y2=2.72
r79 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=3.13 $Y2=2.72
r80 11 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.17 $Y=2.635
+ $X2=4.17 $Y2=2.72
r81 11 13 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.17 $Y=2.635
+ $X2=4.17 $Y2=2
r82 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=2.635 $X2=3.13
+ $Y2=2.72
r83 7 9 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.13 $Y=2.635
+ $X2=3.13 $Y2=2
r84 2 13 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.025
+ $Y=1.485 $X2=4.17 $Y2=2
r85 1 9 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.985
+ $Y=1.485 $X2=3.13 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_2%A_27_47# 1 2 3 10 13 14 19 21
c37 3 0 1.72693e-19 $X=2.005 $Y=0.235
r38 19 21 39.4136 $w=2.48e-07 $l=8.55e-07 $layer=LI1_cond $X=1.285 $Y=0.38
+ $X2=2.14 $Y2=0.38
r39 16 18 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.2 $Y=0.68 $X2=1.2
+ $Y2=0.57
r40 15 19 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.2 $Y=0.505
+ $X2=1.285 $Y2=0.38
r41 15 18 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=1.2 $Y=0.505 $X2=1.2
+ $Y2=0.57
r42 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.115 $Y=0.765
+ $X2=1.2 $Y2=0.68
r43 13 14 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=0.765
+ $X2=0.345 $Y2=0.765
r44 10 14 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.22 $Y=0.68
+ $X2=0.345 $Y2=0.765
r45 10 12 5.368 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=0.22 $Y=0.68 $X2=0.22
+ $Y2=0.57
r46 3 21 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.42
r47 2 18 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.57
r48 1 12 182 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_2%VGND 1 2 9 12 13 14 17 19 32 33 41
r62 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r63 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r64 29 30 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r65 27 30 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=3.91
+ $Y2=0
r66 27 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r67 26 29 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=3.91
+ $Y2=0
r68 26 27 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r69 24 26 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.15
+ $Y2=0
r70 19 21 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r71 17 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r72 17 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r73 14 41 8.0037 $w=5.48e-07 $l=3.15e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.4
r74 14 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r75 14 19 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.705 $Y=0 $X2=0.515
+ $Y2=0
r76 14 24 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.705 $Y=0 $X2=0.895
+ $Y2=0
r77 12 29 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.98 $Y=0 $X2=3.91
+ $Y2=0
r78 12 13 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.98 $Y=0 $X2=4.17
+ $Y2=0
r79 11 32 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=4.36 $Y=0 $X2=4.83
+ $Y2=0
r80 11 13 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.36 $Y=0 $X2=4.17
+ $Y2=0
r81 7 13 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.17 $Y=0.085 $X2=4.17
+ $Y2=0
r82 7 9 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=4.17 $Y=0.085
+ $X2=4.17 $Y2=0.4
r83 2 9 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.985
+ $Y=0.235 $X2=4.17 $Y2=0.4
r84 1 41 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_2%A_507_47# 1 2 3 10 17 18 19 20
r31 20 22 4.19375 $w=3.2e-07 $l=1.1e-07 $layer=LI1_cond $X=4.715 $Y=0.68
+ $X2=4.715 $Y2=0.57
r32 18 20 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=4.555 $Y=0.765
+ $X2=4.715 $Y2=0.68
r33 18 19 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.555 $Y=0.765
+ $X2=3.785 $Y2=0.765
r34 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.7 $Y=0.68
+ $X2=3.785 $Y2=0.765
r35 15 17 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.7 $Y=0.68 $X2=3.7
+ $Y2=0.57
r36 14 17 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.7 $Y=0.505 $X2=3.7
+ $Y2=0.57
r37 10 14 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.615 $Y=0.38
+ $X2=3.7 $Y2=0.505
r38 10 12 44.0233 $w=2.48e-07 $l=9.55e-07 $layer=LI1_cond $X=3.615 $Y=0.38
+ $X2=2.66 $Y2=0.38
r39 3 22 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=4.505
+ $Y=0.235 $X2=4.64 $Y2=0.57
r40 2 17 182 $w=1.7e-07 $l=4.36978e-07 $layer=licon1_NDIFF $count=1 $X=3.465
+ $Y=0.235 $X2=3.7 $Y2=0.57
r41 1 12 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.235 $X2=2.66 $Y2=0.42
.ends

