* NGSPICE file created from sky130_fd_sc_hdll__clkbuf_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__clkbuf_4 A VGND VNB VPB VPWR X
M1000 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=4.011e+11p pd=4.43e+06u as=1.323e+11p ps=1.47e+06u
M1001 X a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=2.982e+11p pd=3.1e+06u as=0p ps=0u
M1002 X a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=9.6e+11p pd=7.92e+06u as=2.75e+11p ps=2.55e+06u
M1004 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=6e+11p ps=5.2e+06u
M1005 VGND a_27_47# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_27_47# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

