* File: sky130_fd_sc_hdll__xnor3_2.pxi.spice
* Created: Thu Aug 27 19:29:30 2020
* 
x_PM_SKY130_FD_SC_HDLL__XNOR3_2%A_79_21# N_A_79_21#_M1007_d N_A_79_21#_M1016_d
+ N_A_79_21#_c_158_n N_A_79_21#_M1002_g N_A_79_21#_c_165_n N_A_79_21#_M1013_g
+ N_A_79_21#_c_166_n N_A_79_21#_M1019_g N_A_79_21#_c_159_n N_A_79_21#_M1023_g
+ N_A_79_21#_c_160_n N_A_79_21#_c_174_p N_A_79_21#_c_246_p N_A_79_21#_c_179_p
+ N_A_79_21#_c_208_p N_A_79_21#_c_161_n N_A_79_21#_c_168_n N_A_79_21#_c_162_n
+ N_A_79_21#_c_169_n N_A_79_21#_c_170_n N_A_79_21#_c_183_p N_A_79_21#_c_193_p
+ N_A_79_21#_c_163_n N_A_79_21#_c_164_n PM_SKY130_FD_SC_HDLL__XNOR3_2%A_79_21#
x_PM_SKY130_FD_SC_HDLL__XNOR3_2%C N_C_c_266_n N_C_M1009_g N_C_M1003_g
+ N_C_c_267_n N_C_M1016_g N_C_c_268_n N_C_M1007_g N_C_c_269_n N_C_c_270_n C
+ PM_SKY130_FD_SC_HDLL__XNOR3_2%C
x_PM_SKY130_FD_SC_HDLL__XNOR3_2%A_328_93# N_A_328_93#_M1009_d
+ N_A_328_93#_M1003_d N_A_328_93#_c_326_n N_A_328_93#_M1000_g
+ N_A_328_93#_c_327_n N_A_328_93#_M1008_g N_A_328_93#_c_342_n
+ N_A_328_93#_c_328_n N_A_328_93#_c_332_n N_A_328_93#_c_333_n
+ N_A_328_93#_c_334_n N_A_328_93#_c_329_n
+ PM_SKY130_FD_SC_HDLL__XNOR3_2%A_328_93#
x_PM_SKY130_FD_SC_HDLL__XNOR3_2%A_885_297# N_A_885_297#_M1022_d
+ N_A_885_297#_M1005_d N_A_885_297#_c_412_n N_A_885_297#_M1017_g
+ N_A_885_297#_M1001_g N_A_885_297#_c_399_n N_A_885_297#_c_414_n
+ N_A_885_297#_M1014_g N_A_885_297#_M1012_g N_A_885_297#_c_400_n
+ N_A_885_297#_c_401_n N_A_885_297#_c_417_n N_A_885_297#_c_402_n
+ N_A_885_297#_c_403_n N_A_885_297#_c_421_p N_A_885_297#_c_404_n
+ N_A_885_297#_c_405_n N_A_885_297#_c_406_n N_A_885_297#_c_407_n
+ N_A_885_297#_c_408_n N_A_885_297#_c_409_n N_A_885_297#_c_410_n
+ N_A_885_297#_c_411_n PM_SKY130_FD_SC_HDLL__XNOR3_2%A_885_297#
x_PM_SKY130_FD_SC_HDLL__XNOR3_2%B N_B_c_589_n N_B_M1005_g N_B_M1022_g
+ N_B_c_582_n N_B_c_583_n N_B_M1010_g N_B_M1015_g N_B_c_592_n N_B_c_593_n
+ N_B_M1004_g N_B_c_594_n N_B_c_595_n N_B_M1006_g N_B_c_585_n N_B_c_586_n
+ N_B_c_587_n N_B_c_600_n B N_B_c_588_n B PM_SKY130_FD_SC_HDLL__XNOR3_2%B
x_PM_SKY130_FD_SC_HDLL__XNOR3_2%A N_A_c_717_n N_A_M1018_g N_A_c_718_n
+ N_A_M1021_g A PM_SKY130_FD_SC_HDLL__XNOR3_2%A
x_PM_SKY130_FD_SC_HDLL__XNOR3_2%A_1003_297# N_A_1003_297#_M1015_s
+ N_A_1003_297#_M1012_d N_A_1003_297#_M1010_s N_A_1003_297#_M1014_d
+ N_A_1003_297#_c_752_n N_A_1003_297#_M1020_g N_A_1003_297#_c_753_n
+ N_A_1003_297#_M1011_g N_A_1003_297#_c_754_n N_A_1003_297#_c_762_n
+ N_A_1003_297#_c_755_n N_A_1003_297#_c_756_n N_A_1003_297#_c_757_n
+ N_A_1003_297#_c_764_n N_A_1003_297#_c_774_n N_A_1003_297#_c_758_n
+ N_A_1003_297#_c_759_n N_A_1003_297#_c_787_n N_A_1003_297#_c_788_n
+ PM_SKY130_FD_SC_HDLL__XNOR3_2%A_1003_297#
x_PM_SKY130_FD_SC_HDLL__XNOR3_2%VPWR N_VPWR_M1013_s N_VPWR_M1019_s
+ N_VPWR_M1005_s N_VPWR_M1018_d N_VPWR_c_885_n N_VPWR_c_886_n N_VPWR_c_887_n
+ N_VPWR_c_888_n N_VPWR_c_889_n N_VPWR_c_890_n N_VPWR_c_891_n VPWR
+ N_VPWR_c_892_n N_VPWR_c_893_n N_VPWR_c_894_n N_VPWR_c_884_n N_VPWR_c_896_n
+ N_VPWR_c_897_n PM_SKY130_FD_SC_HDLL__XNOR3_2%VPWR
x_PM_SKY130_FD_SC_HDLL__XNOR3_2%X N_X_M1002_s N_X_M1013_d X N_X_c_981_n
+ PM_SKY130_FD_SC_HDLL__XNOR3_2%X
x_PM_SKY130_FD_SC_HDLL__XNOR3_2%A_453_325# N_A_453_325#_M1008_d
+ N_A_453_325#_M1015_d N_A_453_325#_M1016_s N_A_453_325#_M1006_d
+ N_A_453_325#_c_1001_n N_A_453_325#_c_995_n N_A_453_325#_c_996_n
+ N_A_453_325#_c_997_n N_A_453_325#_c_1003_n N_A_453_325#_c_1004_n
+ N_A_453_325#_c_1005_n N_A_453_325#_c_1006_n N_A_453_325#_c_998_n
+ N_A_453_325#_c_1008_n N_A_453_325#_c_1046_n N_A_453_325#_c_999_n
+ N_A_453_325#_c_1009_n N_A_453_325#_c_1000_n N_A_453_325#_c_1010_n
+ PM_SKY130_FD_SC_HDLL__XNOR3_2%A_453_325#
x_PM_SKY130_FD_SC_HDLL__XNOR3_2%A_477_49# N_A_477_49#_M1007_s
+ N_A_477_49#_M1004_d N_A_477_49#_M1000_d N_A_477_49#_M1010_d
+ N_A_477_49#_c_1162_n N_A_477_49#_c_1150_n N_A_477_49#_c_1154_n
+ N_A_477_49#_c_1191_n N_A_477_49#_c_1155_n N_A_477_49#_c_1151_n
+ N_A_477_49#_c_1270_p N_A_477_49#_c_1204_n N_A_477_49#_c_1205_n
+ N_A_477_49#_c_1152_n N_A_477_49#_c_1226_n N_A_477_49#_c_1157_n
+ N_A_477_49#_c_1158_n N_A_477_49#_c_1159_n N_A_477_49#_c_1160_n
+ PM_SKY130_FD_SC_HDLL__XNOR3_2%A_477_49#
x_PM_SKY130_FD_SC_HDLL__XNOR3_2%A_1286_297# N_A_1286_297#_M1001_d
+ N_A_1286_297#_M1020_d N_A_1286_297#_M1017_d N_A_1286_297#_M1011_d
+ N_A_1286_297#_c_1286_n N_A_1286_297#_c_1298_n N_A_1286_297#_c_1290_n
+ N_A_1286_297#_c_1287_n N_A_1286_297#_c_1299_n N_A_1286_297#_c_1292_n
+ N_A_1286_297#_c_1288_n PM_SKY130_FD_SC_HDLL__XNOR3_2%A_1286_297#
x_PM_SKY130_FD_SC_HDLL__XNOR3_2%VGND N_VGND_M1002_d N_VGND_M1023_d
+ N_VGND_M1022_s N_VGND_M1021_d N_VGND_c_1353_n N_VGND_c_1354_n N_VGND_c_1355_n
+ N_VGND_c_1356_n N_VGND_c_1357_n N_VGND_c_1358_n N_VGND_c_1359_n
+ N_VGND_c_1360_n N_VGND_c_1361_n VGND N_VGND_c_1362_n N_VGND_c_1363_n
+ N_VGND_c_1364_n N_VGND_c_1365_n PM_SKY130_FD_SC_HDLL__XNOR3_2%VGND
cc_1 VNB N_A_79_21#_c_158_n 0.0228255f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_159_n 0.0187967f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB N_A_79_21#_c_160_n 0.00109568f $X=-0.19 $Y=-0.24 $X2=1.145 $Y2=1.16
cc_4 VNB N_A_79_21#_c_161_n 0.00138296f $X=-0.19 $Y=-0.24 $X2=1.605 $Y2=0.695
cc_5 VNB N_A_79_21#_c_162_n 0.00216404f $X=-0.19 $Y=-0.24 $X2=1.715 $Y2=0.34
cc_6 VNB N_A_79_21#_c_163_n 0.0163054f $X=-0.19 $Y=-0.24 $X2=2.68 $Y2=0.355
cc_7 VNB N_A_79_21#_c_164_n 0.0630256f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.202
cc_8 VNB N_C_c_266_n 0.0199295f $X=-0.19 $Y=-0.24 $X2=2.855 $Y2=0.245
cc_9 VNB N_C_c_267_n 0.0145755f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_10 VNB N_C_c_268_n 0.0213243f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_11 VNB N_C_c_269_n 0.0118432f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.985
cc_12 VNB N_C_c_270_n 0.0544628f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_13 VNB N_A_328_93#_c_326_n 0.0251626f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_14 VNB N_A_328_93#_c_327_n 0.0205014f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_15 VNB N_A_328_93#_c_328_n 0.0026062f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_16 VNB N_A_328_93#_c_329_n 0.00273938f $X=-0.19 $Y=-0.24 $X2=1.605 $Y2=0.425
cc_17 VNB N_A_885_297#_M1001_g 0.0360077f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_18 VNB N_A_885_297#_c_399_n 0.00170012f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.985
cc_19 VNB N_A_885_297#_c_400_n 0.0288368f $X=-0.19 $Y=-0.24 $X2=1.145 $Y2=1.16
cc_20 VNB N_A_885_297#_c_401_n 0.0176837f $X=-0.19 $Y=-0.24 $X2=1.145 $Y2=1.16
cc_21 VNB N_A_885_297#_c_402_n 0.00239744f $X=-0.19 $Y=-0.24 $X2=2.925 $Y2=2.32
cc_22 VNB N_A_885_297#_c_403_n 0.00792514f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_885_297#_c_404_n 0.0128101f $X=-0.19 $Y=-0.24 $X2=3 $Y2=0.355
cc_24 VNB N_A_885_297#_c_405_n 0.00136794f $X=-0.19 $Y=-0.24 $X2=3 $Y2=0.37
cc_25 VNB N_A_885_297#_c_406_n 0.00305152f $X=-0.19 $Y=-0.24 $X2=1.145 $Y2=1.202
cc_26 VNB N_A_885_297#_c_407_n 0.00216737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_885_297#_c_408_n 0.00613074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_885_297#_c_409_n 0.0286378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_885_297#_c_410_n 0.0195573f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_885_297#_c_411_n 0.00256224f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_B_M1022_g 0.0302339f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_B_c_582_n 0.0558482f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_33 VNB N_B_c_583_n 0.0317672f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_34 VNB N_B_M1015_g 0.0287454f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_35 VNB N_B_c_585_n 0.010365f $X=-0.19 $Y=-0.24 $X2=1.72 $Y2=2.235
cc_36 VNB N_B_c_586_n 0.00131136f $X=-0.19 $Y=-0.24 $X2=2.925 $Y2=2.32
cc_37 VNB N_B_c_587_n 0.0298595f $X=-0.19 $Y=-0.24 $X2=2.925 $Y2=2.32
cc_38 VNB N_B_c_588_n 0.0212173f $X=-0.19 $Y=-0.24 $X2=2.68 $Y2=0.355
cc_39 VNB N_A_c_717_n 0.0239526f $X=-0.19 $Y=-0.24 $X2=2.855 $Y2=0.245
cc_40 VNB N_A_c_718_n 0.017807f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB A 0.00586957f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_42 VNB N_A_1003_297#_c_752_n 0.0206212f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.41
cc_43 VNB N_A_1003_297#_c_753_n 0.0371145f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_44 VNB N_A_1003_297#_c_754_n 0.00634916f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.16
cc_45 VNB N_A_1003_297#_c_755_n 0.00288102f $X=-0.19 $Y=-0.24 $X2=1.265 $Y2=1.96
cc_46 VNB N_A_1003_297#_c_756_n 0.00201667f $X=-0.19 $Y=-0.24 $X2=1.605
+ $Y2=0.425
cc_47 VNB N_A_1003_297#_c_757_n 0.00544021f $X=-0.19 $Y=-0.24 $X2=1.605
+ $Y2=0.695
cc_48 VNB N_A_1003_297#_c_758_n 0.00212326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_1003_297#_c_759_n 0.00497895f $X=-0.19 $Y=-0.24 $X2=3 $Y2=0.37
cc_50 VNB N_VPWR_c_884_n 0.402575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_X_c_981_n 0.00171053f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_52 VNB N_A_453_325#_c_995_n 0.0107596f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_53 VNB N_A_453_325#_c_996_n 0.0139216f $X=-0.19 $Y=-0.24 $X2=1.145 $Y2=1.16
cc_54 VNB N_A_453_325#_c_997_n 0.00281469f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=0.78
cc_55 VNB N_A_453_325#_c_998_n 0.00223628f $X=-0.19 $Y=-0.24 $X2=2.68 $Y2=0.34
cc_56 VNB N_A_453_325#_c_999_n 0.0104576f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.202
cc_57 VNB N_A_453_325#_c_1000_n 2.7378e-19 $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.202
cc_58 VNB N_A_477_49#_c_1150_n 0.00895087f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_59 VNB N_A_477_49#_c_1151_n 0.0097913f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=0.78
cc_60 VNB N_A_477_49#_c_1152_n 0.00621279f $X=-0.19 $Y=-0.24 $X2=1.83 $Y2=2.32
cc_61 VNB N_A_1286_297#_c_1286_n 0.00788488f $X=-0.19 $Y=-0.24 $X2=0.985
+ $Y2=1.985
cc_62 VNB N_A_1286_297#_c_1287_n 0.0309074f $X=-0.19 $Y=-0.24 $X2=1.61 $Y2=1.96
cc_63 VNB N_A_1286_297#_c_1288_n 0.0135316f $X=-0.19 $Y=-0.24 $X2=2.925 $Y2=2.32
cc_64 VNB N_VGND_c_1353_n 0.0104904f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.41
cc_65 VNB N_VGND_c_1354_n 0.0259911f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.985
cc_66 VNB N_VGND_c_1355_n 0.00249996f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=0.865
cc_67 VNB N_VGND_c_1356_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=1.145 $Y2=1.16
cc_68 VNB N_VGND_c_1357_n 0.00471543f $X=-0.19 $Y=-0.24 $X2=1.265 $Y2=1.96
cc_69 VNB N_VGND_c_1358_n 0.0677757f $X=-0.19 $Y=-0.24 $X2=1.72 $Y2=2.045
cc_70 VNB N_VGND_c_1359_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=1.72 $Y2=2.235
cc_71 VNB N_VGND_c_1360_n 0.108917f $X=-0.19 $Y=-0.24 $X2=1.715 $Y2=0.34
cc_72 VNB N_VGND_c_1361_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=1.83 $Y2=2.32
cc_73 VNB N_VGND_c_1362_n 0.0173951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1363_n 0.0285145f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1364_n 0.485338f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1365_n 0.00430622f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VPB N_A_79_21#_c_165_n 0.0209226f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_78 VPB N_A_79_21#_c_166_n 0.018106f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_79 VPB N_A_79_21#_c_160_n 0.00159805f $X=-0.19 $Y=1.305 $X2=1.145 $Y2=1.16
cc_80 VPB N_A_79_21#_c_168_n 0.0038652f $X=-0.19 $Y=1.305 $X2=1.72 $Y2=2.235
cc_81 VPB N_A_79_21#_c_169_n 0.00112766f $X=-0.19 $Y=1.305 $X2=1.83 $Y2=2.32
cc_82 VPB N_A_79_21#_c_170_n 0.0124849f $X=-0.19 $Y=1.305 $X2=2.925 $Y2=2.32
cc_83 VPB N_A_79_21#_c_164_n 0.0313336f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.202
cc_84 VPB N_C_M1003_g 0.0318426f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_85 VPB N_C_c_267_n 0.0408591f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_86 VPB N_C_c_269_n 0.00707558f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.985
cc_87 VPB N_C_c_270_n 0.026206f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_88 VPB C 0.00361068f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=0.865
cc_89 VPB N_A_328_93#_c_326_n 0.034375f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_90 VPB N_A_328_93#_c_328_n 0.00441836f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_91 VPB N_A_328_93#_c_332_n 0.00959731f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.875
cc_92 VPB N_A_328_93#_c_333_n 0.00173389f $X=-0.19 $Y=1.305 $X2=1.145 $Y2=1.16
cc_93 VPB N_A_328_93#_c_334_n 0.00184072f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=0.78
cc_94 VPB N_A_328_93#_c_329_n 2.68624e-19 $X=-0.19 $Y=1.305 $X2=1.605 $Y2=0.425
cc_95 VPB N_A_885_297#_c_412_n 0.0182699f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_96 VPB N_A_885_297#_c_399_n 0.0108183f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.985
cc_97 VPB N_A_885_297#_c_414_n 0.0248891f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_98 VPB N_A_885_297#_c_400_n 0.0104543f $X=-0.19 $Y=1.305 $X2=1.145 $Y2=1.16
cc_99 VPB N_A_885_297#_c_401_n 0.00824048f $X=-0.19 $Y=1.305 $X2=1.145 $Y2=1.16
cc_100 VPB N_A_885_297#_c_417_n 0.00601461f $X=-0.19 $Y=1.305 $X2=1.265 $Y2=1.96
cc_101 VPB N_A_885_297#_c_411_n 0.00321756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_B_c_589_n 0.0216593f $X=-0.19 $Y=1.305 $X2=2.855 $Y2=0.245
cc_103 VPB N_B_c_583_n 0.00748587f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_104 VPB N_B_M1010_g 0.0155244f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_105 VPB N_B_c_592_n 0.11933f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_106 VPB N_B_c_593_n 0.0170126f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=0.865
cc_107 VPB N_B_c_594_n 0.00984484f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=0.78
cc_108 VPB N_B_c_595_n 0.00749406f $X=-0.19 $Y=1.305 $X2=1.265 $Y2=0.78
cc_109 VPB N_B_M1006_g 0.0137783f $X=-0.19 $Y=1.305 $X2=1.605 $Y2=0.425
cc_110 VPB N_B_c_585_n 0.00875008f $X=-0.19 $Y=1.305 $X2=1.72 $Y2=2.235
cc_111 VPB N_B_c_586_n 0.00140378f $X=-0.19 $Y=1.305 $X2=2.925 $Y2=2.32
cc_112 VPB N_B_c_587_n 0.00481946f $X=-0.19 $Y=1.305 $X2=2.925 $Y2=2.32
cc_113 VPB N_B_c_600_n 9.50066e-19 $X=-0.19 $Y=1.305 $X2=2.88 $Y2=0.355
cc_114 VPB B 0.0084098f $X=-0.19 $Y=1.305 $X2=3 $Y2=0.355
cc_115 VPB N_A_c_717_n 0.0273239f $X=-0.19 $Y=1.305 $X2=2.855 $Y2=0.245
cc_116 VPB A 0.00309532f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_117 VPB N_A_1003_297#_c_753_n 0.034682f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_118 VPB N_A_1003_297#_c_754_n 0.00274744f $X=-0.19 $Y=1.305 $X2=1.155
+ $Y2=1.16
cc_119 VPB N_A_1003_297#_c_762_n 0.00190108f $X=-0.19 $Y=1.305 $X2=1.145
+ $Y2=1.16
cc_120 VPB N_A_1003_297#_c_757_n 0.00169546f $X=-0.19 $Y=1.305 $X2=1.605
+ $Y2=0.695
cc_121 VPB N_A_1003_297#_c_764_n 0.00176316f $X=-0.19 $Y=1.305 $X2=1.72
+ $Y2=2.045
cc_122 VPB N_VPWR_c_885_n 0.0104612f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_123 VPB N_VPWR_c_886_n 0.0450137f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.985
cc_124 VPB N_VPWR_c_887_n 0.00709021f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.16
cc_125 VPB N_VPWR_c_888_n 0.00743637f $X=-0.19 $Y=1.305 $X2=1.265 $Y2=0.78
cc_126 VPB N_VPWR_c_889_n 4.89207e-19 $X=-0.19 $Y=1.305 $X2=1.605 $Y2=0.695
cc_127 VPB N_VPWR_c_890_n 0.0625838f $X=-0.19 $Y=1.305 $X2=2.68 $Y2=0.34
cc_128 VPB N_VPWR_c_891_n 0.00513206f $X=-0.19 $Y=1.305 $X2=1.715 $Y2=0.34
cc_129 VPB N_VPWR_c_892_n 0.0170895f $X=-0.19 $Y=1.305 $X2=2.925 $Y2=2.32
cc_130 VPB N_VPWR_c_893_n 0.0974174f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_894_n 0.0241631f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_884_n 0.0747448f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_896_n 0.00613115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_897_n 0.00442675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_X_c_981_n 9.42863e-19 $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_136 VPB N_A_453_325#_c_1001_n 0.0110171f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_137 VPB N_A_453_325#_c_997_n 0.00805098f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=0.78
cc_138 VPB N_A_453_325#_c_1003_n 0.00296592f $X=-0.19 $Y=1.305 $X2=1.265
+ $Y2=0.78
cc_139 VPB N_A_453_325#_c_1004_n 0.00293344f $X=-0.19 $Y=1.305 $X2=1.605
+ $Y2=0.425
cc_140 VPB N_A_453_325#_c_1005_n 0.0106403f $X=-0.19 $Y=1.305 $X2=1.605
+ $Y2=0.695
cc_141 VPB N_A_453_325#_c_1006_n 0.00172555f $X=-0.19 $Y=1.305 $X2=1.72
+ $Y2=2.045
cc_142 VPB N_A_453_325#_c_998_n 0.00149669f $X=-0.19 $Y=1.305 $X2=2.68 $Y2=0.34
cc_143 VPB N_A_453_325#_c_1008_n 0.024394f $X=-0.19 $Y=1.305 $X2=2.925 $Y2=2.32
cc_144 VPB N_A_453_325#_c_1009_n 3.60787e-19 $X=-0.19 $Y=1.305 $X2=0.985
+ $Y2=1.202
cc_145 VPB N_A_453_325#_c_1010_n 3.41339e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_477_49#_c_1150_n 0.00148953f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_147 VPB N_A_477_49#_c_1154_n 0.00271724f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_148 VPB N_A_477_49#_c_1155_n 8.50776e-19 $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.16
cc_149 VPB N_A_477_49#_c_1151_n 0.00212375f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=0.78
cc_150 VPB N_A_477_49#_c_1157_n 0.0147524f $X=-0.19 $Y=1.305 $X2=2.925 $Y2=2.32
cc_151 VPB N_A_477_49#_c_1158_n 0.00333347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_477_49#_c_1159_n 0.008761f $X=-0.19 $Y=1.305 $X2=3 $Y2=0.37
cc_153 VPB N_A_477_49#_c_1160_n 0.00154407f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.202
cc_154 VPB N_A_1286_297#_c_1286_n 0.00455825f $X=-0.19 $Y=1.305 $X2=0.985
+ $Y2=1.985
cc_155 VPB N_A_1286_297#_c_1290_n 0.0147295f $X=-0.19 $Y=1.305 $X2=1.145
+ $Y2=1.16
cc_156 VPB N_A_1286_297#_c_1287_n 0.0231133f $X=-0.19 $Y=1.305 $X2=1.61 $Y2=1.96
cc_157 VPB N_A_1286_297#_c_1292_n 0.0101148f $X=-0.19 $Y=1.305 $X2=1.72
+ $Y2=2.235
cc_158 N_A_79_21#_c_159_n N_C_c_266_n 0.0128457f $X=0.99 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_159 N_A_79_21#_c_160_n N_C_c_266_n 0.00138941f $X=1.145 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_160 N_A_79_21#_c_174_p N_C_c_266_n 0.0121405f $X=1.495 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_161 N_A_79_21#_c_161_n N_C_c_266_n 0.0106633f $X=1.605 $Y=0.695 $X2=-0.19
+ $Y2=-0.24
cc_162 N_A_79_21#_c_162_n N_C_c_266_n 0.00609621f $X=1.715 $Y=0.34 $X2=-0.19
+ $Y2=-0.24
cc_163 N_A_79_21#_c_166_n N_C_M1003_g 0.0187374f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_79_21#_c_160_n N_C_M1003_g 0.00567296f $X=1.145 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_79_21#_c_179_p N_C_M1003_g 0.0133831f $X=1.61 $Y=1.96 $X2=0 $Y2=0
cc_166 N_A_79_21#_c_168_n N_C_M1003_g 0.0075271f $X=1.72 $Y=2.235 $X2=0 $Y2=0
cc_167 N_A_79_21#_c_169_n N_C_M1003_g 0.00744783f $X=1.83 $Y=2.32 $X2=0 $Y2=0
cc_168 N_A_79_21#_c_170_n N_C_c_267_n 0.0112964f $X=2.925 $Y=2.32 $X2=0 $Y2=0
cc_169 N_A_79_21#_c_183_p N_C_c_268_n 0.0106037f $X=2.88 $Y=0.355 $X2=0 $Y2=0
cc_170 N_A_79_21#_c_160_n N_C_c_269_n 0.00252367f $X=1.145 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_79_21#_c_164_n N_C_c_269_n 0.0263225f $X=0.99 $Y=1.202 $X2=0 $Y2=0
cc_172 N_A_79_21#_c_163_n N_C_c_270_n 0.011137f $X=2.68 $Y=0.355 $X2=0 $Y2=0
cc_173 N_A_79_21#_c_163_n C 0.00342613f $X=2.68 $Y=0.355 $X2=0 $Y2=0
cc_174 N_A_79_21#_c_174_p N_A_328_93#_M1009_d 0.00226043f $X=1.495 $Y=0.78
+ $X2=-0.19 $Y2=-0.24
cc_175 N_A_79_21#_c_161_n N_A_328_93#_M1009_d 0.00618081f $X=1.605 $Y=0.695
+ $X2=-0.19 $Y2=-0.24
cc_176 N_A_79_21#_c_179_p N_A_328_93#_M1003_d 0.00416203f $X=1.61 $Y=1.96 $X2=0
+ $Y2=0
cc_177 N_A_79_21#_c_168_n N_A_328_93#_M1003_d 0.00266846f $X=1.72 $Y=2.235 $X2=0
+ $Y2=0
cc_178 N_A_79_21#_c_170_n N_A_328_93#_c_326_n 0.0116412f $X=2.925 $Y=2.32 $X2=0
+ $Y2=0
cc_179 N_A_79_21#_c_193_p N_A_328_93#_c_327_n 0.00377914f $X=3 $Y=0.37 $X2=0
+ $Y2=0
cc_180 N_A_79_21#_c_174_p N_A_328_93#_c_342_n 0.00409956f $X=1.495 $Y=0.78 $X2=0
+ $Y2=0
cc_181 N_A_79_21#_c_179_p N_A_328_93#_c_342_n 0.0200253f $X=1.61 $Y=1.96 $X2=0
+ $Y2=0
cc_182 N_A_79_21#_c_170_n N_A_328_93#_c_342_n 0.00176797f $X=2.925 $Y=2.32 $X2=0
+ $Y2=0
cc_183 N_A_79_21#_c_160_n N_A_328_93#_c_328_n 0.018047f $X=1.145 $Y=1.16 $X2=0
+ $Y2=0
cc_184 N_A_79_21#_c_174_p N_A_328_93#_c_328_n 0.0138141f $X=1.495 $Y=0.78 $X2=0
+ $Y2=0
cc_185 N_A_79_21#_c_161_n N_A_328_93#_c_328_n 0.00736858f $X=1.605 $Y=0.695
+ $X2=0 $Y2=0
cc_186 N_A_79_21#_c_163_n N_A_328_93#_c_328_n 0.0130244f $X=2.68 $Y=0.355 $X2=0
+ $Y2=0
cc_187 N_A_79_21#_c_164_n N_A_328_93#_c_328_n 7.42235e-19 $X=0.99 $Y=1.202 $X2=0
+ $Y2=0
cc_188 N_A_79_21#_M1016_d N_A_328_93#_c_332_n 0.00779963f $X=2.78 $Y=1.625 $X2=0
+ $Y2=0
cc_189 N_A_79_21#_c_170_n N_A_328_93#_c_332_n 0.0039224f $X=2.925 $Y=2.32 $X2=0
+ $Y2=0
cc_190 N_A_79_21#_M1016_d N_A_328_93#_c_333_n 5.89264e-19 $X=2.78 $Y=1.625 $X2=0
+ $Y2=0
cc_191 N_A_79_21#_c_170_n N_A_328_93#_c_334_n 0.00633062f $X=2.925 $Y=2.32 $X2=0
+ $Y2=0
cc_192 N_A_79_21#_c_160_n N_VPWR_M1019_s 0.00465367f $X=1.145 $Y=1.16 $X2=0
+ $Y2=0
cc_193 N_A_79_21#_c_179_p N_VPWR_M1019_s 0.00886232f $X=1.61 $Y=1.96 $X2=0 $Y2=0
cc_194 N_A_79_21#_c_208_p N_VPWR_M1019_s 0.00150909f $X=1.265 $Y=1.96 $X2=0
+ $Y2=0
cc_195 N_A_79_21#_c_165_n N_VPWR_c_886_n 0.00341708f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_196 N_A_79_21#_c_165_n N_VPWR_c_887_n 4.59975e-19 $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_197 N_A_79_21#_c_166_n N_VPWR_c_887_n 0.00898123f $X=0.985 $Y=1.41 $X2=0
+ $Y2=0
cc_198 N_A_79_21#_c_179_p N_VPWR_c_887_n 0.0126548f $X=1.61 $Y=1.96 $X2=0 $Y2=0
cc_199 N_A_79_21#_c_208_p N_VPWR_c_887_n 0.0135851f $X=1.265 $Y=1.96 $X2=0 $Y2=0
cc_200 N_A_79_21#_c_168_n N_VPWR_c_887_n 0.00145799f $X=1.72 $Y=2.235 $X2=0
+ $Y2=0
cc_201 N_A_79_21#_c_169_n N_VPWR_c_887_n 0.0137789f $X=1.83 $Y=2.32 $X2=0 $Y2=0
cc_202 N_A_79_21#_c_179_p N_VPWR_c_890_n 0.00233941f $X=1.61 $Y=1.96 $X2=0 $Y2=0
cc_203 N_A_79_21#_c_169_n N_VPWR_c_890_n 0.0109705f $X=1.83 $Y=2.32 $X2=0 $Y2=0
cc_204 N_A_79_21#_c_170_n N_VPWR_c_890_n 0.0597844f $X=2.925 $Y=2.32 $X2=0 $Y2=0
cc_205 N_A_79_21#_c_165_n N_VPWR_c_892_n 0.00643255f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_206 N_A_79_21#_c_166_n N_VPWR_c_892_n 0.00583607f $X=0.985 $Y=1.41 $X2=0
+ $Y2=0
cc_207 N_A_79_21#_c_165_n N_VPWR_c_884_n 0.0119906f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A_79_21#_c_166_n N_VPWR_c_884_n 0.00983716f $X=0.985 $Y=1.41 $X2=0
+ $Y2=0
cc_209 N_A_79_21#_c_179_p N_VPWR_c_884_n 0.00553584f $X=1.61 $Y=1.96 $X2=0 $Y2=0
cc_210 N_A_79_21#_c_208_p N_VPWR_c_884_n 0.00101474f $X=1.265 $Y=1.96 $X2=0
+ $Y2=0
cc_211 N_A_79_21#_c_169_n N_VPWR_c_884_n 0.00809357f $X=1.83 $Y=2.32 $X2=0 $Y2=0
cc_212 N_A_79_21#_c_170_n N_VPWR_c_884_n 0.0473531f $X=2.925 $Y=2.32 $X2=0 $Y2=0
cc_213 N_A_79_21#_c_158_n N_X_c_981_n 0.0064953f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A_79_21#_c_165_n N_X_c_981_n 0.0167863f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A_79_21#_c_166_n N_X_c_981_n 6.38052e-19 $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A_79_21#_c_159_n N_X_c_981_n 0.0017469f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A_79_21#_c_160_n N_X_c_981_n 0.0563142f $X=1.145 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A_79_21#_c_164_n N_X_c_981_n 0.0450472f $X=0.99 $Y=1.202 $X2=0 $Y2=0
cc_219 N_A_79_21#_c_170_n N_A_453_325#_M1016_s 0.00736441f $X=2.925 $Y=2.32
+ $X2=0 $Y2=0
cc_220 N_A_79_21#_M1016_d N_A_453_325#_c_1001_n 0.00510383f $X=2.78 $Y=1.625
+ $X2=0 $Y2=0
cc_221 N_A_79_21#_c_179_p N_A_453_325#_c_1001_n 0.00831987f $X=1.61 $Y=1.96
+ $X2=0 $Y2=0
cc_222 N_A_79_21#_c_168_n N_A_453_325#_c_1001_n 9.56599e-19 $X=1.72 $Y=2.235
+ $X2=0 $Y2=0
cc_223 N_A_79_21#_c_170_n N_A_453_325#_c_1001_n 0.0571361f $X=2.925 $Y=2.32
+ $X2=0 $Y2=0
cc_224 N_A_79_21#_c_193_p N_A_453_325#_c_995_n 0.0118982f $X=3 $Y=0.37 $X2=0
+ $Y2=0
cc_225 N_A_79_21#_c_163_n N_A_477_49#_M1007_s 0.00652268f $X=2.68 $Y=0.355
+ $X2=-0.19 $Y2=-0.24
cc_226 N_A_79_21#_M1007_d N_A_477_49#_c_1162_n 0.00636386f $X=2.855 $Y=0.245
+ $X2=0 $Y2=0
cc_227 N_A_79_21#_c_193_p N_A_477_49#_c_1162_n 0.0116342f $X=3 $Y=0.37 $X2=0
+ $Y2=0
cc_228 N_A_79_21#_c_183_p N_A_477_49#_c_1152_n 0.0116342f $X=2.88 $Y=0.355 $X2=0
+ $Y2=0
cc_229 N_A_79_21#_c_163_n N_A_477_49#_c_1152_n 0.0181831f $X=2.68 $Y=0.355 $X2=0
+ $Y2=0
cc_230 N_A_79_21#_c_160_n N_VGND_M1023_d 2.81692e-19 $X=1.145 $Y=1.16 $X2=0
+ $Y2=0
cc_231 N_A_79_21#_c_174_p N_VGND_M1023_d 0.00889686f $X=1.495 $Y=0.78 $X2=0
+ $Y2=0
cc_232 N_A_79_21#_c_246_p N_VGND_M1023_d 0.00167046f $X=1.265 $Y=0.78 $X2=0
+ $Y2=0
cc_233 N_A_79_21#_c_158_n N_VGND_c_1354_n 0.00599948f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_234 N_A_79_21#_c_158_n N_VGND_c_1355_n 8.28113e-19 $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_235 N_A_79_21#_c_159_n N_VGND_c_1355_n 0.00992764f $X=0.99 $Y=0.995 $X2=0
+ $Y2=0
cc_236 N_A_79_21#_c_174_p N_VGND_c_1355_n 0.0045481f $X=1.495 $Y=0.78 $X2=0
+ $Y2=0
cc_237 N_A_79_21#_c_246_p N_VGND_c_1355_n 0.013837f $X=1.265 $Y=0.78 $X2=0 $Y2=0
cc_238 N_A_79_21#_c_161_n N_VGND_c_1355_n 0.00742455f $X=1.605 $Y=0.695 $X2=0
+ $Y2=0
cc_239 N_A_79_21#_c_162_n N_VGND_c_1355_n 0.0142402f $X=1.715 $Y=0.34 $X2=0
+ $Y2=0
cc_240 N_A_79_21#_c_164_n N_VGND_c_1355_n 7.57381e-19 $X=0.99 $Y=1.202 $X2=0
+ $Y2=0
cc_241 N_A_79_21#_c_174_p N_VGND_c_1358_n 0.00219715f $X=1.495 $Y=0.78 $X2=0
+ $Y2=0
cc_242 N_A_79_21#_c_162_n N_VGND_c_1358_n 0.0156439f $X=1.715 $Y=0.34 $X2=0
+ $Y2=0
cc_243 N_A_79_21#_c_163_n N_VGND_c_1358_n 0.0876356f $X=2.68 $Y=0.355 $X2=0
+ $Y2=0
cc_244 N_A_79_21#_c_158_n N_VGND_c_1362_n 0.00585385f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_A_79_21#_c_159_n N_VGND_c_1362_n 0.0046653f $X=0.99 $Y=0.995 $X2=0
+ $Y2=0
cc_246 N_A_79_21#_c_158_n N_VGND_c_1364_n 0.0118559f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_247 N_A_79_21#_c_159_n N_VGND_c_1364_n 0.00821929f $X=0.99 $Y=0.995 $X2=0
+ $Y2=0
cc_248 N_A_79_21#_c_174_p N_VGND_c_1364_n 0.00486078f $X=1.495 $Y=0.78 $X2=0
+ $Y2=0
cc_249 N_A_79_21#_c_246_p N_VGND_c_1364_n 9.90971e-19 $X=1.265 $Y=0.78 $X2=0
+ $Y2=0
cc_250 N_A_79_21#_c_162_n N_VGND_c_1364_n 0.00844855f $X=1.715 $Y=0.34 $X2=0
+ $Y2=0
cc_251 N_A_79_21#_c_163_n N_VGND_c_1364_n 0.0532675f $X=2.68 $Y=0.355 $X2=0
+ $Y2=0
cc_252 N_C_c_267_n N_A_328_93#_c_326_n 0.0592216f $X=2.69 $Y=1.55 $X2=0 $Y2=0
cc_253 C N_A_328_93#_c_326_n 2.69094e-19 $X=2.44 $Y=1.105 $X2=0 $Y2=0
cc_254 N_C_c_268_n N_A_328_93#_c_327_n 0.0256383f $X=2.78 $Y=0.995 $X2=0 $Y2=0
cc_255 N_C_M1003_g N_A_328_93#_c_342_n 0.0114423f $X=1.59 $Y=1.805 $X2=0 $Y2=0
cc_256 N_C_c_270_n N_A_328_93#_c_342_n 0.00634718f $X=2.59 $Y=1.16 $X2=0 $Y2=0
cc_257 N_C_c_266_n N_A_328_93#_c_328_n 0.0043646f $X=1.565 $Y=0.995 $X2=0 $Y2=0
cc_258 N_C_M1003_g N_A_328_93#_c_328_n 0.00203559f $X=1.59 $Y=1.805 $X2=0 $Y2=0
cc_259 N_C_c_267_n N_A_328_93#_c_328_n 0.00508695f $X=2.69 $Y=1.55 $X2=0 $Y2=0
cc_260 N_C_c_268_n N_A_328_93#_c_328_n 0.00235914f $X=2.78 $Y=0.995 $X2=0 $Y2=0
cc_261 N_C_c_269_n N_A_328_93#_c_328_n 0.0020376f $X=1.59 $Y=1.202 $X2=0 $Y2=0
cc_262 N_C_c_270_n N_A_328_93#_c_328_n 0.0266304f $X=2.59 $Y=1.16 $X2=0 $Y2=0
cc_263 C N_A_328_93#_c_328_n 0.0187897f $X=2.44 $Y=1.105 $X2=0 $Y2=0
cc_264 N_C_c_267_n N_A_328_93#_c_332_n 0.0172192f $X=2.69 $Y=1.55 $X2=0 $Y2=0
cc_265 N_C_c_270_n N_A_328_93#_c_332_n 0.00858517f $X=2.59 $Y=1.16 $X2=0 $Y2=0
cc_266 C N_A_328_93#_c_332_n 0.0378709f $X=2.44 $Y=1.105 $X2=0 $Y2=0
cc_267 N_C_c_267_n N_A_328_93#_c_333_n 0.00427971f $X=2.69 $Y=1.55 $X2=0 $Y2=0
cc_268 N_C_c_267_n N_A_328_93#_c_329_n 0.00351803f $X=2.69 $Y=1.55 $X2=0 $Y2=0
cc_269 C N_A_328_93#_c_329_n 0.0207158f $X=2.44 $Y=1.105 $X2=0 $Y2=0
cc_270 N_C_M1003_g N_VPWR_c_887_n 0.00212825f $X=1.59 $Y=1.805 $X2=0 $Y2=0
cc_271 N_C_M1003_g N_VPWR_c_890_n 0.00514356f $X=1.59 $Y=1.805 $X2=0 $Y2=0
cc_272 N_C_c_267_n N_VPWR_c_890_n 0.00427564f $X=2.69 $Y=1.55 $X2=0 $Y2=0
cc_273 N_C_M1003_g N_VPWR_c_884_n 0.00682402f $X=1.59 $Y=1.805 $X2=0 $Y2=0
cc_274 N_C_c_267_n N_VPWR_c_884_n 0.00784458f $X=2.69 $Y=1.55 $X2=0 $Y2=0
cc_275 N_C_M1003_g N_A_453_325#_c_1001_n 9.4239e-19 $X=1.59 $Y=1.805 $X2=0 $Y2=0
cc_276 N_C_c_267_n N_A_453_325#_c_1001_n 0.0102234f $X=2.69 $Y=1.55 $X2=0 $Y2=0
cc_277 N_C_c_268_n N_A_477_49#_c_1162_n 0.00802637f $X=2.78 $Y=0.995 $X2=0 $Y2=0
cc_278 C N_A_477_49#_c_1162_n 0.00486972f $X=2.44 $Y=1.105 $X2=0 $Y2=0
cc_279 N_C_c_268_n N_A_477_49#_c_1152_n 0.00374405f $X=2.78 $Y=0.995 $X2=0 $Y2=0
cc_280 N_C_c_270_n N_A_477_49#_c_1152_n 0.00655613f $X=2.59 $Y=1.16 $X2=0 $Y2=0
cc_281 C N_A_477_49#_c_1152_n 0.0290801f $X=2.44 $Y=1.105 $X2=0 $Y2=0
cc_282 N_C_c_266_n N_VGND_c_1355_n 0.00139578f $X=1.565 $Y=0.995 $X2=0 $Y2=0
cc_283 N_C_c_266_n N_VGND_c_1358_n 8.79444e-19 $X=1.565 $Y=0.995 $X2=0 $Y2=0
cc_284 N_C_c_268_n N_VGND_c_1358_n 0.00357877f $X=2.78 $Y=0.995 $X2=0 $Y2=0
cc_285 N_C_c_268_n N_VGND_c_1364_n 0.00671982f $X=2.78 $Y=0.995 $X2=0 $Y2=0
cc_286 N_A_328_93#_c_326_n N_VPWR_c_888_n 0.00632978f $X=3.225 $Y=1.41 $X2=0
+ $Y2=0
cc_287 N_A_328_93#_c_326_n N_VPWR_c_890_n 0.00412251f $X=3.225 $Y=1.41 $X2=0
+ $Y2=0
cc_288 N_A_328_93#_c_326_n N_VPWR_c_884_n 0.00595559f $X=3.225 $Y=1.41 $X2=0
+ $Y2=0
cc_289 N_A_328_93#_c_332_n N_A_453_325#_M1016_s 0.00373918f $X=3.01 $Y=1.62
+ $X2=0 $Y2=0
cc_290 N_A_328_93#_c_326_n N_A_453_325#_c_1001_n 0.0182447f $X=3.225 $Y=1.41
+ $X2=0 $Y2=0
cc_291 N_A_328_93#_c_332_n N_A_453_325#_c_1001_n 0.0556467f $X=3.01 $Y=1.62
+ $X2=0 $Y2=0
cc_292 N_A_328_93#_c_329_n N_A_453_325#_c_1001_n 0.00386917f $X=3.2 $Y=1.16
+ $X2=0 $Y2=0
cc_293 N_A_328_93#_c_327_n N_A_453_325#_c_995_n 0.00383691f $X=3.22 $Y=0.995
+ $X2=0 $Y2=0
cc_294 N_A_328_93#_c_327_n N_A_453_325#_c_996_n 0.00468917f $X=3.22 $Y=0.995
+ $X2=0 $Y2=0
cc_295 N_A_328_93#_c_326_n N_A_453_325#_c_997_n 0.00449957f $X=3.225 $Y=1.41
+ $X2=0 $Y2=0
cc_296 N_A_328_93#_c_326_n N_A_477_49#_c_1162_n 0.00407382f $X=3.225 $Y=1.41
+ $X2=0 $Y2=0
cc_297 N_A_328_93#_c_327_n N_A_477_49#_c_1162_n 0.0134027f $X=3.22 $Y=0.995
+ $X2=0 $Y2=0
cc_298 N_A_328_93#_c_329_n N_A_477_49#_c_1162_n 0.017913f $X=3.2 $Y=1.16 $X2=0
+ $Y2=0
cc_299 N_A_328_93#_c_326_n N_A_477_49#_c_1150_n 0.00889685f $X=3.225 $Y=1.41
+ $X2=0 $Y2=0
cc_300 N_A_328_93#_c_327_n N_A_477_49#_c_1150_n 0.00652586f $X=3.22 $Y=0.995
+ $X2=0 $Y2=0
cc_301 N_A_328_93#_c_333_n N_A_477_49#_c_1150_n 0.00218396f $X=3.095 $Y=1.535
+ $X2=0 $Y2=0
cc_302 N_A_328_93#_c_329_n N_A_477_49#_c_1150_n 0.0247426f $X=3.2 $Y=1.16 $X2=0
+ $Y2=0
cc_303 N_A_328_93#_c_327_n N_A_477_49#_c_1152_n 5.34088e-19 $X=3.22 $Y=0.995
+ $X2=0 $Y2=0
cc_304 N_A_328_93#_c_328_n N_A_477_49#_c_1152_n 0.0151384f $X=1.97 $Y=0.76 $X2=0
+ $Y2=0
cc_305 N_A_328_93#_c_332_n N_A_477_49#_c_1158_n 5.94479e-19 $X=3.01 $Y=1.62
+ $X2=0 $Y2=0
cc_306 N_A_328_93#_c_333_n N_A_477_49#_c_1158_n 6.54862e-19 $X=3.095 $Y=1.535
+ $X2=0 $Y2=0
cc_307 N_A_328_93#_c_326_n N_A_477_49#_c_1159_n 0.00719438f $X=3.225 $Y=1.41
+ $X2=0 $Y2=0
cc_308 N_A_328_93#_c_332_n N_A_477_49#_c_1159_n 0.0102953f $X=3.01 $Y=1.62 $X2=0
+ $Y2=0
cc_309 N_A_328_93#_c_333_n N_A_477_49#_c_1159_n 0.00669828f $X=3.095 $Y=1.535
+ $X2=0 $Y2=0
cc_310 N_A_328_93#_c_327_n N_VGND_c_1358_n 0.00414846f $X=3.22 $Y=0.995 $X2=0
+ $Y2=0
cc_311 N_A_328_93#_c_327_n N_VGND_c_1364_n 0.00723015f $X=3.22 $Y=0.995 $X2=0
+ $Y2=0
cc_312 N_A_885_297#_c_417_n N_B_c_589_n 0.00852064f $X=4.73 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_313 N_A_885_297#_c_411_n N_B_c_589_n 8.18494e-19 $X=4.79 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_314 N_A_885_297#_c_421_p N_B_M1022_g 0.00381578f $X=4.815 $Y=0.85 $X2=0 $Y2=0
cc_315 N_A_885_297#_c_411_n N_B_M1022_g 0.0178285f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_316 N_A_885_297#_c_403_n N_B_c_582_n 0.0050801f $X=6.005 $Y=0.85 $X2=0 $Y2=0
cc_317 N_A_885_297#_c_411_n N_B_c_582_n 0.0122706f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A_885_297#_c_417_n N_B_c_583_n 0.00748737f $X=4.73 $Y=1.58 $X2=0 $Y2=0
cc_319 N_A_885_297#_c_411_n N_B_c_583_n 0.00955042f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_320 N_A_885_297#_c_412_n N_B_M1010_g 0.0119272f $X=6.34 $Y=1.41 $X2=0 $Y2=0
cc_321 N_A_885_297#_M1001_g N_B_M1015_g 0.0102876f $X=6.365 $Y=0.455 $X2=0 $Y2=0
cc_322 N_A_885_297#_c_400_n N_B_M1015_g 0.021209f $X=6.24 $Y=1.16 $X2=0 $Y2=0
cc_323 N_A_885_297#_c_402_n N_B_M1015_g 0.00188578f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_324 N_A_885_297#_c_403_n N_B_M1015_g 0.00148554f $X=6.005 $Y=0.85 $X2=0 $Y2=0
cc_325 N_A_885_297#_c_405_n N_B_M1015_g 6.75018e-19 $X=6.295 $Y=0.85 $X2=0 $Y2=0
cc_326 N_A_885_297#_c_406_n N_B_M1015_g 0.00122796f $X=6.15 $Y=0.85 $X2=0 $Y2=0
cc_327 N_A_885_297#_c_412_n N_B_c_592_n 0.0105804f $X=6.34 $Y=1.41 $X2=0 $Y2=0
cc_328 N_A_885_297#_c_414_n N_B_c_592_n 0.0048792f $X=7.83 $Y=1.57 $X2=0 $Y2=0
cc_329 N_A_885_297#_c_412_n N_B_c_594_n 0.00163254f $X=6.34 $Y=1.41 $X2=0 $Y2=0
cc_330 N_A_885_297#_c_399_n N_B_c_594_n 0.0028078f $X=7.83 $Y=1.47 $X2=0 $Y2=0
cc_331 N_A_885_297#_c_414_n N_B_c_595_n 0.0028078f $X=7.83 $Y=1.57 $X2=0 $Y2=0
cc_332 N_A_885_297#_c_412_n N_B_M1006_g 0.00911296f $X=6.34 $Y=1.41 $X2=0 $Y2=0
cc_333 N_A_885_297#_c_414_n N_B_M1006_g 0.0205449f $X=7.83 $Y=1.57 $X2=0 $Y2=0
cc_334 N_A_885_297#_c_401_n N_B_c_585_n 0.00181049f $X=6.34 $Y=1.202 $X2=0 $Y2=0
cc_335 N_A_885_297#_c_399_n N_B_c_586_n 0.00248427f $X=7.83 $Y=1.47 $X2=0 $Y2=0
cc_336 N_A_885_297#_c_404_n N_B_c_586_n 0.00731236f $X=7.485 $Y=0.85 $X2=0 $Y2=0
cc_337 N_A_885_297#_c_408_n N_B_c_586_n 0.021521f $X=7.63 $Y=0.85 $X2=0 $Y2=0
cc_338 N_A_885_297#_c_409_n N_B_c_586_n 2.70696e-19 $X=7.75 $Y=1.11 $X2=0 $Y2=0
cc_339 N_A_885_297#_c_399_n N_B_c_587_n 0.00187722f $X=7.83 $Y=1.47 $X2=0 $Y2=0
cc_340 N_A_885_297#_c_401_n N_B_c_587_n 0.00816231f $X=6.34 $Y=1.202 $X2=0 $Y2=0
cc_341 N_A_885_297#_c_404_n N_B_c_587_n 0.00130216f $X=7.485 $Y=0.85 $X2=0 $Y2=0
cc_342 N_A_885_297#_c_408_n N_B_c_587_n 0.00172718f $X=7.63 $Y=0.85 $X2=0 $Y2=0
cc_343 N_A_885_297#_c_409_n N_B_c_587_n 0.0173414f $X=7.75 $Y=1.11 $X2=0 $Y2=0
cc_344 N_A_885_297#_c_399_n B 0.0013799f $X=7.83 $Y=1.47 $X2=0 $Y2=0
cc_345 N_A_885_297#_c_414_n B 0.00512663f $X=7.83 $Y=1.57 $X2=0 $Y2=0
cc_346 N_A_885_297#_c_404_n B 0.00417695f $X=7.485 $Y=0.85 $X2=0 $Y2=0
cc_347 N_A_885_297#_c_407_n B 0.00235209f $X=7.63 $Y=0.85 $X2=0 $Y2=0
cc_348 N_A_885_297#_c_408_n B 0.0183366f $X=7.63 $Y=0.85 $X2=0 $Y2=0
cc_349 N_A_885_297#_c_409_n B 8.1069e-19 $X=7.75 $Y=1.11 $X2=0 $Y2=0
cc_350 N_A_885_297#_M1001_g N_B_c_588_n 0.00816231f $X=6.365 $Y=0.455 $X2=0
+ $Y2=0
cc_351 N_A_885_297#_c_404_n N_B_c_588_n 0.0076315f $X=7.485 $Y=0.85 $X2=0 $Y2=0
cc_352 N_A_885_297#_c_407_n N_B_c_588_n 0.00141075f $X=7.63 $Y=0.85 $X2=0 $Y2=0
cc_353 N_A_885_297#_c_408_n N_B_c_588_n 0.00206736f $X=7.63 $Y=0.85 $X2=0 $Y2=0
cc_354 N_A_885_297#_c_409_n N_B_c_588_n 0.00135765f $X=7.75 $Y=1.11 $X2=0 $Y2=0
cc_355 N_A_885_297#_c_410_n N_B_c_588_n 0.0136423f $X=7.772 $Y=0.945 $X2=0 $Y2=0
cc_356 N_A_885_297#_c_399_n N_A_c_717_n 0.00765017f $X=7.83 $Y=1.47 $X2=-0.19
+ $Y2=-0.24
cc_357 N_A_885_297#_c_414_n N_A_c_717_n 0.0315678f $X=7.83 $Y=1.57 $X2=-0.19
+ $Y2=-0.24
cc_358 N_A_885_297#_c_408_n N_A_c_717_n 6.51299e-19 $X=7.63 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_359 N_A_885_297#_c_409_n N_A_c_717_n 0.0202732f $X=7.75 $Y=1.11 $X2=-0.19
+ $Y2=-0.24
cc_360 N_A_885_297#_c_408_n N_A_c_718_n 2.39914e-19 $X=7.63 $Y=0.85 $X2=0 $Y2=0
cc_361 N_A_885_297#_c_410_n N_A_c_718_n 0.0185553f $X=7.772 $Y=0.945 $X2=0 $Y2=0
cc_362 N_A_885_297#_c_408_n A 0.0137584f $X=7.63 $Y=0.85 $X2=0 $Y2=0
cc_363 N_A_885_297#_c_409_n A 0.00285423f $X=7.75 $Y=1.11 $X2=0 $Y2=0
cc_364 N_A_885_297#_c_403_n N_A_1003_297#_M1015_s 8.58636e-19 $X=6.005 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_365 N_A_885_297#_c_417_n N_A_1003_297#_c_754_n 0.0194501f $X=4.73 $Y=1.58
+ $X2=0 $Y2=0
cc_366 N_A_885_297#_c_403_n N_A_1003_297#_c_754_n 0.0124002f $X=6.005 $Y=0.85
+ $X2=0 $Y2=0
cc_367 N_A_885_297#_c_421_p N_A_1003_297#_c_754_n 5.77119e-19 $X=4.815 $Y=0.85
+ $X2=0 $Y2=0
cc_368 N_A_885_297#_c_411_n N_A_1003_297#_c_754_n 0.0604107f $X=4.79 $Y=0.74
+ $X2=0 $Y2=0
cc_369 N_A_885_297#_c_414_n N_A_1003_297#_c_762_n 0.00416703f $X=7.83 $Y=1.57
+ $X2=0 $Y2=0
cc_370 N_A_885_297#_c_407_n N_A_1003_297#_c_756_n 0.00537182f $X=7.63 $Y=0.85
+ $X2=0 $Y2=0
cc_371 N_A_885_297#_c_408_n N_A_1003_297#_c_756_n 0.0052004f $X=7.63 $Y=0.85
+ $X2=0 $Y2=0
cc_372 N_A_885_297#_c_410_n N_A_1003_297#_c_756_n 0.00186387f $X=7.772 $Y=0.945
+ $X2=0 $Y2=0
cc_373 N_A_885_297#_M1001_g N_A_1003_297#_c_774_n 0.00613906f $X=6.365 $Y=0.455
+ $X2=0 $Y2=0
cc_374 N_A_885_297#_c_402_n N_A_1003_297#_c_774_n 3.69046e-19 $X=6.13 $Y=0.995
+ $X2=0 $Y2=0
cc_375 N_A_885_297#_c_403_n N_A_1003_297#_c_774_n 0.0529767f $X=6.005 $Y=0.85
+ $X2=0 $Y2=0
cc_376 N_A_885_297#_c_404_n N_A_1003_297#_c_774_n 0.0955498f $X=7.485 $Y=0.85
+ $X2=0 $Y2=0
cc_377 N_A_885_297#_c_405_n N_A_1003_297#_c_774_n 0.026662f $X=6.295 $Y=0.85
+ $X2=0 $Y2=0
cc_378 N_A_885_297#_c_406_n N_A_1003_297#_c_774_n 0.00310602f $X=6.15 $Y=0.85
+ $X2=0 $Y2=0
cc_379 N_A_885_297#_c_407_n N_A_1003_297#_c_774_n 0.0266136f $X=7.63 $Y=0.85
+ $X2=0 $Y2=0
cc_380 N_A_885_297#_c_408_n N_A_1003_297#_c_774_n 0.00475925f $X=7.63 $Y=0.85
+ $X2=0 $Y2=0
cc_381 N_A_885_297#_c_410_n N_A_1003_297#_c_774_n 0.00868614f $X=7.772 $Y=0.945
+ $X2=0 $Y2=0
cc_382 N_A_885_297#_c_403_n N_A_1003_297#_c_758_n 0.0261258f $X=6.005 $Y=0.85
+ $X2=0 $Y2=0
cc_383 N_A_885_297#_c_411_n N_A_1003_297#_c_758_n 0.00683584f $X=4.79 $Y=0.74
+ $X2=0 $Y2=0
cc_384 N_A_885_297#_c_403_n N_A_1003_297#_c_759_n 0.00108548f $X=6.005 $Y=0.85
+ $X2=0 $Y2=0
cc_385 N_A_885_297#_c_411_n N_A_1003_297#_c_759_n 0.01151f $X=4.79 $Y=0.74 $X2=0
+ $Y2=0
cc_386 N_A_885_297#_c_410_n N_A_1003_297#_c_787_n 0.00156339f $X=7.772 $Y=0.945
+ $X2=0 $Y2=0
cc_387 N_A_885_297#_c_410_n N_A_1003_297#_c_788_n 0.00805147f $X=7.772 $Y=0.945
+ $X2=0 $Y2=0
cc_388 N_A_885_297#_c_414_n N_VPWR_c_889_n 0.00118007f $X=7.83 $Y=1.57 $X2=0
+ $Y2=0
cc_389 N_A_885_297#_c_414_n N_VPWR_c_893_n 0.00434439f $X=7.83 $Y=1.57 $X2=0
+ $Y2=0
cc_390 N_A_885_297#_M1005_d N_VPWR_c_884_n 0.00367747f $X=4.425 $Y=1.485 $X2=0
+ $Y2=0
cc_391 N_A_885_297#_c_414_n N_VPWR_c_884_n 0.00665931f $X=7.83 $Y=1.57 $X2=0
+ $Y2=0
cc_392 N_A_885_297#_c_403_n N_A_453_325#_M1015_d 0.00134889f $X=6.005 $Y=0.85
+ $X2=0 $Y2=0
cc_393 N_A_885_297#_c_405_n N_A_453_325#_M1015_d 5.4759e-19 $X=6.295 $Y=0.85
+ $X2=0 $Y2=0
cc_394 N_A_885_297#_c_406_n N_A_453_325#_M1015_d 0.00649965f $X=6.15 $Y=0.85
+ $X2=0 $Y2=0
cc_395 N_A_885_297#_c_421_p N_A_453_325#_c_996_n 0.0023462f $X=4.815 $Y=0.85
+ $X2=0 $Y2=0
cc_396 N_A_885_297#_c_411_n N_A_453_325#_c_996_n 0.00358611f $X=4.79 $Y=0.74
+ $X2=0 $Y2=0
cc_397 N_A_885_297#_c_417_n N_A_453_325#_c_997_n 0.0144171f $X=4.73 $Y=1.58
+ $X2=0 $Y2=0
cc_398 N_A_885_297#_c_411_n N_A_453_325#_c_997_n 0.00928178f $X=4.79 $Y=0.74
+ $X2=0 $Y2=0
cc_399 N_A_885_297#_M1005_d N_A_453_325#_c_1003_n 0.00767171f $X=4.425 $Y=1.485
+ $X2=0 $Y2=0
cc_400 N_A_885_297#_c_417_n N_A_453_325#_c_1003_n 0.0315546f $X=4.73 $Y=1.58
+ $X2=0 $Y2=0
cc_401 N_A_885_297#_M1005_d N_A_453_325#_c_1004_n 0.00313827f $X=4.425 $Y=1.485
+ $X2=0 $Y2=0
cc_402 N_A_885_297#_M1005_d N_A_453_325#_c_1006_n 0.00318432f $X=4.425 $Y=1.485
+ $X2=0 $Y2=0
cc_403 N_A_885_297#_c_412_n N_A_453_325#_c_998_n 0.00131578f $X=6.34 $Y=1.41
+ $X2=0 $Y2=0
cc_404 N_A_885_297#_c_400_n N_A_453_325#_c_998_n 6.52616e-19 $X=6.24 $Y=1.16
+ $X2=0 $Y2=0
cc_405 N_A_885_297#_c_401_n N_A_453_325#_c_998_n 3.9697e-19 $X=6.34 $Y=1.202
+ $X2=0 $Y2=0
cc_406 N_A_885_297#_c_402_n N_A_453_325#_c_998_n 0.0160828f $X=6.13 $Y=0.995
+ $X2=0 $Y2=0
cc_407 N_A_885_297#_c_403_n N_A_453_325#_c_998_n 0.00616329f $X=6.005 $Y=0.85
+ $X2=0 $Y2=0
cc_408 N_A_885_297#_c_405_n N_A_453_325#_c_998_n 0.00105141f $X=6.295 $Y=0.85
+ $X2=0 $Y2=0
cc_409 N_A_885_297#_c_406_n N_A_453_325#_c_998_n 0.00264545f $X=6.15 $Y=0.85
+ $X2=0 $Y2=0
cc_410 N_A_885_297#_c_412_n N_A_453_325#_c_1008_n 0.00258134f $X=6.34 $Y=1.41
+ $X2=0 $Y2=0
cc_411 N_A_885_297#_c_414_n N_A_453_325#_c_1008_n 0.00822576f $X=7.83 $Y=1.57
+ $X2=0 $Y2=0
cc_412 N_A_885_297#_M1001_g N_A_453_325#_c_1046_n 0.00223132f $X=6.365 $Y=0.455
+ $X2=0 $Y2=0
cc_413 N_A_885_297#_c_406_n N_A_453_325#_c_1046_n 0.00180873f $X=6.15 $Y=0.85
+ $X2=0 $Y2=0
cc_414 N_A_885_297#_c_411_n N_A_453_325#_c_999_n 0.00616338f $X=4.79 $Y=0.74
+ $X2=0 $Y2=0
cc_415 N_A_885_297#_c_400_n N_A_453_325#_c_1000_n 2.22283e-19 $X=6.24 $Y=1.16
+ $X2=0 $Y2=0
cc_416 N_A_885_297#_c_402_n N_A_453_325#_c_1000_n 0.00299453f $X=6.13 $Y=0.995
+ $X2=0 $Y2=0
cc_417 N_A_885_297#_c_403_n N_A_453_325#_c_1000_n 0.0171949f $X=6.005 $Y=0.85
+ $X2=0 $Y2=0
cc_418 N_A_885_297#_c_405_n N_A_453_325#_c_1000_n 0.00134696f $X=6.295 $Y=0.85
+ $X2=0 $Y2=0
cc_419 N_A_885_297#_c_406_n N_A_453_325#_c_1000_n 0.0141636f $X=6.15 $Y=0.85
+ $X2=0 $Y2=0
cc_420 N_A_885_297#_c_404_n N_A_477_49#_M1004_d 0.00140408f $X=7.485 $Y=0.85
+ $X2=0 $Y2=0
cc_421 N_A_885_297#_c_407_n N_A_477_49#_M1004_d 0.00214439f $X=7.63 $Y=0.85
+ $X2=0 $Y2=0
cc_422 N_A_885_297#_c_408_n N_A_477_49#_M1004_d 0.0050343f $X=7.63 $Y=0.85 $X2=0
+ $Y2=0
cc_423 N_A_885_297#_c_400_n N_A_477_49#_c_1154_n 0.00881942f $X=6.24 $Y=1.16
+ $X2=0 $Y2=0
cc_424 N_A_885_297#_c_402_n N_A_477_49#_c_1154_n 0.0271004f $X=6.13 $Y=0.995
+ $X2=0 $Y2=0
cc_425 N_A_885_297#_c_403_n N_A_477_49#_c_1154_n 5.63647e-19 $X=6.005 $Y=0.85
+ $X2=0 $Y2=0
cc_426 N_A_885_297#_c_412_n N_A_477_49#_c_1191_n 0.00383389f $X=6.34 $Y=1.41
+ $X2=0 $Y2=0
cc_427 N_A_885_297#_c_412_n N_A_477_49#_c_1155_n 0.0169561f $X=6.34 $Y=1.41
+ $X2=0 $Y2=0
cc_428 N_A_885_297#_c_400_n N_A_477_49#_c_1155_n 7.42472e-19 $X=6.24 $Y=1.16
+ $X2=0 $Y2=0
cc_429 N_A_885_297#_c_401_n N_A_477_49#_c_1155_n 9.0109e-19 $X=6.34 $Y=1.202
+ $X2=0 $Y2=0
cc_430 N_A_885_297#_c_402_n N_A_477_49#_c_1155_n 0.00152864f $X=6.13 $Y=0.995
+ $X2=0 $Y2=0
cc_431 N_A_885_297#_c_404_n N_A_477_49#_c_1155_n 0.00419686f $X=7.485 $Y=0.85
+ $X2=0 $Y2=0
cc_432 N_A_885_297#_c_405_n N_A_477_49#_c_1155_n 6.55203e-19 $X=6.295 $Y=0.85
+ $X2=0 $Y2=0
cc_433 N_A_885_297#_c_412_n N_A_477_49#_c_1151_n 0.00100752f $X=6.34 $Y=1.41
+ $X2=0 $Y2=0
cc_434 N_A_885_297#_M1001_g N_A_477_49#_c_1151_n 0.0154018f $X=6.365 $Y=0.455
+ $X2=0 $Y2=0
cc_435 N_A_885_297#_c_402_n N_A_477_49#_c_1151_n 0.0173003f $X=6.13 $Y=0.995
+ $X2=0 $Y2=0
cc_436 N_A_885_297#_c_404_n N_A_477_49#_c_1151_n 0.0173494f $X=7.485 $Y=0.85
+ $X2=0 $Y2=0
cc_437 N_A_885_297#_c_405_n N_A_477_49#_c_1151_n 0.00232583f $X=6.295 $Y=0.85
+ $X2=0 $Y2=0
cc_438 N_A_885_297#_c_406_n N_A_477_49#_c_1151_n 0.0185267f $X=6.15 $Y=0.85
+ $X2=0 $Y2=0
cc_439 N_A_885_297#_c_404_n N_A_477_49#_c_1204_n 0.00166303f $X=7.485 $Y=0.85
+ $X2=0 $Y2=0
cc_440 N_A_885_297#_c_407_n N_A_477_49#_c_1205_n 3.55136e-19 $X=7.63 $Y=0.85
+ $X2=0 $Y2=0
cc_441 N_A_885_297#_c_408_n N_A_477_49#_c_1205_n 0.00528249f $X=7.63 $Y=0.85
+ $X2=0 $Y2=0
cc_442 N_A_885_297#_c_410_n N_A_477_49#_c_1205_n 0.00335197f $X=7.772 $Y=0.945
+ $X2=0 $Y2=0
cc_443 N_A_885_297#_c_417_n N_A_477_49#_c_1157_n 0.0275977f $X=4.73 $Y=1.58
+ $X2=0 $Y2=0
cc_444 N_A_885_297#_c_402_n N_A_477_49#_c_1157_n 8.40027e-19 $X=6.13 $Y=0.995
+ $X2=0 $Y2=0
cc_445 N_A_885_297#_c_403_n N_A_477_49#_c_1157_n 0.0525103f $X=6.005 $Y=0.85
+ $X2=0 $Y2=0
cc_446 N_A_885_297#_c_421_p N_A_477_49#_c_1157_n 0.0124731f $X=4.815 $Y=0.85
+ $X2=0 $Y2=0
cc_447 N_A_885_297#_c_411_n N_A_477_49#_c_1157_n 0.00234688f $X=4.79 $Y=0.74
+ $X2=0 $Y2=0
cc_448 N_A_885_297#_c_412_n N_A_477_49#_c_1160_n 0.00348376f $X=6.34 $Y=1.41
+ $X2=0 $Y2=0
cc_449 N_A_885_297#_c_400_n N_A_477_49#_c_1160_n 0.00431105f $X=6.24 $Y=1.16
+ $X2=0 $Y2=0
cc_450 N_A_885_297#_c_401_n N_A_477_49#_c_1160_n 2.0806e-19 $X=6.34 $Y=1.202
+ $X2=0 $Y2=0
cc_451 N_A_885_297#_c_402_n N_A_477_49#_c_1160_n 0.00243787f $X=6.13 $Y=0.995
+ $X2=0 $Y2=0
cc_452 N_A_885_297#_c_405_n N_A_477_49#_c_1160_n 0.015476f $X=6.295 $Y=0.85
+ $X2=0 $Y2=0
cc_453 N_A_885_297#_c_404_n N_A_1286_297#_M1001_d 0.00166227f $X=7.485 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_454 N_A_885_297#_c_412_n N_A_1286_297#_c_1286_n 0.00357027f $X=6.34 $Y=1.41
+ $X2=0 $Y2=0
cc_455 N_A_885_297#_c_404_n N_A_1286_297#_c_1286_n 0.0181022f $X=7.485 $Y=0.85
+ $X2=0 $Y2=0
cc_456 N_A_885_297#_c_407_n N_A_1286_297#_c_1286_n 0.0020738f $X=7.63 $Y=0.85
+ $X2=0 $Y2=0
cc_457 N_A_885_297#_c_408_n N_A_1286_297#_c_1286_n 0.00517339f $X=7.63 $Y=0.85
+ $X2=0 $Y2=0
cc_458 N_A_885_297#_c_412_n N_A_1286_297#_c_1298_n 0.0027417f $X=6.34 $Y=1.41
+ $X2=0 $Y2=0
cc_459 N_A_885_297#_c_414_n N_A_1286_297#_c_1299_n 0.0168297f $X=7.83 $Y=1.57
+ $X2=0 $Y2=0
cc_460 N_A_885_297#_c_408_n N_A_1286_297#_c_1299_n 0.00161448f $X=7.63 $Y=0.85
+ $X2=0 $Y2=0
cc_461 N_A_885_297#_c_421_p N_VGND_c_1356_n 0.00371415f $X=4.815 $Y=0.85 $X2=0
+ $Y2=0
cc_462 N_A_885_297#_c_411_n N_VGND_c_1356_n 0.0242428f $X=4.79 $Y=0.74 $X2=0
+ $Y2=0
cc_463 N_A_885_297#_M1001_g N_VGND_c_1360_n 0.00575161f $X=6.365 $Y=0.455 $X2=0
+ $Y2=0
cc_464 N_A_885_297#_c_406_n N_VGND_c_1360_n 0.00340751f $X=6.15 $Y=0.85 $X2=0
+ $Y2=0
cc_465 N_A_885_297#_c_408_n N_VGND_c_1360_n 0.00102193f $X=7.63 $Y=0.85 $X2=0
+ $Y2=0
cc_466 N_A_885_297#_c_410_n N_VGND_c_1360_n 0.00585385f $X=7.772 $Y=0.945 $X2=0
+ $Y2=0
cc_467 N_A_885_297#_c_411_n N_VGND_c_1360_n 0.0088551f $X=4.79 $Y=0.74 $X2=0
+ $Y2=0
cc_468 N_A_885_297#_M1022_d N_VGND_c_1364_n 0.00198811f $X=4.655 $Y=0.235 $X2=0
+ $Y2=0
cc_469 N_A_885_297#_M1001_g N_VGND_c_1364_n 0.00668858f $X=6.365 $Y=0.455 $X2=0
+ $Y2=0
cc_470 N_A_885_297#_c_403_n N_VGND_c_1364_n 0.0112598f $X=6.005 $Y=0.85 $X2=0
+ $Y2=0
cc_471 N_A_885_297#_c_421_p N_VGND_c_1364_n 0.0148172f $X=4.815 $Y=0.85 $X2=0
+ $Y2=0
cc_472 N_A_885_297#_c_410_n N_VGND_c_1364_n 0.00635691f $X=7.772 $Y=0.945 $X2=0
+ $Y2=0
cc_473 N_A_885_297#_c_411_n N_VGND_c_1364_n 0.00448669f $X=4.79 $Y=0.74 $X2=0
+ $Y2=0
cc_474 N_B_c_589_n N_A_1003_297#_c_754_n 0.003607f $X=4.335 $Y=1.41 $X2=0 $Y2=0
cc_475 N_B_M1022_g N_A_1003_297#_c_754_n 0.00120589f $X=4.58 $Y=0.56 $X2=0 $Y2=0
cc_476 N_B_c_582_n N_A_1003_297#_c_754_n 0.014573f $X=5.435 $Y=1.16 $X2=0 $Y2=0
cc_477 N_B_M1010_g N_A_1003_297#_c_754_n 0.00424996f $X=5.535 $Y=1.905 $X2=0
+ $Y2=0
cc_478 N_B_M1015_g N_A_1003_297#_c_754_n 0.0035466f $X=5.56 $Y=0.565 $X2=0 $Y2=0
cc_479 N_B_c_585_n N_A_1003_297#_c_754_n 0.0011146f $X=5.535 $Y=1.16 $X2=0 $Y2=0
cc_480 B N_A_1003_297#_c_762_n 0.008575f $X=7.5 $Y=1.445 $X2=0 $Y2=0
cc_481 N_B_M1015_g N_A_1003_297#_c_774_n 0.00201366f $X=5.56 $Y=0.565 $X2=0
+ $Y2=0
cc_482 N_B_c_588_n N_A_1003_297#_c_774_n 0.0032563f $X=7.245 $Y=0.995 $X2=0
+ $Y2=0
cc_483 N_B_M1022_g N_A_1003_297#_c_758_n 4.212e-19 $X=4.58 $Y=0.56 $X2=0 $Y2=0
cc_484 N_B_M1015_g N_A_1003_297#_c_758_n 9.17075e-19 $X=5.56 $Y=0.565 $X2=0
+ $Y2=0
cc_485 N_B_M1022_g N_A_1003_297#_c_759_n 0.00491597f $X=4.58 $Y=0.56 $X2=0 $Y2=0
cc_486 N_B_c_582_n N_A_1003_297#_c_759_n 0.00309496f $X=5.435 $Y=1.16 $X2=0
+ $Y2=0
cc_487 N_B_c_589_n N_VPWR_c_888_n 0.0113699f $X=4.335 $Y=1.41 $X2=0 $Y2=0
cc_488 N_B_c_589_n N_VPWR_c_893_n 0.00455828f $X=4.335 $Y=1.41 $X2=0 $Y2=0
cc_489 N_B_c_593_n N_VPWR_c_893_n 0.0390761f $X=5.635 $Y=2.54 $X2=0 $Y2=0
cc_490 N_B_c_589_n N_VPWR_c_884_n 0.00656627f $X=4.335 $Y=1.41 $X2=0 $Y2=0
cc_491 N_B_c_592_n N_VPWR_c_884_n 0.0395171f $X=7.085 $Y=2.54 $X2=0 $Y2=0
cc_492 N_B_c_593_n N_VPWR_c_884_n 0.0071208f $X=5.635 $Y=2.54 $X2=0 $Y2=0
cc_493 N_B_M1022_g N_A_453_325#_c_996_n 0.00316063f $X=4.58 $Y=0.56 $X2=0 $Y2=0
cc_494 N_B_c_589_n N_A_453_325#_c_997_n 0.0127882f $X=4.335 $Y=1.41 $X2=0 $Y2=0
cc_495 N_B_c_583_n N_A_453_325#_c_997_n 0.00535881f $X=4.655 $Y=1.16 $X2=0 $Y2=0
cc_496 N_B_c_589_n N_A_453_325#_c_1003_n 0.0175458f $X=4.335 $Y=1.41 $X2=0 $Y2=0
cc_497 N_B_c_589_n N_A_453_325#_c_1004_n 0.00608631f $X=4.335 $Y=1.41 $X2=0
+ $Y2=0
cc_498 N_B_M1010_g N_A_453_325#_c_1004_n 8.94333e-19 $X=5.535 $Y=1.905 $X2=0
+ $Y2=0
cc_499 N_B_c_589_n N_A_453_325#_c_1006_n 0.00366198f $X=4.335 $Y=1.41 $X2=0
+ $Y2=0
cc_500 N_B_c_582_n N_A_453_325#_c_998_n 0.00354518f $X=5.435 $Y=1.16 $X2=0 $Y2=0
cc_501 N_B_M1010_g N_A_453_325#_c_998_n 0.0315935f $X=5.535 $Y=1.905 $X2=0 $Y2=0
cc_502 N_B_M1015_g N_A_453_325#_c_998_n 0.00651676f $X=5.56 $Y=0.565 $X2=0 $Y2=0
cc_503 N_B_c_585_n N_A_453_325#_c_998_n 0.0105369f $X=5.535 $Y=1.16 $X2=0 $Y2=0
cc_504 N_B_M1010_g N_A_453_325#_c_1008_n 0.00817171f $X=5.535 $Y=1.905 $X2=0
+ $Y2=0
cc_505 N_B_c_592_n N_A_453_325#_c_1008_n 0.0346605f $X=7.085 $Y=2.54 $X2=0 $Y2=0
cc_506 N_B_c_593_n N_A_453_325#_c_1008_n 2.38151e-19 $X=5.635 $Y=2.54 $X2=0
+ $Y2=0
cc_507 N_B_M1006_g N_A_453_325#_c_1008_n 0.0104749f $X=7.185 $Y=1.965 $X2=0
+ $Y2=0
cc_508 N_B_M1015_g N_A_453_325#_c_1046_n 5.73691e-19 $X=5.56 $Y=0.565 $X2=0
+ $Y2=0
cc_509 N_B_M1022_g N_A_453_325#_c_999_n 8.48623e-19 $X=4.58 $Y=0.56 $X2=0 $Y2=0
cc_510 N_B_c_583_n N_A_453_325#_c_999_n 0.0038653f $X=4.655 $Y=1.16 $X2=0 $Y2=0
cc_511 N_B_M1015_g N_A_453_325#_c_1000_n 0.0136729f $X=5.56 $Y=0.565 $X2=0 $Y2=0
cc_512 N_B_M1010_g N_A_453_325#_c_1010_n 0.00716396f $X=5.535 $Y=1.905 $X2=0
+ $Y2=0
cc_513 N_B_c_593_n N_A_453_325#_c_1010_n 2.51585e-19 $X=5.635 $Y=2.54 $X2=0
+ $Y2=0
cc_514 N_B_c_583_n N_A_477_49#_c_1150_n 4.44674e-19 $X=4.655 $Y=1.16 $X2=0 $Y2=0
cc_515 N_B_M1010_g N_A_477_49#_c_1154_n 0.00145677f $X=5.535 $Y=1.905 $X2=0
+ $Y2=0
cc_516 N_B_M1010_g N_A_477_49#_c_1191_n 0.00446449f $X=5.535 $Y=1.905 $X2=0
+ $Y2=0
cc_517 N_B_c_588_n N_A_477_49#_c_1151_n 0.00275402f $X=7.245 $Y=0.995 $X2=0
+ $Y2=0
cc_518 N_B_c_586_n N_A_477_49#_c_1204_n 0.0029291f $X=7.22 $Y=1.16 $X2=0 $Y2=0
cc_519 N_B_c_587_n N_A_477_49#_c_1204_n 4.33224e-19 $X=7.22 $Y=1.16 $X2=0 $Y2=0
cc_520 N_B_c_588_n N_A_477_49#_c_1204_n 0.00498906f $X=7.245 $Y=0.995 $X2=0
+ $Y2=0
cc_521 N_B_c_587_n N_A_477_49#_c_1205_n 0.00108686f $X=7.22 $Y=1.16 $X2=0 $Y2=0
cc_522 N_B_c_588_n N_A_477_49#_c_1226_n 0.00521263f $X=7.245 $Y=0.995 $X2=0
+ $Y2=0
cc_523 N_B_c_589_n N_A_477_49#_c_1157_n 0.00469456f $X=4.335 $Y=1.41 $X2=0 $Y2=0
cc_524 N_B_c_582_n N_A_477_49#_c_1157_n 0.00486395f $X=5.435 $Y=1.16 $X2=0 $Y2=0
cc_525 N_B_c_583_n N_A_477_49#_c_1157_n 2.58451e-19 $X=4.655 $Y=1.16 $X2=0 $Y2=0
cc_526 N_B_M1010_g N_A_477_49#_c_1157_n 0.00481446f $X=5.535 $Y=1.905 $X2=0
+ $Y2=0
cc_527 N_B_c_585_n N_A_477_49#_c_1157_n 2.29578e-19 $X=5.535 $Y=1.16 $X2=0 $Y2=0
cc_528 N_B_M1010_g N_A_477_49#_c_1160_n 4.48588e-19 $X=5.535 $Y=1.905 $X2=0
+ $Y2=0
cc_529 N_B_M1006_g N_A_1286_297#_c_1286_n 0.00869344f $X=7.185 $Y=1.965 $X2=0
+ $Y2=0
cc_530 N_B_c_586_n N_A_1286_297#_c_1286_n 0.03273f $X=7.22 $Y=1.16 $X2=0 $Y2=0
cc_531 N_B_c_600_n N_A_1286_297#_c_1286_n 0.0134199f $X=7.355 $Y=1.53 $X2=0
+ $Y2=0
cc_532 N_B_c_588_n N_A_1286_297#_c_1286_n 0.0130696f $X=7.245 $Y=0.995 $X2=0
+ $Y2=0
cc_533 N_B_M1006_g N_A_1286_297#_c_1299_n 0.0153655f $X=7.185 $Y=1.965 $X2=0
+ $Y2=0
cc_534 N_B_c_587_n N_A_1286_297#_c_1299_n 2.73792e-19 $X=7.22 $Y=1.16 $X2=0
+ $Y2=0
cc_535 N_B_c_600_n N_A_1286_297#_c_1299_n 0.00926119f $X=7.355 $Y=1.53 $X2=0
+ $Y2=0
cc_536 B N_A_1286_297#_c_1299_n 0.0178346f $X=7.5 $Y=1.445 $X2=0 $Y2=0
cc_537 N_B_M1022_g N_VGND_c_1356_n 0.0190364f $X=4.58 $Y=0.56 $X2=0 $Y2=0
cc_538 N_B_c_583_n N_VGND_c_1356_n 0.00541821f $X=4.655 $Y=1.16 $X2=0 $Y2=0
cc_539 N_B_M1022_g N_VGND_c_1360_n 0.00494995f $X=4.58 $Y=0.56 $X2=0 $Y2=0
cc_540 N_B_M1015_g N_VGND_c_1360_n 0.00427876f $X=5.56 $Y=0.565 $X2=0 $Y2=0
cc_541 N_B_c_588_n N_VGND_c_1360_n 0.00357877f $X=7.245 $Y=0.995 $X2=0 $Y2=0
cc_542 N_B_M1022_g N_VGND_c_1364_n 0.00918586f $X=4.58 $Y=0.56 $X2=0 $Y2=0
cc_543 N_B_M1015_g N_VGND_c_1364_n 0.00718354f $X=5.56 $Y=0.565 $X2=0 $Y2=0
cc_544 N_B_c_588_n N_VGND_c_1364_n 0.00612424f $X=7.245 $Y=0.995 $X2=0 $Y2=0
cc_545 N_A_c_718_n N_A_1003_297#_c_752_n 0.0228311f $X=8.41 $Y=0.995 $X2=0 $Y2=0
cc_546 N_A_c_717_n N_A_1003_297#_c_753_n 0.0630265f $X=8.385 $Y=1.41 $X2=0 $Y2=0
cc_547 A N_A_1003_297#_c_753_n 0.00219839f $X=8.43 $Y=1.105 $X2=0 $Y2=0
cc_548 N_A_c_717_n N_A_1003_297#_c_762_n 0.0144336f $X=8.385 $Y=1.41 $X2=0 $Y2=0
cc_549 A N_A_1003_297#_c_762_n 0.0434391f $X=8.43 $Y=1.105 $X2=0 $Y2=0
cc_550 N_A_c_717_n N_A_1003_297#_c_755_n 5.76324e-19 $X=8.385 $Y=1.41 $X2=0
+ $Y2=0
cc_551 N_A_c_718_n N_A_1003_297#_c_755_n 0.0111816f $X=8.41 $Y=0.995 $X2=0 $Y2=0
cc_552 A N_A_1003_297#_c_755_n 0.0282016f $X=8.43 $Y=1.105 $X2=0 $Y2=0
cc_553 N_A_c_717_n N_A_1003_297#_c_756_n 0.00444032f $X=8.385 $Y=1.41 $X2=0
+ $Y2=0
cc_554 A N_A_1003_297#_c_756_n 0.0205785f $X=8.43 $Y=1.105 $X2=0 $Y2=0
cc_555 N_A_c_718_n N_A_1003_297#_c_757_n 8.99731e-19 $X=8.41 $Y=0.995 $X2=0
+ $Y2=0
cc_556 A N_A_1003_297#_c_757_n 0.0206762f $X=8.43 $Y=1.105 $X2=0 $Y2=0
cc_557 N_A_c_717_n N_A_1003_297#_c_764_n 8.78751e-19 $X=8.385 $Y=1.41 $X2=0
+ $Y2=0
cc_558 A N_A_1003_297#_c_787_n 9.51454e-19 $X=8.43 $Y=1.105 $X2=0 $Y2=0
cc_559 N_A_c_717_n N_VPWR_c_889_n 0.00866059f $X=8.385 $Y=1.41 $X2=0 $Y2=0
cc_560 N_A_c_717_n N_VPWR_c_893_n 0.00449565f $X=8.385 $Y=1.41 $X2=0 $Y2=0
cc_561 N_A_c_717_n N_VPWR_c_884_n 0.00535272f $X=8.385 $Y=1.41 $X2=0 $Y2=0
cc_562 N_A_c_717_n N_A_453_325#_c_1008_n 0.00156782f $X=8.385 $Y=1.41 $X2=0
+ $Y2=0
cc_563 N_A_c_717_n N_A_1286_297#_c_1299_n 0.0140513f $X=8.385 $Y=1.41 $X2=0
+ $Y2=0
cc_564 N_A_c_718_n N_VGND_c_1357_n 0.00268723f $X=8.41 $Y=0.995 $X2=0 $Y2=0
cc_565 N_A_c_718_n N_VGND_c_1360_n 0.00439206f $X=8.41 $Y=0.995 $X2=0 $Y2=0
cc_566 N_A_c_718_n N_VGND_c_1364_n 0.00631885f $X=8.41 $Y=0.995 $X2=0 $Y2=0
cc_567 N_A_1003_297#_c_762_n N_VPWR_M1018_d 0.00414509f $X=8.865 $Y=1.6 $X2=0
+ $Y2=0
cc_568 N_A_1003_297#_c_753_n N_VPWR_c_889_n 0.00922704f $X=8.855 $Y=1.41 $X2=0
+ $Y2=0
cc_569 N_A_1003_297#_c_753_n N_VPWR_c_894_n 0.00435494f $X=8.855 $Y=1.41 $X2=0
+ $Y2=0
cc_570 N_A_1003_297#_M1014_d N_VPWR_c_884_n 0.00402227f $X=7.92 $Y=1.645 $X2=0
+ $Y2=0
cc_571 N_A_1003_297#_c_753_n N_VPWR_c_884_n 0.00613107f $X=8.855 $Y=1.41 $X2=0
+ $Y2=0
cc_572 N_A_1003_297#_c_774_n N_A_453_325#_M1015_d 0.00599198f $X=7.995 $Y=0.51
+ $X2=0 $Y2=0
cc_573 N_A_1003_297#_c_754_n N_A_453_325#_c_1003_n 0.0132911f $X=5.14 $Y=1.94
+ $X2=0 $Y2=0
cc_574 N_A_1003_297#_c_754_n N_A_453_325#_c_1004_n 0.00274773f $X=5.14 $Y=1.94
+ $X2=0 $Y2=0
cc_575 N_A_1003_297#_M1010_s N_A_453_325#_c_1005_n 0.0102858f $X=5.015 $Y=1.485
+ $X2=0 $Y2=0
cc_576 N_A_1003_297#_c_754_n N_A_453_325#_c_1005_n 0.0128549f $X=5.14 $Y=1.94
+ $X2=0 $Y2=0
cc_577 N_A_1003_297#_c_754_n N_A_453_325#_c_998_n 0.0675972f $X=5.14 $Y=1.94
+ $X2=0 $Y2=0
cc_578 N_A_1003_297#_M1014_d N_A_453_325#_c_1008_n 0.00273002f $X=7.92 $Y=1.645
+ $X2=0 $Y2=0
cc_579 N_A_1003_297#_c_774_n N_A_453_325#_c_1046_n 0.0125715f $X=7.995 $Y=0.51
+ $X2=0 $Y2=0
cc_580 N_A_1003_297#_c_758_n N_A_453_325#_c_1046_n 0.0014251f $X=5.325 $Y=0.51
+ $X2=0 $Y2=0
cc_581 N_A_1003_297#_c_759_n N_A_453_325#_c_1046_n 0.00331722f $X=5.18 $Y=0.51
+ $X2=0 $Y2=0
cc_582 N_A_1003_297#_M1015_s N_A_453_325#_c_1000_n 0.00152093f $X=5.175 $Y=0.245
+ $X2=0 $Y2=0
cc_583 N_A_1003_297#_c_754_n N_A_453_325#_c_1000_n 0.0123119f $X=5.14 $Y=1.94
+ $X2=0 $Y2=0
cc_584 N_A_1003_297#_c_774_n N_A_453_325#_c_1000_n 0.00366657f $X=7.995 $Y=0.51
+ $X2=0 $Y2=0
cc_585 N_A_1003_297#_c_759_n N_A_453_325#_c_1000_n 0.00172491f $X=5.18 $Y=0.51
+ $X2=0 $Y2=0
cc_586 N_A_1003_297#_c_774_n N_A_477_49#_M1004_d 0.00419658f $X=7.995 $Y=0.51
+ $X2=0 $Y2=0
cc_587 N_A_1003_297#_c_774_n N_A_477_49#_c_1151_n 0.0147234f $X=7.995 $Y=0.51
+ $X2=0 $Y2=0
cc_588 N_A_1003_297#_c_774_n N_A_477_49#_c_1204_n 0.00610486f $X=7.995 $Y=0.51
+ $X2=0 $Y2=0
cc_589 N_A_1003_297#_c_774_n N_A_477_49#_c_1205_n 0.00980954f $X=7.995 $Y=0.51
+ $X2=0 $Y2=0
cc_590 N_A_1003_297#_c_787_n N_A_477_49#_c_1205_n 0.0012274f $X=8.14 $Y=0.51
+ $X2=0 $Y2=0
cc_591 N_A_1003_297#_c_788_n N_A_477_49#_c_1205_n 0.00676871f $X=8.14 $Y=0.51
+ $X2=0 $Y2=0
cc_592 N_A_1003_297#_c_774_n N_A_477_49#_c_1226_n 0.0119237f $X=7.995 $Y=0.51
+ $X2=0 $Y2=0
cc_593 N_A_1003_297#_M1010_s N_A_477_49#_c_1157_n 0.00802537f $X=5.015 $Y=1.485
+ $X2=0 $Y2=0
cc_594 N_A_1003_297#_c_754_n N_A_477_49#_c_1157_n 0.0183124f $X=5.14 $Y=1.94
+ $X2=0 $Y2=0
cc_595 N_A_1003_297#_c_774_n N_A_1286_297#_M1001_d 0.00653094f $X=7.995 $Y=0.51
+ $X2=-0.19 $Y2=-0.24
cc_596 N_A_1003_297#_c_757_n N_A_1286_297#_M1020_d 0.00343897f $X=8.95 $Y=1.325
+ $X2=0 $Y2=0
cc_597 N_A_1003_297#_c_762_n N_A_1286_297#_M1011_d 0.00328472f $X=8.865 $Y=1.6
+ $X2=0 $Y2=0
cc_598 N_A_1003_297#_c_774_n N_A_1286_297#_c_1286_n 0.00162336f $X=7.995 $Y=0.51
+ $X2=0 $Y2=0
cc_599 N_A_1003_297#_c_753_n N_A_1286_297#_c_1290_n 0.00981878f $X=8.855 $Y=1.41
+ $X2=0 $Y2=0
cc_600 N_A_1003_297#_c_752_n N_A_1286_297#_c_1287_n 0.0052678f $X=8.83 $Y=0.995
+ $X2=0 $Y2=0
cc_601 N_A_1003_297#_c_753_n N_A_1286_297#_c_1287_n 0.0151795f $X=8.855 $Y=1.41
+ $X2=0 $Y2=0
cc_602 N_A_1003_297#_c_762_n N_A_1286_297#_c_1287_n 0.0118142f $X=8.865 $Y=1.6
+ $X2=0 $Y2=0
cc_603 N_A_1003_297#_c_757_n N_A_1286_297#_c_1287_n 0.0390874f $X=8.95 $Y=1.325
+ $X2=0 $Y2=0
cc_604 N_A_1003_297#_c_764_n N_A_1286_297#_c_1287_n 0.00896957f $X=8.95 $Y=1.495
+ $X2=0 $Y2=0
cc_605 N_A_1003_297#_M1014_d N_A_1286_297#_c_1299_n 0.00774465f $X=7.92 $Y=1.645
+ $X2=0 $Y2=0
cc_606 N_A_1003_297#_c_753_n N_A_1286_297#_c_1299_n 0.0153391f $X=8.855 $Y=1.41
+ $X2=0 $Y2=0
cc_607 N_A_1003_297#_c_762_n N_A_1286_297#_c_1299_n 0.0451449f $X=8.865 $Y=1.6
+ $X2=0 $Y2=0
cc_608 N_A_1003_297#_c_753_n N_A_1286_297#_c_1292_n 0.00211441f $X=8.855 $Y=1.41
+ $X2=0 $Y2=0
cc_609 N_A_1003_297#_c_762_n N_A_1286_297#_c_1292_n 0.00269572f $X=8.865 $Y=1.6
+ $X2=0 $Y2=0
cc_610 N_A_1003_297#_c_757_n N_A_1286_297#_c_1292_n 0.00332545f $X=8.95 $Y=1.325
+ $X2=0 $Y2=0
cc_611 N_A_1003_297#_c_752_n N_A_1286_297#_c_1288_n 0.00684238f $X=8.83 $Y=0.995
+ $X2=0 $Y2=0
cc_612 N_A_1003_297#_c_753_n N_A_1286_297#_c_1288_n 3.13625e-19 $X=8.855 $Y=1.41
+ $X2=0 $Y2=0
cc_613 N_A_1003_297#_c_755_n N_VGND_M1021_d 0.00162006f $X=8.865 $Y=0.82 $X2=0
+ $Y2=0
cc_614 N_A_1003_297#_c_752_n N_VGND_c_1357_n 0.00268723f $X=8.83 $Y=0.995 $X2=0
+ $Y2=0
cc_615 N_A_1003_297#_c_755_n N_VGND_c_1357_n 0.0122414f $X=8.865 $Y=0.82 $X2=0
+ $Y2=0
cc_616 N_A_1003_297#_c_787_n N_VGND_c_1357_n 0.00112928f $X=8.14 $Y=0.51 $X2=0
+ $Y2=0
cc_617 N_A_1003_297#_c_755_n N_VGND_c_1360_n 0.00248202f $X=8.865 $Y=0.82 $X2=0
+ $Y2=0
cc_618 N_A_1003_297#_c_774_n N_VGND_c_1360_n 0.00574592f $X=7.995 $Y=0.51 $X2=0
+ $Y2=0
cc_619 N_A_1003_297#_c_758_n N_VGND_c_1360_n 2.9688e-19 $X=5.325 $Y=0.51 $X2=0
+ $Y2=0
cc_620 N_A_1003_297#_c_759_n N_VGND_c_1360_n 0.0250994f $X=5.18 $Y=0.51 $X2=0
+ $Y2=0
cc_621 N_A_1003_297#_c_787_n N_VGND_c_1360_n 3.63685e-19 $X=8.14 $Y=0.51 $X2=0
+ $Y2=0
cc_622 N_A_1003_297#_c_788_n N_VGND_c_1360_n 0.0149689f $X=8.14 $Y=0.51 $X2=0
+ $Y2=0
cc_623 N_A_1003_297#_c_752_n N_VGND_c_1363_n 0.0043917f $X=8.83 $Y=0.995 $X2=0
+ $Y2=0
cc_624 N_A_1003_297#_c_755_n N_VGND_c_1363_n 0.00180657f $X=8.865 $Y=0.82 $X2=0
+ $Y2=0
cc_625 N_A_1003_297#_c_757_n N_VGND_c_1363_n 0.00215988f $X=8.95 $Y=1.325 $X2=0
+ $Y2=0
cc_626 N_A_1003_297#_M1012_d N_VGND_c_1364_n 0.00244776f $X=7.93 $Y=0.235 $X2=0
+ $Y2=0
cc_627 N_A_1003_297#_c_752_n N_VGND_c_1364_n 0.00735952f $X=8.83 $Y=0.995 $X2=0
+ $Y2=0
cc_628 N_A_1003_297#_c_755_n N_VGND_c_1364_n 0.00919596f $X=8.865 $Y=0.82 $X2=0
+ $Y2=0
cc_629 N_A_1003_297#_c_757_n N_VGND_c_1364_n 0.00454532f $X=8.95 $Y=1.325 $X2=0
+ $Y2=0
cc_630 N_A_1003_297#_c_774_n N_VGND_c_1364_n 0.232931f $X=7.995 $Y=0.51 $X2=0
+ $Y2=0
cc_631 N_A_1003_297#_c_758_n N_VGND_c_1364_n 0.028616f $X=5.325 $Y=0.51 $X2=0
+ $Y2=0
cc_632 N_A_1003_297#_c_759_n N_VGND_c_1364_n 0.00392171f $X=5.18 $Y=0.51 $X2=0
+ $Y2=0
cc_633 N_A_1003_297#_c_787_n N_VGND_c_1364_n 0.0285254f $X=8.14 $Y=0.51 $X2=0
+ $Y2=0
cc_634 N_A_1003_297#_c_788_n N_VGND_c_1364_n 0.0036194f $X=8.14 $Y=0.51 $X2=0
+ $Y2=0
cc_635 N_VPWR_c_884_n N_X_M1013_d 0.00351468f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_636 N_VPWR_c_892_n N_X_c_981_n 0.0193541f $X=1.045 $Y=2.72 $X2=0 $Y2=0
cc_637 N_VPWR_c_884_n N_X_c_981_n 0.0119959f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_638 N_VPWR_c_884_n N_A_453_325#_M1006_d 0.00242686f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_639 N_VPWR_c_888_n N_A_453_325#_c_1001_n 0.00147971f $X=4.1 $Y=2.32 $X2=0
+ $Y2=0
cc_640 N_VPWR_c_890_n N_A_453_325#_c_1001_n 0.012236f $X=3.935 $Y=2.72 $X2=0
+ $Y2=0
cc_641 N_VPWR_c_884_n N_A_453_325#_c_1001_n 0.0223233f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_642 N_VPWR_M1005_s N_A_453_325#_c_997_n 0.00648603f $X=3.975 $Y=2.175 $X2=0
+ $Y2=0
cc_643 N_VPWR_M1005_s N_A_453_325#_c_1003_n 0.00155527f $X=3.975 $Y=2.175 $X2=0
+ $Y2=0
cc_644 N_VPWR_c_888_n N_A_453_325#_c_1003_n 0.00612755f $X=4.1 $Y=2.32 $X2=0
+ $Y2=0
cc_645 N_VPWR_c_893_n N_A_453_325#_c_1003_n 0.00666556f $X=8.455 $Y=2.72 $X2=0
+ $Y2=0
cc_646 N_VPWR_c_884_n N_A_453_325#_c_1003_n 0.0119497f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_647 N_VPWR_c_888_n N_A_453_325#_c_1004_n 0.00140976f $X=4.1 $Y=2.32 $X2=0
+ $Y2=0
cc_648 N_VPWR_c_893_n N_A_453_325#_c_1005_n 0.0300226f $X=8.455 $Y=2.72 $X2=0
+ $Y2=0
cc_649 N_VPWR_c_884_n N_A_453_325#_c_1005_n 0.0193106f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_650 N_VPWR_c_888_n N_A_453_325#_c_1006_n 0.00679194f $X=4.1 $Y=2.32 $X2=0
+ $Y2=0
cc_651 N_VPWR_c_893_n N_A_453_325#_c_1006_n 0.0105925f $X=8.455 $Y=2.72 $X2=0
+ $Y2=0
cc_652 N_VPWR_c_884_n N_A_453_325#_c_1006_n 0.00644598f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_653 N_VPWR_c_889_n N_A_453_325#_c_1008_n 0.00642457f $X=8.62 $Y=2.36 $X2=0
+ $Y2=0
cc_654 N_VPWR_c_893_n N_A_453_325#_c_1008_n 0.134684f $X=8.455 $Y=2.72 $X2=0
+ $Y2=0
cc_655 N_VPWR_c_884_n N_A_453_325#_c_1008_n 0.0814374f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_656 N_VPWR_M1005_s N_A_453_325#_c_1009_n 0.00233831f $X=3.975 $Y=2.175 $X2=0
+ $Y2=0
cc_657 N_VPWR_c_888_n N_A_453_325#_c_1009_n 0.0144069f $X=4.1 $Y=2.32 $X2=0
+ $Y2=0
cc_658 N_VPWR_c_884_n N_A_453_325#_c_1009_n 8.22076e-19 $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_659 N_VPWR_c_893_n N_A_453_325#_c_1010_n 0.0103509f $X=8.455 $Y=2.72 $X2=0
+ $Y2=0
cc_660 N_VPWR_c_884_n N_A_453_325#_c_1010_n 0.00587789f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_661 N_VPWR_M1005_s N_A_477_49#_c_1157_n 0.00109947f $X=3.975 $Y=2.175 $X2=0
+ $Y2=0
cc_662 N_VPWR_c_884_n N_A_1286_297#_M1011_d 0.00469081f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_663 N_VPWR_c_889_n N_A_1286_297#_c_1290_n 0.00757454f $X=8.62 $Y=2.36 $X2=0
+ $Y2=0
cc_664 N_VPWR_c_894_n N_A_1286_297#_c_1290_n 0.0197624f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_665 N_VPWR_c_884_n N_A_1286_297#_c_1290_n 0.0111058f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_666 N_VPWR_M1018_d N_A_1286_297#_c_1299_n 0.00393477f $X=8.475 $Y=1.485 $X2=0
+ $Y2=0
cc_667 N_VPWR_c_889_n N_A_1286_297#_c_1299_n 0.0163118f $X=8.62 $Y=2.36 $X2=0
+ $Y2=0
cc_668 N_VPWR_c_893_n N_A_1286_297#_c_1299_n 0.00776959f $X=8.455 $Y=2.72 $X2=0
+ $Y2=0
cc_669 N_VPWR_c_894_n N_A_1286_297#_c_1299_n 0.00676887f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_670 N_VPWR_c_884_n N_A_1286_297#_c_1299_n 0.0268234f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_671 N_X_c_981_n N_VGND_c_1362_n 0.0125496f $X=0.75 $Y=0.56 $X2=0 $Y2=0
cc_672 N_X_M1002_s N_VGND_c_1364_n 0.00484781f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_673 N_X_c_981_n N_VGND_c_1364_n 0.0116366f $X=0.75 $Y=0.56 $X2=0 $Y2=0
cc_674 N_A_453_325#_c_1001_n N_A_477_49#_M1000_d 0.012215f $X=3.955 $Y=1.98
+ $X2=0 $Y2=0
cc_675 N_A_453_325#_c_1008_n N_A_477_49#_M1010_d 0.00924946f $X=7.585 $Y=2.36
+ $X2=0 $Y2=0
cc_676 N_A_453_325#_M1008_d N_A_477_49#_c_1162_n 0.0122835f $X=3.295 $Y=0.245
+ $X2=0 $Y2=0
cc_677 N_A_453_325#_c_995_n N_A_477_49#_c_1162_n 0.0212586f $X=3.845 $Y=0.37
+ $X2=0 $Y2=0
cc_678 N_A_453_325#_c_996_n N_A_477_49#_c_1162_n 0.0140572f $X=3.93 $Y=1.035
+ $X2=0 $Y2=0
cc_679 N_A_453_325#_M1008_d N_A_477_49#_c_1150_n 0.00280372f $X=3.295 $Y=0.245
+ $X2=0 $Y2=0
cc_680 N_A_453_325#_c_996_n N_A_477_49#_c_1150_n 0.0179158f $X=3.93 $Y=1.035
+ $X2=0 $Y2=0
cc_681 N_A_453_325#_c_997_n N_A_477_49#_c_1150_n 0.00902524f $X=4.04 $Y=1.895
+ $X2=0 $Y2=0
cc_682 N_A_453_325#_c_999_n N_A_477_49#_c_1150_n 0.0132103f $X=4.04 $Y=1.12
+ $X2=0 $Y2=0
cc_683 N_A_453_325#_c_998_n N_A_477_49#_c_1154_n 0.00870819f $X=5.48 $Y=2.275
+ $X2=0 $Y2=0
cc_684 N_A_453_325#_c_1000_n N_A_477_49#_c_1154_n 2.53366e-19 $X=5.48 $Y=0.772
+ $X2=0 $Y2=0
cc_685 N_A_453_325#_c_998_n N_A_477_49#_c_1191_n 0.0255541f $X=5.48 $Y=2.275
+ $X2=0 $Y2=0
cc_686 N_A_453_325#_c_1008_n N_A_477_49#_c_1191_n 0.0238103f $X=7.585 $Y=2.36
+ $X2=0 $Y2=0
cc_687 N_A_453_325#_c_1008_n N_A_477_49#_c_1155_n 0.0100462f $X=7.585 $Y=2.36
+ $X2=0 $Y2=0
cc_688 N_A_453_325#_c_1046_n N_A_477_49#_c_1151_n 0.00253431f $X=5.77 $Y=0.545
+ $X2=0 $Y2=0
cc_689 N_A_453_325#_c_1001_n N_A_477_49#_c_1157_n 0.00437461f $X=3.955 $Y=1.98
+ $X2=0 $Y2=0
cc_690 N_A_453_325#_c_997_n N_A_477_49#_c_1157_n 0.0161183f $X=4.04 $Y=1.895
+ $X2=0 $Y2=0
cc_691 N_A_453_325#_c_1003_n N_A_477_49#_c_1157_n 0.01149f $X=4.7 $Y=1.98 $X2=0
+ $Y2=0
cc_692 N_A_453_325#_c_998_n N_A_477_49#_c_1157_n 0.0194408f $X=5.48 $Y=2.275
+ $X2=0 $Y2=0
cc_693 N_A_453_325#_c_999_n N_A_477_49#_c_1157_n 0.0052436f $X=4.04 $Y=1.12
+ $X2=0 $Y2=0
cc_694 N_A_453_325#_c_1000_n N_A_477_49#_c_1157_n 8.86472e-19 $X=5.48 $Y=0.772
+ $X2=0 $Y2=0
cc_695 N_A_453_325#_c_1001_n N_A_477_49#_c_1158_n 0.00415423f $X=3.955 $Y=1.98
+ $X2=0 $Y2=0
cc_696 N_A_453_325#_c_997_n N_A_477_49#_c_1158_n 0.00275249f $X=4.04 $Y=1.895
+ $X2=0 $Y2=0
cc_697 N_A_453_325#_c_1001_n N_A_477_49#_c_1159_n 0.0251846f $X=3.955 $Y=1.98
+ $X2=0 $Y2=0
cc_698 N_A_453_325#_c_997_n N_A_477_49#_c_1159_n 0.0231767f $X=4.04 $Y=1.895
+ $X2=0 $Y2=0
cc_699 N_A_453_325#_c_998_n N_A_477_49#_c_1160_n 0.00127808f $X=5.48 $Y=2.275
+ $X2=0 $Y2=0
cc_700 N_A_453_325#_c_1008_n N_A_1286_297#_M1017_d 0.00474452f $X=7.585 $Y=2.36
+ $X2=0 $Y2=0
cc_701 N_A_453_325#_c_1008_n N_A_1286_297#_c_1298_n 0.0129278f $X=7.585 $Y=2.36
+ $X2=0 $Y2=0
cc_702 N_A_453_325#_M1006_d N_A_1286_297#_c_1299_n 0.00937242f $X=7.275 $Y=1.645
+ $X2=0 $Y2=0
cc_703 N_A_453_325#_c_1008_n N_A_1286_297#_c_1299_n 0.0533614f $X=7.585 $Y=2.36
+ $X2=0 $Y2=0
cc_704 N_A_453_325#_c_995_n N_VGND_c_1356_n 0.0140424f $X=3.845 $Y=0.37 $X2=0
+ $Y2=0
cc_705 N_A_453_325#_c_996_n N_VGND_c_1356_n 0.0299545f $X=3.93 $Y=1.035 $X2=0
+ $Y2=0
cc_706 N_A_453_325#_c_995_n N_VGND_c_1358_n 0.0348724f $X=3.845 $Y=0.37 $X2=0
+ $Y2=0
cc_707 N_A_453_325#_c_1046_n N_VGND_c_1360_n 0.00800682f $X=5.77 $Y=0.545 $X2=0
+ $Y2=0
cc_708 N_A_453_325#_c_1000_n N_VGND_c_1360_n 0.00283956f $X=5.48 $Y=0.772 $X2=0
+ $Y2=0
cc_709 N_A_453_325#_c_995_n N_VGND_c_1364_n 0.0232692f $X=3.845 $Y=0.37 $X2=0
+ $Y2=0
cc_710 N_A_453_325#_c_1046_n N_VGND_c_1364_n 0.0018012f $X=5.77 $Y=0.545 $X2=0
+ $Y2=0
cc_711 N_A_477_49#_c_1151_n N_A_1286_297#_M1001_d 0.00729398f $X=6.54 $Y=1.445
+ $X2=-0.19 $Y2=-0.24
cc_712 N_A_477_49#_c_1270_p N_A_1286_297#_M1001_d 0.0024562f $X=6.625 $Y=0.34
+ $X2=-0.19 $Y2=-0.24
cc_713 N_A_477_49#_c_1226_n N_A_1286_297#_M1001_d 0.0107136f $X=7.135 $Y=0.36
+ $X2=-0.19 $Y2=-0.24
cc_714 N_A_477_49#_c_1155_n N_A_1286_297#_M1017_d 0.00440874f $X=6.455 $Y=1.53
+ $X2=0 $Y2=0
cc_715 N_A_477_49#_c_1191_n N_A_1286_297#_c_1286_n 0.00453141f $X=5.97 $Y=1.62
+ $X2=0 $Y2=0
cc_716 N_A_477_49#_c_1155_n N_A_1286_297#_c_1286_n 0.013519f $X=6.455 $Y=1.53
+ $X2=0 $Y2=0
cc_717 N_A_477_49#_c_1151_n N_A_1286_297#_c_1286_n 0.0623179f $X=6.54 $Y=1.445
+ $X2=0 $Y2=0
cc_718 N_A_477_49#_c_1226_n N_A_1286_297#_c_1286_n 0.0106102f $X=7.135 $Y=0.36
+ $X2=0 $Y2=0
cc_719 N_A_477_49#_c_1160_n N_A_1286_297#_c_1286_n 0.00130235f $X=6.15 $Y=1.53
+ $X2=0 $Y2=0
cc_720 N_A_477_49#_c_1157_n N_VGND_c_1356_n 0.00557009f $X=6.005 $Y=1.53 $X2=0
+ $Y2=0
cc_721 N_A_477_49#_c_1162_n N_VGND_c_1358_n 0.00334078f $X=3.505 $Y=0.71 $X2=0
+ $Y2=0
cc_722 N_A_477_49#_c_1270_p N_VGND_c_1360_n 0.0104913f $X=6.625 $Y=0.34 $X2=0
+ $Y2=0
cc_723 N_A_477_49#_c_1226_n N_VGND_c_1360_n 0.0617902f $X=7.135 $Y=0.36 $X2=0
+ $Y2=0
cc_724 N_A_477_49#_M1004_d N_VGND_c_1364_n 0.00226821f $X=7.235 $Y=0.245 $X2=0
+ $Y2=0
cc_725 N_A_477_49#_c_1270_p N_VGND_c_1364_n 0.00184693f $X=6.625 $Y=0.34 $X2=0
+ $Y2=0
cc_726 N_A_477_49#_c_1152_n N_VGND_c_1364_n 0.00759655f $X=2.735 $Y=0.765 $X2=0
+ $Y2=0
cc_727 N_A_477_49#_c_1226_n N_VGND_c_1364_n 0.00974346f $X=7.135 $Y=0.36 $X2=0
+ $Y2=0
cc_728 N_A_1286_297#_c_1288_n N_VGND_c_1363_n 0.0199749f $X=9.4 $Y=0.42 $X2=0
+ $Y2=0
cc_729 N_A_1286_297#_M1020_d N_VGND_c_1364_n 0.010063f $X=8.905 $Y=0.235 $X2=0
+ $Y2=0
cc_730 N_A_1286_297#_c_1288_n N_VGND_c_1364_n 0.0113402f $X=9.4 $Y=0.42 $X2=0
+ $Y2=0
