* File: sky130_fd_sc_hdll__a32o_4.spice
* Created: Thu Aug 27 18:56:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a32o_4.pex.spice"
.subckt sky130_fd_sc_hdll__a32o_4  VNB VPB A3 A2 A1 B1 B2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1004 N_X_M1004_d N_A_79_21#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.169 PD=0.97 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1006 N_X_M1004_d N_A_79_21#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1018 N_X_M1018_d N_A_79_21#_M1018_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1025 N_X_M1018_d N_A_79_21#_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1022 N_VGND_M1025_s N_A3_M1022_g N_A_485_47#_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1023 N_VGND_M1023_d N_A3_M1023_g N_A_485_47#_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_A_485_47#_M1001_d N_A2_M1001_g N_A_695_47#_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.2015 PD=0.97 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1020 N_A_485_47#_M1001_d N_A2_M1020_g N_A_695_47#_M1020_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1016 N_A_695_47#_M1020_s N_A1_M1016_g N_A_79_21#_M1016_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1026 N_A_695_47#_M1026_d N_A1_M1026_g N_A_79_21#_M1016_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_A_1194_47#_M1007_d N_B1_M1007_g N_A_79_21#_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1017 N_A_1194_47#_M1017_d N_B1_M1017_g N_A_79_21#_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.102375 AS=0.104 PD=0.965 PS=0.97 NRD=7.38 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1011 N_A_1194_47#_M1017_d N_B2_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.102375 AS=0.104 PD=0.965 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1014 N_A_1194_47#_M1014_d N_B2_M1014_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_A_79_21#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A_79_21#_M1008_g N_X_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1015 N_VPWR_M1008_d N_A_79_21#_M1015_g N_X_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1024 N_VPWR_M1024_d N_A_79_21#_M1024_g N_X_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1024_d N_A3_M1005_g N_A_493_297#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1010_d N_A3_M1010_g N_A_493_297#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1019 N_A_493_297#_M1019_d N_A2_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90004.1 A=0.18 P=2.36 MULT=1
MM1027 N_A_493_297#_M1027_d N_A2_M1027_g N_VPWR_M1019_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003.7 A=0.18 P=2.36 MULT=1
MM1003 N_A_493_297#_M1027_d N_A1_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90003.2 A=0.18 P=2.36 MULT=1
MM1012 N_A_493_297#_M1012_d N_A1_M1012_g N_VPWR_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.475 AS=0.145 PD=1.95 PS=1.29 NRD=130.985 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90002.7 A=0.18 P=2.36 MULT=1
MM1000 N_A_79_21#_M1000_d N_B1_M1000_g N_A_493_297#_M1012_d VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.475 PD=1.29 PS=1.95 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.7 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1021 N_A_79_21#_M1000_d N_B1_M1021_g N_A_493_297#_M1021_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.2 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1009 N_A_493_297#_M1021_s N_B2_M1009_g N_A_79_21#_M1009_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.7 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1013 N_A_493_297#_M1013_d N_B2_M1013_g N_A_79_21#_M1009_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.1 SB=90000.2 A=0.18 P=2.36 MULT=1
DX28_noxref VNB VPB NWDIODE A=13.8993 P=20.53
pX29_noxref noxref_16 N_B1_X29_noxref_CONDUCTOR B1 PROBETYPE=1
pX30_noxref noxref_17 N_B1_X29_noxref_CONDUCTOR B1 PROBETYPE=1
pX31_noxref noxref_18 B2 B2 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__a32o_4.pxi.spice"
*
.ends
*
*
