* File: sky130_fd_sc_hdll__a2bb2oi_2.pex.spice
* Created: Wed Sep  2 08:19:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_2%B1 1 3 4 6 7 9 10 12 13 16 21 22
c74 4 0 1.20797e-19 $X=0.52 $Y=0.995
r75 21 22 8.34998 $w=5.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.375 $Y=1.16
+ $X2=0.375 $Y2=1.53
r76 21 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r77 16 19 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.905 $Y=1.16
+ $X2=1.905 $Y2=1.53
r78 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.16 $X2=1.88 $Y2=1.16
r79 14 22 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=0.64 $Y=1.53
+ $X2=0.375 $Y2=1.53
r80 13 19 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.715 $Y=1.53
+ $X2=1.905 $Y2=1.53
r81 13 14 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=1.715 $Y=1.53
+ $X2=0.64 $Y2=1.53
r82 10 17 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.905 $Y2=1.16
r83 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r84 7 17 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.16
r85 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r86 4 26 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.435 $Y2=1.16
r87 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r88 1 26 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.435 $Y2=1.16
r89 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_2%B2 1 3 4 6 7 9 10 12 13 19 20 23
c44 1 0 6.98311e-20 $X=0.94 $Y=0.995
r45 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.46 $Y2=1.202
r46 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=1.2 $Y=1.202
+ $X2=1.435 $Y2=1.202
r47 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2
+ $Y=1.16 $X2=1.2 $Y2=1.16
r48 16 18 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=1.2 $Y2=1.202
r49 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.202
+ $X2=0.965 $Y2=1.202
r50 13 19 7.48636 $w=1.98e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=1.175
+ $X2=1.2 $Y2=1.175
r51 13 23 2.77273 $w=1.98e-07 $l=5e-08 $layer=LI1_cond $X=1.065 $Y=1.175
+ $X2=1.015 $Y2=1.175
r52 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=1.202
r53 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=0.56
r54 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r55 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r56 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r57 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r58 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=1.202
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995 $X2=0.94
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A_455_21# 1 2 3 10 12 13 15 16 18 19 21
+ 22 24 28 30 34 38 42 45 49
r101 48 49 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.845 $Y2=1.202
r102 47 48 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.82 $Y2=1.202
r103 46 47 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.202
+ $X2=2.375 $Y2=1.202
r104 43 49 31.0329 $w=3.65e-07 $l=2.35e-07 $layer=POLY_cond $X=3.08 $Y=1.202
+ $X2=2.845 $Y2=1.202
r105 42 44 21.0935 $w=2.14e-07 $l=3.7e-07 $layer=LI1_cond $X=3.14 $Y=1.16
+ $X2=3.14 $Y2=1.53
r106 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.08
+ $Y=1.16 $X2=3.08 $Y2=1.16
r107 40 42 19.6682 $w=2.14e-07 $l=3.45e-07 $layer=LI1_cond $X=3.14 $Y=0.815
+ $X2=3.14 $Y2=1.16
r108 36 38 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=5.01 $Y=1.615
+ $X2=5.01 $Y2=1.62
r109 32 34 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.985 $Y=0.725
+ $X2=4.985 $Y2=0.39
r110 31 45 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.235 $Y=0.815
+ $X2=4.045 $Y2=0.815
r111 30 32 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=4.795 $Y=0.815
+ $X2=4.985 $Y2=0.725
r112 30 31 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.795 $Y=0.815
+ $X2=4.235 $Y2=0.815
r113 26 45 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=4.045 $Y=0.725
+ $X2=4.045 $Y2=0.815
r114 26 28 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.045 $Y=0.725
+ $X2=4.045 $Y2=0.39
r115 25 44 2.08775 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.285 $Y=1.53
+ $X2=3.14 $Y2=1.53
r116 24 36 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.885 $Y=1.53
+ $X2=5.01 $Y2=1.615
r117 24 25 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=4.885 $Y=1.53
+ $X2=3.285 $Y2=1.53
r118 23 40 1.75188 $w=1.8e-07 $l=1.45e-07 $layer=LI1_cond $X=3.285 $Y=0.815
+ $X2=3.14 $Y2=0.815
r119 22 45 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.855 $Y=0.815
+ $X2=4.045 $Y2=0.815
r120 22 23 35.1212 $w=1.78e-07 $l=5.7e-07 $layer=LI1_cond $X=3.855 $Y=0.815
+ $X2=3.285 $Y2=0.815
r121 19 49 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r122 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r123 16 48 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=1.202
r124 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=0.56
r125 13 47 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r126 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r127 10 46 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.202
r128 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=0.56
r129 3 38 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=1.62
r130 2 34 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.825
+ $Y=0.235 $X2=5.01 $Y2=0.39
r131 1 28 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.885
+ $Y=0.235 $X2=4.07 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A1_N 1 3 4 6 7 9 10 12 13 20 23
r45 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.305 $Y=1.202
+ $X2=4.33 $Y2=1.202
r46 18 20 31.0763 $w=3.8e-07 $l=2.45e-07 $layer=POLY_cond $X=4.06 $Y=1.202
+ $X2=4.305 $Y2=1.202
r47 16 18 28.5395 $w=3.8e-07 $l=2.25e-07 $layer=POLY_cond $X=3.835 $Y=1.202
+ $X2=4.06 $Y2=1.202
r48 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.81 $Y=1.202
+ $X2=3.835 $Y2=1.202
r49 13 23 14.6955 $w=1.98e-07 $l=2.65e-07 $layer=LI1_cond $X=4.06 $Y=1.175
+ $X2=3.795 $Y2=1.175
r50 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.06
+ $Y=1.16 $X2=4.06 $Y2=1.16
r51 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.33 $Y=0.995
+ $X2=4.33 $Y2=1.202
r52 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.33 $Y=0.995
+ $X2=4.33 $Y2=0.56
r53 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.202
r54 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.985
r55 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.202
r56 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.985
r57 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=1.202
r58 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.81 $Y=0.995 $X2=3.81
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A2_N 1 3 4 6 7 9 10 12 13 20 25
r37 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=5.245 $Y=1.202
+ $X2=5.27 $Y2=1.202
r38 19 25 5.82273 $w=1.98e-07 $l=1.05e-07 $layer=LI1_cond $X=5.02 $Y=1.175
+ $X2=5.125 $Y2=1.175
r39 18 20 28.5395 $w=3.8e-07 $l=2.25e-07 $layer=POLY_cond $X=5.02 $Y=1.202
+ $X2=5.245 $Y2=1.202
r40 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.02
+ $Y=1.16 $X2=5.02 $Y2=1.16
r41 16 18 31.0763 $w=3.8e-07 $l=2.45e-07 $layer=POLY_cond $X=4.775 $Y=1.202
+ $X2=5.02 $Y2=1.202
r42 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.75 $Y=1.202
+ $X2=4.775 $Y2=1.202
r43 13 25 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=5.165 $Y=1.175
+ $X2=5.125 $Y2=1.175
r44 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.27 $Y=0.995
+ $X2=5.27 $Y2=1.202
r45 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.27 $Y=0.995
+ $X2=5.27 $Y2=0.56
r46 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.202
r47 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.985
r48 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.202
r49 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
r50 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.75 $Y=0.995
+ $X2=4.75 $Y2=1.202
r51 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.75 $Y=0.995 $X2=4.75
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A_27_297# 1 2 3 4 15 17 18 21 23 29 30
+ 33 35
r43 31 33 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.08 $Y=2.295
+ $X2=3.08 $Y2=1.96
r44 29 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.955 $Y=2.38
+ $X2=3.08 $Y2=2.295
r45 29 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.955 $Y=2.38
+ $X2=2.265 $Y2=2.38
r46 26 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.14 $Y=2.295
+ $X2=2.265 $Y2=2.38
r47 26 28 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.14 $Y=2.295
+ $X2=2.14 $Y2=1.96
r48 25 28 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=2.14 $Y=1.955
+ $X2=2.14 $Y2=1.96
r49 24 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.325 $Y=1.87
+ $X2=1.2 $Y2=1.87
r50 23 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.015 $Y=1.87
+ $X2=2.14 $Y2=1.955
r51 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.015 $Y=1.87
+ $X2=1.325 $Y2=1.87
r52 19 35 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=1.955
+ $X2=1.2 $Y2=1.87
r53 19 21 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.2 $Y=1.955 $X2=1.2
+ $Y2=1.96
r54 17 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.075 $Y=1.87
+ $X2=1.2 $Y2=1.87
r55 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.075 $Y=1.87
+ $X2=0.385 $Y2=1.87
r56 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.26 $Y=1.955
+ $X2=0.385 $Y2=1.87
r57 13 15 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.26 $Y=1.955
+ $X2=0.26 $Y2=1.96
r58 4 33 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=1.96
r59 3 28 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.96
r60 2 21 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.96
r61 1 15 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_2%VPWR 1 2 3 12 14 18 22 25 26 27 29 45 46
+ 49 52
r78 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r79 50 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r80 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r81 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r82 43 46 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.75 $Y2=2.72
r83 42 45 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=5.75 $Y2=2.72
r84 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r85 40 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r86 39 40 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r87 37 40 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.91 $Y2=2.72
r88 37 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r89 36 39 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.91 $Y2=2.72
r90 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r91 34 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.795 $Y=2.72
+ $X2=1.67 $Y2=2.72
r92 34 36 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.795 $Y=2.72
+ $X2=2.07 $Y2=2.72
r93 29 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.605 $Y=2.72
+ $X2=0.73 $Y2=2.72
r94 29 31 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.605 $Y=2.72
+ $X2=0.23 $Y2=2.72
r95 27 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r96 27 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r97 25 39 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.945 $Y=2.72
+ $X2=3.91 $Y2=2.72
r98 25 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.945 $Y=2.72
+ $X2=4.07 $Y2=2.72
r99 24 42 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.195 $Y=2.72
+ $X2=4.37 $Y2=2.72
r100 24 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.195 $Y=2.72
+ $X2=4.07 $Y2=2.72
r101 20 26 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=2.635
+ $X2=4.07 $Y2=2.72
r102 20 22 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.07 $Y=2.635
+ $X2=4.07 $Y2=2.3
r103 16 52 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.72
r104 16 18 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.3
r105 15 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=0.73 $Y2=2.72
r106 14 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.545 $Y=2.72
+ $X2=1.67 $Y2=2.72
r107 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.545 $Y=2.72
+ $X2=0.855 $Y2=2.72
r108 10 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.72
r109 10 12 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.3
r110 3 22 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=2.3
r111 2 18 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.3
r112 1 12 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_2%Y 1 2 3 10 14 19 21 22 23
c45 19 0 1.20797e-19 $X=1.365 $Y=0.775
r46 23 30 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.61 $Y=1.53 $X2=2.61
+ $Y2=1.62
r47 22 23 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.61 $Y=1.19
+ $X2=2.61 $Y2=1.53
r48 20 22 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.61 $Y=0.905
+ $X2=2.61 $Y2=1.19
r49 20 21 2.84597 $w=3.55e-07 $l=1.01735e-07 $layer=LI1_cond $X=2.61 $Y=0.905
+ $X2=2.585 $Y2=0.815
r50 17 19 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.2 $Y=0.775
+ $X2=1.365 $Y2=0.775
r51 12 21 2.84597 $w=3.55e-07 $l=9e-08 $layer=LI1_cond $X=2.585 $Y=0.725
+ $X2=2.585 $Y2=0.815
r52 12 14 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.585 $Y=0.725
+ $X2=2.585 $Y2=0.39
r53 10 21 3.86989 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=0.815
+ $X2=2.585 $Y2=0.815
r54 10 19 63.4646 $w=1.78e-07 $l=1.03e-06 $layer=LI1_cond $X=2.395 $Y=0.815
+ $X2=1.365 $Y2=0.815
r55 3 30 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.62
r56 2 14 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.39
r57 1 17 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A_695_297# 1 2 3 12 14 16 17 18 20 23
r35 18 27 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=2.295
+ $X2=5.48 $Y2=2.38
r36 18 20 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.48 $Y=2.295
+ $X2=5.48 $Y2=1.62
r37 16 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.355 $Y=2.38
+ $X2=5.48 $Y2=2.38
r38 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.355 $Y=2.38
+ $X2=4.665 $Y2=2.38
r39 15 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.54 $Y=2.295
+ $X2=4.665 $Y2=2.38
r40 14 25 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=4.54 $Y=1.965 $X2=4.54
+ $Y2=1.875
r41 14 15 15.2122 $w=2.48e-07 $l=3.3e-07 $layer=LI1_cond $X=4.54 $Y=1.965
+ $X2=4.54 $Y2=2.295
r42 13 23 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.725 $Y=1.875
+ $X2=3.6 $Y2=1.875
r43 12 25 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.415 $Y=1.875
+ $X2=4.54 $Y2=1.875
r44 12 13 42.5152 $w=1.78e-07 $l=6.9e-07 $layer=LI1_cond $X=4.415 $Y=1.875
+ $X2=3.725 $Y2=1.875
r45 3 27 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=2.3
r46 3 20 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=1.62
r47 2 25 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.395
+ $Y=1.485 $X2=4.54 $Y2=1.96
r48 1 23 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=3.475
+ $Y=1.485 $X2=3.6 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_2%VGND 1 2 3 4 5 16 18 22 26 30 33 34 36
+ 37 38 40 58 59 65 70 73
r85 72 73 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=0.235
+ $X2=3.685 $Y2=0.235
r86 68 72 2.80331 $w=6.38e-07 $l=1.5e-07 $layer=LI1_cond $X=3.45 $Y=0.235
+ $X2=3.6 $Y2=0.235
r87 68 70 15.8366 $w=6.38e-07 $l=4.55e-07 $layer=LI1_cond $X=3.45 $Y=0.235
+ $X2=2.995 $Y2=0.235
r88 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r89 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r90 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r91 56 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r92 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r93 53 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r94 53 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.45
+ $Y2=0
r95 52 73 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=4.37 $Y=0 $X2=3.685
+ $Y2=0
r96 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r97 49 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r98 49 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r99 48 70 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.99 $Y=0 $X2=2.995
+ $Y2=0
r100 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r101 46 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=0 $X2=2.14
+ $Y2=0
r102 46 48 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.225 $Y=0
+ $X2=2.99 $Y2=0
r103 44 66 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=2.07 $Y2=0
r104 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r105 41 62 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r106 41 43 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r107 40 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0 $X2=2.14
+ $Y2=0
r108 40 43 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=2.055 $Y=0
+ $X2=0.69 $Y2=0
r109 38 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r110 38 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r111 36 55 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=5.395 $Y=0
+ $X2=5.29 $Y2=0
r112 36 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=0 $X2=5.48
+ $Y2=0
r113 35 58 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.565 $Y=0
+ $X2=5.75 $Y2=0
r114 35 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=0 $X2=5.48
+ $Y2=0
r115 33 52 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=0 $X2=4.37
+ $Y2=0
r116 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=0 $X2=4.54
+ $Y2=0
r117 32 55 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.625 $Y=0 $X2=5.29
+ $Y2=0
r118 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=0 $X2=4.54
+ $Y2=0
r119 28 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0
r120 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.39
r121 24 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0
r122 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0.39
r123 20 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0
r124 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0.39
r125 16 62 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r126 16 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.39
r127 5 30 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.345
+ $Y=0.235 $X2=5.48 $Y2=0.39
r128 4 26 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.405
+ $Y=0.235 $X2=4.54 $Y2=0.39
r129 3 72 91 $w=1.7e-07 $l=7.78653e-07 $layer=licon1_NDIFF $count=2 $X=2.895
+ $Y=0.235 $X2=3.6 $Y2=0.39
r130 2 22 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.39
r131 1 18 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A_119_47# 1 2 7 9 13
c21 9 0 6.98311e-20 $X=0.73 $Y=0.73
r22 11 16 4.05488 $w=2.2e-07 $l=1.5e-07 $layer=LI1_cond $X=0.815 $Y=0.365
+ $X2=0.665 $Y2=0.365
r23 11 13 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=0.815 $Y=0.365
+ $X2=1.67 $Y2=0.365
r24 7 16 2.97358 $w=3e-07 $l=1.1e-07 $layer=LI1_cond $X=0.665 $Y=0.475 $X2=0.665
+ $Y2=0.365
r25 7 9 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=0.665 $Y=0.475
+ $X2=0.665 $Y2=0.73
r26 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.39
r27 1 16 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.39
r28 1 9 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.73
.ends

