* File: sky130_fd_sc_hdll__isobufsrc_1.pex.spice
* Created: Thu Aug 27 19:09:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%A 3 5 7 8 9 10 11
r30 11 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r31 10 11 15.8781 $w=2.23e-07 $l=3.1e-07 $layer=LI1_cond $X=0.212 $Y=0.85
+ $X2=0.212 $Y2=1.16
r32 8 15 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=0.63 $Y=1.16 $X2=0.24
+ $Y2=1.16
r33 8 9 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.63 $Y=1.16 $X2=0.63
+ $Y2=0.995
r34 5 9 34.7346 $w=1.65e-07 $l=4.64543e-07 $layer=POLY_cond $X=0.735 $Y=1.41
+ $X2=0.63 $Y2=0.995
r35 5 7 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.735 $Y=1.41
+ $X2=0.735 $Y2=1.695
r36 1 9 34.7346 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=0.705 $Y=0.995
+ $X2=0.63 $Y2=0.995
r37 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.705 $Y=0.995
+ $X2=0.705 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%SLEEP 1 3 4 6 7 13
c33 1 0 5.50183e-20 $X=1.24 $Y=0.995
r34 7 13 2.21624 $w=2.58e-07 $l=5e-08 $layer=LI1_cond $X=1.2 $Y=1.195 $X2=1.15
+ $Y2=1.195
r35 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.21
+ $Y=1.16 $X2=1.21 $Y2=1.16
r36 4 10 45.964 $w=3.43e-07 $l=2.91548e-07 $layer=POLY_cond $X=1.325 $Y=1.41
+ $X2=1.235 $Y2=1.16
r37 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.325 $Y=1.41
+ $X2=1.325 $Y2=1.985
r38 1 10 38.7084 $w=3.43e-07 $l=1.67481e-07 $layer=POLY_cond $X=1.24 $Y=0.995
+ $X2=1.235 $Y2=1.16
r39 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.24 $Y=0.995 $X2=1.24
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%A_74_47# 1 2 7 9 10 12 15 19 25 27 28
c55 19 0 5.50183e-20 $X=1.77 $Y=1.16
r56 27 30 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.545 $Y=1.595
+ $X2=0.545 $Y2=1.73
r57 27 28 4.86943 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=0.545 $Y=1.595
+ $X2=0.545 $Y2=1.51
r58 23 25 5.7039 $w=1.73e-07 $l=9e-08 $layer=LI1_cond $X=0.495 $Y=0.457
+ $X2=0.585 $Y2=0.457
r59 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.77
+ $Y=1.16 $X2=1.77 $Y2=1.16
r60 17 19 18.3343 $w=2.18e-07 $l=3.5e-07 $layer=LI1_cond $X=1.745 $Y=1.51
+ $X2=1.745 $Y2=1.16
r61 16 27 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.675 $Y=1.595
+ $X2=0.545 $Y2=1.595
r62 15 17 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.635 $Y=1.595
+ $X2=1.745 $Y2=1.51
r63 15 16 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.635 $Y=1.595
+ $X2=0.675 $Y2=1.595
r64 13 25 0.543965 $w=1.8e-07 $l=8.8e-08 $layer=LI1_cond $X=0.585 $Y=0.545
+ $X2=0.585 $Y2=0.457
r65 13 28 59.4596 $w=1.78e-07 $l=9.65e-07 $layer=LI1_cond $X=0.585 $Y=0.545
+ $X2=0.585 $Y2=1.51
r66 10 20 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=1.735 $Y=1.41
+ $X2=1.795 $Y2=1.16
r67 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.735 $Y=1.41
+ $X2=1.735 $Y2=1.985
r68 7 20 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.71 $Y=0.995
+ $X2=1.795 $Y2=1.16
r69 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.71 $Y=0.995 $X2=1.71
+ $Y2=0.56
r70 2 30 600 $w=1.7e-07 $l=3.01081e-07 $layer=licon1_PDIFF $count=1 $X=0.375
+ $Y=1.485 $X2=0.5 $Y2=1.73
r71 1 23 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=0.37
+ $Y=0.235 $X2=0.495 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%VPWR 1 6 8 10 17 18 21
r24 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r25 18 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r26 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r27 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.255 $Y=2.72
+ $X2=1.09 $Y2=2.72
r28 15 17 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=1.255 $Y=2.72
+ $X2=2.07 $Y2=2.72
r29 13 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r30 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r31 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=1.09 $Y2=2.72
r32 10 12 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=0.69 $Y2=2.72
r33 8 13 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r34 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.09 $Y=2.635 $X2=1.09
+ $Y2=2.72
r35 4 6 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.09 $Y=2.635
+ $X2=1.09 $Y2=2
r36 1 6 300 $w=1.7e-07 $l=6.33798e-07 $layer=licon1_PDIFF $count=2 $X=0.825
+ $Y=1.485 $X2=1.09 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%X 1 2 9 11 12 15 18 19
r30 18 19 8.43549 $w=4.48e-07 $l=1.5e-07 $layer=LI1_cond $X=1.98 $Y=2 $X2=1.98
+ $Y2=1.85
r31 15 18 5.5817 $w=4.48e-07 $l=2.1e-07 $layer=LI1_cond $X=1.98 $Y=2.21 $X2=1.98
+ $Y2=2
r32 13 19 63.7727 $w=1.78e-07 $l=1.035e-06 $layer=LI1_cond $X=2.115 $Y=0.815
+ $X2=2.115 $Y2=1.85
r33 11 13 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.025 $Y=0.73
+ $X2=2.115 $Y2=0.815
r34 11 12 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.025 $Y=0.73
+ $X2=1.635 $Y2=0.73
r35 7 12 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=1.46 $Y=0.645
+ $X2=1.635 $Y2=0.73
r36 7 9 8.39637 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=1.46 $Y=0.645
+ $X2=1.46 $Y2=0.39
r37 2 18 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.825
+ $Y=1.485 $X2=1.97 $Y2=2
r38 1 9 91 $w=1.7e-07 $l=2.19203e-07 $layer=licon1_NDIFF $count=2 $X=1.315
+ $Y=0.235 $X2=1.47 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%VGND 1 2 9 11 13 16 17 18 24 30
r35 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r36 27 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r37 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r38 24 29 4.63344 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=1.805 $Y=0 $X2=2.052
+ $Y2=0
r39 24 26 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.805 $Y=0 $X2=1.61
+ $Y2=0
r40 22 27 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r41 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r42 18 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r43 16 21 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.69
+ $Y2=0
r44 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.01
+ $Y2=0
r45 15 26 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.61
+ $Y2=0
r46 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.01
+ $Y2=0
r47 11 29 3.13273 $w=3.3e-07 $l=1.19143e-07 $layer=LI1_cond $X=1.97 $Y=0.085
+ $X2=2.052 $Y2=0
r48 11 13 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.97 $Y=0.085
+ $X2=1.97 $Y2=0.39
r49 7 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.01 $Y=0.085
+ $X2=1.01 $Y2=0
r50 7 9 16.1082 $w=2.08e-07 $l=3.05e-07 $layer=LI1_cond $X=1.01 $Y=0.085
+ $X2=1.01 $Y2=0.39
r51 2 13 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.785
+ $Y=0.235 $X2=1.97 $Y2=0.39
r52 1 9 91 $w=1.7e-07 $l=3.18198e-07 $layer=licon1_NDIFF $count=2 $X=0.78
+ $Y=0.235 $X2=1.03 $Y2=0.39
.ends

