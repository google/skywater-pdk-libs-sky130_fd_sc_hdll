# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__muxb16to1_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__muxb16to1_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  17.02000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D[0]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.335000 1.055000 0.730000 1.325000 ;
        RECT 0.560000 0.395000 0.835000 0.625000 ;
        RECT 0.560000 0.625000 0.730000 1.055000 ;
    END
  END D[0]
  PIN D[1]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765000 0.395000 4.040000 0.625000 ;
        RECT 3.870000 0.625000 4.040000 1.055000 ;
        RECT 3.870000 1.055000 4.265000 1.325000 ;
    END
  END D[1]
  PIN D[2]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.475000 1.055000 4.870000 1.325000 ;
        RECT 4.700000 0.395000 4.975000 0.625000 ;
        RECT 4.700000 0.625000 4.870000 1.055000 ;
    END
  END D[2]
  PIN D[3]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.905000 0.395000 8.180000 0.625000 ;
        RECT 8.010000 0.625000 8.180000 1.055000 ;
        RECT 8.010000 1.055000 8.405000 1.325000 ;
    END
  END D[3]
  PIN D[4]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.615000 1.055000 9.010000 1.325000 ;
        RECT 8.840000 0.395000 9.115000 0.625000 ;
        RECT 8.840000 0.625000 9.010000 1.055000 ;
    END
  END D[4]
  PIN D[5]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.045000 0.395000 12.320000 0.625000 ;
        RECT 12.150000 0.625000 12.320000 1.055000 ;
        RECT 12.150000 1.055000 12.545000 1.325000 ;
    END
  END D[5]
  PIN D[6]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.755000 1.055000 13.150000 1.325000 ;
        RECT 12.980000 0.395000 13.255000 0.625000 ;
        RECT 12.980000 0.625000 13.150000 1.055000 ;
    END
  END D[6]
  PIN D[7]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.185000 0.395000 16.460000 0.625000 ;
        RECT 16.290000 0.625000 16.460000 1.055000 ;
        RECT 16.290000 1.055000 16.685000 1.325000 ;
    END
  END D[7]
  PIN D[8]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.335000 4.115000 0.730000 4.385000 ;
        RECT 0.560000 4.385000 0.730000 4.815000 ;
        RECT 0.560000 4.815000 0.835000 5.045000 ;
    END
  END D[8]
  PIN D[9]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765000 4.815000 4.040000 5.045000 ;
        RECT 3.870000 4.115000 4.265000 4.385000 ;
        RECT 3.870000 4.385000 4.040000 4.815000 ;
    END
  END D[9]
  PIN D[10]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.475000 4.115000 4.870000 4.385000 ;
        RECT 4.700000 4.385000 4.870000 4.815000 ;
        RECT 4.700000 4.815000 4.975000 5.045000 ;
    END
  END D[10]
  PIN D[11]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.905000 4.815000 8.180000 5.045000 ;
        RECT 8.010000 4.115000 8.405000 4.385000 ;
        RECT 8.010000 4.385000 8.180000 4.815000 ;
    END
  END D[11]
  PIN D[12]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.615000 4.115000 9.010000 4.385000 ;
        RECT 8.840000 4.385000 9.010000 4.815000 ;
        RECT 8.840000 4.815000 9.115000 5.045000 ;
    END
  END D[12]
  PIN D[13]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.045000 4.815000 12.320000 5.045000 ;
        RECT 12.150000 4.115000 12.545000 4.385000 ;
        RECT 12.150000 4.385000 12.320000 4.815000 ;
    END
  END D[13]
  PIN D[14]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.755000 4.115000 13.150000 4.385000 ;
        RECT 12.980000 4.385000 13.150000 4.815000 ;
        RECT 12.980000 4.815000 13.255000 5.045000 ;
    END
  END D[14]
  PIN D[15]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.185000 4.815000 16.460000 5.045000 ;
        RECT 16.290000 4.115000 16.685000 4.385000 ;
        RECT 16.290000 4.385000 16.460000 4.815000 ;
    END
  END D[15]
  PIN S[0]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805000 0.945000 2.205000 1.295000 ;
    END
  END S[0]
  PIN S[1]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.395000 0.945000 2.795000 1.295000 ;
    END
  END S[1]
  PIN S[2]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.945000 0.945000 6.345000 1.295000 ;
    END
  END S[2]
  PIN S[3]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.535000 0.945000 6.935000 1.295000 ;
    END
  END S[3]
  PIN S[4]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.085000 0.945000 10.485000 1.295000 ;
    END
  END S[4]
  PIN S[5]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.675000 0.945000 11.075000 1.295000 ;
    END
  END S[5]
  PIN S[6]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.225000 0.945000 14.625000 1.295000 ;
    END
  END S[6]
  PIN S[7]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.815000 0.945000 15.215000 1.295000 ;
    END
  END S[7]
  PIN S[8]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805000 4.145000 2.205000 4.495000 ;
    END
  END S[8]
  PIN S[9]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.395000 4.145000 2.795000 4.495000 ;
    END
  END S[9]
  PIN S[10]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.945000 4.145000 6.345000 4.495000 ;
    END
  END S[10]
  PIN S[11]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.535000 4.145000 6.935000 4.495000 ;
    END
  END S[11]
  PIN S[12]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.085000 4.145000 10.485000 4.495000 ;
    END
  END S[12]
  PIN S[13]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.675000 4.145000 11.075000 4.495000 ;
    END
  END S[13]
  PIN S[14]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.225000 4.145000 14.625000 4.495000 ;
    END
  END S[14]
  PIN S[15]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.815000 4.145000 15.215000 4.495000 ;
    END
  END S[15]
  PIN VGND
    ANTENNADIFFAREA  1.875900 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 17.020000 0.085000 ;
        RECT  0.130000  0.085000  0.390000 0.885000 ;
        RECT  2.135000  0.085000  2.465000 0.660000 ;
        RECT  4.210000  0.085000  4.530000 0.885000 ;
        RECT  6.275000  0.085000  6.605000 0.660000 ;
        RECT  8.350000  0.085000  8.670000 0.885000 ;
        RECT 10.415000  0.085000 10.745000 0.660000 ;
        RECT 12.490000  0.085000 12.810000 0.885000 ;
        RECT 14.555000  0.085000 14.885000 0.660000 ;
        RECT 16.630000  0.085000 16.890000 0.885000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
        RECT 10.725000 -0.085000 10.895000 0.085000 ;
        RECT 11.185000 -0.085000 11.355000 0.085000 ;
        RECT 11.645000 -0.085000 11.815000 0.085000 ;
        RECT 12.105000 -0.085000 12.275000 0.085000 ;
        RECT 12.565000 -0.085000 12.735000 0.085000 ;
        RECT 13.025000 -0.085000 13.195000 0.085000 ;
        RECT 13.485000 -0.085000 13.655000 0.085000 ;
        RECT 13.945000 -0.085000 14.115000 0.085000 ;
        RECT 14.405000 -0.085000 14.575000 0.085000 ;
        RECT 14.865000 -0.085000 15.035000 0.085000 ;
        RECT 15.325000 -0.085000 15.495000 0.085000 ;
        RECT 15.785000 -0.085000 15.955000 0.085000 ;
        RECT 16.245000 -0.085000 16.415000 0.085000 ;
        RECT 16.705000 -0.085000 16.875000 0.085000 ;
    END
    PORT
      LAYER li1 ;
        RECT  0.000000 5.355000 17.020000 5.525000 ;
        RECT  0.130000 4.555000  0.390000 5.355000 ;
        RECT  2.135000 4.780000  2.465000 5.355000 ;
        RECT  4.210000 4.555000  4.530000 5.355000 ;
        RECT  6.275000 4.780000  6.605000 5.355000 ;
        RECT  8.350000 4.555000  8.670000 5.355000 ;
        RECT 10.415000 4.780000 10.745000 5.355000 ;
        RECT 12.490000 4.555000 12.810000 5.355000 ;
        RECT 14.555000 4.780000 14.885000 5.355000 ;
        RECT 16.630000 4.555000 16.890000 5.355000 ;
      LAYER mcon ;
        RECT  0.145000 5.355000  0.315000 5.525000 ;
        RECT  0.605000 5.355000  0.775000 5.525000 ;
        RECT  1.065000 5.355000  1.235000 5.525000 ;
        RECT  1.525000 5.355000  1.695000 5.525000 ;
        RECT  1.985000 5.355000  2.155000 5.525000 ;
        RECT  2.445000 5.355000  2.615000 5.525000 ;
        RECT  2.905000 5.355000  3.075000 5.525000 ;
        RECT  3.365000 5.355000  3.535000 5.525000 ;
        RECT  3.825000 5.355000  3.995000 5.525000 ;
        RECT  4.285000 5.355000  4.455000 5.525000 ;
        RECT  4.745000 5.355000  4.915000 5.525000 ;
        RECT  5.205000 5.355000  5.375000 5.525000 ;
        RECT  5.665000 5.355000  5.835000 5.525000 ;
        RECT  6.125000 5.355000  6.295000 5.525000 ;
        RECT  6.585000 5.355000  6.755000 5.525000 ;
        RECT  7.045000 5.355000  7.215000 5.525000 ;
        RECT  7.505000 5.355000  7.675000 5.525000 ;
        RECT  7.965000 5.355000  8.135000 5.525000 ;
        RECT  8.425000 5.355000  8.595000 5.525000 ;
        RECT  8.885000 5.355000  9.055000 5.525000 ;
        RECT  9.345000 5.355000  9.515000 5.525000 ;
        RECT  9.805000 5.355000  9.975000 5.525000 ;
        RECT 10.265000 5.355000 10.435000 5.525000 ;
        RECT 10.725000 5.355000 10.895000 5.525000 ;
        RECT 11.185000 5.355000 11.355000 5.525000 ;
        RECT 11.645000 5.355000 11.815000 5.525000 ;
        RECT 12.105000 5.355000 12.275000 5.525000 ;
        RECT 12.565000 5.355000 12.735000 5.525000 ;
        RECT 13.025000 5.355000 13.195000 5.525000 ;
        RECT 13.485000 5.355000 13.655000 5.525000 ;
        RECT 13.945000 5.355000 14.115000 5.525000 ;
        RECT 14.405000 5.355000 14.575000 5.525000 ;
        RECT 14.865000 5.355000 15.035000 5.525000 ;
        RECT 15.325000 5.355000 15.495000 5.525000 ;
        RECT 15.785000 5.355000 15.955000 5.525000 ;
        RECT 16.245000 5.355000 16.415000 5.525000 ;
        RECT 16.705000 5.355000 16.875000 5.525000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 17.020000 0.240000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 17.020000 5.680000 ;
    END
  END VGND
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
    PORT
      LAYER pwell ;
        RECT 0.145000 5.355000 0.315000 5.525000 ;
    END
    PORT
      LAYER pwell ;
        RECT 12.565000 -0.085000 12.735000 0.085000 ;
    END
    PORT
      LAYER pwell ;
        RECT 12.565000 5.355000 12.735000 5.525000 ;
    END
    PORT
      LAYER pwell ;
        RECT 16.705000 -0.085000 16.875000 0.085000 ;
    END
    PORT
      LAYER pwell ;
        RECT 16.705000 5.355000 16.875000 5.525000 ;
    END
    PORT
      LAYER pwell ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
    END
    PORT
      LAYER pwell ;
        RECT 4.285000 5.355000 4.455000 5.525000 ;
    END
    PORT
      LAYER pwell ;
        RECT 8.425000 -0.085000 8.595000 0.085000 ;
    END
    PORT
      LAYER pwell ;
        RECT 8.425000 5.355000 8.595000 5.525000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 17.210000 4.135000 ;
    END
  END VPB
  PIN VPWR
    ANTENNADIFFAREA  6.380000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 0.920000 2.805000 ;
        RECT 0.095000 1.495000 0.425000 2.635000 ;
        RECT 0.095000 2.805000 0.425000 3.945000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
    END
    PORT
      LAYER li1 ;
        RECT 11.960000 2.635000 13.340000 2.805000 ;
        RECT 12.455000 1.495000 12.845000 2.635000 ;
        RECT 12.455000 2.805000 12.845000 3.945000 ;
      LAYER mcon ;
        RECT 12.105000 2.635000 12.275000 2.805000 ;
        RECT 12.565000 2.635000 12.735000 2.805000 ;
        RECT 13.025000 2.635000 13.195000 2.805000 ;
    END
    PORT
      LAYER li1 ;
        RECT 16.100000 2.635000 17.020000 2.805000 ;
        RECT 16.595000 1.495000 16.925000 2.635000 ;
        RECT 16.595000 2.805000 16.925000 3.945000 ;
      LAYER mcon ;
        RECT 16.245000 2.635000 16.415000 2.805000 ;
        RECT 16.705000 2.635000 16.875000 2.805000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.680000 2.635000 5.060000 2.805000 ;
        RECT 4.175000 1.495000 4.565000 2.635000 ;
        RECT 4.175000 2.805000 4.565000 3.945000 ;
      LAYER mcon ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.820000 2.635000 9.200000 2.805000 ;
        RECT 8.315000 1.495000 8.705000 2.635000 ;
        RECT 8.315000 2.805000 8.705000 3.945000 ;
      LAYER mcon ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
        RECT 8.425000 2.635000 8.595000 2.805000 ;
        RECT 8.885000 2.635000 9.055000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 17.020000 2.960000 ;
    END
  END VPWR
  PIN Z
    ANTENNADIFFAREA  5.705600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.900000 0.835000 1.290000 1.005000 ;
        RECT 0.900000 1.005000 1.070000 1.755000 ;
        RECT 0.900000 1.755000 1.295000 1.805000 ;
        RECT 0.900000 1.805000 1.420000 1.985000 ;
        RECT 0.900000 3.455000 1.420000 3.635000 ;
        RECT 0.900000 3.635000 1.295000 3.685000 ;
        RECT 0.900000 3.685000 1.070000 4.435000 ;
        RECT 0.900000 4.435000 1.290000 4.605000 ;
        RECT 1.045000 0.330000 1.290000 0.835000 ;
        RECT 1.045000 4.605000 1.290000 5.110000 ;
        RECT 1.090000 1.985000 1.420000 2.465000 ;
        RECT 1.090000 2.465000 1.295000 2.975000 ;
        RECT 1.090000 2.975000 1.420000 3.455000 ;
      LAYER mcon ;
        RECT 1.065000 1.785000 1.235000 1.955000 ;
        RECT 1.065000 3.485000 1.235000 3.655000 ;
    END
    PORT
      LAYER li1 ;
        RECT 11.460000 1.805000 11.980000 1.985000 ;
        RECT 11.460000 1.985000 11.790000 2.465000 ;
        RECT 11.460000 2.975000 11.790000 3.455000 ;
        RECT 11.460000 3.455000 11.980000 3.635000 ;
        RECT 11.585000 1.755000 11.980000 1.805000 ;
        RECT 11.585000 2.465000 11.790000 2.975000 ;
        RECT 11.585000 3.635000 11.980000 3.685000 ;
        RECT 11.590000 0.330000 11.835000 0.835000 ;
        RECT 11.590000 0.835000 11.980000 1.005000 ;
        RECT 11.590000 4.435000 11.980000 4.605000 ;
        RECT 11.590000 4.605000 11.835000 5.110000 ;
        RECT 11.810000 1.005000 11.980000 1.755000 ;
        RECT 11.810000 3.685000 11.980000 4.435000 ;
      LAYER mcon ;
        RECT 11.645000 1.785000 11.815000 1.955000 ;
        RECT 11.645000 3.485000 11.815000 3.655000 ;
    END
    PORT
      LAYER li1 ;
        RECT 13.320000 0.835000 13.710000 1.005000 ;
        RECT 13.320000 1.005000 13.490000 1.755000 ;
        RECT 13.320000 1.755000 13.715000 1.805000 ;
        RECT 13.320000 1.805000 13.840000 1.985000 ;
        RECT 13.320000 3.455000 13.840000 3.635000 ;
        RECT 13.320000 3.635000 13.715000 3.685000 ;
        RECT 13.320000 3.685000 13.490000 4.435000 ;
        RECT 13.320000 4.435000 13.710000 4.605000 ;
        RECT 13.465000 0.330000 13.710000 0.835000 ;
        RECT 13.465000 4.605000 13.710000 5.110000 ;
        RECT 13.510000 1.985000 13.840000 2.465000 ;
        RECT 13.510000 2.465000 13.715000 2.975000 ;
        RECT 13.510000 2.975000 13.840000 3.455000 ;
      LAYER mcon ;
        RECT 13.485000 1.785000 13.655000 1.955000 ;
        RECT 13.485000 3.485000 13.655000 3.655000 ;
    END
    PORT
      LAYER li1 ;
        RECT 15.600000 1.805000 16.120000 1.985000 ;
        RECT 15.600000 1.985000 15.930000 2.465000 ;
        RECT 15.600000 2.975000 15.930000 3.455000 ;
        RECT 15.600000 3.455000 16.120000 3.635000 ;
        RECT 15.725000 1.755000 16.120000 1.805000 ;
        RECT 15.725000 2.465000 15.930000 2.975000 ;
        RECT 15.725000 3.635000 16.120000 3.685000 ;
        RECT 15.730000 0.330000 15.975000 0.835000 ;
        RECT 15.730000 0.835000 16.120000 1.005000 ;
        RECT 15.730000 4.435000 16.120000 4.605000 ;
        RECT 15.730000 4.605000 15.975000 5.110000 ;
        RECT 15.950000 1.005000 16.120000 1.755000 ;
        RECT 15.950000 3.685000 16.120000 4.435000 ;
      LAYER mcon ;
        RECT 15.785000 1.785000 15.955000 1.955000 ;
        RECT 15.785000 3.485000 15.955000 3.655000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.180000 1.805000 3.700000 1.985000 ;
        RECT 3.180000 1.985000 3.510000 2.465000 ;
        RECT 3.180000 2.975000 3.510000 3.455000 ;
        RECT 3.180000 3.455000 3.700000 3.635000 ;
        RECT 3.305000 1.755000 3.700000 1.805000 ;
        RECT 3.305000 2.465000 3.510000 2.975000 ;
        RECT 3.305000 3.635000 3.700000 3.685000 ;
        RECT 3.310000 0.330000 3.555000 0.835000 ;
        RECT 3.310000 0.835000 3.700000 1.005000 ;
        RECT 3.310000 4.435000 3.700000 4.605000 ;
        RECT 3.310000 4.605000 3.555000 5.110000 ;
        RECT 3.530000 1.005000 3.700000 1.755000 ;
        RECT 3.530000 3.685000 3.700000 4.435000 ;
      LAYER mcon ;
        RECT 3.365000 1.785000 3.535000 1.955000 ;
        RECT 3.365000 3.485000 3.535000 3.655000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.040000 0.835000 5.430000 1.005000 ;
        RECT 5.040000 1.005000 5.210000 1.755000 ;
        RECT 5.040000 1.755000 5.435000 1.805000 ;
        RECT 5.040000 1.805000 5.560000 1.985000 ;
        RECT 5.040000 3.455000 5.560000 3.635000 ;
        RECT 5.040000 3.635000 5.435000 3.685000 ;
        RECT 5.040000 3.685000 5.210000 4.435000 ;
        RECT 5.040000 4.435000 5.430000 4.605000 ;
        RECT 5.185000 0.330000 5.430000 0.835000 ;
        RECT 5.185000 4.605000 5.430000 5.110000 ;
        RECT 5.230000 1.985000 5.560000 2.465000 ;
        RECT 5.230000 2.465000 5.435000 2.975000 ;
        RECT 5.230000 2.975000 5.560000 3.455000 ;
      LAYER mcon ;
        RECT 5.205000 1.785000 5.375000 1.955000 ;
        RECT 5.205000 3.485000 5.375000 3.655000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.320000 1.805000 7.840000 1.985000 ;
        RECT 7.320000 1.985000 7.650000 2.465000 ;
        RECT 7.320000 2.975000 7.650000 3.455000 ;
        RECT 7.320000 3.455000 7.840000 3.635000 ;
        RECT 7.445000 1.755000 7.840000 1.805000 ;
        RECT 7.445000 2.465000 7.650000 2.975000 ;
        RECT 7.445000 3.635000 7.840000 3.685000 ;
        RECT 7.450000 0.330000 7.695000 0.835000 ;
        RECT 7.450000 0.835000 7.840000 1.005000 ;
        RECT 7.450000 4.435000 7.840000 4.605000 ;
        RECT 7.450000 4.605000 7.695000 5.110000 ;
        RECT 7.670000 1.005000 7.840000 1.755000 ;
        RECT 7.670000 3.685000 7.840000 4.435000 ;
      LAYER mcon ;
        RECT 7.505000 1.785000 7.675000 1.955000 ;
        RECT 7.505000 3.485000 7.675000 3.655000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.180000 0.835000 9.570000 1.005000 ;
        RECT 9.180000 1.005000 9.350000 1.755000 ;
        RECT 9.180000 1.755000 9.575000 1.805000 ;
        RECT 9.180000 1.805000 9.700000 1.985000 ;
        RECT 9.180000 3.455000 9.700000 3.635000 ;
        RECT 9.180000 3.635000 9.575000 3.685000 ;
        RECT 9.180000 3.685000 9.350000 4.435000 ;
        RECT 9.180000 4.435000 9.570000 4.605000 ;
        RECT 9.325000 0.330000 9.570000 0.835000 ;
        RECT 9.325000 4.605000 9.570000 5.110000 ;
        RECT 9.370000 1.985000 9.700000 2.465000 ;
        RECT 9.370000 2.465000 9.575000 2.975000 ;
        RECT 9.370000 2.975000 9.700000 3.455000 ;
      LAYER mcon ;
        RECT 9.345000 1.785000 9.515000 1.955000 ;
        RECT 9.345000 3.485000 9.515000 3.655000 ;
    END
    PORT
      LAYER met1 ;
        RECT  1.005000 1.755000  1.295000 1.800000 ;
        RECT  1.005000 1.800000 16.015000 1.940000 ;
        RECT  1.005000 1.940000  1.295000 1.985000 ;
        RECT  1.005000 3.455000  1.295000 3.500000 ;
        RECT  1.005000 3.500000 16.015000 3.640000 ;
        RECT  1.005000 3.640000  1.295000 3.685000 ;
        RECT  3.305000 1.755000  3.595000 1.800000 ;
        RECT  3.305000 1.940000  3.595000 1.985000 ;
        RECT  3.305000 3.455000  3.595000 3.500000 ;
        RECT  3.305000 3.640000  3.595000 3.685000 ;
        RECT  5.145000 1.755000  5.435000 1.800000 ;
        RECT  5.145000 1.940000  5.435000 1.985000 ;
        RECT  5.145000 3.455000  5.435000 3.500000 ;
        RECT  5.145000 3.640000  5.435000 3.685000 ;
        RECT  7.445000 1.755000  7.735000 1.800000 ;
        RECT  7.445000 1.940000  7.735000 1.985000 ;
        RECT  7.445000 3.455000  7.735000 3.500000 ;
        RECT  7.445000 3.640000  7.735000 3.685000 ;
        RECT  9.285000 1.755000  9.575000 1.800000 ;
        RECT  9.285000 1.940000  9.575000 1.985000 ;
        RECT  9.285000 3.455000  9.575000 3.500000 ;
        RECT  9.285000 3.640000  9.575000 3.685000 ;
        RECT 11.585000 1.755000 11.875000 1.800000 ;
        RECT 11.585000 1.940000 11.875000 1.985000 ;
        RECT 11.585000 3.455000 11.875000 3.500000 ;
        RECT 11.585000 3.640000 11.875000 3.685000 ;
        RECT 13.425000 1.755000 13.715000 1.800000 ;
        RECT 13.425000 1.940000 13.715000 1.985000 ;
        RECT 13.425000 3.455000 13.715000 3.500000 ;
        RECT 13.425000 3.640000 13.715000 3.685000 ;
        RECT 15.725000 1.755000 16.015000 1.800000 ;
        RECT 15.725000 1.940000 16.015000 1.985000 ;
        RECT 15.725000 3.455000 16.015000 3.500000 ;
        RECT 15.725000 3.640000 16.015000 3.685000 ;
    END
  END Z
  OBS
    LAYER li1 ;
      RECT  1.240000 1.175000  1.630000 1.465000 ;
      RECT  1.240000 1.465000  1.940000 1.505000 ;
      RECT  1.240000 3.935000  1.940000 3.975000 ;
      RECT  1.240000 3.975000  1.630000 4.265000 ;
      RECT  1.460000 0.585000  1.900000 0.755000 ;
      RECT  1.460000 0.755000  1.630000 1.175000 ;
      RECT  1.460000 1.505000  1.940000 1.635000 ;
      RECT  1.460000 3.805000  1.940000 3.935000 ;
      RECT  1.460000 4.265000  1.630000 4.685000 ;
      RECT  1.460000 4.685000  1.900000 4.855000 ;
      RECT  1.465000 2.635000  3.135000 2.805000 ;
      RECT  1.610000 1.635000  1.940000 2.465000 ;
      RECT  1.610000 2.975000  1.940000 3.805000 ;
      RECT  1.650000 0.330000  1.900000 0.585000 ;
      RECT  1.650000 4.855000  1.900000 5.110000 ;
      RECT  2.135000 1.465000  2.465000 2.635000 ;
      RECT  2.135000 2.805000  2.465000 3.975000 ;
      RECT  2.660000 1.465000  3.360000 1.505000 ;
      RECT  2.660000 1.505000  3.140000 1.635000 ;
      RECT  2.660000 1.635000  2.990000 2.465000 ;
      RECT  2.660000 2.975000  2.990000 3.805000 ;
      RECT  2.660000 3.805000  3.140000 3.935000 ;
      RECT  2.660000 3.935000  3.360000 3.975000 ;
      RECT  2.700000 0.330000  2.950000 0.585000 ;
      RECT  2.700000 0.585000  3.140000 0.755000 ;
      RECT  2.700000 4.685000  3.140000 4.855000 ;
      RECT  2.700000 4.855000  2.950000 5.110000 ;
      RECT  2.970000 0.755000  3.140000 1.175000 ;
      RECT  2.970000 1.175000  3.360000 1.465000 ;
      RECT  2.970000 3.975000  3.360000 4.265000 ;
      RECT  2.970000 4.265000  3.140000 4.685000 ;
      RECT  5.380000 1.175000  5.770000 1.465000 ;
      RECT  5.380000 1.465000  6.080000 1.505000 ;
      RECT  5.380000 3.935000  6.080000 3.975000 ;
      RECT  5.380000 3.975000  5.770000 4.265000 ;
      RECT  5.600000 0.585000  6.040000 0.755000 ;
      RECT  5.600000 0.755000  5.770000 1.175000 ;
      RECT  5.600000 1.505000  6.080000 1.635000 ;
      RECT  5.600000 3.805000  6.080000 3.935000 ;
      RECT  5.600000 4.265000  5.770000 4.685000 ;
      RECT  5.600000 4.685000  6.040000 4.855000 ;
      RECT  5.605000 2.635000  7.275000 2.805000 ;
      RECT  5.750000 1.635000  6.080000 2.465000 ;
      RECT  5.750000 2.975000  6.080000 3.805000 ;
      RECT  5.790000 0.330000  6.040000 0.585000 ;
      RECT  5.790000 4.855000  6.040000 5.110000 ;
      RECT  6.275000 1.465000  6.605000 2.635000 ;
      RECT  6.275000 2.805000  6.605000 3.975000 ;
      RECT  6.800000 1.465000  7.500000 1.505000 ;
      RECT  6.800000 1.505000  7.280000 1.635000 ;
      RECT  6.800000 1.635000  7.130000 2.465000 ;
      RECT  6.800000 2.975000  7.130000 3.805000 ;
      RECT  6.800000 3.805000  7.280000 3.935000 ;
      RECT  6.800000 3.935000  7.500000 3.975000 ;
      RECT  6.840000 0.330000  7.090000 0.585000 ;
      RECT  6.840000 0.585000  7.280000 0.755000 ;
      RECT  6.840000 4.685000  7.280000 4.855000 ;
      RECT  6.840000 4.855000  7.090000 5.110000 ;
      RECT  7.110000 0.755000  7.280000 1.175000 ;
      RECT  7.110000 1.175000  7.500000 1.465000 ;
      RECT  7.110000 3.975000  7.500000 4.265000 ;
      RECT  7.110000 4.265000  7.280000 4.685000 ;
      RECT  9.520000 1.175000  9.910000 1.465000 ;
      RECT  9.520000 1.465000 10.220000 1.505000 ;
      RECT  9.520000 3.935000 10.220000 3.975000 ;
      RECT  9.520000 3.975000  9.910000 4.265000 ;
      RECT  9.740000 0.585000 10.180000 0.755000 ;
      RECT  9.740000 0.755000  9.910000 1.175000 ;
      RECT  9.740000 1.505000 10.220000 1.635000 ;
      RECT  9.740000 3.805000 10.220000 3.935000 ;
      RECT  9.740000 4.265000  9.910000 4.685000 ;
      RECT  9.740000 4.685000 10.180000 4.855000 ;
      RECT  9.745000 2.635000 11.415000 2.805000 ;
      RECT  9.890000 1.635000 10.220000 2.465000 ;
      RECT  9.890000 2.975000 10.220000 3.805000 ;
      RECT  9.930000 0.330000 10.180000 0.585000 ;
      RECT  9.930000 4.855000 10.180000 5.110000 ;
      RECT 10.415000 1.465000 10.745000 2.635000 ;
      RECT 10.415000 2.805000 10.745000 3.975000 ;
      RECT 10.940000 1.465000 11.640000 1.505000 ;
      RECT 10.940000 1.505000 11.420000 1.635000 ;
      RECT 10.940000 1.635000 11.270000 2.465000 ;
      RECT 10.940000 2.975000 11.270000 3.805000 ;
      RECT 10.940000 3.805000 11.420000 3.935000 ;
      RECT 10.940000 3.935000 11.640000 3.975000 ;
      RECT 10.980000 0.330000 11.230000 0.585000 ;
      RECT 10.980000 0.585000 11.420000 0.755000 ;
      RECT 10.980000 4.685000 11.420000 4.855000 ;
      RECT 10.980000 4.855000 11.230000 5.110000 ;
      RECT 11.250000 0.755000 11.420000 1.175000 ;
      RECT 11.250000 1.175000 11.640000 1.465000 ;
      RECT 11.250000 3.975000 11.640000 4.265000 ;
      RECT 11.250000 4.265000 11.420000 4.685000 ;
      RECT 13.660000 1.175000 14.050000 1.465000 ;
      RECT 13.660000 1.465000 14.360000 1.505000 ;
      RECT 13.660000 3.935000 14.360000 3.975000 ;
      RECT 13.660000 3.975000 14.050000 4.265000 ;
      RECT 13.880000 0.585000 14.320000 0.755000 ;
      RECT 13.880000 0.755000 14.050000 1.175000 ;
      RECT 13.880000 1.505000 14.360000 1.635000 ;
      RECT 13.880000 3.805000 14.360000 3.935000 ;
      RECT 13.880000 4.265000 14.050000 4.685000 ;
      RECT 13.880000 4.685000 14.320000 4.855000 ;
      RECT 13.885000 2.635000 15.555000 2.805000 ;
      RECT 14.030000 1.635000 14.360000 2.465000 ;
      RECT 14.030000 2.975000 14.360000 3.805000 ;
      RECT 14.070000 0.330000 14.320000 0.585000 ;
      RECT 14.070000 4.855000 14.320000 5.110000 ;
      RECT 14.555000 1.465000 14.885000 2.635000 ;
      RECT 14.555000 2.805000 14.885000 3.975000 ;
      RECT 15.080000 1.465000 15.780000 1.505000 ;
      RECT 15.080000 1.505000 15.560000 1.635000 ;
      RECT 15.080000 1.635000 15.410000 2.465000 ;
      RECT 15.080000 2.975000 15.410000 3.805000 ;
      RECT 15.080000 3.805000 15.560000 3.935000 ;
      RECT 15.080000 3.935000 15.780000 3.975000 ;
      RECT 15.120000 0.330000 15.370000 0.585000 ;
      RECT 15.120000 0.585000 15.560000 0.755000 ;
      RECT 15.120000 4.685000 15.560000 4.855000 ;
      RECT 15.120000 4.855000 15.370000 5.110000 ;
      RECT 15.390000 0.755000 15.560000 1.175000 ;
      RECT 15.390000 1.175000 15.780000 1.465000 ;
      RECT 15.390000 3.975000 15.780000 4.265000 ;
      RECT 15.390000 4.265000 15.560000 4.685000 ;
    LAYER mcon ;
      RECT  1.525000 2.635000  1.695000 2.805000 ;
      RECT  1.985000 2.635000  2.155000 2.805000 ;
      RECT  2.445000 2.635000  2.615000 2.805000 ;
      RECT  2.905000 2.635000  3.075000 2.805000 ;
      RECT  5.665000 2.635000  5.835000 2.805000 ;
      RECT  6.125000 2.635000  6.295000 2.805000 ;
      RECT  6.585000 2.635000  6.755000 2.805000 ;
      RECT  7.045000 2.635000  7.215000 2.805000 ;
      RECT  9.805000 2.635000  9.975000 2.805000 ;
      RECT 10.265000 2.635000 10.435000 2.805000 ;
      RECT 10.725000 2.635000 10.895000 2.805000 ;
      RECT 11.185000 2.635000 11.355000 2.805000 ;
      RECT 13.945000 2.635000 14.115000 2.805000 ;
      RECT 14.405000 2.635000 14.575000 2.805000 ;
      RECT 14.865000 2.635000 15.035000 2.805000 ;
      RECT 15.325000 2.635000 15.495000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb16to1_1
END LIBRARY
