* File: sky130_fd_sc_hdll__o211a_1.pex.spice
* Created: Thu Aug 27 19:18:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O211A_1%A_79_21# 1 2 3 12 14 16 17 23 24 25 28 30
+ 33 36 39 41 45
c82 23 0 1.32642e-19 $X=1.09 $Y=1.495
r83 41 43 14.9958 $w=5.48e-07 $l=4.85e-07 $layer=LI1_cond $X=3.525 $Y=0.38
+ $X2=3.525 $Y2=0.865
r84 34 45 3.40559 $w=2.75e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.635 $Y=1.665
+ $X2=3.525 $Y2=1.58
r85 34 36 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.635 $Y=1.665
+ $X2=3.635 $Y2=2.34
r86 33 45 3.40559 $w=2.75e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.36 $Y=1.495
+ $X2=3.525 $Y2=1.58
r87 33 43 33.0018 $w=2.18e-07 $l=6.3e-07 $layer=LI1_cond $X=3.36 $Y=1.495
+ $X2=3.36 $Y2=0.865
r88 31 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.465 $Y=1.58
+ $X2=2.275 $Y2=1.58
r89 30 45 3.11956 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.25 $Y=1.58
+ $X2=3.525 $Y2=1.58
r90 30 31 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=3.25 $Y=1.58
+ $X2=2.465 $Y2=1.58
r91 26 39 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=1.665
+ $X2=2.275 $Y2=1.58
r92 26 28 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=2.275 $Y=1.665
+ $X2=2.275 $Y2=2.34
r93 24 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.085 $Y=1.58
+ $X2=2.275 $Y2=1.58
r94 24 25 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=2.085 $Y=1.58
+ $X2=1.175 $Y2=1.58
r95 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.09 $Y=1.495
+ $X2=1.175 $Y2=1.58
r96 22 23 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.09 $Y=1.245
+ $X2=1.09 $Y2=1.495
r97 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.595
+ $Y=1.16 $X2=0.595 $Y2=1.16
r98 17 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.005 $Y=1.16
+ $X2=1.09 $Y2=1.245
r99 17 19 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.005 $Y=1.16
+ $X2=0.595 $Y2=1.16
r100 14 20 45.7629 $w=3.5e-07 $l=2.98747e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.602 $Y2=1.16
r101 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r102 10 20 34.6525 $w=3.5e-07 $l=1.89855e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.602 $Y2=1.16
r103 10 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=0.56
r104 3 45 400 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_PDIFF $count=1 $X=3.45
+ $Y=1.485 $X2=3.635 $Y2=1.66
r105 3 36 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=3.45
+ $Y=1.485 $X2=3.635 $Y2=2.34
r106 2 39 400 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=1.485 $X2=2.3 $Y2=1.66
r107 2 28 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=1.485 $X2=2.3 $Y2=2.34
r108 1 41 91 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=2 $X=3.41
+ $Y=0.235 $X2=3.635 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_1%A1 1 3 4 6 7 15
c32 4 0 1.75245e-19 $X=1.485 $Y=1.41
r33 7 15 6.1 $w=1.98e-07 $l=1.1e-07 $layer=LI1_cond $X=1.525 $Y=1.175 $X2=1.635
+ $Y2=1.175
r34 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.525
+ $Y=1.16 $X2=1.525 $Y2=1.16
r35 4 10 48.3784 $w=2.91e-07 $l=2.77038e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.542 $Y2=1.16
r36 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.985
r37 1 10 38.6072 $w=2.91e-07 $l=2.01879e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.542 $Y2=1.16
r38 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.46 $Y=0.995 $X2=1.46
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_1%A2 1 3 4 6 7 14
c29 7 0 1.75245e-19 $X=2.16 $Y=1.105
r30 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.205
+ $Y=1.16 $X2=2.205 $Y2=1.16
r31 7 14 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=2.245 $Y=1.175
+ $X2=2.205 $Y2=1.175
r32 4 10 45.1054 $w=3.82e-07 $l=3.02076e-07 $layer=POLY_cond $X=2.01 $Y=1.41
+ $X2=2.125 $Y2=1.16
r33 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.01 $Y=1.41 $X2=2.01
+ $Y2=1.985
r34 1 10 39.2524 $w=3.82e-07 $l=2.24332e-07 $layer=POLY_cond $X=1.985 $Y=0.995
+ $X2=2.125 $Y2=1.16
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.985 $Y=0.995
+ $X2=1.985 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_1%B1 1 3 4 6 9 15 19
r35 15 19 3.60455 $w=1.98e-07 $l=6.5e-08 $layer=LI1_cond $X=2.815 $Y=1.175
+ $X2=2.75 $Y2=1.175
r36 9 15 3.97773 $w=2e-07 $l=1.32e-07 $layer=LI1_cond $X=2.947 $Y=1.175
+ $X2=2.815 $Y2=1.175
r37 9 19 2.49545 $w=1.98e-07 $l=4.5e-08 $layer=LI1_cond $X=2.705 $Y=1.175
+ $X2=2.75 $Y2=1.175
r38 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.705
+ $Y=1.16 $X2=2.705 $Y2=1.16
r39 4 13 47.2262 $w=3.11e-07 $l=2.82843e-07 $layer=POLY_cond $X=2.65 $Y=1.41
+ $X2=2.72 $Y2=1.16
r40 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.65 $Y=1.41 $X2=2.65
+ $Y2=1.985
r41 1 13 38.532 $w=3.11e-07 $l=2.07123e-07 $layer=POLY_cond $X=2.625 $Y=0.995
+ $X2=2.72 $Y2=1.16
r42 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.625 $Y=0.995
+ $X2=2.625 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_1%C1 1 3 4 6 8 9 12 17
r29 12 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.82
+ $Y=1.16 $X2=3.82 $Y2=1.16
r30 9 17 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=3.86 $Y=1.2 $X2=3.82
+ $Y2=1.2
r31 7 12 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=3.46 $Y=1.16 $X2=3.82
+ $Y2=1.16
r32 7 8 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=3.46 $Y=1.16
+ $X2=3.36 $Y2=1.202
r33 4 8 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=3.36 $Y=1.41
+ $X2=3.36 $Y2=1.202
r34 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.36 $Y=1.41 $X2=3.36
+ $Y2=1.985
r35 1 8 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=3.335 $Y=0.995
+ $X2=3.36 $Y2=1.202
r36 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.335 $Y=0.995
+ $X2=3.335 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_1%X 1 2 10 13 14 15 16 17 22
r21 17 31 4.4064 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=0.255 $Y=2.21
+ $X2=0.255 $Y2=2.34
r22 16 17 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.255 $Y=1.87
+ $X2=0.255 $Y2=2.21
r23 15 22 4.4064 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=0.255 $Y=0.51
+ $X2=0.255 $Y2=0.38
r24 13 14 8.29786 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.255 $Y=1.66
+ $X2=0.255 $Y2=1.495
r25 11 16 6.94855 $w=3.38e-07 $l=2.05e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=1.87
r26 11 13 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=1.66
r27 10 14 38.6597 $w=1.73e-07 $l=6.1e-07 $layer=LI1_cond $X=0.172 $Y=0.885
+ $X2=0.172 $Y2=1.495
r28 9 15 6.94855 $w=3.38e-07 $l=2.05e-07 $layer=LI1_cond $X=0.255 $Y=0.715
+ $X2=0.255 $Y2=0.51
r29 9 10 8.46734 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.255 $Y=0.715
+ $X2=0.255 $Y2=0.885
r30 2 31 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r31 2 13 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r32 1 22 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_1%VPWR 1 2 3 14 18 22 26 28 30 40 41 44 47
+ 50 53
c45 2 0 1.32642e-19 $X=1.125 $Y=1.485
r46 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r47 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r48 45 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r49 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 41 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=2.99 $Y2=2.72
r51 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r52 38 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.09 $Y=2.72
+ $X2=2.925 $Y2=2.72
r53 38 40 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=3.09 $Y=2.72
+ $X2=3.91 $Y2=2.72
r54 37 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r55 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r56 34 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r57 34 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r58 33 36 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r59 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r60 31 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.21 $Y2=2.72
r61 31 33 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.61 $Y2=2.72
r62 30 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.76 $Y=2.72
+ $X2=2.925 $Y2=2.72
r63 30 36 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.76 $Y=2.72
+ $X2=2.53 $Y2=2.72
r64 28 45 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 28 53 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r66 24 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=2.635
+ $X2=2.925 $Y2=2.72
r67 24 26 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.925 $Y=2.635
+ $X2=2.925 $Y2=2
r68 20 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=2.635
+ $X2=1.21 $Y2=2.72
r69 20 22 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.21 $Y=2.635
+ $X2=1.21 $Y2=2
r70 19 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=2.72
+ $X2=0.73 $Y2=2.72
r71 18 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.085 $Y=2.72
+ $X2=1.21 $Y2=2.72
r72 18 19 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.085 $Y=2.72
+ $X2=0.815 $Y2=2.72
r73 14 17 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.73 $Y=1.66
+ $X2=0.73 $Y2=2.34
r74 12 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.72
r75 12 17 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.34
r76 3 26 300 $w=1.7e-07 $l=6.00417e-07 $layer=licon1_PDIFF $count=2 $X=2.74
+ $Y=1.485 $X2=2.925 $Y2=2
r77 2 22 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=1.125
+ $Y=1.485 $X2=1.25 $Y2=2
r78 1 17 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r79 1 14 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_1%VGND 1 2 11 15 18 19 20 30 31 34 37
r47 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r48 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r49 28 31 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=3.91
+ $Y2=0
r50 27 30 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.91
+ $Y2=0
r51 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r52 25 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r53 25 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r54 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r55 22 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.77
+ $Y2=0
r56 22 24 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.61
+ $Y2=0
r57 20 35 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r58 20 37 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r59 18 24 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.635 $Y=0 $X2=1.61
+ $Y2=0
r60 18 19 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=1.635 $Y=0 $X2=1.747
+ $Y2=0
r61 17 27 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=2.07
+ $Y2=0
r62 17 19 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=1.747
+ $Y2=0
r63 13 19 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.747 $Y=0.085
+ $X2=1.747 $Y2=0
r64 13 15 15.1098 $w=2.23e-07 $l=2.95e-07 $layer=LI1_cond $X=1.747 $Y=0.085
+ $X2=1.747 $Y2=0.38
r65 9 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=0.085
+ $X2=0.77 $Y2=0
r66 9 11 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.77 $Y=0.085
+ $X2=0.77 $Y2=0.38
r67 2 15 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.75 $Y2=0.38
r68 1 11 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_1%A_225_47# 1 2 9 11 12 15
r38 13 15 10.7662 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=2.22 $Y=0.735
+ $X2=2.22 $Y2=0.38
r39 11 13 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=2.03 $Y=0.82
+ $X2=2.22 $Y2=0.735
r40 11 12 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.03 $Y=0.82
+ $X2=1.415 $Y2=0.82
r41 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.25 $Y=0.735
+ $X2=1.415 $Y2=0.82
r42 7 9 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.25 $Y=0.735
+ $X2=1.25 $Y2=0.38
r43 2 15 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=2.06
+ $Y=0.235 $X2=2.245 $Y2=0.38
r44 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.125
+ $Y=0.235 $X2=1.25 $Y2=0.38
.ends

