* File: sky130_fd_sc_hdll__o211ai_1.spice
* Created: Wed Sep  2 08:42:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o211ai_1.pex.spice"
.subckt sky130_fd_sc_hdll__o211ai_1  VNB VPB A1 A2 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A1_M1000_g N_A_27_47#_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.20475 PD=0.98 PS=1.93 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75000.2
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1001 N_A_27_47#_M1001_d N_A2_M1001_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.09425 AS=0.10725 PD=0.94 PS=0.98 NRD=2.76 NRS=10.152 M=1 R=4.33333
+ SA=75000.7 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1007 A_304_47# N_B1_M1007_g N_A_27_47#_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.121875 AS=0.09425 PD=1.025 PS=0.94 NRD=24.456 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75001 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_C1_M1004_g A_304_47# VNB NSHORT L=0.15 W=0.65 AD=0.377
+ AS=0.121875 PD=2.46 PS=1.025 NRD=45.228 NRS=24.456 M=1 R=4.33333 SA=75001.7
+ SB=75000.5 A=0.0975 P=1.6 MULT=1
MM1005 A_118_297# N_A1_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1 AD=0.115
+ AS=0.275 PD=1.23 PS=2.55 NRD=11.8003 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90001.9 A=0.18 P=2.36 MULT=1
MM1002 N_Y_M1002_d N_A2_M1002_g A_118_297# VPB PHIGHVT L=0.18 W=1 AD=0.19
+ AS=0.115 PD=1.38 PS=1.23 NRD=3.9203 NRS=11.8003 M=1 R=5.55556 SA=90000.6
+ SB=90001.5 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_B1_M1003_g N_Y_M1002_d VPB PHIGHVT L=0.18 W=1 AD=0.1725
+ AS=0.19 PD=1.345 PS=1.38 NRD=0.9653 NRS=15.7403 M=1 R=5.55556 SA=90001.2
+ SB=90001 A=0.18 P=2.36 MULT=1
MM1006 N_Y_M1006_d N_C1_M1006_g N_VPWR_M1003_d VPB PHIGHVT L=0.18 W=1 AD=0.54
+ AS=0.1725 PD=3.08 PS=1.345 NRD=42.3353 NRS=11.8003 M=1 R=5.55556 SA=90001.7
+ SB=90000.4 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hdll__o211ai_1.pxi.spice"
*
.ends
*
*
