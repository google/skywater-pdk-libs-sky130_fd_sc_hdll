* File: sky130_fd_sc_hdll__diode_8.spice
* Created: Thu Aug 27 19:05:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__diode_8.pex.spice"
.subckt sky130_fd_sc_hdll__diode_8  VNB VPB DIODE VGND VPWR
* 
* DIODE	DIODE
* VPB	VPB
* VNB	VNB
D0_noxref VNB N_DIODE_D0_noxref_neg NDIODE  AREA=3.5464 PJ=9.74 M=1
+ AHFTEMPPERIM=9.74
DX1_noxref VNB VPB NWDIODE A=4.6956 P=12.86
*
.include "sky130_fd_sc_hdll__diode_8.pxi.spice"
*
.ends
*
*
