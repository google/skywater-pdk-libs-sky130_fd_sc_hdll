# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__probe_p_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.832500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 1.075000 1.240000 1.275000 ;
    END
  END A
  PIN VGND
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.980000 0.085000 ;
        RECT 0.615000  0.085000 0.895000 0.565000 ;
        RECT 1.505000  0.085000 1.805000 0.565000 ;
        RECT 2.475000  0.085000 2.745000 0.565000 ;
        RECT 3.415000  0.085000 3.685000 0.565000 ;
        RECT 4.355000  0.085000 4.625000 0.565000 ;
        RECT 5.295000  0.085000 5.545000 0.885000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.980000 2.805000 ;
        RECT 0.595000 1.835000 0.865000 2.635000 ;
        RECT 1.535000 1.835000 1.805000 2.635000 ;
        RECT 2.475000 1.835000 2.745000 2.635000 ;
        RECT 3.415000 1.835000 3.685000 2.635000 ;
        RECT 4.355000 1.835000 4.625000 2.635000 ;
        RECT 5.295000 1.485000 5.595000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1.250000 0.560000 4.270000 2.160000 ;
      LAYER via4 ;
        RECT 1.560000 0.870000 2.360000 1.670000 ;
        RECT 3.160000 0.870000 3.960000 1.670000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.095000 1.445000 1.595000 1.615000 ;
      RECT 0.095000 1.615000 0.425000 2.465000 ;
      RECT 0.145000 0.255000 0.445000 0.735000 ;
      RECT 0.145000 0.735000 1.595000 0.905000 ;
      RECT 1.035000 1.615000 1.365000 2.465000 ;
      RECT 1.065000 0.255000 1.335000 0.735000 ;
      RECT 1.420000 0.905000 1.595000 1.075000 ;
      RECT 1.420000 1.075000 4.045000 1.245000 ;
      RECT 1.420000 1.245000 1.595000 1.445000 ;
      RECT 1.975000 0.255000 2.305000 0.735000 ;
      RECT 1.975000 0.735000 5.125000 0.905000 ;
      RECT 1.975000 1.445000 5.125000 1.615000 ;
      RECT 1.975000 1.615000 2.305000 2.465000 ;
      RECT 2.915000 0.255000 3.245000 0.735000 ;
      RECT 2.915000 1.615000 3.245000 2.465000 ;
      RECT 3.855000 0.255000 4.185000 0.735000 ;
      RECT 3.855000 1.615000 4.185000 2.465000 ;
      RECT 4.290000 0.905000 5.125000 1.445000 ;
      RECT 4.795000 0.255000 5.125000 0.735000 ;
      RECT 4.795000 1.615000 5.125000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.560000  1.105000 4.730000 1.275000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 4.920000  1.105000 5.090000 1.275000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 3.465000 1.060000 4.105000 1.320000 ;
      RECT 4.105000 1.075000 5.150000 1.305000 ;
    LAYER met2 ;
      RECT 3.445000 1.005000 4.125000 1.375000 ;
      RECT 3.465000 1.060000 4.105000 1.320000 ;
    LAYER met3 ;
      RECT 3.395000 1.025000 3.420000 1.355000 ;
      RECT 3.395000 1.030000 4.175000 1.350000 ;
      RECT 3.420000 1.025000 4.150000 1.355000 ;
      RECT 4.150000 1.025000 4.175000 1.355000 ;
    LAYER met4 ;
      RECT 1.370000 0.680000 4.150000 1.860000 ;
      RECT 3.420000 1.025000 4.150000 1.355000 ;
    LAYER via ;
      RECT 3.550000 1.115000 3.700000 1.265000 ;
      RECT 3.870000 1.115000 4.020000 1.265000 ;
    LAYER via2 ;
      RECT 3.485000 1.090000 3.685000 1.290000 ;
      RECT 3.885000 1.090000 4.085000 1.290000 ;
    LAYER via3 ;
      RECT 3.485000 1.090000 3.685000 1.290000 ;
      RECT 3.885000 1.090000 4.085000 1.290000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__probe_p_8
