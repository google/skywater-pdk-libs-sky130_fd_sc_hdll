* File: sky130_fd_sc_hdll__or2_8.pxi.spice
* Created: Thu Aug 27 19:23:36 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR2_8%A N_A_c_106_n N_A_M1000_g N_A_c_102_n N_A_M1001_g
+ N_A_c_103_n N_A_M1004_g N_A_c_107_n N_A_M1014_g A N_A_c_104_n N_A_c_105_n A
+ PM_SKY130_FD_SC_HDLL__OR2_8%A
x_PM_SKY130_FD_SC_HDLL__OR2_8%B N_B_c_145_n N_B_M1006_g N_B_c_141_n N_B_M1012_g
+ N_B_c_142_n N_B_M1016_g N_B_c_146_n N_B_M1008_g B N_B_c_143_n N_B_c_144_n B
+ PM_SKY130_FD_SC_HDLL__OR2_8%B
x_PM_SKY130_FD_SC_HDLL__OR2_8%A_123_47# N_A_123_47#_M1001_s N_A_123_47#_M1012_d
+ N_A_123_47#_M1006_s N_A_123_47#_c_213_n N_A_123_47#_M1002_g
+ N_A_123_47#_c_196_n N_A_123_47#_M1003_g N_A_123_47#_c_197_n
+ N_A_123_47#_M1005_g N_A_123_47#_c_214_n N_A_123_47#_M1007_g
+ N_A_123_47#_c_215_n N_A_123_47#_M1009_g N_A_123_47#_c_198_n
+ N_A_123_47#_M1010_g N_A_123_47#_c_199_n N_A_123_47#_M1013_g
+ N_A_123_47#_c_216_n N_A_123_47#_M1011_g N_A_123_47#_c_217_n
+ N_A_123_47#_M1015_g N_A_123_47#_c_200_n N_A_123_47#_M1018_g
+ N_A_123_47#_c_201_n N_A_123_47#_M1021_g N_A_123_47#_c_218_n
+ N_A_123_47#_M1017_g N_A_123_47#_c_219_n N_A_123_47#_M1019_g
+ N_A_123_47#_c_202_n N_A_123_47#_M1022_g N_A_123_47#_c_203_n
+ N_A_123_47#_M1023_g N_A_123_47#_c_220_n N_A_123_47#_M1020_g
+ N_A_123_47#_c_225_n N_A_123_47#_c_204_n N_A_123_47#_c_205_n
+ N_A_123_47#_c_234_n N_A_123_47#_c_206_n N_A_123_47#_c_221_n
+ N_A_123_47#_c_207_n N_A_123_47#_c_208_n N_A_123_47#_c_209_n
+ N_A_123_47#_c_210_n N_A_123_47#_c_223_n N_A_123_47#_c_211_n
+ N_A_123_47#_c_212_n PM_SKY130_FD_SC_HDLL__OR2_8%A_123_47#
x_PM_SKY130_FD_SC_HDLL__OR2_8%A_27_297# N_A_27_297#_M1000_s N_A_27_297#_M1014_s
+ N_A_27_297#_M1008_d N_A_27_297#_c_414_n N_A_27_297#_c_415_n
+ N_A_27_297#_c_416_n N_A_27_297#_c_417_n N_A_27_297#_c_438_p
+ N_A_27_297#_c_418_n N_A_27_297#_c_419_n PM_SKY130_FD_SC_HDLL__OR2_8%A_27_297#
x_PM_SKY130_FD_SC_HDLL__OR2_8%VPWR N_VPWR_M1000_d N_VPWR_M1002_s N_VPWR_M1007_s
+ N_VPWR_M1011_s N_VPWR_M1017_s N_VPWR_M1020_s N_VPWR_c_449_n N_VPWR_c_450_n
+ N_VPWR_c_451_n N_VPWR_c_452_n N_VPWR_c_453_n N_VPWR_c_454_n N_VPWR_c_455_n
+ N_VPWR_c_456_n N_VPWR_c_457_n N_VPWR_c_458_n N_VPWR_c_459_n N_VPWR_c_460_n
+ N_VPWR_c_461_n N_VPWR_c_462_n N_VPWR_c_463_n N_VPWR_c_464_n VPWR
+ N_VPWR_c_465_n N_VPWR_c_466_n N_VPWR_c_448_n N_VPWR_c_468_n
+ PM_SKY130_FD_SC_HDLL__OR2_8%VPWR
x_PM_SKY130_FD_SC_HDLL__OR2_8%X N_X_M1003_s N_X_M1010_s N_X_M1018_s N_X_M1022_s
+ N_X_M1002_d N_X_M1009_d N_X_M1015_d N_X_M1019_d N_X_c_548_n N_X_c_549_n
+ N_X_c_553_n N_X_c_539_n N_X_c_540_n N_X_c_564_n N_X_c_568_n N_X_c_653_p
+ N_X_c_541_n N_X_c_576_n N_X_c_580_n N_X_c_656_p N_X_c_542_n N_X_c_588_n
+ N_X_c_592_n N_X_c_659_p N_X_c_595_n N_X_c_543_n N_X_c_603_n N_X_c_544_n
+ N_X_c_611_n N_X_c_545_n X PM_SKY130_FD_SC_HDLL__OR2_8%X
x_PM_SKY130_FD_SC_HDLL__OR2_8%VGND N_VGND_M1001_d N_VGND_M1004_d N_VGND_M1016_s
+ N_VGND_M1005_d N_VGND_M1013_d N_VGND_M1021_d N_VGND_M1023_d N_VGND_c_673_n
+ N_VGND_c_674_n N_VGND_c_675_n N_VGND_c_676_n N_VGND_c_677_n N_VGND_c_678_n
+ N_VGND_c_679_n N_VGND_c_680_n N_VGND_c_681_n N_VGND_c_682_n N_VGND_c_683_n
+ N_VGND_c_684_n N_VGND_c_685_n N_VGND_c_686_n N_VGND_c_687_n N_VGND_c_688_n
+ N_VGND_c_689_n VGND N_VGND_c_690_n N_VGND_c_691_n N_VGND_c_692_n
+ N_VGND_c_693_n N_VGND_c_694_n PM_SKY130_FD_SC_HDLL__OR2_8%VGND
cc_1 VNB N_A_c_102_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_2 VNB N_A_c_103_n 0.0168874f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_3 VNB N_A_c_104_n 0.00954103f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=1.16
cc_4 VNB N_A_c_105_n 0.0446632f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=1.202
cc_5 VNB N_B_c_141_n 0.0168863f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_6 VNB N_B_c_142_n 0.0192987f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_7 VNB N_B_c_143_n 0.00334669f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=1.16
cc_8 VNB N_B_c_144_n 0.0398898f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=1.202
cc_9 VNB N_A_123_47#_c_196_n 0.0196693f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_10 VNB N_A_123_47#_c_197_n 0.0167085f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.202
cc_11 VNB N_A_123_47#_c_198_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_12 VNB N_A_123_47#_c_199_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_123_47#_c_200_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_123_47#_c_201_n 0.0167199f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_123_47#_c_202_n 0.0166979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_123_47#_c_203_n 0.019415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_123_47#_c_204_n 0.00468914f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_123_47#_c_205_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_123_47#_c_206_n 0.00282074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_123_47#_c_207_n 0.00481184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_123_47#_c_208_n 8.16212e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_123_47#_c_209_n 0.015542f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_123_47#_c_210_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_123_47#_c_211_n 0.00247108f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_123_47#_c_212_n 0.159021f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_448_n 0.288713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_539_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_X_c_540_n 0.00221586f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_X_c_541_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_X_c_542_n 0.00335912f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_X_c_543_n 0.00220648f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_X_c_544_n 0.00220648f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_X_c_545_n 0.00214047f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB X 0.0157603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_673_n 0.0120163f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.175
cc_36 VNB N_VGND_c_674_n 0.00988966f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.175
cc_37 VNB N_VGND_c_675_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=1.175
cc_38 VNB N_VGND_c_676_n 0.00413904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_677_n 0.00286952f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_678_n 0.00445447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_679_n 0.00442069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_680_n 0.00442069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_681_n 0.0183517f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_682_n 0.0167328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_683_n 0.00631953f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_684_n 0.0155459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_685_n 0.00631953f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_686_n 0.0155459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_687_n 0.00631953f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_688_n 0.0155446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_689_n 0.00631953f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_690_n 0.0115308f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_691_n 0.342161f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_692_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_693_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_694_n 0.0221721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VPB N_A_c_106_n 0.0201729f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_58 VPB N_A_c_107_n 0.0159343f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_59 VPB N_A_c_105_n 0.0228641f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.202
cc_60 VPB N_B_c_145_n 0.01625f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_61 VPB N_B_c_146_n 0.0192027f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_62 VPB N_B_c_144_n 0.0203675f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.202
cc_63 VPB N_A_123_47#_c_213_n 0.0195908f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_64 VPB N_A_123_47#_c_214_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0.92 $Y2=1.16
cc_65 VPB N_A_123_47#_c_215_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.175
cc_66 VPB N_A_123_47#_c_216_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_123_47#_c_217_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_123_47#_c_218_n 0.0162627f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_123_47#_c_219_n 0.016253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_123_47#_c_220_n 0.0192858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_123_47#_c_221_n 0.0074991f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_123_47#_c_208_n 0.00391833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_123_47#_c_223_n 0.00174301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_123_47#_c_212_n 0.100092f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_297#_c_414_n 0.0154985f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_76 VPB N_A_27_297#_c_415_n 0.0313426f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.985
cc_77 VPB N_A_27_297#_c_416_n 0.00185333f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_297#_c_417_n 0.00449763f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.202
cc_79 VPB N_A_27_297#_c_418_n 0.00188991f $X=-0.19 $Y=1.305 $X2=0.92 $Y2=1.16
cc_80 VPB N_A_27_297#_c_419_n 0.00463934f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.175
cc_81 VPB N_VPWR_c_449_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_82 VPB N_VPWR_c_450_n 0.014029f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.19
cc_83 VPB N_VPWR_c_451_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_452_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_453_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_454_n 0.00472202f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_455_n 0.038808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_456_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_457_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_458_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_459_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_460_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_461_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_462_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_463_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_464_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_465_n 0.0166737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_466_n 0.0124854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_448_n 0.062942f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_468_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB X 0.00816161f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 N_A_c_107_n N_B_c_145_n 0.00966038f $X=0.985 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_103 N_A_c_103_n N_B_c_141_n 0.0179509f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A_c_104_n N_B_c_143_n 0.0115142f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_c_105_n N_B_c_143_n 2.50364e-19 $X=0.96 $Y=1.202 $X2=0 $Y2=0
cc_106 N_A_c_104_n N_B_c_144_n 2.50364e-19 $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_c_105_n N_B_c_144_n 0.0228273f $X=0.96 $Y=1.202 $X2=0 $Y2=0
cc_108 N_A_c_102_n N_A_123_47#_c_225_n 0.00539651f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_c_103_n N_A_123_47#_c_225_n 0.00671723f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_110 N_A_c_103_n N_A_123_47#_c_204_n 0.00922411f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A_c_104_n N_A_123_47#_c_204_n 0.0118735f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_c_105_n N_A_123_47#_c_204_n 0.00141784f $X=0.96 $Y=1.202 $X2=0 $Y2=0
cc_113 N_A_c_102_n N_A_123_47#_c_205_n 0.00262807f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A_c_103_n N_A_123_47#_c_205_n 0.00113286f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A_c_104_n N_A_123_47#_c_205_n 0.0265405f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_c_105_n N_A_123_47#_c_205_n 0.00230339f $X=0.96 $Y=1.202 $X2=0 $Y2=0
cc_117 N_A_c_103_n N_A_123_47#_c_234_n 5.24636e-19 $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A_c_106_n N_A_27_297#_c_416_n 0.0167211f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_c_107_n N_A_27_297#_c_416_n 0.0164317f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_c_104_n N_A_27_297#_c_416_n 0.0457717f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_c_105_n N_A_27_297#_c_416_n 0.00831613f $X=0.96 $Y=1.202 $X2=0 $Y2=0
cc_122 N_A_c_106_n N_VPWR_c_449_n 0.0127203f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A_c_107_n N_VPWR_c_449_n 0.0120006f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A_c_107_n N_VPWR_c_455_n 0.00622633f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A_c_106_n N_VPWR_c_465_n 0.00622633f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A_c_106_n N_VPWR_c_448_n 0.0113307f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A_c_107_n N_VPWR_c_448_n 0.0104264f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A_c_102_n N_VGND_c_674_n 0.00366701f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_c_102_n N_VGND_c_675_n 0.00541359f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_c_103_n N_VGND_c_675_n 0.00423334f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_c_103_n N_VGND_c_676_n 0.00166854f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_c_102_n N_VGND_c_691_n 0.0105165f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_c_103_n N_VGND_c_691_n 0.00596967f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_134 N_B_c_141_n N_A_123_47#_c_225_n 5.24636e-19 $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_135 N_B_c_141_n N_A_123_47#_c_204_n 0.00922411f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_136 N_B_c_143_n N_A_123_47#_c_204_n 0.0118735f $X=1.86 $Y=1.16 $X2=0 $Y2=0
cc_137 N_B_c_144_n N_A_123_47#_c_204_n 0.00141784f $X=1.9 $Y=1.202 $X2=0 $Y2=0
cc_138 N_B_c_141_n N_A_123_47#_c_234_n 0.00671723f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_139 N_B_c_142_n N_A_123_47#_c_234_n 0.0109565f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_140 N_B_c_142_n N_A_123_47#_c_206_n 0.0101683f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_141 N_B_c_143_n N_A_123_47#_c_206_n 0.0118215f $X=1.86 $Y=1.16 $X2=0 $Y2=0
cc_142 N_B_c_144_n N_A_123_47#_c_206_n 0.00141613f $X=1.9 $Y=1.202 $X2=0 $Y2=0
cc_143 N_B_c_146_n N_A_123_47#_c_221_n 0.0145448f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_144 N_B_c_143_n N_A_123_47#_c_221_n 0.0119049f $X=1.86 $Y=1.16 $X2=0 $Y2=0
cc_145 N_B_c_144_n N_A_123_47#_c_221_n 2.7776e-19 $X=1.9 $Y=1.202 $X2=0 $Y2=0
cc_146 N_B_c_142_n N_A_123_47#_c_207_n 0.00290689f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_147 N_B_c_144_n N_A_123_47#_c_207_n 0.00328986f $X=1.9 $Y=1.202 $X2=0 $Y2=0
cc_148 N_B_c_146_n N_A_123_47#_c_208_n 0.00118343f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_149 N_B_c_144_n N_A_123_47#_c_208_n 0.00507668f $X=1.9 $Y=1.202 $X2=0 $Y2=0
cc_150 N_B_c_141_n N_A_123_47#_c_210_n 0.00113286f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_151 N_B_c_142_n N_A_123_47#_c_210_n 0.00158032f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_152 N_B_c_143_n N_A_123_47#_c_210_n 0.0265405f $X=1.86 $Y=1.16 $X2=0 $Y2=0
cc_153 N_B_c_144_n N_A_123_47#_c_210_n 0.00230339f $X=1.9 $Y=1.202 $X2=0 $Y2=0
cc_154 N_B_c_145_n N_A_123_47#_c_223_n 0.00824242f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_155 N_B_c_146_n N_A_123_47#_c_223_n 0.0119312f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_156 N_B_c_143_n N_A_123_47#_c_223_n 0.0267279f $X=1.86 $Y=1.16 $X2=0 $Y2=0
cc_157 N_B_c_144_n N_A_123_47#_c_223_n 0.00806013f $X=1.9 $Y=1.202 $X2=0 $Y2=0
cc_158 N_B_c_143_n N_A_123_47#_c_211_n 0.0176337f $X=1.86 $Y=1.16 $X2=0 $Y2=0
cc_159 N_B_c_144_n N_A_123_47#_c_211_n 0.00155012f $X=1.9 $Y=1.202 $X2=0 $Y2=0
cc_160 N_B_c_145_n N_A_27_297#_c_417_n 2.72094e-19 $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_161 N_B_c_145_n N_A_27_297#_c_418_n 0.0137768f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_162 N_B_c_146_n N_A_27_297#_c_418_n 0.0111504f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_163 N_B_c_145_n N_VPWR_c_449_n 9.95594e-19 $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_164 N_B_c_146_n N_VPWR_c_450_n 0.00746267f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_165 N_B_c_145_n N_VPWR_c_455_n 0.00429453f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_166 N_B_c_146_n N_VPWR_c_455_n 0.00429453f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_167 N_B_c_145_n N_VPWR_c_448_n 0.00609021f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_168 N_B_c_146_n N_VPWR_c_448_n 0.00734734f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_169 N_B_c_141_n N_VGND_c_676_n 0.00166738f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_170 N_B_c_142_n N_VGND_c_677_n 0.00451653f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_171 N_B_c_141_n N_VGND_c_691_n 0.00596967f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B_c_142_n N_VGND_c_691_n 0.00705967f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_173 N_B_c_141_n N_VGND_c_693_n 0.00423334f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_174 N_B_c_142_n N_VGND_c_693_n 0.00424416f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_175 N_B_c_142_n N_VGND_c_694_n 0.00336547f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_123_47#_c_221_n N_A_27_297#_M1008_d 0.00319987f $X=2.195 $Y=1.555
+ $X2=0 $Y2=0
cc_177 N_A_123_47#_c_204_n N_A_27_297#_c_417_n 0.0101144f $X=1.525 $Y=0.815
+ $X2=0 $Y2=0
cc_178 N_A_123_47#_c_223_n N_A_27_297#_c_417_n 0.010246f $X=1.69 $Y=1.62 $X2=0
+ $Y2=0
cc_179 N_A_123_47#_M1006_s N_A_27_297#_c_418_n 0.00352392f $X=1.545 $Y=1.485
+ $X2=0 $Y2=0
cc_180 N_A_123_47#_c_221_n N_A_27_297#_c_418_n 0.00370305f $X=2.195 $Y=1.555
+ $X2=0 $Y2=0
cc_181 N_A_123_47#_c_223_n N_A_27_297#_c_418_n 0.0160463f $X=1.69 $Y=1.62 $X2=0
+ $Y2=0
cc_182 N_A_123_47#_c_221_n N_A_27_297#_c_419_n 0.021786f $X=2.195 $Y=1.555 $X2=0
+ $Y2=0
cc_183 N_A_123_47#_c_213_n N_VPWR_c_450_n 0.00354866f $X=2.915 $Y=1.41 $X2=0
+ $Y2=0
cc_184 N_A_123_47#_c_221_n N_VPWR_c_450_n 0.0148255f $X=2.195 $Y=1.555 $X2=0
+ $Y2=0
cc_185 N_A_123_47#_c_209_n N_VPWR_c_450_n 0.0169062f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_123_47#_c_214_n N_VPWR_c_451_n 0.00173895f $X=3.385 $Y=1.41 $X2=0
+ $Y2=0
cc_187 N_A_123_47#_c_215_n N_VPWR_c_451_n 0.00173895f $X=3.855 $Y=1.41 $X2=0
+ $Y2=0
cc_188 N_A_123_47#_c_216_n N_VPWR_c_452_n 0.00173895f $X=4.325 $Y=1.41 $X2=0
+ $Y2=0
cc_189 N_A_123_47#_c_217_n N_VPWR_c_452_n 0.00173895f $X=4.795 $Y=1.41 $X2=0
+ $Y2=0
cc_190 N_A_123_47#_c_218_n N_VPWR_c_453_n 0.00173895f $X=5.265 $Y=1.41 $X2=0
+ $Y2=0
cc_191 N_A_123_47#_c_219_n N_VPWR_c_453_n 0.00173895f $X=5.735 $Y=1.41 $X2=0
+ $Y2=0
cc_192 N_A_123_47#_c_220_n N_VPWR_c_454_n 0.00354866f $X=6.205 $Y=1.41 $X2=0
+ $Y2=0
cc_193 N_A_123_47#_c_213_n N_VPWR_c_457_n 0.00673617f $X=2.915 $Y=1.41 $X2=0
+ $Y2=0
cc_194 N_A_123_47#_c_214_n N_VPWR_c_457_n 0.00673617f $X=3.385 $Y=1.41 $X2=0
+ $Y2=0
cc_195 N_A_123_47#_c_215_n N_VPWR_c_459_n 0.00673617f $X=3.855 $Y=1.41 $X2=0
+ $Y2=0
cc_196 N_A_123_47#_c_216_n N_VPWR_c_459_n 0.00673617f $X=4.325 $Y=1.41 $X2=0
+ $Y2=0
cc_197 N_A_123_47#_c_217_n N_VPWR_c_461_n 0.00673617f $X=4.795 $Y=1.41 $X2=0
+ $Y2=0
cc_198 N_A_123_47#_c_218_n N_VPWR_c_461_n 0.00673617f $X=5.265 $Y=1.41 $X2=0
+ $Y2=0
cc_199 N_A_123_47#_c_219_n N_VPWR_c_463_n 0.00673617f $X=5.735 $Y=1.41 $X2=0
+ $Y2=0
cc_200 N_A_123_47#_c_220_n N_VPWR_c_463_n 0.00673617f $X=6.205 $Y=1.41 $X2=0
+ $Y2=0
cc_201 N_A_123_47#_M1006_s N_VPWR_c_448_n 0.00232895f $X=1.545 $Y=1.485 $X2=0
+ $Y2=0
cc_202 N_A_123_47#_c_213_n N_VPWR_c_448_n 0.0130007f $X=2.915 $Y=1.41 $X2=0
+ $Y2=0
cc_203 N_A_123_47#_c_214_n N_VPWR_c_448_n 0.0117184f $X=3.385 $Y=1.41 $X2=0
+ $Y2=0
cc_204 N_A_123_47#_c_215_n N_VPWR_c_448_n 0.0117184f $X=3.855 $Y=1.41 $X2=0
+ $Y2=0
cc_205 N_A_123_47#_c_216_n N_VPWR_c_448_n 0.0117184f $X=4.325 $Y=1.41 $X2=0
+ $Y2=0
cc_206 N_A_123_47#_c_217_n N_VPWR_c_448_n 0.0117184f $X=4.795 $Y=1.41 $X2=0
+ $Y2=0
cc_207 N_A_123_47#_c_218_n N_VPWR_c_448_n 0.0117184f $X=5.265 $Y=1.41 $X2=0
+ $Y2=0
cc_208 N_A_123_47#_c_219_n N_VPWR_c_448_n 0.0117184f $X=5.735 $Y=1.41 $X2=0
+ $Y2=0
cc_209 N_A_123_47#_c_220_n N_VPWR_c_448_n 0.0127698f $X=6.205 $Y=1.41 $X2=0
+ $Y2=0
cc_210 N_A_123_47#_c_196_n N_X_c_548_n 0.00538045f $X=2.94 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A_123_47#_c_213_n N_X_c_549_n 0.00220007f $X=2.915 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A_123_47#_c_214_n N_X_c_549_n 6.2e-19 $X=3.385 $Y=1.41 $X2=0 $Y2=0
cc_213 N_A_123_47#_c_209_n N_X_c_549_n 0.017187f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_214 N_A_123_47#_c_212_n N_X_c_549_n 0.006857f $X=6.18 $Y=1.202 $X2=0 $Y2=0
cc_215 N_A_123_47#_c_213_n N_X_c_553_n 0.00897418f $X=2.915 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A_123_47#_c_214_n N_X_c_553_n 0.0100233f $X=3.385 $Y=1.41 $X2=0 $Y2=0
cc_217 N_A_123_47#_c_215_n N_X_c_553_n 5.91934e-19 $X=3.855 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A_123_47#_c_197_n N_X_c_539_n 0.0109667f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A_123_47#_c_198_n N_X_c_539_n 0.0109667f $X=3.88 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_123_47#_c_209_n N_X_c_539_n 0.0475176f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A_123_47#_c_212_n N_X_c_539_n 0.00468948f $X=6.18 $Y=1.202 $X2=0 $Y2=0
cc_222 N_A_123_47#_c_196_n N_X_c_540_n 0.00262807f $X=2.94 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A_123_47#_c_197_n N_X_c_540_n 2.083e-19 $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A_123_47#_c_209_n N_X_c_540_n 0.0242381f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_225 N_A_123_47#_c_212_n N_X_c_540_n 0.00230339f $X=6.18 $Y=1.202 $X2=0 $Y2=0
cc_226 N_A_123_47#_c_214_n N_X_c_564_n 0.0141085f $X=3.385 $Y=1.41 $X2=0 $Y2=0
cc_227 N_A_123_47#_c_215_n N_X_c_564_n 0.0141085f $X=3.855 $Y=1.41 $X2=0 $Y2=0
cc_228 N_A_123_47#_c_209_n N_X_c_564_n 0.0312997f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A_123_47#_c_212_n N_X_c_564_n 0.00626531f $X=6.18 $Y=1.202 $X2=0 $Y2=0
cc_230 N_A_123_47#_c_214_n N_X_c_568_n 5.91934e-19 $X=3.385 $Y=1.41 $X2=0 $Y2=0
cc_231 N_A_123_47#_c_215_n N_X_c_568_n 0.0100233f $X=3.855 $Y=1.41 $X2=0 $Y2=0
cc_232 N_A_123_47#_c_216_n N_X_c_568_n 0.0100233f $X=4.325 $Y=1.41 $X2=0 $Y2=0
cc_233 N_A_123_47#_c_217_n N_X_c_568_n 5.91934e-19 $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_234 N_A_123_47#_c_199_n N_X_c_541_n 0.0109667f $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A_123_47#_c_200_n N_X_c_541_n 0.0109667f $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A_123_47#_c_209_n N_X_c_541_n 0.0475176f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A_123_47#_c_212_n N_X_c_541_n 0.00468948f $X=6.18 $Y=1.202 $X2=0 $Y2=0
cc_238 N_A_123_47#_c_216_n N_X_c_576_n 0.0141085f $X=4.325 $Y=1.41 $X2=0 $Y2=0
cc_239 N_A_123_47#_c_217_n N_X_c_576_n 0.0141085f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_240 N_A_123_47#_c_209_n N_X_c_576_n 0.0312997f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A_123_47#_c_212_n N_X_c_576_n 0.00626531f $X=6.18 $Y=1.202 $X2=0 $Y2=0
cc_242 N_A_123_47#_c_216_n N_X_c_580_n 5.91934e-19 $X=4.325 $Y=1.41 $X2=0 $Y2=0
cc_243 N_A_123_47#_c_217_n N_X_c_580_n 0.0100233f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_244 N_A_123_47#_c_218_n N_X_c_580_n 0.0100233f $X=5.265 $Y=1.41 $X2=0 $Y2=0
cc_245 N_A_123_47#_c_219_n N_X_c_580_n 5.91934e-19 $X=5.735 $Y=1.41 $X2=0 $Y2=0
cc_246 N_A_123_47#_c_201_n N_X_c_542_n 0.0109667f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A_123_47#_c_202_n N_X_c_542_n 0.0128442f $X=5.76 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A_123_47#_c_209_n N_X_c_542_n 0.0255764f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_249 N_A_123_47#_c_212_n N_X_c_542_n 0.0050384f $X=6.18 $Y=1.202 $X2=0 $Y2=0
cc_250 N_A_123_47#_c_218_n N_X_c_588_n 0.0141085f $X=5.265 $Y=1.41 $X2=0 $Y2=0
cc_251 N_A_123_47#_c_219_n N_X_c_588_n 0.0158202f $X=5.735 $Y=1.41 $X2=0 $Y2=0
cc_252 N_A_123_47#_c_209_n N_X_c_588_n 0.017107f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_253 N_A_123_47#_c_212_n N_X_c_588_n 0.00649693f $X=6.18 $Y=1.202 $X2=0 $Y2=0
cc_254 N_A_123_47#_c_218_n N_X_c_592_n 5.91934e-19 $X=5.265 $Y=1.41 $X2=0 $Y2=0
cc_255 N_A_123_47#_c_219_n N_X_c_592_n 0.0100233f $X=5.735 $Y=1.41 $X2=0 $Y2=0
cc_256 N_A_123_47#_c_220_n N_X_c_592_n 0.0144287f $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_257 N_A_123_47#_c_215_n N_X_c_595_n 6.2e-19 $X=3.855 $Y=1.41 $X2=0 $Y2=0
cc_258 N_A_123_47#_c_216_n N_X_c_595_n 6.2e-19 $X=4.325 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A_123_47#_c_209_n N_X_c_595_n 0.017187f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_260 N_A_123_47#_c_212_n N_X_c_595_n 0.006857f $X=6.18 $Y=1.202 $X2=0 $Y2=0
cc_261 N_A_123_47#_c_198_n N_X_c_543_n 2.19873e-19 $X=3.88 $Y=0.995 $X2=0 $Y2=0
cc_262 N_A_123_47#_c_199_n N_X_c_543_n 2.19873e-19 $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A_123_47#_c_209_n N_X_c_543_n 0.0219356f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A_123_47#_c_212_n N_X_c_543_n 0.00230339f $X=6.18 $Y=1.202 $X2=0 $Y2=0
cc_265 N_A_123_47#_c_217_n N_X_c_603_n 6.2e-19 $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A_123_47#_c_218_n N_X_c_603_n 6.2e-19 $X=5.265 $Y=1.41 $X2=0 $Y2=0
cc_267 N_A_123_47#_c_209_n N_X_c_603_n 0.017187f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_268 N_A_123_47#_c_212_n N_X_c_603_n 0.006857f $X=6.18 $Y=1.202 $X2=0 $Y2=0
cc_269 N_A_123_47#_c_200_n N_X_c_544_n 2.19873e-19 $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_270 N_A_123_47#_c_201_n N_X_c_544_n 2.19873e-19 $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A_123_47#_c_209_n N_X_c_544_n 0.0219356f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_272 N_A_123_47#_c_212_n N_X_c_544_n 0.00230339f $X=6.18 $Y=1.202 $X2=0 $Y2=0
cc_273 N_A_123_47#_c_219_n N_X_c_611_n 8.06138e-19 $X=5.735 $Y=1.41 $X2=0 $Y2=0
cc_274 N_A_123_47#_c_220_n N_X_c_611_n 0.0136833f $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_275 N_A_123_47#_c_212_n N_X_c_611_n 0.00285622f $X=6.18 $Y=1.202 $X2=0 $Y2=0
cc_276 N_A_123_47#_c_202_n N_X_c_545_n 2.0357e-19 $X=5.76 $Y=0.995 $X2=0 $Y2=0
cc_277 N_A_123_47#_c_203_n N_X_c_545_n 0.00935833f $X=6.18 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A_123_47#_c_212_n N_X_c_545_n 3.22957e-19 $X=6.18 $Y=1.202 $X2=0 $Y2=0
cc_279 N_A_123_47#_c_219_n X 9.26126e-19 $X=5.735 $Y=1.41 $X2=0 $Y2=0
cc_280 N_A_123_47#_c_202_n X 0.00105608f $X=5.76 $Y=0.995 $X2=0 $Y2=0
cc_281 N_A_123_47#_c_203_n X 0.00349337f $X=6.18 $Y=0.995 $X2=0 $Y2=0
cc_282 N_A_123_47#_c_220_n X 0.00339336f $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_283 N_A_123_47#_c_209_n X 0.00785868f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_284 N_A_123_47#_c_212_n X 0.040587f $X=6.18 $Y=1.202 $X2=0 $Y2=0
cc_285 N_A_123_47#_c_204_n N_VGND_M1004_d 0.00274794f $X=1.525 $Y=0.815 $X2=0
+ $Y2=0
cc_286 N_A_123_47#_c_206_n N_VGND_M1016_s 0.00701263f $X=2.195 $Y=0.82 $X2=0
+ $Y2=0
cc_287 N_A_123_47#_c_205_n N_VGND_c_674_n 0.00835241f $X=0.915 $Y=0.815 $X2=0
+ $Y2=0
cc_288 N_A_123_47#_c_225_n N_VGND_c_675_n 0.0188551f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_289 N_A_123_47#_c_204_n N_VGND_c_675_n 0.00198695f $X=1.525 $Y=0.815 $X2=0
+ $Y2=0
cc_290 N_A_123_47#_c_204_n N_VGND_c_676_n 0.0201123f $X=1.525 $Y=0.815 $X2=0
+ $Y2=0
cc_291 N_A_123_47#_c_196_n N_VGND_c_677_n 4.44251e-19 $X=2.94 $Y=0.995 $X2=0
+ $Y2=0
cc_292 N_A_123_47#_c_206_n N_VGND_c_677_n 0.0143404f $X=2.195 $Y=0.82 $X2=0
+ $Y2=0
cc_293 N_A_123_47#_c_209_n N_VGND_c_677_n 0.0217006f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_294 N_A_123_47#_c_197_n N_VGND_c_678_n 0.00179446f $X=3.36 $Y=0.995 $X2=0
+ $Y2=0
cc_295 N_A_123_47#_c_198_n N_VGND_c_678_n 0.00175624f $X=3.88 $Y=0.995 $X2=0
+ $Y2=0
cc_296 N_A_123_47#_c_199_n N_VGND_c_679_n 0.00175624f $X=4.3 $Y=0.995 $X2=0
+ $Y2=0
cc_297 N_A_123_47#_c_200_n N_VGND_c_679_n 0.00175624f $X=4.82 $Y=0.995 $X2=0
+ $Y2=0
cc_298 N_A_123_47#_c_201_n N_VGND_c_680_n 0.00175624f $X=5.24 $Y=0.995 $X2=0
+ $Y2=0
cc_299 N_A_123_47#_c_202_n N_VGND_c_680_n 0.00175624f $X=5.76 $Y=0.995 $X2=0
+ $Y2=0
cc_300 N_A_123_47#_c_203_n N_VGND_c_681_n 0.00337638f $X=6.18 $Y=0.995 $X2=0
+ $Y2=0
cc_301 N_A_123_47#_c_196_n N_VGND_c_682_n 0.00541359f $X=2.94 $Y=0.995 $X2=0
+ $Y2=0
cc_302 N_A_123_47#_c_197_n N_VGND_c_682_n 0.00437852f $X=3.36 $Y=0.995 $X2=0
+ $Y2=0
cc_303 N_A_123_47#_c_198_n N_VGND_c_684_n 0.00437852f $X=3.88 $Y=0.995 $X2=0
+ $Y2=0
cc_304 N_A_123_47#_c_199_n N_VGND_c_684_n 0.00437852f $X=4.3 $Y=0.995 $X2=0
+ $Y2=0
cc_305 N_A_123_47#_c_200_n N_VGND_c_686_n 0.00437852f $X=4.82 $Y=0.995 $X2=0
+ $Y2=0
cc_306 N_A_123_47#_c_201_n N_VGND_c_686_n 0.00437852f $X=5.24 $Y=0.995 $X2=0
+ $Y2=0
cc_307 N_A_123_47#_c_202_n N_VGND_c_688_n 0.00437852f $X=5.76 $Y=0.995 $X2=0
+ $Y2=0
cc_308 N_A_123_47#_c_203_n N_VGND_c_688_n 0.00437716f $X=6.18 $Y=0.995 $X2=0
+ $Y2=0
cc_309 N_A_123_47#_M1001_s N_VGND_c_691_n 0.00215201f $X=0.615 $Y=0.235 $X2=0
+ $Y2=0
cc_310 N_A_123_47#_M1012_d N_VGND_c_691_n 0.00215201f $X=1.555 $Y=0.235 $X2=0
+ $Y2=0
cc_311 N_A_123_47#_c_196_n N_VGND_c_691_n 0.0108251f $X=2.94 $Y=0.995 $X2=0
+ $Y2=0
cc_312 N_A_123_47#_c_197_n N_VGND_c_691_n 0.00605375f $X=3.36 $Y=0.995 $X2=0
+ $Y2=0
cc_313 N_A_123_47#_c_198_n N_VGND_c_691_n 0.00605375f $X=3.88 $Y=0.995 $X2=0
+ $Y2=0
cc_314 N_A_123_47#_c_199_n N_VGND_c_691_n 0.00605375f $X=4.3 $Y=0.995 $X2=0
+ $Y2=0
cc_315 N_A_123_47#_c_200_n N_VGND_c_691_n 0.00605375f $X=4.82 $Y=0.995 $X2=0
+ $Y2=0
cc_316 N_A_123_47#_c_201_n N_VGND_c_691_n 0.00605375f $X=5.24 $Y=0.995 $X2=0
+ $Y2=0
cc_317 N_A_123_47#_c_202_n N_VGND_c_691_n 0.00605375f $X=5.76 $Y=0.995 $X2=0
+ $Y2=0
cc_318 N_A_123_47#_c_203_n N_VGND_c_691_n 0.00693179f $X=6.18 $Y=0.995 $X2=0
+ $Y2=0
cc_319 N_A_123_47#_c_225_n N_VGND_c_691_n 0.0122069f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_320 N_A_123_47#_c_204_n N_VGND_c_691_n 0.00874058f $X=1.525 $Y=0.815 $X2=0
+ $Y2=0
cc_321 N_A_123_47#_c_234_n N_VGND_c_691_n 0.0122069f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_322 N_A_123_47#_c_206_n N_VGND_c_691_n 0.00523777f $X=2.195 $Y=0.82 $X2=0
+ $Y2=0
cc_323 N_A_123_47#_c_204_n N_VGND_c_693_n 0.00198695f $X=1.525 $Y=0.815 $X2=0
+ $Y2=0
cc_324 N_A_123_47#_c_234_n N_VGND_c_693_n 0.0188551f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_325 N_A_123_47#_c_206_n N_VGND_c_693_n 0.00193763f $X=2.195 $Y=0.82 $X2=0
+ $Y2=0
cc_326 N_A_123_47#_c_196_n N_VGND_c_694_n 0.00332573f $X=2.94 $Y=0.995 $X2=0
+ $Y2=0
cc_327 N_A_123_47#_c_206_n N_VGND_c_694_n 0.0268543f $X=2.195 $Y=0.82 $X2=0
+ $Y2=0
cc_328 N_A_123_47#_c_209_n N_VGND_c_694_n 0.00634565f $X=5.36 $Y=1.16 $X2=0
+ $Y2=0
cc_329 N_A_27_297#_c_416_n N_VPWR_M1000_d 0.00188315f $X=1.085 $Y=1.56 $X2=-0.19
+ $Y2=1.305
cc_330 N_A_27_297#_c_416_n N_VPWR_c_449_n 0.0173789f $X=1.085 $Y=1.56 $X2=0
+ $Y2=0
cc_331 N_A_27_297#_c_418_n N_VPWR_c_450_n 0.0123662f $X=2.025 $Y=2.38 $X2=0
+ $Y2=0
cc_332 N_A_27_297#_c_419_n N_VPWR_c_450_n 0.03124f $X=2.16 $Y=2 $X2=0 $Y2=0
cc_333 N_A_27_297#_c_438_p N_VPWR_c_455_n 0.0157117f $X=1.22 $Y=2.295 $X2=0
+ $Y2=0
cc_334 N_A_27_297#_c_418_n N_VPWR_c_455_n 0.0573901f $X=2.025 $Y=2.38 $X2=0
+ $Y2=0
cc_335 N_A_27_297#_c_415_n N_VPWR_c_465_n 0.0211714f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_336 N_A_27_297#_M1000_s N_VPWR_c_448_n 0.00268629f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_337 N_A_27_297#_M1014_s N_VPWR_c_448_n 0.00262506f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_338 N_A_27_297#_M1008_d N_VPWR_c_448_n 0.00217518f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_339 N_A_27_297#_c_415_n N_VPWR_c_448_n 0.0124393f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_340 N_A_27_297#_c_438_p N_VPWR_c_448_n 0.0103877f $X=1.22 $Y=2.295 $X2=0
+ $Y2=0
cc_341 N_A_27_297#_c_418_n N_VPWR_c_448_n 0.0347001f $X=2.025 $Y=2.38 $X2=0
+ $Y2=0
cc_342 N_A_27_297#_c_414_n N_VGND_c_674_n 0.0110621f $X=0.252 $Y=1.665 $X2=0
+ $Y2=0
cc_343 N_VPWR_c_448_n N_X_M1002_d 0.00231261f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_344 N_VPWR_c_448_n N_X_M1009_d 0.00231261f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_345 N_VPWR_c_448_n N_X_M1015_d 0.00231261f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_346 N_VPWR_c_448_n N_X_M1019_d 0.00231261f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_347 N_VPWR_c_457_n N_X_c_553_n 0.0189467f $X=3.485 $Y=2.72 $X2=0 $Y2=0
cc_348 N_VPWR_c_448_n N_X_c_553_n 0.0123132f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_349 N_VPWR_M1007_s N_X_c_564_n 0.00349981f $X=3.475 $Y=1.485 $X2=0 $Y2=0
cc_350 N_VPWR_c_451_n N_X_c_564_n 0.0143191f $X=3.62 $Y=2 $X2=0 $Y2=0
cc_351 N_VPWR_c_459_n N_X_c_568_n 0.0189467f $X=4.425 $Y=2.72 $X2=0 $Y2=0
cc_352 N_VPWR_c_448_n N_X_c_568_n 0.0123132f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_353 N_VPWR_M1011_s N_X_c_576_n 0.00349981f $X=4.415 $Y=1.485 $X2=0 $Y2=0
cc_354 N_VPWR_c_452_n N_X_c_576_n 0.0143191f $X=4.56 $Y=2 $X2=0 $Y2=0
cc_355 N_VPWR_c_461_n N_X_c_580_n 0.0189467f $X=5.365 $Y=2.72 $X2=0 $Y2=0
cc_356 N_VPWR_c_448_n N_X_c_580_n 0.0123132f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_357 N_VPWR_M1017_s N_X_c_588_n 0.00374786f $X=5.355 $Y=1.485 $X2=0 $Y2=0
cc_358 N_VPWR_c_453_n N_X_c_588_n 0.0143191f $X=5.5 $Y=2 $X2=0 $Y2=0
cc_359 N_VPWR_c_463_n N_X_c_592_n 0.0189467f $X=6.305 $Y=2.72 $X2=0 $Y2=0
cc_360 N_VPWR_c_448_n N_X_c_592_n 0.0123132f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_361 N_X_c_539_n N_VGND_M1005_d 0.00274794f $X=3.955 $Y=0.815 $X2=0 $Y2=0
cc_362 N_X_c_541_n N_VGND_M1013_d 0.00274794f $X=4.895 $Y=0.815 $X2=0 $Y2=0
cc_363 N_X_c_542_n N_VGND_M1021_d 0.00274794f $X=5.835 $Y=0.815 $X2=0 $Y2=0
cc_364 N_X_c_545_n N_VGND_M1023_d 0.00746601f $X=6.085 $Y=0.815 $X2=0 $Y2=0
cc_365 N_X_c_540_n N_VGND_c_677_n 0.00835241f $X=3.285 $Y=0.815 $X2=0 $Y2=0
cc_366 N_X_c_539_n N_VGND_c_678_n 0.0201123f $X=3.955 $Y=0.815 $X2=0 $Y2=0
cc_367 N_X_c_541_n N_VGND_c_679_n 0.0201123f $X=4.895 $Y=0.815 $X2=0 $Y2=0
cc_368 N_X_c_542_n N_VGND_c_680_n 0.0201123f $X=5.835 $Y=0.815 $X2=0 $Y2=0
cc_369 N_X_c_545_n N_VGND_c_681_n 0.00198903f $X=6.085 $Y=0.815 $X2=0 $Y2=0
cc_370 N_X_c_548_n N_VGND_c_682_n 0.0168814f $X=3.15 $Y=0.42 $X2=0 $Y2=0
cc_371 N_X_c_539_n N_VGND_c_682_n 0.00215746f $X=3.955 $Y=0.815 $X2=0 $Y2=0
cc_372 N_X_c_539_n N_VGND_c_684_n 0.00215746f $X=3.955 $Y=0.815 $X2=0 $Y2=0
cc_373 N_X_c_653_p N_VGND_c_684_n 0.0149077f $X=4.09 $Y=0.42 $X2=0 $Y2=0
cc_374 N_X_c_541_n N_VGND_c_684_n 0.00215746f $X=4.895 $Y=0.815 $X2=0 $Y2=0
cc_375 N_X_c_541_n N_VGND_c_686_n 0.00215746f $X=4.895 $Y=0.815 $X2=0 $Y2=0
cc_376 N_X_c_656_p N_VGND_c_686_n 0.0149077f $X=5.03 $Y=0.42 $X2=0 $Y2=0
cc_377 N_X_c_542_n N_VGND_c_686_n 0.00215746f $X=5.835 $Y=0.815 $X2=0 $Y2=0
cc_378 N_X_c_542_n N_VGND_c_688_n 0.00215746f $X=5.835 $Y=0.815 $X2=0 $Y2=0
cc_379 N_X_c_659_p N_VGND_c_688_n 0.0149339f $X=5.97 $Y=0.42 $X2=0 $Y2=0
cc_380 N_X_c_545_n N_VGND_c_688_n 0.00235405f $X=6.085 $Y=0.815 $X2=0 $Y2=0
cc_381 N_X_M1003_s N_VGND_c_691_n 0.00215201f $X=3.015 $Y=0.235 $X2=0 $Y2=0
cc_382 N_X_M1010_s N_VGND_c_691_n 0.00215201f $X=3.955 $Y=0.235 $X2=0 $Y2=0
cc_383 N_X_M1018_s N_VGND_c_691_n 0.00215201f $X=4.895 $Y=0.235 $X2=0 $Y2=0
cc_384 N_X_M1022_s N_VGND_c_691_n 0.00215201f $X=5.835 $Y=0.235 $X2=0 $Y2=0
cc_385 N_X_c_548_n N_VGND_c_691_n 0.0112579f $X=3.15 $Y=0.42 $X2=0 $Y2=0
cc_386 N_X_c_539_n N_VGND_c_691_n 0.00863654f $X=3.955 $Y=0.815 $X2=0 $Y2=0
cc_387 N_X_c_653_p N_VGND_c_691_n 0.0103089f $X=4.09 $Y=0.42 $X2=0 $Y2=0
cc_388 N_X_c_541_n N_VGND_c_691_n 0.00863654f $X=4.895 $Y=0.815 $X2=0 $Y2=0
cc_389 N_X_c_656_p N_VGND_c_691_n 0.0103089f $X=5.03 $Y=0.42 $X2=0 $Y2=0
cc_390 N_X_c_542_n N_VGND_c_691_n 0.00863654f $X=5.835 $Y=0.815 $X2=0 $Y2=0
cc_391 N_X_c_659_p N_VGND_c_691_n 0.0103166f $X=5.97 $Y=0.42 $X2=0 $Y2=0
cc_392 N_X_c_545_n N_VGND_c_691_n 0.00421024f $X=6.085 $Y=0.815 $X2=0 $Y2=0
