* File: sky130_fd_sc_hdll__xnor2_2.spice
* Created: Thu Aug 27 19:29:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__xnor2_2.pex.spice"
.subckt sky130_fd_sc_hdll__xnor2_2  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1007 N_A_27_47#_M1007_d N_B_M1007_g N_A_27_297#_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.17875 AS=0.12025 PD=1.85 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1017 N_A_27_47#_M1017_d N_B_M1017_g N_A_27_297#_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1002 N_A_27_47#_M1017_d N_A_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1003 N_A_27_47#_M1003_d N_A_M1003_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2145 AS=0.104 PD=1.96 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A_M1011_g N_A_600_47#_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.12025 PD=1.86 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1018_d N_A_M1018_g N_A_600_47#_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1018_d N_B_M1004_g N_A_600_47#_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.131625 PD=0.92 PS=1.055 NRD=0 NRS=14.76 M=1 R=4.33333
+ SA=75001.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1014_d N_B_M1014_g N_A_600_47#_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.131625 PD=1.82 PS=1.055 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_Y_M1001_d N_A_27_297#_M1001_g N_A_600_47#_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1013 N_Y_M1013_d N_A_27_297#_M1013_g N_A_600_47#_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=17.532 M=1 R=4.33333
+ SA=75000.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_B_M1005_g N_A_27_297#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.285 PD=1.29 PS=2.57 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1016 N_VPWR_M1005_d N_B_M1016_g N_A_27_297#_M1016_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1009 N_A_27_297#_M1016_s N_A_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1012 N_A_27_297#_M1012_d N_A_M1012_g N_VPWR_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.29 AS=0.145 PD=2.58 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1000 N_A_514_297#_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.29 AS=0.145 PD=2.58 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1006 N_A_514_297#_M1006_d N_A_M1006_g N_VPWR_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1015 N_Y_M1015_d N_B_M1015_g N_A_514_297#_M1006_d VPB PHIGHVT L=0.18 W=1
+ AD=0.1625 AS=0.145 PD=1.325 PS=1.29 NRD=7.8603 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1019 N_Y_M1015_d N_B_M1019_g N_A_514_297#_M1019_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1625 AS=0.27 PD=1.325 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A_27_297#_M1008_g N_Y_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1010_d N_A_27_297#_M1010_g N_Y_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.29 AS=0.145 PD=2.58 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.9461 P=16.85
*
.include "sky130_fd_sc_hdll__xnor2_2.pxi.spice"
*
.ends
*
*
