* File: sky130_fd_sc_hdll__and4b_2.pex.spice
* Created: Wed Sep  2 08:23:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND4B_2%A_N 2 3 5 8 10 11 12 21
r33 20 21 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r34 17 20 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.495 $Y2=1.16
r35 11 12 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.16
+ $X2=0.235 $Y2=1.53
r36 11 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r37 10 11 17.1909 $w=1.98e-07 $l=3.1e-07 $layer=LI1_cond $X=0.235 $Y=0.85
+ $X2=0.235 $Y2=1.16
r38 6 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.16
r39 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r40 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r41 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.89 $X2=0.495
+ $Y2=1.99
r42 1 20 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r43 1 2 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_2%A_27_413# 1 2 7 8 9 11 12 14 16 19 21 22
+ 24 26 28 34
r66 35 37 64.3271 $w=2.66e-07 $l=3.55e-07 $layer=POLY_cond $X=0.965 $Y=1.16
+ $X2=0.965 $Y2=0.805
r67 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r68 31 34 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=0.77 $Y=1.16
+ $X2=0.94 $Y2=1.16
r69 28 30 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=0.42
+ $X2=0.75 $Y2=0.585
r70 25 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=1.325
+ $X2=0.77 $Y2=1.16
r71 25 26 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=0.77 $Y=1.325
+ $X2=0.77 $Y2=1.83
r72 24 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=0.995
+ $X2=0.77 $Y2=1.16
r73 24 30 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=0.77 $Y=0.995
+ $X2=0.77 $Y2=0.585
r74 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.685 $Y=1.915
+ $X2=0.77 $Y2=1.83
r75 21 22 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.685 $Y=1.915
+ $X2=0.345 $Y2=1.915
r76 17 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=2
+ $X2=0.345 $Y2=1.915
r77 17 19 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.26 $Y=2 $X2=0.26
+ $Y2=2.3
r78 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.51 $Y=0.73 $X2=1.51
+ $Y2=0.445
r79 13 37 16.1576 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.125 $Y=0.805
+ $X2=0.965 $Y2=0.805
r80 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.435 $Y=0.805
+ $X2=1.51 $Y2=0.73
r81 12 13 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=1.435 $Y=0.805
+ $X2=1.125 $Y2=0.805
r82 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.965 $Y=1.99
+ $X2=0.965 $Y2=2.275
r83 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.89 $X2=0.965
+ $Y2=1.99
r84 7 35 32.9756 $w=2.66e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.325
+ $X2=0.965 $Y2=1.16
r85 7 8 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.965 $Y=1.325
+ $X2=0.965 $Y2=1.89
r86 2 19 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
r87 1 28 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_2%B 3 6 7 9 10 13 14 15 16 17 23
r39 16 17 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=2.025 $Y=1.19
+ $X2=2.025 $Y2=1.53
r40 16 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.98
+ $Y=1.24 $X2=1.98 $Y2=1.24
r41 15 16 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=2.025 $Y=0.85
+ $X2=2.025 $Y2=1.19
r42 14 15 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=2.025 $Y=0.51
+ $X2=2.025 $Y2=0.85
r43 12 23 82.2043 $w=2.7e-07 $l=3.7e-07 $layer=POLY_cond $X=1.98 $Y=1.61
+ $X2=1.98 $Y2=1.24
r44 12 13 34.1495 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=1.98 $Y=1.61
+ $X2=1.98 $Y2=1.745
r45 10 23 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=1.98 $Y=1.21 $X2=1.98
+ $Y2=1.24
r46 10 11 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=1.98 $Y=1.21
+ $X2=1.98 $Y2=1.075
r47 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.945 $Y=1.99
+ $X2=1.945 $Y2=2.275
r48 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.945 $Y=1.89 $X2=1.945
+ $Y2=1.99
r49 6 13 48.0787 $w=2e-07 $l=1.45e-07 $layer=POLY_cond $X=1.945 $Y=1.89
+ $X2=1.945 $Y2=1.745
r50 3 11 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.92 $Y=0.445
+ $X2=1.92 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_2%C 2 3 5 8 10 11 12 13 19
r43 19 22 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.46 $Y=1.16
+ $X2=2.46 $Y2=1.325
r44 19 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.46 $Y=1.16
+ $X2=2.46 $Y2=0.995
r45 12 13 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.495 $Y=0.85
+ $X2=2.495 $Y2=0.51
r46 11 12 14.8857 $w=2.38e-07 $l=3.1e-07 $layer=LI1_cond $X=2.495 $Y=1.16
+ $X2=2.495 $Y2=0.85
r47 11 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.46
+ $Y=1.16 $X2=2.46 $Y2=1.16
r48 10 11 16.0862 $w=2.38e-07 $l=3.35e-07 $layer=LI1_cond $X=2.495 $Y=1.495
+ $X2=2.495 $Y2=1.16
r49 8 21 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.52 $Y=0.445
+ $X2=2.52 $Y2=0.995
r50 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.495 $Y=1.99
+ $X2=2.495 $Y2=2.275
r51 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.495 $Y=1.89 $X2=2.495
+ $Y2=1.99
r52 2 22 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=2.495 $Y=1.89
+ $X2=2.495 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_2%D 2 3 5 8 10 11 12 17
c47 17 0 3.39525e-19 $X=2.955 $Y=1.16
c48 8 0 1.96288e-19 $X=3.015 $Y=0.445
r49 17 20 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.955 $Y=1.16
+ $X2=2.955 $Y2=1.325
r50 17 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.955 $Y=1.16
+ $X2=2.955 $Y2=0.995
r51 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.95 $Y=1.16
+ $X2=2.95 $Y2=1.53
r52 11 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.955
+ $Y=1.16 $X2=2.955 $Y2=1.16
r53 10 11 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.95 $Y=0.85 $X2=2.95
+ $Y2=1.16
r54 8 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.015 $Y=0.445
+ $X2=3.015 $Y2=0.995
r55 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.99 $Y=1.99 $X2=2.99
+ $Y2=2.275
r56 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.99 $Y=1.89 $X2=2.99
+ $Y2=1.99
r57 2 20 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=2.99 $Y=1.89 $X2=2.99
+ $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_2%A_211_413# 1 2 3 10 12 13 15 16 18 19 21
+ 24 28 30 32 34 37 38 39 42 50 56
c118 34 0 1.10344e-19 $X=3.295 $Y=1.88
c119 30 0 1.684e-19 $X=2.765 $Y=2.085
r120 56 57 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=4.045 $Y=1.202
+ $X2=4.07 $Y2=1.202
r121 55 56 62.3612 $w=3.71e-07 $l=4.8e-07 $layer=POLY_cond $X=3.565 $Y=1.202
+ $X2=4.045 $Y2=1.202
r122 54 55 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=3.54 $Y=1.202
+ $X2=3.565 $Y2=1.202
r123 51 54 9.09434 $w=3.71e-07 $l=7e-08 $layer=POLY_cond $X=3.47 $Y=1.202
+ $X2=3.54 $Y2=1.202
r124 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.47
+ $Y=1.16 $X2=3.47 $Y2=1.16
r125 47 50 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.38 $Y=1.16 $X2=3.47
+ $Y2=1.16
r126 45 46 8.0884 $w=1.81e-07 $l=1.2e-07 $layer=LI1_cond $X=2.765 $Y=1.88
+ $X2=2.765 $Y2=2
r127 42 44 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0.42
+ $X2=1.305 $Y2=0.585
r128 39 44 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=1.33 $Y=1.66
+ $X2=1.33 $Y2=0.585
r129 38 40 5.41145 $w=2.98e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=2
+ $X2=1.265 $Y2=2.085
r130 38 39 15.2072 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=1.265 $Y=2
+ $X2=1.265 $Y2=1.66
r131 36 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.38 $Y=1.325
+ $X2=3.38 $Y2=1.16
r132 36 37 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=3.38 $Y=1.325
+ $X2=3.38 $Y2=1.795
r133 35 45 1.09592 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.86 $Y=1.88
+ $X2=2.765 $Y2=1.88
r134 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.295 $Y=1.88
+ $X2=3.38 $Y2=1.795
r135 34 35 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.295 $Y=1.88
+ $X2=2.86 $Y2=1.88
r136 30 46 5.45789 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.765 $Y=2.085
+ $X2=2.765 $Y2=2
r137 30 32 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=2.765 $Y=2.085
+ $X2=2.765 $Y2=2.3
r138 29 38 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.415 $Y=2 $X2=1.265
+ $Y2=2
r139 28 46 1.09592 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.67 $Y=2 $X2=2.765
+ $Y2=2
r140 28 29 81.877 $w=1.68e-07 $l=1.255e-06 $layer=LI1_cond $X=2.67 $Y=2
+ $X2=1.415 $Y2=2
r141 24 40 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.2 $Y=2.3 $X2=1.2
+ $Y2=2.085
r142 19 57 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.07 $Y=0.995
+ $X2=4.07 $Y2=1.202
r143 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.07 $Y=0.995
+ $X2=4.07 $Y2=0.56
r144 16 56 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.045 $Y=1.41
+ $X2=4.045 $Y2=1.202
r145 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.045 $Y=1.41
+ $X2=4.045 $Y2=1.985
r146 13 55 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.565 $Y=0.995
+ $X2=3.565 $Y2=1.202
r147 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.565 $Y=0.995
+ $X2=3.565 $Y2=0.56
r148 10 54 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.54 $Y=1.41
+ $X2=3.54 $Y2=1.202
r149 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.54 $Y=1.41
+ $X2=3.54 $Y2=1.985
r150 3 32 600 $w=1.7e-07 $l=3.08504e-07 $layer=licon1_PDIFF $count=1 $X=2.585
+ $Y=2.065 $X2=2.755 $Y2=2.3
r151 2 24 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=2.065 $X2=1.2 $Y2=2.3
r152 1 42 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.175
+ $Y=0.235 $X2=1.3 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_2%VPWR 1 2 3 4 15 19 21 23 26 27 28 30 44 49
+ 54 57 60
r72 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r73 56 57 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=2.53
+ $X2=2.425 $Y2=2.53
r74 52 56 4.13191 $w=5.48e-07 $l=1.9e-07 $layer=LI1_cond $X=2.07 $Y=2.53
+ $X2=2.26 $Y2=2.53
r75 52 54 14.1814 $w=5.48e-07 $l=3.65e-07 $layer=LI1_cond $X=2.07 $Y=2.53
+ $X2=1.705 $Y2=2.53
r76 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r77 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r78 47 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r79 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r80 44 59 4.00497 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=4.195 $Y=2.72
+ $X2=4.397 $Y2=2.72
r81 44 46 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.195 $Y=2.72
+ $X2=3.91 $Y2=2.72
r82 43 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r83 43 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r84 42 57 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=2.425 $Y2=2.72
r85 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r86 39 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r87 39 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r88 38 54 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=1.705 $Y2=2.72
r89 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r90 36 49 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r91 36 38 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r92 30 49 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r93 30 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r94 28 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r95 28 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r96 26 42 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.14 $Y=2.72 $X2=2.99
+ $Y2=2.72
r97 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=2.72
+ $X2=3.305 $Y2=2.72
r98 25 46 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.47 $Y=2.72
+ $X2=3.91 $Y2=2.72
r99 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.47 $Y=2.72
+ $X2=3.305 $Y2=2.72
r100 21 59 3.17226 $w=2.55e-07 $l=1.16619e-07 $layer=LI1_cond $X=4.322 $Y=2.635
+ $X2=4.397 $Y2=2.72
r101 21 23 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=4.322 $Y=2.635
+ $X2=4.322 $Y2=2
r102 17 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=2.635
+ $X2=3.305 $Y2=2.72
r103 17 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.305 $Y=2.635
+ $X2=3.305 $Y2=2.34
r104 13 49 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r105 13 15 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.34
r106 4 23 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.135
+ $Y=1.485 $X2=4.28 $Y2=2
r107 3 19 600 $w=1.7e-07 $l=3.7081e-07 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=2.065 $X2=3.305 $Y2=2.34
r108 2 56 600 $w=1.7e-07 $l=3.7081e-07 $layer=licon1_PDIFF $count=1 $X=2.035
+ $Y=2.065 $X2=2.26 $Y2=2.34
r109 1 15 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.065 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_2%X 1 2 7 8 9 10 11 12 23 38 46
c43 38 0 6.07816e-20 $X=3.905 $Y=0.85
c44 10 0 1.96288e-19 $X=4.22 $Y=0.765
r45 46 52 0.0879469 $w=6.78e-07 $l=5e-09 $layer=LI1_cond $X=4.115 $Y=1.53
+ $X2=4.115 $Y2=1.535
r46 38 50 0.439735 $w=6.78e-07 $l=2.5e-08 $layer=LI1_cond $X=4.115 $Y=0.85
+ $X2=4.115 $Y2=0.825
r47 12 53 5.8779 $w=7.63e-07 $l=9e-08 $layer=LI1_cond $X=4.072 $Y=1.575
+ $X2=4.072 $Y2=1.665
r48 12 52 0.801609 $w=7.63e-07 $l=4e-08 $layer=LI1_cond $X=4.072 $Y=1.575
+ $X2=4.072 $Y2=1.535
r49 12 46 0.703576 $w=6.78e-07 $l=4e-08 $layer=LI1_cond $X=4.115 $Y=1.49
+ $X2=4.115 $Y2=1.53
r50 11 12 5.27682 $w=6.78e-07 $l=3e-07 $layer=LI1_cond $X=4.115 $Y=1.19
+ $X2=4.115 $Y2=1.49
r51 10 50 1.1424 $w=8.93e-07 $l=3e-08 $layer=LI1_cond $X=4.007 $Y=0.795
+ $X2=4.007 $Y2=0.825
r52 10 49 7.11295 $w=8.93e-07 $l=1.55e-07 $layer=LI1_cond $X=4.007 $Y=0.795
+ $X2=4.007 $Y2=0.64
r53 10 11 5.45271 $w=6.78e-07 $l=3.1e-07 $layer=LI1_cond $X=4.115 $Y=0.88
+ $X2=4.115 $Y2=1.19
r54 10 38 0.527682 $w=6.78e-07 $l=3e-08 $layer=LI1_cond $X=4.115 $Y=0.88
+ $X2=4.115 $Y2=0.85
r55 9 31 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=3.842 $Y=2.21
+ $X2=3.842 $Y2=1.96
r56 8 31 3.40065 $w=3.03e-07 $l=9e-08 $layer=LI1_cond $X=3.842 $Y=1.87 $X2=3.842
+ $Y2=1.96
r57 8 53 7.74593 $w=3.03e-07 $l=2.05e-07 $layer=LI1_cond $X=3.842 $Y=1.87
+ $X2=3.842 $Y2=1.665
r58 7 49 4.47217 $w=3.33e-07 $l=1.3e-07 $layer=LI1_cond $X=3.727 $Y=0.51
+ $X2=3.727 $Y2=0.64
r59 7 23 3.09612 $w=3.33e-07 $l=9e-08 $layer=LI1_cond $X=3.727 $Y=0.51 $X2=3.727
+ $Y2=0.42
r60 2 31 300 $w=1.7e-07 $l=5.57786e-07 $layer=licon1_PDIFF $count=2 $X=3.63
+ $Y=1.485 $X2=3.81 $Y2=1.96
r61 1 23 182 $w=1.7e-07 $l=2.56271e-07 $layer=licon1_NDIFF $count=1 $X=3.64
+ $Y=0.235 $X2=3.81 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_2%VGND 1 2 3 10 12 14 15 21 30 38 39
r61 38 41 10.7564 $w=4.31e-07 $l=3.8e-07 $layer=LI1_cond $X=4.332 $Y=0 $X2=4.332
+ $Y2=0.38
r62 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r63 33 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r64 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r65 30 38 6.2345 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=4.065 $Y=0 $X2=4.332
+ $Y2=0
r66 30 32 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.065 $Y=0 $X2=3.91
+ $Y2=0
r67 29 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r68 28 29 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r69 26 29 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.99
+ $Y2=0
r70 25 28 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.99
+ $Y2=0
r71 25 26 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r72 23 35 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r73 23 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r74 21 26 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r75 21 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r76 17 32 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.39 $Y=0 $X2=3.91
+ $Y2=0
r77 15 28 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.01 $Y=0 $X2=2.99
+ $Y2=0
r78 14 19 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.2 $Y=0 $X2=3.2
+ $Y2=0.38
r79 14 17 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.2 $Y=0 $X2=3.39
+ $Y2=0
r80 14 15 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.2 $Y=0 $X2=3.01
+ $Y2=0
r81 10 35 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r82 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r83 3 41 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.145
+ $Y=0.235 $X2=4.28 $Y2=0.38
r84 2 19 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.09
+ $Y=0.235 $X2=3.225 $Y2=0.38
r85 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

