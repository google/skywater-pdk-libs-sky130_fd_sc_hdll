* File: sky130_fd_sc_hdll__inputiso0n_1.pex.spice
* Created: Wed Sep  2 08:32:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%A 2 3 5 8 10 11 15 16
r32 19 25 0.382416 $w=2.65e-07 $l=1.25e-07 $layer=LI1_cond $X=0.232 $Y=1.325
+ $X2=0.232 $Y2=1.2
r33 16 25 8.89686 $w=2.48e-07 $l=1.93e-07 $layer=LI1_cond $X=0.425 $Y=1.2
+ $X2=0.232 $Y2=1.2
r34 15 18 37.7763 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.452 $Y=1.16
+ $X2=0.452 $Y2=1.325
r35 15 17 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.452 $Y=1.16
+ $X2=0.452 $Y2=0.995
r36 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.425
+ $Y=1.16 $X2=0.425 $Y2=1.16
r37 11 19 8.91512 $w=2.63e-07 $l=2.05e-07 $layer=LI1_cond $X=0.232 $Y=1.53
+ $X2=0.232 $Y2=1.325
r38 10 25 0.0921954 $w=2.48e-07 $l=2e-09 $layer=LI1_cond $X=0.23 $Y=1.2
+ $X2=0.232 $Y2=1.2
r39 8 17 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.54 $Y=0.585
+ $X2=0.54 $Y2=0.995
r40 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.515 $Y=1.78
+ $X2=0.515 $Y2=2.065
r41 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.515 $Y=1.68 $X2=0.515
+ $Y2=1.78
r42 2 18 117.71 $w=2e-07 $l=3.55e-07 $layer=POLY_cond $X=0.515 $Y=1.68 $X2=0.515
+ $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%SLEEP_B 3 6 7 9 10 13 20
r40 13 16 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.02 $Y=1.16
+ $X2=1.02 $Y2=1.325
r41 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.02 $Y=1.16
+ $X2=1.02 $Y2=0.995
r42 10 20 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=1.02 $Y=1.2 $X2=1.1
+ $Y2=1.2
r43 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.02
+ $Y=1.16 $X2=1.02 $Y2=1.16
r44 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.985 $Y=1.78
+ $X2=0.985 $Y2=2.065
r45 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.985 $Y=1.68 $X2=0.985
+ $Y2=1.78
r46 6 16 117.71 $w=2e-07 $l=3.55e-07 $layer=POLY_cond $X=0.985 $Y=1.68 $X2=0.985
+ $Y2=1.325
r47 3 15 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.96 $Y=0.585
+ $X2=0.96 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%A_27_75# 1 2 7 9 10 12 15 17 18 21 23
+ 24 28
r69 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.16 $X2=1.61 $Y2=1.16
r70 26 28 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.61 $Y=1.575
+ $X2=1.61 $Y2=1.16
r71 25 28 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.61 $Y=0.905
+ $X2=1.61 $Y2=1.16
r72 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.525 $Y=1.66
+ $X2=1.61 $Y2=1.575
r73 23 24 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.525 $Y=1.66
+ $X2=0.925 $Y2=1.66
r74 19 24 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=0.775 $Y=1.745
+ $X2=0.925 $Y2=1.66
r75 19 21 14.7897 $w=2.98e-07 $l=3.85e-07 $layer=LI1_cond $X=0.775 $Y=1.745
+ $X2=0.775 $Y2=2.13
r76 17 25 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.525 $Y=0.81
+ $X2=1.61 $Y2=0.905
r77 17 18 62.4593 $w=1.88e-07 $l=1.07e-06 $layer=LI1_cond $X=1.525 $Y=0.81
+ $X2=0.455 $Y2=0.81
r78 13 18 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=0.29 $Y=0.715
+ $X2=0.455 $Y2=0.81
r79 13 15 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.29 $Y=0.715
+ $X2=0.29 $Y2=0.52
r80 10 29 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.575 $Y=1.41
+ $X2=1.61 $Y2=1.16
r81 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.575 $Y=1.41
+ $X2=1.575 $Y2=1.985
r82 7 29 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.55 $Y=0.995
+ $X2=1.61 $Y2=1.16
r83 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.55 $Y=0.995 $X2=1.55
+ $Y2=0.56
r84 2 21 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.855 $X2=0.75 $Y2=2.13
r85 1 15 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.375 $X2=0.28 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%VPWR 1 2 7 9 13 16 17 18 25 26
r30 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r31 23 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r32 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r33 20 29 4.25667 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=2.72
+ $X2=0.202 $Y2=2.72
r34 20 22 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=0.405 $Y=2.72
+ $X2=1.15 $Y2=2.72
r35 18 23 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r36 18 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r37 16 22 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.175 $Y=2.72
+ $X2=1.15 $Y2=2.72
r38 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.175 $Y=2.72
+ $X2=1.34 $Y2=2.72
r39 15 25 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.505 $Y=2.72
+ $X2=2.07 $Y2=2.72
r40 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=2.72
+ $X2=1.34 $Y2=2.72
r41 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.34 $Y=2.635
+ $X2=1.34 $Y2=2.72
r42 11 13 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.34 $Y=2.635
+ $X2=1.34 $Y2=2
r43 7 29 3.10338 $w=2.8e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.202 $Y2=2.72
r44 7 9 20.7851 $w=2.78e-07 $l=5.05e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.265 $Y2=2.13
r45 2 13 300 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_PDIFF $count=2 $X=1.075
+ $Y=1.855 $X2=1.34 $Y2=2
r46 1 9 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.855 $X2=0.28 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%X 1 2 7 11 12 13 14 15 16 25 36
r23 36 40 2.0744 $w=2.48e-07 $l=4.5e-08 $layer=LI1_cond $X=2.08 $Y=1.87 $X2=2.08
+ $Y2=1.915
r24 16 42 5.46036 $w=4.58e-07 $l=2.1e-07 $layer=LI1_cond $X=1.975 $Y=2.21
+ $X2=1.975 $Y2=2
r25 15 42 1.69011 $w=4.58e-07 $l=6.5e-08 $layer=LI1_cond $X=1.975 $Y=1.935
+ $X2=1.975 $Y2=2
r26 15 40 2.99563 $w=4.58e-07 $l=2e-08 $layer=LI1_cond $X=1.975 $Y=1.935
+ $X2=1.975 $Y2=1.915
r27 15 36 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=2.08 $Y=1.85 $X2=2.08
+ $Y2=1.87
r28 14 15 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=2.08 $Y=1.53
+ $X2=2.08 $Y2=1.85
r29 13 14 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=2.08 $Y=1.19
+ $X2=2.08 $Y2=1.53
r30 12 13 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=2.08 $Y=0.85
+ $X2=2.08 $Y2=1.19
r31 11 25 3.6869 $w=2.5e-07 $l=1.45e-07 $layer=LI1_cond $X=2.08 $Y=0.4 $X2=2.08
+ $Y2=0.545
r32 11 12 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=2.08 $Y=0.57
+ $X2=2.08 $Y2=0.85
r33 11 25 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=2.08 $Y=0.57
+ $X2=2.08 $Y2=0.545
r34 7 11 3.17836 $w=2.9e-07 $l=1.25e-07 $layer=LI1_cond $X=1.955 $Y=0.4 $X2=2.08
+ $Y2=0.4
r35 7 9 7.74919 $w=2.88e-07 $l=1.95e-07 $layer=LI1_cond $X=1.955 $Y=0.4 $X2=1.76
+ $Y2=0.4
r36 2 42 300 $w=1.7e-07 $l=6.2562e-07 $layer=licon1_PDIFF $count=2 $X=1.665
+ $Y=1.485 $X2=1.91 $Y2=2
r37 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.625
+ $Y=0.235 $X2=1.76 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%VGND 1 6 9 10 11 21 22
r25 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r26 19 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r27 18 19 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r28 14 18 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r29 11 19 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r30 11 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r31 9 18 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.175 $Y=0 $X2=1.15
+ $Y2=0
r32 9 10 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.175 $Y=0 $X2=1.3
+ $Y2=0
r33 8 21 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=2.07
+ $Y2=0
r34 8 10 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=1.3
+ $Y2=0
r35 4 10 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=0.085
+ $X2=1.3 $Y2=0
r36 4 6 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.3 $Y=0.085 $X2=1.3
+ $Y2=0.38
r37 1 6 182 $w=1.7e-07 $l=3.0749e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.375 $X2=1.34 $Y2=0.38
.ends

