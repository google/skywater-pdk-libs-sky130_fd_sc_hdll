* File: sky130_fd_sc_hdll__inputiso1p_1.pex.spice
* Created: Wed Sep  2 08:32:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%A 1 3 6 8 9
r23 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.355
+ $Y=1.16 $X2=0.355 $Y2=1.16
r24 9 14 0.973895 $w=3.53e-07 $l=3e-08 $layer=LI1_cond $X=0.262 $Y=1.19
+ $X2=0.262 $Y2=1.16
r25 8 14 10.0636 $w=3.53e-07 $l=3.1e-07 $layer=LI1_cond $X=0.262 $Y=0.85
+ $X2=0.262 $Y2=1.16
r26 4 13 40.2182 $w=4.3e-07 $l=2.38642e-07 $layer=POLY_cond $X=0.605 $Y=0.995
+ $X2=0.435 $Y2=1.16
r27 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.605 $Y=0.995
+ $X2=0.605 $Y2=0.445
r28 1 13 44.7166 $w=4.3e-07 $l=3.14245e-07 $layer=POLY_cond $X=0.58 $Y=1.41
+ $X2=0.435 $Y2=1.16
r29 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.58 $Y=1.41 $X2=0.58
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%SLEEP 3 5 7 8 9
r30 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.085
+ $Y=1.16 $X2=1.085 $Y2=1.16
r31 8 9 11.3415 $w=3.13e-07 $l=3.1e-07 $layer=LI1_cond $X=1.157 $Y=0.85
+ $X2=1.157 $Y2=1.16
r32 5 13 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=1.05 $Y=1.41
+ $X2=1.11 $Y2=1.16
r33 5 7 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.05 $Y=1.41 $X2=1.05
+ $Y2=1.695
r34 1 13 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.025 $Y=0.995
+ $X2=1.11 $Y2=1.16
r35 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.025 $Y=0.995
+ $X2=1.025 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%A_44_297# 1 2 7 9 10 12 14 15 16 19
+ 26
c45 14 0 1.05122e-19 $X=0.72 $Y=1.495
r46 26 28 7.04571 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.775 $Y=0.43
+ $X2=0.775 $Y2=0.595
r47 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.62
+ $Y=1.16 $X2=1.62 $Y2=1.16
r48 17 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.62 $Y=1.495
+ $X2=1.62 $Y2=1.16
r49 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.535 $Y=1.58
+ $X2=1.62 $Y2=1.495
r50 15 16 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=1.535 $Y=1.58
+ $X2=0.83 $Y2=1.58
r51 14 16 6.63579 $w=2.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.72 $Y=1.495
+ $X2=0.83 $Y2=1.58
r52 14 23 16.9444 $w=2.7e-07 $l=4.52907e-07 $layer=LI1_cond $X=0.72 $Y=1.495
+ $X2=0.345 $Y2=1.667
r53 14 28 47.1454 $w=2.18e-07 $l=9e-07 $layer=LI1_cond $X=0.72 $Y=1.495 $X2=0.72
+ $Y2=0.595
r54 10 20 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.585 $Y=1.41
+ $X2=1.62 $Y2=1.16
r55 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.585 $Y=1.41
+ $X2=1.585 $Y2=1.985
r56 7 20 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.56 $Y=0.995
+ $X2=1.62 $Y2=1.16
r57 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.56 $Y=0.995 $X2=1.56
+ $Y2=0.56
r58 2 23 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.22
+ $Y=1.485 $X2=0.345 $Y2=1.66
r59 1 26 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=0.68
+ $Y=0.235 $X2=0.815 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%VPWR 1 6 9 10 11 21 22
r20 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r21 19 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r22 18 19 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r23 14 18 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r24 11 19 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r25 11 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r26 9 18 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.15 $Y2=2.72
r27 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.35 $Y2=2.72
r28 8 21 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.515 $Y=2.72
+ $X2=2.07 $Y2=2.72
r29 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=2.72
+ $X2=1.35 $Y2=2.72
r30 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=2.635 $X2=1.35
+ $Y2=2.72
r31 4 6 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=1.35 $Y=2.635
+ $X2=1.35 $Y2=1.92
r32 1 6 300 $w=1.7e-07 $l=5.29693e-07 $layer=licon1_PDIFF $count=2 $X=1.14
+ $Y=1.485 $X2=1.35 $Y2=1.92
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%X 1 2 9 12 18
r18 18 19 1.43211 $w=4.18e-07 $l=2.5e-08 $layer=LI1_cond $X=2.005 $Y=1.87
+ $X2=2.005 $Y2=1.845
r19 12 22 2.74391 $w=4.18e-07 $l=1e-07 $layer=LI1_cond $X=2.005 $Y=1.9 $X2=2.005
+ $Y2=2
r20 12 18 0.823174 $w=4.18e-07 $l=3e-08 $layer=LI1_cond $X=2.005 $Y=1.9
+ $X2=2.005 $Y2=1.87
r21 12 19 1.09756 $w=3.13e-07 $l=3e-08 $layer=LI1_cond $X=2.057 $Y=1.815
+ $X2=2.057 $Y2=1.845
r22 11 12 36.2196 $w=3.13e-07 $l=9.9e-07 $layer=LI1_cond $X=2.057 $Y=0.825
+ $X2=2.057 $Y2=1.815
r23 9 11 11.6252 $w=5.48e-07 $l=4.35e-07 $layer=LI1_cond $X=1.94 $Y=0.39
+ $X2=1.94 $Y2=0.825
r24 2 22 300 $w=1.7e-07 $l=6.41872e-07 $layer=licon1_PDIFF $count=2 $X=1.675
+ $Y=1.485 $X2=1.96 $Y2=2
r25 1 9 91 $w=1.7e-07 $l=3.1305e-07 $layer=licon1_NDIFF $count=2 $X=1.635
+ $Y=0.235 $X2=1.88 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%VGND 1 2 7 9 13 16 17 18 25 26
r31 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r32 23 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r33 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r34 20 29 3.85266 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.215
+ $Y2=0
r35 20 22 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=1.15
+ $Y2=0
r36 18 23 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r37 18 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r38 16 22 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=1.22 $Y=0 $X2=1.15
+ $Y2=0
r39 16 17 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=1.327
+ $Y2=0
r40 15 25 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.435 $Y=0 $X2=2.07
+ $Y2=0
r41 15 17 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.327
+ $Y2=0
r42 11 17 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.327 $Y=0.085
+ $X2=1.327 $Y2=0
r43 11 13 18.4927 $w=2.13e-07 $l=3.45e-07 $layer=LI1_cond $X=1.327 $Y=0.085
+ $X2=1.327 $Y2=0.43
r44 7 29 3.22548 $w=2.4e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.31 $Y=0.085
+ $X2=0.215 $Y2=0
r45 7 9 16.5664 $w=2.38e-07 $l=3.45e-07 $layer=LI1_cond $X=0.31 $Y=0.085
+ $X2=0.31 $Y2=0.43
r46 2 13 182 $w=1.7e-07 $l=3.28329e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.235 $X2=1.345 $Y2=0.43
r47 1 9 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.22
+ $Y=0.235 $X2=0.345 $Y2=0.43
.ends

