* File: sky130_fd_sc_hdll__nor4bb_4.pex.spice
* Created: Wed Sep  2 08:42:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_4%C_N 1 3 4 6 7 12 15
c26 4 0 1.23817e-19 $X=0.54 $Y=0.995
c27 1 0 1.26528e-19 $X=0.515 $Y=1.41
r28 12 13 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.54 $Y2=1.202
r29 10 12 30.9481 $w=3.66e-07 $l=2.35e-07 $layer=POLY_cond $X=0.28 $Y=1.202
+ $X2=0.515 $Y2=1.202
r30 7 15 0.198697 $w=2.88e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=1.22 $X2=0.23
+ $Y2=1.22
r31 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.28
+ $Y=1.16 $X2=0.28 $Y2=1.16
r32 4 13 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.54 $Y2=1.202
r33 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.54 $Y=0.995 $X2=0.54
+ $Y2=0.56
r34 1 12 19.3576 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r35 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_4%D_N 1 3 4 6 7 10 15
r40 10 12 31.1181 $w=3.64e-07 $l=2.35e-07 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.22 $Y2=1.202
r41 9 10 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=0.96 $Y=1.202
+ $X2=0.985 $Y2=1.202
r42 7 15 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=1.16 $Y=1.2 $X2=1.15
+ $Y2=1.2
r43 7 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.22
+ $Y=1.16 $X2=1.22 $Y2=1.16
r44 4 10 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r45 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r46 1 9 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.96 $Y=0.995 $X2=0.96
+ $Y2=1.202
r47 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.96 $Y=0.995 $X2=0.96
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_4%A_207_47# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 33 35 39 40 42 44 50 53 62
c124 40 0 1.23817e-19 $X=1.385 $Y=0.82
c125 35 0 1.26528e-19 $X=1.565 $Y=1.62
c126 25 0 2.79668e-20 $X=3.425 $Y=1.41
c127 22 0 7.87746e-20 $X=2.955 $Y=1.41
r128 62 63 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.425 $Y=1.202
+ $X2=3.45 $Y2=1.202
r129 61 62 60.8979 $w=3.72e-07 $l=4.7e-07 $layer=POLY_cond $X=2.955 $Y=1.202
+ $X2=3.425 $Y2=1.202
r130 60 61 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.93 $Y=1.202
+ $X2=2.955 $Y2=1.202
r131 57 58 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.46 $Y=1.202
+ $X2=2.485 $Y2=1.202
r132 54 55 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.99 $Y=1.202
+ $X2=2.015 $Y2=1.202
r133 51 60 6.47849 $w=3.72e-07 $l=5e-08 $layer=POLY_cond $X=2.88 $Y=1.202
+ $X2=2.93 $Y2=1.202
r134 51 58 51.1801 $w=3.72e-07 $l=3.95e-07 $layer=POLY_cond $X=2.88 $Y=1.202
+ $X2=2.485 $Y2=1.202
r135 50 51 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.88
+ $Y=1.16 $X2=2.88 $Y2=1.16
r136 48 57 46.6452 $w=3.72e-07 $l=3.6e-07 $layer=POLY_cond $X=2.1 $Y=1.202
+ $X2=2.46 $Y2=1.202
r137 48 55 11.0134 $w=3.72e-07 $l=8.5e-08 $layer=POLY_cond $X=2.1 $Y=1.202
+ $X2=2.015 $Y2=1.202
r138 47 50 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=2.1 $Y=1.16
+ $X2=2.88 $Y2=1.16
r139 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.1
+ $Y=1.16 $X2=2.1 $Y2=1.16
r140 45 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.735 $Y=1.16
+ $X2=1.65 $Y2=1.16
r141 45 47 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.735 $Y=1.16
+ $X2=2.1 $Y2=1.16
r142 43 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=1.245
+ $X2=1.65 $Y2=1.16
r143 43 44 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.65 $Y=1.245
+ $X2=1.65 $Y2=1.535
r144 42 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=1.075
+ $X2=1.65 $Y2=1.16
r145 41 42 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.65 $Y=0.905
+ $X2=1.65 $Y2=1.075
r146 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.565 $Y=0.82
+ $X2=1.65 $Y2=0.905
r147 39 40 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.565 $Y=0.82
+ $X2=1.385 $Y2=0.82
r148 35 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.565 $Y=1.62
+ $X2=1.65 $Y2=1.535
r149 35 37 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.565 $Y=1.62
+ $X2=1.22 $Y2=1.62
r150 31 40 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=1.195 $Y=0.735
+ $X2=1.385 $Y2=0.82
r151 31 33 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=1.195 $Y=0.735
+ $X2=1.195 $Y2=0.39
r152 28 63 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.45 $Y=0.995
+ $X2=3.45 $Y2=1.202
r153 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.45 $Y=0.995
+ $X2=3.45 $Y2=0.56
r154 25 62 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.425 $Y=1.41
+ $X2=3.425 $Y2=1.202
r155 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.425 $Y=1.41
+ $X2=3.425 $Y2=1.985
r156 22 61 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.955 $Y=1.41
+ $X2=2.955 $Y2=1.202
r157 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.955 $Y=1.41
+ $X2=2.955 $Y2=1.985
r158 19 60 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.93 $Y=0.995
+ $X2=2.93 $Y2=1.202
r159 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.93 $Y=0.995
+ $X2=2.93 $Y2=0.56
r160 16 58 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.485 $Y=1.41
+ $X2=2.485 $Y2=1.202
r161 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.485 $Y=1.41
+ $X2=2.485 $Y2=1.985
r162 13 57 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.46 $Y=0.995
+ $X2=2.46 $Y2=1.202
r163 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.46 $Y=0.995
+ $X2=2.46 $Y2=0.56
r164 10 55 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.015 $Y=1.41
+ $X2=2.015 $Y2=1.202
r165 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.015 $Y=1.41
+ $X2=2.015 $Y2=1.985
r166 7 54 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.99 $Y=0.995
+ $X2=1.99 $Y2=1.202
r167 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.99 $Y=0.995
+ $X2=1.99 $Y2=0.56
r168 2 37 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.62
r169 1 33 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.035
+ $Y=0.235 $X2=1.22 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_4%A_27_297# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 33 37 39 40 42 43 46 47 52 60 69
c149 46 0 1.21732e-19 $X=3.74 $Y=1.875
c150 10 0 3.26191e-21 $X=3.895 $Y=1.41
r151 69 70 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.305 $Y=1.202
+ $X2=5.33 $Y2=1.202
r152 66 67 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.81 $Y=1.202
+ $X2=4.835 $Y2=1.202
r153 65 66 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=4.365 $Y=1.202
+ $X2=4.81 $Y2=1.202
r154 64 65 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.34 $Y=1.202
+ $X2=4.365 $Y2=1.202
r155 61 62 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.87 $Y=1.202
+ $X2=3.895 $Y2=1.202
r156 59 60 7.70264 $w=5.08e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=1.79
+ $X2=0.835 $Y2=1.79
r157 58 59 11.0227 $w=5.08e-07 $l=4.7e-07 $layer=LI1_cond $X=0.28 $Y=1.79
+ $X2=0.75 $Y2=1.79
r158 55 58 1.28989 $w=5.08e-07 $l=5.5e-08 $layer=LI1_cond $X=0.225 $Y=1.79
+ $X2=0.28 $Y2=1.79
r159 53 69 14.9005 $w=3.72e-07 $l=1.15e-07 $layer=POLY_cond $X=5.19 $Y=1.202
+ $X2=5.305 $Y2=1.202
r160 53 67 45.9973 $w=3.72e-07 $l=3.55e-07 $layer=POLY_cond $X=5.19 $Y=1.202
+ $X2=4.835 $Y2=1.202
r161 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.19
+ $Y=1.16 $X2=5.19 $Y2=1.16
r162 50 64 41.4624 $w=3.72e-07 $l=3.2e-07 $layer=POLY_cond $X=4.02 $Y=1.202
+ $X2=4.34 $Y2=1.202
r163 50 62 16.1962 $w=3.72e-07 $l=1.25e-07 $layer=POLY_cond $X=4.02 $Y=1.202
+ $X2=3.895 $Y2=1.202
r164 49 52 61.7922 $w=2.08e-07 $l=1.17e-06 $layer=LI1_cond $X=4.02 $Y=1.18
+ $X2=5.19 $Y2=1.18
r165 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.02
+ $Y=1.16 $X2=4.02 $Y2=1.16
r166 47 49 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=3.825 $Y=1.18
+ $X2=4.02 $Y2=1.18
r167 45 47 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.74 $Y=1.285
+ $X2=3.825 $Y2=1.18
r168 45 46 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.74 $Y=1.285
+ $X2=3.74 $Y2=1.875
r169 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.655 $Y=1.96
+ $X2=3.74 $Y2=1.875
r170 43 60 183.979 $w=1.68e-07 $l=2.82e-06 $layer=LI1_cond $X=3.655 $Y=1.96
+ $X2=0.835 $Y2=1.96
r171 42 59 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.75 $Y=1.535
+ $X2=0.75 $Y2=1.79
r172 41 42 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.75 $Y=0.895
+ $X2=0.75 $Y2=1.535
r173 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=0.81
+ $X2=0.75 $Y2=0.895
r174 39 40 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.665 $Y=0.81
+ $X2=0.445 $Y2=0.81
r175 35 55 4.24724 $w=2.8e-07 $l=2.55e-07 $layer=LI1_cond $X=0.225 $Y=2.045
+ $X2=0.225 $Y2=1.79
r176 35 37 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=0.225 $Y=2.045
+ $X2=0.225 $Y2=2.3
r177 31 40 8.02311 $w=1.7e-07 $l=2.18403e-07 $layer=LI1_cond $X=0.265 $Y=0.725
+ $X2=0.445 $Y2=0.81
r178 31 33 10.7241 $w=3.58e-07 $l=3.35e-07 $layer=LI1_cond $X=0.265 $Y=0.725
+ $X2=0.265 $Y2=0.39
r179 28 70 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.33 $Y=0.995
+ $X2=5.33 $Y2=1.202
r180 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.33 $Y=0.995
+ $X2=5.33 $Y2=0.56
r181 25 69 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.305 $Y=1.41
+ $X2=5.305 $Y2=1.202
r182 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.305 $Y=1.41
+ $X2=5.305 $Y2=1.985
r183 22 67 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.835 $Y=1.41
+ $X2=4.835 $Y2=1.202
r184 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.835 $Y=1.41
+ $X2=4.835 $Y2=1.985
r185 19 66 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.81 $Y=0.995
+ $X2=4.81 $Y2=1.202
r186 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.81 $Y=0.995
+ $X2=4.81 $Y2=0.56
r187 16 65 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.365 $Y=1.41
+ $X2=4.365 $Y2=1.202
r188 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.365 $Y=1.41
+ $X2=4.365 $Y2=1.985
r189 13 64 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.34 $Y=0.995
+ $X2=4.34 $Y2=1.202
r190 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.34 $Y=0.995
+ $X2=4.34 $Y2=0.56
r191 10 62 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.895 $Y=1.41
+ $X2=3.895 $Y2=1.202
r192 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.895 $Y=1.41
+ $X2=3.895 $Y2=1.985
r193 7 61 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.87 $Y=0.995
+ $X2=3.87 $Y2=1.202
r194 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.87 $Y=0.995
+ $X2=3.87 $Y2=0.56
r195 2 58 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r196 2 37 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r197 1 33 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_4%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39 44
r77 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.705 $Y=1.202
+ $X2=7.73 $Y2=1.202
r78 37 39 14.9005 $w=3.72e-07 $l=1.15e-07 $layer=POLY_cond $X=7.59 $Y=1.202
+ $X2=7.705 $Y2=1.202
r79 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.59
+ $Y=1.16 $X2=7.59 $Y2=1.16
r80 35 37 45.9973 $w=3.72e-07 $l=3.55e-07 $layer=POLY_cond $X=7.235 $Y=1.202
+ $X2=7.59 $Y2=1.202
r81 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.21 $Y=1.202
+ $X2=7.235 $Y2=1.202
r82 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=6.765 $Y=1.202
+ $X2=7.21 $Y2=1.202
r83 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.74 $Y=1.202
+ $X2=6.765 $Y2=1.202
r84 31 44 5.54545 $w=2.08e-07 $l=1.05e-07 $layer=LI1_cond $X=6.42 $Y=1.18
+ $X2=6.525 $Y2=1.18
r85 30 32 41.4624 $w=3.72e-07 $l=3.2e-07 $layer=POLY_cond $X=6.42 $Y=1.202
+ $X2=6.74 $Y2=1.202
r86 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.42
+ $Y=1.16 $X2=6.42 $Y2=1.16
r87 28 30 16.1962 $w=3.72e-07 $l=1.25e-07 $layer=POLY_cond $X=6.295 $Y=1.202
+ $X2=6.42 $Y2=1.202
r88 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.27 $Y=1.202
+ $X2=6.295 $Y2=1.202
r89 25 38 48.0606 $w=2.08e-07 $l=9.1e-07 $layer=LI1_cond $X=6.68 $Y=1.18
+ $X2=7.59 $Y2=1.18
r90 25 44 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=6.68 $Y=1.18
+ $X2=6.525 $Y2=1.18
r91 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.73 $Y=0.995
+ $X2=7.73 $Y2=1.202
r92 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.73 $Y=0.995
+ $X2=7.73 $Y2=0.56
r93 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.705 $Y=1.41
+ $X2=7.705 $Y2=1.202
r94 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.705 $Y=1.41
+ $X2=7.705 $Y2=1.985
r95 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.235 $Y=1.41
+ $X2=7.235 $Y2=1.202
r96 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.235 $Y=1.41
+ $X2=7.235 $Y2=1.985
r97 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.21 $Y=0.995
+ $X2=7.21 $Y2=1.202
r98 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.21 $Y=0.995
+ $X2=7.21 $Y2=0.56
r99 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.765 $Y=1.41
+ $X2=6.765 $Y2=1.202
r100 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.765 $Y=1.41
+ $X2=6.765 $Y2=1.985
r101 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.74 $Y=0.995
+ $X2=6.74 $Y2=1.202
r102 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.74 $Y=0.995
+ $X2=6.74 $Y2=0.56
r103 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.295 $Y=1.41
+ $X2=6.295 $Y2=1.202
r104 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.295 $Y=1.41
+ $X2=6.295 $Y2=1.985
r105 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.27 $Y=0.995
+ $X2=6.27 $Y2=1.202
r106 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.27 $Y=0.995
+ $X2=6.27 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39 44
r69 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=9.585 $Y=1.202
+ $X2=9.61 $Y2=1.202
r70 37 39 14.9005 $w=3.72e-07 $l=1.15e-07 $layer=POLY_cond $X=9.47 $Y=1.202
+ $X2=9.585 $Y2=1.202
r71 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.47
+ $Y=1.16 $X2=9.47 $Y2=1.16
r72 35 37 45.9973 $w=3.72e-07 $l=3.55e-07 $layer=POLY_cond $X=9.115 $Y=1.202
+ $X2=9.47 $Y2=1.202
r73 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=9.09 $Y=1.202
+ $X2=9.115 $Y2=1.202
r74 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=8.645 $Y=1.202
+ $X2=9.09 $Y2=1.202
r75 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.62 $Y=1.202
+ $X2=8.645 $Y2=1.202
r76 31 44 29.0476 $w=2.08e-07 $l=5.5e-07 $layer=LI1_cond $X=8.3 $Y=1.18 $X2=8.85
+ $Y2=1.18
r77 30 32 41.4624 $w=3.72e-07 $l=3.2e-07 $layer=POLY_cond $X=8.3 $Y=1.202
+ $X2=8.62 $Y2=1.202
r78 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.3 $Y=1.16
+ $X2=8.3 $Y2=1.16
r79 28 30 16.1962 $w=3.72e-07 $l=1.25e-07 $layer=POLY_cond $X=8.175 $Y=1.202
+ $X2=8.3 $Y2=1.202
r80 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.15 $Y=1.202
+ $X2=8.175 $Y2=1.202
r81 25 38 26.4069 $w=2.08e-07 $l=5e-07 $layer=LI1_cond $X=8.97 $Y=1.18 $X2=9.47
+ $Y2=1.18
r82 25 44 6.33766 $w=2.08e-07 $l=1.2e-07 $layer=LI1_cond $X=8.97 $Y=1.18
+ $X2=8.85 $Y2=1.18
r83 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.61 $Y=0.995
+ $X2=9.61 $Y2=1.202
r84 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.61 $Y=0.995
+ $X2=9.61 $Y2=0.56
r85 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.585 $Y=1.41
+ $X2=9.585 $Y2=1.202
r86 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.585 $Y=1.41
+ $X2=9.585 $Y2=1.985
r87 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.115 $Y=1.41
+ $X2=9.115 $Y2=1.202
r88 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.115 $Y=1.41
+ $X2=9.115 $Y2=1.985
r89 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.09 $Y=0.995
+ $X2=9.09 $Y2=1.202
r90 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.09 $Y=0.995
+ $X2=9.09 $Y2=0.56
r91 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.645 $Y=1.41
+ $X2=8.645 $Y2=1.202
r92 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.645 $Y=1.41
+ $X2=8.645 $Y2=1.985
r93 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.62 $Y=0.995
+ $X2=8.62 $Y2=1.202
r94 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.62 $Y=0.995 $X2=8.62
+ $Y2=0.56
r95 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.175 $Y=1.41
+ $X2=8.175 $Y2=1.202
r96 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.175 $Y=1.41
+ $X2=8.175 $Y2=1.985
r97 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.15 $Y=0.995
+ $X2=8.15 $Y2=1.202
r98 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.15 $Y=0.995 $X2=8.15
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_4%VPWR 1 2 3 12 16 20 23 24 26 27 28 30 46
+ 47 50
r106 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r107 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r108 44 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r109 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r110 41 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r111 40 41 1.1625 $w=1.7e-07 $l=1.36e-06 $layer=mcon $count=8 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r112 38 41 1.96334 $w=4.8e-07 $l=6.9e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=8.05 $Y2=2.72
r113 38 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r114 37 40 450.16 $w=1.68e-07 $l=6.9e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=8.05 $Y2=2.72
r115 37 38 1.1625 $w=1.7e-07 $l=1.36e-06 $layer=mcon $count=8 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r116 35 50 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.915 $Y=2.72
+ $X2=0.725 $Y2=2.72
r117 35 37 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.915 $Y=2.72
+ $X2=1.15 $Y2=2.72
r118 30 50 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.725 $Y2=2.72
r119 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.23 $Y2=2.72
r120 28 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r121 28 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r122 26 43 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=9.225 $Y=2.72
+ $X2=8.97 $Y2=2.72
r123 26 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.225 $Y=2.72
+ $X2=9.35 $Y2=2.72
r124 25 46 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.475 $Y=2.72
+ $X2=9.89 $Y2=2.72
r125 25 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.475 $Y=2.72
+ $X2=9.35 $Y2=2.72
r126 23 40 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=8.285 $Y=2.72
+ $X2=8.05 $Y2=2.72
r127 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.285 $Y=2.72
+ $X2=8.41 $Y2=2.72
r128 22 43 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=8.535 $Y=2.72
+ $X2=8.97 $Y2=2.72
r129 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.535 $Y=2.72
+ $X2=8.41 $Y2=2.72
r130 18 27 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.35 $Y=2.635
+ $X2=9.35 $Y2=2.72
r131 18 20 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=9.35 $Y=2.635
+ $X2=9.35 $Y2=1.96
r132 14 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.41 $Y=2.635
+ $X2=8.41 $Y2=2.72
r133 14 16 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=8.41 $Y=2.635
+ $X2=8.41 $Y2=1.96
r134 10 50 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=2.635
+ $X2=0.725 $Y2=2.72
r135 10 12 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.725 $Y=2.635
+ $X2=0.725 $Y2=2.3
r136 3 20 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=9.205
+ $Y=1.485 $X2=9.35 $Y2=1.96
r137 2 16 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=8.265
+ $Y=1.485 $X2=8.41 $Y2=1.96
r138 1 12 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_4%A_331_297# 1 2 3 4 5 16 24 28 30 34 36 37
r48 32 34 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.555 $Y=2.295
+ $X2=5.555 $Y2=1.96
r49 31 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.725 $Y=2.38
+ $X2=4.6 $Y2=2.38
r50 30 32 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=5.415 $Y=2.38
+ $X2=5.555 $Y2=2.295
r51 30 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.415 $Y=2.38
+ $X2=4.725 $Y2=2.38
r52 26 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.6 $Y=2.295
+ $X2=4.6 $Y2=2.38
r53 26 28 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.6 $Y=2.295
+ $X2=4.6 $Y2=1.96
r54 24 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.475 $Y=2.38
+ $X2=4.6 $Y2=2.38
r55 24 36 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.475 $Y=2.38
+ $X2=3.825 $Y2=2.38
r56 21 23 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=2.72 $Y=2.34
+ $X2=3.66 $Y2=2.34
r57 18 21 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=1.78 $Y=2.34
+ $X2=2.72 $Y2=2.34
r58 16 36 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.7 $Y=2.34
+ $X2=3.825 $Y2=2.34
r59 16 23 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=3.7 $Y=2.34 $X2=3.66
+ $Y2=2.34
r60 5 34 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.395
+ $Y=1.485 $X2=5.54 $Y2=1.96
r61 4 28 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.455
+ $Y=1.485 $X2=4.6 $Y2=1.96
r62 3 23 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.485 $X2=3.66 $Y2=2.3
r63 2 21 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.575
+ $Y=1.485 $X2=2.72 $Y2=2.3
r64 1 18 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=1.655
+ $Y=1.485 $X2=1.78 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_4%Y 1 2 3 4 5 6 7 8 9 10 33 35 36 39 42 43
+ 47 49 53 55 59 61 65 67 71 73 77 79 80 81 82 83 84 85 86 92
c192 42 0 1.10003e-19 $X=3.35 $Y=1.415
r193 89 92 29.2085 $w=2.88e-07 $l=7.35e-07 $layer=LI1_cond $X=2.25 $Y=1.56
+ $X2=2.985 $Y2=1.56
r194 86 95 7.74919 $w=2.88e-07 $l=1.95e-07 $layer=LI1_cond $X=2.995 $Y=1.56
+ $X2=3.19 $Y2=1.56
r195 86 92 0.397394 $w=2.88e-07 $l=1e-08 $layer=LI1_cond $X=2.995 $Y=1.56
+ $X2=2.985 $Y2=1.56
r196 80 95 2.98046 $w=2.88e-07 $l=7.5e-08 $layer=LI1_cond $X=3.265 $Y=1.56
+ $X2=3.19 $Y2=1.56
r197 75 77 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=9.325 $Y=0.725
+ $X2=9.325 $Y2=0.39
r198 74 85 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=8.575 $Y=0.815
+ $X2=8.385 $Y2=0.815
r199 73 75 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=9.135 $Y=0.815
+ $X2=9.325 $Y2=0.725
r200 73 74 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=9.135 $Y=0.815
+ $X2=8.575 $Y2=0.815
r201 69 85 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=8.385 $Y=0.725
+ $X2=8.385 $Y2=0.815
r202 69 71 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=8.385 $Y=0.725
+ $X2=8.385 $Y2=0.39
r203 68 84 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=7.635 $Y=0.815
+ $X2=7.445 $Y2=0.815
r204 67 85 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=8.195 $Y=0.815
+ $X2=8.385 $Y2=0.815
r205 67 68 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=8.195 $Y=0.815
+ $X2=7.635 $Y2=0.815
r206 63 84 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=7.445 $Y=0.725
+ $X2=7.445 $Y2=0.815
r207 63 65 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.445 $Y=0.725
+ $X2=7.445 $Y2=0.39
r208 62 83 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.695 $Y=0.815
+ $X2=6.505 $Y2=0.815
r209 61 84 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=7.255 $Y=0.815
+ $X2=7.445 $Y2=0.815
r210 61 62 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=7.255 $Y=0.815
+ $X2=6.695 $Y2=0.815
r211 57 83 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=6.505 $Y=0.725
+ $X2=6.505 $Y2=0.815
r212 57 59 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.505 $Y=0.725
+ $X2=6.505 $Y2=0.39
r213 56 82 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.235 $Y=0.815
+ $X2=5.045 $Y2=0.815
r214 55 83 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.315 $Y=0.815
+ $X2=6.505 $Y2=0.815
r215 55 56 66.5455 $w=1.78e-07 $l=1.08e-06 $layer=LI1_cond $X=6.315 $Y=0.815
+ $X2=5.235 $Y2=0.815
r216 51 82 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=5.045 $Y=0.725
+ $X2=5.045 $Y2=0.815
r217 51 53 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.045 $Y=0.725
+ $X2=5.045 $Y2=0.39
r218 50 81 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.295 $Y=0.815
+ $X2=4.105 $Y2=0.815
r219 49 82 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.855 $Y=0.815
+ $X2=5.045 $Y2=0.815
r220 49 50 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.855 $Y=0.815
+ $X2=4.295 $Y2=0.815
r221 45 81 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=4.105 $Y=0.725
+ $X2=4.105 $Y2=0.815
r222 45 47 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.105 $Y=0.725
+ $X2=4.105 $Y2=0.39
r223 44 79 4.43084 $w=1.8e-07 $l=2.3e-07 $layer=LI1_cond $X=3.435 $Y=0.815
+ $X2=3.205 $Y2=0.815
r224 43 81 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.915 $Y=0.815
+ $X2=4.105 $Y2=0.815
r225 43 44 29.5758 $w=1.78e-07 $l=4.8e-07 $layer=LI1_cond $X=3.915 $Y=0.815
+ $X2=3.435 $Y2=0.815
r226 42 80 7.43784 $w=2.9e-07 $l=1.8262e-07 $layer=LI1_cond $X=3.35 $Y=1.415
+ $X2=3.265 $Y2=1.56
r227 41 79 1.86605 $w=1.7e-07 $l=1.84594e-07 $layer=LI1_cond $X=3.35 $Y=0.905
+ $X2=3.205 $Y2=0.815
r228 41 42 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.35 $Y=0.905
+ $X2=3.35 $Y2=1.415
r229 37 79 1.86605 $w=3.8e-07 $l=1.08167e-07 $layer=LI1_cond $X=3.165 $Y=0.725
+ $X2=3.205 $Y2=0.815
r230 37 39 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.165 $Y=0.725
+ $X2=3.165 $Y2=0.39
r231 35 79 4.43084 $w=1.8e-07 $l=2.3e-07 $layer=LI1_cond $X=2.975 $Y=0.815
+ $X2=3.205 $Y2=0.815
r232 35 36 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=2.975 $Y=0.815
+ $X2=2.415 $Y2=0.815
r233 31 36 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=2.225 $Y=0.725
+ $X2=2.415 $Y2=0.815
r234 31 33 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.225 $Y=0.725
+ $X2=2.225 $Y2=0.39
r235 10 95 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.045
+ $Y=1.485 $X2=3.19 $Y2=1.62
r236 9 89 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.105
+ $Y=1.485 $X2=2.25 $Y2=1.62
r237 8 77 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=9.165
+ $Y=0.235 $X2=9.35 $Y2=0.39
r238 7 71 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=8.225
+ $Y=0.235 $X2=8.41 $Y2=0.39
r239 6 65 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=7.285
+ $Y=0.235 $X2=7.47 $Y2=0.39
r240 5 59 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=6.345
+ $Y=0.235 $X2=6.53 $Y2=0.39
r241 4 53 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.885
+ $Y=0.235 $X2=5.07 $Y2=0.39
r242 3 47 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.945
+ $Y=0.235 $X2=4.13 $Y2=0.39
r243 2 39 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.005
+ $Y=0.235 $X2=3.19 $Y2=0.39
r244 1 33 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=2.065
+ $Y=0.235 $X2=2.25 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_4%A_797_297# 1 2 3 4 15 19 23 28 30 32 34
r61 24 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.655 $Y=1.54
+ $X2=6.53 $Y2=1.54
r62 23 34 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.345 $Y=1.54
+ $X2=7.47 $Y2=1.54
r63 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.345 $Y=1.54
+ $X2=6.655 $Y2=1.54
r64 20 30 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.195 $Y=1.54
+ $X2=5.07 $Y2=1.54
r65 19 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.405 $Y=1.54
+ $X2=6.53 $Y2=1.54
r66 19 20 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=6.405 $Y=1.54
+ $X2=5.195 $Y2=1.54
r67 16 28 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.255 $Y=1.54
+ $X2=4.15 $Y2=1.54
r68 15 30 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.945 $Y=1.54
+ $X2=5.07 $Y2=1.54
r69 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.945 $Y=1.54
+ $X2=4.255 $Y2=1.54
r70 4 34 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=7.325
+ $Y=1.485 $X2=7.47 $Y2=1.62
r71 3 32 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.385
+ $Y=1.485 $X2=6.53 $Y2=1.62
r72 2 30 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=4.925
+ $Y=1.485 $X2=5.07 $Y2=1.62
r73 1 28 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.985
+ $Y=1.485 $X2=4.13 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_4%A_1187_297# 1 2 3 4 5 18 20 21 24 26 28
+ 29 30 34 36 38 40 42 48
r63 38 50 2.68365 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=9.852 $Y=1.625
+ $X2=9.852 $Y2=1.54
r64 38 40 24.6952 $w=3.13e-07 $l=6.75e-07 $layer=LI1_cond $X=9.852 $Y=1.625
+ $X2=9.852 $Y2=2.3
r65 37 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.005 $Y=1.54
+ $X2=8.88 $Y2=1.54
r66 36 50 4.95685 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=9.695 $Y=1.54
+ $X2=9.852 $Y2=1.54
r67 36 37 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.695 $Y=1.54
+ $X2=9.005 $Y2=1.54
r68 32 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.88 $Y=1.625
+ $X2=8.88 $Y2=1.54
r69 32 34 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=8.88 $Y=1.625
+ $X2=8.88 $Y2=2.3
r70 31 44 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.065 $Y=1.54
+ $X2=7.94 $Y2=1.54
r71 30 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.755 $Y=1.54
+ $X2=8.88 $Y2=1.54
r72 30 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.755 $Y=1.54
+ $X2=8.065 $Y2=1.54
r73 29 46 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.94 $Y=2.295
+ $X2=7.94 $Y2=2.38
r74 28 44 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.94 $Y=1.625
+ $X2=7.94 $Y2=1.54
r75 28 29 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=7.94 $Y=1.625
+ $X2=7.94 $Y2=2.295
r76 27 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.125 $Y=2.38 $X2=7
+ $Y2=2.38
r77 26 46 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.815 $Y=2.38
+ $X2=7.94 $Y2=2.38
r78 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.815 $Y=2.38
+ $X2=7.125 $Y2=2.38
r79 22 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7 $Y=2.295 $X2=7
+ $Y2=2.38
r80 22 24 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=7 $Y=2.295 $X2=7
+ $Y2=1.96
r81 20 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.875 $Y=2.38 $X2=7
+ $Y2=2.38
r82 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.875 $Y=2.38
+ $X2=6.185 $Y2=2.38
r83 16 21 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=6.032 $Y=2.295
+ $X2=6.185 $Y2=2.38
r84 16 18 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=6.032 $Y=2.295
+ $X2=6.032 $Y2=1.96
r85 5 50 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.675
+ $Y=1.485 $X2=9.82 $Y2=1.62
r86 5 40 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=9.675
+ $Y=1.485 $X2=9.82 $Y2=2.3
r87 4 48 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.735
+ $Y=1.485 $X2=8.88 $Y2=1.62
r88 4 34 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=8.735
+ $Y=1.485 $X2=8.88 $Y2=2.3
r89 3 46 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=7.795
+ $Y=1.485 $X2=7.94 $Y2=2.3
r90 3 44 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.795
+ $Y=1.485 $X2=7.94 $Y2=1.62
r91 2 24 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.855
+ $Y=1.485 $X2=7 $Y2=1.96
r92 1 18 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=5.935
+ $Y=1.485 $X2=6.06 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_4%VGND 1 2 3 4 5 6 7 8 9 10 35 39 43 47 51
+ 55 59 63 65 67 70 71 73 74 76 77 79 80 82 83 85 86 88 89 90 119 124 129 132
+ 135 137
r167 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r168 131 132 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=6.06 $Y=0.235
+ $X2=6.145 $Y2=0.235
r169 127 131 5.7935 $w=6.38e-07 $l=3.1e-07 $layer=LI1_cond $X=5.75 $Y=0.235
+ $X2=6.06 $Y2=0.235
r170 127 129 12.8464 $w=6.38e-07 $l=2.95e-07 $layer=LI1_cond $X=5.75 $Y=0.235
+ $X2=5.455 $Y2=0.235
r171 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r172 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r173 122 135 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=9.89 $Y2=0
r174 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r175 119 134 4.23443 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=9.735 $Y=0
+ $X2=9.927 $Y2=0
r176 119 121 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.735 $Y=0
+ $X2=9.43 $Y2=0
r177 118 122 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=9.43 $Y2=0
r178 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r179 115 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.51 $Y2=0
r180 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r181 112 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r182 112 128 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=5.75 $Y2=0
r183 111 132 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=6.67 $Y=0
+ $X2=6.145 $Y2=0
r184 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r185 108 128 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=5.75 $Y2=0
r186 107 129 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.29 $Y=0
+ $X2=5.455 $Y2=0
r187 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r188 104 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.29 $Y2=0
r189 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r190 101 104 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.37 $Y2=0
r191 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r192 98 101 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.45 $Y2=0
r193 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r194 95 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r195 95 125 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=0.69 $Y2=0
r196 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r197 92 124 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=0 $X2=0.75
+ $Y2=0
r198 92 94 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.835 $Y=0
+ $X2=1.61 $Y2=0
r199 90 125 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r200 90 137 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r201 88 117 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.795 $Y=0
+ $X2=8.51 $Y2=0
r202 88 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.795 $Y=0 $X2=8.88
+ $Y2=0
r203 87 121 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=8.965 $Y=0
+ $X2=9.43 $Y2=0
r204 87 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.965 $Y=0 $X2=8.88
+ $Y2=0
r205 85 114 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.855 $Y=0
+ $X2=7.59 $Y2=0
r206 85 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.855 $Y=0 $X2=7.94
+ $Y2=0
r207 84 117 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=8.025 $Y=0
+ $X2=8.51 $Y2=0
r208 84 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.025 $Y=0 $X2=7.94
+ $Y2=0
r209 82 111 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.915 $Y=0
+ $X2=6.67 $Y2=0
r210 82 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.915 $Y=0 $X2=7
+ $Y2=0
r211 81 114 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=7.085 $Y=0
+ $X2=7.59 $Y2=0
r212 81 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.085 $Y=0 $X2=7
+ $Y2=0
r213 79 103 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.515 $Y=0
+ $X2=4.37 $Y2=0
r214 79 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.515 $Y=0 $X2=4.6
+ $Y2=0
r215 78 107 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.685 $Y=0
+ $X2=5.29 $Y2=0
r216 78 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.685 $Y=0 $X2=4.6
+ $Y2=0
r217 76 100 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.575 $Y=0
+ $X2=3.45 $Y2=0
r218 76 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.575 $Y=0 $X2=3.66
+ $Y2=0
r219 75 103 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.745 $Y=0
+ $X2=4.37 $Y2=0
r220 75 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.745 $Y=0 $X2=3.66
+ $Y2=0
r221 73 97 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.635 $Y=0
+ $X2=2.53 $Y2=0
r222 73 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=0 $X2=2.72
+ $Y2=0
r223 72 100 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=2.805 $Y=0
+ $X2=3.45 $Y2=0
r224 72 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.805 $Y=0 $X2=2.72
+ $Y2=0
r225 70 94 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=0 $X2=1.61
+ $Y2=0
r226 70 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=0 $X2=1.78
+ $Y2=0
r227 69 97 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.53
+ $Y2=0
r228 69 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.78
+ $Y2=0
r229 65 134 3.08761 $w=2.75e-07 $l=1.09087e-07 $layer=LI1_cond $X=9.872 $Y=0.085
+ $X2=9.927 $Y2=0
r230 65 67 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=9.872 $Y=0.085
+ $X2=9.872 $Y2=0.39
r231 61 89 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.88 $Y=0.085
+ $X2=8.88 $Y2=0
r232 61 63 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.88 $Y=0.085
+ $X2=8.88 $Y2=0.39
r233 57 86 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.94 $Y=0.085
+ $X2=7.94 $Y2=0
r234 57 59 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.94 $Y=0.085
+ $X2=7.94 $Y2=0.39
r235 53 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7 $Y=0.085 $X2=7
+ $Y2=0
r236 53 55 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7 $Y=0.085 $X2=7
+ $Y2=0.39
r237 49 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.6 $Y=0.085 $X2=4.6
+ $Y2=0
r238 49 51 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.6 $Y=0.085
+ $X2=4.6 $Y2=0.39
r239 45 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.66 $Y=0.085
+ $X2=3.66 $Y2=0
r240 45 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.66 $Y=0.085
+ $X2=3.66 $Y2=0.39
r241 41 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.72 $Y=0.085
+ $X2=2.72 $Y2=0
r242 41 43 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.72 $Y=0.085
+ $X2=2.72 $Y2=0.39
r243 37 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0
r244 37 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0.39
r245 33 124 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r246 33 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.39
r247 10 67 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=9.685
+ $Y=0.235 $X2=9.82 $Y2=0.39
r248 9 63 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=8.695
+ $Y=0.235 $X2=8.88 $Y2=0.39
r249 8 59 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.805
+ $Y=0.235 $X2=7.94 $Y2=0.39
r250 7 55 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=6.815
+ $Y=0.235 $X2=7 $Y2=0.39
r251 6 131 91 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_NDIFF $count=2 $X=5.405
+ $Y=0.235 $X2=6.06 $Y2=0.39
r252 5 51 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.415
+ $Y=0.235 $X2=4.6 $Y2=0.39
r253 4 47 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.525
+ $Y=0.235 $X2=3.66 $Y2=0.39
r254 3 43 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.235 $X2=2.72 $Y2=0.39
r255 2 39 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.655
+ $Y=0.235 $X2=1.78 $Y2=0.39
r256 1 35 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

