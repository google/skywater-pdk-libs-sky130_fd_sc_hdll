* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_455_21# a_211_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VPWR A1_N a_455_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_211_297# a_455_21# a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 X a_211_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 a_787_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR B1 a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 a_455_21# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 a_27_47# a_455_21# a_211_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_117_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_787_47# A2_N a_455_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 X a_211_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_211_297# B2 a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 X a_211_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR a_211_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 VGND B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 X a_211_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VPWR A2_N a_455_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 a_27_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_117_297# B2 a_211_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 VGND A1_N a_787_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VGND a_211_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR a_211_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 a_455_21# A2_N a_787_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VGND a_211_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_211_297# a_455_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X27 a_455_21# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
