* File: sky130_fd_sc_hdll__a21boi_2.spice
* Created: Thu Aug 27 18:52:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a21boi_2.pex.spice"
.subckt sky130_fd_sc_hdll__a21boi_2  VNB VPB B1_N A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_B1_N_M1010_g N_A_61_47#_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.164762 AS=0.147 PD=1.05196 PS=1.54 NRD=74.988 NRS=24.276 M=1 R=2.8
+ SA=75000.3 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1010_d N_A_61_47#_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.254988 AS=0.104 PD=1.62804 PS=0.97 NRD=27.684 NRS=0 M=1 R=4.33333
+ SA=75000.9 SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_A_61_47#_M1012_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.104 PD=1.03 PS=0.97 NRD=9.228 NRS=8.304 M=1 R=4.33333
+ SA=75001.4 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1012_d N_A2_M1009_g A_529_47# VNB NSHORT L=0.15 W=0.65 AD=0.1235
+ AS=0.06825 PD=1.03 PS=0.86 NRD=9.228 NRS=9.228 M=1 R=4.33333 SA=75001.9
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1004 A_529_47# N_A1_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65 AD=0.06825
+ AS=0.10725 PD=0.86 PS=0.98 NRD=9.228 NRS=9.228 M=1 R=4.33333 SA=75002.3
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1011 A_697_47# N_A1_M1011_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65 AD=0.10725
+ AS=0.10725 PD=0.98 PS=0.98 NRD=20.304 NRS=0 M=1 R=4.33333 SA=75002.7
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_A2_M1013_g A_697_47# VNB NSHORT L=0.15 W=0.65 AD=0.21775
+ AS=0.10725 PD=1.97 PS=0.98 NRD=9.228 NRS=20.304 M=1 R=4.33333 SA=75003.2
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1007 N_A_61_47#_M1007_d N_B1_N_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1155 AS=0.1155 PD=1.39 PS=1.39 NRD=4.6886 NRS=4.6886 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1003 N_A_228_297#_M1003_d N_A_61_47#_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.18
+ W=1 AD=0.315 AS=0.145 PD=2.63 PS=1.29 NRD=9.8303 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1005 N_A_228_297#_M1005_d N_A_61_47#_M1005_g N_Y_M1003_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A2_M1001_g N_A_228_297#_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1000 N_A_228_297#_M1000_d N_A1_M1000_g N_VPWR_M1001_d VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.145 PD=1.3 PS=1.29 NRD=1.9503 NRS=0.9653 M=1 R=5.55556 SA=90001.6
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1008 N_A_228_297#_M1000_d N_A1_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.1
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1008_s N_A2_M1002_g N_A_228_297#_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
pX15_noxref noxref_13 Y Y PROBETYPE=1
pX16_noxref noxref_14 A1 A1 PROBETYPE=1
pX17_noxref noxref_15 A2 A2 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__a21boi_2.pxi.spice"
*
.ends
*
*
