* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 a_121_297# B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=5.75e+11p pd=5.15e+06u as=2.75e+11p ps=2.55e+06u
M1001 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=4.095e+11p ps=3.86e+06u
M1002 a_219_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u
M1003 VPWR A1 a_121_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.15e+11p pd=2.63e+06u as=0p ps=0u
M1004 a_121_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A2 a_219_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
