* File: sky130_fd_sc_hdll__muxb16to1_1.pxi.spice
* Created: Wed Sep  2 08:35:15 2020
* 
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[0] N_D[0]_c_548_n N_D[0]_M1086_g
+ N_D[0]_c_549_n N_D[0]_M1027_g N_D[0]_c_550_n N_D[0]_c_551_n D[0]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[0]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[8] N_D[8]_c_577_n N_D[8]_M1025_g
+ N_D[8]_c_581_n N_D[8]_M1032_g N_D[8]_c_578_n N_D[8]_c_579_n D[8]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[8]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_184_265# N_A_184_265#_M1058_s
+ N_A_184_265#_M1045_s N_A_184_265#_M1036_g N_A_184_265#_c_608_n
+ N_A_184_265#_c_609_n N_A_184_265#_c_613_n N_A_184_265#_c_610_n
+ N_A_184_265#_c_611_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_184_265#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_184_793# N_A_184_793#_M1067_s
+ N_A_184_793#_M1048_s N_A_184_793#_M1090_g N_A_184_793#_c_666_n
+ N_A_184_793#_c_667_n N_A_184_793#_c_671_n N_A_184_793#_c_668_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_184_793#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[0] N_S[0]_c_722_n N_S[0]_M1092_g
+ N_S[0]_c_723_n N_S[0]_c_724_n N_S[0]_c_725_n N_S[0]_M1045_g N_S[0]_c_726_n
+ N_S[0]_M1058_g S[0] N_S[0]_c_727_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[0]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[8] N_S[8]_c_771_n N_S[8]_M1056_g
+ N_S[8]_c_772_n N_S[8]_c_773_n N_S[8]_c_776_n N_S[8]_M1048_g N_S[8]_c_774_n
+ N_S[8]_M1067_g S[8] PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[8]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[1] N_S[1]_c_819_n N_S[1]_M1039_g
+ N_S[1]_c_820_n N_S[1]_M1055_g N_S[1]_c_821_n N_S[1]_c_822_n N_S[1]_M1023_g
+ S[1] N_S[1]_c_823_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[1]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[9] N_S[9]_c_869_n N_S[9]_M1042_g
+ N_S[9]_c_865_n N_S[9]_M1031_g N_S[9]_c_866_n N_S[9]_c_867_n N_S[9]_M1047_g
+ S[9] PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[9]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_533_47# N_A_533_47#_M1055_d
+ N_A_533_47#_M1039_d N_A_533_47#_M1017_g N_A_533_47#_c_917_n
+ N_A_533_47#_c_912_n N_A_533_47#_c_913_n N_A_533_47#_c_914_n
+ N_A_533_47#_c_915_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_533_47#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_533_937# N_A_533_937#_M1031_d
+ N_A_533_937#_M1042_d N_A_533_937#_M1071_g N_A_533_937#_c_974_n
+ N_A_533_937#_c_969_n N_A_533_937#_c_970_n N_A_533_937#_c_971_n
+ N_A_533_937#_c_972_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_533_937#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[1] N_D[1]_c_1028_n N_D[1]_M1075_g
+ N_D[1]_c_1029_n N_D[1]_M1062_g N_D[1]_c_1030_n N_D[1]_c_1031_n D[1]
+ N_D[1]_c_1061_p PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[1]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[9] N_D[9]_c_1069_n N_D[9]_M1076_g
+ N_D[9]_c_1066_n N_D[9]_M1057_g N_D[9]_c_1067_n N_D[9]_c_1068_n D[9]
+ N_D[9]_c_1102_p PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[9]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[2] N_D[2]_c_1107_n N_D[2]_M1002_g
+ N_D[2]_c_1108_n N_D[2]_M1040_g N_D[2]_c_1109_n N_D[2]_c_1110_n D[2]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[2]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[10] N_D[10]_c_1145_n N_D[10]_M1011_g
+ N_D[10]_c_1149_n N_D[10]_M1044_g N_D[10]_c_1146_n N_D[10]_c_1147_n D[10]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[10]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1012_265# N_A_1012_265#_M1088_s
+ N_A_1012_265#_M1050_s N_A_1012_265#_M1041_g N_A_1012_265#_c_1186_n
+ N_A_1012_265#_c_1187_n N_A_1012_265#_c_1191_n N_A_1012_265#_c_1188_n
+ N_A_1012_265#_c_1189_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1012_265#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1012_793# N_A_1012_793#_M1082_s
+ N_A_1012_793#_M1053_s N_A_1012_793#_M1000_g N_A_1012_793#_c_1244_n
+ N_A_1012_793#_c_1245_n N_A_1012_793#_c_1249_n N_A_1012_793#_c_1246_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1012_793#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[2] N_S[2]_c_1300_n N_S[2]_M1018_g
+ N_S[2]_c_1301_n N_S[2]_c_1302_n N_S[2]_c_1303_n N_S[2]_M1050_g N_S[2]_c_1304_n
+ N_S[2]_M1088_g S[2] N_S[2]_c_1305_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[2]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[10] N_S[10]_c_1349_n N_S[10]_M1065_g
+ N_S[10]_c_1350_n N_S[10]_c_1351_n N_S[10]_c_1354_n N_S[10]_M1053_g
+ N_S[10]_c_1352_n N_S[10]_M1082_g S[10] PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[10]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[3] N_S[3]_c_1397_n N_S[3]_M1009_g
+ N_S[3]_c_1398_n N_S[3]_M1052_g N_S[3]_c_1399_n N_S[3]_c_1400_n N_S[3]_M1015_g
+ S[3] N_S[3]_c_1401_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[3]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[11] N_S[11]_c_1447_n N_S[11]_M1012_g
+ N_S[11]_c_1443_n N_S[11]_M1061_g N_S[11]_c_1444_n N_S[11]_c_1445_n
+ N_S[11]_M1068_g S[11] PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[11]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1361_47# N_A_1361_47#_M1052_d
+ N_A_1361_47#_M1009_d N_A_1361_47#_M1022_g N_A_1361_47#_c_1495_n
+ N_A_1361_47#_c_1490_n N_A_1361_47#_c_1491_n N_A_1361_47#_c_1492_n
+ N_A_1361_47#_c_1493_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1361_47#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1361_937# N_A_1361_937#_M1061_d
+ N_A_1361_937#_M1012_d N_A_1361_937#_M1074_g N_A_1361_937#_c_1552_n
+ N_A_1361_937#_c_1547_n N_A_1361_937#_c_1548_n N_A_1361_937#_c_1549_n
+ N_A_1361_937#_c_1550_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1361_937#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[3] N_D[3]_c_1606_n N_D[3]_M1028_g
+ N_D[3]_c_1607_n N_D[3]_M1081_g N_D[3]_c_1608_n N_D[3]_c_1609_n D[3]
+ N_D[3]_c_1639_p PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[3]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[11] N_D[11]_c_1647_n N_D[11]_M1033_g
+ N_D[11]_c_1644_n N_D[11]_M1043_g N_D[11]_c_1645_n N_D[11]_c_1646_n D[11]
+ N_D[11]_c_1680_p PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[11]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[4] N_D[4]_c_1685_n N_D[4]_M1001_g
+ N_D[4]_c_1686_n N_D[4]_M1005_g N_D[4]_c_1687_n N_D[4]_c_1688_n D[4]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[4]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[12] N_D[12]_c_1723_n N_D[12]_M1037_g
+ N_D[12]_c_1727_n N_D[12]_M1006_g N_D[12]_c_1724_n N_D[12]_c_1725_n D[12]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[12]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1840_265# N_A_1840_265#_M1094_s
+ N_A_1840_265#_M1080_s N_A_1840_265#_M1014_g N_A_1840_265#_c_1764_n
+ N_A_1840_265#_c_1765_n N_A_1840_265#_c_1769_n N_A_1840_265#_c_1766_n
+ N_A_1840_265#_c_1767_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1840_265#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1840_793# N_A_1840_793#_M1024_s
+ N_A_1840_793#_M1085_s N_A_1840_793#_M1064_g N_A_1840_793#_c_1822_n
+ N_A_1840_793#_c_1823_n N_A_1840_793#_c_1827_n N_A_1840_793#_c_1824_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1840_793#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[4] N_S[4]_c_1878_n N_S[4]_M1030_g
+ N_S[4]_c_1879_n N_S[4]_c_1880_n N_S[4]_c_1881_n N_S[4]_M1080_g N_S[4]_c_1882_n
+ N_S[4]_M1094_g S[4] N_S[4]_c_1883_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[4]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[12] N_S[12]_c_1927_n N_S[12]_M1069_g
+ N_S[12]_c_1928_n N_S[12]_c_1929_n N_S[12]_c_1932_n N_S[12]_M1085_g
+ N_S[12]_c_1930_n N_S[12]_M1024_g S[12] PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[12]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[5] N_S[5]_c_1975_n N_S[5]_M1046_g
+ N_S[5]_c_1976_n N_S[5]_M1078_g N_S[5]_c_1977_n N_S[5]_c_1978_n N_S[5]_M1020_g
+ S[5] N_S[5]_c_1979_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[5]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[13] N_S[13]_c_2025_n N_S[13]_M1049_g
+ N_S[13]_c_2021_n N_S[13]_M1070_g N_S[13]_c_2022_n N_S[13]_c_2023_n
+ N_S[13]_M1016_g S[13] PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[13]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_2189_47# N_A_2189_47#_M1078_d
+ N_A_2189_47#_M1046_d N_A_2189_47#_M1059_g N_A_2189_47#_c_2073_n
+ N_A_2189_47#_c_2068_n N_A_2189_47#_c_2069_n N_A_2189_47#_c_2070_n
+ N_A_2189_47#_c_2071_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_2189_47#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_2189_937# N_A_2189_937#_M1070_d
+ N_A_2189_937#_M1049_d N_A_2189_937#_M1008_g N_A_2189_937#_c_2130_n
+ N_A_2189_937#_c_2125_n N_A_2189_937#_c_2126_n N_A_2189_937#_c_2127_n
+ N_A_2189_937#_c_2128_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_2189_937#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[5] N_D[5]_c_2184_n N_D[5]_M1077_g
+ N_D[5]_c_2185_n N_D[5]_M1087_g N_D[5]_c_2186_n N_D[5]_c_2187_n D[5]
+ N_D[5]_c_2217_p PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[5]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[13] N_D[13]_c_2225_n N_D[13]_M1079_g
+ N_D[13]_c_2222_n N_D[13]_M1091_g N_D[13]_c_2223_n N_D[13]_c_2224_n D[13]
+ N_D[13]_c_2258_p PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[13]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[6] N_D[6]_c_2263_n N_D[6]_M1003_g
+ N_D[6]_c_2264_n N_D[6]_M1029_g N_D[6]_c_2265_n N_D[6]_c_2266_n D[6]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[6]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[14] N_D[14]_c_2301_n N_D[14]_M1083_g
+ N_D[14]_c_2305_n N_D[14]_M1035_g N_D[14]_c_2302_n N_D[14]_c_2303_n D[14]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[14]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_2668_265# N_A_2668_265#_M1007_s
+ N_A_2668_265#_M1066_s N_A_2668_265#_M1051_g N_A_2668_265#_c_2342_n
+ N_A_2668_265#_c_2343_n N_A_2668_265#_c_2347_n N_A_2668_265#_c_2344_n
+ N_A_2668_265#_c_2345_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_2668_265#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_2668_793# N_A_2668_793#_M1026_s
+ N_A_2668_793#_M1072_s N_A_2668_793#_M1004_g N_A_2668_793#_c_2400_n
+ N_A_2668_793#_c_2401_n N_A_2668_793#_c_2405_n N_A_2668_793#_c_2402_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_2668_793#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[6] N_S[6]_c_2456_n N_S[6]_M1063_g
+ N_S[6]_c_2457_n N_S[6]_c_2458_n N_S[6]_c_2459_n N_S[6]_M1066_g N_S[6]_c_2460_n
+ N_S[6]_M1007_g S[6] N_S[6]_c_2461_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[6]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[14] N_S[14]_c_2505_n N_S[14]_M1084_g
+ N_S[14]_c_2506_n N_S[14]_c_2507_n N_S[14]_c_2510_n N_S[14]_M1072_g
+ N_S[14]_c_2508_n N_S[14]_M1026_g S[14] PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[14]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[7] N_S[7]_c_2553_n N_S[7]_M1019_g
+ N_S[7]_c_2554_n N_S[7]_M1095_g N_S[7]_c_2555_n N_S[7]_c_2556_n N_S[7]_M1060_g
+ S[7] N_S[7]_c_2557_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[7]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[15] N_S[15]_c_2603_n N_S[15]_M1021_g
+ N_S[15]_c_2599_n N_S[15]_M1073_g N_S[15]_c_2600_n N_S[15]_c_2601_n
+ N_S[15]_M1054_g S[15] PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[15]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_3017_47# N_A_3017_47#_M1095_d
+ N_A_3017_47#_M1019_d N_A_3017_47#_M1093_g N_A_3017_47#_c_2651_n
+ N_A_3017_47#_c_2646_n N_A_3017_47#_c_2647_n N_A_3017_47#_c_2648_n
+ N_A_3017_47#_c_2649_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_3017_47#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_3017_937# N_A_3017_937#_M1073_d
+ N_A_3017_937#_M1021_d N_A_3017_937#_M1038_g N_A_3017_937#_c_2708_n
+ N_A_3017_937#_c_2703_n N_A_3017_937#_c_2704_n N_A_3017_937#_c_2705_n
+ N_A_3017_937#_c_2706_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_3017_937#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[7] N_D[7]_c_2762_n N_D[7]_M1010_g
+ N_D[7]_c_2763_n N_D[7]_M1089_g N_D[7]_c_2764_n N_D[7]_c_2765_n D[7]
+ N_D[7]_c_2786_p PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[7]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[15] N_D[15]_c_2794_n N_D[15]_M1013_g
+ N_D[15]_c_2791_n N_D[15]_M1034_g N_D[15]_c_2792_n N_D[15]_c_2793_n D[15]
+ N_D[15]_c_2817_p PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[15]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%VPWR N_VPWR_M1027_s N_VPWR_M1032_s
+ N_VPWR_M1045_d N_VPWR_M1048_d N_VPWR_M1075_d N_VPWR_M1076_d N_VPWR_M1050_d
+ N_VPWR_M1053_d N_VPWR_M1028_d N_VPWR_M1033_d N_VPWR_M1080_d N_VPWR_M1085_d
+ N_VPWR_M1077_d N_VPWR_M1079_d N_VPWR_M1066_d N_VPWR_M1072_d N_VPWR_M1010_d
+ N_VPWR_M1013_d N_VPWR_c_2822_n N_VPWR_c_2823_n N_VPWR_c_2824_n N_VPWR_c_2825_n
+ N_VPWR_c_2826_n N_VPWR_c_2827_n N_VPWR_c_2828_n N_VPWR_c_2829_n
+ N_VPWR_c_2830_n N_VPWR_c_2831_n N_VPWR_c_2832_n N_VPWR_c_2833_n
+ N_VPWR_c_2834_n N_VPWR_c_2835_n N_VPWR_c_2836_n N_VPWR_c_2837_n
+ N_VPWR_c_2838_n N_VPWR_c_2839_n N_VPWR_c_2840_n N_VPWR_c_2841_n
+ N_VPWR_c_2842_n N_VPWR_c_2843_n N_VPWR_c_2844_n N_VPWR_c_2845_n
+ N_VPWR_c_2846_n N_VPWR_c_2847_n VPWR VPWR VPWR VPWR VPWR N_VPWR_c_2849_n
+ N_VPWR_c_2850_n N_VPWR_c_2851_n N_VPWR_c_2852_n N_VPWR_c_2853_n
+ N_VPWR_c_2854_n N_VPWR_c_2855_n N_VPWR_c_2856_n N_VPWR_c_2857_n
+ N_VPWR_c_2858_n N_VPWR_c_2859_n N_VPWR_c_2860_n N_VPWR_c_2861_n
+ N_VPWR_c_2862_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%VPWR
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%Z N_Z_M1092_d N_Z_M1056_d N_Z_M1023_s
+ N_Z_M1047_s N_Z_M1018_d N_Z_M1065_d N_Z_M1015_s N_Z_M1068_s N_Z_M1030_d
+ N_Z_M1069_d N_Z_M1020_s N_Z_M1016_s N_Z_M1063_d N_Z_M1084_d N_Z_M1060_s
+ N_Z_M1054_s N_Z_M1036_d N_Z_M1090_d N_Z_M1017_s N_Z_M1071_s N_Z_M1041_d
+ N_Z_M1000_d N_Z_M1022_s N_Z_M1074_s N_Z_M1014_d N_Z_M1064_d N_Z_M1059_s
+ N_Z_M1008_s N_Z_M1051_d N_Z_M1004_d N_Z_M1093_s N_Z_M1038_s N_Z_c_3315_n
+ N_Z_c_3316_n N_Z_c_3317_n N_Z_c_3318_n N_Z_c_3319_n N_Z_c_3320_n N_Z_c_3365_n
+ N_Z_c_3366_n N_Z_c_3367_n N_Z_c_3368_n N_Z_c_3321_n N_Z_c_3322_n N_Z_c_3323_n
+ N_Z_c_3324_n N_Z_c_3325_n N_Z_c_3326_n N_Z_c_3327_n N_Z_c_3328_n N_Z_c_3329_n
+ N_Z_c_3330_n N_Z_c_3373_n N_Z_c_3374_n N_Z_c_3375_n N_Z_c_3376_n N_Z_c_3331_n
+ N_Z_c_3332_n N_Z_c_3333_n N_Z_c_3334_n N_Z_c_3335_n N_Z_c_3336_n N_Z_c_3337_n
+ N_Z_c_3338_n N_Z_c_3339_n N_Z_c_3340_n N_Z_c_3381_n N_Z_c_3382_n N_Z_c_3383_n
+ N_Z_c_3384_n N_Z_c_3341_n N_Z_c_3342_n N_Z_c_3343_n N_Z_c_3344_n N_Z_c_3345_n
+ N_Z_c_3346_n N_Z_c_3347_n N_Z_c_3348_n N_Z_c_3349_n N_Z_c_3350_n N_Z_c_3389_n
+ N_Z_c_3390_n N_Z_c_3391_n N_Z_c_3392_n N_Z_c_3351_n N_Z_c_3352_n N_Z_c_3353_n
+ N_Z_c_3354_n N_Z_c_3395_n N_Z_c_3396_n N_Z_c_3397_n N_Z_c_3398_n N_Z_c_3399_n
+ N_Z_c_3400_n N_Z_c_3355_n N_Z_c_3356_n N_Z_c_3401_n N_Z_c_3402_n N_Z_c_3403_n
+ N_Z_c_3404_n N_Z_c_3405_n N_Z_c_3406_n N_Z_c_3357_n N_Z_c_3358_n N_Z_c_3407_n
+ N_Z_c_3408_n N_Z_c_3409_n N_Z_c_3410_n N_Z_c_3411_n N_Z_c_3412_n N_Z_c_3359_n
+ N_Z_c_3360_n N_Z_c_3413_n N_Z_c_3414_n N_Z_c_3415_n N_Z_c_3416_n N_Z_c_3417_n
+ N_Z_c_3418_n N_Z_c_3361_n N_Z_c_3362_n N_Z_c_3419_n N_Z_c_3472_n N_Z_c_3420_n
+ N_Z_c_3494_n N_Z_c_3585_n N_Z_c_3549_n N_Z_c_3595_n N_Z_c_3572_n N_Z_c_3421_n
+ N_Z_c_3635_n N_Z_c_3422_n N_Z_c_3657_n N_Z_c_3748_n N_Z_c_3712_n N_Z_c_3758_n
+ N_Z_c_3735_n N_Z_c_3423_n N_Z_c_3798_n N_Z_c_3424_n N_Z_c_3820_n N_Z_c_3911_n
+ N_Z_c_3875_n N_Z_c_3921_n N_Z_c_3898_n N_Z_c_3425_n N_Z_c_3961_n N_Z_c_3426_n
+ N_Z_c_3983_n Z Z Z Z Z Z Z Z Z Z Z Z Z Z Z Z N_Z_c_3427_n N_Z_c_3428_n
+ N_Z_c_3429_n N_Z_c_3430_n N_Z_c_3431_n N_Z_c_3432_n N_Z_c_3433_n N_Z_c_3434_n
+ N_Z_c_3435_n N_Z_c_3436_n N_Z_c_3437_n N_Z_c_3438_n N_Z_c_3439_n N_Z_c_3440_n
+ N_Z_c_3441_n N_Z_c_3442_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%Z
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%VGND N_VGND_M1086_s N_VGND_M1025_s
+ N_VGND_M1058_d N_VGND_M1067_d N_VGND_M1062_d N_VGND_M1057_d N_VGND_M1088_d
+ N_VGND_M1082_d N_VGND_M1081_d N_VGND_M1043_d N_VGND_M1094_d N_VGND_M1024_d
+ N_VGND_M1087_d N_VGND_M1091_d N_VGND_M1007_d N_VGND_M1026_d N_VGND_M1089_d
+ N_VGND_M1034_d N_VGND_c_4367_n N_VGND_c_4368_n N_VGND_c_4369_n N_VGND_c_4370_n
+ N_VGND_c_4371_n N_VGND_c_4372_n N_VGND_c_4373_n N_VGND_c_4374_n
+ N_VGND_c_4375_n N_VGND_c_4376_n N_VGND_c_4377_n N_VGND_c_4378_n
+ N_VGND_c_4379_n N_VGND_c_4380_n N_VGND_c_4381_n N_VGND_c_4382_n
+ N_VGND_c_4383_n N_VGND_c_4384_n N_VGND_c_4385_n N_VGND_c_4386_n
+ N_VGND_c_4387_n N_VGND_c_4388_n N_VGND_c_4389_n N_VGND_c_4390_n
+ N_VGND_c_4391_n N_VGND_c_4392_n N_VGND_c_4393_n N_VGND_c_4394_n
+ N_VGND_c_4395_n N_VGND_c_4396_n N_VGND_c_4397_n N_VGND_c_4398_n
+ N_VGND_c_4399_n N_VGND_c_4400_n N_VGND_c_4401_n N_VGND_c_4402_n
+ N_VGND_c_4403_n N_VGND_c_4404_n VGND VGND VGND VGND VGND VGND VGND VGND VGND
+ VGND N_VGND_c_4407_n N_VGND_c_4408_n N_VGND_c_4409_n N_VGND_c_4410_n
+ N_VGND_c_4411_n N_VGND_c_4412_n N_VGND_c_4413_n N_VGND_c_4414_n
+ N_VGND_c_4415_n N_VGND_c_4416_n N_VGND_c_4417_n N_VGND_c_4418_n
+ N_VGND_c_4419_n N_VGND_c_4420_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%VGND
cc_1 VNB N_D[0]_c_548_n 0.0226847f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_D[0]_c_549_n 0.0309471f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_3 VNB N_D[0]_c_550_n 0.00249376f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_4 VNB N_D[0]_c_551_n 0.012124f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.19
cc_5 VNB N_D[8]_c_577_n 0.0536318f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_6 VNB N_D[8]_c_578_n 0.00249376f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_7 VNB N_D[8]_c_579_n 0.012124f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.19
cc_8 VNB N_A_184_265#_c_608_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_9 VNB N_A_184_265#_c_609_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_184_265#_c_610_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_184_265#_c_611_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_184_793#_c_666_n 0.013798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_184_793#_c_667_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.19
cc_14 VNB N_A_184_793#_c_668_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_S[0]_c_722_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_16 VNB N_S[0]_c_723_n 0.0502713f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_17 VNB N_S[0]_c_724_n 0.00937382f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_18 VNB N_S[0]_c_725_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_19 VNB N_S[0]_c_726_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_20 VNB N_S[0]_c_727_n 0.00873659f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_21 VNB N_S[8]_c_771_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_22 VNB N_S[8]_c_772_n 0.0502713f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_23 VNB N_S[8]_c_773_n 0.00937382f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_24 VNB N_S[8]_c_774_n 0.051972f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_25 VNB S[8] 0.00873659f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_S[1]_c_819_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_27 VNB N_S[1]_c_820_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_28 VNB N_S[1]_c_821_n 0.0596452f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.625
cc_29 VNB N_S[1]_c_822_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_30 VNB N_S[1]_c_823_n 0.00873659f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_31 VNB N_S[9]_c_865_n 0.051972f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_32 VNB N_S[9]_c_866_n 0.0596452f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.625
cc_33 VNB N_S[9]_c_867_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_34 VNB S[9] 0.00873659f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_533_47#_c_912_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_533_47#_c_913_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_533_47#_c_914_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_533_47#_c_915_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_533_937#_c_969_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_533_937#_c_970_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_533_937#_c_971_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_533_937#_c_972_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_D[1]_c_1028_n 0.0251359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_44 VNB N_D[1]_c_1029_n 0.0174886f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_45 VNB N_D[1]_c_1030_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_46 VNB N_D[1]_c_1031_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_D[9]_c_1066_n 0.0426246f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_48 VNB N_D[9]_c_1067_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_49 VNB N_D[9]_c_1068_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_D[2]_c_1107_n 0.0174886f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_51 VNB N_D[2]_c_1108_n 0.0251359f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_52 VNB N_D[2]_c_1109_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_53 VNB N_D[2]_c_1110_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.19
cc_54 VNB N_D[10]_c_1145_n 0.0426246f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_55 VNB N_D[10]_c_1146_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_56 VNB N_D[10]_c_1147_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.19
cc_57 VNB N_A_1012_265#_c_1186_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_58 VNB N_A_1012_265#_c_1187_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_1012_265#_c_1188_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_1012_265#_c_1189_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_1012_793#_c_1244_n 0.013798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_1012_793#_c_1245_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0.645
+ $Y2=1.19
cc_63 VNB N_A_1012_793#_c_1246_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_S[2]_c_1300_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_65 VNB N_S[2]_c_1301_n 0.0502713f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_66 VNB N_S[2]_c_1302_n 0.00937382f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_67 VNB N_S[2]_c_1303_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_68 VNB N_S[2]_c_1304_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_69 VNB N_S[2]_c_1305_n 0.00873659f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_70 VNB N_S[10]_c_1349_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_71 VNB N_S[10]_c_1350_n 0.0502713f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_72 VNB N_S[10]_c_1351_n 0.00937382f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_73 VNB N_S[10]_c_1352_n 0.051972f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_74 VNB S[10] 0.00873659f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_S[3]_c_1397_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_76 VNB N_S[3]_c_1398_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_77 VNB N_S[3]_c_1399_n 0.0596452f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.625
cc_78 VNB N_S[3]_c_1400_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_79 VNB N_S[3]_c_1401_n 0.00873659f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_80 VNB N_S[11]_c_1443_n 0.051972f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_81 VNB N_S[11]_c_1444_n 0.0596452f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.625
cc_82 VNB N_S[11]_c_1445_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_83 VNB S[11] 0.00873659f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1361_47#_c_1490_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_1361_47#_c_1491_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_1361_47#_c_1492_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_1361_47#_c_1493_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_1361_937#_c_1547_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_1361_937#_c_1548_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_1361_937#_c_1549_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_1361_937#_c_1550_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_D[3]_c_1606_n 0.0251359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_93 VNB N_D[3]_c_1607_n 0.0174886f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_94 VNB N_D[3]_c_1608_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_95 VNB N_D[3]_c_1609_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_D[11]_c_1644_n 0.0426246f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_97 VNB N_D[11]_c_1645_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_98 VNB N_D[11]_c_1646_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_D[4]_c_1685_n 0.0174886f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_100 VNB N_D[4]_c_1686_n 0.0251359f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_101 VNB N_D[4]_c_1687_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_102 VNB N_D[4]_c_1688_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.19
cc_103 VNB N_D[12]_c_1723_n 0.0426246f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_104 VNB N_D[12]_c_1724_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_105 VNB N_D[12]_c_1725_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.19
cc_106 VNB N_A_1840_265#_c_1764_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_107 VNB N_A_1840_265#_c_1765_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_A_1840_265#_c_1766_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_A_1840_265#_c_1767_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_A_1840_793#_c_1822_n 0.013798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_A_1840_793#_c_1823_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0.645
+ $Y2=1.19
cc_112 VNB N_A_1840_793#_c_1824_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_S[4]_c_1878_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_114 VNB N_S[4]_c_1879_n 0.0502713f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_115 VNB N_S[4]_c_1880_n 0.00937382f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_116 VNB N_S[4]_c_1881_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_117 VNB N_S[4]_c_1882_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_118 VNB N_S[4]_c_1883_n 0.00873659f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_119 VNB N_S[12]_c_1927_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_120 VNB N_S[12]_c_1928_n 0.0502713f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_121 VNB N_S[12]_c_1929_n 0.00937382f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_122 VNB N_S[12]_c_1930_n 0.051972f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_123 VNB S[12] 0.00873659f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_S[5]_c_1975_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_125 VNB N_S[5]_c_1976_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_126 VNB N_S[5]_c_1977_n 0.0596452f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.625
cc_127 VNB N_S[5]_c_1978_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_128 VNB N_S[5]_c_1979_n 0.00873659f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_129 VNB N_S[13]_c_2021_n 0.051972f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_130 VNB N_S[13]_c_2022_n 0.0596452f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.625
cc_131 VNB N_S[13]_c_2023_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_132 VNB S[13] 0.00873659f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_133 VNB N_A_2189_47#_c_2068_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_134 VNB N_A_2189_47#_c_2069_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_135 VNB N_A_2189_47#_c_2070_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_136 VNB N_A_2189_47#_c_2071_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_137 VNB N_A_2189_937#_c_2125_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_138 VNB N_A_2189_937#_c_2126_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_139 VNB N_A_2189_937#_c_2127_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_140 VNB N_A_2189_937#_c_2128_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_141 VNB N_D[5]_c_2184_n 0.0251359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_142 VNB N_D[5]_c_2185_n 0.0174886f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_143 VNB N_D[5]_c_2186_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_144 VNB N_D[5]_c_2187_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_145 VNB N_D[13]_c_2222_n 0.0426246f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_146 VNB N_D[13]_c_2223_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_147 VNB N_D[13]_c_2224_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_148 VNB N_D[6]_c_2263_n 0.0174886f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_149 VNB N_D[6]_c_2264_n 0.0251359f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_150 VNB N_D[6]_c_2265_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_151 VNB N_D[6]_c_2266_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.19
cc_152 VNB N_D[14]_c_2301_n 0.0426246f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_153 VNB N_D[14]_c_2302_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_154 VNB N_D[14]_c_2303_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.19
cc_155 VNB N_A_2668_265#_c_2342_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_156 VNB N_A_2668_265#_c_2343_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_157 VNB N_A_2668_265#_c_2344_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_158 VNB N_A_2668_265#_c_2345_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_159 VNB N_A_2668_793#_c_2400_n 0.013798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_160 VNB N_A_2668_793#_c_2401_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0.645
+ $Y2=1.19
cc_161 VNB N_A_2668_793#_c_2402_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_162 VNB N_S[6]_c_2456_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_163 VNB N_S[6]_c_2457_n 0.0502713f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_164 VNB N_S[6]_c_2458_n 0.00937382f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_165 VNB N_S[6]_c_2459_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_166 VNB N_S[6]_c_2460_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_167 VNB N_S[6]_c_2461_n 0.00873659f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_168 VNB N_S[14]_c_2505_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_169 VNB N_S[14]_c_2506_n 0.0502713f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_170 VNB N_S[14]_c_2507_n 0.00937382f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_171 VNB N_S[14]_c_2508_n 0.051972f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_172 VNB S[14] 0.00873659f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_173 VNB N_S[7]_c_2553_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_174 VNB N_S[7]_c_2554_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_175 VNB N_S[7]_c_2555_n 0.0596452f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.625
cc_176 VNB N_S[7]_c_2556_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_177 VNB N_S[7]_c_2557_n 0.00873659f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_178 VNB N_S[15]_c_2599_n 0.051972f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_179 VNB N_S[15]_c_2600_n 0.0596452f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.625
cc_180 VNB N_S[15]_c_2601_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_181 VNB S[15] 0.00873659f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_182 VNB N_A_3017_47#_c_2646_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_183 VNB N_A_3017_47#_c_2647_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_184 VNB N_A_3017_47#_c_2648_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_185 VNB N_A_3017_47#_c_2649_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_186 VNB N_A_3017_937#_c_2703_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_187 VNB N_A_3017_937#_c_2704_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_188 VNB N_A_3017_937#_c_2705_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_189 VNB N_A_3017_937#_c_2706_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_190 VNB N_D[7]_c_2762_n 0.0309471f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_191 VNB N_D[7]_c_2763_n 0.0226847f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_192 VNB N_D[7]_c_2764_n 0.00249376f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_193 VNB N_D[7]_c_2765_n 0.012124f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_194 VNB N_D[15]_c_2791_n 0.0536318f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_195 VNB N_D[15]_c_2792_n 0.00249376f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_196 VNB N_D[15]_c_2793_n 0.012124f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_197 VNB N_Z_c_3315_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_198 VNB N_Z_c_3316_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_199 VNB N_Z_c_3317_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_200 VNB N_Z_c_3318_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_201 VNB N_Z_c_3319_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_202 VNB N_Z_c_3320_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_203 VNB N_Z_c_3321_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_204 VNB N_Z_c_3322_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_205 VNB N_Z_c_3323_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_206 VNB N_Z_c_3324_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_207 VNB N_Z_c_3325_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_208 VNB N_Z_c_3326_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_209 VNB N_Z_c_3327_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_210 VNB N_Z_c_3328_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_211 VNB N_Z_c_3329_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_212 VNB N_Z_c_3330_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_213 VNB N_Z_c_3331_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_214 VNB N_Z_c_3332_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_215 VNB N_Z_c_3333_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_216 VNB N_Z_c_3334_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_217 VNB N_Z_c_3335_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_218 VNB N_Z_c_3336_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_219 VNB N_Z_c_3337_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_220 VNB N_Z_c_3338_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_221 VNB N_Z_c_3339_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_222 VNB N_Z_c_3340_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_223 VNB N_Z_c_3341_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_224 VNB N_Z_c_3342_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_225 VNB N_Z_c_3343_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_226 VNB N_Z_c_3344_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_227 VNB N_Z_c_3345_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_228 VNB N_Z_c_3346_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_229 VNB N_Z_c_3347_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_230 VNB N_Z_c_3348_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_231 VNB N_Z_c_3349_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_232 VNB N_Z_c_3350_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_233 VNB N_Z_c_3351_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_234 VNB N_Z_c_3352_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_235 VNB N_Z_c_3353_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_236 VNB N_Z_c_3354_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_237 VNB N_Z_c_3355_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_238 VNB N_Z_c_3356_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_239 VNB N_Z_c_3357_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_240 VNB N_Z_c_3358_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_241 VNB N_Z_c_3359_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_242 VNB N_Z_c_3360_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_243 VNB N_Z_c_3361_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_244 VNB N_Z_c_3362_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_245 VNB N_VGND_c_4367_n 0.0113488f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_246 VNB N_VGND_c_4368_n 0.0320435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_247 VNB N_VGND_c_4369_n 0.0113229f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_248 VNB N_VGND_c_4370_n 0.0320435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_249 VNB N_VGND_c_4371_n 0.00561737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_250 VNB N_VGND_c_4372_n 0.00561737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_251 VNB N_VGND_c_4373_n 0.00902444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_252 VNB N_VGND_c_4374_n 0.00902444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_253 VNB N_VGND_c_4375_n 0.00561737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_254 VNB N_VGND_c_4376_n 0.00561737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_255 VNB N_VGND_c_4377_n 0.00902444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_256 VNB N_VGND_c_4378_n 0.00902444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_257 VNB N_VGND_c_4379_n 0.00561737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_258 VNB N_VGND_c_4380_n 0.00561737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_259 VNB N_VGND_c_4381_n 0.00902444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_260 VNB N_VGND_c_4382_n 0.00902444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_261 VNB N_VGND_c_4383_n 0.00561737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_262 VNB N_VGND_c_4384_n 0.00561737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_263 VNB N_VGND_c_4385_n 0.0113488f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_264 VNB N_VGND_c_4386_n 0.0320435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_265 VNB N_VGND_c_4387_n 0.0113229f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_266 VNB N_VGND_c_4388_n 0.0320435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_267 VNB N_VGND_c_4389_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_268 VNB N_VGND_c_4390_n 0.00634747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_269 VNB N_VGND_c_4391_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_270 VNB N_VGND_c_4392_n 0.00632158f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_271 VNB N_VGND_c_4393_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_272 VNB N_VGND_c_4394_n 0.00634747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_273 VNB N_VGND_c_4395_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_274 VNB N_VGND_c_4396_n 0.00632158f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_275 VNB N_VGND_c_4397_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_276 VNB N_VGND_c_4398_n 0.00634747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_277 VNB N_VGND_c_4399_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_278 VNB N_VGND_c_4400_n 0.00632158f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_279 VNB N_VGND_c_4401_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_280 VNB N_VGND_c_4402_n 0.00634747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_281 VNB N_VGND_c_4403_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_282 VNB N_VGND_c_4404_n 0.00632158f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_283 VNB VGND 0.799771f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_284 VNB VGND 0.799771f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_285 VNB N_VGND_c_4407_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_286 VNB N_VGND_c_4408_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_287 VNB N_VGND_c_4409_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_288 VNB N_VGND_c_4410_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_289 VNB N_VGND_c_4411_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_290 VNB N_VGND_c_4412_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_291 VNB N_VGND_c_4413_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_292 VNB N_VGND_c_4414_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_293 VNB N_VGND_c_4415_n 0.00615512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_294 VNB N_VGND_c_4416_n 0.00612923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_295 VNB N_VGND_c_4417_n 0.00615512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_296 VNB N_VGND_c_4418_n 0.00612923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_297 VNB N_VGND_c_4419_n 0.00615512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_298 VNB N_VGND_c_4420_n 0.00612923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_299 VPB N_D[0]_c_549_n 0.0294852f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_300 VPB N_D[0]_c_551_n 0.00458905f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_301 VPB N_D[8]_c_577_n 0.012746f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_302 VPB N_D[8]_c_581_n 0.0167392f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_303 VPB N_D[8]_c_579_n 0.00458905f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_304 VPB N_A_184_265#_M1036_g 0.0216418f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_305 VPB N_A_184_265#_c_613_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.425
cc_306 VPB N_A_184_265#_c_610_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_307 VPB N_A_184_265#_c_611_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_308 VPB N_A_184_793#_M1090_g 0.0216418f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_309 VPB N_A_184_793#_c_667_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_310 VPB N_A_184_793#_c_671_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.425
cc_311 VPB N_A_184_793#_c_668_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_312 VPB N_S[0]_c_725_n 0.0238468f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_313 VPB N_S[8]_c_776_n 0.01606f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_314 VPB N_S[8]_c_774_n 0.00778682f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_315 VPB N_S[1]_c_819_n 0.0238468f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_316 VPB N_S[9]_c_869_n 0.01606f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_317 VPB N_S[9]_c_865_n 0.00778682f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_318 VPB N_A_533_47#_M1017_g 0.0216418f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_319 VPB N_A_533_47#_c_917_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_320 VPB N_A_533_47#_c_913_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_321 VPB N_A_533_47#_c_914_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_322 VPB N_A_533_937#_M1071_g 0.0216418f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_323 VPB N_A_533_937#_c_974_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_324 VPB N_A_533_937#_c_970_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_325 VPB N_A_533_937#_c_971_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_326 VPB N_D[1]_c_1028_n 0.0226466f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_327 VPB N_D[1]_c_1031_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_328 VPB N_D[9]_c_1069_n 0.0131744f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_329 VPB N_D[9]_c_1066_n 0.00947228f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_330 VPB N_D[9]_c_1068_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_331 VPB N_D[2]_c_1108_n 0.0226466f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_332 VPB N_D[2]_c_1110_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_333 VPB N_D[10]_c_1145_n 0.00947228f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_334 VPB N_D[10]_c_1149_n 0.0131744f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_335 VPB N_D[10]_c_1147_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_336 VPB N_A_1012_265#_M1041_g 0.0216418f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_337 VPB N_A_1012_265#_c_1191_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.605
+ $Y2=0.425
cc_338 VPB N_A_1012_265#_c_1188_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_339 VPB N_A_1012_265#_c_1189_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_340 VPB N_A_1012_793#_M1000_g 0.0216418f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_341 VPB N_A_1012_793#_c_1245_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0.645
+ $Y2=1.19
cc_342 VPB N_A_1012_793#_c_1249_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.605
+ $Y2=0.425
cc_343 VPB N_A_1012_793#_c_1246_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_344 VPB N_S[2]_c_1303_n 0.0238468f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_345 VPB N_S[10]_c_1354_n 0.01606f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_346 VPB N_S[10]_c_1352_n 0.00778682f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_347 VPB N_S[3]_c_1397_n 0.0238468f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_348 VPB N_S[11]_c_1447_n 0.01606f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_349 VPB N_S[11]_c_1443_n 0.00778682f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_350 VPB N_A_1361_47#_M1022_g 0.0216418f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_351 VPB N_A_1361_47#_c_1495_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_352 VPB N_A_1361_47#_c_1491_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_353 VPB N_A_1361_47#_c_1492_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_354 VPB N_A_1361_937#_M1074_g 0.0216418f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_355 VPB N_A_1361_937#_c_1552_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.645
+ $Y2=1.19
cc_356 VPB N_A_1361_937#_c_1548_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_357 VPB N_A_1361_937#_c_1549_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_358 VPB N_D[3]_c_1606_n 0.0226466f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_359 VPB N_D[3]_c_1609_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_360 VPB N_D[11]_c_1647_n 0.0131744f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_361 VPB N_D[11]_c_1644_n 0.00947228f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_362 VPB N_D[11]_c_1646_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_363 VPB N_D[4]_c_1686_n 0.0226466f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_364 VPB N_D[4]_c_1688_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_365 VPB N_D[12]_c_1723_n 0.00947228f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_366 VPB N_D[12]_c_1727_n 0.0131744f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_367 VPB N_D[12]_c_1725_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_368 VPB N_A_1840_265#_M1014_g 0.0216418f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_369 VPB N_A_1840_265#_c_1769_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.605
+ $Y2=0.425
cc_370 VPB N_A_1840_265#_c_1766_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_371 VPB N_A_1840_265#_c_1767_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_372 VPB N_A_1840_793#_M1064_g 0.0216418f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_373 VPB N_A_1840_793#_c_1823_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0.645
+ $Y2=1.19
cc_374 VPB N_A_1840_793#_c_1827_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.605
+ $Y2=0.425
cc_375 VPB N_A_1840_793#_c_1824_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_376 VPB N_S[4]_c_1881_n 0.0238468f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_377 VPB N_S[12]_c_1932_n 0.01606f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_378 VPB N_S[12]_c_1930_n 0.00778682f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_379 VPB N_S[5]_c_1975_n 0.0238468f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_380 VPB N_S[13]_c_2025_n 0.01606f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_381 VPB N_S[13]_c_2021_n 0.00778682f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_382 VPB N_A_2189_47#_M1059_g 0.0216418f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_383 VPB N_A_2189_47#_c_2073_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_384 VPB N_A_2189_47#_c_2069_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_385 VPB N_A_2189_47#_c_2070_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_386 VPB N_A_2189_937#_M1008_g 0.0216418f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_387 VPB N_A_2189_937#_c_2130_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.645
+ $Y2=1.19
cc_388 VPB N_A_2189_937#_c_2126_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_389 VPB N_A_2189_937#_c_2127_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_390 VPB N_D[5]_c_2184_n 0.0226466f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_391 VPB N_D[5]_c_2187_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_392 VPB N_D[13]_c_2225_n 0.0131744f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_393 VPB N_D[13]_c_2222_n 0.00947228f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_394 VPB N_D[13]_c_2224_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_395 VPB N_D[6]_c_2264_n 0.0226466f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_396 VPB N_D[6]_c_2266_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_397 VPB N_D[14]_c_2301_n 0.00947228f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_398 VPB N_D[14]_c_2305_n 0.0131744f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_399 VPB N_D[14]_c_2303_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_400 VPB N_A_2668_265#_M1051_g 0.0216418f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_401 VPB N_A_2668_265#_c_2347_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.605
+ $Y2=0.425
cc_402 VPB N_A_2668_265#_c_2344_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_403 VPB N_A_2668_265#_c_2345_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_404 VPB N_A_2668_793#_M1004_g 0.0216418f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_405 VPB N_A_2668_793#_c_2401_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0.645
+ $Y2=1.19
cc_406 VPB N_A_2668_793#_c_2405_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.605
+ $Y2=0.425
cc_407 VPB N_A_2668_793#_c_2402_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_408 VPB N_S[6]_c_2459_n 0.0238468f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_409 VPB N_S[14]_c_2510_n 0.01606f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_410 VPB N_S[14]_c_2508_n 0.00778682f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_411 VPB N_S[7]_c_2553_n 0.0238468f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_412 VPB N_S[15]_c_2603_n 0.01606f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_413 VPB N_S[15]_c_2599_n 0.00778682f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_414 VPB N_A_3017_47#_M1093_g 0.0216418f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_415 VPB N_A_3017_47#_c_2651_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_416 VPB N_A_3017_47#_c_2647_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_417 VPB N_A_3017_47#_c_2648_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_418 VPB N_A_3017_937#_M1038_g 0.0216418f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_419 VPB N_A_3017_937#_c_2708_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.645
+ $Y2=1.19
cc_420 VPB N_A_3017_937#_c_2704_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_421 VPB N_A_3017_937#_c_2705_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_422 VPB N_D[7]_c_2762_n 0.0294852f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_423 VPB N_D[7]_c_2765_n 0.00458905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_424 VPB N_D[15]_c_2794_n 0.0167392f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_425 VPB N_D[15]_c_2791_n 0.012746f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_426 VPB N_D[15]_c_2793_n 0.00458905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_427 VPB N_VPWR_c_2822_n 0.0424332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_428 VPB N_VPWR_c_2823_n 0.0424332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_429 VPB N_VPWR_c_2824_n 0.0150686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_430 VPB N_VPWR_c_2825_n 0.0150686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_431 VPB N_VPWR_c_2826_n 3.54074e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_432 VPB N_VPWR_c_2827_n 3.54074e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_433 VPB N_VPWR_c_2828_n 0.0150686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_434 VPB N_VPWR_c_2829_n 0.0150686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_435 VPB N_VPWR_c_2830_n 3.54074e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_436 VPB N_VPWR_c_2831_n 3.54074e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_437 VPB N_VPWR_c_2832_n 0.0150686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_438 VPB N_VPWR_c_2833_n 0.0150686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_439 VPB N_VPWR_c_2834_n 3.54074e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_440 VPB N_VPWR_c_2835_n 3.54074e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_441 VPB N_VPWR_c_2836_n 0.0150686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_442 VPB N_VPWR_c_2837_n 0.0150686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_443 VPB N_VPWR_c_2838_n 0.0424332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_444 VPB N_VPWR_c_2839_n 0.0424332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_445 VPB N_VPWR_c_2840_n 0.0154398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_446 VPB N_VPWR_c_2841_n 0.00207495f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_447 VPB N_VPWR_c_2842_n 0.0154398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_448 VPB N_VPWR_c_2843_n 0.00207495f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_449 VPB N_VPWR_c_2844_n 0.0154398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_450 VPB N_VPWR_c_2845_n 0.00207495f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_451 VPB N_VPWR_c_2846_n 0.0154398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_452 VPB N_VPWR_c_2847_n 0.00207495f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_453 VPB VPWR 0.10678f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_454 VPB N_VPWR_c_2849_n 0.0149679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_455 VPB N_VPWR_c_2850_n 0.0154398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_456 VPB N_VPWR_c_2851_n 0.0149679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_457 VPB N_VPWR_c_2852_n 0.0149679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_458 VPB N_VPWR_c_2853_n 0.0154398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_459 VPB N_VPWR_c_2854_n 0.0149679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_460 VPB N_VPWR_c_2855_n 0.0149679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_461 VPB N_VPWR_c_2856_n 0.0154398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_462 VPB N_VPWR_c_2857_n 0.0149679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_463 VPB N_VPWR_c_2858_n 0.0149679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_464 VPB N_VPWR_c_2859_n 0.0154398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_465 VPB N_VPWR_c_2860_n 0.0149679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_466 VPB N_VPWR_c_2861_n 0.00604875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_467 VPB N_VPWR_c_2862_n 0.00604875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_468 VPB N_Z_c_3315_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_469 VPB N_Z_c_3316_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_470 VPB N_Z_c_3365_n 0.00280567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_471 VPB N_Z_c_3366_n 0.00280567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_472 VPB N_Z_c_3367_n 0.00280567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_473 VPB N_Z_c_3368_n 0.00280567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_474 VPB N_Z_c_3323_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_475 VPB N_Z_c_3324_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_476 VPB N_Z_c_3325_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_477 VPB N_Z_c_3326_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_478 VPB N_Z_c_3373_n 0.00280567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_479 VPB N_Z_c_3374_n 0.00280567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_480 VPB N_Z_c_3375_n 0.00280567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_481 VPB N_Z_c_3376_n 0.00280567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_482 VPB N_Z_c_3333_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_483 VPB N_Z_c_3334_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_484 VPB N_Z_c_3335_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_485 VPB N_Z_c_3336_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_486 VPB N_Z_c_3381_n 0.00280567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_487 VPB N_Z_c_3382_n 0.00280567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_488 VPB N_Z_c_3383_n 0.00280567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_489 VPB N_Z_c_3384_n 0.00280567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_490 VPB N_Z_c_3343_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_491 VPB N_Z_c_3344_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_492 VPB N_Z_c_3345_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_493 VPB N_Z_c_3346_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_494 VPB N_Z_c_3389_n 0.00280567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_495 VPB N_Z_c_3390_n 0.00280567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_496 VPB N_Z_c_3391_n 0.00280567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_497 VPB N_Z_c_3392_n 0.00280567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_498 VPB N_Z_c_3353_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_499 VPB N_Z_c_3354_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_500 VPB N_Z_c_3395_n 0.00183099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_501 VPB N_Z_c_3396_n 0.00183099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_502 VPB N_Z_c_3397_n 0.00468622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_503 VPB N_Z_c_3398_n 0.00183099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_504 VPB N_Z_c_3399_n 0.00183099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_505 VPB N_Z_c_3400_n 0.00468622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_506 VPB N_Z_c_3401_n 0.00183099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_507 VPB N_Z_c_3402_n 0.00183099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_508 VPB N_Z_c_3403_n 0.00468622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_509 VPB N_Z_c_3404_n 0.00183099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_510 VPB N_Z_c_3405_n 0.00183099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_511 VPB N_Z_c_3406_n 0.00468622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_512 VPB N_Z_c_3407_n 0.00183099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_513 VPB N_Z_c_3408_n 0.00183099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_514 VPB N_Z_c_3409_n 0.00468622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_515 VPB N_Z_c_3410_n 0.00183099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_516 VPB N_Z_c_3411_n 0.00183099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_517 VPB N_Z_c_3412_n 0.00468622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_518 VPB N_Z_c_3413_n 0.00183099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_519 VPB N_Z_c_3414_n 0.00183099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_520 VPB N_Z_c_3415_n 0.00468622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_521 VPB N_Z_c_3416_n 0.00183099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_522 VPB N_Z_c_3417_n 0.00183099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_523 VPB N_Z_c_3418_n 0.00468622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_524 VPB N_Z_c_3419_n 0.00809084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_525 VPB N_Z_c_3420_n 0.00809084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_526 VPB N_Z_c_3421_n 0.00809084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_527 VPB N_Z_c_3422_n 0.00809084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_528 VPB N_Z_c_3423_n 0.00809084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_529 VPB N_Z_c_3424_n 0.00809084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_530 VPB N_Z_c_3425_n 0.00809084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_531 VPB N_Z_c_3426_n 0.00809084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_532 VPB N_Z_c_3427_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_533 VPB N_Z_c_3428_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_534 VPB N_Z_c_3429_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_535 VPB N_Z_c_3430_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_536 VPB N_Z_c_3431_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_537 VPB N_Z_c_3432_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_538 VPB N_Z_c_3433_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_539 VPB N_Z_c_3434_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_540 VPB N_Z_c_3435_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_541 VPB N_Z_c_3436_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_542 VPB N_Z_c_3437_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_543 VPB N_Z_c_3438_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_544 VPB N_Z_c_3439_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_545 VPB N_Z_c_3440_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_546 VPB N_Z_c_3441_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_547 VPB N_Z_c_3442_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_548 N_D[0]_c_549_n N_D[8]_c_581_n 0.0129371f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_549 N_D[0]_c_549_n N_A_184_265#_M1036_g 0.0383393f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_550 N_D[0]_c_549_n N_A_184_265#_c_611_n 0.00712672f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_551 N_D[0]_c_548_n N_S[0]_c_722_n 0.0286599f $X=0.47 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_552 N_D[0]_c_550_n N_S[0]_c_722_n 0.00289497f $X=0.645 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_553 N_D[0]_c_549_n N_VPWR_c_2822_n 0.0235f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_554 N_D[0]_c_551_n N_VPWR_c_2822_n 0.00471543f $X=0.645 $Y=1.19 $X2=0 $Y2=0
cc_555 N_D[0]_c_549_n VPWR 0.00937833f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_556 N_D[0]_c_549_n N_VPWR_c_2849_n 0.00342413f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_557 N_D[0]_c_549_n N_Z_c_3315_n 0.00605747f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_558 N_D[0]_c_550_n N_Z_c_3315_n 0.00376465f $X=0.645 $Y=1.055 $X2=0 $Y2=0
cc_559 N_D[0]_c_551_n N_Z_c_3315_n 0.0216525f $X=0.645 $Y=1.19 $X2=0 $Y2=0
cc_560 N_D[0]_c_550_n N_Z_c_3317_n 0.0128881f $X=0.645 $Y=1.055 $X2=0 $Y2=0
cc_561 N_D[0]_c_550_n N_Z_c_3318_n 0.00686805f $X=0.645 $Y=1.055 $X2=0 $Y2=0
cc_562 N_D[0]_c_549_n N_Z_c_3365_n 0.00176496f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_563 N_D[0]_c_548_n N_VGND_c_4368_n 0.00487865f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_564 N_D[0]_c_551_n N_VGND_c_4368_n 0.00222881f $X=0.645 $Y=1.19 $X2=0 $Y2=0
cc_565 N_D[0]_c_548_n N_VGND_c_4389_n 0.00585385f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_566 D[0] N_VGND_c_4389_n 0.00842546f $X=0.605 $Y=0.425 $X2=0 $Y2=0
cc_567 N_D[0]_c_548_n VGND 0.011617f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_568 D[0] VGND 0.00942277f $X=0.605 $Y=0.425 $X2=0 $Y2=0
cc_569 N_D[0]_c_550_n A_109_47# 0.00426617f $X=0.645 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_570 D[0] A_109_47# 0.00894235f $X=0.605 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_571 N_D[8]_c_581_n N_A_184_793#_M1090_g 0.0383393f $X=0.495 $Y=4.03 $X2=0
+ $Y2=0
cc_572 N_D[8]_c_577_n N_A_184_793#_c_668_n 0.00496096f $X=0.47 $Y=4.445 $X2=0
+ $Y2=0
cc_573 N_D[8]_c_581_n N_A_184_793#_c_668_n 0.00216577f $X=0.495 $Y=4.03 $X2=0
+ $Y2=0
cc_574 N_D[8]_c_577_n N_S[8]_c_773_n 0.0286599f $X=0.47 $Y=4.445 $X2=0 $Y2=0
cc_575 N_D[8]_c_578_n N_S[8]_c_773_n 0.00289497f $X=0.645 $Y=4.815 $X2=0 $Y2=0
cc_576 N_D[8]_c_581_n N_VPWR_c_2823_n 0.0235f $X=0.495 $Y=4.03 $X2=0 $Y2=0
cc_577 N_D[8]_c_579_n N_VPWR_c_2823_n 0.00471543f $X=0.645 $Y=4.25 $X2=0 $Y2=0
cc_578 N_D[8]_c_581_n VPWR 0.00937833f $X=0.495 $Y=4.03 $X2=0 $Y2=0
cc_579 N_D[8]_c_581_n N_VPWR_c_2849_n 0.00342413f $X=0.495 $Y=4.03 $X2=0 $Y2=0
cc_580 N_D[8]_c_577_n N_Z_c_3316_n 0.00299906f $X=0.47 $Y=4.445 $X2=0 $Y2=0
cc_581 N_D[8]_c_581_n N_Z_c_3316_n 0.00305841f $X=0.495 $Y=4.03 $X2=0 $Y2=0
cc_582 N_D[8]_c_578_n N_Z_c_3316_n 0.00376465f $X=0.645 $Y=4.815 $X2=0 $Y2=0
cc_583 N_D[8]_c_579_n N_Z_c_3316_n 0.0216525f $X=0.645 $Y=4.25 $X2=0 $Y2=0
cc_584 N_D[8]_c_578_n N_Z_c_3319_n 0.0128881f $X=0.645 $Y=4.815 $X2=0 $Y2=0
cc_585 N_D[8]_c_578_n N_Z_c_3320_n 0.00686805f $X=0.645 $Y=4.815 $X2=0 $Y2=0
cc_586 N_D[8]_c_581_n N_Z_c_3397_n 0.00176496f $X=0.495 $Y=4.03 $X2=0 $Y2=0
cc_587 N_D[8]_c_577_n N_VGND_c_4370_n 0.00487865f $X=0.47 $Y=4.445 $X2=0 $Y2=0
cc_588 N_D[8]_c_579_n N_VGND_c_4370_n 0.00222881f $X=0.645 $Y=4.25 $X2=0 $Y2=0
cc_589 N_D[8]_c_577_n N_VGND_c_4391_n 0.00585385f $X=0.47 $Y=4.445 $X2=0 $Y2=0
cc_590 D[8] N_VGND_c_4391_n 0.00842546f $X=0.605 $Y=4.845 $X2=0 $Y2=0
cc_591 N_D[8]_c_577_n VGND 0.011617f $X=0.47 $Y=4.445 $X2=0 $Y2=0
cc_592 D[8] VGND 0.00941728f $X=0.605 $Y=4.845 $X2=0 $Y2=0
cc_593 N_D[8]_c_578_n A_109_911# 0.00426617f $X=0.645 $Y=4.815 $X2=-0.19
+ $Y2=-0.24
cc_594 D[8] A_109_911# 0.00894235f $X=0.605 $Y=4.845 $X2=-0.19 $Y2=-0.24
cc_595 N_A_184_265#_M1036_g N_A_184_793#_M1090_g 0.0129371f $X=1.02 $Y=2.075
+ $X2=0 $Y2=0
cc_596 N_A_184_265#_c_608_n N_S[0]_c_723_n 0.00827389f $X=1.545 $Y=0.755 $X2=0
+ $Y2=0
cc_597 N_A_184_265#_c_609_n N_S[0]_c_723_n 0.0164662f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_598 N_A_184_265#_c_610_n N_S[0]_c_723_n 0.00928634f $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_599 N_A_184_265#_c_611_n N_S[0]_c_723_n 0.0184911f $X=1.02 $Y=1.34 $X2=0
+ $Y2=0
cc_600 N_A_184_265#_c_611_n N_S[0]_c_724_n 0.00820745f $X=1.02 $Y=1.34 $X2=0
+ $Y2=0
cc_601 N_A_184_265#_c_609_n N_S[0]_c_725_n 0.0012443f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_602 N_A_184_265#_c_613_n N_S[0]_c_725_n 0.00902681f $X=1.775 $Y=2.31 $X2=0
+ $Y2=0
cc_603 N_A_184_265#_c_610_n N_S[0]_c_725_n 0.00767015f $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_604 N_A_184_265#_c_611_n N_S[0]_c_725_n 0.00659591f $X=1.02 $Y=1.34 $X2=0
+ $Y2=0
cc_605 N_A_184_265#_c_609_n N_S[0]_c_726_n 0.00219336f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_606 N_A_184_265#_c_608_n N_S[0]_c_727_n 0.00603567f $X=1.545 $Y=0.755 $X2=0
+ $Y2=0
cc_607 N_A_184_265#_c_609_n N_S[0]_c_727_n 0.0178233f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_608 N_A_184_265#_c_610_n N_S[0]_c_727_n 0.0214702f $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_609 N_A_184_265#_c_611_n N_S[0]_c_727_n 2.59957e-19 $X=1.02 $Y=1.34 $X2=0
+ $Y2=0
cc_610 N_A_184_265#_M1036_g N_VPWR_c_2822_n 0.00247893f $X=1.02 $Y=2.075 $X2=0
+ $Y2=0
cc_611 N_A_184_265#_c_613_n N_VPWR_c_2824_n 0.0292866f $X=1.775 $Y=2.31 $X2=0
+ $Y2=0
cc_612 N_A_184_265#_c_610_n N_VPWR_c_2824_n 0.00688579f $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_613 N_A_184_265#_c_613_n N_VPWR_c_2840_n 0.0210596f $X=1.775 $Y=2.31 $X2=0
+ $Y2=0
cc_614 N_A_184_265#_M1045_s VPWR 0.00179197f $X=1.65 $Y=1.485 $X2=0 $Y2=0
cc_615 N_A_184_265#_M1036_g VPWR 0.00407291f $X=1.02 $Y=2.075 $X2=0 $Y2=0
cc_616 N_A_184_265#_c_613_n VPWR 0.00594162f $X=1.775 $Y=2.31 $X2=0 $Y2=0
cc_617 N_A_184_265#_M1036_g N_Z_c_3315_n 0.00862328f $X=1.02 $Y=2.075 $X2=0
+ $Y2=0
cc_618 N_A_184_265#_c_609_n N_Z_c_3315_n 0.00719188f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_619 N_A_184_265#_c_613_n N_Z_c_3315_n 0.00378484f $X=1.775 $Y=2.31 $X2=0
+ $Y2=0
cc_620 N_A_184_265#_c_610_n N_Z_c_3315_n 0.0304368f $X=1.775 $Y=1.63 $X2=0 $Y2=0
cc_621 N_A_184_265#_c_611_n N_Z_c_3315_n 0.00814206f $X=1.02 $Y=1.34 $X2=0 $Y2=0
cc_622 N_A_184_265#_c_609_n N_Z_c_3317_n 0.0124144f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_623 N_A_184_265#_c_610_n N_Z_c_3317_n 0.00398133f $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_624 N_A_184_265#_c_611_n N_Z_c_3317_n 0.00349316f $X=1.02 $Y=1.34 $X2=0 $Y2=0
cc_625 N_A_184_265#_c_608_n N_Z_c_3318_n 0.0259454f $X=1.545 $Y=0.755 $X2=0
+ $Y2=0
cc_626 N_A_184_265#_c_609_n N_Z_c_3318_n 0.00611965f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_627 N_A_184_265#_M1036_g N_Z_c_3365_n 0.00544362f $X=1.02 $Y=2.075 $X2=0
+ $Y2=0
cc_628 N_A_184_265#_c_613_n N_Z_c_3365_n 0.0371028f $X=1.775 $Y=2.31 $X2=0 $Y2=0
cc_629 N_A_184_265#_M1036_g N_Z_c_3395_n 0.00335035f $X=1.02 $Y=2.075 $X2=0
+ $Y2=0
cc_630 N_A_184_265#_M1036_g N_Z_c_3397_n 0.00502861f $X=1.02 $Y=2.075 $X2=0
+ $Y2=0
cc_631 N_A_184_265#_c_613_n N_Z_c_3419_n 0.0291787f $X=1.775 $Y=2.31 $X2=0 $Y2=0
cc_632 N_A_184_265#_c_610_n N_Z_c_3419_n 0.0126642f $X=1.775 $Y=1.63 $X2=0 $Y2=0
cc_633 N_A_184_265#_M1036_g N_Z_c_3472_n 0.00289142f $X=1.02 $Y=2.075 $X2=0
+ $Y2=0
cc_634 N_A_184_265#_c_613_n N_Z_c_3472_n 6.03258e-19 $X=1.775 $Y=2.31 $X2=0
+ $Y2=0
cc_635 N_A_184_265#_c_610_n N_Z_c_3472_n 4.25753e-19 $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_636 N_A_184_265#_M1036_g N_Z_c_3427_n 0.0107335f $X=1.02 $Y=2.075 $X2=0 $Y2=0
cc_637 N_A_184_265#_c_613_n N_Z_c_3427_n 0.0139746f $X=1.775 $Y=2.31 $X2=0 $Y2=0
cc_638 N_A_184_265#_c_610_n N_Z_c_3427_n 0.00749574f $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_639 N_A_184_265#_c_611_n N_Z_c_3427_n 0.00449418f $X=1.02 $Y=1.34 $X2=0 $Y2=0
cc_640 N_A_184_265#_c_608_n N_VGND_c_4389_n 0.015238f $X=1.545 $Y=0.755 $X2=0
+ $Y2=0
cc_641 N_A_184_265#_M1058_s VGND 0.00358139f $X=1.65 $Y=0.235 $X2=0 $Y2=0
cc_642 N_A_184_265#_c_608_n VGND 0.0150148f $X=1.545 $Y=0.755 $X2=0 $Y2=0
cc_643 N_A_184_793#_c_666_n N_S[8]_c_772_n 0.0247401f $X=1.545 $Y=4.685 $X2=0
+ $Y2=0
cc_644 N_A_184_793#_c_667_n N_S[8]_c_772_n 0.00928634f $X=1.775 $Y=3.805 $X2=0
+ $Y2=0
cc_645 N_A_184_793#_c_668_n N_S[8]_c_772_n 0.0184911f $X=1.02 $Y=4.1 $X2=0 $Y2=0
cc_646 N_A_184_793#_c_668_n N_S[8]_c_773_n 0.00820745f $X=1.02 $Y=4.1 $X2=0
+ $Y2=0
cc_647 N_A_184_793#_c_667_n N_S[8]_c_776_n 0.00382813f $X=1.775 $Y=3.805 $X2=0
+ $Y2=0
cc_648 N_A_184_793#_c_671_n N_S[8]_c_776_n 0.00902681f $X=1.775 $Y=3.13 $X2=0
+ $Y2=0
cc_649 N_A_184_793#_c_668_n N_S[8]_c_776_n 0.00150889f $X=1.02 $Y=4.1 $X2=0
+ $Y2=0
cc_650 N_A_184_793#_c_666_n N_S[8]_c_774_n 0.00343766f $X=1.545 $Y=4.685 $X2=0
+ $Y2=0
cc_651 N_A_184_793#_c_667_n N_S[8]_c_774_n 0.00384202f $X=1.775 $Y=3.805 $X2=0
+ $Y2=0
cc_652 N_A_184_793#_c_668_n N_S[8]_c_774_n 0.00508702f $X=1.02 $Y=4.1 $X2=0
+ $Y2=0
cc_653 N_A_184_793#_c_666_n S[8] 0.023859f $X=1.545 $Y=4.685 $X2=0 $Y2=0
cc_654 N_A_184_793#_c_667_n S[8] 0.0214702f $X=1.775 $Y=3.805 $X2=0 $Y2=0
cc_655 N_A_184_793#_c_668_n S[8] 2.59957e-19 $X=1.02 $Y=4.1 $X2=0 $Y2=0
cc_656 N_A_184_793#_M1090_g N_VPWR_c_2823_n 0.00247893f $X=1.02 $Y=3.365 $X2=0
+ $Y2=0
cc_657 N_A_184_793#_c_667_n N_VPWR_c_2825_n 0.00688579f $X=1.775 $Y=3.805 $X2=0
+ $Y2=0
cc_658 N_A_184_793#_c_671_n N_VPWR_c_2825_n 0.0292866f $X=1.775 $Y=3.13 $X2=0
+ $Y2=0
cc_659 N_A_184_793#_c_671_n N_VPWR_c_2840_n 0.0210596f $X=1.775 $Y=3.13 $X2=0
+ $Y2=0
cc_660 N_A_184_793#_M1048_s VPWR 0.00179197f $X=1.65 $Y=2.955 $X2=0 $Y2=0
cc_661 N_A_184_793#_M1090_g VPWR 0.00407291f $X=1.02 $Y=3.365 $X2=0 $Y2=0
cc_662 N_A_184_793#_c_671_n VPWR 0.00594162f $X=1.775 $Y=3.13 $X2=0 $Y2=0
cc_663 N_A_184_793#_M1090_g N_Z_c_3316_n 0.00862328f $X=1.02 $Y=3.365 $X2=0
+ $Y2=0
cc_664 N_A_184_793#_c_666_n N_Z_c_3316_n 0.00719188f $X=1.545 $Y=4.685 $X2=0
+ $Y2=0
cc_665 N_A_184_793#_c_667_n N_Z_c_3316_n 0.0304368f $X=1.775 $Y=3.805 $X2=0
+ $Y2=0
cc_666 N_A_184_793#_c_671_n N_Z_c_3316_n 0.00378484f $X=1.775 $Y=3.13 $X2=0
+ $Y2=0
cc_667 N_A_184_793#_c_668_n N_Z_c_3316_n 0.00814206f $X=1.02 $Y=4.1 $X2=0 $Y2=0
cc_668 N_A_184_793#_c_666_n N_Z_c_3319_n 0.0124144f $X=1.545 $Y=4.685 $X2=0
+ $Y2=0
cc_669 N_A_184_793#_c_667_n N_Z_c_3319_n 0.00398133f $X=1.775 $Y=3.805 $X2=0
+ $Y2=0
cc_670 N_A_184_793#_c_668_n N_Z_c_3319_n 0.00349316f $X=1.02 $Y=4.1 $X2=0 $Y2=0
cc_671 N_A_184_793#_c_666_n N_Z_c_3320_n 0.032065f $X=1.545 $Y=4.685 $X2=0 $Y2=0
cc_672 N_A_184_793#_M1090_g N_Z_c_3366_n 0.00544362f $X=1.02 $Y=3.365 $X2=0
+ $Y2=0
cc_673 N_A_184_793#_M1090_g N_Z_c_3396_n 0.00335035f $X=1.02 $Y=3.365 $X2=0
+ $Y2=0
cc_674 N_A_184_793#_c_671_n N_Z_c_3396_n 0.0371028f $X=1.775 $Y=3.13 $X2=0 $Y2=0
cc_675 N_A_184_793#_M1090_g N_Z_c_3397_n 0.00502861f $X=1.02 $Y=3.365 $X2=0
+ $Y2=0
cc_676 N_A_184_793#_c_667_n N_Z_c_3420_n 0.0126642f $X=1.775 $Y=3.805 $X2=0
+ $Y2=0
cc_677 N_A_184_793#_c_671_n N_Z_c_3420_n 0.0291787f $X=1.775 $Y=3.13 $X2=0 $Y2=0
cc_678 N_A_184_793#_M1090_g N_Z_c_3494_n 0.00289142f $X=1.02 $Y=3.365 $X2=0
+ $Y2=0
cc_679 N_A_184_793#_c_667_n N_Z_c_3494_n 4.25753e-19 $X=1.775 $Y=3.805 $X2=0
+ $Y2=0
cc_680 N_A_184_793#_c_671_n N_Z_c_3494_n 6.03258e-19 $X=1.775 $Y=3.13 $X2=0
+ $Y2=0
cc_681 N_A_184_793#_M1090_g N_Z_c_3428_n 0.0107344f $X=1.02 $Y=3.365 $X2=0 $Y2=0
cc_682 N_A_184_793#_c_667_n N_Z_c_3428_n 0.00749574f $X=1.775 $Y=3.805 $X2=0
+ $Y2=0
cc_683 N_A_184_793#_c_671_n N_Z_c_3428_n 0.0139746f $X=1.775 $Y=3.13 $X2=0 $Y2=0
cc_684 N_A_184_793#_c_668_n N_Z_c_3428_n 0.00449418f $X=1.02 $Y=4.1 $X2=0 $Y2=0
cc_685 N_A_184_793#_c_666_n N_VGND_c_4391_n 0.015238f $X=1.545 $Y=4.685 $X2=0
+ $Y2=0
cc_686 N_A_184_793#_M1067_s VGND 0.00358139f $X=1.65 $Y=4.685 $X2=0 $Y2=0
cc_687 N_A_184_793#_c_666_n VGND 0.0150148f $X=1.545 $Y=4.685 $X2=0 $Y2=0
cc_688 N_S[0]_c_725_n N_S[8]_c_776_n 0.0130744f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_689 N_S[0]_c_725_n N_S[1]_c_819_n 0.0578733f $X=2.01 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_690 N_S[0]_c_727_n N_S[1]_c_819_n 0.00112057f $X=1.975 $Y=1.03 $X2=-0.19
+ $Y2=-0.24
cc_691 N_S[0]_c_726_n N_S[1]_c_820_n 0.0091402f $X=2.01 $Y=0.83 $X2=0 $Y2=0
cc_692 N_S[0]_c_725_n N_S[1]_c_823_n 0.00112057f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_693 N_S[0]_c_727_n N_S[1]_c_823_n 0.0277403f $X=1.975 $Y=1.03 $X2=0 $Y2=0
cc_694 N_S[0]_c_725_n N_VPWR_c_2824_n 0.00965725f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_695 N_S[0]_c_727_n N_VPWR_c_2824_n 0.00587376f $X=1.975 $Y=1.03 $X2=0 $Y2=0
cc_696 N_S[0]_c_725_n N_VPWR_c_2840_n 0.0035837f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_697 N_S[0]_c_725_n VPWR 0.0072999f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_698 N_S[0]_c_724_n N_Z_c_3315_n 7.46972e-19 $X=1.02 $Y=0.905 $X2=0 $Y2=0
cc_699 N_S[0]_c_723_n N_Z_c_3317_n 0.00806549f $X=1.84 $Y=0.905 $X2=0 $Y2=0
cc_700 N_S[0]_c_724_n N_Z_c_3317_n 0.00605736f $X=1.02 $Y=0.905 $X2=0 $Y2=0
cc_701 N_S[0]_c_722_n N_Z_c_3318_n 0.00316445f $X=0.945 $Y=0.83 $X2=0 $Y2=0
cc_702 N_S[0]_c_723_n N_Z_c_3318_n 0.00501353f $X=1.84 $Y=0.905 $X2=0 $Y2=0
cc_703 N_S[0]_c_725_n N_Z_c_3397_n 0.00124373f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_704 N_S[0]_c_725_n N_Z_c_3419_n 0.0062071f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_705 N_S[0]_c_727_n N_Z_c_3419_n 0.00659242f $X=1.975 $Y=1.03 $X2=0 $Y2=0
cc_706 N_S[0]_c_726_n N_VGND_c_4371_n 0.00570474f $X=2.01 $Y=0.83 $X2=0 $Y2=0
cc_707 N_S[0]_c_727_n N_VGND_c_4371_n 0.00391126f $X=1.975 $Y=1.03 $X2=0 $Y2=0
cc_708 N_S[0]_c_722_n N_VGND_c_4389_n 0.00585385f $X=0.945 $Y=0.83 $X2=0 $Y2=0
cc_709 N_S[0]_c_726_n N_VGND_c_4389_n 0.00585385f $X=2.01 $Y=0.83 $X2=0 $Y2=0
cc_710 N_S[0]_c_722_n VGND 0.00880034f $X=0.945 $Y=0.83 $X2=0 $Y2=0
cc_711 N_S[0]_c_723_n VGND 0.00349917f $X=1.84 $Y=0.905 $X2=0 $Y2=0
cc_712 N_S[0]_c_725_n VGND 6.15795e-19 $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_713 N_S[0]_c_726_n VGND 0.0124506f $X=2.01 $Y=0.83 $X2=0 $Y2=0
cc_714 N_S[8]_c_776_n N_S[9]_c_869_n 0.0296874f $X=2.01 $Y=4.03 $X2=-0.19
+ $Y2=-0.24
cc_715 N_S[8]_c_774_n N_S[9]_c_865_n 0.0373261f $X=2.01 $Y=4.61 $X2=0 $Y2=0
cc_716 S[8] N_S[9]_c_865_n 0.00112057f $X=1.985 $Y=4.165 $X2=0 $Y2=0
cc_717 N_S[8]_c_774_n S[9] 0.00112057f $X=2.01 $Y=4.61 $X2=0 $Y2=0
cc_718 S[8] S[9] 0.0277403f $X=1.985 $Y=4.165 $X2=0 $Y2=0
cc_719 N_S[8]_c_776_n N_VPWR_c_2825_n 0.00965725f $X=2.01 $Y=4.03 $X2=0 $Y2=0
cc_720 S[8] N_VPWR_c_2825_n 0.00587376f $X=1.985 $Y=4.165 $X2=0 $Y2=0
cc_721 N_S[8]_c_776_n N_VPWR_c_2840_n 0.0035837f $X=2.01 $Y=4.03 $X2=0 $Y2=0
cc_722 N_S[8]_c_776_n VPWR 0.0072999f $X=2.01 $Y=4.03 $X2=0 $Y2=0
cc_723 N_S[8]_c_773_n N_Z_c_3316_n 7.46972e-19 $X=1.02 $Y=4.535 $X2=0 $Y2=0
cc_724 N_S[8]_c_772_n N_Z_c_3319_n 0.00806549f $X=1.84 $Y=4.535 $X2=0 $Y2=0
cc_725 N_S[8]_c_773_n N_Z_c_3319_n 0.00605736f $X=1.02 $Y=4.535 $X2=0 $Y2=0
cc_726 N_S[8]_c_771_n N_Z_c_3320_n 0.00316445f $X=0.945 $Y=4.61 $X2=0 $Y2=0
cc_727 N_S[8]_c_772_n N_Z_c_3320_n 0.00501353f $X=1.84 $Y=4.535 $X2=0 $Y2=0
cc_728 N_S[8]_c_776_n N_Z_c_3397_n 0.00124373f $X=2.01 $Y=4.03 $X2=0 $Y2=0
cc_729 N_S[8]_c_776_n N_Z_c_3420_n 0.00597491f $X=2.01 $Y=4.03 $X2=0 $Y2=0
cc_730 N_S[8]_c_774_n N_Z_c_3420_n 2.32192e-19 $X=2.01 $Y=4.61 $X2=0 $Y2=0
cc_731 S[8] N_Z_c_3420_n 0.00659242f $X=1.985 $Y=4.165 $X2=0 $Y2=0
cc_732 N_S[8]_c_774_n N_VGND_c_4372_n 0.00570474f $X=2.01 $Y=4.61 $X2=0 $Y2=0
cc_733 S[8] N_VGND_c_4372_n 0.00391126f $X=1.985 $Y=4.165 $X2=0 $Y2=0
cc_734 N_S[8]_c_771_n N_VGND_c_4391_n 0.00585385f $X=0.945 $Y=4.61 $X2=0 $Y2=0
cc_735 N_S[8]_c_774_n N_VGND_c_4391_n 0.00585385f $X=2.01 $Y=4.61 $X2=0 $Y2=0
cc_736 N_S[8]_c_771_n VGND 0.00880034f $X=0.945 $Y=4.61 $X2=0 $Y2=0
cc_737 N_S[8]_c_772_n VGND 0.00349917f $X=1.84 $Y=4.535 $X2=0 $Y2=0
cc_738 N_S[8]_c_774_n VGND 0.0130664f $X=2.01 $Y=4.61 $X2=0 $Y2=0
cc_739 N_S[1]_c_819_n N_S[9]_c_869_n 0.0130744f $X=2.59 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_740 N_S[1]_c_819_n N_A_533_47#_c_917_n 0.00902681f $X=2.59 $Y=1.41 $X2=0
+ $Y2=0
cc_741 N_S[1]_c_819_n N_A_533_47#_c_912_n 0.0012443f $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_742 N_S[1]_c_820_n N_A_533_47#_c_912_n 0.00219336f $X=2.59 $Y=0.83 $X2=0
+ $Y2=0
cc_743 N_S[1]_c_821_n N_A_533_47#_c_912_n 0.0164662f $X=3.58 $Y=0.905 $X2=0
+ $Y2=0
cc_744 N_S[1]_c_823_n N_A_533_47#_c_912_n 0.0178233f $X=2.625 $Y=1.03 $X2=0
+ $Y2=0
cc_745 N_S[1]_c_819_n N_A_533_47#_c_913_n 0.00767015f $X=2.59 $Y=1.41 $X2=0
+ $Y2=0
cc_746 N_S[1]_c_821_n N_A_533_47#_c_913_n 0.00928634f $X=3.58 $Y=0.905 $X2=0
+ $Y2=0
cc_747 N_S[1]_c_823_n N_A_533_47#_c_913_n 0.0214702f $X=2.625 $Y=1.03 $X2=0
+ $Y2=0
cc_748 N_S[1]_c_819_n N_A_533_47#_c_914_n 0.00659591f $X=2.59 $Y=1.41 $X2=0
+ $Y2=0
cc_749 N_S[1]_c_821_n N_A_533_47#_c_914_n 0.0266986f $X=3.58 $Y=0.905 $X2=0
+ $Y2=0
cc_750 N_S[1]_c_823_n N_A_533_47#_c_914_n 2.59957e-19 $X=2.625 $Y=1.03 $X2=0
+ $Y2=0
cc_751 N_S[1]_c_819_n N_A_533_47#_c_915_n 0.00827389f $X=2.59 $Y=1.41 $X2=0
+ $Y2=0
cc_752 N_S[1]_c_823_n N_A_533_47#_c_915_n 0.00603567f $X=2.625 $Y=1.03 $X2=0
+ $Y2=0
cc_753 N_S[1]_c_822_n N_D[1]_c_1029_n 0.0286599f $X=3.655 $Y=0.83 $X2=0 $Y2=0
cc_754 N_S[1]_c_822_n N_D[1]_c_1030_n 0.00289497f $X=3.655 $Y=0.83 $X2=0 $Y2=0
cc_755 N_S[1]_c_819_n N_VPWR_c_2824_n 0.00965725f $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_756 N_S[1]_c_823_n N_VPWR_c_2824_n 0.00587376f $X=2.625 $Y=1.03 $X2=0 $Y2=0
cc_757 N_S[1]_c_819_n VPWR 0.0072999f $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_758 N_S[1]_c_819_n N_VPWR_c_2850_n 0.0035837f $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_759 N_S[1]_c_821_n N_Z_c_3321_n 0.00501353f $X=3.58 $Y=0.905 $X2=0 $Y2=0
cc_760 N_S[1]_c_822_n N_Z_c_3321_n 0.00316445f $X=3.655 $Y=0.83 $X2=0 $Y2=0
cc_761 N_S[1]_c_821_n N_Z_c_3323_n 7.46972e-19 $X=3.58 $Y=0.905 $X2=0 $Y2=0
cc_762 N_S[1]_c_819_n N_Z_c_3400_n 0.00124373f $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_763 N_S[1]_c_821_n N_Z_c_3355_n 0.0141229f $X=3.58 $Y=0.905 $X2=0 $Y2=0
cc_764 N_S[1]_c_819_n N_Z_c_3419_n 0.0062071f $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_765 N_S[1]_c_823_n N_Z_c_3419_n 0.00659242f $X=2.625 $Y=1.03 $X2=0 $Y2=0
cc_766 N_S[1]_c_820_n N_VGND_c_4371_n 0.00570474f $X=2.59 $Y=0.83 $X2=0 $Y2=0
cc_767 N_S[1]_c_823_n N_VGND_c_4371_n 0.00391126f $X=2.625 $Y=1.03 $X2=0 $Y2=0
cc_768 N_S[1]_c_819_n VGND 6.15795e-19 $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_769 N_S[1]_c_820_n VGND 0.0124506f $X=2.59 $Y=0.83 $X2=0 $Y2=0
cc_770 N_S[1]_c_821_n VGND 0.00349917f $X=3.58 $Y=0.905 $X2=0 $Y2=0
cc_771 N_S[1]_c_822_n VGND 0.00880034f $X=3.655 $Y=0.83 $X2=0 $Y2=0
cc_772 N_S[1]_c_820_n N_VGND_c_4407_n 0.00585385f $X=2.59 $Y=0.83 $X2=0 $Y2=0
cc_773 N_S[1]_c_822_n N_VGND_c_4407_n 0.00585385f $X=3.655 $Y=0.83 $X2=0 $Y2=0
cc_774 N_S[9]_c_869_n N_A_533_937#_c_974_n 0.00902681f $X=2.59 $Y=4.03 $X2=0
+ $Y2=0
cc_775 N_S[9]_c_865_n N_A_533_937#_c_969_n 0.00343766f $X=2.59 $Y=4.61 $X2=0
+ $Y2=0
cc_776 N_S[9]_c_866_n N_A_533_937#_c_969_n 0.0164662f $X=3.58 $Y=4.535 $X2=0
+ $Y2=0
cc_777 S[9] N_A_533_937#_c_969_n 0.0178233f $X=2.445 $Y=4.165 $X2=0 $Y2=0
cc_778 N_S[9]_c_869_n N_A_533_937#_c_970_n 0.00382813f $X=2.59 $Y=4.03 $X2=0
+ $Y2=0
cc_779 N_S[9]_c_865_n N_A_533_937#_c_970_n 0.00384202f $X=2.59 $Y=4.61 $X2=0
+ $Y2=0
cc_780 N_S[9]_c_866_n N_A_533_937#_c_970_n 0.00928634f $X=3.58 $Y=4.535 $X2=0
+ $Y2=0
cc_781 S[9] N_A_533_937#_c_970_n 0.0214702f $X=2.445 $Y=4.165 $X2=0 $Y2=0
cc_782 N_S[9]_c_869_n N_A_533_937#_c_971_n 0.00150889f $X=2.59 $Y=4.03 $X2=0
+ $Y2=0
cc_783 N_S[9]_c_865_n N_A_533_937#_c_971_n 0.00508702f $X=2.59 $Y=4.61 $X2=0
+ $Y2=0
cc_784 N_S[9]_c_866_n N_A_533_937#_c_971_n 0.0266986f $X=3.58 $Y=4.535 $X2=0
+ $Y2=0
cc_785 S[9] N_A_533_937#_c_971_n 2.59957e-19 $X=2.445 $Y=4.165 $X2=0 $Y2=0
cc_786 N_S[9]_c_865_n N_A_533_937#_c_972_n 0.00827389f $X=2.59 $Y=4.61 $X2=0
+ $Y2=0
cc_787 S[9] N_A_533_937#_c_972_n 0.00603567f $X=2.445 $Y=4.165 $X2=0 $Y2=0
cc_788 N_S[9]_c_866_n N_D[9]_c_1066_n 0.0286599f $X=3.58 $Y=4.535 $X2=0 $Y2=0
cc_789 N_S[9]_c_866_n N_D[9]_c_1067_n 0.00289497f $X=3.58 $Y=4.535 $X2=0 $Y2=0
cc_790 N_S[9]_c_869_n N_VPWR_c_2825_n 0.00965725f $X=2.59 $Y=4.03 $X2=0 $Y2=0
cc_791 S[9] N_VPWR_c_2825_n 0.00587376f $X=2.445 $Y=4.165 $X2=0 $Y2=0
cc_792 N_S[9]_c_869_n VPWR 0.0072999f $X=2.59 $Y=4.03 $X2=0 $Y2=0
cc_793 N_S[9]_c_869_n N_VPWR_c_2850_n 0.0035837f $X=2.59 $Y=4.03 $X2=0 $Y2=0
cc_794 N_S[9]_c_866_n N_Z_c_3322_n 0.00501353f $X=3.58 $Y=4.535 $X2=0 $Y2=0
cc_795 N_S[9]_c_867_n N_Z_c_3322_n 0.00316445f $X=3.655 $Y=4.61 $X2=0 $Y2=0
cc_796 N_S[9]_c_866_n N_Z_c_3324_n 7.46972e-19 $X=3.58 $Y=4.535 $X2=0 $Y2=0
cc_797 N_S[9]_c_869_n N_Z_c_3400_n 0.00124373f $X=2.59 $Y=4.03 $X2=0 $Y2=0
cc_798 N_S[9]_c_866_n N_Z_c_3356_n 0.0141229f $X=3.58 $Y=4.535 $X2=0 $Y2=0
cc_799 N_S[9]_c_869_n N_Z_c_3420_n 0.00597491f $X=2.59 $Y=4.03 $X2=0 $Y2=0
cc_800 N_S[9]_c_865_n N_Z_c_3420_n 2.32192e-19 $X=2.59 $Y=4.61 $X2=0 $Y2=0
cc_801 S[9] N_Z_c_3420_n 0.00659242f $X=2.445 $Y=4.165 $X2=0 $Y2=0
cc_802 N_S[9]_c_865_n N_VGND_c_4372_n 0.00570474f $X=2.59 $Y=4.61 $X2=0 $Y2=0
cc_803 S[9] N_VGND_c_4372_n 0.00391126f $X=2.445 $Y=4.165 $X2=0 $Y2=0
cc_804 N_S[9]_c_865_n VGND 0.0130664f $X=2.59 $Y=4.61 $X2=0 $Y2=0
cc_805 N_S[9]_c_866_n VGND 0.00349917f $X=3.58 $Y=4.535 $X2=0 $Y2=0
cc_806 N_S[9]_c_867_n VGND 0.00880034f $X=3.655 $Y=4.61 $X2=0 $Y2=0
cc_807 N_S[9]_c_865_n N_VGND_c_4408_n 0.00585385f $X=2.59 $Y=4.61 $X2=0 $Y2=0
cc_808 N_S[9]_c_867_n N_VGND_c_4408_n 0.00585385f $X=3.655 $Y=4.61 $X2=0 $Y2=0
cc_809 N_A_533_47#_M1017_g N_A_533_937#_M1071_g 0.0129371f $X=3.58 $Y=2.075
+ $X2=0 $Y2=0
cc_810 N_A_533_47#_M1017_g N_D[1]_c_1028_n 0.0390641f $X=3.58 $Y=2.075 $X2=-0.19
+ $Y2=-0.24
cc_811 N_A_533_47#_c_914_n N_D[1]_c_1028_n 0.00712672f $X=3.275 $Y=1.34
+ $X2=-0.19 $Y2=-0.24
cc_812 N_A_533_47#_c_917_n N_VPWR_c_2824_n 0.0292866f $X=2.825 $Y=2.31 $X2=0
+ $Y2=0
cc_813 N_A_533_47#_c_913_n N_VPWR_c_2824_n 0.00688579f $X=3.055 $Y=1.405 $X2=0
+ $Y2=0
cc_814 N_A_533_47#_M1017_g N_VPWR_c_2826_n 0.00258498f $X=3.58 $Y=2.075 $X2=0
+ $Y2=0
cc_815 N_A_533_47#_M1039_d VPWR 0.00179197f $X=2.68 $Y=1.485 $X2=0 $Y2=0
cc_816 N_A_533_47#_M1017_g VPWR 0.00387928f $X=3.58 $Y=2.075 $X2=0 $Y2=0
cc_817 N_A_533_47#_c_917_n VPWR 0.00594162f $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_818 N_A_533_47#_c_917_n N_VPWR_c_2850_n 0.0210596f $X=2.825 $Y=2.31 $X2=0
+ $Y2=0
cc_819 N_A_533_47#_M1017_g N_Z_c_3367_n 0.00544362f $X=3.58 $Y=2.075 $X2=0 $Y2=0
cc_820 N_A_533_47#_c_917_n N_Z_c_3367_n 0.0371028f $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_821 N_A_533_47#_c_912_n N_Z_c_3321_n 0.00611965f $X=3.055 $Y=1.175 $X2=0
+ $Y2=0
cc_822 N_A_533_47#_c_915_n N_Z_c_3321_n 0.0259454f $X=2.825 $Y=0.495 $X2=0 $Y2=0
cc_823 N_A_533_47#_M1017_g N_Z_c_3323_n 0.00862328f $X=3.58 $Y=2.075 $X2=0 $Y2=0
cc_824 N_A_533_47#_c_917_n N_Z_c_3323_n 0.00378484f $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_825 N_A_533_47#_c_912_n N_Z_c_3323_n 0.00719188f $X=3.055 $Y=1.175 $X2=0
+ $Y2=0
cc_826 N_A_533_47#_c_913_n N_Z_c_3323_n 0.0304368f $X=3.055 $Y=1.405 $X2=0 $Y2=0
cc_827 N_A_533_47#_c_914_n N_Z_c_3323_n 0.00814206f $X=3.275 $Y=1.34 $X2=0 $Y2=0
cc_828 N_A_533_47#_M1017_g N_Z_c_3398_n 0.00335035f $X=3.58 $Y=2.075 $X2=0 $Y2=0
cc_829 N_A_533_47#_M1017_g N_Z_c_3400_n 0.00502861f $X=3.58 $Y=2.075 $X2=0 $Y2=0
cc_830 N_A_533_47#_c_912_n N_Z_c_3355_n 0.0124144f $X=3.055 $Y=1.175 $X2=0 $Y2=0
cc_831 N_A_533_47#_c_913_n N_Z_c_3355_n 0.00398133f $X=3.055 $Y=1.405 $X2=0
+ $Y2=0
cc_832 N_A_533_47#_c_914_n N_Z_c_3355_n 0.00349316f $X=3.275 $Y=1.34 $X2=0 $Y2=0
cc_833 N_A_533_47#_c_917_n N_Z_c_3419_n 0.0291787f $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_834 N_A_533_47#_c_913_n N_Z_c_3419_n 0.0126642f $X=3.055 $Y=1.405 $X2=0 $Y2=0
cc_835 N_A_533_47#_M1017_g N_Z_c_3549_n 0.00289142f $X=3.58 $Y=2.075 $X2=0 $Y2=0
cc_836 N_A_533_47#_c_917_n N_Z_c_3549_n 6.03258e-19 $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_837 N_A_533_47#_c_913_n N_Z_c_3549_n 4.25753e-19 $X=3.055 $Y=1.405 $X2=0
+ $Y2=0
cc_838 N_A_533_47#_M1017_g N_Z_c_3429_n 0.0107335f $X=3.58 $Y=2.075 $X2=0 $Y2=0
cc_839 N_A_533_47#_c_917_n N_Z_c_3429_n 0.0139746f $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_840 N_A_533_47#_c_913_n N_Z_c_3429_n 0.00749574f $X=3.055 $Y=1.405 $X2=0
+ $Y2=0
cc_841 N_A_533_47#_c_914_n N_Z_c_3429_n 0.00449418f $X=3.275 $Y=1.34 $X2=0 $Y2=0
cc_842 N_A_533_47#_M1055_d VGND 0.00358139f $X=2.665 $Y=0.235 $X2=0 $Y2=0
cc_843 N_A_533_47#_c_915_n VGND 0.0150148f $X=2.825 $Y=0.495 $X2=0 $Y2=0
cc_844 N_A_533_47#_c_915_n N_VGND_c_4407_n 0.015238f $X=2.825 $Y=0.495 $X2=0
+ $Y2=0
cc_845 N_A_533_937#_M1071_g N_D[9]_c_1069_n 0.0390641f $X=3.58 $Y=3.365
+ $X2=-0.19 $Y2=-0.24
cc_846 N_A_533_937#_c_971_n N_D[9]_c_1069_n 0.00216577f $X=3.275 $Y=4.1
+ $X2=-0.19 $Y2=-0.24
cc_847 N_A_533_937#_c_971_n N_D[9]_c_1066_n 0.00496096f $X=3.275 $Y=4.1 $X2=0
+ $Y2=0
cc_848 N_A_533_937#_c_974_n N_VPWR_c_2825_n 0.0292866f $X=2.825 $Y=3.13 $X2=0
+ $Y2=0
cc_849 N_A_533_937#_c_970_n N_VPWR_c_2825_n 0.00688579f $X=3.055 $Y=4.035 $X2=0
+ $Y2=0
cc_850 N_A_533_937#_M1071_g N_VPWR_c_2827_n 0.00258498f $X=3.58 $Y=3.365 $X2=0
+ $Y2=0
cc_851 N_A_533_937#_M1042_d VPWR 0.00179197f $X=2.68 $Y=2.955 $X2=0 $Y2=0
cc_852 N_A_533_937#_M1071_g VPWR 0.00387928f $X=3.58 $Y=3.365 $X2=0 $Y2=0
cc_853 N_A_533_937#_c_974_n VPWR 0.00594162f $X=2.825 $Y=3.13 $X2=0 $Y2=0
cc_854 N_A_533_937#_c_974_n N_VPWR_c_2850_n 0.0210596f $X=2.825 $Y=3.13 $X2=0
+ $Y2=0
cc_855 N_A_533_937#_M1071_g N_Z_c_3368_n 0.00544362f $X=3.58 $Y=3.365 $X2=0
+ $Y2=0
cc_856 N_A_533_937#_c_969_n N_Z_c_3322_n 0.00611965f $X=3.055 $Y=4.685 $X2=0
+ $Y2=0
cc_857 N_A_533_937#_c_972_n N_Z_c_3322_n 0.0259454f $X=2.825 $Y=4.945 $X2=0
+ $Y2=0
cc_858 N_A_533_937#_M1071_g N_Z_c_3324_n 0.00862328f $X=3.58 $Y=3.365 $X2=0
+ $Y2=0
cc_859 N_A_533_937#_c_974_n N_Z_c_3324_n 0.00378484f $X=2.825 $Y=3.13 $X2=0
+ $Y2=0
cc_860 N_A_533_937#_c_969_n N_Z_c_3324_n 0.00719188f $X=3.055 $Y=4.685 $X2=0
+ $Y2=0
cc_861 N_A_533_937#_c_970_n N_Z_c_3324_n 0.0304368f $X=3.055 $Y=4.035 $X2=0
+ $Y2=0
cc_862 N_A_533_937#_c_971_n N_Z_c_3324_n 0.00814206f $X=3.275 $Y=4.1 $X2=0 $Y2=0
cc_863 N_A_533_937#_M1071_g N_Z_c_3399_n 0.00335035f $X=3.58 $Y=3.365 $X2=0
+ $Y2=0
cc_864 N_A_533_937#_c_974_n N_Z_c_3399_n 0.0371028f $X=2.825 $Y=3.13 $X2=0 $Y2=0
cc_865 N_A_533_937#_M1071_g N_Z_c_3400_n 0.00502861f $X=3.58 $Y=3.365 $X2=0
+ $Y2=0
cc_866 N_A_533_937#_c_969_n N_Z_c_3356_n 0.0124144f $X=3.055 $Y=4.685 $X2=0
+ $Y2=0
cc_867 N_A_533_937#_c_970_n N_Z_c_3356_n 0.00398133f $X=3.055 $Y=4.035 $X2=0
+ $Y2=0
cc_868 N_A_533_937#_c_971_n N_Z_c_3356_n 0.00349316f $X=3.275 $Y=4.1 $X2=0 $Y2=0
cc_869 N_A_533_937#_c_974_n N_Z_c_3420_n 0.0291787f $X=2.825 $Y=3.13 $X2=0 $Y2=0
cc_870 N_A_533_937#_c_970_n N_Z_c_3420_n 0.0126642f $X=3.055 $Y=4.035 $X2=0
+ $Y2=0
cc_871 N_A_533_937#_M1071_g N_Z_c_3572_n 0.00289142f $X=3.58 $Y=3.365 $X2=0
+ $Y2=0
cc_872 N_A_533_937#_c_974_n N_Z_c_3572_n 6.03258e-19 $X=2.825 $Y=3.13 $X2=0
+ $Y2=0
cc_873 N_A_533_937#_c_970_n N_Z_c_3572_n 4.25753e-19 $X=3.055 $Y=4.035 $X2=0
+ $Y2=0
cc_874 N_A_533_937#_M1071_g N_Z_c_3430_n 0.0107344f $X=3.58 $Y=3.365 $X2=0 $Y2=0
cc_875 N_A_533_937#_c_974_n N_Z_c_3430_n 0.0139746f $X=2.825 $Y=3.13 $X2=0 $Y2=0
cc_876 N_A_533_937#_c_970_n N_Z_c_3430_n 0.00749574f $X=3.055 $Y=4.035 $X2=0
+ $Y2=0
cc_877 N_A_533_937#_c_971_n N_Z_c_3430_n 0.00449418f $X=3.275 $Y=4.1 $X2=0 $Y2=0
cc_878 N_A_533_937#_M1031_d VGND 0.00358139f $X=2.665 $Y=4.685 $X2=0 $Y2=0
cc_879 N_A_533_937#_c_972_n VGND 0.0150148f $X=2.825 $Y=4.945 $X2=0 $Y2=0
cc_880 N_A_533_937#_c_972_n N_VGND_c_4408_n 0.015238f $X=2.825 $Y=4.945 $X2=0
+ $Y2=0
cc_881 N_D[1]_c_1028_n N_D[9]_c_1069_n 0.0129371f $X=4.105 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_882 N_D[1]_c_1029_n N_D[2]_c_1107_n 0.00915308f $X=4.13 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_883 N_D[1]_c_1028_n N_D[2]_c_1108_n 0.0270908f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_884 N_D[1]_c_1031_n N_D[2]_c_1108_n 9.4377e-19 $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_885 N_D[1]_c_1030_n N_D[2]_c_1109_n 0.00442615f $X=3.955 $Y=1.055 $X2=0 $Y2=0
cc_886 N_D[1]_c_1028_n N_D[2]_c_1110_n 9.4377e-19 $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_887 N_D[1]_c_1031_n N_D[2]_c_1110_n 0.0199139f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_888 N_D[1]_c_1028_n N_VPWR_c_2826_n 0.0220781f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_889 N_D[1]_c_1031_n N_VPWR_c_2826_n 0.0044581f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_890 N_D[1]_c_1028_n VPWR 0.00468368f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_891 N_D[1]_c_1028_n N_VPWR_c_2851_n 0.00342413f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_892 N_D[1]_c_1028_n N_Z_c_3367_n 0.00176496f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_893 N_D[1]_c_1030_n N_Z_c_3321_n 0.00686805f $X=3.955 $Y=1.055 $X2=0 $Y2=0
cc_894 N_D[1]_c_1028_n N_Z_c_3323_n 0.00605747f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_895 N_D[1]_c_1030_n N_Z_c_3323_n 0.00376465f $X=3.955 $Y=1.055 $X2=0 $Y2=0
cc_896 N_D[1]_c_1031_n N_Z_c_3323_n 0.0216525f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_897 N_D[1]_c_1030_n N_Z_c_3355_n 0.0128881f $X=3.955 $Y=1.055 $X2=0 $Y2=0
cc_898 N_D[1]_c_1028_n N_Z_c_3585_n 0.00719456f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_899 N_D[1]_c_1031_n N_Z_c_3585_n 0.00989895f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_900 N_D[1]_c_1028_n N_Z_c_3429_n 8.42164e-19 $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_901 N_D[1]_c_1029_n N_VGND_c_4373_n 0.00322791f $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_902 N_D[1]_c_1031_n N_VGND_c_4373_n 0.00222881f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_903 N_D[1]_c_1029_n VGND 0.0108306f $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_904 N_D[1]_c_1061_p VGND 0.00942277f $X=3.955 $Y=0.51 $X2=0 $Y2=0
cc_905 N_D[1]_c_1029_n N_VGND_c_4407_n 0.00585385f $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_906 N_D[1]_c_1061_p N_VGND_c_4407_n 0.00842546f $X=3.955 $Y=0.51 $X2=0 $Y2=0
cc_907 N_D[1]_c_1030_n A_746_47# 0.00426617f $X=3.955 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_908 N_D[1]_c_1061_p A_746_47# 0.00894235f $X=3.955 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_909 N_D[9]_c_1066_n N_D[10]_c_1145_n 0.0287172f $X=4.13 $Y=4.445 $X2=-0.19
+ $Y2=-0.24
cc_910 N_D[9]_c_1068_n N_D[10]_c_1145_n 9.4377e-19 $X=4.1 $Y=4.28 $X2=-0.19
+ $Y2=-0.24
cc_911 N_D[9]_c_1069_n N_D[10]_c_1149_n 0.00752667f $X=4.105 $Y=4.03 $X2=0 $Y2=0
cc_912 N_D[9]_c_1067_n N_D[10]_c_1146_n 0.00442615f $X=3.955 $Y=4.815 $X2=0
+ $Y2=0
cc_913 N_D[9]_c_1066_n N_D[10]_c_1147_n 9.4377e-19 $X=4.13 $Y=4.445 $X2=0 $Y2=0
cc_914 N_D[9]_c_1068_n N_D[10]_c_1147_n 0.0199139f $X=4.1 $Y=4.28 $X2=0 $Y2=0
cc_915 N_D[9]_c_1069_n N_VPWR_c_2827_n 0.0220781f $X=4.105 $Y=4.03 $X2=0 $Y2=0
cc_916 N_D[9]_c_1068_n N_VPWR_c_2827_n 0.0044581f $X=4.1 $Y=4.28 $X2=0 $Y2=0
cc_917 N_D[9]_c_1069_n VPWR 0.00468368f $X=4.105 $Y=4.03 $X2=0 $Y2=0
cc_918 N_D[9]_c_1069_n N_VPWR_c_2851_n 0.00342413f $X=4.105 $Y=4.03 $X2=0 $Y2=0
cc_919 N_D[9]_c_1067_n N_Z_c_3322_n 0.00686805f $X=3.955 $Y=4.815 $X2=0 $Y2=0
cc_920 N_D[9]_c_1069_n N_Z_c_3324_n 0.00305841f $X=4.105 $Y=4.03 $X2=0 $Y2=0
cc_921 N_D[9]_c_1066_n N_Z_c_3324_n 0.00299906f $X=4.13 $Y=4.445 $X2=0 $Y2=0
cc_922 N_D[9]_c_1067_n N_Z_c_3324_n 0.00376465f $X=3.955 $Y=4.815 $X2=0 $Y2=0
cc_923 N_D[9]_c_1068_n N_Z_c_3324_n 0.0216525f $X=4.1 $Y=4.28 $X2=0 $Y2=0
cc_924 N_D[9]_c_1069_n N_Z_c_3400_n 0.00176496f $X=4.105 $Y=4.03 $X2=0 $Y2=0
cc_925 N_D[9]_c_1067_n N_Z_c_3356_n 0.0128881f $X=3.955 $Y=4.815 $X2=0 $Y2=0
cc_926 N_D[9]_c_1069_n N_Z_c_3595_n 0.0061664f $X=4.105 $Y=4.03 $X2=0 $Y2=0
cc_927 N_D[9]_c_1066_n N_Z_c_3595_n 0.00102816f $X=4.13 $Y=4.445 $X2=0 $Y2=0
cc_928 N_D[9]_c_1068_n N_Z_c_3595_n 0.00989895f $X=4.1 $Y=4.28 $X2=0 $Y2=0
cc_929 N_D[9]_c_1069_n N_Z_c_3430_n 8.42164e-19 $X=4.105 $Y=4.03 $X2=0 $Y2=0
cc_930 N_D[9]_c_1066_n N_VGND_c_4374_n 0.00322791f $X=4.13 $Y=4.445 $X2=0 $Y2=0
cc_931 N_D[9]_c_1068_n N_VGND_c_4374_n 0.00222881f $X=4.1 $Y=4.28 $X2=0 $Y2=0
cc_932 N_D[9]_c_1066_n VGND 0.0108306f $X=4.13 $Y=4.445 $X2=0 $Y2=0
cc_933 N_D[9]_c_1102_p VGND 0.00941728f $X=3.955 $Y=4.93 $X2=0 $Y2=0
cc_934 N_D[9]_c_1066_n N_VGND_c_4408_n 0.00585385f $X=4.13 $Y=4.445 $X2=0 $Y2=0
cc_935 N_D[9]_c_1102_p N_VGND_c_4408_n 0.00842546f $X=3.955 $Y=4.93 $X2=0 $Y2=0
cc_936 N_D[9]_c_1067_n A_746_937# 0.00426617f $X=3.955 $Y=4.815 $X2=-0.19
+ $Y2=-0.24
cc_937 N_D[9]_c_1102_p A_746_937# 0.00894235f $X=3.955 $Y=4.93 $X2=-0.19
+ $Y2=-0.24
cc_938 N_D[2]_c_1108_n N_D[10]_c_1149_n 0.0129371f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_939 N_D[2]_c_1108_n N_A_1012_265#_M1041_g 0.0390641f $X=4.635 $Y=1.41 $X2=0
+ $Y2=0
cc_940 N_D[2]_c_1108_n N_A_1012_265#_c_1189_n 0.00712672f $X=4.635 $Y=1.41 $X2=0
+ $Y2=0
cc_941 N_D[2]_c_1107_n N_S[2]_c_1300_n 0.0286599f $X=4.61 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_942 N_D[2]_c_1109_n N_S[2]_c_1300_n 0.00289497f $X=4.785 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_943 N_D[2]_c_1108_n N_VPWR_c_2826_n 0.0220781f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_944 N_D[2]_c_1110_n N_VPWR_c_2826_n 0.0044581f $X=4.785 $Y=1.19 $X2=0 $Y2=0
cc_945 N_D[2]_c_1108_n VPWR 0.00468368f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_946 N_D[2]_c_1108_n N_VPWR_c_2852_n 0.00342413f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_947 N_D[2]_c_1108_n N_Z_c_3325_n 0.00605747f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_948 N_D[2]_c_1109_n N_Z_c_3325_n 0.00376465f $X=4.785 $Y=1.055 $X2=0 $Y2=0
cc_949 N_D[2]_c_1110_n N_Z_c_3325_n 0.0216525f $X=4.785 $Y=1.19 $X2=0 $Y2=0
cc_950 N_D[2]_c_1109_n N_Z_c_3327_n 0.0128881f $X=4.785 $Y=1.055 $X2=0 $Y2=0
cc_951 N_D[2]_c_1109_n N_Z_c_3328_n 0.00686805f $X=4.785 $Y=1.055 $X2=0 $Y2=0
cc_952 N_D[2]_c_1108_n N_Z_c_3373_n 0.00176496f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_953 N_D[2]_c_1108_n N_Z_c_3585_n 0.00719456f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_954 N_D[2]_c_1110_n N_Z_c_3585_n 0.00989895f $X=4.785 $Y=1.19 $X2=0 $Y2=0
cc_955 N_D[2]_c_1108_n N_Z_c_3431_n 8.42164e-19 $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_956 N_D[2]_c_1107_n N_VGND_c_4373_n 0.00322791f $X=4.61 $Y=0.995 $X2=0 $Y2=0
cc_957 N_D[2]_c_1110_n N_VGND_c_4373_n 0.00222881f $X=4.785 $Y=1.19 $X2=0 $Y2=0
cc_958 N_D[2]_c_1107_n N_VGND_c_4393_n 0.00585385f $X=4.61 $Y=0.995 $X2=0 $Y2=0
cc_959 D[2] N_VGND_c_4393_n 0.00842546f $X=4.745 $Y=0.425 $X2=0 $Y2=0
cc_960 N_D[2]_c_1107_n VGND 0.0108306f $X=4.61 $Y=0.995 $X2=0 $Y2=0
cc_961 D[2] VGND 0.00942277f $X=4.745 $Y=0.425 $X2=0 $Y2=0
cc_962 N_D[2]_c_1109_n A_937_47# 0.00426617f $X=4.785 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_963 D[2] A_937_47# 0.00894235f $X=4.745 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_964 N_D[10]_c_1149_n N_A_1012_793#_M1000_g 0.0390641f $X=4.635 $Y=4.03 $X2=0
+ $Y2=0
cc_965 N_D[10]_c_1145_n N_A_1012_793#_c_1246_n 0.00496096f $X=4.61 $Y=4.445
+ $X2=0 $Y2=0
cc_966 N_D[10]_c_1149_n N_A_1012_793#_c_1246_n 0.00216577f $X=4.635 $Y=4.03
+ $X2=0 $Y2=0
cc_967 N_D[10]_c_1145_n N_S[10]_c_1351_n 0.0286599f $X=4.61 $Y=4.445 $X2=0 $Y2=0
cc_968 N_D[10]_c_1146_n N_S[10]_c_1351_n 0.00289497f $X=4.785 $Y=4.815 $X2=0
+ $Y2=0
cc_969 N_D[10]_c_1149_n N_VPWR_c_2827_n 0.0220781f $X=4.635 $Y=4.03 $X2=0 $Y2=0
cc_970 N_D[10]_c_1147_n N_VPWR_c_2827_n 0.0044581f $X=4.785 $Y=4.25 $X2=0 $Y2=0
cc_971 N_D[10]_c_1149_n VPWR 0.00468368f $X=4.635 $Y=4.03 $X2=0 $Y2=0
cc_972 N_D[10]_c_1149_n N_VPWR_c_2852_n 0.00342413f $X=4.635 $Y=4.03 $X2=0 $Y2=0
cc_973 N_D[10]_c_1145_n N_Z_c_3326_n 0.00299906f $X=4.61 $Y=4.445 $X2=0 $Y2=0
cc_974 N_D[10]_c_1149_n N_Z_c_3326_n 0.00305841f $X=4.635 $Y=4.03 $X2=0 $Y2=0
cc_975 N_D[10]_c_1146_n N_Z_c_3326_n 0.00376465f $X=4.785 $Y=4.815 $X2=0 $Y2=0
cc_976 N_D[10]_c_1147_n N_Z_c_3326_n 0.0216525f $X=4.785 $Y=4.25 $X2=0 $Y2=0
cc_977 N_D[10]_c_1146_n N_Z_c_3329_n 0.0128881f $X=4.785 $Y=4.815 $X2=0 $Y2=0
cc_978 N_D[10]_c_1146_n N_Z_c_3330_n 0.00686805f $X=4.785 $Y=4.815 $X2=0 $Y2=0
cc_979 N_D[10]_c_1149_n N_Z_c_3403_n 0.00176496f $X=4.635 $Y=4.03 $X2=0 $Y2=0
cc_980 N_D[10]_c_1145_n N_Z_c_3595_n 0.00102816f $X=4.61 $Y=4.445 $X2=0 $Y2=0
cc_981 N_D[10]_c_1149_n N_Z_c_3595_n 0.0061664f $X=4.635 $Y=4.03 $X2=0 $Y2=0
cc_982 N_D[10]_c_1147_n N_Z_c_3595_n 0.00989895f $X=4.785 $Y=4.25 $X2=0 $Y2=0
cc_983 N_D[10]_c_1149_n N_Z_c_3432_n 8.42164e-19 $X=4.635 $Y=4.03 $X2=0 $Y2=0
cc_984 N_D[10]_c_1145_n N_VGND_c_4374_n 0.00322791f $X=4.61 $Y=4.445 $X2=0 $Y2=0
cc_985 N_D[10]_c_1147_n N_VGND_c_4374_n 0.00222881f $X=4.785 $Y=4.25 $X2=0 $Y2=0
cc_986 N_D[10]_c_1145_n N_VGND_c_4395_n 0.00585385f $X=4.61 $Y=4.445 $X2=0 $Y2=0
cc_987 D[10] N_VGND_c_4395_n 0.00842546f $X=4.745 $Y=4.845 $X2=0 $Y2=0
cc_988 N_D[10]_c_1145_n VGND 0.0108306f $X=4.61 $Y=4.445 $X2=0 $Y2=0
cc_989 D[10] VGND 0.00941728f $X=4.745 $Y=4.845 $X2=0 $Y2=0
cc_990 N_D[10]_c_1146_n A_937_911# 0.00426617f $X=4.785 $Y=4.815 $X2=-0.19
+ $Y2=-0.24
cc_991 D[10] A_937_911# 0.00894235f $X=4.745 $Y=4.845 $X2=-0.19 $Y2=-0.24
cc_992 N_A_1012_265#_M1041_g N_A_1012_793#_M1000_g 0.0129371f $X=5.16 $Y=2.075
+ $X2=0 $Y2=0
cc_993 N_A_1012_265#_c_1186_n N_S[2]_c_1301_n 0.00827389f $X=5.685 $Y=0.755
+ $X2=0 $Y2=0
cc_994 N_A_1012_265#_c_1187_n N_S[2]_c_1301_n 0.0164662f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_995 N_A_1012_265#_c_1188_n N_S[2]_c_1301_n 0.00928634f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_996 N_A_1012_265#_c_1189_n N_S[2]_c_1301_n 0.0184911f $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_997 N_A_1012_265#_c_1189_n N_S[2]_c_1302_n 0.00820745f $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_998 N_A_1012_265#_c_1187_n N_S[2]_c_1303_n 0.0012443f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_999 N_A_1012_265#_c_1191_n N_S[2]_c_1303_n 0.00902681f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_1000 N_A_1012_265#_c_1188_n N_S[2]_c_1303_n 0.00767015f $X=5.915 $Y=1.63
+ $X2=0 $Y2=0
cc_1001 N_A_1012_265#_c_1189_n N_S[2]_c_1303_n 0.00659591f $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_1002 N_A_1012_265#_c_1187_n N_S[2]_c_1304_n 0.00219336f $X=5.685 $Y=1.175
+ $X2=0 $Y2=0
cc_1003 N_A_1012_265#_c_1186_n N_S[2]_c_1305_n 0.00603567f $X=5.685 $Y=0.755
+ $X2=0 $Y2=0
cc_1004 N_A_1012_265#_c_1187_n N_S[2]_c_1305_n 0.0178233f $X=5.685 $Y=1.175
+ $X2=0 $Y2=0
cc_1005 N_A_1012_265#_c_1188_n N_S[2]_c_1305_n 0.0214702f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_1006 N_A_1012_265#_c_1189_n N_S[2]_c_1305_n 2.59957e-19 $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_1007 N_A_1012_265#_M1041_g N_VPWR_c_2826_n 0.00258498f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_1008 N_A_1012_265#_c_1191_n N_VPWR_c_2828_n 0.0292866f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_1009 N_A_1012_265#_c_1188_n N_VPWR_c_2828_n 0.00688579f $X=5.915 $Y=1.63
+ $X2=0 $Y2=0
cc_1010 N_A_1012_265#_c_1191_n N_VPWR_c_2842_n 0.0210596f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_1011 N_A_1012_265#_M1050_s VPWR 0.00179197f $X=5.79 $Y=1.485 $X2=0 $Y2=0
cc_1012 N_A_1012_265#_M1041_g VPWR 0.00387928f $X=5.16 $Y=2.075 $X2=0 $Y2=0
cc_1013 N_A_1012_265#_c_1191_n VPWR 0.00594162f $X=5.915 $Y=2.31 $X2=0 $Y2=0
cc_1014 N_A_1012_265#_M1041_g N_Z_c_3325_n 0.00862328f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_1015 N_A_1012_265#_c_1187_n N_Z_c_3325_n 0.00719188f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_1016 N_A_1012_265#_c_1191_n N_Z_c_3325_n 0.00378484f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_1017 N_A_1012_265#_c_1188_n N_Z_c_3325_n 0.0304368f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_1018 N_A_1012_265#_c_1189_n N_Z_c_3325_n 0.00814206f $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_1019 N_A_1012_265#_c_1187_n N_Z_c_3327_n 0.0124144f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_1020 N_A_1012_265#_c_1188_n N_Z_c_3327_n 0.00398133f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_1021 N_A_1012_265#_c_1189_n N_Z_c_3327_n 0.00349316f $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_1022 N_A_1012_265#_c_1186_n N_Z_c_3328_n 0.0259454f $X=5.685 $Y=0.755 $X2=0
+ $Y2=0
cc_1023 N_A_1012_265#_c_1187_n N_Z_c_3328_n 0.00611965f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_1024 N_A_1012_265#_M1041_g N_Z_c_3373_n 0.00544362f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_1025 N_A_1012_265#_c_1191_n N_Z_c_3373_n 0.0371028f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_1026 N_A_1012_265#_M1041_g N_Z_c_3401_n 0.00335035f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_1027 N_A_1012_265#_M1041_g N_Z_c_3403_n 0.00502861f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_1028 N_A_1012_265#_c_1191_n N_Z_c_3421_n 0.0291787f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_1029 N_A_1012_265#_c_1188_n N_Z_c_3421_n 0.0126642f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_1030 N_A_1012_265#_M1041_g N_Z_c_3635_n 0.00289142f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_1031 N_A_1012_265#_c_1191_n N_Z_c_3635_n 6.03258e-19 $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_1032 N_A_1012_265#_c_1188_n N_Z_c_3635_n 4.25753e-19 $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_1033 N_A_1012_265#_M1041_g N_Z_c_3431_n 0.0107335f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_1034 N_A_1012_265#_c_1191_n N_Z_c_3431_n 0.0139746f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_1035 N_A_1012_265#_c_1188_n N_Z_c_3431_n 0.00749574f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_1036 N_A_1012_265#_c_1189_n N_Z_c_3431_n 0.00449418f $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_1037 N_A_1012_265#_c_1186_n N_VGND_c_4393_n 0.015238f $X=5.685 $Y=0.755 $X2=0
+ $Y2=0
cc_1038 N_A_1012_265#_M1088_s VGND 0.00358139f $X=5.79 $Y=0.235 $X2=0 $Y2=0
cc_1039 N_A_1012_265#_c_1186_n VGND 0.0150148f $X=5.685 $Y=0.755 $X2=0 $Y2=0
cc_1040 N_A_1012_793#_c_1244_n N_S[10]_c_1350_n 0.0247401f $X=5.685 $Y=4.685
+ $X2=0 $Y2=0
cc_1041 N_A_1012_793#_c_1245_n N_S[10]_c_1350_n 0.00928634f $X=5.915 $Y=3.805
+ $X2=0 $Y2=0
cc_1042 N_A_1012_793#_c_1246_n N_S[10]_c_1350_n 0.0184911f $X=5.16 $Y=4.1 $X2=0
+ $Y2=0
cc_1043 N_A_1012_793#_c_1246_n N_S[10]_c_1351_n 0.00820745f $X=5.16 $Y=4.1 $X2=0
+ $Y2=0
cc_1044 N_A_1012_793#_c_1245_n N_S[10]_c_1354_n 0.00382813f $X=5.915 $Y=3.805
+ $X2=0 $Y2=0
cc_1045 N_A_1012_793#_c_1249_n N_S[10]_c_1354_n 0.00902681f $X=5.915 $Y=3.13
+ $X2=0 $Y2=0
cc_1046 N_A_1012_793#_c_1246_n N_S[10]_c_1354_n 0.00150889f $X=5.16 $Y=4.1 $X2=0
+ $Y2=0
cc_1047 N_A_1012_793#_c_1244_n N_S[10]_c_1352_n 0.00343766f $X=5.685 $Y=4.685
+ $X2=0 $Y2=0
cc_1048 N_A_1012_793#_c_1245_n N_S[10]_c_1352_n 0.00384202f $X=5.915 $Y=3.805
+ $X2=0 $Y2=0
cc_1049 N_A_1012_793#_c_1246_n N_S[10]_c_1352_n 0.00508702f $X=5.16 $Y=4.1 $X2=0
+ $Y2=0
cc_1050 N_A_1012_793#_c_1244_n S[10] 0.023859f $X=5.685 $Y=4.685 $X2=0 $Y2=0
cc_1051 N_A_1012_793#_c_1245_n S[10] 0.0214702f $X=5.915 $Y=3.805 $X2=0 $Y2=0
cc_1052 N_A_1012_793#_c_1246_n S[10] 2.59957e-19 $X=5.16 $Y=4.1 $X2=0 $Y2=0
cc_1053 N_A_1012_793#_M1000_g N_VPWR_c_2827_n 0.00258498f $X=5.16 $Y=3.365 $X2=0
+ $Y2=0
cc_1054 N_A_1012_793#_c_1245_n N_VPWR_c_2829_n 0.00688579f $X=5.915 $Y=3.805
+ $X2=0 $Y2=0
cc_1055 N_A_1012_793#_c_1249_n N_VPWR_c_2829_n 0.0292866f $X=5.915 $Y=3.13 $X2=0
+ $Y2=0
cc_1056 N_A_1012_793#_c_1249_n N_VPWR_c_2842_n 0.0210596f $X=5.915 $Y=3.13 $X2=0
+ $Y2=0
cc_1057 N_A_1012_793#_M1053_s VPWR 0.00179197f $X=5.79 $Y=2.955 $X2=0 $Y2=0
cc_1058 N_A_1012_793#_M1000_g VPWR 0.00387928f $X=5.16 $Y=3.365 $X2=0 $Y2=0
cc_1059 N_A_1012_793#_c_1249_n VPWR 0.00594162f $X=5.915 $Y=3.13 $X2=0 $Y2=0
cc_1060 N_A_1012_793#_M1000_g N_Z_c_3326_n 0.00862328f $X=5.16 $Y=3.365 $X2=0
+ $Y2=0
cc_1061 N_A_1012_793#_c_1244_n N_Z_c_3326_n 0.00719188f $X=5.685 $Y=4.685 $X2=0
+ $Y2=0
cc_1062 N_A_1012_793#_c_1245_n N_Z_c_3326_n 0.0304368f $X=5.915 $Y=3.805 $X2=0
+ $Y2=0
cc_1063 N_A_1012_793#_c_1249_n N_Z_c_3326_n 0.00378484f $X=5.915 $Y=3.13 $X2=0
+ $Y2=0
cc_1064 N_A_1012_793#_c_1246_n N_Z_c_3326_n 0.00814206f $X=5.16 $Y=4.1 $X2=0
+ $Y2=0
cc_1065 N_A_1012_793#_c_1244_n N_Z_c_3329_n 0.0124144f $X=5.685 $Y=4.685 $X2=0
+ $Y2=0
cc_1066 N_A_1012_793#_c_1245_n N_Z_c_3329_n 0.00398133f $X=5.915 $Y=3.805 $X2=0
+ $Y2=0
cc_1067 N_A_1012_793#_c_1246_n N_Z_c_3329_n 0.00349316f $X=5.16 $Y=4.1 $X2=0
+ $Y2=0
cc_1068 N_A_1012_793#_c_1244_n N_Z_c_3330_n 0.032065f $X=5.685 $Y=4.685 $X2=0
+ $Y2=0
cc_1069 N_A_1012_793#_M1000_g N_Z_c_3374_n 0.00544362f $X=5.16 $Y=3.365 $X2=0
+ $Y2=0
cc_1070 N_A_1012_793#_M1000_g N_Z_c_3402_n 0.00335035f $X=5.16 $Y=3.365 $X2=0
+ $Y2=0
cc_1071 N_A_1012_793#_c_1249_n N_Z_c_3402_n 0.0371028f $X=5.915 $Y=3.13 $X2=0
+ $Y2=0
cc_1072 N_A_1012_793#_M1000_g N_Z_c_3403_n 0.00502861f $X=5.16 $Y=3.365 $X2=0
+ $Y2=0
cc_1073 N_A_1012_793#_c_1245_n N_Z_c_3422_n 0.0126642f $X=5.915 $Y=3.805 $X2=0
+ $Y2=0
cc_1074 N_A_1012_793#_c_1249_n N_Z_c_3422_n 0.0291787f $X=5.915 $Y=3.13 $X2=0
+ $Y2=0
cc_1075 N_A_1012_793#_M1000_g N_Z_c_3657_n 0.00289142f $X=5.16 $Y=3.365 $X2=0
+ $Y2=0
cc_1076 N_A_1012_793#_c_1245_n N_Z_c_3657_n 4.25753e-19 $X=5.915 $Y=3.805 $X2=0
+ $Y2=0
cc_1077 N_A_1012_793#_c_1249_n N_Z_c_3657_n 6.03258e-19 $X=5.915 $Y=3.13 $X2=0
+ $Y2=0
cc_1078 N_A_1012_793#_M1000_g N_Z_c_3432_n 0.0107344f $X=5.16 $Y=3.365 $X2=0
+ $Y2=0
cc_1079 N_A_1012_793#_c_1245_n N_Z_c_3432_n 0.00749574f $X=5.915 $Y=3.805 $X2=0
+ $Y2=0
cc_1080 N_A_1012_793#_c_1249_n N_Z_c_3432_n 0.0139746f $X=5.915 $Y=3.13 $X2=0
+ $Y2=0
cc_1081 N_A_1012_793#_c_1246_n N_Z_c_3432_n 0.00449418f $X=5.16 $Y=4.1 $X2=0
+ $Y2=0
cc_1082 N_A_1012_793#_c_1244_n N_VGND_c_4395_n 0.015238f $X=5.685 $Y=4.685 $X2=0
+ $Y2=0
cc_1083 N_A_1012_793#_M1082_s VGND 0.00358139f $X=5.79 $Y=4.685 $X2=0 $Y2=0
cc_1084 N_A_1012_793#_c_1244_n VGND 0.0150148f $X=5.685 $Y=4.685 $X2=0 $Y2=0
cc_1085 N_S[2]_c_1303_n N_S[10]_c_1354_n 0.0130744f $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_1086 N_S[2]_c_1303_n N_S[3]_c_1397_n 0.0578733f $X=6.15 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_1087 N_S[2]_c_1305_n N_S[3]_c_1397_n 0.00112057f $X=6.115 $Y=1.03 $X2=-0.19
+ $Y2=-0.24
cc_1088 N_S[2]_c_1304_n N_S[3]_c_1398_n 0.0091402f $X=6.15 $Y=0.83 $X2=0 $Y2=0
cc_1089 N_S[2]_c_1303_n N_S[3]_c_1401_n 0.00112057f $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_1090 N_S[2]_c_1305_n N_S[3]_c_1401_n 0.0277403f $X=6.115 $Y=1.03 $X2=0 $Y2=0
cc_1091 N_S[2]_c_1303_n N_VPWR_c_2828_n 0.00965725f $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_1092 N_S[2]_c_1305_n N_VPWR_c_2828_n 0.00587376f $X=6.115 $Y=1.03 $X2=0 $Y2=0
cc_1093 N_S[2]_c_1303_n N_VPWR_c_2842_n 0.0035837f $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_1094 N_S[2]_c_1303_n VPWR 0.0072999f $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_1095 N_S[2]_c_1302_n N_Z_c_3325_n 7.46972e-19 $X=5.16 $Y=0.905 $X2=0 $Y2=0
cc_1096 N_S[2]_c_1301_n N_Z_c_3327_n 0.00806549f $X=5.98 $Y=0.905 $X2=0 $Y2=0
cc_1097 N_S[2]_c_1302_n N_Z_c_3327_n 0.00605736f $X=5.16 $Y=0.905 $X2=0 $Y2=0
cc_1098 N_S[2]_c_1300_n N_Z_c_3328_n 0.00316445f $X=5.085 $Y=0.83 $X2=0 $Y2=0
cc_1099 N_S[2]_c_1301_n N_Z_c_3328_n 0.00501353f $X=5.98 $Y=0.905 $X2=0 $Y2=0
cc_1100 N_S[2]_c_1303_n N_Z_c_3403_n 0.00124373f $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_1101 N_S[2]_c_1303_n N_Z_c_3421_n 0.0062071f $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_1102 N_S[2]_c_1305_n N_Z_c_3421_n 0.00659242f $X=6.115 $Y=1.03 $X2=0 $Y2=0
cc_1103 N_S[2]_c_1304_n N_VGND_c_4375_n 0.00570474f $X=6.15 $Y=0.83 $X2=0 $Y2=0
cc_1104 N_S[2]_c_1305_n N_VGND_c_4375_n 0.00391126f $X=6.115 $Y=1.03 $X2=0 $Y2=0
cc_1105 N_S[2]_c_1300_n N_VGND_c_4393_n 0.00585385f $X=5.085 $Y=0.83 $X2=0 $Y2=0
cc_1106 N_S[2]_c_1304_n N_VGND_c_4393_n 0.00585385f $X=6.15 $Y=0.83 $X2=0 $Y2=0
cc_1107 N_S[2]_c_1300_n VGND 0.00880034f $X=5.085 $Y=0.83 $X2=0 $Y2=0
cc_1108 N_S[2]_c_1301_n VGND 0.00349917f $X=5.98 $Y=0.905 $X2=0 $Y2=0
cc_1109 N_S[2]_c_1303_n VGND 6.15795e-19 $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_1110 N_S[2]_c_1304_n VGND 0.0124506f $X=6.15 $Y=0.83 $X2=0 $Y2=0
cc_1111 N_S[10]_c_1354_n N_S[11]_c_1447_n 0.0296874f $X=6.15 $Y=4.03 $X2=-0.19
+ $Y2=-0.24
cc_1112 N_S[10]_c_1352_n N_S[11]_c_1443_n 0.0373261f $X=6.15 $Y=4.61 $X2=0 $Y2=0
cc_1113 S[10] N_S[11]_c_1443_n 0.00112057f $X=6.125 $Y=4.165 $X2=0 $Y2=0
cc_1114 N_S[10]_c_1352_n S[11] 0.00112057f $X=6.15 $Y=4.61 $X2=0 $Y2=0
cc_1115 S[10] S[11] 0.0277403f $X=6.125 $Y=4.165 $X2=0 $Y2=0
cc_1116 N_S[10]_c_1354_n N_VPWR_c_2829_n 0.00965725f $X=6.15 $Y=4.03 $X2=0 $Y2=0
cc_1117 S[10] N_VPWR_c_2829_n 0.00587376f $X=6.125 $Y=4.165 $X2=0 $Y2=0
cc_1118 N_S[10]_c_1354_n N_VPWR_c_2842_n 0.0035837f $X=6.15 $Y=4.03 $X2=0 $Y2=0
cc_1119 N_S[10]_c_1354_n VPWR 0.0072999f $X=6.15 $Y=4.03 $X2=0 $Y2=0
cc_1120 N_S[10]_c_1351_n N_Z_c_3326_n 7.46972e-19 $X=5.16 $Y=4.535 $X2=0 $Y2=0
cc_1121 N_S[10]_c_1350_n N_Z_c_3329_n 0.00806549f $X=5.98 $Y=4.535 $X2=0 $Y2=0
cc_1122 N_S[10]_c_1351_n N_Z_c_3329_n 0.00605736f $X=5.16 $Y=4.535 $X2=0 $Y2=0
cc_1123 N_S[10]_c_1349_n N_Z_c_3330_n 0.00316445f $X=5.085 $Y=4.61 $X2=0 $Y2=0
cc_1124 N_S[10]_c_1350_n N_Z_c_3330_n 0.00501353f $X=5.98 $Y=4.535 $X2=0 $Y2=0
cc_1125 N_S[10]_c_1354_n N_Z_c_3403_n 0.00124373f $X=6.15 $Y=4.03 $X2=0 $Y2=0
cc_1126 N_S[10]_c_1354_n N_Z_c_3422_n 0.00597491f $X=6.15 $Y=4.03 $X2=0 $Y2=0
cc_1127 N_S[10]_c_1352_n N_Z_c_3422_n 2.32192e-19 $X=6.15 $Y=4.61 $X2=0 $Y2=0
cc_1128 S[10] N_Z_c_3422_n 0.00659242f $X=6.125 $Y=4.165 $X2=0 $Y2=0
cc_1129 N_S[10]_c_1352_n N_VGND_c_4376_n 0.00570474f $X=6.15 $Y=4.61 $X2=0 $Y2=0
cc_1130 S[10] N_VGND_c_4376_n 0.00391126f $X=6.125 $Y=4.165 $X2=0 $Y2=0
cc_1131 N_S[10]_c_1349_n N_VGND_c_4395_n 0.00585385f $X=5.085 $Y=4.61 $X2=0
+ $Y2=0
cc_1132 N_S[10]_c_1352_n N_VGND_c_4395_n 0.00585385f $X=6.15 $Y=4.61 $X2=0 $Y2=0
cc_1133 N_S[10]_c_1349_n VGND 0.00880034f $X=5.085 $Y=4.61 $X2=0 $Y2=0
cc_1134 N_S[10]_c_1350_n VGND 0.00349917f $X=5.98 $Y=4.535 $X2=0 $Y2=0
cc_1135 N_S[10]_c_1352_n VGND 0.0130664f $X=6.15 $Y=4.61 $X2=0 $Y2=0
cc_1136 N_S[3]_c_1397_n N_S[11]_c_1447_n 0.0130744f $X=6.73 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_1137 N_S[3]_c_1397_n N_A_1361_47#_c_1495_n 0.00902681f $X=6.73 $Y=1.41 $X2=0
+ $Y2=0
cc_1138 N_S[3]_c_1397_n N_A_1361_47#_c_1490_n 0.0012443f $X=6.73 $Y=1.41 $X2=0
+ $Y2=0
cc_1139 N_S[3]_c_1398_n N_A_1361_47#_c_1490_n 0.00219336f $X=6.73 $Y=0.83 $X2=0
+ $Y2=0
cc_1140 N_S[3]_c_1399_n N_A_1361_47#_c_1490_n 0.0164662f $X=7.72 $Y=0.905 $X2=0
+ $Y2=0
cc_1141 N_S[3]_c_1401_n N_A_1361_47#_c_1490_n 0.0178233f $X=6.765 $Y=1.03 $X2=0
+ $Y2=0
cc_1142 N_S[3]_c_1397_n N_A_1361_47#_c_1491_n 0.00767015f $X=6.73 $Y=1.41 $X2=0
+ $Y2=0
cc_1143 N_S[3]_c_1399_n N_A_1361_47#_c_1491_n 0.00928634f $X=7.72 $Y=0.905 $X2=0
+ $Y2=0
cc_1144 N_S[3]_c_1401_n N_A_1361_47#_c_1491_n 0.0214702f $X=6.765 $Y=1.03 $X2=0
+ $Y2=0
cc_1145 N_S[3]_c_1397_n N_A_1361_47#_c_1492_n 0.00659591f $X=6.73 $Y=1.41 $X2=0
+ $Y2=0
cc_1146 N_S[3]_c_1399_n N_A_1361_47#_c_1492_n 0.0266986f $X=7.72 $Y=0.905 $X2=0
+ $Y2=0
cc_1147 N_S[3]_c_1401_n N_A_1361_47#_c_1492_n 2.59957e-19 $X=6.765 $Y=1.03 $X2=0
+ $Y2=0
cc_1148 N_S[3]_c_1397_n N_A_1361_47#_c_1493_n 0.00827389f $X=6.73 $Y=1.41 $X2=0
+ $Y2=0
cc_1149 N_S[3]_c_1401_n N_A_1361_47#_c_1493_n 0.00603567f $X=6.765 $Y=1.03 $X2=0
+ $Y2=0
cc_1150 N_S[3]_c_1400_n N_D[3]_c_1607_n 0.0286599f $X=7.795 $Y=0.83 $X2=0 $Y2=0
cc_1151 N_S[3]_c_1400_n N_D[3]_c_1608_n 0.00289497f $X=7.795 $Y=0.83 $X2=0 $Y2=0
cc_1152 N_S[3]_c_1397_n N_VPWR_c_2828_n 0.00965725f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_1153 N_S[3]_c_1401_n N_VPWR_c_2828_n 0.00587376f $X=6.765 $Y=1.03 $X2=0 $Y2=0
cc_1154 N_S[3]_c_1397_n VPWR 0.0072999f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_1155 N_S[3]_c_1397_n N_VPWR_c_2853_n 0.0035837f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_1156 N_S[3]_c_1399_n N_Z_c_3331_n 0.00501353f $X=7.72 $Y=0.905 $X2=0 $Y2=0
cc_1157 N_S[3]_c_1400_n N_Z_c_3331_n 0.00316445f $X=7.795 $Y=0.83 $X2=0 $Y2=0
cc_1158 N_S[3]_c_1399_n N_Z_c_3333_n 7.46972e-19 $X=7.72 $Y=0.905 $X2=0 $Y2=0
cc_1159 N_S[3]_c_1397_n N_Z_c_3406_n 0.00124373f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_1160 N_S[3]_c_1399_n N_Z_c_3357_n 0.0141229f $X=7.72 $Y=0.905 $X2=0 $Y2=0
cc_1161 N_S[3]_c_1397_n N_Z_c_3421_n 0.0062071f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_1162 N_S[3]_c_1401_n N_Z_c_3421_n 0.00659242f $X=6.765 $Y=1.03 $X2=0 $Y2=0
cc_1163 N_S[3]_c_1398_n N_VGND_c_4375_n 0.00570474f $X=6.73 $Y=0.83 $X2=0 $Y2=0
cc_1164 N_S[3]_c_1401_n N_VGND_c_4375_n 0.00391126f $X=6.765 $Y=1.03 $X2=0 $Y2=0
cc_1165 N_S[3]_c_1397_n VGND 6.15795e-19 $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_1166 N_S[3]_c_1398_n VGND 0.0124506f $X=6.73 $Y=0.83 $X2=0 $Y2=0
cc_1167 N_S[3]_c_1399_n VGND 0.00349917f $X=7.72 $Y=0.905 $X2=0 $Y2=0
cc_1168 N_S[3]_c_1400_n VGND 0.00880034f $X=7.795 $Y=0.83 $X2=0 $Y2=0
cc_1169 N_S[3]_c_1398_n N_VGND_c_4409_n 0.00585385f $X=6.73 $Y=0.83 $X2=0 $Y2=0
cc_1170 N_S[3]_c_1400_n N_VGND_c_4409_n 0.00585385f $X=7.795 $Y=0.83 $X2=0 $Y2=0
cc_1171 N_S[11]_c_1447_n N_A_1361_937#_c_1552_n 0.00902681f $X=6.73 $Y=4.03
+ $X2=0 $Y2=0
cc_1172 N_S[11]_c_1443_n N_A_1361_937#_c_1547_n 0.00343766f $X=6.73 $Y=4.61
+ $X2=0 $Y2=0
cc_1173 N_S[11]_c_1444_n N_A_1361_937#_c_1547_n 0.0164662f $X=7.72 $Y=4.535
+ $X2=0 $Y2=0
cc_1174 S[11] N_A_1361_937#_c_1547_n 0.0178233f $X=6.585 $Y=4.165 $X2=0 $Y2=0
cc_1175 N_S[11]_c_1447_n N_A_1361_937#_c_1548_n 0.00382813f $X=6.73 $Y=4.03
+ $X2=0 $Y2=0
cc_1176 N_S[11]_c_1443_n N_A_1361_937#_c_1548_n 0.00384202f $X=6.73 $Y=4.61
+ $X2=0 $Y2=0
cc_1177 N_S[11]_c_1444_n N_A_1361_937#_c_1548_n 0.00928634f $X=7.72 $Y=4.535
+ $X2=0 $Y2=0
cc_1178 S[11] N_A_1361_937#_c_1548_n 0.0214702f $X=6.585 $Y=4.165 $X2=0 $Y2=0
cc_1179 N_S[11]_c_1447_n N_A_1361_937#_c_1549_n 0.00150889f $X=6.73 $Y=4.03
+ $X2=0 $Y2=0
cc_1180 N_S[11]_c_1443_n N_A_1361_937#_c_1549_n 0.00508702f $X=6.73 $Y=4.61
+ $X2=0 $Y2=0
cc_1181 N_S[11]_c_1444_n N_A_1361_937#_c_1549_n 0.0266986f $X=7.72 $Y=4.535
+ $X2=0 $Y2=0
cc_1182 S[11] N_A_1361_937#_c_1549_n 2.59957e-19 $X=6.585 $Y=4.165 $X2=0 $Y2=0
cc_1183 N_S[11]_c_1443_n N_A_1361_937#_c_1550_n 0.00827389f $X=6.73 $Y=4.61
+ $X2=0 $Y2=0
cc_1184 S[11] N_A_1361_937#_c_1550_n 0.00603567f $X=6.585 $Y=4.165 $X2=0 $Y2=0
cc_1185 N_S[11]_c_1444_n N_D[11]_c_1644_n 0.0286599f $X=7.72 $Y=4.535 $X2=0
+ $Y2=0
cc_1186 N_S[11]_c_1444_n N_D[11]_c_1645_n 0.00289497f $X=7.72 $Y=4.535 $X2=0
+ $Y2=0
cc_1187 N_S[11]_c_1447_n N_VPWR_c_2829_n 0.00965725f $X=6.73 $Y=4.03 $X2=0 $Y2=0
cc_1188 S[11] N_VPWR_c_2829_n 0.00587376f $X=6.585 $Y=4.165 $X2=0 $Y2=0
cc_1189 N_S[11]_c_1447_n VPWR 0.0072999f $X=6.73 $Y=4.03 $X2=0 $Y2=0
cc_1190 N_S[11]_c_1447_n N_VPWR_c_2853_n 0.0035837f $X=6.73 $Y=4.03 $X2=0 $Y2=0
cc_1191 N_S[11]_c_1444_n N_Z_c_3332_n 0.00501353f $X=7.72 $Y=4.535 $X2=0 $Y2=0
cc_1192 N_S[11]_c_1445_n N_Z_c_3332_n 0.00316445f $X=7.795 $Y=4.61 $X2=0 $Y2=0
cc_1193 N_S[11]_c_1444_n N_Z_c_3334_n 7.46972e-19 $X=7.72 $Y=4.535 $X2=0 $Y2=0
cc_1194 N_S[11]_c_1447_n N_Z_c_3406_n 0.00124373f $X=6.73 $Y=4.03 $X2=0 $Y2=0
cc_1195 N_S[11]_c_1444_n N_Z_c_3358_n 0.0141229f $X=7.72 $Y=4.535 $X2=0 $Y2=0
cc_1196 N_S[11]_c_1447_n N_Z_c_3422_n 0.00597491f $X=6.73 $Y=4.03 $X2=0 $Y2=0
cc_1197 N_S[11]_c_1443_n N_Z_c_3422_n 2.32192e-19 $X=6.73 $Y=4.61 $X2=0 $Y2=0
cc_1198 S[11] N_Z_c_3422_n 0.00659242f $X=6.585 $Y=4.165 $X2=0 $Y2=0
cc_1199 N_S[11]_c_1443_n N_VGND_c_4376_n 0.00570474f $X=6.73 $Y=4.61 $X2=0 $Y2=0
cc_1200 S[11] N_VGND_c_4376_n 0.00391126f $X=6.585 $Y=4.165 $X2=0 $Y2=0
cc_1201 N_S[11]_c_1443_n VGND 0.0130664f $X=6.73 $Y=4.61 $X2=0 $Y2=0
cc_1202 N_S[11]_c_1444_n VGND 0.00349917f $X=7.72 $Y=4.535 $X2=0 $Y2=0
cc_1203 N_S[11]_c_1445_n VGND 0.00880034f $X=7.795 $Y=4.61 $X2=0 $Y2=0
cc_1204 N_S[11]_c_1443_n N_VGND_c_4410_n 0.00585385f $X=6.73 $Y=4.61 $X2=0 $Y2=0
cc_1205 N_S[11]_c_1445_n N_VGND_c_4410_n 0.00585385f $X=7.795 $Y=4.61 $X2=0
+ $Y2=0
cc_1206 N_A_1361_47#_M1022_g N_A_1361_937#_M1074_g 0.0129371f $X=7.72 $Y=2.075
+ $X2=0 $Y2=0
cc_1207 N_A_1361_47#_M1022_g N_D[3]_c_1606_n 0.0390641f $X=7.72 $Y=2.075
+ $X2=-0.19 $Y2=-0.24
cc_1208 N_A_1361_47#_c_1492_n N_D[3]_c_1606_n 0.00712672f $X=7.415 $Y=1.34
+ $X2=-0.19 $Y2=-0.24
cc_1209 N_A_1361_47#_c_1495_n N_VPWR_c_2828_n 0.0292866f $X=6.965 $Y=2.31 $X2=0
+ $Y2=0
cc_1210 N_A_1361_47#_c_1491_n N_VPWR_c_2828_n 0.00688579f $X=7.195 $Y=1.405
+ $X2=0 $Y2=0
cc_1211 N_A_1361_47#_M1022_g N_VPWR_c_2830_n 0.00258498f $X=7.72 $Y=2.075 $X2=0
+ $Y2=0
cc_1212 N_A_1361_47#_M1009_d VPWR 0.00179197f $X=6.82 $Y=1.485 $X2=0 $Y2=0
cc_1213 N_A_1361_47#_M1022_g VPWR 0.00387928f $X=7.72 $Y=2.075 $X2=0 $Y2=0
cc_1214 N_A_1361_47#_c_1495_n VPWR 0.00594162f $X=6.965 $Y=2.31 $X2=0 $Y2=0
cc_1215 N_A_1361_47#_c_1495_n N_VPWR_c_2853_n 0.0210596f $X=6.965 $Y=2.31 $X2=0
+ $Y2=0
cc_1216 N_A_1361_47#_M1022_g N_Z_c_3375_n 0.00544362f $X=7.72 $Y=2.075 $X2=0
+ $Y2=0
cc_1217 N_A_1361_47#_c_1495_n N_Z_c_3375_n 0.0371028f $X=6.965 $Y=2.31 $X2=0
+ $Y2=0
cc_1218 N_A_1361_47#_c_1490_n N_Z_c_3331_n 0.00611965f $X=7.195 $Y=1.175 $X2=0
+ $Y2=0
cc_1219 N_A_1361_47#_c_1493_n N_Z_c_3331_n 0.0259454f $X=6.965 $Y=0.495 $X2=0
+ $Y2=0
cc_1220 N_A_1361_47#_M1022_g N_Z_c_3333_n 0.00862328f $X=7.72 $Y=2.075 $X2=0
+ $Y2=0
cc_1221 N_A_1361_47#_c_1495_n N_Z_c_3333_n 0.00378484f $X=6.965 $Y=2.31 $X2=0
+ $Y2=0
cc_1222 N_A_1361_47#_c_1490_n N_Z_c_3333_n 0.00719188f $X=7.195 $Y=1.175 $X2=0
+ $Y2=0
cc_1223 N_A_1361_47#_c_1491_n N_Z_c_3333_n 0.0304368f $X=7.195 $Y=1.405 $X2=0
+ $Y2=0
cc_1224 N_A_1361_47#_c_1492_n N_Z_c_3333_n 0.00814206f $X=7.415 $Y=1.34 $X2=0
+ $Y2=0
cc_1225 N_A_1361_47#_M1022_g N_Z_c_3404_n 0.00335035f $X=7.72 $Y=2.075 $X2=0
+ $Y2=0
cc_1226 N_A_1361_47#_M1022_g N_Z_c_3406_n 0.00502861f $X=7.72 $Y=2.075 $X2=0
+ $Y2=0
cc_1227 N_A_1361_47#_c_1490_n N_Z_c_3357_n 0.0124144f $X=7.195 $Y=1.175 $X2=0
+ $Y2=0
cc_1228 N_A_1361_47#_c_1491_n N_Z_c_3357_n 0.00398133f $X=7.195 $Y=1.405 $X2=0
+ $Y2=0
cc_1229 N_A_1361_47#_c_1492_n N_Z_c_3357_n 0.00349316f $X=7.415 $Y=1.34 $X2=0
+ $Y2=0
cc_1230 N_A_1361_47#_c_1495_n N_Z_c_3421_n 0.0291787f $X=6.965 $Y=2.31 $X2=0
+ $Y2=0
cc_1231 N_A_1361_47#_c_1491_n N_Z_c_3421_n 0.0126642f $X=7.195 $Y=1.405 $X2=0
+ $Y2=0
cc_1232 N_A_1361_47#_M1022_g N_Z_c_3712_n 0.00289142f $X=7.72 $Y=2.075 $X2=0
+ $Y2=0
cc_1233 N_A_1361_47#_c_1495_n N_Z_c_3712_n 6.03258e-19 $X=6.965 $Y=2.31 $X2=0
+ $Y2=0
cc_1234 N_A_1361_47#_c_1491_n N_Z_c_3712_n 4.25753e-19 $X=7.195 $Y=1.405 $X2=0
+ $Y2=0
cc_1235 N_A_1361_47#_M1022_g N_Z_c_3433_n 0.0107335f $X=7.72 $Y=2.075 $X2=0
+ $Y2=0
cc_1236 N_A_1361_47#_c_1495_n N_Z_c_3433_n 0.0139746f $X=6.965 $Y=2.31 $X2=0
+ $Y2=0
cc_1237 N_A_1361_47#_c_1491_n N_Z_c_3433_n 0.00749574f $X=7.195 $Y=1.405 $X2=0
+ $Y2=0
cc_1238 N_A_1361_47#_c_1492_n N_Z_c_3433_n 0.00449418f $X=7.415 $Y=1.34 $X2=0
+ $Y2=0
cc_1239 N_A_1361_47#_M1052_d VGND 0.00358139f $X=6.805 $Y=0.235 $X2=0 $Y2=0
cc_1240 N_A_1361_47#_c_1493_n VGND 0.0150148f $X=6.965 $Y=0.495 $X2=0 $Y2=0
cc_1241 N_A_1361_47#_c_1493_n N_VGND_c_4409_n 0.015238f $X=6.965 $Y=0.495 $X2=0
+ $Y2=0
cc_1242 N_A_1361_937#_M1074_g N_D[11]_c_1647_n 0.0390641f $X=7.72 $Y=3.365
+ $X2=-0.19 $Y2=-0.24
cc_1243 N_A_1361_937#_c_1549_n N_D[11]_c_1647_n 0.00216577f $X=7.415 $Y=4.1
+ $X2=-0.19 $Y2=-0.24
cc_1244 N_A_1361_937#_c_1549_n N_D[11]_c_1644_n 0.00496096f $X=7.415 $Y=4.1
+ $X2=0 $Y2=0
cc_1245 N_A_1361_937#_c_1552_n N_VPWR_c_2829_n 0.0292866f $X=6.965 $Y=3.13 $X2=0
+ $Y2=0
cc_1246 N_A_1361_937#_c_1548_n N_VPWR_c_2829_n 0.00688579f $X=7.195 $Y=4.035
+ $X2=0 $Y2=0
cc_1247 N_A_1361_937#_M1074_g N_VPWR_c_2831_n 0.00258498f $X=7.72 $Y=3.365 $X2=0
+ $Y2=0
cc_1248 N_A_1361_937#_M1012_d VPWR 0.00179197f $X=6.82 $Y=2.955 $X2=0 $Y2=0
cc_1249 N_A_1361_937#_M1074_g VPWR 0.00387928f $X=7.72 $Y=3.365 $X2=0 $Y2=0
cc_1250 N_A_1361_937#_c_1552_n VPWR 0.00594162f $X=6.965 $Y=3.13 $X2=0 $Y2=0
cc_1251 N_A_1361_937#_c_1552_n N_VPWR_c_2853_n 0.0210596f $X=6.965 $Y=3.13 $X2=0
+ $Y2=0
cc_1252 N_A_1361_937#_M1074_g N_Z_c_3376_n 0.00544362f $X=7.72 $Y=3.365 $X2=0
+ $Y2=0
cc_1253 N_A_1361_937#_c_1547_n N_Z_c_3332_n 0.00611965f $X=7.195 $Y=4.685 $X2=0
+ $Y2=0
cc_1254 N_A_1361_937#_c_1550_n N_Z_c_3332_n 0.0259454f $X=6.965 $Y=4.945 $X2=0
+ $Y2=0
cc_1255 N_A_1361_937#_M1074_g N_Z_c_3334_n 0.00862328f $X=7.72 $Y=3.365 $X2=0
+ $Y2=0
cc_1256 N_A_1361_937#_c_1552_n N_Z_c_3334_n 0.00378484f $X=6.965 $Y=3.13 $X2=0
+ $Y2=0
cc_1257 N_A_1361_937#_c_1547_n N_Z_c_3334_n 0.00719188f $X=7.195 $Y=4.685 $X2=0
+ $Y2=0
cc_1258 N_A_1361_937#_c_1548_n N_Z_c_3334_n 0.0304368f $X=7.195 $Y=4.035 $X2=0
+ $Y2=0
cc_1259 N_A_1361_937#_c_1549_n N_Z_c_3334_n 0.00814206f $X=7.415 $Y=4.1 $X2=0
+ $Y2=0
cc_1260 N_A_1361_937#_M1074_g N_Z_c_3405_n 0.00335035f $X=7.72 $Y=3.365 $X2=0
+ $Y2=0
cc_1261 N_A_1361_937#_c_1552_n N_Z_c_3405_n 0.0371028f $X=6.965 $Y=3.13 $X2=0
+ $Y2=0
cc_1262 N_A_1361_937#_M1074_g N_Z_c_3406_n 0.00502861f $X=7.72 $Y=3.365 $X2=0
+ $Y2=0
cc_1263 N_A_1361_937#_c_1547_n N_Z_c_3358_n 0.0124144f $X=7.195 $Y=4.685 $X2=0
+ $Y2=0
cc_1264 N_A_1361_937#_c_1548_n N_Z_c_3358_n 0.00398133f $X=7.195 $Y=4.035 $X2=0
+ $Y2=0
cc_1265 N_A_1361_937#_c_1549_n N_Z_c_3358_n 0.00349316f $X=7.415 $Y=4.1 $X2=0
+ $Y2=0
cc_1266 N_A_1361_937#_c_1552_n N_Z_c_3422_n 0.0291787f $X=6.965 $Y=3.13 $X2=0
+ $Y2=0
cc_1267 N_A_1361_937#_c_1548_n N_Z_c_3422_n 0.0126642f $X=7.195 $Y=4.035 $X2=0
+ $Y2=0
cc_1268 N_A_1361_937#_M1074_g N_Z_c_3735_n 0.00289142f $X=7.72 $Y=3.365 $X2=0
+ $Y2=0
cc_1269 N_A_1361_937#_c_1552_n N_Z_c_3735_n 6.03258e-19 $X=6.965 $Y=3.13 $X2=0
+ $Y2=0
cc_1270 N_A_1361_937#_c_1548_n N_Z_c_3735_n 4.25753e-19 $X=7.195 $Y=4.035 $X2=0
+ $Y2=0
cc_1271 N_A_1361_937#_M1074_g N_Z_c_3434_n 0.0107344f $X=7.72 $Y=3.365 $X2=0
+ $Y2=0
cc_1272 N_A_1361_937#_c_1552_n N_Z_c_3434_n 0.0139746f $X=6.965 $Y=3.13 $X2=0
+ $Y2=0
cc_1273 N_A_1361_937#_c_1548_n N_Z_c_3434_n 0.00749574f $X=7.195 $Y=4.035 $X2=0
+ $Y2=0
cc_1274 N_A_1361_937#_c_1549_n N_Z_c_3434_n 0.00449418f $X=7.415 $Y=4.1 $X2=0
+ $Y2=0
cc_1275 N_A_1361_937#_M1061_d VGND 0.00358139f $X=6.805 $Y=4.685 $X2=0 $Y2=0
cc_1276 N_A_1361_937#_c_1550_n VGND 0.0150148f $X=6.965 $Y=4.945 $X2=0 $Y2=0
cc_1277 N_A_1361_937#_c_1550_n N_VGND_c_4410_n 0.015238f $X=6.965 $Y=4.945 $X2=0
+ $Y2=0
cc_1278 N_D[3]_c_1606_n N_D[11]_c_1647_n 0.0129371f $X=8.245 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_1279 N_D[3]_c_1607_n N_D[4]_c_1685_n 0.00915308f $X=8.27 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_1280 N_D[3]_c_1606_n N_D[4]_c_1686_n 0.0270908f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_1281 N_D[3]_c_1609_n N_D[4]_c_1686_n 9.4377e-19 $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_1282 N_D[3]_c_1608_n N_D[4]_c_1687_n 0.00442615f $X=8.095 $Y=1.055 $X2=0
+ $Y2=0
cc_1283 N_D[3]_c_1606_n N_D[4]_c_1688_n 9.4377e-19 $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_1284 N_D[3]_c_1609_n N_D[4]_c_1688_n 0.0199139f $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_1285 N_D[3]_c_1606_n N_VPWR_c_2830_n 0.0220781f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_1286 N_D[3]_c_1609_n N_VPWR_c_2830_n 0.0044581f $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_1287 N_D[3]_c_1606_n VPWR 0.00468368f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_1288 N_D[3]_c_1606_n N_VPWR_c_2854_n 0.00342413f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_1289 N_D[3]_c_1606_n N_Z_c_3375_n 0.00176496f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_1290 N_D[3]_c_1608_n N_Z_c_3331_n 0.00686805f $X=8.095 $Y=1.055 $X2=0 $Y2=0
cc_1291 N_D[3]_c_1606_n N_Z_c_3333_n 0.00605747f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_1292 N_D[3]_c_1608_n N_Z_c_3333_n 0.00376465f $X=8.095 $Y=1.055 $X2=0 $Y2=0
cc_1293 N_D[3]_c_1609_n N_Z_c_3333_n 0.0216525f $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_1294 N_D[3]_c_1608_n N_Z_c_3357_n 0.0128881f $X=8.095 $Y=1.055 $X2=0 $Y2=0
cc_1295 N_D[3]_c_1606_n N_Z_c_3748_n 0.00719456f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_1296 N_D[3]_c_1609_n N_Z_c_3748_n 0.00989895f $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_1297 N_D[3]_c_1606_n N_Z_c_3433_n 8.42164e-19 $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_1298 N_D[3]_c_1607_n N_VGND_c_4377_n 0.00322791f $X=8.27 $Y=0.995 $X2=0 $Y2=0
cc_1299 N_D[3]_c_1609_n N_VGND_c_4377_n 0.00222881f $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_1300 N_D[3]_c_1607_n VGND 0.0108306f $X=8.27 $Y=0.995 $X2=0 $Y2=0
cc_1301 N_D[3]_c_1639_p VGND 0.00942277f $X=8.095 $Y=0.51 $X2=0 $Y2=0
cc_1302 N_D[3]_c_1607_n N_VGND_c_4409_n 0.00585385f $X=8.27 $Y=0.995 $X2=0 $Y2=0
cc_1303 N_D[3]_c_1639_p N_VGND_c_4409_n 0.00842546f $X=8.095 $Y=0.51 $X2=0 $Y2=0
cc_1304 N_D[3]_c_1608_n A_1574_47# 0.00426617f $X=8.095 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_1305 N_D[3]_c_1639_p A_1574_47# 0.00894235f $X=8.095 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_1306 N_D[11]_c_1644_n N_D[12]_c_1723_n 0.0287172f $X=8.27 $Y=4.445 $X2=-0.19
+ $Y2=-0.24
cc_1307 N_D[11]_c_1646_n N_D[12]_c_1723_n 9.4377e-19 $X=8.24 $Y=4.28 $X2=-0.19
+ $Y2=-0.24
cc_1308 N_D[11]_c_1647_n N_D[12]_c_1727_n 0.00752667f $X=8.245 $Y=4.03 $X2=0
+ $Y2=0
cc_1309 N_D[11]_c_1645_n N_D[12]_c_1724_n 0.00442615f $X=8.095 $Y=4.815 $X2=0
+ $Y2=0
cc_1310 N_D[11]_c_1644_n N_D[12]_c_1725_n 9.4377e-19 $X=8.27 $Y=4.445 $X2=0
+ $Y2=0
cc_1311 N_D[11]_c_1646_n N_D[12]_c_1725_n 0.0199139f $X=8.24 $Y=4.28 $X2=0 $Y2=0
cc_1312 N_D[11]_c_1647_n N_VPWR_c_2831_n 0.0220781f $X=8.245 $Y=4.03 $X2=0 $Y2=0
cc_1313 N_D[11]_c_1646_n N_VPWR_c_2831_n 0.0044581f $X=8.24 $Y=4.28 $X2=0 $Y2=0
cc_1314 N_D[11]_c_1647_n VPWR 0.00468368f $X=8.245 $Y=4.03 $X2=0 $Y2=0
cc_1315 N_D[11]_c_1647_n N_VPWR_c_2854_n 0.00342413f $X=8.245 $Y=4.03 $X2=0
+ $Y2=0
cc_1316 N_D[11]_c_1645_n N_Z_c_3332_n 0.00686805f $X=8.095 $Y=4.815 $X2=0 $Y2=0
cc_1317 N_D[11]_c_1647_n N_Z_c_3334_n 0.00305841f $X=8.245 $Y=4.03 $X2=0 $Y2=0
cc_1318 N_D[11]_c_1644_n N_Z_c_3334_n 0.00299906f $X=8.27 $Y=4.445 $X2=0 $Y2=0
cc_1319 N_D[11]_c_1645_n N_Z_c_3334_n 0.00376465f $X=8.095 $Y=4.815 $X2=0 $Y2=0
cc_1320 N_D[11]_c_1646_n N_Z_c_3334_n 0.0216525f $X=8.24 $Y=4.28 $X2=0 $Y2=0
cc_1321 N_D[11]_c_1647_n N_Z_c_3406_n 0.00176496f $X=8.245 $Y=4.03 $X2=0 $Y2=0
cc_1322 N_D[11]_c_1645_n N_Z_c_3358_n 0.0128881f $X=8.095 $Y=4.815 $X2=0 $Y2=0
cc_1323 N_D[11]_c_1647_n N_Z_c_3758_n 0.0061664f $X=8.245 $Y=4.03 $X2=0 $Y2=0
cc_1324 N_D[11]_c_1644_n N_Z_c_3758_n 0.00102816f $X=8.27 $Y=4.445 $X2=0 $Y2=0
cc_1325 N_D[11]_c_1646_n N_Z_c_3758_n 0.00989895f $X=8.24 $Y=4.28 $X2=0 $Y2=0
cc_1326 N_D[11]_c_1647_n N_Z_c_3434_n 8.42164e-19 $X=8.245 $Y=4.03 $X2=0 $Y2=0
cc_1327 N_D[11]_c_1644_n N_VGND_c_4378_n 0.00322791f $X=8.27 $Y=4.445 $X2=0
+ $Y2=0
cc_1328 N_D[11]_c_1646_n N_VGND_c_4378_n 0.00222881f $X=8.24 $Y=4.28 $X2=0 $Y2=0
cc_1329 N_D[11]_c_1644_n VGND 0.0108306f $X=8.27 $Y=4.445 $X2=0 $Y2=0
cc_1330 N_D[11]_c_1680_p VGND 0.00941728f $X=8.095 $Y=4.93 $X2=0 $Y2=0
cc_1331 N_D[11]_c_1644_n N_VGND_c_4410_n 0.00585385f $X=8.27 $Y=4.445 $X2=0
+ $Y2=0
cc_1332 N_D[11]_c_1680_p N_VGND_c_4410_n 0.00842546f $X=8.095 $Y=4.93 $X2=0
+ $Y2=0
cc_1333 N_D[11]_c_1645_n A_1574_937# 0.00426617f $X=8.095 $Y=4.815 $X2=-0.19
+ $Y2=-0.24
cc_1334 N_D[11]_c_1680_p A_1574_937# 0.00894235f $X=8.095 $Y=4.93 $X2=-0.19
+ $Y2=-0.24
cc_1335 N_D[4]_c_1686_n N_D[12]_c_1727_n 0.0129371f $X=8.775 $Y=1.41 $X2=0 $Y2=0
cc_1336 N_D[4]_c_1686_n N_A_1840_265#_M1014_g 0.0390641f $X=8.775 $Y=1.41 $X2=0
+ $Y2=0
cc_1337 N_D[4]_c_1686_n N_A_1840_265#_c_1767_n 0.00712672f $X=8.775 $Y=1.41
+ $X2=0 $Y2=0
cc_1338 N_D[4]_c_1685_n N_S[4]_c_1878_n 0.0286599f $X=8.75 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_1339 N_D[4]_c_1687_n N_S[4]_c_1878_n 0.00289497f $X=8.925 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_1340 N_D[4]_c_1686_n N_VPWR_c_2830_n 0.0220781f $X=8.775 $Y=1.41 $X2=0 $Y2=0
cc_1341 N_D[4]_c_1688_n N_VPWR_c_2830_n 0.0044581f $X=8.925 $Y=1.19 $X2=0 $Y2=0
cc_1342 N_D[4]_c_1686_n VPWR 0.00468368f $X=8.775 $Y=1.41 $X2=0 $Y2=0
cc_1343 N_D[4]_c_1686_n N_VPWR_c_2855_n 0.00342413f $X=8.775 $Y=1.41 $X2=0 $Y2=0
cc_1344 N_D[4]_c_1686_n N_Z_c_3335_n 0.00605747f $X=8.775 $Y=1.41 $X2=0 $Y2=0
cc_1345 N_D[4]_c_1687_n N_Z_c_3335_n 0.00376465f $X=8.925 $Y=1.055 $X2=0 $Y2=0
cc_1346 N_D[4]_c_1688_n N_Z_c_3335_n 0.0216525f $X=8.925 $Y=1.19 $X2=0 $Y2=0
cc_1347 N_D[4]_c_1687_n N_Z_c_3337_n 0.0128881f $X=8.925 $Y=1.055 $X2=0 $Y2=0
cc_1348 N_D[4]_c_1687_n N_Z_c_3338_n 0.00686805f $X=8.925 $Y=1.055 $X2=0 $Y2=0
cc_1349 N_D[4]_c_1686_n N_Z_c_3381_n 0.00176496f $X=8.775 $Y=1.41 $X2=0 $Y2=0
cc_1350 N_D[4]_c_1686_n N_Z_c_3748_n 0.00719456f $X=8.775 $Y=1.41 $X2=0 $Y2=0
cc_1351 N_D[4]_c_1688_n N_Z_c_3748_n 0.00989895f $X=8.925 $Y=1.19 $X2=0 $Y2=0
cc_1352 N_D[4]_c_1686_n N_Z_c_3435_n 8.42164e-19 $X=8.775 $Y=1.41 $X2=0 $Y2=0
cc_1353 N_D[4]_c_1685_n N_VGND_c_4377_n 0.00322791f $X=8.75 $Y=0.995 $X2=0 $Y2=0
cc_1354 N_D[4]_c_1688_n N_VGND_c_4377_n 0.00222881f $X=8.925 $Y=1.19 $X2=0 $Y2=0
cc_1355 N_D[4]_c_1685_n N_VGND_c_4397_n 0.00585385f $X=8.75 $Y=0.995 $X2=0 $Y2=0
cc_1356 D[4] N_VGND_c_4397_n 0.00842546f $X=8.885 $Y=0.425 $X2=0 $Y2=0
cc_1357 N_D[4]_c_1685_n VGND 0.0108306f $X=8.75 $Y=0.995 $X2=0 $Y2=0
cc_1358 D[4] VGND 0.00942277f $X=8.885 $Y=0.425 $X2=0 $Y2=0
cc_1359 N_D[4]_c_1687_n A_1765_47# 0.00426617f $X=8.925 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_1360 D[4] A_1765_47# 0.00894235f $X=8.885 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_1361 N_D[12]_c_1727_n N_A_1840_793#_M1064_g 0.0390641f $X=8.775 $Y=4.03 $X2=0
+ $Y2=0
cc_1362 N_D[12]_c_1723_n N_A_1840_793#_c_1824_n 0.00496096f $X=8.75 $Y=4.445
+ $X2=0 $Y2=0
cc_1363 N_D[12]_c_1727_n N_A_1840_793#_c_1824_n 0.00216577f $X=8.775 $Y=4.03
+ $X2=0 $Y2=0
cc_1364 N_D[12]_c_1723_n N_S[12]_c_1929_n 0.0286599f $X=8.75 $Y=4.445 $X2=0
+ $Y2=0
cc_1365 N_D[12]_c_1724_n N_S[12]_c_1929_n 0.00289497f $X=8.925 $Y=4.815 $X2=0
+ $Y2=0
cc_1366 N_D[12]_c_1727_n N_VPWR_c_2831_n 0.0220781f $X=8.775 $Y=4.03 $X2=0 $Y2=0
cc_1367 N_D[12]_c_1725_n N_VPWR_c_2831_n 0.0044581f $X=8.925 $Y=4.25 $X2=0 $Y2=0
cc_1368 N_D[12]_c_1727_n VPWR 0.00468368f $X=8.775 $Y=4.03 $X2=0 $Y2=0
cc_1369 N_D[12]_c_1727_n N_VPWR_c_2855_n 0.00342413f $X=8.775 $Y=4.03 $X2=0
+ $Y2=0
cc_1370 N_D[12]_c_1723_n N_Z_c_3336_n 0.00299906f $X=8.75 $Y=4.445 $X2=0 $Y2=0
cc_1371 N_D[12]_c_1727_n N_Z_c_3336_n 0.00305841f $X=8.775 $Y=4.03 $X2=0 $Y2=0
cc_1372 N_D[12]_c_1724_n N_Z_c_3336_n 0.00376465f $X=8.925 $Y=4.815 $X2=0 $Y2=0
cc_1373 N_D[12]_c_1725_n N_Z_c_3336_n 0.0216525f $X=8.925 $Y=4.25 $X2=0 $Y2=0
cc_1374 N_D[12]_c_1724_n N_Z_c_3339_n 0.0128881f $X=8.925 $Y=4.815 $X2=0 $Y2=0
cc_1375 N_D[12]_c_1724_n N_Z_c_3340_n 0.00686805f $X=8.925 $Y=4.815 $X2=0 $Y2=0
cc_1376 N_D[12]_c_1727_n N_Z_c_3409_n 0.00176496f $X=8.775 $Y=4.03 $X2=0 $Y2=0
cc_1377 N_D[12]_c_1723_n N_Z_c_3758_n 0.00102816f $X=8.75 $Y=4.445 $X2=0 $Y2=0
cc_1378 N_D[12]_c_1727_n N_Z_c_3758_n 0.0061664f $X=8.775 $Y=4.03 $X2=0 $Y2=0
cc_1379 N_D[12]_c_1725_n N_Z_c_3758_n 0.00989895f $X=8.925 $Y=4.25 $X2=0 $Y2=0
cc_1380 N_D[12]_c_1727_n N_Z_c_3436_n 8.42164e-19 $X=8.775 $Y=4.03 $X2=0 $Y2=0
cc_1381 N_D[12]_c_1723_n N_VGND_c_4378_n 0.00322791f $X=8.75 $Y=4.445 $X2=0
+ $Y2=0
cc_1382 N_D[12]_c_1725_n N_VGND_c_4378_n 0.00222881f $X=8.925 $Y=4.25 $X2=0
+ $Y2=0
cc_1383 N_D[12]_c_1723_n N_VGND_c_4399_n 0.00585385f $X=8.75 $Y=4.445 $X2=0
+ $Y2=0
cc_1384 D[12] N_VGND_c_4399_n 0.00842546f $X=8.885 $Y=4.845 $X2=0 $Y2=0
cc_1385 N_D[12]_c_1723_n VGND 0.0108306f $X=8.75 $Y=4.445 $X2=0 $Y2=0
cc_1386 D[12] VGND 0.00941728f $X=8.885 $Y=4.845 $X2=0 $Y2=0
cc_1387 N_D[12]_c_1724_n A_1765_911# 0.00426617f $X=8.925 $Y=4.815 $X2=-0.19
+ $Y2=-0.24
cc_1388 D[12] A_1765_911# 0.00894235f $X=8.885 $Y=4.845 $X2=-0.19 $Y2=-0.24
cc_1389 N_A_1840_265#_M1014_g N_A_1840_793#_M1064_g 0.0129371f $X=9.3 $Y=2.075
+ $X2=0 $Y2=0
cc_1390 N_A_1840_265#_c_1764_n N_S[4]_c_1879_n 0.00827389f $X=9.825 $Y=0.755
+ $X2=0 $Y2=0
cc_1391 N_A_1840_265#_c_1765_n N_S[4]_c_1879_n 0.0164662f $X=9.825 $Y=1.175
+ $X2=0 $Y2=0
cc_1392 N_A_1840_265#_c_1766_n N_S[4]_c_1879_n 0.00928634f $X=10.055 $Y=1.63
+ $X2=0 $Y2=0
cc_1393 N_A_1840_265#_c_1767_n N_S[4]_c_1879_n 0.0184911f $X=9.3 $Y=1.34 $X2=0
+ $Y2=0
cc_1394 N_A_1840_265#_c_1767_n N_S[4]_c_1880_n 0.00820745f $X=9.3 $Y=1.34 $X2=0
+ $Y2=0
cc_1395 N_A_1840_265#_c_1765_n N_S[4]_c_1881_n 0.0012443f $X=9.825 $Y=1.175
+ $X2=0 $Y2=0
cc_1396 N_A_1840_265#_c_1769_n N_S[4]_c_1881_n 0.00902681f $X=10.055 $Y=2.31
+ $X2=0 $Y2=0
cc_1397 N_A_1840_265#_c_1766_n N_S[4]_c_1881_n 0.00767015f $X=10.055 $Y=1.63
+ $X2=0 $Y2=0
cc_1398 N_A_1840_265#_c_1767_n N_S[4]_c_1881_n 0.00659591f $X=9.3 $Y=1.34 $X2=0
+ $Y2=0
cc_1399 N_A_1840_265#_c_1765_n N_S[4]_c_1882_n 0.00219336f $X=9.825 $Y=1.175
+ $X2=0 $Y2=0
cc_1400 N_A_1840_265#_c_1764_n N_S[4]_c_1883_n 0.00603567f $X=9.825 $Y=0.755
+ $X2=0 $Y2=0
cc_1401 N_A_1840_265#_c_1765_n N_S[4]_c_1883_n 0.0178233f $X=9.825 $Y=1.175
+ $X2=0 $Y2=0
cc_1402 N_A_1840_265#_c_1766_n N_S[4]_c_1883_n 0.0214702f $X=10.055 $Y=1.63
+ $X2=0 $Y2=0
cc_1403 N_A_1840_265#_c_1767_n N_S[4]_c_1883_n 2.59957e-19 $X=9.3 $Y=1.34 $X2=0
+ $Y2=0
cc_1404 N_A_1840_265#_M1014_g N_VPWR_c_2830_n 0.00258498f $X=9.3 $Y=2.075 $X2=0
+ $Y2=0
cc_1405 N_A_1840_265#_c_1769_n N_VPWR_c_2832_n 0.0292866f $X=10.055 $Y=2.31
+ $X2=0 $Y2=0
cc_1406 N_A_1840_265#_c_1766_n N_VPWR_c_2832_n 0.00688579f $X=10.055 $Y=1.63
+ $X2=0 $Y2=0
cc_1407 N_A_1840_265#_c_1769_n N_VPWR_c_2844_n 0.0210596f $X=10.055 $Y=2.31
+ $X2=0 $Y2=0
cc_1408 N_A_1840_265#_M1080_s VPWR 0.00179197f $X=9.93 $Y=1.485 $X2=0 $Y2=0
cc_1409 N_A_1840_265#_M1014_g VPWR 0.00387928f $X=9.3 $Y=2.075 $X2=0 $Y2=0
cc_1410 N_A_1840_265#_c_1769_n VPWR 0.00594162f $X=10.055 $Y=2.31 $X2=0 $Y2=0
cc_1411 N_A_1840_265#_M1014_g N_Z_c_3335_n 0.00862328f $X=9.3 $Y=2.075 $X2=0
+ $Y2=0
cc_1412 N_A_1840_265#_c_1765_n N_Z_c_3335_n 0.00719188f $X=9.825 $Y=1.175 $X2=0
+ $Y2=0
cc_1413 N_A_1840_265#_c_1769_n N_Z_c_3335_n 0.00378484f $X=10.055 $Y=2.31 $X2=0
+ $Y2=0
cc_1414 N_A_1840_265#_c_1766_n N_Z_c_3335_n 0.0304368f $X=10.055 $Y=1.63 $X2=0
+ $Y2=0
cc_1415 N_A_1840_265#_c_1767_n N_Z_c_3335_n 0.00814206f $X=9.3 $Y=1.34 $X2=0
+ $Y2=0
cc_1416 N_A_1840_265#_c_1765_n N_Z_c_3337_n 0.0124144f $X=9.825 $Y=1.175 $X2=0
+ $Y2=0
cc_1417 N_A_1840_265#_c_1766_n N_Z_c_3337_n 0.00398133f $X=10.055 $Y=1.63 $X2=0
+ $Y2=0
cc_1418 N_A_1840_265#_c_1767_n N_Z_c_3337_n 0.00349316f $X=9.3 $Y=1.34 $X2=0
+ $Y2=0
cc_1419 N_A_1840_265#_c_1764_n N_Z_c_3338_n 0.0259454f $X=9.825 $Y=0.755 $X2=0
+ $Y2=0
cc_1420 N_A_1840_265#_c_1765_n N_Z_c_3338_n 0.00611965f $X=9.825 $Y=1.175 $X2=0
+ $Y2=0
cc_1421 N_A_1840_265#_M1014_g N_Z_c_3381_n 0.00544362f $X=9.3 $Y=2.075 $X2=0
+ $Y2=0
cc_1422 N_A_1840_265#_c_1769_n N_Z_c_3381_n 0.0371028f $X=10.055 $Y=2.31 $X2=0
+ $Y2=0
cc_1423 N_A_1840_265#_M1014_g N_Z_c_3407_n 0.00335035f $X=9.3 $Y=2.075 $X2=0
+ $Y2=0
cc_1424 N_A_1840_265#_M1014_g N_Z_c_3409_n 0.00502861f $X=9.3 $Y=2.075 $X2=0
+ $Y2=0
cc_1425 N_A_1840_265#_c_1769_n N_Z_c_3423_n 0.0291787f $X=10.055 $Y=2.31 $X2=0
+ $Y2=0
cc_1426 N_A_1840_265#_c_1766_n N_Z_c_3423_n 0.0126642f $X=10.055 $Y=1.63 $X2=0
+ $Y2=0
cc_1427 N_A_1840_265#_M1014_g N_Z_c_3798_n 0.00289142f $X=9.3 $Y=2.075 $X2=0
+ $Y2=0
cc_1428 N_A_1840_265#_c_1769_n N_Z_c_3798_n 6.03258e-19 $X=10.055 $Y=2.31 $X2=0
+ $Y2=0
cc_1429 N_A_1840_265#_c_1766_n N_Z_c_3798_n 4.25753e-19 $X=10.055 $Y=1.63 $X2=0
+ $Y2=0
cc_1430 N_A_1840_265#_M1014_g N_Z_c_3435_n 0.0107335f $X=9.3 $Y=2.075 $X2=0
+ $Y2=0
cc_1431 N_A_1840_265#_c_1769_n N_Z_c_3435_n 0.0139746f $X=10.055 $Y=2.31 $X2=0
+ $Y2=0
cc_1432 N_A_1840_265#_c_1766_n N_Z_c_3435_n 0.00749574f $X=10.055 $Y=1.63 $X2=0
+ $Y2=0
cc_1433 N_A_1840_265#_c_1767_n N_Z_c_3435_n 0.00449418f $X=9.3 $Y=1.34 $X2=0
+ $Y2=0
cc_1434 N_A_1840_265#_c_1764_n N_VGND_c_4397_n 0.015238f $X=9.825 $Y=0.755 $X2=0
+ $Y2=0
cc_1435 N_A_1840_265#_M1094_s VGND 0.00358139f $X=9.93 $Y=0.235 $X2=0 $Y2=0
cc_1436 N_A_1840_265#_c_1764_n VGND 0.0150148f $X=9.825 $Y=0.755 $X2=0 $Y2=0
cc_1437 N_A_1840_793#_c_1822_n N_S[12]_c_1928_n 0.0247401f $X=9.825 $Y=4.685
+ $X2=0 $Y2=0
cc_1438 N_A_1840_793#_c_1823_n N_S[12]_c_1928_n 0.00928634f $X=10.055 $Y=3.805
+ $X2=0 $Y2=0
cc_1439 N_A_1840_793#_c_1824_n N_S[12]_c_1928_n 0.0184911f $X=9.3 $Y=4.1 $X2=0
+ $Y2=0
cc_1440 N_A_1840_793#_c_1824_n N_S[12]_c_1929_n 0.00820745f $X=9.3 $Y=4.1 $X2=0
+ $Y2=0
cc_1441 N_A_1840_793#_c_1823_n N_S[12]_c_1932_n 0.00382813f $X=10.055 $Y=3.805
+ $X2=0 $Y2=0
cc_1442 N_A_1840_793#_c_1827_n N_S[12]_c_1932_n 0.00902681f $X=10.055 $Y=3.13
+ $X2=0 $Y2=0
cc_1443 N_A_1840_793#_c_1824_n N_S[12]_c_1932_n 0.00150889f $X=9.3 $Y=4.1 $X2=0
+ $Y2=0
cc_1444 N_A_1840_793#_c_1822_n N_S[12]_c_1930_n 0.00343766f $X=9.825 $Y=4.685
+ $X2=0 $Y2=0
cc_1445 N_A_1840_793#_c_1823_n N_S[12]_c_1930_n 0.00384202f $X=10.055 $Y=3.805
+ $X2=0 $Y2=0
cc_1446 N_A_1840_793#_c_1824_n N_S[12]_c_1930_n 0.00508702f $X=9.3 $Y=4.1 $X2=0
+ $Y2=0
cc_1447 N_A_1840_793#_c_1822_n S[12] 0.023859f $X=9.825 $Y=4.685 $X2=0 $Y2=0
cc_1448 N_A_1840_793#_c_1823_n S[12] 0.0214702f $X=10.055 $Y=3.805 $X2=0 $Y2=0
cc_1449 N_A_1840_793#_c_1824_n S[12] 2.59957e-19 $X=9.3 $Y=4.1 $X2=0 $Y2=0
cc_1450 N_A_1840_793#_M1064_g N_VPWR_c_2831_n 0.00258498f $X=9.3 $Y=3.365 $X2=0
+ $Y2=0
cc_1451 N_A_1840_793#_c_1823_n N_VPWR_c_2833_n 0.00688579f $X=10.055 $Y=3.805
+ $X2=0 $Y2=0
cc_1452 N_A_1840_793#_c_1827_n N_VPWR_c_2833_n 0.0292866f $X=10.055 $Y=3.13
+ $X2=0 $Y2=0
cc_1453 N_A_1840_793#_c_1827_n N_VPWR_c_2844_n 0.0210596f $X=10.055 $Y=3.13
+ $X2=0 $Y2=0
cc_1454 N_A_1840_793#_M1085_s VPWR 0.00179197f $X=9.93 $Y=2.955 $X2=0 $Y2=0
cc_1455 N_A_1840_793#_M1064_g VPWR 0.00387928f $X=9.3 $Y=3.365 $X2=0 $Y2=0
cc_1456 N_A_1840_793#_c_1827_n VPWR 0.00594162f $X=10.055 $Y=3.13 $X2=0 $Y2=0
cc_1457 N_A_1840_793#_M1064_g N_Z_c_3336_n 0.00862328f $X=9.3 $Y=3.365 $X2=0
+ $Y2=0
cc_1458 N_A_1840_793#_c_1822_n N_Z_c_3336_n 0.00719188f $X=9.825 $Y=4.685 $X2=0
+ $Y2=0
cc_1459 N_A_1840_793#_c_1823_n N_Z_c_3336_n 0.0304368f $X=10.055 $Y=3.805 $X2=0
+ $Y2=0
cc_1460 N_A_1840_793#_c_1827_n N_Z_c_3336_n 0.00378484f $X=10.055 $Y=3.13 $X2=0
+ $Y2=0
cc_1461 N_A_1840_793#_c_1824_n N_Z_c_3336_n 0.00814206f $X=9.3 $Y=4.1 $X2=0
+ $Y2=0
cc_1462 N_A_1840_793#_c_1822_n N_Z_c_3339_n 0.0124144f $X=9.825 $Y=4.685 $X2=0
+ $Y2=0
cc_1463 N_A_1840_793#_c_1823_n N_Z_c_3339_n 0.00398133f $X=10.055 $Y=3.805 $X2=0
+ $Y2=0
cc_1464 N_A_1840_793#_c_1824_n N_Z_c_3339_n 0.00349316f $X=9.3 $Y=4.1 $X2=0
+ $Y2=0
cc_1465 N_A_1840_793#_c_1822_n N_Z_c_3340_n 0.032065f $X=9.825 $Y=4.685 $X2=0
+ $Y2=0
cc_1466 N_A_1840_793#_M1064_g N_Z_c_3382_n 0.00544362f $X=9.3 $Y=3.365 $X2=0
+ $Y2=0
cc_1467 N_A_1840_793#_M1064_g N_Z_c_3408_n 0.00335035f $X=9.3 $Y=3.365 $X2=0
+ $Y2=0
cc_1468 N_A_1840_793#_c_1827_n N_Z_c_3408_n 0.0371028f $X=10.055 $Y=3.13 $X2=0
+ $Y2=0
cc_1469 N_A_1840_793#_M1064_g N_Z_c_3409_n 0.00502861f $X=9.3 $Y=3.365 $X2=0
+ $Y2=0
cc_1470 N_A_1840_793#_c_1823_n N_Z_c_3424_n 0.0126642f $X=10.055 $Y=3.805 $X2=0
+ $Y2=0
cc_1471 N_A_1840_793#_c_1827_n N_Z_c_3424_n 0.0291787f $X=10.055 $Y=3.13 $X2=0
+ $Y2=0
cc_1472 N_A_1840_793#_M1064_g N_Z_c_3820_n 0.00289142f $X=9.3 $Y=3.365 $X2=0
+ $Y2=0
cc_1473 N_A_1840_793#_c_1823_n N_Z_c_3820_n 4.25753e-19 $X=10.055 $Y=3.805 $X2=0
+ $Y2=0
cc_1474 N_A_1840_793#_c_1827_n N_Z_c_3820_n 6.03258e-19 $X=10.055 $Y=3.13 $X2=0
+ $Y2=0
cc_1475 N_A_1840_793#_M1064_g N_Z_c_3436_n 0.0107344f $X=9.3 $Y=3.365 $X2=0
+ $Y2=0
cc_1476 N_A_1840_793#_c_1823_n N_Z_c_3436_n 0.00749574f $X=10.055 $Y=3.805 $X2=0
+ $Y2=0
cc_1477 N_A_1840_793#_c_1827_n N_Z_c_3436_n 0.0139746f $X=10.055 $Y=3.13 $X2=0
+ $Y2=0
cc_1478 N_A_1840_793#_c_1824_n N_Z_c_3436_n 0.00449418f $X=9.3 $Y=4.1 $X2=0
+ $Y2=0
cc_1479 N_A_1840_793#_c_1822_n N_VGND_c_4399_n 0.015238f $X=9.825 $Y=4.685 $X2=0
+ $Y2=0
cc_1480 N_A_1840_793#_M1024_s VGND 0.00358139f $X=9.93 $Y=4.685 $X2=0 $Y2=0
cc_1481 N_A_1840_793#_c_1822_n VGND 0.0150148f $X=9.825 $Y=4.685 $X2=0 $Y2=0
cc_1482 N_S[4]_c_1881_n N_S[12]_c_1932_n 0.0130744f $X=10.29 $Y=1.41 $X2=0 $Y2=0
cc_1483 N_S[4]_c_1881_n N_S[5]_c_1975_n 0.0578733f $X=10.29 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_1484 N_S[4]_c_1883_n N_S[5]_c_1975_n 0.00112057f $X=10.255 $Y=1.03 $X2=-0.19
+ $Y2=-0.24
cc_1485 N_S[4]_c_1882_n N_S[5]_c_1976_n 0.0091402f $X=10.29 $Y=0.83 $X2=0 $Y2=0
cc_1486 N_S[4]_c_1881_n N_S[5]_c_1979_n 0.00112057f $X=10.29 $Y=1.41 $X2=0 $Y2=0
cc_1487 N_S[4]_c_1883_n N_S[5]_c_1979_n 0.0277403f $X=10.255 $Y=1.03 $X2=0 $Y2=0
cc_1488 N_S[4]_c_1881_n N_VPWR_c_2832_n 0.00965725f $X=10.29 $Y=1.41 $X2=0 $Y2=0
cc_1489 N_S[4]_c_1883_n N_VPWR_c_2832_n 0.00587376f $X=10.255 $Y=1.03 $X2=0
+ $Y2=0
cc_1490 N_S[4]_c_1881_n N_VPWR_c_2844_n 0.0035837f $X=10.29 $Y=1.41 $X2=0 $Y2=0
cc_1491 N_S[4]_c_1881_n VPWR 0.0072999f $X=10.29 $Y=1.41 $X2=0 $Y2=0
cc_1492 N_S[4]_c_1880_n N_Z_c_3335_n 7.46972e-19 $X=9.3 $Y=0.905 $X2=0 $Y2=0
cc_1493 N_S[4]_c_1879_n N_Z_c_3337_n 0.00806549f $X=10.12 $Y=0.905 $X2=0 $Y2=0
cc_1494 N_S[4]_c_1880_n N_Z_c_3337_n 0.00605736f $X=9.3 $Y=0.905 $X2=0 $Y2=0
cc_1495 N_S[4]_c_1878_n N_Z_c_3338_n 0.00316445f $X=9.225 $Y=0.83 $X2=0 $Y2=0
cc_1496 N_S[4]_c_1879_n N_Z_c_3338_n 0.00501353f $X=10.12 $Y=0.905 $X2=0 $Y2=0
cc_1497 N_S[4]_c_1881_n N_Z_c_3409_n 0.00124373f $X=10.29 $Y=1.41 $X2=0 $Y2=0
cc_1498 N_S[4]_c_1881_n N_Z_c_3423_n 0.0062071f $X=10.29 $Y=1.41 $X2=0 $Y2=0
cc_1499 N_S[4]_c_1883_n N_Z_c_3423_n 0.00659242f $X=10.255 $Y=1.03 $X2=0 $Y2=0
cc_1500 N_S[4]_c_1882_n N_VGND_c_4379_n 0.00570474f $X=10.29 $Y=0.83 $X2=0 $Y2=0
cc_1501 N_S[4]_c_1883_n N_VGND_c_4379_n 0.00391126f $X=10.255 $Y=1.03 $X2=0
+ $Y2=0
cc_1502 N_S[4]_c_1878_n N_VGND_c_4397_n 0.00585385f $X=9.225 $Y=0.83 $X2=0 $Y2=0
cc_1503 N_S[4]_c_1882_n N_VGND_c_4397_n 0.00585385f $X=10.29 $Y=0.83 $X2=0 $Y2=0
cc_1504 N_S[4]_c_1878_n VGND 0.00880034f $X=9.225 $Y=0.83 $X2=0 $Y2=0
cc_1505 N_S[4]_c_1879_n VGND 0.00349917f $X=10.12 $Y=0.905 $X2=0 $Y2=0
cc_1506 N_S[4]_c_1881_n VGND 6.15795e-19 $X=10.29 $Y=1.41 $X2=0 $Y2=0
cc_1507 N_S[4]_c_1882_n VGND 0.0124506f $X=10.29 $Y=0.83 $X2=0 $Y2=0
cc_1508 N_S[12]_c_1932_n N_S[13]_c_2025_n 0.0296874f $X=10.29 $Y=4.03 $X2=-0.19
+ $Y2=-0.24
cc_1509 N_S[12]_c_1930_n N_S[13]_c_2021_n 0.0373261f $X=10.29 $Y=4.61 $X2=0
+ $Y2=0
cc_1510 S[12] N_S[13]_c_2021_n 0.00112057f $X=10.265 $Y=4.165 $X2=0 $Y2=0
cc_1511 N_S[12]_c_1930_n S[13] 0.00112057f $X=10.29 $Y=4.61 $X2=0 $Y2=0
cc_1512 S[12] S[13] 0.0277403f $X=10.265 $Y=4.165 $X2=0 $Y2=0
cc_1513 N_S[12]_c_1932_n N_VPWR_c_2833_n 0.00965725f $X=10.29 $Y=4.03 $X2=0
+ $Y2=0
cc_1514 S[12] N_VPWR_c_2833_n 0.00587376f $X=10.265 $Y=4.165 $X2=0 $Y2=0
cc_1515 N_S[12]_c_1932_n N_VPWR_c_2844_n 0.0035837f $X=10.29 $Y=4.03 $X2=0 $Y2=0
cc_1516 N_S[12]_c_1932_n VPWR 0.0072999f $X=10.29 $Y=4.03 $X2=0 $Y2=0
cc_1517 N_S[12]_c_1929_n N_Z_c_3336_n 7.46972e-19 $X=9.3 $Y=4.535 $X2=0 $Y2=0
cc_1518 N_S[12]_c_1928_n N_Z_c_3339_n 0.00806549f $X=10.12 $Y=4.535 $X2=0 $Y2=0
cc_1519 N_S[12]_c_1929_n N_Z_c_3339_n 0.00605736f $X=9.3 $Y=4.535 $X2=0 $Y2=0
cc_1520 N_S[12]_c_1927_n N_Z_c_3340_n 0.00316445f $X=9.225 $Y=4.61 $X2=0 $Y2=0
cc_1521 N_S[12]_c_1928_n N_Z_c_3340_n 0.00501353f $X=10.12 $Y=4.535 $X2=0 $Y2=0
cc_1522 N_S[12]_c_1932_n N_Z_c_3409_n 0.00124373f $X=10.29 $Y=4.03 $X2=0 $Y2=0
cc_1523 N_S[12]_c_1932_n N_Z_c_3424_n 0.00597491f $X=10.29 $Y=4.03 $X2=0 $Y2=0
cc_1524 N_S[12]_c_1930_n N_Z_c_3424_n 2.32192e-19 $X=10.29 $Y=4.61 $X2=0 $Y2=0
cc_1525 S[12] N_Z_c_3424_n 0.00659242f $X=10.265 $Y=4.165 $X2=0 $Y2=0
cc_1526 N_S[12]_c_1930_n N_VGND_c_4380_n 0.00570474f $X=10.29 $Y=4.61 $X2=0
+ $Y2=0
cc_1527 S[12] N_VGND_c_4380_n 0.00391126f $X=10.265 $Y=4.165 $X2=0 $Y2=0
cc_1528 N_S[12]_c_1927_n N_VGND_c_4399_n 0.00585385f $X=9.225 $Y=4.61 $X2=0
+ $Y2=0
cc_1529 N_S[12]_c_1930_n N_VGND_c_4399_n 0.00585385f $X=10.29 $Y=4.61 $X2=0
+ $Y2=0
cc_1530 N_S[12]_c_1927_n VGND 0.00880034f $X=9.225 $Y=4.61 $X2=0 $Y2=0
cc_1531 N_S[12]_c_1928_n VGND 0.00349917f $X=10.12 $Y=4.535 $X2=0 $Y2=0
cc_1532 N_S[12]_c_1930_n VGND 0.0130664f $X=10.29 $Y=4.61 $X2=0 $Y2=0
cc_1533 N_S[5]_c_1975_n N_S[13]_c_2025_n 0.0130744f $X=10.87 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_1534 N_S[5]_c_1975_n N_A_2189_47#_c_2073_n 0.00902681f $X=10.87 $Y=1.41 $X2=0
+ $Y2=0
cc_1535 N_S[5]_c_1975_n N_A_2189_47#_c_2068_n 0.0012443f $X=10.87 $Y=1.41 $X2=0
+ $Y2=0
cc_1536 N_S[5]_c_1976_n N_A_2189_47#_c_2068_n 0.00219336f $X=10.87 $Y=0.83 $X2=0
+ $Y2=0
cc_1537 N_S[5]_c_1977_n N_A_2189_47#_c_2068_n 0.0164662f $X=11.86 $Y=0.905 $X2=0
+ $Y2=0
cc_1538 N_S[5]_c_1979_n N_A_2189_47#_c_2068_n 0.0178233f $X=10.905 $Y=1.03 $X2=0
+ $Y2=0
cc_1539 N_S[5]_c_1975_n N_A_2189_47#_c_2069_n 0.00767015f $X=10.87 $Y=1.41 $X2=0
+ $Y2=0
cc_1540 N_S[5]_c_1977_n N_A_2189_47#_c_2069_n 0.00928634f $X=11.86 $Y=0.905
+ $X2=0 $Y2=0
cc_1541 N_S[5]_c_1979_n N_A_2189_47#_c_2069_n 0.0214702f $X=10.905 $Y=1.03 $X2=0
+ $Y2=0
cc_1542 N_S[5]_c_1975_n N_A_2189_47#_c_2070_n 0.00659591f $X=10.87 $Y=1.41 $X2=0
+ $Y2=0
cc_1543 N_S[5]_c_1977_n N_A_2189_47#_c_2070_n 0.0266986f $X=11.86 $Y=0.905 $X2=0
+ $Y2=0
cc_1544 N_S[5]_c_1979_n N_A_2189_47#_c_2070_n 2.59957e-19 $X=10.905 $Y=1.03
+ $X2=0 $Y2=0
cc_1545 N_S[5]_c_1975_n N_A_2189_47#_c_2071_n 0.00827389f $X=10.87 $Y=1.41 $X2=0
+ $Y2=0
cc_1546 N_S[5]_c_1979_n N_A_2189_47#_c_2071_n 0.00603567f $X=10.905 $Y=1.03
+ $X2=0 $Y2=0
cc_1547 N_S[5]_c_1978_n N_D[5]_c_2185_n 0.0286599f $X=11.935 $Y=0.83 $X2=0 $Y2=0
cc_1548 N_S[5]_c_1978_n N_D[5]_c_2186_n 0.00289497f $X=11.935 $Y=0.83 $X2=0
+ $Y2=0
cc_1549 N_S[5]_c_1975_n N_VPWR_c_2832_n 0.00965725f $X=10.87 $Y=1.41 $X2=0 $Y2=0
cc_1550 N_S[5]_c_1979_n N_VPWR_c_2832_n 0.00587376f $X=10.905 $Y=1.03 $X2=0
+ $Y2=0
cc_1551 N_S[5]_c_1975_n VPWR 0.0072999f $X=10.87 $Y=1.41 $X2=0 $Y2=0
cc_1552 N_S[5]_c_1975_n N_VPWR_c_2856_n 0.0035837f $X=10.87 $Y=1.41 $X2=0 $Y2=0
cc_1553 N_S[5]_c_1977_n N_Z_c_3341_n 0.00501353f $X=11.86 $Y=0.905 $X2=0 $Y2=0
cc_1554 N_S[5]_c_1978_n N_Z_c_3341_n 0.00316445f $X=11.935 $Y=0.83 $X2=0 $Y2=0
cc_1555 N_S[5]_c_1977_n N_Z_c_3343_n 7.46972e-19 $X=11.86 $Y=0.905 $X2=0 $Y2=0
cc_1556 N_S[5]_c_1975_n N_Z_c_3412_n 0.00124373f $X=10.87 $Y=1.41 $X2=0 $Y2=0
cc_1557 N_S[5]_c_1977_n N_Z_c_3359_n 0.0141229f $X=11.86 $Y=0.905 $X2=0 $Y2=0
cc_1558 N_S[5]_c_1975_n N_Z_c_3423_n 0.0062071f $X=10.87 $Y=1.41 $X2=0 $Y2=0
cc_1559 N_S[5]_c_1979_n N_Z_c_3423_n 0.00659242f $X=10.905 $Y=1.03 $X2=0 $Y2=0
cc_1560 N_S[5]_c_1976_n N_VGND_c_4379_n 0.00570474f $X=10.87 $Y=0.83 $X2=0 $Y2=0
cc_1561 N_S[5]_c_1979_n N_VGND_c_4379_n 0.00391126f $X=10.905 $Y=1.03 $X2=0
+ $Y2=0
cc_1562 N_S[5]_c_1975_n VGND 6.15795e-19 $X=10.87 $Y=1.41 $X2=0 $Y2=0
cc_1563 N_S[5]_c_1976_n VGND 0.0124506f $X=10.87 $Y=0.83 $X2=0 $Y2=0
cc_1564 N_S[5]_c_1977_n VGND 0.00349917f $X=11.86 $Y=0.905 $X2=0 $Y2=0
cc_1565 N_S[5]_c_1978_n VGND 0.00880034f $X=11.935 $Y=0.83 $X2=0 $Y2=0
cc_1566 N_S[5]_c_1976_n N_VGND_c_4411_n 0.00585385f $X=10.87 $Y=0.83 $X2=0 $Y2=0
cc_1567 N_S[5]_c_1978_n N_VGND_c_4411_n 0.00585385f $X=11.935 $Y=0.83 $X2=0
+ $Y2=0
cc_1568 N_S[13]_c_2025_n N_A_2189_937#_c_2130_n 0.00902681f $X=10.87 $Y=4.03
+ $X2=0 $Y2=0
cc_1569 N_S[13]_c_2021_n N_A_2189_937#_c_2125_n 0.00343766f $X=10.87 $Y=4.61
+ $X2=0 $Y2=0
cc_1570 N_S[13]_c_2022_n N_A_2189_937#_c_2125_n 0.0164662f $X=11.86 $Y=4.535
+ $X2=0 $Y2=0
cc_1571 S[13] N_A_2189_937#_c_2125_n 0.0178233f $X=10.725 $Y=4.165 $X2=0 $Y2=0
cc_1572 N_S[13]_c_2025_n N_A_2189_937#_c_2126_n 0.00382813f $X=10.87 $Y=4.03
+ $X2=0 $Y2=0
cc_1573 N_S[13]_c_2021_n N_A_2189_937#_c_2126_n 0.00384202f $X=10.87 $Y=4.61
+ $X2=0 $Y2=0
cc_1574 N_S[13]_c_2022_n N_A_2189_937#_c_2126_n 0.00928634f $X=11.86 $Y=4.535
+ $X2=0 $Y2=0
cc_1575 S[13] N_A_2189_937#_c_2126_n 0.0214702f $X=10.725 $Y=4.165 $X2=0 $Y2=0
cc_1576 N_S[13]_c_2025_n N_A_2189_937#_c_2127_n 0.00150889f $X=10.87 $Y=4.03
+ $X2=0 $Y2=0
cc_1577 N_S[13]_c_2021_n N_A_2189_937#_c_2127_n 0.00508702f $X=10.87 $Y=4.61
+ $X2=0 $Y2=0
cc_1578 N_S[13]_c_2022_n N_A_2189_937#_c_2127_n 0.0266986f $X=11.86 $Y=4.535
+ $X2=0 $Y2=0
cc_1579 S[13] N_A_2189_937#_c_2127_n 2.59957e-19 $X=10.725 $Y=4.165 $X2=0 $Y2=0
cc_1580 N_S[13]_c_2021_n N_A_2189_937#_c_2128_n 0.00827389f $X=10.87 $Y=4.61
+ $X2=0 $Y2=0
cc_1581 S[13] N_A_2189_937#_c_2128_n 0.00603567f $X=10.725 $Y=4.165 $X2=0 $Y2=0
cc_1582 N_S[13]_c_2022_n N_D[13]_c_2222_n 0.0286599f $X=11.86 $Y=4.535 $X2=0
+ $Y2=0
cc_1583 N_S[13]_c_2022_n N_D[13]_c_2223_n 0.00289497f $X=11.86 $Y=4.535 $X2=0
+ $Y2=0
cc_1584 N_S[13]_c_2025_n N_VPWR_c_2833_n 0.00965725f $X=10.87 $Y=4.03 $X2=0
+ $Y2=0
cc_1585 S[13] N_VPWR_c_2833_n 0.00587376f $X=10.725 $Y=4.165 $X2=0 $Y2=0
cc_1586 N_S[13]_c_2025_n VPWR 0.0072999f $X=10.87 $Y=4.03 $X2=0 $Y2=0
cc_1587 N_S[13]_c_2025_n N_VPWR_c_2856_n 0.0035837f $X=10.87 $Y=4.03 $X2=0 $Y2=0
cc_1588 N_S[13]_c_2022_n N_Z_c_3342_n 0.00501353f $X=11.86 $Y=4.535 $X2=0 $Y2=0
cc_1589 N_S[13]_c_2023_n N_Z_c_3342_n 0.00316445f $X=11.935 $Y=4.61 $X2=0 $Y2=0
cc_1590 N_S[13]_c_2022_n N_Z_c_3344_n 7.46972e-19 $X=11.86 $Y=4.535 $X2=0 $Y2=0
cc_1591 N_S[13]_c_2025_n N_Z_c_3412_n 0.00124373f $X=10.87 $Y=4.03 $X2=0 $Y2=0
cc_1592 N_S[13]_c_2022_n N_Z_c_3360_n 0.0141229f $X=11.86 $Y=4.535 $X2=0 $Y2=0
cc_1593 N_S[13]_c_2025_n N_Z_c_3424_n 0.00597491f $X=10.87 $Y=4.03 $X2=0 $Y2=0
cc_1594 N_S[13]_c_2021_n N_Z_c_3424_n 2.32192e-19 $X=10.87 $Y=4.61 $X2=0 $Y2=0
cc_1595 S[13] N_Z_c_3424_n 0.00659242f $X=10.725 $Y=4.165 $X2=0 $Y2=0
cc_1596 N_S[13]_c_2021_n N_VGND_c_4380_n 0.00570474f $X=10.87 $Y=4.61 $X2=0
+ $Y2=0
cc_1597 S[13] N_VGND_c_4380_n 0.00391126f $X=10.725 $Y=4.165 $X2=0 $Y2=0
cc_1598 N_S[13]_c_2021_n VGND 0.0130664f $X=10.87 $Y=4.61 $X2=0 $Y2=0
cc_1599 N_S[13]_c_2022_n VGND 0.00349917f $X=11.86 $Y=4.535 $X2=0 $Y2=0
cc_1600 N_S[13]_c_2023_n VGND 0.00880034f $X=11.935 $Y=4.61 $X2=0 $Y2=0
cc_1601 N_S[13]_c_2021_n N_VGND_c_4412_n 0.00585385f $X=10.87 $Y=4.61 $X2=0
+ $Y2=0
cc_1602 N_S[13]_c_2023_n N_VGND_c_4412_n 0.00585385f $X=11.935 $Y=4.61 $X2=0
+ $Y2=0
cc_1603 N_A_2189_47#_M1059_g N_A_2189_937#_M1008_g 0.0129371f $X=11.86 $Y=2.075
+ $X2=0 $Y2=0
cc_1604 N_A_2189_47#_M1059_g N_D[5]_c_2184_n 0.0390641f $X=11.86 $Y=2.075
+ $X2=-0.19 $Y2=-0.24
cc_1605 N_A_2189_47#_c_2070_n N_D[5]_c_2184_n 0.00712672f $X=11.555 $Y=1.34
+ $X2=-0.19 $Y2=-0.24
cc_1606 N_A_2189_47#_c_2073_n N_VPWR_c_2832_n 0.0292866f $X=11.105 $Y=2.31 $X2=0
+ $Y2=0
cc_1607 N_A_2189_47#_c_2069_n N_VPWR_c_2832_n 0.00688579f $X=11.335 $Y=1.405
+ $X2=0 $Y2=0
cc_1608 N_A_2189_47#_M1059_g N_VPWR_c_2834_n 0.00258498f $X=11.86 $Y=2.075 $X2=0
+ $Y2=0
cc_1609 N_A_2189_47#_M1046_d VPWR 0.00179197f $X=10.96 $Y=1.485 $X2=0 $Y2=0
cc_1610 N_A_2189_47#_M1059_g VPWR 0.00387928f $X=11.86 $Y=2.075 $X2=0 $Y2=0
cc_1611 N_A_2189_47#_c_2073_n VPWR 0.00594162f $X=11.105 $Y=2.31 $X2=0 $Y2=0
cc_1612 N_A_2189_47#_c_2073_n N_VPWR_c_2856_n 0.0210596f $X=11.105 $Y=2.31 $X2=0
+ $Y2=0
cc_1613 N_A_2189_47#_M1059_g N_Z_c_3383_n 0.00544362f $X=11.86 $Y=2.075 $X2=0
+ $Y2=0
cc_1614 N_A_2189_47#_c_2073_n N_Z_c_3383_n 0.0371028f $X=11.105 $Y=2.31 $X2=0
+ $Y2=0
cc_1615 N_A_2189_47#_c_2068_n N_Z_c_3341_n 0.00611965f $X=11.335 $Y=1.175 $X2=0
+ $Y2=0
cc_1616 N_A_2189_47#_c_2071_n N_Z_c_3341_n 0.0259454f $X=11.105 $Y=0.495 $X2=0
+ $Y2=0
cc_1617 N_A_2189_47#_M1059_g N_Z_c_3343_n 0.00862328f $X=11.86 $Y=2.075 $X2=0
+ $Y2=0
cc_1618 N_A_2189_47#_c_2073_n N_Z_c_3343_n 0.00378484f $X=11.105 $Y=2.31 $X2=0
+ $Y2=0
cc_1619 N_A_2189_47#_c_2068_n N_Z_c_3343_n 0.00719188f $X=11.335 $Y=1.175 $X2=0
+ $Y2=0
cc_1620 N_A_2189_47#_c_2069_n N_Z_c_3343_n 0.0304368f $X=11.335 $Y=1.405 $X2=0
+ $Y2=0
cc_1621 N_A_2189_47#_c_2070_n N_Z_c_3343_n 0.00814206f $X=11.555 $Y=1.34 $X2=0
+ $Y2=0
cc_1622 N_A_2189_47#_M1059_g N_Z_c_3410_n 0.00335035f $X=11.86 $Y=2.075 $X2=0
+ $Y2=0
cc_1623 N_A_2189_47#_M1059_g N_Z_c_3412_n 0.00502861f $X=11.86 $Y=2.075 $X2=0
+ $Y2=0
cc_1624 N_A_2189_47#_c_2068_n N_Z_c_3359_n 0.0124144f $X=11.335 $Y=1.175 $X2=0
+ $Y2=0
cc_1625 N_A_2189_47#_c_2069_n N_Z_c_3359_n 0.00398133f $X=11.335 $Y=1.405 $X2=0
+ $Y2=0
cc_1626 N_A_2189_47#_c_2070_n N_Z_c_3359_n 0.00349316f $X=11.555 $Y=1.34 $X2=0
+ $Y2=0
cc_1627 N_A_2189_47#_c_2073_n N_Z_c_3423_n 0.0291787f $X=11.105 $Y=2.31 $X2=0
+ $Y2=0
cc_1628 N_A_2189_47#_c_2069_n N_Z_c_3423_n 0.0126642f $X=11.335 $Y=1.405 $X2=0
+ $Y2=0
cc_1629 N_A_2189_47#_M1059_g N_Z_c_3875_n 0.00289142f $X=11.86 $Y=2.075 $X2=0
+ $Y2=0
cc_1630 N_A_2189_47#_c_2073_n N_Z_c_3875_n 6.03258e-19 $X=11.105 $Y=2.31 $X2=0
+ $Y2=0
cc_1631 N_A_2189_47#_c_2069_n N_Z_c_3875_n 4.25753e-19 $X=11.335 $Y=1.405 $X2=0
+ $Y2=0
cc_1632 N_A_2189_47#_M1059_g N_Z_c_3437_n 0.0107335f $X=11.86 $Y=2.075 $X2=0
+ $Y2=0
cc_1633 N_A_2189_47#_c_2073_n N_Z_c_3437_n 0.0139746f $X=11.105 $Y=2.31 $X2=0
+ $Y2=0
cc_1634 N_A_2189_47#_c_2069_n N_Z_c_3437_n 0.00749574f $X=11.335 $Y=1.405 $X2=0
+ $Y2=0
cc_1635 N_A_2189_47#_c_2070_n N_Z_c_3437_n 0.00449418f $X=11.555 $Y=1.34 $X2=0
+ $Y2=0
cc_1636 N_A_2189_47#_M1078_d VGND 0.00358139f $X=10.945 $Y=0.235 $X2=0 $Y2=0
cc_1637 N_A_2189_47#_c_2071_n VGND 0.0150148f $X=11.105 $Y=0.495 $X2=0 $Y2=0
cc_1638 N_A_2189_47#_c_2071_n N_VGND_c_4411_n 0.015238f $X=11.105 $Y=0.495 $X2=0
+ $Y2=0
cc_1639 N_A_2189_937#_M1008_g N_D[13]_c_2225_n 0.0390641f $X=11.86 $Y=3.365
+ $X2=-0.19 $Y2=-0.24
cc_1640 N_A_2189_937#_c_2127_n N_D[13]_c_2225_n 0.00216577f $X=11.555 $Y=4.1
+ $X2=-0.19 $Y2=-0.24
cc_1641 N_A_2189_937#_c_2127_n N_D[13]_c_2222_n 0.00496096f $X=11.555 $Y=4.1
+ $X2=0 $Y2=0
cc_1642 N_A_2189_937#_c_2130_n N_VPWR_c_2833_n 0.0292866f $X=11.105 $Y=3.13
+ $X2=0 $Y2=0
cc_1643 N_A_2189_937#_c_2126_n N_VPWR_c_2833_n 0.00688579f $X=11.335 $Y=4.035
+ $X2=0 $Y2=0
cc_1644 N_A_2189_937#_M1008_g N_VPWR_c_2835_n 0.00258498f $X=11.86 $Y=3.365
+ $X2=0 $Y2=0
cc_1645 N_A_2189_937#_M1049_d VPWR 0.00179197f $X=10.96 $Y=2.955 $X2=0 $Y2=0
cc_1646 N_A_2189_937#_M1008_g VPWR 0.00387928f $X=11.86 $Y=3.365 $X2=0 $Y2=0
cc_1647 N_A_2189_937#_c_2130_n VPWR 0.00594162f $X=11.105 $Y=3.13 $X2=0 $Y2=0
cc_1648 N_A_2189_937#_c_2130_n N_VPWR_c_2856_n 0.0210596f $X=11.105 $Y=3.13
+ $X2=0 $Y2=0
cc_1649 N_A_2189_937#_M1008_g N_Z_c_3384_n 0.00544362f $X=11.86 $Y=3.365 $X2=0
+ $Y2=0
cc_1650 N_A_2189_937#_c_2125_n N_Z_c_3342_n 0.00611965f $X=11.335 $Y=4.685 $X2=0
+ $Y2=0
cc_1651 N_A_2189_937#_c_2128_n N_Z_c_3342_n 0.0259454f $X=11.105 $Y=4.945 $X2=0
+ $Y2=0
cc_1652 N_A_2189_937#_M1008_g N_Z_c_3344_n 0.00862328f $X=11.86 $Y=3.365 $X2=0
+ $Y2=0
cc_1653 N_A_2189_937#_c_2130_n N_Z_c_3344_n 0.00378484f $X=11.105 $Y=3.13 $X2=0
+ $Y2=0
cc_1654 N_A_2189_937#_c_2125_n N_Z_c_3344_n 0.00719188f $X=11.335 $Y=4.685 $X2=0
+ $Y2=0
cc_1655 N_A_2189_937#_c_2126_n N_Z_c_3344_n 0.0304368f $X=11.335 $Y=4.035 $X2=0
+ $Y2=0
cc_1656 N_A_2189_937#_c_2127_n N_Z_c_3344_n 0.00814206f $X=11.555 $Y=4.1 $X2=0
+ $Y2=0
cc_1657 N_A_2189_937#_M1008_g N_Z_c_3411_n 0.00335035f $X=11.86 $Y=3.365 $X2=0
+ $Y2=0
cc_1658 N_A_2189_937#_c_2130_n N_Z_c_3411_n 0.0371028f $X=11.105 $Y=3.13 $X2=0
+ $Y2=0
cc_1659 N_A_2189_937#_M1008_g N_Z_c_3412_n 0.00502861f $X=11.86 $Y=3.365 $X2=0
+ $Y2=0
cc_1660 N_A_2189_937#_c_2125_n N_Z_c_3360_n 0.0124144f $X=11.335 $Y=4.685 $X2=0
+ $Y2=0
cc_1661 N_A_2189_937#_c_2126_n N_Z_c_3360_n 0.00398133f $X=11.335 $Y=4.035 $X2=0
+ $Y2=0
cc_1662 N_A_2189_937#_c_2127_n N_Z_c_3360_n 0.00349316f $X=11.555 $Y=4.1 $X2=0
+ $Y2=0
cc_1663 N_A_2189_937#_c_2130_n N_Z_c_3424_n 0.0291787f $X=11.105 $Y=3.13 $X2=0
+ $Y2=0
cc_1664 N_A_2189_937#_c_2126_n N_Z_c_3424_n 0.0126642f $X=11.335 $Y=4.035 $X2=0
+ $Y2=0
cc_1665 N_A_2189_937#_M1008_g N_Z_c_3898_n 0.00289142f $X=11.86 $Y=3.365 $X2=0
+ $Y2=0
cc_1666 N_A_2189_937#_c_2130_n N_Z_c_3898_n 6.03258e-19 $X=11.105 $Y=3.13 $X2=0
+ $Y2=0
cc_1667 N_A_2189_937#_c_2126_n N_Z_c_3898_n 4.25753e-19 $X=11.335 $Y=4.035 $X2=0
+ $Y2=0
cc_1668 N_A_2189_937#_M1008_g N_Z_c_3438_n 0.0107344f $X=11.86 $Y=3.365 $X2=0
+ $Y2=0
cc_1669 N_A_2189_937#_c_2130_n N_Z_c_3438_n 0.0139746f $X=11.105 $Y=3.13 $X2=0
+ $Y2=0
cc_1670 N_A_2189_937#_c_2126_n N_Z_c_3438_n 0.00749574f $X=11.335 $Y=4.035 $X2=0
+ $Y2=0
cc_1671 N_A_2189_937#_c_2127_n N_Z_c_3438_n 0.00449418f $X=11.555 $Y=4.1 $X2=0
+ $Y2=0
cc_1672 N_A_2189_937#_M1070_d VGND 0.00358139f $X=10.945 $Y=4.685 $X2=0 $Y2=0
cc_1673 N_A_2189_937#_c_2128_n VGND 0.0150148f $X=11.105 $Y=4.945 $X2=0 $Y2=0
cc_1674 N_A_2189_937#_c_2128_n N_VGND_c_4412_n 0.015238f $X=11.105 $Y=4.945
+ $X2=0 $Y2=0
cc_1675 N_D[5]_c_2184_n N_D[13]_c_2225_n 0.0129371f $X=12.385 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_1676 N_D[5]_c_2185_n N_D[6]_c_2263_n 0.00915308f $X=12.41 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_1677 N_D[5]_c_2184_n N_D[6]_c_2264_n 0.0270908f $X=12.385 $Y=1.41 $X2=0 $Y2=0
cc_1678 N_D[5]_c_2187_n N_D[6]_c_2264_n 9.4377e-19 $X=12.38 $Y=1.16 $X2=0 $Y2=0
cc_1679 N_D[5]_c_2186_n N_D[6]_c_2265_n 0.00442615f $X=12.235 $Y=1.055 $X2=0
+ $Y2=0
cc_1680 N_D[5]_c_2184_n N_D[6]_c_2266_n 9.4377e-19 $X=12.385 $Y=1.41 $X2=0 $Y2=0
cc_1681 N_D[5]_c_2187_n N_D[6]_c_2266_n 0.0199139f $X=12.38 $Y=1.16 $X2=0 $Y2=0
cc_1682 N_D[5]_c_2184_n N_VPWR_c_2834_n 0.0220781f $X=12.385 $Y=1.41 $X2=0 $Y2=0
cc_1683 N_D[5]_c_2187_n N_VPWR_c_2834_n 0.0044581f $X=12.38 $Y=1.16 $X2=0 $Y2=0
cc_1684 N_D[5]_c_2184_n VPWR 0.00468368f $X=12.385 $Y=1.41 $X2=0 $Y2=0
cc_1685 N_D[5]_c_2184_n N_VPWR_c_2857_n 0.00342413f $X=12.385 $Y=1.41 $X2=0
+ $Y2=0
cc_1686 N_D[5]_c_2184_n N_Z_c_3383_n 0.00176496f $X=12.385 $Y=1.41 $X2=0 $Y2=0
cc_1687 N_D[5]_c_2186_n N_Z_c_3341_n 0.00686805f $X=12.235 $Y=1.055 $X2=0 $Y2=0
cc_1688 N_D[5]_c_2184_n N_Z_c_3343_n 0.00605747f $X=12.385 $Y=1.41 $X2=0 $Y2=0
cc_1689 N_D[5]_c_2186_n N_Z_c_3343_n 0.00376465f $X=12.235 $Y=1.055 $X2=0 $Y2=0
cc_1690 N_D[5]_c_2187_n N_Z_c_3343_n 0.0216525f $X=12.38 $Y=1.16 $X2=0 $Y2=0
cc_1691 N_D[5]_c_2186_n N_Z_c_3359_n 0.0128881f $X=12.235 $Y=1.055 $X2=0 $Y2=0
cc_1692 N_D[5]_c_2184_n N_Z_c_3911_n 0.00719456f $X=12.385 $Y=1.41 $X2=0 $Y2=0
cc_1693 N_D[5]_c_2187_n N_Z_c_3911_n 0.00989895f $X=12.38 $Y=1.16 $X2=0 $Y2=0
cc_1694 N_D[5]_c_2184_n N_Z_c_3437_n 8.42164e-19 $X=12.385 $Y=1.41 $X2=0 $Y2=0
cc_1695 N_D[5]_c_2185_n N_VGND_c_4381_n 0.00322791f $X=12.41 $Y=0.995 $X2=0
+ $Y2=0
cc_1696 N_D[5]_c_2187_n N_VGND_c_4381_n 0.00222881f $X=12.38 $Y=1.16 $X2=0 $Y2=0
cc_1697 N_D[5]_c_2185_n VGND 0.0108306f $X=12.41 $Y=0.995 $X2=0 $Y2=0
cc_1698 N_D[5]_c_2217_p VGND 0.00942277f $X=12.235 $Y=0.51 $X2=0 $Y2=0
cc_1699 N_D[5]_c_2185_n N_VGND_c_4411_n 0.00585385f $X=12.41 $Y=0.995 $X2=0
+ $Y2=0
cc_1700 N_D[5]_c_2217_p N_VGND_c_4411_n 0.00842546f $X=12.235 $Y=0.51 $X2=0
+ $Y2=0
cc_1701 N_D[5]_c_2186_n A_2402_47# 0.00426617f $X=12.235 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_1702 N_D[5]_c_2217_p A_2402_47# 0.00894235f $X=12.235 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_1703 N_D[13]_c_2222_n N_D[14]_c_2301_n 0.0287172f $X=12.41 $Y=4.445 $X2=-0.19
+ $Y2=-0.24
cc_1704 N_D[13]_c_2224_n N_D[14]_c_2301_n 9.4377e-19 $X=12.38 $Y=4.28 $X2=-0.19
+ $Y2=-0.24
cc_1705 N_D[13]_c_2225_n N_D[14]_c_2305_n 0.00752667f $X=12.385 $Y=4.03 $X2=0
+ $Y2=0
cc_1706 N_D[13]_c_2223_n N_D[14]_c_2302_n 0.00442615f $X=12.235 $Y=4.815 $X2=0
+ $Y2=0
cc_1707 N_D[13]_c_2222_n N_D[14]_c_2303_n 9.4377e-19 $X=12.41 $Y=4.445 $X2=0
+ $Y2=0
cc_1708 N_D[13]_c_2224_n N_D[14]_c_2303_n 0.0199139f $X=12.38 $Y=4.28 $X2=0
+ $Y2=0
cc_1709 N_D[13]_c_2225_n N_VPWR_c_2835_n 0.0220781f $X=12.385 $Y=4.03 $X2=0
+ $Y2=0
cc_1710 N_D[13]_c_2224_n N_VPWR_c_2835_n 0.0044581f $X=12.38 $Y=4.28 $X2=0 $Y2=0
cc_1711 N_D[13]_c_2225_n VPWR 0.00468368f $X=12.385 $Y=4.03 $X2=0 $Y2=0
cc_1712 N_D[13]_c_2225_n N_VPWR_c_2857_n 0.00342413f $X=12.385 $Y=4.03 $X2=0
+ $Y2=0
cc_1713 N_D[13]_c_2223_n N_Z_c_3342_n 0.00686805f $X=12.235 $Y=4.815 $X2=0 $Y2=0
cc_1714 N_D[13]_c_2225_n N_Z_c_3344_n 0.00305841f $X=12.385 $Y=4.03 $X2=0 $Y2=0
cc_1715 N_D[13]_c_2222_n N_Z_c_3344_n 0.00299906f $X=12.41 $Y=4.445 $X2=0 $Y2=0
cc_1716 N_D[13]_c_2223_n N_Z_c_3344_n 0.00376465f $X=12.235 $Y=4.815 $X2=0 $Y2=0
cc_1717 N_D[13]_c_2224_n N_Z_c_3344_n 0.0216525f $X=12.38 $Y=4.28 $X2=0 $Y2=0
cc_1718 N_D[13]_c_2225_n N_Z_c_3412_n 0.00176496f $X=12.385 $Y=4.03 $X2=0 $Y2=0
cc_1719 N_D[13]_c_2223_n N_Z_c_3360_n 0.0128881f $X=12.235 $Y=4.815 $X2=0 $Y2=0
cc_1720 N_D[13]_c_2225_n N_Z_c_3921_n 0.0061664f $X=12.385 $Y=4.03 $X2=0 $Y2=0
cc_1721 N_D[13]_c_2222_n N_Z_c_3921_n 0.00102816f $X=12.41 $Y=4.445 $X2=0 $Y2=0
cc_1722 N_D[13]_c_2224_n N_Z_c_3921_n 0.00989895f $X=12.38 $Y=4.28 $X2=0 $Y2=0
cc_1723 N_D[13]_c_2225_n N_Z_c_3438_n 8.42164e-19 $X=12.385 $Y=4.03 $X2=0 $Y2=0
cc_1724 N_D[13]_c_2222_n N_VGND_c_4382_n 0.00322791f $X=12.41 $Y=4.445 $X2=0
+ $Y2=0
cc_1725 N_D[13]_c_2224_n N_VGND_c_4382_n 0.00222881f $X=12.38 $Y=4.28 $X2=0
+ $Y2=0
cc_1726 N_D[13]_c_2222_n VGND 0.0108306f $X=12.41 $Y=4.445 $X2=0 $Y2=0
cc_1727 N_D[13]_c_2258_p VGND 0.00941728f $X=12.235 $Y=4.93 $X2=0 $Y2=0
cc_1728 N_D[13]_c_2222_n N_VGND_c_4412_n 0.00585385f $X=12.41 $Y=4.445 $X2=0
+ $Y2=0
cc_1729 N_D[13]_c_2258_p N_VGND_c_4412_n 0.00842546f $X=12.235 $Y=4.93 $X2=0
+ $Y2=0
cc_1730 N_D[13]_c_2223_n A_2402_937# 0.00426617f $X=12.235 $Y=4.815 $X2=-0.19
+ $Y2=-0.24
cc_1731 N_D[13]_c_2258_p A_2402_937# 0.00894235f $X=12.235 $Y=4.93 $X2=-0.19
+ $Y2=-0.24
cc_1732 N_D[6]_c_2264_n N_D[14]_c_2305_n 0.0129371f $X=12.915 $Y=1.41 $X2=0
+ $Y2=0
cc_1733 N_D[6]_c_2264_n N_A_2668_265#_M1051_g 0.0390641f $X=12.915 $Y=1.41 $X2=0
+ $Y2=0
cc_1734 N_D[6]_c_2264_n N_A_2668_265#_c_2345_n 0.00712672f $X=12.915 $Y=1.41
+ $X2=0 $Y2=0
cc_1735 N_D[6]_c_2263_n N_S[6]_c_2456_n 0.0286599f $X=12.89 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_1736 N_D[6]_c_2265_n N_S[6]_c_2456_n 0.00289497f $X=13.065 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_1737 N_D[6]_c_2264_n N_VPWR_c_2834_n 0.0220781f $X=12.915 $Y=1.41 $X2=0 $Y2=0
cc_1738 N_D[6]_c_2266_n N_VPWR_c_2834_n 0.0044581f $X=13.065 $Y=1.19 $X2=0 $Y2=0
cc_1739 N_D[6]_c_2264_n VPWR 0.00468368f $X=12.915 $Y=1.41 $X2=0 $Y2=0
cc_1740 N_D[6]_c_2264_n N_VPWR_c_2858_n 0.00342413f $X=12.915 $Y=1.41 $X2=0
+ $Y2=0
cc_1741 N_D[6]_c_2264_n N_Z_c_3345_n 0.00605747f $X=12.915 $Y=1.41 $X2=0 $Y2=0
cc_1742 N_D[6]_c_2265_n N_Z_c_3345_n 0.00376465f $X=13.065 $Y=1.055 $X2=0 $Y2=0
cc_1743 N_D[6]_c_2266_n N_Z_c_3345_n 0.0216525f $X=13.065 $Y=1.19 $X2=0 $Y2=0
cc_1744 N_D[6]_c_2265_n N_Z_c_3347_n 0.0128881f $X=13.065 $Y=1.055 $X2=0 $Y2=0
cc_1745 N_D[6]_c_2265_n N_Z_c_3348_n 0.00686805f $X=13.065 $Y=1.055 $X2=0 $Y2=0
cc_1746 N_D[6]_c_2264_n N_Z_c_3389_n 0.00176496f $X=12.915 $Y=1.41 $X2=0 $Y2=0
cc_1747 N_D[6]_c_2264_n N_Z_c_3911_n 0.00719456f $X=12.915 $Y=1.41 $X2=0 $Y2=0
cc_1748 N_D[6]_c_2266_n N_Z_c_3911_n 0.00989895f $X=13.065 $Y=1.19 $X2=0 $Y2=0
cc_1749 N_D[6]_c_2264_n N_Z_c_3439_n 8.42164e-19 $X=12.915 $Y=1.41 $X2=0 $Y2=0
cc_1750 N_D[6]_c_2263_n N_VGND_c_4381_n 0.00322791f $X=12.89 $Y=0.995 $X2=0
+ $Y2=0
cc_1751 N_D[6]_c_2266_n N_VGND_c_4381_n 0.00222881f $X=13.065 $Y=1.19 $X2=0
+ $Y2=0
cc_1752 N_D[6]_c_2263_n N_VGND_c_4401_n 0.00585385f $X=12.89 $Y=0.995 $X2=0
+ $Y2=0
cc_1753 D[6] N_VGND_c_4401_n 0.00842546f $X=13.025 $Y=0.425 $X2=0 $Y2=0
cc_1754 N_D[6]_c_2263_n VGND 0.0108306f $X=12.89 $Y=0.995 $X2=0 $Y2=0
cc_1755 D[6] VGND 0.00942277f $X=13.025 $Y=0.425 $X2=0 $Y2=0
cc_1756 N_D[6]_c_2265_n A_2593_47# 0.00426617f $X=13.065 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_1757 D[6] A_2593_47# 0.00894235f $X=13.025 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_1758 N_D[14]_c_2305_n N_A_2668_793#_M1004_g 0.0390641f $X=12.915 $Y=4.03
+ $X2=0 $Y2=0
cc_1759 N_D[14]_c_2301_n N_A_2668_793#_c_2402_n 0.00496096f $X=12.89 $Y=4.445
+ $X2=0 $Y2=0
cc_1760 N_D[14]_c_2305_n N_A_2668_793#_c_2402_n 0.00216577f $X=12.915 $Y=4.03
+ $X2=0 $Y2=0
cc_1761 N_D[14]_c_2301_n N_S[14]_c_2507_n 0.0286599f $X=12.89 $Y=4.445 $X2=0
+ $Y2=0
cc_1762 N_D[14]_c_2302_n N_S[14]_c_2507_n 0.00289497f $X=13.065 $Y=4.815 $X2=0
+ $Y2=0
cc_1763 N_D[14]_c_2305_n N_VPWR_c_2835_n 0.0220781f $X=12.915 $Y=4.03 $X2=0
+ $Y2=0
cc_1764 N_D[14]_c_2303_n N_VPWR_c_2835_n 0.0044581f $X=13.065 $Y=4.25 $X2=0
+ $Y2=0
cc_1765 N_D[14]_c_2305_n VPWR 0.00468368f $X=12.915 $Y=4.03 $X2=0 $Y2=0
cc_1766 N_D[14]_c_2305_n N_VPWR_c_2858_n 0.00342413f $X=12.915 $Y=4.03 $X2=0
+ $Y2=0
cc_1767 N_D[14]_c_2301_n N_Z_c_3346_n 0.00299906f $X=12.89 $Y=4.445 $X2=0 $Y2=0
cc_1768 N_D[14]_c_2305_n N_Z_c_3346_n 0.00305841f $X=12.915 $Y=4.03 $X2=0 $Y2=0
cc_1769 N_D[14]_c_2302_n N_Z_c_3346_n 0.00376465f $X=13.065 $Y=4.815 $X2=0 $Y2=0
cc_1770 N_D[14]_c_2303_n N_Z_c_3346_n 0.0216525f $X=13.065 $Y=4.25 $X2=0 $Y2=0
cc_1771 N_D[14]_c_2302_n N_Z_c_3349_n 0.0128881f $X=13.065 $Y=4.815 $X2=0 $Y2=0
cc_1772 N_D[14]_c_2302_n N_Z_c_3350_n 0.00686805f $X=13.065 $Y=4.815 $X2=0 $Y2=0
cc_1773 N_D[14]_c_2305_n N_Z_c_3415_n 0.00176496f $X=12.915 $Y=4.03 $X2=0 $Y2=0
cc_1774 N_D[14]_c_2301_n N_Z_c_3921_n 0.00102816f $X=12.89 $Y=4.445 $X2=0 $Y2=0
cc_1775 N_D[14]_c_2305_n N_Z_c_3921_n 0.0061664f $X=12.915 $Y=4.03 $X2=0 $Y2=0
cc_1776 N_D[14]_c_2303_n N_Z_c_3921_n 0.00989895f $X=13.065 $Y=4.25 $X2=0 $Y2=0
cc_1777 N_D[14]_c_2305_n N_Z_c_3440_n 8.42164e-19 $X=12.915 $Y=4.03 $X2=0 $Y2=0
cc_1778 N_D[14]_c_2301_n N_VGND_c_4382_n 0.00322791f $X=12.89 $Y=4.445 $X2=0
+ $Y2=0
cc_1779 N_D[14]_c_2303_n N_VGND_c_4382_n 0.00222881f $X=13.065 $Y=4.25 $X2=0
+ $Y2=0
cc_1780 N_D[14]_c_2301_n N_VGND_c_4403_n 0.00585385f $X=12.89 $Y=4.445 $X2=0
+ $Y2=0
cc_1781 D[14] N_VGND_c_4403_n 0.00842546f $X=13.025 $Y=4.845 $X2=0 $Y2=0
cc_1782 N_D[14]_c_2301_n VGND 0.0108306f $X=12.89 $Y=4.445 $X2=0 $Y2=0
cc_1783 D[14] VGND 0.00941728f $X=13.025 $Y=4.845 $X2=0 $Y2=0
cc_1784 N_D[14]_c_2302_n A_2593_911# 0.00426617f $X=13.065 $Y=4.815 $X2=-0.19
+ $Y2=-0.24
cc_1785 D[14] A_2593_911# 0.00894235f $X=13.025 $Y=4.845 $X2=-0.19 $Y2=-0.24
cc_1786 N_A_2668_265#_M1051_g N_A_2668_793#_M1004_g 0.0129371f $X=13.44 $Y=2.075
+ $X2=0 $Y2=0
cc_1787 N_A_2668_265#_c_2342_n N_S[6]_c_2457_n 0.00827389f $X=13.965 $Y=0.755
+ $X2=0 $Y2=0
cc_1788 N_A_2668_265#_c_2343_n N_S[6]_c_2457_n 0.0164662f $X=13.965 $Y=1.175
+ $X2=0 $Y2=0
cc_1789 N_A_2668_265#_c_2344_n N_S[6]_c_2457_n 0.00928634f $X=14.195 $Y=1.63
+ $X2=0 $Y2=0
cc_1790 N_A_2668_265#_c_2345_n N_S[6]_c_2457_n 0.0184911f $X=13.44 $Y=1.34 $X2=0
+ $Y2=0
cc_1791 N_A_2668_265#_c_2345_n N_S[6]_c_2458_n 0.00820745f $X=13.44 $Y=1.34
+ $X2=0 $Y2=0
cc_1792 N_A_2668_265#_c_2343_n N_S[6]_c_2459_n 0.0012443f $X=13.965 $Y=1.175
+ $X2=0 $Y2=0
cc_1793 N_A_2668_265#_c_2347_n N_S[6]_c_2459_n 0.00902681f $X=14.195 $Y=2.31
+ $X2=0 $Y2=0
cc_1794 N_A_2668_265#_c_2344_n N_S[6]_c_2459_n 0.00767015f $X=14.195 $Y=1.63
+ $X2=0 $Y2=0
cc_1795 N_A_2668_265#_c_2345_n N_S[6]_c_2459_n 0.00659591f $X=13.44 $Y=1.34
+ $X2=0 $Y2=0
cc_1796 N_A_2668_265#_c_2343_n N_S[6]_c_2460_n 0.00219336f $X=13.965 $Y=1.175
+ $X2=0 $Y2=0
cc_1797 N_A_2668_265#_c_2342_n N_S[6]_c_2461_n 0.00603567f $X=13.965 $Y=0.755
+ $X2=0 $Y2=0
cc_1798 N_A_2668_265#_c_2343_n N_S[6]_c_2461_n 0.0178233f $X=13.965 $Y=1.175
+ $X2=0 $Y2=0
cc_1799 N_A_2668_265#_c_2344_n N_S[6]_c_2461_n 0.0214702f $X=14.195 $Y=1.63
+ $X2=0 $Y2=0
cc_1800 N_A_2668_265#_c_2345_n N_S[6]_c_2461_n 2.59957e-19 $X=13.44 $Y=1.34
+ $X2=0 $Y2=0
cc_1801 N_A_2668_265#_M1051_g N_VPWR_c_2834_n 0.00258498f $X=13.44 $Y=2.075
+ $X2=0 $Y2=0
cc_1802 N_A_2668_265#_c_2347_n N_VPWR_c_2836_n 0.0292866f $X=14.195 $Y=2.31
+ $X2=0 $Y2=0
cc_1803 N_A_2668_265#_c_2344_n N_VPWR_c_2836_n 0.00688579f $X=14.195 $Y=1.63
+ $X2=0 $Y2=0
cc_1804 N_A_2668_265#_c_2347_n N_VPWR_c_2846_n 0.0210596f $X=14.195 $Y=2.31
+ $X2=0 $Y2=0
cc_1805 N_A_2668_265#_M1066_s VPWR 0.00179197f $X=14.07 $Y=1.485 $X2=0 $Y2=0
cc_1806 N_A_2668_265#_M1051_g VPWR 0.00387928f $X=13.44 $Y=2.075 $X2=0 $Y2=0
cc_1807 N_A_2668_265#_c_2347_n VPWR 0.00594162f $X=14.195 $Y=2.31 $X2=0 $Y2=0
cc_1808 N_A_2668_265#_M1051_g N_Z_c_3345_n 0.00862328f $X=13.44 $Y=2.075 $X2=0
+ $Y2=0
cc_1809 N_A_2668_265#_c_2343_n N_Z_c_3345_n 0.00719188f $X=13.965 $Y=1.175 $X2=0
+ $Y2=0
cc_1810 N_A_2668_265#_c_2347_n N_Z_c_3345_n 0.00378484f $X=14.195 $Y=2.31 $X2=0
+ $Y2=0
cc_1811 N_A_2668_265#_c_2344_n N_Z_c_3345_n 0.0304368f $X=14.195 $Y=1.63 $X2=0
+ $Y2=0
cc_1812 N_A_2668_265#_c_2345_n N_Z_c_3345_n 0.00814206f $X=13.44 $Y=1.34 $X2=0
+ $Y2=0
cc_1813 N_A_2668_265#_c_2343_n N_Z_c_3347_n 0.0124144f $X=13.965 $Y=1.175 $X2=0
+ $Y2=0
cc_1814 N_A_2668_265#_c_2344_n N_Z_c_3347_n 0.00398133f $X=14.195 $Y=1.63 $X2=0
+ $Y2=0
cc_1815 N_A_2668_265#_c_2345_n N_Z_c_3347_n 0.00349316f $X=13.44 $Y=1.34 $X2=0
+ $Y2=0
cc_1816 N_A_2668_265#_c_2342_n N_Z_c_3348_n 0.0259454f $X=13.965 $Y=0.755 $X2=0
+ $Y2=0
cc_1817 N_A_2668_265#_c_2343_n N_Z_c_3348_n 0.00611965f $X=13.965 $Y=1.175 $X2=0
+ $Y2=0
cc_1818 N_A_2668_265#_M1051_g N_Z_c_3389_n 0.00544362f $X=13.44 $Y=2.075 $X2=0
+ $Y2=0
cc_1819 N_A_2668_265#_c_2347_n N_Z_c_3389_n 0.0371028f $X=14.195 $Y=2.31 $X2=0
+ $Y2=0
cc_1820 N_A_2668_265#_M1051_g N_Z_c_3413_n 0.00335035f $X=13.44 $Y=2.075 $X2=0
+ $Y2=0
cc_1821 N_A_2668_265#_M1051_g N_Z_c_3415_n 0.00502861f $X=13.44 $Y=2.075 $X2=0
+ $Y2=0
cc_1822 N_A_2668_265#_c_2347_n N_Z_c_3425_n 0.0291787f $X=14.195 $Y=2.31 $X2=0
+ $Y2=0
cc_1823 N_A_2668_265#_c_2344_n N_Z_c_3425_n 0.0126642f $X=14.195 $Y=1.63 $X2=0
+ $Y2=0
cc_1824 N_A_2668_265#_M1051_g N_Z_c_3961_n 0.00289142f $X=13.44 $Y=2.075 $X2=0
+ $Y2=0
cc_1825 N_A_2668_265#_c_2347_n N_Z_c_3961_n 6.03258e-19 $X=14.195 $Y=2.31 $X2=0
+ $Y2=0
cc_1826 N_A_2668_265#_c_2344_n N_Z_c_3961_n 4.25753e-19 $X=14.195 $Y=1.63 $X2=0
+ $Y2=0
cc_1827 N_A_2668_265#_M1051_g N_Z_c_3439_n 0.0107335f $X=13.44 $Y=2.075 $X2=0
+ $Y2=0
cc_1828 N_A_2668_265#_c_2347_n N_Z_c_3439_n 0.0139746f $X=14.195 $Y=2.31 $X2=0
+ $Y2=0
cc_1829 N_A_2668_265#_c_2344_n N_Z_c_3439_n 0.00749574f $X=14.195 $Y=1.63 $X2=0
+ $Y2=0
cc_1830 N_A_2668_265#_c_2345_n N_Z_c_3439_n 0.00449418f $X=13.44 $Y=1.34 $X2=0
+ $Y2=0
cc_1831 N_A_2668_265#_c_2342_n N_VGND_c_4401_n 0.015238f $X=13.965 $Y=0.755
+ $X2=0 $Y2=0
cc_1832 N_A_2668_265#_M1007_s VGND 0.00358139f $X=14.07 $Y=0.235 $X2=0 $Y2=0
cc_1833 N_A_2668_265#_c_2342_n VGND 0.0150148f $X=13.965 $Y=0.755 $X2=0 $Y2=0
cc_1834 N_A_2668_793#_c_2400_n N_S[14]_c_2506_n 0.0247401f $X=13.965 $Y=4.685
+ $X2=0 $Y2=0
cc_1835 N_A_2668_793#_c_2401_n N_S[14]_c_2506_n 0.00928634f $X=14.195 $Y=3.805
+ $X2=0 $Y2=0
cc_1836 N_A_2668_793#_c_2402_n N_S[14]_c_2506_n 0.0184911f $X=13.44 $Y=4.1 $X2=0
+ $Y2=0
cc_1837 N_A_2668_793#_c_2402_n N_S[14]_c_2507_n 0.00820745f $X=13.44 $Y=4.1
+ $X2=0 $Y2=0
cc_1838 N_A_2668_793#_c_2401_n N_S[14]_c_2510_n 0.00382813f $X=14.195 $Y=3.805
+ $X2=0 $Y2=0
cc_1839 N_A_2668_793#_c_2405_n N_S[14]_c_2510_n 0.00902681f $X=14.195 $Y=3.13
+ $X2=0 $Y2=0
cc_1840 N_A_2668_793#_c_2402_n N_S[14]_c_2510_n 0.00150889f $X=13.44 $Y=4.1
+ $X2=0 $Y2=0
cc_1841 N_A_2668_793#_c_2400_n N_S[14]_c_2508_n 0.00343766f $X=13.965 $Y=4.685
+ $X2=0 $Y2=0
cc_1842 N_A_2668_793#_c_2401_n N_S[14]_c_2508_n 0.00384202f $X=14.195 $Y=3.805
+ $X2=0 $Y2=0
cc_1843 N_A_2668_793#_c_2402_n N_S[14]_c_2508_n 0.00508702f $X=13.44 $Y=4.1
+ $X2=0 $Y2=0
cc_1844 N_A_2668_793#_c_2400_n S[14] 0.023859f $X=13.965 $Y=4.685 $X2=0 $Y2=0
cc_1845 N_A_2668_793#_c_2401_n S[14] 0.0214702f $X=14.195 $Y=3.805 $X2=0 $Y2=0
cc_1846 N_A_2668_793#_c_2402_n S[14] 2.59957e-19 $X=13.44 $Y=4.1 $X2=0 $Y2=0
cc_1847 N_A_2668_793#_M1004_g N_VPWR_c_2835_n 0.00258498f $X=13.44 $Y=3.365
+ $X2=0 $Y2=0
cc_1848 N_A_2668_793#_c_2401_n N_VPWR_c_2837_n 0.00688579f $X=14.195 $Y=3.805
+ $X2=0 $Y2=0
cc_1849 N_A_2668_793#_c_2405_n N_VPWR_c_2837_n 0.0292866f $X=14.195 $Y=3.13
+ $X2=0 $Y2=0
cc_1850 N_A_2668_793#_c_2405_n N_VPWR_c_2846_n 0.0210596f $X=14.195 $Y=3.13
+ $X2=0 $Y2=0
cc_1851 N_A_2668_793#_M1072_s VPWR 0.00179197f $X=14.07 $Y=2.955 $X2=0 $Y2=0
cc_1852 N_A_2668_793#_M1004_g VPWR 0.00387928f $X=13.44 $Y=3.365 $X2=0 $Y2=0
cc_1853 N_A_2668_793#_c_2405_n VPWR 0.00594162f $X=14.195 $Y=3.13 $X2=0 $Y2=0
cc_1854 N_A_2668_793#_M1004_g N_Z_c_3346_n 0.00862328f $X=13.44 $Y=3.365 $X2=0
+ $Y2=0
cc_1855 N_A_2668_793#_c_2400_n N_Z_c_3346_n 0.00719188f $X=13.965 $Y=4.685 $X2=0
+ $Y2=0
cc_1856 N_A_2668_793#_c_2401_n N_Z_c_3346_n 0.0304368f $X=14.195 $Y=3.805 $X2=0
+ $Y2=0
cc_1857 N_A_2668_793#_c_2405_n N_Z_c_3346_n 0.00378484f $X=14.195 $Y=3.13 $X2=0
+ $Y2=0
cc_1858 N_A_2668_793#_c_2402_n N_Z_c_3346_n 0.00814206f $X=13.44 $Y=4.1 $X2=0
+ $Y2=0
cc_1859 N_A_2668_793#_c_2400_n N_Z_c_3349_n 0.0124144f $X=13.965 $Y=4.685 $X2=0
+ $Y2=0
cc_1860 N_A_2668_793#_c_2401_n N_Z_c_3349_n 0.00398133f $X=14.195 $Y=3.805 $X2=0
+ $Y2=0
cc_1861 N_A_2668_793#_c_2402_n N_Z_c_3349_n 0.00349316f $X=13.44 $Y=4.1 $X2=0
+ $Y2=0
cc_1862 N_A_2668_793#_c_2400_n N_Z_c_3350_n 0.032065f $X=13.965 $Y=4.685 $X2=0
+ $Y2=0
cc_1863 N_A_2668_793#_M1004_g N_Z_c_3390_n 0.00544362f $X=13.44 $Y=3.365 $X2=0
+ $Y2=0
cc_1864 N_A_2668_793#_M1004_g N_Z_c_3414_n 0.00335035f $X=13.44 $Y=3.365 $X2=0
+ $Y2=0
cc_1865 N_A_2668_793#_c_2405_n N_Z_c_3414_n 0.0371028f $X=14.195 $Y=3.13 $X2=0
+ $Y2=0
cc_1866 N_A_2668_793#_M1004_g N_Z_c_3415_n 0.00502861f $X=13.44 $Y=3.365 $X2=0
+ $Y2=0
cc_1867 N_A_2668_793#_c_2401_n N_Z_c_3426_n 0.0126642f $X=14.195 $Y=3.805 $X2=0
+ $Y2=0
cc_1868 N_A_2668_793#_c_2405_n N_Z_c_3426_n 0.0291787f $X=14.195 $Y=3.13 $X2=0
+ $Y2=0
cc_1869 N_A_2668_793#_M1004_g N_Z_c_3983_n 0.00289142f $X=13.44 $Y=3.365 $X2=0
+ $Y2=0
cc_1870 N_A_2668_793#_c_2401_n N_Z_c_3983_n 4.25753e-19 $X=14.195 $Y=3.805 $X2=0
+ $Y2=0
cc_1871 N_A_2668_793#_c_2405_n N_Z_c_3983_n 6.03258e-19 $X=14.195 $Y=3.13 $X2=0
+ $Y2=0
cc_1872 N_A_2668_793#_M1004_g N_Z_c_3440_n 0.0107344f $X=13.44 $Y=3.365 $X2=0
+ $Y2=0
cc_1873 N_A_2668_793#_c_2401_n N_Z_c_3440_n 0.00749574f $X=14.195 $Y=3.805 $X2=0
+ $Y2=0
cc_1874 N_A_2668_793#_c_2405_n N_Z_c_3440_n 0.0139746f $X=14.195 $Y=3.13 $X2=0
+ $Y2=0
cc_1875 N_A_2668_793#_c_2402_n N_Z_c_3440_n 0.00449418f $X=13.44 $Y=4.1 $X2=0
+ $Y2=0
cc_1876 N_A_2668_793#_c_2400_n N_VGND_c_4403_n 0.015238f $X=13.965 $Y=4.685
+ $X2=0 $Y2=0
cc_1877 N_A_2668_793#_M1026_s VGND 0.00358139f $X=14.07 $Y=4.685 $X2=0 $Y2=0
cc_1878 N_A_2668_793#_c_2400_n VGND 0.0150148f $X=13.965 $Y=4.685 $X2=0 $Y2=0
cc_1879 N_S[6]_c_2459_n N_S[14]_c_2510_n 0.0130744f $X=14.43 $Y=1.41 $X2=0 $Y2=0
cc_1880 N_S[6]_c_2459_n N_S[7]_c_2553_n 0.0578733f $X=14.43 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_1881 N_S[6]_c_2461_n N_S[7]_c_2553_n 0.00112057f $X=14.395 $Y=1.03 $X2=-0.19
+ $Y2=-0.24
cc_1882 N_S[6]_c_2460_n N_S[7]_c_2554_n 0.0091402f $X=14.43 $Y=0.83 $X2=0 $Y2=0
cc_1883 N_S[6]_c_2459_n N_S[7]_c_2557_n 0.00112057f $X=14.43 $Y=1.41 $X2=0 $Y2=0
cc_1884 N_S[6]_c_2461_n N_S[7]_c_2557_n 0.0277403f $X=14.395 $Y=1.03 $X2=0 $Y2=0
cc_1885 N_S[6]_c_2459_n N_VPWR_c_2836_n 0.00965725f $X=14.43 $Y=1.41 $X2=0 $Y2=0
cc_1886 N_S[6]_c_2461_n N_VPWR_c_2836_n 0.00587376f $X=14.395 $Y=1.03 $X2=0
+ $Y2=0
cc_1887 N_S[6]_c_2459_n N_VPWR_c_2846_n 0.0035837f $X=14.43 $Y=1.41 $X2=0 $Y2=0
cc_1888 N_S[6]_c_2459_n VPWR 0.0072999f $X=14.43 $Y=1.41 $X2=0 $Y2=0
cc_1889 N_S[6]_c_2458_n N_Z_c_3345_n 7.46972e-19 $X=13.44 $Y=0.905 $X2=0 $Y2=0
cc_1890 N_S[6]_c_2457_n N_Z_c_3347_n 0.00806549f $X=14.26 $Y=0.905 $X2=0 $Y2=0
cc_1891 N_S[6]_c_2458_n N_Z_c_3347_n 0.00605736f $X=13.44 $Y=0.905 $X2=0 $Y2=0
cc_1892 N_S[6]_c_2456_n N_Z_c_3348_n 0.00316445f $X=13.365 $Y=0.83 $X2=0 $Y2=0
cc_1893 N_S[6]_c_2457_n N_Z_c_3348_n 0.00501353f $X=14.26 $Y=0.905 $X2=0 $Y2=0
cc_1894 N_S[6]_c_2459_n N_Z_c_3415_n 0.00124373f $X=14.43 $Y=1.41 $X2=0 $Y2=0
cc_1895 N_S[6]_c_2459_n N_Z_c_3425_n 0.0062071f $X=14.43 $Y=1.41 $X2=0 $Y2=0
cc_1896 N_S[6]_c_2461_n N_Z_c_3425_n 0.00659242f $X=14.395 $Y=1.03 $X2=0 $Y2=0
cc_1897 N_S[6]_c_2460_n N_VGND_c_4383_n 0.00570474f $X=14.43 $Y=0.83 $X2=0 $Y2=0
cc_1898 N_S[6]_c_2461_n N_VGND_c_4383_n 0.00391126f $X=14.395 $Y=1.03 $X2=0
+ $Y2=0
cc_1899 N_S[6]_c_2456_n N_VGND_c_4401_n 0.00585385f $X=13.365 $Y=0.83 $X2=0
+ $Y2=0
cc_1900 N_S[6]_c_2460_n N_VGND_c_4401_n 0.00585385f $X=14.43 $Y=0.83 $X2=0 $Y2=0
cc_1901 N_S[6]_c_2456_n VGND 0.00880034f $X=13.365 $Y=0.83 $X2=0 $Y2=0
cc_1902 N_S[6]_c_2457_n VGND 0.00349917f $X=14.26 $Y=0.905 $X2=0 $Y2=0
cc_1903 N_S[6]_c_2459_n VGND 6.15795e-19 $X=14.43 $Y=1.41 $X2=0 $Y2=0
cc_1904 N_S[6]_c_2460_n VGND 0.0124506f $X=14.43 $Y=0.83 $X2=0 $Y2=0
cc_1905 N_S[14]_c_2510_n N_S[15]_c_2603_n 0.0296874f $X=14.43 $Y=4.03 $X2=-0.19
+ $Y2=-0.24
cc_1906 N_S[14]_c_2508_n N_S[15]_c_2599_n 0.0373261f $X=14.43 $Y=4.61 $X2=0
+ $Y2=0
cc_1907 S[14] N_S[15]_c_2599_n 0.00112057f $X=14.405 $Y=4.165 $X2=0 $Y2=0
cc_1908 N_S[14]_c_2508_n S[15] 0.00112057f $X=14.43 $Y=4.61 $X2=0 $Y2=0
cc_1909 S[14] S[15] 0.0277403f $X=14.405 $Y=4.165 $X2=0 $Y2=0
cc_1910 N_S[14]_c_2510_n N_VPWR_c_2837_n 0.00965725f $X=14.43 $Y=4.03 $X2=0
+ $Y2=0
cc_1911 S[14] N_VPWR_c_2837_n 0.00587376f $X=14.405 $Y=4.165 $X2=0 $Y2=0
cc_1912 N_S[14]_c_2510_n N_VPWR_c_2846_n 0.0035837f $X=14.43 $Y=4.03 $X2=0 $Y2=0
cc_1913 N_S[14]_c_2510_n VPWR 0.0072999f $X=14.43 $Y=4.03 $X2=0 $Y2=0
cc_1914 N_S[14]_c_2507_n N_Z_c_3346_n 7.46972e-19 $X=13.44 $Y=4.535 $X2=0 $Y2=0
cc_1915 N_S[14]_c_2506_n N_Z_c_3349_n 0.00806549f $X=14.26 $Y=4.535 $X2=0 $Y2=0
cc_1916 N_S[14]_c_2507_n N_Z_c_3349_n 0.00605736f $X=13.44 $Y=4.535 $X2=0 $Y2=0
cc_1917 N_S[14]_c_2505_n N_Z_c_3350_n 0.00316445f $X=13.365 $Y=4.61 $X2=0 $Y2=0
cc_1918 N_S[14]_c_2506_n N_Z_c_3350_n 0.00501353f $X=14.26 $Y=4.535 $X2=0 $Y2=0
cc_1919 N_S[14]_c_2510_n N_Z_c_3415_n 0.00124373f $X=14.43 $Y=4.03 $X2=0 $Y2=0
cc_1920 N_S[14]_c_2510_n N_Z_c_3426_n 0.00597491f $X=14.43 $Y=4.03 $X2=0 $Y2=0
cc_1921 N_S[14]_c_2508_n N_Z_c_3426_n 2.32192e-19 $X=14.43 $Y=4.61 $X2=0 $Y2=0
cc_1922 S[14] N_Z_c_3426_n 0.00659242f $X=14.405 $Y=4.165 $X2=0 $Y2=0
cc_1923 N_S[14]_c_2508_n N_VGND_c_4384_n 0.00570474f $X=14.43 $Y=4.61 $X2=0
+ $Y2=0
cc_1924 S[14] N_VGND_c_4384_n 0.00391126f $X=14.405 $Y=4.165 $X2=0 $Y2=0
cc_1925 N_S[14]_c_2505_n N_VGND_c_4403_n 0.00585385f $X=13.365 $Y=4.61 $X2=0
+ $Y2=0
cc_1926 N_S[14]_c_2508_n N_VGND_c_4403_n 0.00585385f $X=14.43 $Y=4.61 $X2=0
+ $Y2=0
cc_1927 N_S[14]_c_2505_n VGND 0.00880034f $X=13.365 $Y=4.61 $X2=0 $Y2=0
cc_1928 N_S[14]_c_2506_n VGND 0.00349917f $X=14.26 $Y=4.535 $X2=0 $Y2=0
cc_1929 N_S[14]_c_2508_n VGND 0.0130664f $X=14.43 $Y=4.61 $X2=0 $Y2=0
cc_1930 N_S[7]_c_2553_n N_S[15]_c_2603_n 0.0130744f $X=15.01 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_1931 N_S[7]_c_2553_n N_A_3017_47#_c_2651_n 0.00902681f $X=15.01 $Y=1.41 $X2=0
+ $Y2=0
cc_1932 N_S[7]_c_2553_n N_A_3017_47#_c_2646_n 0.0012443f $X=15.01 $Y=1.41 $X2=0
+ $Y2=0
cc_1933 N_S[7]_c_2554_n N_A_3017_47#_c_2646_n 0.00219336f $X=15.01 $Y=0.83 $X2=0
+ $Y2=0
cc_1934 N_S[7]_c_2555_n N_A_3017_47#_c_2646_n 0.0164662f $X=16 $Y=0.905 $X2=0
+ $Y2=0
cc_1935 N_S[7]_c_2557_n N_A_3017_47#_c_2646_n 0.0178233f $X=15.045 $Y=1.03 $X2=0
+ $Y2=0
cc_1936 N_S[7]_c_2553_n N_A_3017_47#_c_2647_n 0.00767015f $X=15.01 $Y=1.41 $X2=0
+ $Y2=0
cc_1937 N_S[7]_c_2555_n N_A_3017_47#_c_2647_n 0.00928634f $X=16 $Y=0.905 $X2=0
+ $Y2=0
cc_1938 N_S[7]_c_2557_n N_A_3017_47#_c_2647_n 0.0214702f $X=15.045 $Y=1.03 $X2=0
+ $Y2=0
cc_1939 N_S[7]_c_2553_n N_A_3017_47#_c_2648_n 0.00659591f $X=15.01 $Y=1.41 $X2=0
+ $Y2=0
cc_1940 N_S[7]_c_2555_n N_A_3017_47#_c_2648_n 0.0266986f $X=16 $Y=0.905 $X2=0
+ $Y2=0
cc_1941 N_S[7]_c_2557_n N_A_3017_47#_c_2648_n 2.59957e-19 $X=15.045 $Y=1.03
+ $X2=0 $Y2=0
cc_1942 N_S[7]_c_2553_n N_A_3017_47#_c_2649_n 0.00827389f $X=15.01 $Y=1.41 $X2=0
+ $Y2=0
cc_1943 N_S[7]_c_2557_n N_A_3017_47#_c_2649_n 0.00603567f $X=15.045 $Y=1.03
+ $X2=0 $Y2=0
cc_1944 N_S[7]_c_2556_n N_D[7]_c_2763_n 0.0286599f $X=16.075 $Y=0.83 $X2=0 $Y2=0
cc_1945 N_S[7]_c_2556_n N_D[7]_c_2764_n 0.00289497f $X=16.075 $Y=0.83 $X2=0
+ $Y2=0
cc_1946 N_S[7]_c_2553_n N_VPWR_c_2836_n 0.00965725f $X=15.01 $Y=1.41 $X2=0 $Y2=0
cc_1947 N_S[7]_c_2557_n N_VPWR_c_2836_n 0.00587376f $X=15.045 $Y=1.03 $X2=0
+ $Y2=0
cc_1948 N_S[7]_c_2553_n VPWR 0.0072999f $X=15.01 $Y=1.41 $X2=0 $Y2=0
cc_1949 N_S[7]_c_2553_n N_VPWR_c_2859_n 0.0035837f $X=15.01 $Y=1.41 $X2=0 $Y2=0
cc_1950 N_S[7]_c_2555_n N_Z_c_3351_n 0.00501353f $X=16 $Y=0.905 $X2=0 $Y2=0
cc_1951 N_S[7]_c_2556_n N_Z_c_3351_n 0.00316445f $X=16.075 $Y=0.83 $X2=0 $Y2=0
cc_1952 N_S[7]_c_2555_n N_Z_c_3353_n 7.46972e-19 $X=16 $Y=0.905 $X2=0 $Y2=0
cc_1953 N_S[7]_c_2553_n N_Z_c_3418_n 0.00124373f $X=15.01 $Y=1.41 $X2=0 $Y2=0
cc_1954 N_S[7]_c_2555_n N_Z_c_3361_n 0.0141229f $X=16 $Y=0.905 $X2=0 $Y2=0
cc_1955 N_S[7]_c_2553_n N_Z_c_3425_n 0.0062071f $X=15.01 $Y=1.41 $X2=0 $Y2=0
cc_1956 N_S[7]_c_2557_n N_Z_c_3425_n 0.00659242f $X=15.045 $Y=1.03 $X2=0 $Y2=0
cc_1957 N_S[7]_c_2554_n N_VGND_c_4383_n 0.00570474f $X=15.01 $Y=0.83 $X2=0 $Y2=0
cc_1958 N_S[7]_c_2557_n N_VGND_c_4383_n 0.00391126f $X=15.045 $Y=1.03 $X2=0
+ $Y2=0
cc_1959 N_S[7]_c_2553_n VGND 6.15795e-19 $X=15.01 $Y=1.41 $X2=0 $Y2=0
cc_1960 N_S[7]_c_2554_n VGND 0.0124506f $X=15.01 $Y=0.83 $X2=0 $Y2=0
cc_1961 N_S[7]_c_2555_n VGND 0.00349917f $X=16 $Y=0.905 $X2=0 $Y2=0
cc_1962 N_S[7]_c_2556_n VGND 0.00880034f $X=16.075 $Y=0.83 $X2=0 $Y2=0
cc_1963 N_S[7]_c_2554_n N_VGND_c_4413_n 0.00585385f $X=15.01 $Y=0.83 $X2=0 $Y2=0
cc_1964 N_S[7]_c_2556_n N_VGND_c_4413_n 0.00585385f $X=16.075 $Y=0.83 $X2=0
+ $Y2=0
cc_1965 N_S[15]_c_2603_n N_A_3017_937#_c_2708_n 0.00902681f $X=15.01 $Y=4.03
+ $X2=0 $Y2=0
cc_1966 N_S[15]_c_2599_n N_A_3017_937#_c_2703_n 0.00343766f $X=15.01 $Y=4.61
+ $X2=0 $Y2=0
cc_1967 N_S[15]_c_2600_n N_A_3017_937#_c_2703_n 0.0164662f $X=16 $Y=4.535 $X2=0
+ $Y2=0
cc_1968 S[15] N_A_3017_937#_c_2703_n 0.0178233f $X=14.865 $Y=4.165 $X2=0 $Y2=0
cc_1969 N_S[15]_c_2603_n N_A_3017_937#_c_2704_n 0.00382813f $X=15.01 $Y=4.03
+ $X2=0 $Y2=0
cc_1970 N_S[15]_c_2599_n N_A_3017_937#_c_2704_n 0.00384202f $X=15.01 $Y=4.61
+ $X2=0 $Y2=0
cc_1971 N_S[15]_c_2600_n N_A_3017_937#_c_2704_n 0.00928634f $X=16 $Y=4.535 $X2=0
+ $Y2=0
cc_1972 S[15] N_A_3017_937#_c_2704_n 0.0214702f $X=14.865 $Y=4.165 $X2=0 $Y2=0
cc_1973 N_S[15]_c_2603_n N_A_3017_937#_c_2705_n 0.00150889f $X=15.01 $Y=4.03
+ $X2=0 $Y2=0
cc_1974 N_S[15]_c_2599_n N_A_3017_937#_c_2705_n 0.00508702f $X=15.01 $Y=4.61
+ $X2=0 $Y2=0
cc_1975 N_S[15]_c_2600_n N_A_3017_937#_c_2705_n 0.0266986f $X=16 $Y=4.535 $X2=0
+ $Y2=0
cc_1976 S[15] N_A_3017_937#_c_2705_n 2.59957e-19 $X=14.865 $Y=4.165 $X2=0 $Y2=0
cc_1977 N_S[15]_c_2599_n N_A_3017_937#_c_2706_n 0.00827389f $X=15.01 $Y=4.61
+ $X2=0 $Y2=0
cc_1978 S[15] N_A_3017_937#_c_2706_n 0.00603567f $X=14.865 $Y=4.165 $X2=0 $Y2=0
cc_1979 N_S[15]_c_2600_n N_D[15]_c_2791_n 0.0286599f $X=16 $Y=4.535 $X2=0 $Y2=0
cc_1980 N_S[15]_c_2600_n N_D[15]_c_2792_n 0.00289497f $X=16 $Y=4.535 $X2=0 $Y2=0
cc_1981 N_S[15]_c_2603_n N_VPWR_c_2837_n 0.00965725f $X=15.01 $Y=4.03 $X2=0
+ $Y2=0
cc_1982 S[15] N_VPWR_c_2837_n 0.00587376f $X=14.865 $Y=4.165 $X2=0 $Y2=0
cc_1983 N_S[15]_c_2603_n VPWR 0.0072999f $X=15.01 $Y=4.03 $X2=0 $Y2=0
cc_1984 N_S[15]_c_2603_n N_VPWR_c_2859_n 0.0035837f $X=15.01 $Y=4.03 $X2=0 $Y2=0
cc_1985 N_S[15]_c_2600_n N_Z_c_3352_n 0.00501353f $X=16 $Y=4.535 $X2=0 $Y2=0
cc_1986 N_S[15]_c_2601_n N_Z_c_3352_n 0.00316445f $X=16.075 $Y=4.61 $X2=0 $Y2=0
cc_1987 N_S[15]_c_2600_n N_Z_c_3354_n 7.46972e-19 $X=16 $Y=4.535 $X2=0 $Y2=0
cc_1988 N_S[15]_c_2603_n N_Z_c_3418_n 0.00124373f $X=15.01 $Y=4.03 $X2=0 $Y2=0
cc_1989 N_S[15]_c_2600_n N_Z_c_3362_n 0.0141229f $X=16 $Y=4.535 $X2=0 $Y2=0
cc_1990 N_S[15]_c_2603_n N_Z_c_3426_n 0.00597491f $X=15.01 $Y=4.03 $X2=0 $Y2=0
cc_1991 N_S[15]_c_2599_n N_Z_c_3426_n 2.32192e-19 $X=15.01 $Y=4.61 $X2=0 $Y2=0
cc_1992 S[15] N_Z_c_3426_n 0.00659242f $X=14.865 $Y=4.165 $X2=0 $Y2=0
cc_1993 N_S[15]_c_2599_n N_VGND_c_4384_n 0.00570474f $X=15.01 $Y=4.61 $X2=0
+ $Y2=0
cc_1994 S[15] N_VGND_c_4384_n 0.00391126f $X=14.865 $Y=4.165 $X2=0 $Y2=0
cc_1995 N_S[15]_c_2599_n VGND 0.0130664f $X=15.01 $Y=4.61 $X2=0 $Y2=0
cc_1996 N_S[15]_c_2600_n VGND 0.00349917f $X=16 $Y=4.535 $X2=0 $Y2=0
cc_1997 N_S[15]_c_2601_n VGND 0.00880034f $X=16.075 $Y=4.61 $X2=0 $Y2=0
cc_1998 N_S[15]_c_2599_n N_VGND_c_4414_n 0.00585385f $X=15.01 $Y=4.61 $X2=0
+ $Y2=0
cc_1999 N_S[15]_c_2601_n N_VGND_c_4414_n 0.00585385f $X=16.075 $Y=4.61 $X2=0
+ $Y2=0
cc_2000 N_A_3017_47#_M1093_g N_A_3017_937#_M1038_g 0.0129371f $X=16 $Y=2.075
+ $X2=0 $Y2=0
cc_2001 N_A_3017_47#_M1093_g N_D[7]_c_2762_n 0.0383393f $X=16 $Y=2.075 $X2=-0.19
+ $Y2=-0.24
cc_2002 N_A_3017_47#_c_2648_n N_D[7]_c_2762_n 0.00712672f $X=15.695 $Y=1.34
+ $X2=-0.19 $Y2=-0.24
cc_2003 N_A_3017_47#_c_2651_n N_VPWR_c_2836_n 0.0292866f $X=15.245 $Y=2.31 $X2=0
+ $Y2=0
cc_2004 N_A_3017_47#_c_2647_n N_VPWR_c_2836_n 0.00688579f $X=15.475 $Y=1.405
+ $X2=0 $Y2=0
cc_2005 N_A_3017_47#_M1093_g N_VPWR_c_2838_n 0.00247893f $X=16 $Y=2.075 $X2=0
+ $Y2=0
cc_2006 N_A_3017_47#_M1019_d VPWR 0.00179197f $X=15.1 $Y=1.485 $X2=0 $Y2=0
cc_2007 N_A_3017_47#_M1093_g VPWR 0.00407291f $X=16 $Y=2.075 $X2=0 $Y2=0
cc_2008 N_A_3017_47#_c_2651_n VPWR 0.00594162f $X=15.245 $Y=2.31 $X2=0 $Y2=0
cc_2009 N_A_3017_47#_c_2651_n N_VPWR_c_2859_n 0.0210596f $X=15.245 $Y=2.31 $X2=0
+ $Y2=0
cc_2010 N_A_3017_47#_M1093_g N_Z_c_3391_n 0.00544362f $X=16 $Y=2.075 $X2=0 $Y2=0
cc_2011 N_A_3017_47#_c_2651_n N_Z_c_3391_n 0.0371028f $X=15.245 $Y=2.31 $X2=0
+ $Y2=0
cc_2012 N_A_3017_47#_c_2646_n N_Z_c_3351_n 0.00611965f $X=15.475 $Y=1.175 $X2=0
+ $Y2=0
cc_2013 N_A_3017_47#_c_2649_n N_Z_c_3351_n 0.0259454f $X=15.245 $Y=0.495 $X2=0
+ $Y2=0
cc_2014 N_A_3017_47#_M1093_g N_Z_c_3353_n 0.00862328f $X=16 $Y=2.075 $X2=0 $Y2=0
cc_2015 N_A_3017_47#_c_2651_n N_Z_c_3353_n 0.00378484f $X=15.245 $Y=2.31 $X2=0
+ $Y2=0
cc_2016 N_A_3017_47#_c_2646_n N_Z_c_3353_n 0.00719188f $X=15.475 $Y=1.175 $X2=0
+ $Y2=0
cc_2017 N_A_3017_47#_c_2647_n N_Z_c_3353_n 0.0304368f $X=15.475 $Y=1.405 $X2=0
+ $Y2=0
cc_2018 N_A_3017_47#_c_2648_n N_Z_c_3353_n 0.00814206f $X=15.695 $Y=1.34 $X2=0
+ $Y2=0
cc_2019 N_A_3017_47#_M1093_g N_Z_c_3416_n 0.00335035f $X=16 $Y=2.075 $X2=0 $Y2=0
cc_2020 N_A_3017_47#_M1093_g N_Z_c_3418_n 0.00502861f $X=16 $Y=2.075 $X2=0 $Y2=0
cc_2021 N_A_3017_47#_c_2646_n N_Z_c_3361_n 0.0124144f $X=15.475 $Y=1.175 $X2=0
+ $Y2=0
cc_2022 N_A_3017_47#_c_2647_n N_Z_c_3361_n 0.00398133f $X=15.475 $Y=1.405 $X2=0
+ $Y2=0
cc_2023 N_A_3017_47#_c_2648_n N_Z_c_3361_n 0.00349316f $X=15.695 $Y=1.34 $X2=0
+ $Y2=0
cc_2024 N_A_3017_47#_c_2651_n N_Z_c_3425_n 0.0291787f $X=15.245 $Y=2.31 $X2=0
+ $Y2=0
cc_2025 N_A_3017_47#_c_2647_n N_Z_c_3425_n 0.0126642f $X=15.475 $Y=1.405 $X2=0
+ $Y2=0
cc_2026 N_A_3017_47#_M1093_g Z 0.00289142f $X=16 $Y=2.075 $X2=0 $Y2=0
cc_2027 N_A_3017_47#_c_2651_n Z 6.03258e-19 $X=15.245 $Y=2.31 $X2=0 $Y2=0
cc_2028 N_A_3017_47#_c_2647_n Z 4.25753e-19 $X=15.475 $Y=1.405 $X2=0 $Y2=0
cc_2029 N_A_3017_47#_M1093_g N_Z_c_3441_n 0.0107335f $X=16 $Y=2.075 $X2=0 $Y2=0
cc_2030 N_A_3017_47#_c_2651_n N_Z_c_3441_n 0.0139746f $X=15.245 $Y=2.31 $X2=0
+ $Y2=0
cc_2031 N_A_3017_47#_c_2647_n N_Z_c_3441_n 0.00749574f $X=15.475 $Y=1.405 $X2=0
+ $Y2=0
cc_2032 N_A_3017_47#_c_2648_n N_Z_c_3441_n 0.00449418f $X=15.695 $Y=1.34 $X2=0
+ $Y2=0
cc_2033 N_A_3017_47#_M1095_d VGND 0.00358139f $X=15.085 $Y=0.235 $X2=0 $Y2=0
cc_2034 N_A_3017_47#_c_2649_n VGND 0.0150148f $X=15.245 $Y=0.495 $X2=0 $Y2=0
cc_2035 N_A_3017_47#_c_2649_n N_VGND_c_4413_n 0.015238f $X=15.245 $Y=0.495 $X2=0
+ $Y2=0
cc_2036 N_A_3017_937#_M1038_g N_D[15]_c_2794_n 0.0383393f $X=16 $Y=3.365
+ $X2=-0.19 $Y2=-0.24
cc_2037 N_A_3017_937#_c_2705_n N_D[15]_c_2794_n 0.00216577f $X=15.695 $Y=4.1
+ $X2=-0.19 $Y2=-0.24
cc_2038 N_A_3017_937#_c_2705_n N_D[15]_c_2791_n 0.00496096f $X=15.695 $Y=4.1
+ $X2=0 $Y2=0
cc_2039 N_A_3017_937#_c_2708_n N_VPWR_c_2837_n 0.0292866f $X=15.245 $Y=3.13
+ $X2=0 $Y2=0
cc_2040 N_A_3017_937#_c_2704_n N_VPWR_c_2837_n 0.00688579f $X=15.475 $Y=4.035
+ $X2=0 $Y2=0
cc_2041 N_A_3017_937#_M1038_g N_VPWR_c_2839_n 0.00247893f $X=16 $Y=3.365 $X2=0
+ $Y2=0
cc_2042 N_A_3017_937#_M1021_d VPWR 0.00179197f $X=15.1 $Y=2.955 $X2=0 $Y2=0
cc_2043 N_A_3017_937#_M1038_g VPWR 0.00407291f $X=16 $Y=3.365 $X2=0 $Y2=0
cc_2044 N_A_3017_937#_c_2708_n VPWR 0.00594162f $X=15.245 $Y=3.13 $X2=0 $Y2=0
cc_2045 N_A_3017_937#_c_2708_n N_VPWR_c_2859_n 0.0210596f $X=15.245 $Y=3.13
+ $X2=0 $Y2=0
cc_2046 N_A_3017_937#_M1038_g N_Z_c_3392_n 0.00544362f $X=16 $Y=3.365 $X2=0
+ $Y2=0
cc_2047 N_A_3017_937#_c_2703_n N_Z_c_3352_n 0.00611965f $X=15.475 $Y=4.685 $X2=0
+ $Y2=0
cc_2048 N_A_3017_937#_c_2706_n N_Z_c_3352_n 0.0259454f $X=15.245 $Y=4.945 $X2=0
+ $Y2=0
cc_2049 N_A_3017_937#_M1038_g N_Z_c_3354_n 0.00862328f $X=16 $Y=3.365 $X2=0
+ $Y2=0
cc_2050 N_A_3017_937#_c_2708_n N_Z_c_3354_n 0.00378484f $X=15.245 $Y=3.13 $X2=0
+ $Y2=0
cc_2051 N_A_3017_937#_c_2703_n N_Z_c_3354_n 0.00719188f $X=15.475 $Y=4.685 $X2=0
+ $Y2=0
cc_2052 N_A_3017_937#_c_2704_n N_Z_c_3354_n 0.0304368f $X=15.475 $Y=4.035 $X2=0
+ $Y2=0
cc_2053 N_A_3017_937#_c_2705_n N_Z_c_3354_n 0.00814206f $X=15.695 $Y=4.1 $X2=0
+ $Y2=0
cc_2054 N_A_3017_937#_M1038_g N_Z_c_3417_n 0.00335035f $X=16 $Y=3.365 $X2=0
+ $Y2=0
cc_2055 N_A_3017_937#_c_2708_n N_Z_c_3417_n 0.0371028f $X=15.245 $Y=3.13 $X2=0
+ $Y2=0
cc_2056 N_A_3017_937#_M1038_g N_Z_c_3418_n 0.00502861f $X=16 $Y=3.365 $X2=0
+ $Y2=0
cc_2057 N_A_3017_937#_c_2703_n N_Z_c_3362_n 0.0124144f $X=15.475 $Y=4.685 $X2=0
+ $Y2=0
cc_2058 N_A_3017_937#_c_2704_n N_Z_c_3362_n 0.00398133f $X=15.475 $Y=4.035 $X2=0
+ $Y2=0
cc_2059 N_A_3017_937#_c_2705_n N_Z_c_3362_n 0.00349316f $X=15.695 $Y=4.1 $X2=0
+ $Y2=0
cc_2060 N_A_3017_937#_c_2708_n N_Z_c_3426_n 0.0291787f $X=15.245 $Y=3.13 $X2=0
+ $Y2=0
cc_2061 N_A_3017_937#_c_2704_n N_Z_c_3426_n 0.0126642f $X=15.475 $Y=4.035 $X2=0
+ $Y2=0
cc_2062 N_A_3017_937#_M1038_g Z 0.00289142f $X=16 $Y=3.365 $X2=0 $Y2=0
cc_2063 N_A_3017_937#_c_2708_n Z 6.03258e-19 $X=15.245 $Y=3.13 $X2=0 $Y2=0
cc_2064 N_A_3017_937#_c_2704_n Z 4.25753e-19 $X=15.475 $Y=4.035 $X2=0 $Y2=0
cc_2065 N_A_3017_937#_M1038_g N_Z_c_3442_n 0.0107344f $X=16 $Y=3.365 $X2=0 $Y2=0
cc_2066 N_A_3017_937#_c_2708_n N_Z_c_3442_n 0.0139746f $X=15.245 $Y=3.13 $X2=0
+ $Y2=0
cc_2067 N_A_3017_937#_c_2704_n N_Z_c_3442_n 0.00749574f $X=15.475 $Y=4.035 $X2=0
+ $Y2=0
cc_2068 N_A_3017_937#_c_2705_n N_Z_c_3442_n 0.00449418f $X=15.695 $Y=4.1 $X2=0
+ $Y2=0
cc_2069 N_A_3017_937#_M1073_d VGND 0.00358139f $X=15.085 $Y=4.685 $X2=0 $Y2=0
cc_2070 N_A_3017_937#_c_2706_n VGND 0.0150148f $X=15.245 $Y=4.945 $X2=0 $Y2=0
cc_2071 N_A_3017_937#_c_2706_n N_VGND_c_4414_n 0.015238f $X=15.245 $Y=4.945
+ $X2=0 $Y2=0
cc_2072 N_D[7]_c_2762_n N_D[15]_c_2794_n 0.0129371f $X=16.525 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_2073 N_D[7]_c_2762_n N_VPWR_c_2838_n 0.0235f $X=16.525 $Y=1.41 $X2=0 $Y2=0
cc_2074 N_D[7]_c_2765_n N_VPWR_c_2838_n 0.00471543f $X=16.52 $Y=1.16 $X2=0 $Y2=0
cc_2075 N_D[7]_c_2762_n VPWR 0.00937833f $X=16.525 $Y=1.41 $X2=0 $Y2=0
cc_2076 N_D[7]_c_2762_n N_VPWR_c_2860_n 0.00342413f $X=16.525 $Y=1.41 $X2=0
+ $Y2=0
cc_2077 N_D[7]_c_2762_n N_Z_c_3391_n 0.00176496f $X=16.525 $Y=1.41 $X2=0 $Y2=0
cc_2078 N_D[7]_c_2764_n N_Z_c_3351_n 0.00686805f $X=16.375 $Y=1.055 $X2=0 $Y2=0
cc_2079 N_D[7]_c_2762_n N_Z_c_3353_n 0.00605747f $X=16.525 $Y=1.41 $X2=0 $Y2=0
cc_2080 N_D[7]_c_2764_n N_Z_c_3353_n 0.00376465f $X=16.375 $Y=1.055 $X2=0 $Y2=0
cc_2081 N_D[7]_c_2765_n N_Z_c_3353_n 0.0216525f $X=16.52 $Y=1.16 $X2=0 $Y2=0
cc_2082 N_D[7]_c_2764_n N_Z_c_3361_n 0.0128881f $X=16.375 $Y=1.055 $X2=0 $Y2=0
cc_2083 N_D[7]_c_2763_n N_VGND_c_4386_n 0.00487865f $X=16.55 $Y=0.995 $X2=0
+ $Y2=0
cc_2084 N_D[7]_c_2765_n N_VGND_c_4386_n 0.00222881f $X=16.52 $Y=1.16 $X2=0 $Y2=0
cc_2085 N_D[7]_c_2763_n VGND 0.011617f $X=16.55 $Y=0.995 $X2=0 $Y2=0
cc_2086 N_D[7]_c_2786_p VGND 0.00942277f $X=16.375 $Y=0.51 $X2=0 $Y2=0
cc_2087 N_D[7]_c_2763_n N_VGND_c_4413_n 0.00585385f $X=16.55 $Y=0.995 $X2=0
+ $Y2=0
cc_2088 N_D[7]_c_2786_p N_VGND_c_4413_n 0.00842546f $X=16.375 $Y=0.51 $X2=0
+ $Y2=0
cc_2089 N_D[7]_c_2764_n A_3230_47# 0.00426617f $X=16.375 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_2090 N_D[7]_c_2786_p A_3230_47# 0.00894235f $X=16.375 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_2091 N_D[15]_c_2794_n N_VPWR_c_2839_n 0.0235f $X=16.525 $Y=4.03 $X2=0 $Y2=0
cc_2092 N_D[15]_c_2793_n N_VPWR_c_2839_n 0.00471543f $X=16.52 $Y=4.28 $X2=0
+ $Y2=0
cc_2093 N_D[15]_c_2794_n VPWR 0.00937833f $X=16.525 $Y=4.03 $X2=0 $Y2=0
cc_2094 N_D[15]_c_2794_n N_VPWR_c_2860_n 0.00342413f $X=16.525 $Y=4.03 $X2=0
+ $Y2=0
cc_2095 N_D[15]_c_2792_n N_Z_c_3352_n 0.00686805f $X=16.375 $Y=4.815 $X2=0 $Y2=0
cc_2096 N_D[15]_c_2794_n N_Z_c_3354_n 0.00305841f $X=16.525 $Y=4.03 $X2=0 $Y2=0
cc_2097 N_D[15]_c_2791_n N_Z_c_3354_n 0.00299906f $X=16.55 $Y=4.445 $X2=0 $Y2=0
cc_2098 N_D[15]_c_2792_n N_Z_c_3354_n 0.00376465f $X=16.375 $Y=4.815 $X2=0 $Y2=0
cc_2099 N_D[15]_c_2793_n N_Z_c_3354_n 0.0216525f $X=16.52 $Y=4.28 $X2=0 $Y2=0
cc_2100 N_D[15]_c_2794_n N_Z_c_3418_n 0.00176496f $X=16.525 $Y=4.03 $X2=0 $Y2=0
cc_2101 N_D[15]_c_2792_n N_Z_c_3362_n 0.0128881f $X=16.375 $Y=4.815 $X2=0 $Y2=0
cc_2102 N_D[15]_c_2791_n N_VGND_c_4388_n 0.00487865f $X=16.55 $Y=4.445 $X2=0
+ $Y2=0
cc_2103 N_D[15]_c_2793_n N_VGND_c_4388_n 0.00222881f $X=16.52 $Y=4.28 $X2=0
+ $Y2=0
cc_2104 N_D[15]_c_2791_n VGND 0.011617f $X=16.55 $Y=4.445 $X2=0 $Y2=0
cc_2105 N_D[15]_c_2817_p VGND 0.00941728f $X=16.375 $Y=4.93 $X2=0 $Y2=0
cc_2106 N_D[15]_c_2791_n N_VGND_c_4414_n 0.00585385f $X=16.55 $Y=4.445 $X2=0
+ $Y2=0
cc_2107 N_D[15]_c_2817_p N_VGND_c_4414_n 0.00842546f $X=16.375 $Y=4.93 $X2=0
+ $Y2=0
cc_2108 N_D[15]_c_2792_n A_3230_937# 0.00426617f $X=16.375 $Y=4.815 $X2=-0.19
+ $Y2=-0.24
cc_2109 N_D[15]_c_2817_p A_3230_937# 0.00894235f $X=16.375 $Y=4.93 $X2=-0.19
+ $Y2=-0.24
cc_2110 VPWR A_117_297# 0.0138589f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=1.305
cc_2111 VPWR A_117_591# 0.0138589f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=1.305
cc_2112 VPWR N_Z_M1036_d 5.61457e-19 $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2113 VPWR N_Z_M1090_d 5.61457e-19 $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2114 VPWR N_Z_M1017_s 5.61457e-19 $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2115 VPWR N_Z_M1071_s 5.61457e-19 $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2116 VPWR N_Z_M1041_d 5.61457e-19 $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2117 VPWR N_Z_M1000_d 5.61457e-19 $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2118 VPWR N_Z_M1022_s 5.61457e-19 $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2119 VPWR N_Z_M1074_s 5.61457e-19 $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2120 VPWR N_Z_M1014_d 5.61457e-19 $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2121 VPWR N_Z_M1064_d 5.61457e-19 $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2122 VPWR N_Z_M1059_s 5.61457e-19 $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2123 VPWR N_Z_M1008_s 5.61457e-19 $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2124 VPWR N_Z_M1051_d 5.61457e-19 $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2125 VPWR N_Z_M1004_d 5.61457e-19 $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2126 VPWR N_Z_M1093_s 5.61457e-19 $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2127 VPWR N_Z_M1038_s 5.61457e-19 $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2128 N_VPWR_c_2822_n N_Z_c_3315_n 0.00734981f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_2129 N_VPWR_c_2823_n N_Z_c_3316_n 0.00734981f $X=0.26 $Y=3.1 $X2=0 $Y2=0
cc_2130 N_VPWR_c_2822_n N_Z_c_3365_n 0.012112f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_2131 N_VPWR_c_2826_n N_Z_c_3367_n 0.0122518f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_2132 N_VPWR_c_2826_n N_Z_c_3323_n 0.0074594f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_2133 N_VPWR_c_2827_n N_Z_c_3324_n 0.0074594f $X=4.37 $Y=3.1 $X2=0 $Y2=0
cc_2134 N_VPWR_c_2826_n N_Z_c_3325_n 0.0074594f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_2135 N_VPWR_c_2827_n N_Z_c_3326_n 0.0074594f $X=4.37 $Y=3.1 $X2=0 $Y2=0
cc_2136 N_VPWR_c_2826_n N_Z_c_3373_n 0.0122518f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_2137 N_VPWR_c_2830_n N_Z_c_3375_n 0.0122518f $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_2138 N_VPWR_c_2830_n N_Z_c_3333_n 0.0074594f $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_2139 N_VPWR_c_2831_n N_Z_c_3334_n 0.0074594f $X=8.51 $Y=3.1 $X2=0 $Y2=0
cc_2140 N_VPWR_c_2830_n N_Z_c_3335_n 0.0074594f $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_2141 N_VPWR_c_2831_n N_Z_c_3336_n 0.0074594f $X=8.51 $Y=3.1 $X2=0 $Y2=0
cc_2142 N_VPWR_c_2830_n N_Z_c_3381_n 0.0122518f $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_2143 N_VPWR_c_2834_n N_Z_c_3383_n 0.0122518f $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_2144 N_VPWR_c_2834_n N_Z_c_3343_n 0.0074594f $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_2145 N_VPWR_c_2835_n N_Z_c_3344_n 0.0074594f $X=12.65 $Y=3.1 $X2=0 $Y2=0
cc_2146 N_VPWR_c_2834_n N_Z_c_3345_n 0.0074594f $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_2147 N_VPWR_c_2835_n N_Z_c_3346_n 0.0074594f $X=12.65 $Y=3.1 $X2=0 $Y2=0
cc_2148 N_VPWR_c_2834_n N_Z_c_3389_n 0.0122518f $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_2149 N_VPWR_c_2838_n N_Z_c_3391_n 0.012112f $X=16.76 $Y=1.66 $X2=0 $Y2=0
cc_2150 N_VPWR_c_2838_n N_Z_c_3353_n 0.00734981f $X=16.76 $Y=1.66 $X2=0 $Y2=0
cc_2151 N_VPWR_c_2839_n N_Z_c_3354_n 0.00734981f $X=16.76 $Y=3.1 $X2=0 $Y2=0
cc_2152 VPWR N_Z_c_3395_n 0.00328229f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2153 VPWR N_Z_c_3396_n 0.00328229f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2154 N_VPWR_c_2823_n N_Z_c_3397_n 0.012112f $X=0.26 $Y=3.1 $X2=0 $Y2=0
cc_2155 N_VPWR_c_2840_n N_Z_c_3397_n 0.0122229f $X=2.135 $Y=2.72 $X2=0 $Y2=0
cc_2156 VPWR N_Z_c_3397_n 0.0412991f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2157 N_VPWR_c_2849_n N_Z_c_3397_n 0.0122229f $X=0.69 $Y=2.72 $X2=0 $Y2=0
cc_2158 VPWR N_Z_c_3398_n 0.00328229f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2159 VPWR N_Z_c_3399_n 0.00328229f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2160 N_VPWR_c_2827_n N_Z_c_3400_n 0.0122518f $X=4.37 $Y=3.1 $X2=0 $Y2=0
cc_2161 VPWR N_Z_c_3400_n 0.0412991f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2162 N_VPWR_c_2850_n N_Z_c_3400_n 0.0122229f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_2163 N_VPWR_c_2851_n N_Z_c_3400_n 0.0122229f $X=4.175 $Y=2.72 $X2=0 $Y2=0
cc_2164 VPWR N_Z_c_3401_n 0.00328229f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2165 VPWR N_Z_c_3402_n 0.00328229f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2166 N_VPWR_c_2827_n N_Z_c_3403_n 0.0122518f $X=4.37 $Y=3.1 $X2=0 $Y2=0
cc_2167 N_VPWR_c_2842_n N_Z_c_3403_n 0.0122229f $X=6.275 $Y=2.72 $X2=0 $Y2=0
cc_2168 VPWR N_Z_c_3403_n 0.0412991f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2169 N_VPWR_c_2852_n N_Z_c_3403_n 0.0122229f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_2170 VPWR N_Z_c_3404_n 0.00328229f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2171 VPWR N_Z_c_3405_n 0.00328229f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2172 N_VPWR_c_2831_n N_Z_c_3406_n 0.0122518f $X=8.51 $Y=3.1 $X2=0 $Y2=0
cc_2173 VPWR N_Z_c_3406_n 0.0412991f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2174 N_VPWR_c_2853_n N_Z_c_3406_n 0.0122229f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_2175 N_VPWR_c_2854_n N_Z_c_3406_n 0.0122229f $X=8.315 $Y=2.72 $X2=0 $Y2=0
cc_2176 VPWR N_Z_c_3407_n 0.00328229f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2177 VPWR N_Z_c_3408_n 0.00328229f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2178 N_VPWR_c_2831_n N_Z_c_3409_n 0.0122518f $X=8.51 $Y=3.1 $X2=0 $Y2=0
cc_2179 N_VPWR_c_2844_n N_Z_c_3409_n 0.0122229f $X=10.415 $Y=2.72 $X2=0 $Y2=0
cc_2180 VPWR N_Z_c_3409_n 0.0412991f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2181 N_VPWR_c_2855_n N_Z_c_3409_n 0.0122229f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_2182 VPWR N_Z_c_3410_n 0.00328229f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2183 VPWR N_Z_c_3411_n 0.00328229f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2184 N_VPWR_c_2835_n N_Z_c_3412_n 0.0122518f $X=12.65 $Y=3.1 $X2=0 $Y2=0
cc_2185 VPWR N_Z_c_3412_n 0.0412991f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2186 N_VPWR_c_2856_n N_Z_c_3412_n 0.0122229f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_2187 N_VPWR_c_2857_n N_Z_c_3412_n 0.0122229f $X=12.455 $Y=2.72 $X2=0 $Y2=0
cc_2188 VPWR N_Z_c_3413_n 0.00328229f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2189 VPWR N_Z_c_3414_n 0.00328229f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2190 N_VPWR_c_2835_n N_Z_c_3415_n 0.0122518f $X=12.65 $Y=3.1 $X2=0 $Y2=0
cc_2191 N_VPWR_c_2846_n N_Z_c_3415_n 0.0122229f $X=14.555 $Y=2.72 $X2=0 $Y2=0
cc_2192 VPWR N_Z_c_3415_n 0.0412991f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2193 N_VPWR_c_2858_n N_Z_c_3415_n 0.0122229f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_2194 VPWR N_Z_c_3416_n 0.00328229f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2195 VPWR N_Z_c_3417_n 0.00328229f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2196 N_VPWR_c_2839_n N_Z_c_3418_n 0.012112f $X=16.76 $Y=3.1 $X2=0 $Y2=0
cc_2197 VPWR N_Z_c_3418_n 0.0412991f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2198 N_VPWR_c_2859_n N_Z_c_3418_n 0.0122229f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_2199 N_VPWR_c_2860_n N_Z_c_3418_n 0.0122229f $X=16.595 $Y=2.72 $X2=0 $Y2=0
cc_2200 N_VPWR_M1045_d N_Z_c_3419_n 0.001769f $X=2.1 $Y=1.485 $X2=0 $Y2=0
cc_2201 N_VPWR_c_2824_n N_Z_c_3419_n 0.0291114f $X=2.3 $Y=1.63 $X2=0 $Y2=0
cc_2202 VPWR N_Z_c_3419_n 0.094685f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2203 N_VPWR_c_2822_n N_Z_c_3472_n 0.00119119f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_2204 VPWR N_Z_c_3472_n 0.0135621f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2205 N_VPWR_M1048_d N_Z_c_3420_n 0.001769f $X=2.1 $Y=2.955 $X2=0 $Y2=0
cc_2206 N_VPWR_c_2825_n N_Z_c_3420_n 0.0291114f $X=2.3 $Y=3.13 $X2=0 $Y2=0
cc_2207 VPWR N_Z_c_3420_n 0.094685f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2208 N_VPWR_c_2823_n N_Z_c_3494_n 0.00119119f $X=0.26 $Y=3.1 $X2=0 $Y2=0
cc_2209 VPWR N_Z_c_3494_n 0.0135621f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2210 N_VPWR_c_2826_n N_Z_c_3585_n 0.0355595f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_2211 VPWR N_Z_c_3585_n 0.0739714f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2212 N_VPWR_c_2826_n N_Z_c_3549_n 4.83404e-19 $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_2213 VPWR N_Z_c_3549_n 0.0135621f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2214 N_VPWR_c_2827_n N_Z_c_3595_n 0.0355595f $X=4.37 $Y=3.1 $X2=0 $Y2=0
cc_2215 VPWR N_Z_c_3595_n 0.0739714f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2216 N_VPWR_c_2827_n N_Z_c_3572_n 4.83404e-19 $X=4.37 $Y=3.1 $X2=0 $Y2=0
cc_2217 VPWR N_Z_c_3572_n 0.0135621f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2218 N_VPWR_M1050_d N_Z_c_3421_n 0.001769f $X=6.24 $Y=1.485 $X2=0 $Y2=0
cc_2219 N_VPWR_c_2828_n N_Z_c_3421_n 0.0291114f $X=6.44 $Y=1.63 $X2=0 $Y2=0
cc_2220 VPWR N_Z_c_3421_n 0.094685f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2221 N_VPWR_c_2826_n N_Z_c_3635_n 4.83404e-19 $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_2222 VPWR N_Z_c_3635_n 0.0135621f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2223 N_VPWR_M1053_d N_Z_c_3422_n 0.001769f $X=6.24 $Y=2.955 $X2=0 $Y2=0
cc_2224 N_VPWR_c_2829_n N_Z_c_3422_n 0.0291114f $X=6.44 $Y=3.13 $X2=0 $Y2=0
cc_2225 VPWR N_Z_c_3422_n 0.094685f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2226 N_VPWR_c_2827_n N_Z_c_3657_n 4.83404e-19 $X=4.37 $Y=3.1 $X2=0 $Y2=0
cc_2227 VPWR N_Z_c_3657_n 0.0135621f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2228 N_VPWR_c_2830_n N_Z_c_3748_n 0.0355595f $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_2229 VPWR N_Z_c_3748_n 0.0739714f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2230 N_VPWR_c_2830_n N_Z_c_3712_n 4.83404e-19 $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_2231 VPWR N_Z_c_3712_n 0.0135621f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2232 N_VPWR_c_2831_n N_Z_c_3758_n 0.0355595f $X=8.51 $Y=3.1 $X2=0 $Y2=0
cc_2233 VPWR N_Z_c_3758_n 0.0739714f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2234 N_VPWR_c_2831_n N_Z_c_3735_n 4.83404e-19 $X=8.51 $Y=3.1 $X2=0 $Y2=0
cc_2235 VPWR N_Z_c_3735_n 0.0135621f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2236 N_VPWR_M1080_d N_Z_c_3423_n 0.001769f $X=10.38 $Y=1.485 $X2=0 $Y2=0
cc_2237 N_VPWR_c_2832_n N_Z_c_3423_n 0.0291114f $X=10.58 $Y=1.63 $X2=0 $Y2=0
cc_2238 VPWR N_Z_c_3423_n 0.094685f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2239 N_VPWR_c_2830_n N_Z_c_3798_n 4.83404e-19 $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_2240 VPWR N_Z_c_3798_n 0.0135621f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2241 N_VPWR_M1085_d N_Z_c_3424_n 0.001769f $X=10.38 $Y=2.955 $X2=0 $Y2=0
cc_2242 N_VPWR_c_2833_n N_Z_c_3424_n 0.0291114f $X=10.58 $Y=3.13 $X2=0 $Y2=0
cc_2243 VPWR N_Z_c_3424_n 0.094685f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2244 N_VPWR_c_2831_n N_Z_c_3820_n 4.83404e-19 $X=8.51 $Y=3.1 $X2=0 $Y2=0
cc_2245 VPWR N_Z_c_3820_n 0.0135621f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2246 N_VPWR_c_2834_n N_Z_c_3911_n 0.0355595f $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_2247 VPWR N_Z_c_3911_n 0.0739714f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2248 N_VPWR_c_2834_n N_Z_c_3875_n 4.83404e-19 $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_2249 VPWR N_Z_c_3875_n 0.0135621f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2250 N_VPWR_c_2835_n N_Z_c_3921_n 0.0355595f $X=12.65 $Y=3.1 $X2=0 $Y2=0
cc_2251 VPWR N_Z_c_3921_n 0.0739714f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2252 N_VPWR_c_2835_n N_Z_c_3898_n 4.83404e-19 $X=12.65 $Y=3.1 $X2=0 $Y2=0
cc_2253 VPWR N_Z_c_3898_n 0.0135621f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2254 N_VPWR_M1066_d N_Z_c_3425_n 0.001769f $X=14.52 $Y=1.485 $X2=0 $Y2=0
cc_2255 N_VPWR_c_2836_n N_Z_c_3425_n 0.0291114f $X=14.72 $Y=1.63 $X2=0 $Y2=0
cc_2256 VPWR N_Z_c_3425_n 0.094685f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2257 N_VPWR_c_2834_n N_Z_c_3961_n 4.83404e-19 $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_2258 VPWR N_Z_c_3961_n 0.0135621f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2259 N_VPWR_M1072_d N_Z_c_3426_n 0.001769f $X=14.52 $Y=2.955 $X2=0 $Y2=0
cc_2260 N_VPWR_c_2837_n N_Z_c_3426_n 0.0291114f $X=14.72 $Y=3.13 $X2=0 $Y2=0
cc_2261 VPWR N_Z_c_3426_n 0.094685f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2262 N_VPWR_c_2835_n N_Z_c_3983_n 4.83404e-19 $X=12.65 $Y=3.1 $X2=0 $Y2=0
cc_2263 VPWR N_Z_c_3983_n 0.0135621f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2264 N_VPWR_c_2838_n Z 0.00119119f $X=16.76 $Y=1.66 $X2=0 $Y2=0
cc_2265 VPWR Z 0.0135621f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2266 N_VPWR_c_2839_n Z 0.00119119f $X=16.76 $Y=3.1 $X2=0 $Y2=0
cc_2267 VPWR Z 0.0135621f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2268 VPWR N_Z_c_3427_n 0.00481505f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2269 VPWR N_Z_c_3428_n 0.00482221f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2270 N_VPWR_c_2826_n N_Z_c_3429_n 0.00305596f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_2271 VPWR N_Z_c_3429_n 0.00344415f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2272 N_VPWR_c_2827_n N_Z_c_3430_n 0.00305596f $X=4.37 $Y=3.1 $X2=0 $Y2=0
cc_2273 VPWR N_Z_c_3430_n 0.00345131f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2274 N_VPWR_c_2826_n N_Z_c_3431_n 0.00305596f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_2275 VPWR N_Z_c_3431_n 0.00344415f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2276 N_VPWR_c_2827_n N_Z_c_3432_n 0.00305596f $X=4.37 $Y=3.1 $X2=0 $Y2=0
cc_2277 VPWR N_Z_c_3432_n 0.00345131f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2278 N_VPWR_c_2830_n N_Z_c_3433_n 0.00305596f $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_2279 VPWR N_Z_c_3433_n 0.00344415f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2280 N_VPWR_c_2831_n N_Z_c_3434_n 0.00305596f $X=8.51 $Y=3.1 $X2=0 $Y2=0
cc_2281 VPWR N_Z_c_3434_n 0.00345131f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2282 N_VPWR_c_2830_n N_Z_c_3435_n 0.00305596f $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_2283 VPWR N_Z_c_3435_n 0.00344415f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2284 N_VPWR_c_2831_n N_Z_c_3436_n 0.00305596f $X=8.51 $Y=3.1 $X2=0 $Y2=0
cc_2285 VPWR N_Z_c_3436_n 0.00345131f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2286 N_VPWR_c_2834_n N_Z_c_3437_n 0.00305596f $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_2287 VPWR N_Z_c_3437_n 0.00344415f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2288 N_VPWR_c_2835_n N_Z_c_3438_n 0.00305596f $X=12.65 $Y=3.1 $X2=0 $Y2=0
cc_2289 VPWR N_Z_c_3438_n 0.00345131f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2290 N_VPWR_c_2834_n N_Z_c_3439_n 0.00305596f $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_2291 VPWR N_Z_c_3439_n 0.00344415f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2292 N_VPWR_c_2835_n N_Z_c_3440_n 0.00305596f $X=12.65 $Y=3.1 $X2=0 $Y2=0
cc_2293 VPWR N_Z_c_3440_n 0.00345131f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2294 VPWR N_Z_c_3441_n 0.00481505f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2295 VPWR N_Z_c_3442_n 0.00482221f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_2296 VPWR A_734_333# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=1.305
cc_2297 VPWR A_734_591# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=1.305
cc_2298 VPWR A_945_297# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=1.305
cc_2299 VPWR A_945_591# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=1.305
cc_2300 VPWR A_1562_333# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=1.305
cc_2301 VPWR A_1562_591# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=1.305
cc_2302 VPWR A_1773_297# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=1.305
cc_2303 VPWR A_1773_591# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=1.305
cc_2304 VPWR A_2390_333# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=1.305
cc_2305 VPWR A_2390_591# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=1.305
cc_2306 VPWR A_2601_297# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=1.305
cc_2307 VPWR A_2601_591# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=1.305
cc_2308 VPWR A_3218_333# 0.0138589f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=1.305
cc_2309 VPWR A_3218_591# 0.0138589f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=1.305
cc_2310 N_VPWR_c_2822_n N_VGND_c_4368_n 0.00704239f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_2311 N_VPWR_c_2823_n N_VGND_c_4370_n 0.00704239f $X=0.26 $Y=3.1 $X2=0 $Y2=0
cc_2312 N_VPWR_c_2826_n N_VGND_c_4373_n 0.00723368f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_2313 N_VPWR_c_2827_n N_VGND_c_4374_n 0.00723368f $X=4.37 $Y=3.1 $X2=0 $Y2=0
cc_2314 N_VPWR_c_2830_n N_VGND_c_4377_n 0.00723368f $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_2315 N_VPWR_c_2831_n N_VGND_c_4378_n 0.00723368f $X=8.51 $Y=3.1 $X2=0 $Y2=0
cc_2316 N_VPWR_c_2834_n N_VGND_c_4381_n 0.00723368f $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_2317 N_VPWR_c_2835_n N_VGND_c_4382_n 0.00723368f $X=12.65 $Y=3.1 $X2=0 $Y2=0
cc_2318 N_VPWR_c_2838_n N_VGND_c_4386_n 0.00704239f $X=16.76 $Y=1.66 $X2=0 $Y2=0
cc_2319 N_VPWR_c_2839_n N_VGND_c_4388_n 0.00704239f $X=16.76 $Y=3.1 $X2=0 $Y2=0
cc_2320 N_Z_c_3585_n A_734_333# 0.0127078f $X=5.145 $Y=1.87 $X2=-0.19 $Y2=-0.24
cc_2321 N_Z_c_3595_n A_734_591# 0.0127078f $X=5.145 $Y=3.57 $X2=-0.19 $Y2=-0.24
cc_2322 N_Z_c_3585_n A_945_297# 0.0127078f $X=5.145 $Y=1.87 $X2=-0.19 $Y2=-0.24
cc_2323 N_Z_c_3595_n A_945_591# 0.0127078f $X=5.145 $Y=3.57 $X2=-0.19 $Y2=-0.24
cc_2324 N_Z_c_3748_n A_1562_333# 0.0127078f $X=9.285 $Y=1.87 $X2=-0.19 $Y2=-0.24
cc_2325 N_Z_c_3758_n A_1562_591# 0.0127078f $X=9.285 $Y=3.57 $X2=-0.19 $Y2=-0.24
cc_2326 N_Z_c_3748_n A_1773_297# 0.0127078f $X=9.285 $Y=1.87 $X2=-0.19 $Y2=-0.24
cc_2327 N_Z_c_3758_n A_1773_591# 0.0127078f $X=9.285 $Y=3.57 $X2=-0.19 $Y2=-0.24
cc_2328 N_Z_c_3911_n A_2390_333# 0.0127078f $X=13.425 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_2329 N_Z_c_3921_n A_2390_591# 0.0127078f $X=13.425 $Y=3.57 $X2=-0.19
+ $Y2=-0.24
cc_2330 N_Z_c_3911_n A_2601_297# 0.0127078f $X=13.425 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_2331 N_Z_c_3921_n A_2601_591# 0.0127078f $X=13.425 $Y=3.57 $X2=-0.19
+ $Y2=-0.24
cc_2332 N_Z_c_3318_n N_VGND_c_4389_n 0.0106022f $X=1.155 $Y=0.495 $X2=0 $Y2=0
cc_2333 N_Z_c_3320_n N_VGND_c_4391_n 0.0106022f $X=1.155 $Y=4.945 $X2=0 $Y2=0
cc_2334 N_Z_c_3328_n N_VGND_c_4393_n 0.0106022f $X=5.295 $Y=0.495 $X2=0 $Y2=0
cc_2335 N_Z_c_3330_n N_VGND_c_4395_n 0.0106022f $X=5.295 $Y=4.945 $X2=0 $Y2=0
cc_2336 N_Z_c_3338_n N_VGND_c_4397_n 0.0106022f $X=9.435 $Y=0.495 $X2=0 $Y2=0
cc_2337 N_Z_c_3340_n N_VGND_c_4399_n 0.0106022f $X=9.435 $Y=4.945 $X2=0 $Y2=0
cc_2338 N_Z_c_3348_n N_VGND_c_4401_n 0.0106022f $X=13.575 $Y=0.495 $X2=0 $Y2=0
cc_2339 N_Z_c_3350_n N_VGND_c_4403_n 0.0106022f $X=13.575 $Y=4.945 $X2=0 $Y2=0
cc_2340 N_Z_M1092_d VGND 0.00232956f $X=1.02 $Y=0.235 $X2=0 $Y2=0
cc_2341 N_Z_M1023_s VGND 0.00232956f $X=3.32 $Y=0.235 $X2=0 $Y2=0
cc_2342 N_Z_M1018_d VGND 0.00232956f $X=5.16 $Y=0.235 $X2=0 $Y2=0
cc_2343 N_Z_M1015_s VGND 0.00232956f $X=7.46 $Y=0.235 $X2=0 $Y2=0
cc_2344 N_Z_M1030_d VGND 0.00232956f $X=9.3 $Y=0.235 $X2=0 $Y2=0
cc_2345 N_Z_M1020_s VGND 0.00232956f $X=11.6 $Y=0.235 $X2=0 $Y2=0
cc_2346 N_Z_M1063_d VGND 0.00232956f $X=13.44 $Y=0.235 $X2=0 $Y2=0
cc_2347 N_Z_M1060_s VGND 0.00232956f $X=15.74 $Y=0.235 $X2=0 $Y2=0
cc_2348 N_Z_c_3317_n VGND 0.00409585f $X=1.167 $Y=0.835 $X2=0 $Y2=0
cc_2349 N_Z_c_3318_n VGND 0.00891193f $X=1.155 $Y=0.495 $X2=0 $Y2=0
cc_2350 N_Z_c_3321_n VGND 0.00891193f $X=3.445 $Y=0.495 $X2=0 $Y2=0
cc_2351 N_Z_c_3327_n VGND 0.00409585f $X=5.307 $Y=0.835 $X2=0 $Y2=0
cc_2352 N_Z_c_3328_n VGND 0.00891193f $X=5.295 $Y=0.495 $X2=0 $Y2=0
cc_2353 N_Z_c_3331_n VGND 0.00891193f $X=7.585 $Y=0.495 $X2=0 $Y2=0
cc_2354 N_Z_c_3337_n VGND 0.00409585f $X=9.447 $Y=0.835 $X2=0 $Y2=0
cc_2355 N_Z_c_3338_n VGND 0.00891193f $X=9.435 $Y=0.495 $X2=0 $Y2=0
cc_2356 N_Z_c_3341_n VGND 0.00891193f $X=11.725 $Y=0.495 $X2=0 $Y2=0
cc_2357 N_Z_c_3347_n VGND 0.00409585f $X=13.587 $Y=0.835 $X2=0 $Y2=0
cc_2358 N_Z_c_3348_n VGND 0.00891193f $X=13.575 $Y=0.495 $X2=0 $Y2=0
cc_2359 N_Z_c_3351_n VGND 0.00891193f $X=15.865 $Y=0.495 $X2=0 $Y2=0
cc_2360 N_Z_c_3355_n VGND 0.00409585f $X=3.615 $Y=0.92 $X2=0 $Y2=0
cc_2361 N_Z_c_3357_n VGND 0.00409585f $X=7.755 $Y=0.92 $X2=0 $Y2=0
cc_2362 N_Z_c_3359_n VGND 0.00409585f $X=11.895 $Y=0.92 $X2=0 $Y2=0
cc_2363 N_Z_c_3361_n VGND 0.00409585f $X=16.035 $Y=0.92 $X2=0 $Y2=0
cc_2364 N_Z_M1056_d VGND 0.00232956f $X=1.02 $Y=4.685 $X2=0 $Y2=0
cc_2365 N_Z_M1047_s VGND 0.00232956f $X=3.32 $Y=4.685 $X2=0 $Y2=0
cc_2366 N_Z_M1065_d VGND 0.00232956f $X=5.16 $Y=4.685 $X2=0 $Y2=0
cc_2367 N_Z_M1068_s VGND 0.00232956f $X=7.46 $Y=4.685 $X2=0 $Y2=0
cc_2368 N_Z_M1069_d VGND 0.00232956f $X=9.3 $Y=4.685 $X2=0 $Y2=0
cc_2369 N_Z_M1016_s VGND 0.00232956f $X=11.6 $Y=4.685 $X2=0 $Y2=0
cc_2370 N_Z_M1084_d VGND 0.00232956f $X=13.44 $Y=4.685 $X2=0 $Y2=0
cc_2371 N_Z_M1054_s VGND 0.00232956f $X=15.74 $Y=4.685 $X2=0 $Y2=0
cc_2372 N_Z_c_3319_n VGND 0.00410796f $X=1.167 $Y=4.605 $X2=0 $Y2=0
cc_2373 N_Z_c_3320_n VGND 0.00891193f $X=1.155 $Y=4.945 $X2=0 $Y2=0
cc_2374 N_Z_c_3322_n VGND 0.00891193f $X=3.445 $Y=4.945 $X2=0 $Y2=0
cc_2375 N_Z_c_3329_n VGND 0.00410796f $X=5.307 $Y=4.605 $X2=0 $Y2=0
cc_2376 N_Z_c_3330_n VGND 0.00891193f $X=5.295 $Y=4.945 $X2=0 $Y2=0
cc_2377 N_Z_c_3332_n VGND 0.00891193f $X=7.585 $Y=4.945 $X2=0 $Y2=0
cc_2378 N_Z_c_3339_n VGND 0.00410796f $X=9.447 $Y=4.605 $X2=0 $Y2=0
cc_2379 N_Z_c_3340_n VGND 0.00891193f $X=9.435 $Y=4.945 $X2=0 $Y2=0
cc_2380 N_Z_c_3342_n VGND 0.00891193f $X=11.725 $Y=4.945 $X2=0 $Y2=0
cc_2381 N_Z_c_3349_n VGND 0.00410796f $X=13.587 $Y=4.605 $X2=0 $Y2=0
cc_2382 N_Z_c_3350_n VGND 0.00891193f $X=13.575 $Y=4.945 $X2=0 $Y2=0
cc_2383 N_Z_c_3352_n VGND 0.00891193f $X=15.865 $Y=4.945 $X2=0 $Y2=0
cc_2384 N_Z_c_3356_n VGND 0.00410796f $X=3.615 $Y=4.52 $X2=0 $Y2=0
cc_2385 N_Z_c_3358_n VGND 0.00410796f $X=7.755 $Y=4.52 $X2=0 $Y2=0
cc_2386 N_Z_c_3360_n VGND 0.00410796f $X=11.895 $Y=4.52 $X2=0 $Y2=0
cc_2387 N_Z_c_3362_n VGND 0.00410796f $X=16.035 $Y=4.52 $X2=0 $Y2=0
cc_2388 N_Z_c_3321_n N_VGND_c_4407_n 0.0106022f $X=3.445 $Y=0.495 $X2=0 $Y2=0
cc_2389 N_Z_c_3322_n N_VGND_c_4408_n 0.0106022f $X=3.445 $Y=4.945 $X2=0 $Y2=0
cc_2390 N_Z_c_3331_n N_VGND_c_4409_n 0.0106022f $X=7.585 $Y=0.495 $X2=0 $Y2=0
cc_2391 N_Z_c_3332_n N_VGND_c_4410_n 0.0106022f $X=7.585 $Y=4.945 $X2=0 $Y2=0
cc_2392 N_Z_c_3341_n N_VGND_c_4411_n 0.0106022f $X=11.725 $Y=0.495 $X2=0 $Y2=0
cc_2393 N_Z_c_3342_n N_VGND_c_4412_n 0.0106022f $X=11.725 $Y=4.945 $X2=0 $Y2=0
cc_2394 N_Z_c_3351_n N_VGND_c_4413_n 0.0106022f $X=15.865 $Y=0.495 $X2=0 $Y2=0
cc_2395 N_Z_c_3352_n N_VGND_c_4414_n 0.0106022f $X=15.865 $Y=4.945 $X2=0 $Y2=0
cc_2396 VGND A_109_47# 0.00453173f $X=16.705 $Y=-0.085 $X2=-0.19 $Y2=-0.24
cc_2397 VGND A_109_911# 0.00453173f $X=16.705 $Y=5.355 $X2=-0.19 $Y2=-0.24
cc_2398 VGND A_746_47# 0.00453173f $X=16.705 $Y=-0.085 $X2=-0.19 $Y2=-0.24
cc_2399 VGND A_746_937# 0.00453173f $X=16.705 $Y=5.355 $X2=-0.19 $Y2=-0.24
cc_2400 VGND A_937_47# 0.00453173f $X=16.705 $Y=-0.085 $X2=-0.19 $Y2=-0.24
cc_2401 VGND A_937_911# 0.00453173f $X=16.705 $Y=5.355 $X2=-0.19 $Y2=-0.24
cc_2402 VGND A_1574_47# 0.00453173f $X=16.705 $Y=-0.085 $X2=-0.19 $Y2=-0.24
cc_2403 VGND A_1574_937# 0.00453173f $X=16.705 $Y=5.355 $X2=-0.19 $Y2=-0.24
cc_2404 VGND A_1765_47# 0.00453173f $X=16.705 $Y=-0.085 $X2=-0.19 $Y2=-0.24
cc_2405 VGND A_1765_911# 0.00453173f $X=16.705 $Y=5.355 $X2=-0.19 $Y2=-0.24
cc_2406 VGND A_2402_47# 0.00453173f $X=16.705 $Y=-0.085 $X2=-0.19 $Y2=-0.24
cc_2407 VGND A_2402_937# 0.00453173f $X=16.705 $Y=5.355 $X2=-0.19 $Y2=-0.24
cc_2408 VGND A_2593_47# 0.00453173f $X=16.705 $Y=-0.085 $X2=-0.19 $Y2=-0.24
cc_2409 VGND A_2593_911# 0.00453173f $X=16.705 $Y=5.355 $X2=-0.19 $Y2=-0.24
cc_2410 VGND A_3230_47# 0.00453173f $X=16.705 $Y=-0.085 $X2=-0.19 $Y2=-0.24
cc_2411 VGND A_3230_937# 0.00453173f $X=16.705 $Y=5.355 $X2=-0.19 $Y2=-0.24
