* File: sky130_fd_sc_hdll__dlxtn_2.pxi.spice
* Created: Thu Aug 27 19:06:20 2020
* 
x_PM_SKY130_FD_SC_HDLL__DLXTN_2%GATE_N N_GATE_N_c_136_n N_GATE_N_c_137_n
+ N_GATE_N_M1002_g N_GATE_N_c_131_n N_GATE_N_M1015_g N_GATE_N_c_132_n GATE_N
+ GATE_N N_GATE_N_c_134_n N_GATE_N_c_135_n PM_SKY130_FD_SC_HDLL__DLXTN_2%GATE_N
x_PM_SKY130_FD_SC_HDLL__DLXTN_2%A_27_47# N_A_27_47#_M1015_s N_A_27_47#_M1002_s
+ N_A_27_47#_c_182_n N_A_27_47#_c_183_n N_A_27_47#_M1016_g N_A_27_47#_M1000_g
+ N_A_27_47#_M1013_g N_A_27_47#_c_184_n N_A_27_47#_M1005_g N_A_27_47#_c_323_p
+ N_A_27_47#_c_173_n N_A_27_47#_c_174_n N_A_27_47#_c_185_n N_A_27_47#_c_186_n
+ N_A_27_47#_c_187_n N_A_27_47#_c_188_n N_A_27_47#_c_175_n N_A_27_47#_c_176_n
+ N_A_27_47#_c_177_n N_A_27_47#_c_178_n N_A_27_47#_c_190_n N_A_27_47#_c_191_n
+ N_A_27_47#_c_192_n N_A_27_47#_c_193_n N_A_27_47#_c_194_n N_A_27_47#_c_179_n
+ N_A_27_47#_c_180_n N_A_27_47#_c_181_n PM_SKY130_FD_SC_HDLL__DLXTN_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__DLXTN_2%D N_D_c_338_n N_D_c_343_n N_D_M1010_g
+ N_D_M1009_g D N_D_c_340_n N_D_c_341_n PM_SKY130_FD_SC_HDLL__DLXTN_2%D
x_PM_SKY130_FD_SC_HDLL__DLXTN_2%A_319_47# N_A_319_47#_M1009_s
+ N_A_319_47#_M1010_s N_A_319_47#_c_381_n N_A_319_47#_c_389_n
+ N_A_319_47#_M1003_g N_A_319_47#_M1006_g N_A_319_47#_c_390_n
+ N_A_319_47#_c_382_n N_A_319_47#_c_391_n N_A_319_47#_c_392_n
+ N_A_319_47#_c_383_n N_A_319_47#_c_384_n N_A_319_47#_c_385_n
+ N_A_319_47#_c_386_n N_A_319_47#_c_387_n
+ PM_SKY130_FD_SC_HDLL__DLXTN_2%A_319_47#
x_PM_SKY130_FD_SC_HDLL__DLXTN_2%A_211_363# N_A_211_363#_M1000_d
+ N_A_211_363#_M1016_d N_A_211_363#_c_470_n N_A_211_363#_c_475_n
+ N_A_211_363#_c_476_n N_A_211_363#_M1018_g N_A_211_363#_c_471_n
+ N_A_211_363#_M1001_g N_A_211_363#_c_473_n N_A_211_363#_c_479_n
+ N_A_211_363#_c_480_n N_A_211_363#_c_481_n N_A_211_363#_c_482_n
+ N_A_211_363#_c_483_n N_A_211_363#_c_484_n
+ PM_SKY130_FD_SC_HDLL__DLXTN_2%A_211_363#
x_PM_SKY130_FD_SC_HDLL__DLXTN_2%A_783_21# N_A_783_21#_M1014_s
+ N_A_783_21#_M1017_s N_A_783_21#_M1011_g N_A_783_21#_c_588_n
+ N_A_783_21#_M1019_g N_A_783_21#_c_589_n N_A_783_21#_M1004_g
+ N_A_783_21#_c_582_n N_A_783_21#_M1007_g N_A_783_21#_c_590_n
+ N_A_783_21#_M1012_g N_A_783_21#_c_583_n N_A_783_21#_M1008_g
+ N_A_783_21#_c_591_n N_A_783_21#_c_659_p N_A_783_21#_c_628_p
+ N_A_783_21#_c_584_n N_A_783_21#_c_592_n N_A_783_21#_c_585_n
+ N_A_783_21#_c_609_p N_A_783_21#_c_610_p N_A_783_21#_c_611_p
+ N_A_783_21#_c_586_n PM_SKY130_FD_SC_HDLL__DLXTN_2%A_783_21#
x_PM_SKY130_FD_SC_HDLL__DLXTN_2%A_608_413# N_A_608_413#_M1013_d
+ N_A_608_413#_M1018_d N_A_608_413#_c_679_n N_A_608_413#_M1017_g
+ N_A_608_413#_c_673_n N_A_608_413#_M1014_g N_A_608_413#_c_674_n
+ N_A_608_413#_c_675_n N_A_608_413#_c_684_n N_A_608_413#_c_686_n
+ N_A_608_413#_c_676_n N_A_608_413#_c_677_n N_A_608_413#_c_682_n
+ N_A_608_413#_c_678_n PM_SKY130_FD_SC_HDLL__DLXTN_2%A_608_413#
x_PM_SKY130_FD_SC_HDLL__DLXTN_2%VPWR N_VPWR_M1002_d N_VPWR_M1010_d
+ N_VPWR_M1019_d N_VPWR_M1017_d N_VPWR_M1012_d N_VPWR_c_754_n N_VPWR_c_755_n
+ N_VPWR_c_756_n N_VPWR_c_757_n N_VPWR_c_758_n N_VPWR_c_759_n N_VPWR_c_760_n
+ N_VPWR_c_761_n VPWR N_VPWR_c_762_n N_VPWR_c_763_n N_VPWR_c_764_n
+ N_VPWR_c_765_n N_VPWR_c_766_n N_VPWR_c_767_n N_VPWR_c_768_n N_VPWR_c_753_n
+ PM_SKY130_FD_SC_HDLL__DLXTN_2%VPWR
x_PM_SKY130_FD_SC_HDLL__DLXTN_2%Q N_Q_M1007_s N_Q_M1004_s N_Q_c_855_n
+ N_Q_c_862_n N_Q_c_857_n Q Q Q Q PM_SKY130_FD_SC_HDLL__DLXTN_2%Q
x_PM_SKY130_FD_SC_HDLL__DLXTN_2%VGND N_VGND_M1015_d N_VGND_M1009_d
+ N_VGND_M1011_d N_VGND_M1014_d N_VGND_M1008_d N_VGND_c_883_n N_VGND_c_884_n
+ N_VGND_c_885_n N_VGND_c_886_n N_VGND_c_887_n N_VGND_c_888_n VGND
+ N_VGND_c_889_n N_VGND_c_890_n N_VGND_c_891_n N_VGND_c_892_n N_VGND_c_893_n
+ N_VGND_c_894_n N_VGND_c_895_n N_VGND_c_896_n
+ PM_SKY130_FD_SC_HDLL__DLXTN_2%VGND
cc_1 VNB N_GATE_N_c_131_n 0.0173562f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_2 VNB N_GATE_N_c_132_n 0.0272334f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_3 VNB GATE_N 0.0156215f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_GATE_N_c_134_n 0.0217779f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_GATE_N_c_135_n 0.0136718f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_6 VNB N_A_27_47#_M1000_g 0.0409859f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_173_n 0.00233896f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.19
cc_8 VNB N_A_27_47#_c_174_n 0.00643242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_175_n 0.0013847f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_176_n 0.00663785f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_177_n 0.0317895f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_178_n 0.0039153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_179_n 0.0266603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_180_n 0.0184345f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_181_n 0.00490716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_D_c_338_n 0.00677792f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.07
cc_17 VNB N_D_M1009_g 0.0261824f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_18 VNB N_D_c_340_n 0.00715095f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_D_c_341_n 0.0452157f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.665
cc_20 VNB N_A_319_47#_c_381_n 0.014357f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_21 VNB N_A_319_47#_c_382_n 0.00320313f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_22 VNB N_A_319_47#_c_383_n 0.00579201f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_23 VNB N_A_319_47#_c_384_n 0.00340984f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_24 VNB N_A_319_47#_c_385_n 0.00287801f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_25 VNB N_A_319_47#_c_386_n 0.0307009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_319_47#_c_387_n 0.0178076f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_211_363#_c_470_n 0.00625798f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_28 VNB N_A_211_363#_c_471_n 0.0159234f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_211_363#_M1001_g 0.047874f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_211_363#_c_473_n 0.01415f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_31 VNB N_A_783_21#_M1011_g 0.04871f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_32 VNB N_A_783_21#_c_582_n 0.0171483f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.665
cc_33 VNB N_A_783_21#_c_583_n 0.0219903f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_34 VNB N_A_783_21#_c_584_n 0.00259455f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_783_21#_c_585_n 0.00281539f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_783_21#_c_586_n 0.0429675f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_608_413#_c_673_n 0.0198635f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_38 VNB N_A_608_413#_c_674_n 0.0449172f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_39 VNB N_A_608_413#_c_675_n 0.0124501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_608_413#_c_676_n 0.00704689f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_41 VNB N_A_608_413#_c_677_n 0.0119787f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_42 VNB N_A_608_413#_c_678_n 0.00241127f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VPWR_c_753_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_Q_c_855_n 0.00105223f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_45 VNB Q 0.0191317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_883_n 0.0138864f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_884_n 0.00527876f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_885_n 0.00988569f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_49 VNB N_VGND_c_886_n 0.0180189f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_50 VNB N_VGND_c_887_n 0.0463477f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_888_n 0.00606646f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_889_n 0.0154125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_890_n 0.0298657f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_891_n 0.0213492f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_892_n 0.0199476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_893_n 0.0085923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_894_n 0.00859087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_895_n 0.00519339f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_896_n 0.336145f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VPB N_GATE_N_c_136_n 0.0108902f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_61 VPB N_GATE_N_c_137_n 0.0470277f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.74
cc_62 VPB GATE_N 0.0156114f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_63 VPB N_GATE_N_c_134_n 0.0110489f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_64 VPB N_A_27_47#_c_182_n 0.0196311f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_65 VPB N_A_27_47#_c_183_n 0.0261759f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_66 VPB N_A_27_47#_c_184_n 0.0172576f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_67 VPB N_A_27_47#_c_185_n 0.00146141f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_27_47#_c_186_n 0.00585397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_27_47#_c_187_n 0.042255f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_27_47#_c_188_n 0.00363222f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_47#_c_175_n 6.22232e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_47#_c_190_n 0.0253302f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_47#_c_191_n 0.00387417f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_47#_c_192_n 0.00593858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_47#_c_193_n 0.00354884f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_47#_c_194_n 0.00401103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_47#_c_179_n 0.0120947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_47#_c_181_n 3.20024e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_D_c_338_n 0.0240874f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.07
cc_80 VPB N_D_c_343_n 0.0271119f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.4
cc_81 VPB N_D_c_340_n 0.00340154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_319_47#_c_381_n 0.0191152f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_83 VPB N_A_319_47#_c_389_n 0.0225552f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_84 VPB N_A_319_47#_c_390_n 0.00714124f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.665
cc_85 VPB N_A_319_47#_c_391_n 0.00424606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_319_47#_c_392_n 0.00286464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_319_47#_c_384_n 0.00369206f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_88 VPB N_A_211_363#_c_470_n 0.0309494f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_89 VPB N_A_211_363#_c_475_n 0.0108433f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_90 VPB N_A_211_363#_c_476_n 0.024873f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_91 VPB N_A_211_363#_c_471_n 0.0185364f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_211_363#_c_473_n 0.00827089f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_93 VPB N_A_211_363#_c_479_n 0.00300202f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_211_363#_c_480_n 0.00507872f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_95 VPB N_A_211_363#_c_481_n 0.00241696f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_96 VPB N_A_211_363#_c_482_n 0.0071704f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.19
cc_97 VPB N_A_211_363#_c_483_n 0.00114173f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_98 VPB N_A_211_363#_c_484_n 0.0129315f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_783_21#_M1011_g 0.0157901f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_100 VPB N_A_783_21#_c_588_n 0.071851f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_101 VPB N_A_783_21#_c_589_n 0.0162079f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_783_21#_c_590_n 0.020759f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_103 VPB N_A_783_21#_c_591_n 0.00678594f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_104 VPB N_A_783_21#_c_592_n 0.00378052f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_783_21#_c_585_n 0.00281539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_783_21#_c_586_n 0.0258435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_608_413#_c_679_n 0.0193127f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_108 VPB N_A_608_413#_c_674_n 0.0157968f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.805
cc_109 VPB N_A_608_413#_c_675_n 0.00695624f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_608_413#_c_682_n 0.00588113f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_111 VPB N_A_608_413#_c_678_n 0.00221288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_754_n 0.00126291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_755_n 0.00367613f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_756_n 0.00980734f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_115 VPB N_VPWR_c_757_n 0.00199952f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_758_n 0.0100141f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_759_n 0.0329668f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_760_n 0.0326954f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_761_n 0.00446482f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_762_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_763_n 0.0463954f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_764_n 0.019323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_765_n 0.0182359f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_766_n 0.0054556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_767_n 0.00574408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_768_n 0.00398392f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_753_n 0.0587147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_Q_c_857_n 0.00153538f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB Q 0.00612965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 N_GATE_N_c_137_n N_A_27_47#_c_182_n 0.00641193f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_131 N_GATE_N_c_134_n N_A_27_47#_c_182_n 0.00265145f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_132 N_GATE_N_c_137_n N_A_27_47#_c_183_n 0.0182633f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_133 N_GATE_N_c_131_n N_A_27_47#_M1000_g 0.015454f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_134 N_GATE_N_c_135_n N_A_27_47#_M1000_g 0.00178537f $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_135 N_GATE_N_c_131_n N_A_27_47#_c_173_n 0.00633651f $X=0.52 $Y=0.73 $X2=0
+ $Y2=0
cc_136 N_GATE_N_c_132_n N_A_27_47#_c_173_n 0.0136405f $X=0.52 $Y=0.805 $X2=0
+ $Y2=0
cc_137 N_GATE_N_c_132_n N_A_27_47#_c_174_n 0.00657185f $X=0.52 $Y=0.805 $X2=0
+ $Y2=0
cc_138 GATE_N N_A_27_47#_c_174_n 0.0125186f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_139 N_GATE_N_c_134_n N_A_27_47#_c_174_n 3.35813e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_140 N_GATE_N_c_137_n N_A_27_47#_c_185_n 0.0185787f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_141 N_GATE_N_c_137_n N_A_27_47#_c_188_n 0.00836964f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_142 GATE_N N_A_27_47#_c_188_n 0.0139005f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_143 N_GATE_N_c_134_n N_A_27_47#_c_188_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_144 N_GATE_N_c_134_n N_A_27_47#_c_175_n 0.00207629f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_145 N_GATE_N_c_132_n N_A_27_47#_c_176_n 0.00186433f $X=0.52 $Y=0.805 $X2=0
+ $Y2=0
cc_146 GATE_N N_A_27_47#_c_176_n 0.0250709f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_147 N_GATE_N_c_135_n N_A_27_47#_c_176_n 6.20429e-19 $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_148 N_GATE_N_c_136_n N_A_27_47#_c_191_n 0.0015178f $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_149 N_GATE_N_c_137_n N_A_27_47#_c_191_n 0.00103413f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_150 GATE_N N_A_27_47#_c_191_n 0.00630136f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_151 N_GATE_N_c_136_n N_A_27_47#_c_192_n 4.6708e-19 $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_152 N_GATE_N_c_137_n N_A_27_47#_c_192_n 0.00432676f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_153 GATE_N N_A_27_47#_c_179_n 0.00100538f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_154 N_GATE_N_c_134_n N_A_27_47#_c_179_n 0.0129544f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_155 N_GATE_N_c_137_n N_VPWR_c_754_n 0.0125197f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_156 N_GATE_N_c_137_n N_VPWR_c_762_n 0.00304525f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_157 N_GATE_N_c_137_n N_VPWR_c_753_n 0.00454898f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_158 N_GATE_N_c_131_n N_VGND_c_889_n 0.00198377f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_159 N_GATE_N_c_132_n N_VGND_c_889_n 6.41851e-19 $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_160 N_GATE_N_c_131_n N_VGND_c_893_n 0.0142867f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_161 N_GATE_N_c_131_n N_VGND_c_896_n 0.00367064f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_190_n N_D_c_338_n 0.00789696f $X=3.115 $Y=1.53 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_190_n N_D_c_340_n 0.0134197f $X=3.115 $Y=1.53 $X2=0 $Y2=0
cc_164 N_A_27_47#_M1000_g N_D_c_341_n 0.00523969f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_190_n N_A_319_47#_c_381_n 0.00625272f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_c_181_n N_A_319_47#_c_381_n 0.00364423f $X=3.34 $Y=1.415 $X2=0
+ $Y2=0
cc_167 N_A_27_47#_c_190_n N_A_319_47#_c_391_n 0.0135374f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_168 N_A_27_47#_c_190_n N_A_319_47#_c_392_n 0.0114021f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_169 N_A_27_47#_c_177_n N_A_319_47#_c_383_n 9.85912e-19 $X=3 $Y=0.87 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_c_178_n N_A_319_47#_c_383_n 0.013007f $X=3.255 $Y=0.87 $X2=0
+ $Y2=0
cc_171 N_A_27_47#_c_190_n N_A_319_47#_c_383_n 0.00840141f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_172 N_A_27_47#_c_181_n N_A_319_47#_c_383_n 0.00169547f $X=3.34 $Y=1.415 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_c_190_n N_A_319_47#_c_384_n 0.0109087f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_c_177_n N_A_319_47#_c_386_n 0.0120615f $X=3 $Y=0.87 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_c_178_n N_A_319_47#_c_386_n 9.79934e-19 $X=3.255 $Y=0.87 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_c_190_n N_A_319_47#_c_386_n 0.00107604f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_181_n N_A_319_47#_c_386_n 9.89334e-19 $X=3.34 $Y=1.415 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_177_n N_A_319_47#_c_387_n 0.0020564f $X=3 $Y=0.87 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_178_n N_A_319_47#_c_387_n 2.08319e-19 $X=3.255 $Y=0.87 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_180_n N_A_319_47#_c_387_n 0.0199591f $X=3.025 $Y=0.705 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_187_n N_A_211_363#_c_470_n 0.0163374f $X=3.425 $Y=1.74 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_177_n N_A_211_363#_c_470_n 0.0221522f $X=3 $Y=0.87 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_178_n N_A_211_363#_c_470_n 0.0017113f $X=3.255 $Y=0.87 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_190_n N_A_211_363#_c_470_n 0.00674363f $X=3.115 $Y=1.53
+ $X2=0 $Y2=0
cc_185 N_A_27_47#_c_193_n N_A_211_363#_c_470_n 0.00206946f $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_181_n N_A_211_363#_c_470_n 0.00238057f $X=3.34 $Y=1.415
+ $X2=0 $Y2=0
cc_187 N_A_27_47#_c_187_n N_A_211_363#_c_475_n 0.00231825f $X=3.425 $Y=1.74
+ $X2=0 $Y2=0
cc_188 N_A_27_47#_c_194_n N_A_211_363#_c_475_n 0.00238057f $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_184_n N_A_211_363#_c_476_n 0.0170396f $X=3.605 $Y=1.99 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_186_n N_A_211_363#_c_476_n 0.00242155f $X=3.425 $Y=1.74
+ $X2=0 $Y2=0
cc_191 N_A_27_47#_c_187_n N_A_211_363#_c_471_n 0.022219f $X=3.425 $Y=1.74 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_178_n N_A_211_363#_c_471_n 6.84765e-19 $X=3.255 $Y=0.87
+ $X2=0 $Y2=0
cc_193 N_A_27_47#_c_190_n N_A_211_363#_c_471_n 0.00144279f $X=3.115 $Y=1.53
+ $X2=0 $Y2=0
cc_194 N_A_27_47#_c_193_n N_A_211_363#_c_471_n 0.00140497f $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_194_n N_A_211_363#_c_471_n 0.00486358f $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_181_n N_A_211_363#_c_471_n 0.0133603f $X=3.34 $Y=1.415 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_177_n N_A_211_363#_M1001_g 0.0150841f $X=3 $Y=0.87 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_178_n N_A_211_363#_M1001_g 0.00279019f $X=3.255 $Y=0.87
+ $X2=0 $Y2=0
cc_199 N_A_27_47#_c_180_n N_A_211_363#_M1001_g 0.00922417f $X=3.025 $Y=0.705
+ $X2=0 $Y2=0
cc_200 N_A_27_47#_c_181_n N_A_211_363#_M1001_g 0.00479331f $X=3.34 $Y=1.415
+ $X2=0 $Y2=0
cc_201 N_A_27_47#_M1000_g N_A_211_363#_c_473_n 0.0112065f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_173_n N_A_211_363#_c_473_n 0.00937011f $X=0.66 $Y=0.72 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_175_n N_A_211_363#_c_473_n 0.0196553f $X=0.805 $Y=1.235
+ $X2=0 $Y2=0
cc_204 N_A_27_47#_c_176_n N_A_211_363#_c_473_n 0.0138555f $X=0.775 $Y=1.07 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_c_190_n N_A_211_363#_c_473_n 0.0187427f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_191_n N_A_211_363#_c_473_n 0.00220079f $X=0.89 $Y=1.53 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_192_n N_A_211_363#_c_473_n 0.0175551f $X=0.745 $Y=1.53 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_c_182_n N_A_211_363#_c_479_n 0.0112065f $X=0.965 $Y=1.64 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_183_n N_A_211_363#_c_479_n 0.00723076f $X=0.965 $Y=1.74
+ $X2=0 $Y2=0
cc_210 N_A_27_47#_c_185_n N_A_211_363#_c_479_n 0.00387314f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_c_190_n N_A_211_363#_c_479_n 0.00195186f $X=3.115 $Y=1.53
+ $X2=0 $Y2=0
cc_212 N_A_27_47#_c_190_n N_A_211_363#_c_480_n 0.0950762f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_183_n N_A_211_363#_c_481_n 0.00459592f $X=0.965 $Y=1.74
+ $X2=0 $Y2=0
cc_214 N_A_27_47#_c_185_n N_A_211_363#_c_481_n 0.00534864f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_190_n N_A_211_363#_c_481_n 0.0259095f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_192_n N_A_211_363#_c_481_n 0.00107077f $X=0.745 $Y=1.53
+ $X2=0 $Y2=0
cc_217 N_A_27_47#_c_186_n N_A_211_363#_c_483_n 0.00155242f $X=3.425 $Y=1.74
+ $X2=0 $Y2=0
cc_218 N_A_27_47#_c_190_n N_A_211_363#_c_483_n 0.0255946f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_c_187_n N_A_211_363#_c_484_n 3.3276e-19 $X=3.425 $Y=1.74 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_177_n N_A_211_363#_c_484_n 4.0812e-19 $X=3 $Y=0.87 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_c_178_n N_A_211_363#_c_484_n 0.00161882f $X=3.255 $Y=0.87
+ $X2=0 $Y2=0
cc_222 N_A_27_47#_c_190_n N_A_211_363#_c_484_n 0.0245865f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_193_n N_A_211_363#_c_484_n 0.00264902f $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_181_n N_A_211_363#_c_484_n 0.0367681f $X=3.34 $Y=1.415 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_194_n N_A_783_21#_M1011_g 4.94163e-19 $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_181_n N_A_783_21#_M1011_g 2.07812e-19 $X=3.34 $Y=1.415 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_184_n N_A_783_21#_c_588_n 0.0353715f $X=3.605 $Y=1.99 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_c_186_n N_A_783_21#_c_588_n 7.89228e-19 $X=3.425 $Y=1.74 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_c_187_n N_A_783_21#_c_588_n 0.0239253f $X=3.425 $Y=1.74 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_177_n N_A_608_413#_c_684_n 0.00216088f $X=3 $Y=0.87 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_178_n N_A_608_413#_c_684_n 0.0173039f $X=3.255 $Y=0.87 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_184_n N_A_608_413#_c_686_n 0.016617f $X=3.605 $Y=1.99 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_186_n N_A_608_413#_c_686_n 0.0162898f $X=3.425 $Y=1.74 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_187_n N_A_608_413#_c_686_n 0.00113296f $X=3.425 $Y=1.74
+ $X2=0 $Y2=0
cc_235 N_A_27_47#_c_193_n N_A_608_413#_c_686_n 0.00173361f $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_178_n N_A_608_413#_c_676_n 0.0163172f $X=3.255 $Y=0.87 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_c_187_n N_A_608_413#_c_677_n 0.00288725f $X=3.425 $Y=1.74
+ $X2=0 $Y2=0
cc_238 N_A_27_47#_c_178_n N_A_608_413#_c_677_n 0.00245146f $X=3.255 $Y=0.87
+ $X2=0 $Y2=0
cc_239 N_A_27_47#_c_181_n N_A_608_413#_c_677_n 0.0143477f $X=3.34 $Y=1.415 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_c_184_n N_A_608_413#_c_682_n 0.00589555f $X=3.605 $Y=1.99
+ $X2=0 $Y2=0
cc_241 N_A_27_47#_c_187_n N_A_608_413#_c_682_n 0.00302322f $X=3.425 $Y=1.74
+ $X2=0 $Y2=0
cc_242 N_A_27_47#_c_193_n N_A_608_413#_c_682_n 0.00130594f $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_194_n N_A_608_413#_c_682_n 0.0306117f $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_c_181_n N_A_608_413#_c_682_n 0.00322764f $X=3.34 $Y=1.415
+ $X2=0 $Y2=0
cc_245 N_A_27_47#_c_185_n N_VPWR_M1002_d 0.0022997f $X=0.66 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_246 N_A_27_47#_c_183_n N_VPWR_c_754_n 0.00977612f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_185_n N_VPWR_c_754_n 0.0196375f $X=0.66 $Y=1.88 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_188_n N_VPWR_c_754_n 0.0246493f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_249 N_A_27_47#_c_191_n N_VPWR_c_754_n 0.00314061f $X=0.89 $Y=1.53 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_190_n N_VPWR_c_755_n 0.0018348f $X=3.115 $Y=1.53 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_183_n N_VPWR_c_760_n 0.00590576f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_c_185_n N_VPWR_c_762_n 0.00180073f $X=0.66 $Y=1.88 $X2=0 $Y2=0
cc_253 N_A_27_47#_c_188_n N_VPWR_c_762_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_184_n N_VPWR_c_763_n 0.00439333f $X=3.605 $Y=1.99 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_183_n N_VPWR_c_753_n 0.0113647f $X=0.965 $Y=1.74 $X2=0 $Y2=0
cc_256 N_A_27_47#_c_184_n N_VPWR_c_753_n 0.00640904f $X=3.605 $Y=1.99 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_185_n N_VPWR_c_753_n 0.00504362f $X=0.66 $Y=1.88 $X2=0 $Y2=0
cc_258 N_A_27_47#_c_188_n N_VPWR_c_753_n 0.00646745f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_259 N_A_27_47#_c_173_n N_VGND_M1015_d 0.00215196f $X=0.66 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_260 N_A_27_47#_c_177_n N_VGND_c_887_n 0.0013208f $X=3 $Y=0.87 $X2=0 $Y2=0
cc_261 N_A_27_47#_c_178_n N_VGND_c_887_n 0.00248266f $X=3.255 $Y=0.87 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_180_n N_VGND_c_887_n 0.00435108f $X=3.025 $Y=0.705 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_c_323_p N_VGND_c_889_n 0.00725596f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_173_n N_VGND_c_889_n 0.00244154f $X=0.66 $Y=0.72 $X2=0 $Y2=0
cc_265 N_A_27_47#_M1000_g N_VGND_c_890_n 0.00585385f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_M1000_g N_VGND_c_893_n 0.00317372f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_323_p N_VGND_c_893_n 0.00895866f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_268 N_A_27_47#_c_173_n N_VGND_c_893_n 0.0205047f $X=0.66 $Y=0.72 $X2=0 $Y2=0
cc_269 N_A_27_47#_c_175_n N_VGND_c_893_n 0.00148975f $X=0.805 $Y=1.235 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_179_n N_VGND_c_893_n 7.59537e-19 $X=0.99 $Y=1.235 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_M1015_s N_VGND_c_896_n 0.00437169f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_M1000_g N_VGND_c_896_n 0.0120602f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_273 N_A_27_47#_c_323_p N_VGND_c_896_n 0.00608739f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_274 N_A_27_47#_c_173_n N_VGND_c_896_n 0.00595002f $X=0.66 $Y=0.72 $X2=0 $Y2=0
cc_275 N_A_27_47#_c_177_n N_VGND_c_896_n 0.00170666f $X=3 $Y=0.87 $X2=0 $Y2=0
cc_276 N_A_27_47#_c_178_n N_VGND_c_896_n 0.00437549f $X=3.255 $Y=0.87 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_180_n N_VGND_c_896_n 0.0066276f $X=3.025 $Y=0.705 $X2=0
+ $Y2=0
cc_278 N_D_c_341_n N_A_319_47#_c_381_n 0.0145035f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_279 N_D_c_338_n N_A_319_47#_c_389_n 0.0145035f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_280 N_D_c_343_n N_A_319_47#_c_389_n 0.00935018f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_281 N_D_c_343_n N_A_319_47#_c_390_n 0.0136011f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_282 N_D_M1009_g N_A_319_47#_c_382_n 0.0153745f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_283 N_D_c_340_n N_A_319_47#_c_382_n 0.00639931f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_284 N_D_c_341_n N_A_319_47#_c_382_n 0.0029398f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_285 N_D_c_338_n N_A_319_47#_c_391_n 0.0106635f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_286 N_D_c_338_n N_A_319_47#_c_392_n 0.00412429f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_287 N_D_c_340_n N_A_319_47#_c_392_n 0.0233961f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_288 N_D_c_341_n N_A_319_47#_c_392_n 0.00131849f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_289 N_D_M1009_g N_A_319_47#_c_383_n 0.00591272f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_290 N_D_c_340_n N_A_319_47#_c_383_n 0.00920968f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_291 N_D_c_340_n N_A_319_47#_c_384_n 0.013986f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_292 N_D_c_341_n N_A_319_47#_c_384_n 0.0057769f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_293 N_D_M1009_g N_A_319_47#_c_385_n 8.59557e-19 $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_294 N_D_c_340_n N_A_319_47#_c_385_n 0.0138491f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_295 N_D_c_341_n N_A_319_47#_c_385_n 0.0042466f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_296 N_D_M1009_g N_A_319_47#_c_386_n 0.0198512f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_297 N_D_M1009_g N_A_319_47#_c_387_n 0.0127335f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_298 N_D_c_338_n N_A_211_363#_c_473_n 0.00463913f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_299 N_D_M1009_g N_A_211_363#_c_473_n 0.00193515f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_300 N_D_c_340_n N_A_211_363#_c_473_n 0.0287516f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_301 N_D_c_341_n N_A_211_363#_c_473_n 0.00236382f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_302 N_D_c_343_n N_A_211_363#_c_479_n 0.00132248f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_303 N_D_c_343_n N_A_211_363#_c_480_n 0.00420236f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_304 N_D_c_343_n N_VPWR_c_755_n 0.00664063f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_305 N_D_c_343_n N_VPWR_c_760_n 0.00674916f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_306 N_D_c_343_n N_VPWR_c_753_n 0.00848136f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_307 N_D_M1009_g N_VGND_c_890_n 0.00196986f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_308 N_D_M1009_g N_VGND_c_894_n 0.0139983f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_309 N_D_M1009_g N_VGND_c_896_n 0.00398772f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_310 N_D_c_341_n N_VGND_c_896_n 0.00103829f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_311 N_A_319_47#_c_381_n N_A_211_363#_c_470_n 0.0253663f $X=2.425 $Y=1.67
+ $X2=0 $Y2=0
cc_312 N_A_319_47#_c_389_n N_A_211_363#_c_475_n 0.0107827f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_313 N_A_319_47#_c_389_n N_A_211_363#_c_476_n 0.0230246f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_314 N_A_319_47#_c_390_n N_A_211_363#_c_473_n 0.0010921f $X=1.72 $Y=1.99 $X2=0
+ $Y2=0
cc_315 N_A_319_47#_c_392_n N_A_211_363#_c_473_n 0.00880329f $X=1.885 $Y=1.58
+ $X2=0 $Y2=0
cc_316 N_A_319_47#_c_385_n N_A_211_363#_c_473_n 0.0191835f $X=1.72 $Y=0.51 $X2=0
+ $Y2=0
cc_317 N_A_319_47#_c_390_n N_A_211_363#_c_479_n 0.0471073f $X=1.72 $Y=1.99 $X2=0
+ $Y2=0
cc_318 N_A_319_47#_c_389_n N_A_211_363#_c_480_n 0.00505686f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_319 N_A_319_47#_c_390_n N_A_211_363#_c_480_n 0.0230027f $X=1.72 $Y=1.99 $X2=0
+ $Y2=0
cc_320 N_A_319_47#_c_391_n N_A_211_363#_c_480_n 0.00667484f $X=2.12 $Y=1.58
+ $X2=0 $Y2=0
cc_321 N_A_319_47#_c_390_n N_A_211_363#_c_481_n 0.00273055f $X=1.72 $Y=1.99
+ $X2=0 $Y2=0
cc_322 N_A_319_47#_c_389_n N_A_211_363#_c_483_n 0.00149778f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_323 N_A_319_47#_c_381_n N_A_211_363#_c_484_n 0.00472707f $X=2.425 $Y=1.67
+ $X2=0 $Y2=0
cc_324 N_A_319_47#_c_389_n N_A_211_363#_c_484_n 0.00231211f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_325 N_A_319_47#_c_391_n N_A_211_363#_c_484_n 0.00664087f $X=2.12 $Y=1.58
+ $X2=0 $Y2=0
cc_326 N_A_319_47#_c_384_n N_A_211_363#_c_484_n 0.00578855f $X=2.205 $Y=1.495
+ $X2=0 $Y2=0
cc_327 N_A_319_47#_c_389_n N_VPWR_c_755_n 0.0228103f $X=2.425 $Y=1.77 $X2=0
+ $Y2=0
cc_328 N_A_319_47#_c_390_n N_VPWR_c_755_n 0.0355228f $X=1.72 $Y=1.99 $X2=0 $Y2=0
cc_329 N_A_319_47#_c_391_n N_VPWR_c_755_n 0.013562f $X=2.12 $Y=1.58 $X2=0 $Y2=0
cc_330 N_A_319_47#_c_390_n N_VPWR_c_760_n 0.0159613f $X=1.72 $Y=1.99 $X2=0 $Y2=0
cc_331 N_A_319_47#_c_389_n N_VPWR_c_763_n 0.00368966f $X=2.425 $Y=1.77 $X2=0
+ $Y2=0
cc_332 N_A_319_47#_M1010_s N_VPWR_c_753_n 0.00181388f $X=1.595 $Y=1.845 $X2=0
+ $Y2=0
cc_333 N_A_319_47#_c_389_n N_VPWR_c_753_n 0.00385316f $X=2.425 $Y=1.77 $X2=0
+ $Y2=0
cc_334 N_A_319_47#_c_390_n N_VPWR_c_753_n 0.0057885f $X=1.72 $Y=1.99 $X2=0 $Y2=0
cc_335 N_A_319_47#_c_383_n N_VGND_M1009_d 0.00229352f $X=2.205 $Y=1.095 $X2=0
+ $Y2=0
cc_336 N_A_319_47#_c_386_n N_VGND_c_887_n 0.00112938f $X=2.405 $Y=0.93 $X2=0
+ $Y2=0
cc_337 N_A_319_47#_c_387_n N_VGND_c_887_n 0.00585385f $X=2.43 $Y=0.765 $X2=0
+ $Y2=0
cc_338 N_A_319_47#_c_382_n N_VGND_c_890_n 0.00256875f $X=2.12 $Y=0.7 $X2=0 $Y2=0
cc_339 N_A_319_47#_c_385_n N_VGND_c_890_n 0.00723406f $X=1.72 $Y=0.51 $X2=0
+ $Y2=0
cc_340 N_A_319_47#_c_382_n N_VGND_c_894_n 0.00613814f $X=2.12 $Y=0.7 $X2=0 $Y2=0
cc_341 N_A_319_47#_c_383_n N_VGND_c_894_n 0.0161158f $X=2.205 $Y=1.095 $X2=0
+ $Y2=0
cc_342 N_A_319_47#_c_385_n N_VGND_c_894_n 0.00746555f $X=1.72 $Y=0.51 $X2=0
+ $Y2=0
cc_343 N_A_319_47#_c_386_n N_VGND_c_894_n 4.19595e-19 $X=2.405 $Y=0.93 $X2=0
+ $Y2=0
cc_344 N_A_319_47#_c_387_n N_VGND_c_894_n 0.00317372f $X=2.43 $Y=0.765 $X2=0
+ $Y2=0
cc_345 N_A_319_47#_M1009_s N_VGND_c_896_n 0.00343585f $X=1.595 $Y=0.235 $X2=0
+ $Y2=0
cc_346 N_A_319_47#_c_382_n N_VGND_c_896_n 0.0051978f $X=2.12 $Y=0.7 $X2=0 $Y2=0
cc_347 N_A_319_47#_c_383_n N_VGND_c_896_n 0.00710218f $X=2.205 $Y=1.095 $X2=0
+ $Y2=0
cc_348 N_A_319_47#_c_385_n N_VGND_c_896_n 0.00607883f $X=1.72 $Y=0.51 $X2=0
+ $Y2=0
cc_349 N_A_319_47#_c_386_n N_VGND_c_896_n 0.00117722f $X=2.405 $Y=0.93 $X2=0
+ $Y2=0
cc_350 N_A_319_47#_c_387_n N_VGND_c_896_n 0.0064032f $X=2.43 $Y=0.765 $X2=0
+ $Y2=0
cc_351 N_A_211_363#_M1001_g N_A_783_21#_M1011_g 0.0430128f $X=3.515 $Y=0.415
+ $X2=0 $Y2=0
cc_352 N_A_211_363#_M1001_g N_A_608_413#_c_684_n 0.0125662f $X=3.515 $Y=0.415
+ $X2=0 $Y2=0
cc_353 N_A_211_363#_c_476_n N_A_608_413#_c_686_n 0.0054085f $X=2.95 $Y=1.99
+ $X2=0 $Y2=0
cc_354 N_A_211_363#_M1001_g N_A_608_413#_c_676_n 0.00582899f $X=3.515 $Y=0.415
+ $X2=0 $Y2=0
cc_355 N_A_211_363#_M1001_g N_A_608_413#_c_677_n 0.00377136f $X=3.515 $Y=0.415
+ $X2=0 $Y2=0
cc_356 N_A_211_363#_c_471_n N_A_608_413#_c_682_n 7.08904e-19 $X=3.44 $Y=1.32
+ $X2=0 $Y2=0
cc_357 N_A_211_363#_c_480_n N_VPWR_M1010_d 8.51638e-19 $X=2.61 $Y=1.87 $X2=0
+ $Y2=0
cc_358 N_A_211_363#_c_482_n N_VPWR_c_754_n 0.0206383f $X=1.255 $Y=1.87 $X2=0
+ $Y2=0
cc_359 N_A_211_363#_c_476_n N_VPWR_c_755_n 0.003449f $X=2.95 $Y=1.99 $X2=0 $Y2=0
cc_360 N_A_211_363#_c_480_n N_VPWR_c_755_n 0.017675f $X=2.61 $Y=1.87 $X2=0 $Y2=0
cc_361 N_A_211_363#_c_483_n N_VPWR_c_755_n 0.00130564f $X=2.755 $Y=1.87 $X2=0
+ $Y2=0
cc_362 N_A_211_363#_c_484_n N_VPWR_c_755_n 0.00772079f $X=2.87 $Y=1.52 $X2=0
+ $Y2=0
cc_363 N_A_211_363#_c_482_n N_VPWR_c_760_n 0.015988f $X=1.255 $Y=1.87 $X2=0
+ $Y2=0
cc_364 N_A_211_363#_c_476_n N_VPWR_c_763_n 0.00633231f $X=2.95 $Y=1.99 $X2=0
+ $Y2=0
cc_365 N_A_211_363#_c_484_n N_VPWR_c_763_n 0.00457854f $X=2.87 $Y=1.52 $X2=0
+ $Y2=0
cc_366 N_A_211_363#_c_476_n N_VPWR_c_753_n 0.0105199f $X=2.95 $Y=1.99 $X2=0
+ $Y2=0
cc_367 N_A_211_363#_c_480_n N_VPWR_c_753_n 0.0567835f $X=2.61 $Y=1.87 $X2=0
+ $Y2=0
cc_368 N_A_211_363#_c_481_n N_VPWR_c_753_n 0.0152065f $X=1.4 $Y=1.87 $X2=0 $Y2=0
cc_369 N_A_211_363#_c_482_n N_VPWR_c_753_n 0.00389918f $X=1.255 $Y=1.87 $X2=0
+ $Y2=0
cc_370 N_A_211_363#_c_483_n N_VPWR_c_753_n 0.0151073f $X=2.755 $Y=1.87 $X2=0
+ $Y2=0
cc_371 N_A_211_363#_c_484_n N_VPWR_c_753_n 0.00405108f $X=2.87 $Y=1.52 $X2=0
+ $Y2=0
cc_372 N_A_211_363#_c_480_n A_503_369# 0.00150032f $X=2.61 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_373 N_A_211_363#_c_483_n A_503_369# 0.00122092f $X=2.755 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_374 N_A_211_363#_c_484_n A_503_369# 0.0032229f $X=2.87 $Y=1.52 $X2=-0.19
+ $Y2=-0.24
cc_375 N_A_211_363#_M1001_g N_VGND_c_883_n 0.00184584f $X=3.515 $Y=0.415 $X2=0
+ $Y2=0
cc_376 N_A_211_363#_M1001_g N_VGND_c_887_n 0.0037981f $X=3.515 $Y=0.415 $X2=0
+ $Y2=0
cc_377 N_A_211_363#_c_473_n N_VGND_c_890_n 0.00732874f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_378 N_A_211_363#_M1000_d N_VGND_c_896_n 0.00535012f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_379 N_A_211_363#_M1001_g N_VGND_c_896_n 0.00577943f $X=3.515 $Y=0.415 $X2=0
+ $Y2=0
cc_380 N_A_211_363#_c_473_n N_VGND_c_896_n 0.00616598f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_381 N_A_783_21#_c_588_n N_A_608_413#_c_679_n 0.00329184f $X=4.015 $Y=1.99
+ $X2=0 $Y2=0
cc_382 N_A_783_21#_c_589_n N_A_608_413#_c_679_n 0.0193811f $X=5.475 $Y=1.41
+ $X2=0 $Y2=0
cc_383 N_A_783_21#_c_592_n N_A_608_413#_c_679_n 0.00413095f $X=4.82 $Y=1.535
+ $X2=0 $Y2=0
cc_384 N_A_783_21#_c_582_n N_A_608_413#_c_673_n 0.0176547f $X=5.5 $Y=0.995 $X2=0
+ $Y2=0
cc_385 N_A_783_21#_c_584_n N_A_608_413#_c_673_n 0.00635275f $X=4.82 $Y=0.995
+ $X2=0 $Y2=0
cc_386 N_A_783_21#_M1011_g N_A_608_413#_c_674_n 0.01646f $X=3.99 $Y=0.445 $X2=0
+ $Y2=0
cc_387 N_A_783_21#_c_588_n N_A_608_413#_c_674_n 0.00487525f $X=4.015 $Y=1.99
+ $X2=0 $Y2=0
cc_388 N_A_783_21#_c_591_n N_A_608_413#_c_674_n 0.00879412f $X=4.685 $Y=1.7
+ $X2=0 $Y2=0
cc_389 N_A_783_21#_c_609_p N_A_608_413#_c_674_n 0.00203472f $X=4.795 $Y=0.825
+ $X2=0 $Y2=0
cc_390 N_A_783_21#_c_610_p N_A_608_413#_c_674_n 0.00212837f $X=4.77 $Y=1.755
+ $X2=0 $Y2=0
cc_391 N_A_783_21#_c_611_p N_A_608_413#_c_674_n 0.0181912f $X=4.82 $Y=1.16 $X2=0
+ $Y2=0
cc_392 N_A_783_21#_c_592_n N_A_608_413#_c_675_n 0.0036022f $X=4.82 $Y=1.535
+ $X2=0 $Y2=0
cc_393 N_A_783_21#_c_585_n N_A_608_413#_c_675_n 0.0276191f $X=5.45 $Y=1.16 $X2=0
+ $Y2=0
cc_394 N_A_783_21#_c_586_n N_A_608_413#_c_675_n 0.0256136f $X=5.945 $Y=1.202
+ $X2=0 $Y2=0
cc_395 N_A_783_21#_M1011_g N_A_608_413#_c_684_n 0.00149885f $X=3.99 $Y=0.445
+ $X2=0 $Y2=0
cc_396 N_A_783_21#_c_588_n N_A_608_413#_c_686_n 0.00398626f $X=4.015 $Y=1.99
+ $X2=0 $Y2=0
cc_397 N_A_783_21#_M1011_g N_A_608_413#_c_676_n 0.00598699f $X=3.99 $Y=0.445
+ $X2=0 $Y2=0
cc_398 N_A_783_21#_M1011_g N_A_608_413#_c_677_n 0.00570022f $X=3.99 $Y=0.445
+ $X2=0 $Y2=0
cc_399 N_A_783_21#_M1011_g N_A_608_413#_c_682_n 0.0114233f $X=3.99 $Y=0.445
+ $X2=0 $Y2=0
cc_400 N_A_783_21#_c_588_n N_A_608_413#_c_682_n 0.0238269f $X=4.015 $Y=1.99
+ $X2=0 $Y2=0
cc_401 N_A_783_21#_c_591_n N_A_608_413#_c_682_n 0.019033f $X=4.685 $Y=1.7 $X2=0
+ $Y2=0
cc_402 N_A_783_21#_M1011_g N_A_608_413#_c_678_n 0.0176525f $X=3.99 $Y=0.445
+ $X2=0 $Y2=0
cc_403 N_A_783_21#_c_588_n N_A_608_413#_c_678_n 0.00820473f $X=4.015 $Y=1.99
+ $X2=0 $Y2=0
cc_404 N_A_783_21#_c_591_n N_A_608_413#_c_678_n 0.02399f $X=4.685 $Y=1.7 $X2=0
+ $Y2=0
cc_405 N_A_783_21#_c_611_p N_A_608_413#_c_678_n 0.0253721f $X=4.82 $Y=1.16 $X2=0
+ $Y2=0
cc_406 N_A_783_21#_c_588_n N_VPWR_c_756_n 0.012526f $X=4.015 $Y=1.99 $X2=0 $Y2=0
cc_407 N_A_783_21#_c_591_n N_VPWR_c_756_n 0.0154822f $X=4.685 $Y=1.7 $X2=0 $Y2=0
cc_408 N_A_783_21#_c_628_p N_VPWR_c_756_n 0.0196385f $X=4.77 $Y=2.27 $X2=0 $Y2=0
cc_409 N_A_783_21#_c_589_n N_VPWR_c_757_n 0.0189852f $X=5.475 $Y=1.41 $X2=0
+ $Y2=0
cc_410 N_A_783_21#_c_590_n N_VPWR_c_757_n 0.00140703f $X=5.945 $Y=1.41 $X2=0
+ $Y2=0
cc_411 N_A_783_21#_c_585_n N_VPWR_c_757_n 0.0195387f $X=5.45 $Y=1.16 $X2=0 $Y2=0
cc_412 N_A_783_21#_c_586_n N_VPWR_c_757_n 0.00125453f $X=5.945 $Y=1.202 $X2=0
+ $Y2=0
cc_413 N_A_783_21#_c_590_n N_VPWR_c_759_n 0.00831633f $X=5.945 $Y=1.41 $X2=0
+ $Y2=0
cc_414 N_A_783_21#_c_588_n N_VPWR_c_763_n 0.00694824f $X=4.015 $Y=1.99 $X2=0
+ $Y2=0
cc_415 N_A_783_21#_c_628_p N_VPWR_c_764_n 0.0115253f $X=4.77 $Y=2.27 $X2=0 $Y2=0
cc_416 N_A_783_21#_c_589_n N_VPWR_c_765_n 0.00622633f $X=5.475 $Y=1.41 $X2=0
+ $Y2=0
cc_417 N_A_783_21#_c_590_n N_VPWR_c_765_n 0.00621235f $X=5.945 $Y=1.41 $X2=0
+ $Y2=0
cc_418 N_A_783_21#_M1017_s N_VPWR_c_753_n 0.00284579f $X=4.645 $Y=1.485 $X2=0
+ $Y2=0
cc_419 N_A_783_21#_c_588_n N_VPWR_c_753_n 0.01438f $X=4.015 $Y=1.99 $X2=0 $Y2=0
cc_420 N_A_783_21#_c_589_n N_VPWR_c_753_n 0.0104011f $X=5.475 $Y=1.41 $X2=0
+ $Y2=0
cc_421 N_A_783_21#_c_590_n N_VPWR_c_753_n 0.0114615f $X=5.945 $Y=1.41 $X2=0
+ $Y2=0
cc_422 N_A_783_21#_c_591_n N_VPWR_c_753_n 0.00898578f $X=4.685 $Y=1.7 $X2=0
+ $Y2=0
cc_423 N_A_783_21#_c_628_p N_VPWR_c_753_n 0.00827281f $X=4.77 $Y=2.27 $X2=0
+ $Y2=0
cc_424 N_A_783_21#_c_582_n N_Q_c_855_n 0.00358785f $X=5.5 $Y=0.995 $X2=0 $Y2=0
cc_425 N_A_783_21#_c_583_n N_Q_c_855_n 0.00805744f $X=5.97 $Y=0.995 $X2=0 $Y2=0
cc_426 N_A_783_21#_c_586_n N_Q_c_855_n 0.00232072f $X=5.945 $Y=1.202 $X2=0 $Y2=0
cc_427 N_A_783_21#_c_589_n N_Q_c_862_n 0.00469231f $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_428 N_A_783_21#_c_590_n N_Q_c_862_n 0.0078022f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_429 N_A_783_21#_c_586_n N_Q_c_862_n 0.00359264f $X=5.945 $Y=1.202 $X2=0 $Y2=0
cc_430 N_A_783_21#_c_589_n N_Q_c_857_n 0.00174751f $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_431 N_A_783_21#_c_590_n N_Q_c_857_n 0.00414246f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_432 N_A_783_21#_c_586_n N_Q_c_857_n 0.00923077f $X=5.945 $Y=1.202 $X2=0 $Y2=0
cc_433 N_A_783_21#_c_583_n Q 0.0136435f $X=5.97 $Y=0.995 $X2=0 $Y2=0
cc_434 N_A_783_21#_c_586_n Q 0.00217272f $X=5.945 $Y=1.202 $X2=0 $Y2=0
cc_435 N_A_783_21#_c_590_n Q 0.0161201f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_436 N_A_783_21#_c_585_n Q 0.0236524f $X=5.45 $Y=1.16 $X2=0 $Y2=0
cc_437 N_A_783_21#_c_586_n Q 0.0355201f $X=5.945 $Y=1.202 $X2=0 $Y2=0
cc_438 N_A_783_21#_M1011_g N_VGND_c_883_n 0.0188178f $X=3.99 $Y=0.445 $X2=0
+ $Y2=0
cc_439 N_A_783_21#_c_659_p N_VGND_c_883_n 0.0236254f $X=4.77 $Y=0.58 $X2=0 $Y2=0
cc_440 N_A_783_21#_c_582_n N_VGND_c_884_n 0.00408035f $X=5.5 $Y=0.995 $X2=0
+ $Y2=0
cc_441 N_A_783_21#_c_585_n N_VGND_c_884_n 0.0200847f $X=5.45 $Y=1.16 $X2=0 $Y2=0
cc_442 N_A_783_21#_c_586_n N_VGND_c_884_n 0.00204942f $X=5.945 $Y=1.202 $X2=0
+ $Y2=0
cc_443 N_A_783_21#_c_583_n N_VGND_c_886_n 0.00450677f $X=5.97 $Y=0.995 $X2=0
+ $Y2=0
cc_444 N_A_783_21#_M1011_g N_VGND_c_887_n 0.0046653f $X=3.99 $Y=0.445 $X2=0
+ $Y2=0
cc_445 N_A_783_21#_c_659_p N_VGND_c_891_n 0.00732441f $X=4.77 $Y=0.58 $X2=0
+ $Y2=0
cc_446 N_A_783_21#_c_582_n N_VGND_c_892_n 0.00585385f $X=5.5 $Y=0.995 $X2=0
+ $Y2=0
cc_447 N_A_783_21#_c_583_n N_VGND_c_892_n 0.00567045f $X=5.97 $Y=0.995 $X2=0
+ $Y2=0
cc_448 N_A_783_21#_M1014_s N_VGND_c_896_n 0.00589711f $X=4.645 $Y=0.235 $X2=0
+ $Y2=0
cc_449 N_A_783_21#_M1011_g N_VGND_c_896_n 0.00813035f $X=3.99 $Y=0.445 $X2=0
+ $Y2=0
cc_450 N_A_783_21#_c_582_n N_VGND_c_896_n 0.0108962f $X=5.5 $Y=0.995 $X2=0 $Y2=0
cc_451 N_A_783_21#_c_583_n N_VGND_c_896_n 0.0111951f $X=5.97 $Y=0.995 $X2=0
+ $Y2=0
cc_452 N_A_783_21#_c_659_p N_VGND_c_896_n 0.00762661f $X=4.77 $Y=0.58 $X2=0
+ $Y2=0
cc_453 N_A_608_413#_c_679_n N_VPWR_c_756_n 0.00253117f $X=5.005 $Y=1.41 $X2=0
+ $Y2=0
cc_454 N_A_608_413#_c_686_n N_VPWR_c_756_n 0.0113935f $X=3.775 $Y=2.34 $X2=0
+ $Y2=0
cc_455 N_A_608_413#_c_682_n N_VPWR_c_756_n 0.00720228f $X=3.86 $Y=2.255 $X2=0
+ $Y2=0
cc_456 N_A_608_413#_c_679_n N_VPWR_c_757_n 0.0027968f $X=5.005 $Y=1.41 $X2=0
+ $Y2=0
cc_457 N_A_608_413#_c_686_n N_VPWR_c_763_n 0.0368884f $X=3.775 $Y=2.34 $X2=0
+ $Y2=0
cc_458 N_A_608_413#_c_679_n N_VPWR_c_764_n 0.00702461f $X=5.005 $Y=1.41 $X2=0
+ $Y2=0
cc_459 N_A_608_413#_M1018_d N_VPWR_c_753_n 0.00724737f $X=3.04 $Y=2.065 $X2=0
+ $Y2=0
cc_460 N_A_608_413#_c_679_n N_VPWR_c_753_n 0.0138941f $X=5.005 $Y=1.41 $X2=0
+ $Y2=0
cc_461 N_A_608_413#_c_686_n N_VPWR_c_753_n 0.0283655f $X=3.775 $Y=2.34 $X2=0
+ $Y2=0
cc_462 N_A_608_413#_c_686_n A_739_413# 0.00204526f $X=3.775 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_463 N_A_608_413#_c_682_n A_739_413# 0.00209205f $X=3.86 $Y=2.255 $X2=-0.19
+ $Y2=-0.24
cc_464 N_A_608_413#_c_673_n N_VGND_c_883_n 0.00699752f $X=5.03 $Y=0.995 $X2=0
+ $Y2=0
cc_465 N_A_608_413#_c_674_n N_VGND_c_883_n 0.00207331f $X=4.905 $Y=1.16 $X2=0
+ $Y2=0
cc_466 N_A_608_413#_c_684_n N_VGND_c_883_n 0.0109093f $X=3.625 $Y=0.45 $X2=0
+ $Y2=0
cc_467 N_A_608_413#_c_676_n N_VGND_c_883_n 0.0168172f $X=3.71 $Y=0.995 $X2=0
+ $Y2=0
cc_468 N_A_608_413#_c_678_n N_VGND_c_883_n 0.0328206f $X=4.46 $Y=1.16 $X2=0
+ $Y2=0
cc_469 N_A_608_413#_c_673_n N_VGND_c_884_n 0.00400015f $X=5.03 $Y=0.995 $X2=0
+ $Y2=0
cc_470 N_A_608_413#_c_684_n N_VGND_c_887_n 0.0243846f $X=3.625 $Y=0.45 $X2=0
+ $Y2=0
cc_471 N_A_608_413#_c_673_n N_VGND_c_891_n 0.00585385f $X=5.03 $Y=0.995 $X2=0
+ $Y2=0
cc_472 N_A_608_413#_M1013_d N_VGND_c_896_n 0.00327132f $X=3.065 $Y=0.235 $X2=0
+ $Y2=0
cc_473 N_A_608_413#_c_673_n N_VGND_c_896_n 0.0121665f $X=5.03 $Y=0.995 $X2=0
+ $Y2=0
cc_474 N_A_608_413#_c_684_n N_VGND_c_896_n 0.0241568f $X=3.625 $Y=0.45 $X2=0
+ $Y2=0
cc_475 N_A_608_413#_c_684_n A_718_47# 0.00369918f $X=3.625 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_476 N_A_608_413#_c_676_n A_718_47# 0.00128174f $X=3.71 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_477 N_VPWR_c_753_n A_503_369# 0.00393797f $X=6.21 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_478 N_VPWR_c_753_n A_739_413# 0.00186708f $X=6.21 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_479 N_VPWR_c_753_n N_Q_M1004_s 0.00439839f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_480 N_VPWR_c_757_n N_Q_c_862_n 0.0595171f $X=5.24 $Y=1.735 $X2=0 $Y2=0
cc_481 N_VPWR_c_759_n Q 0.0492906f $X=6.18 $Y=2 $X2=0 $Y2=0
cc_482 N_VPWR_c_765_n Q 0.0166993f $X=6.095 $Y=2.72 $X2=0 $Y2=0
cc_483 N_VPWR_c_753_n Q 0.0105267f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_484 N_VPWR_c_759_n Q 0.0111243f $X=6.18 $Y=2 $X2=0 $Y2=0
cc_485 Q N_VGND_c_886_n 0.0107109f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_486 Q N_VGND_c_892_n 0.00849755f $X=5.68 $Y=0.425 $X2=0 $Y2=0
cc_487 N_Q_M1007_s N_VGND_c_896_n 0.00457716f $X=5.575 $Y=0.235 $X2=0 $Y2=0
cc_488 Q N_VGND_c_896_n 0.00975124f $X=5.68 $Y=0.425 $X2=0 $Y2=0
cc_489 N_VGND_c_896_n A_505_47# 0.0139156f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_490 N_VGND_c_896_n A_718_47# 0.00687059f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
