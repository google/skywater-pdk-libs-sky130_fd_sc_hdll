* File: sky130_fd_sc_hdll__o211a_4.pex.spice
* Created: Wed Sep  2 08:42:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O211A_4%A_80_21# 1 2 3 4 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 37 44 46 48 49 51 53 54 57 59 63 65 69 70 71 73
c161 70 0 1.2412e-19 $X=3.18 $Y=1.94
c162 44 0 1.11396e-19 $X=2.26 $Y=1.16
c163 34 0 3.24388e-20 $X=2.38 $Y=1.41
r164 80 81 1.99724 $w=3.62e-07 $l=1.5e-08 $layer=POLY_cond $X=1.885 $Y=1.202
+ $X2=1.9 $Y2=1.202
r165 79 80 61.9144 $w=3.62e-07 $l=4.65e-07 $layer=POLY_cond $X=1.42 $Y=1.202
+ $X2=1.885 $Y2=1.202
r166 78 79 0.665746 $w=3.62e-07 $l=5e-09 $layer=POLY_cond $X=1.415 $Y=1.202
+ $X2=1.42 $Y2=1.202
r167 77 78 62.5801 $w=3.62e-07 $l=4.7e-07 $layer=POLY_cond $X=0.945 $Y=1.202
+ $X2=1.415 $Y2=1.202
r168 76 77 0.665746 $w=3.62e-07 $l=5e-09 $layer=POLY_cond $X=0.94 $Y=1.202
+ $X2=0.945 $Y2=1.202
r169 66 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.415 $Y=1.94
+ $X2=4.25 $Y2=1.94
r170 65 73 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.465 $Y=1.94
+ $X2=5.655 $Y2=1.94
r171 65 66 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=5.465 $Y=1.94
+ $X2=4.415 $Y2=1.94
r172 61 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.25 $Y=2.025
+ $X2=4.25 $Y2=1.94
r173 61 63 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.25 $Y=2.025
+ $X2=4.25 $Y2=2.3
r174 60 70 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.36 $Y=1.94
+ $X2=3.18 $Y2=1.94
r175 59 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.085 $Y=1.94
+ $X2=4.25 $Y2=1.94
r176 59 60 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=4.085 $Y=1.94
+ $X2=3.36 $Y2=1.94
r177 55 70 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.18 $Y=2.025
+ $X2=3.18 $Y2=1.94
r178 55 57 8.80338 $w=3.58e-07 $l=2.75e-07 $layer=LI1_cond $X=3.18 $Y=2.025
+ $X2=3.18 $Y2=2.3
r179 53 70 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3 $Y=1.94 $X2=3.18
+ $Y2=1.94
r180 53 54 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3 $Y=1.94 $X2=2.62
+ $Y2=1.94
r181 49 51 60.6919 $w=1.78e-07 $l=9.85e-07 $layer=LI1_cond $X=2.62 $Y=0.725
+ $X2=3.605 $Y2=0.725
r182 48 54 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.51 $Y=1.855
+ $X2=2.62 $Y2=1.94
r183 47 69 4.76867 $w=2.2e-07 $l=1e-07 $layer=LI1_cond $X=2.51 $Y=1.265 $X2=2.51
+ $Y2=1.165
r184 47 48 30.9064 $w=2.18e-07 $l=5.9e-07 $layer=LI1_cond $X=2.51 $Y=1.265
+ $X2=2.51 $Y2=1.855
r185 46 69 4.76867 $w=2.2e-07 $l=1e-07 $layer=LI1_cond $X=2.51 $Y=1.065 $X2=2.51
+ $Y2=1.165
r186 45 49 6.90553 $w=1.8e-07 $l=1.48324e-07 $layer=LI1_cond $X=2.51 $Y=0.815
+ $X2=2.62 $Y2=0.725
r187 45 46 13.0959 $w=2.18e-07 $l=2.5e-07 $layer=LI1_cond $X=2.51 $Y=0.815
+ $X2=2.51 $Y2=1.065
r188 44 83 15.9779 $w=3.62e-07 $l=1.2e-07 $layer=POLY_cond $X=2.26 $Y=1.202
+ $X2=2.38 $Y2=1.202
r189 44 81 47.9337 $w=3.62e-07 $l=3.6e-07 $layer=POLY_cond $X=2.26 $Y=1.202
+ $X2=1.9 $Y2=1.202
r190 43 44 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.26
+ $Y=1.16 $X2=2.26 $Y2=1.16
r191 40 76 25.2983 $w=3.62e-07 $l=1.9e-07 $layer=POLY_cond $X=0.75 $Y=1.202
+ $X2=0.94 $Y2=1.202
r192 40 74 36.616 $w=3.62e-07 $l=2.75e-07 $layer=POLY_cond $X=0.75 $Y=1.202
+ $X2=0.475 $Y2=1.202
r193 39 43 83.7364 $w=1.98e-07 $l=1.51e-06 $layer=LI1_cond $X=0.75 $Y=1.165
+ $X2=2.26 $Y2=1.165
r194 39 40 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.75
+ $Y=1.16 $X2=0.75 $Y2=1.16
r195 37 69 1.68792 $w=2e-07 $l=1.1e-07 $layer=LI1_cond $X=2.4 $Y=1.165 $X2=2.51
+ $Y2=1.165
r196 37 43 7.76364 $w=1.98e-07 $l=1.4e-07 $layer=LI1_cond $X=2.4 $Y=1.165
+ $X2=2.26 $Y2=1.165
r197 34 83 19.0988 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.38 $Y=1.41
+ $X2=2.38 $Y2=1.202
r198 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.38 $Y=1.41
+ $X2=2.38 $Y2=1.985
r199 31 81 19.0988 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.9 $Y=1.41
+ $X2=1.9 $Y2=1.202
r200 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.9 $Y=1.41
+ $X2=1.9 $Y2=1.985
r201 28 80 23.4391 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.885 $Y=0.995
+ $X2=1.885 $Y2=1.202
r202 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.885 $Y=0.995
+ $X2=1.885 $Y2=0.56
r203 25 78 23.4391 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.415 $Y=0.995
+ $X2=1.415 $Y2=1.202
r204 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.415 $Y=0.995
+ $X2=1.415 $Y2=0.56
r205 22 79 19.0988 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.42 $Y=1.41
+ $X2=1.42 $Y2=1.202
r206 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.42 $Y=1.41
+ $X2=1.42 $Y2=1.985
r207 19 77 23.4391 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.945 $Y=0.995
+ $X2=0.945 $Y2=1.202
r208 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.945 $Y=0.995
+ $X2=0.945 $Y2=0.56
r209 16 76 19.0988 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.94 $Y=1.41
+ $X2=0.94 $Y2=1.202
r210 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.94 $Y=1.41
+ $X2=0.94 $Y2=1.985
r211 13 74 23.4391 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=1.202
r212 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=0.56
r213 4 73 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=5.53
+ $Y=1.485 $X2=5.68 $Y2=2.02
r214 3 63 600 $w=1.7e-07 $l=8.95977e-07 $layer=licon1_PDIFF $count=1 $X=4.08
+ $Y=1.485 $X2=4.25 $Y2=2.3
r215 2 57 600 $w=1.7e-07 $l=9.31652e-07 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.485 $X2=3.195 $Y2=2.3
r216 1 51 182 $w=1.7e-07 $l=5.90741e-07 $layer=licon1_NDIFF $count=1 $X=3.395
+ $Y=0.235 $X2=3.605 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_4%B1 1 3 4 6 7 9 10 12 15 18 19 26
c84 15 0 3.24388e-20 $X=2.875 $Y=1.16
c85 1 0 1.2412e-19 $X=2.855 $Y=1.41
r86 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.435
+ $Y=1.16 $X2=4.435 $Y2=1.16
r87 19 26 8.20134 $w=4.98e-07 $l=2.85e-07 $layer=LI1_cond $X=4.435 $Y=1.445
+ $X2=4.435 $Y2=1.16
r88 18 19 34.5455 $w=4.08e-07 $l=1.185e-06 $layer=LI1_cond $X=3.085 $Y=1.565
+ $X2=4.27 $Y2=1.565
r89 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.875
+ $Y=1.16 $X2=2.875 $Y2=1.16
r90 13 18 6.91061 $w=2.4e-07 $l=1.99158e-07 $layer=LI1_cond $X=2.937 $Y=1.445
+ $X2=3.085 $Y2=1.565
r91 13 15 11.1338 $w=2.93e-07 $l=2.85e-07 $layer=LI1_cond $X=2.937 $Y=1.445
+ $X2=2.937 $Y2=1.16
r92 10 25 50.2707 $w=2.67e-07 $l=2.70647e-07 $layer=POLY_cond $X=4.485 $Y=1.41
+ $X2=4.442 $Y2=1.16
r93 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.485 $Y=1.41
+ $X2=4.485 $Y2=1.985
r94 7 25 38.9672 $w=2.67e-07 $l=1.84811e-07 $layer=POLY_cond $X=4.4 $Y=0.995
+ $X2=4.442 $Y2=1.16
r95 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.4 $Y=0.995 $X2=4.4
+ $Y2=0.56
r96 4 16 38.8084 $w=2.75e-07 $l=1.98167e-07 $layer=POLY_cond $X=2.96 $Y=0.995
+ $X2=2.887 $Y2=1.16
r97 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.96 $Y=0.995 $X2=2.96
+ $Y2=0.56
r98 1 16 49.5676 $w=2.75e-07 $l=2.65518e-07 $layer=POLY_cond $X=2.855 $Y=1.41
+ $X2=2.887 $Y2=1.16
r99 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.855 $Y=1.41
+ $X2=2.855 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_4%C1 1 3 4 6 7 9 10 12 13 19 20 25
r47 20 21 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=3.99 $Y=1.202
+ $X2=4.015 $Y2=1.202
r48 19 25 20.6479 $w=2.38e-07 $l=4.3e-07 $layer=LI1_cond $X=3.875 $Y=1.155
+ $X2=3.445 $Y2=1.155
r49 18 20 14.9811 $w=3.7e-07 $l=1.15e-07 $layer=POLY_cond $X=3.875 $Y=1.202
+ $X2=3.99 $Y2=1.202
r50 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.875
+ $Y=1.16 $X2=3.875 $Y2=1.16
r51 16 18 47.5486 $w=3.7e-07 $l=3.65e-07 $layer=POLY_cond $X=3.51 $Y=1.202
+ $X2=3.875 $Y2=1.202
r52 15 16 24.7514 $w=3.7e-07 $l=1.9e-07 $layer=POLY_cond $X=3.32 $Y=1.202
+ $X2=3.51 $Y2=1.202
r53 13 25 0.240092 $w=2.38e-07 $l=5e-09 $layer=LI1_cond $X=3.44 $Y=1.155
+ $X2=3.445 $Y2=1.155
r54 10 21 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.015 $Y=0.995
+ $X2=4.015 $Y2=1.202
r55 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.015 $Y=0.995
+ $X2=4.015 $Y2=0.56
r56 7 20 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.99 $Y=1.41
+ $X2=3.99 $Y2=1.202
r57 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.99 $Y=1.41 $X2=3.99
+ $Y2=1.985
r58 4 16 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.51 $Y=1.41
+ $X2=3.51 $Y2=1.202
r59 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.51 $Y=1.41 $X2=3.51
+ $Y2=1.985
r60 1 15 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.32 $Y=0.995
+ $X2=3.32 $Y2=1.202
r61 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.32 $Y=0.995 $X2=3.32
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_4%A1 1 3 4 6 7 9 10 12 15 18 19 20 25
c73 15 0 1.15076e-19 $X=4.99 $Y=1.16
c74 1 0 6.40318e-20 $X=4.875 $Y=0.995
r75 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.495
+ $Y=1.16 $X2=6.495 $Y2=1.16
r76 20 25 8.59318 $w=5.13e-07 $l=3.7e-07 $layer=LI1_cond $X=6.557 $Y=1.53
+ $X2=6.557 $Y2=1.16
r77 18 20 1.39349 $w=5.13e-07 $l=6e-08 $layer=LI1_cond $X=6.557 $Y=1.59
+ $X2=6.557 $Y2=1.53
r78 18 19 66.8373 $w=1.88e-07 $l=1.145e-06 $layer=LI1_cond $X=6.3 $Y=1.59
+ $X2=5.155 $Y2=1.59
r79 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.99
+ $Y=1.16 $X2=4.99 $Y2=1.16
r80 13 19 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=4.99 $Y=1.495
+ $X2=5.155 $Y2=1.59
r81 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.99 $Y=1.495
+ $X2=4.99 $Y2=1.16
r82 10 24 44.909 $w=3.98e-07 $l=3.06186e-07 $layer=POLY_cond $X=6.4 $Y=1.41
+ $X2=6.525 $Y2=1.16
r83 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.4 $Y=1.41 $X2=6.4
+ $Y2=1.985
r84 7 24 39.5463 $w=3.98e-07 $l=2.2798e-07 $layer=POLY_cond $X=6.375 $Y=0.995
+ $X2=6.525 $Y2=1.16
r85 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.375 $Y=0.995
+ $X2=6.375 $Y2=0.56
r86 4 16 47.6478 $w=3.03e-07 $l=2.52488e-07 $layer=POLY_cond $X=4.96 $Y=1.41
+ $X2=4.965 $Y2=1.16
r87 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.96 $Y=1.41 $X2=4.96
+ $Y2=1.985
r88 1 16 38.5416 $w=3.03e-07 $l=2.05122e-07 $layer=POLY_cond $X=4.875 $Y=0.995
+ $X2=4.965 $Y2=1.16
r89 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.875 $Y=0.995
+ $X2=4.875 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_4%A2 1 3 4 6 7 9 10 12 13 18 19 22
r53 18 20 3.21333 $w=3.75e-07 $l=2.5e-08 $layer=POLY_cond $X=5.895 $Y=1.202
+ $X2=5.92 $Y2=1.202
r54 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.895
+ $Y=1.16 $X2=5.895 $Y2=1.16
r55 16 18 58.4827 $w=3.75e-07 $l=4.55e-07 $layer=POLY_cond $X=5.44 $Y=1.202
+ $X2=5.895 $Y2=1.202
r56 15 16 3.21333 $w=3.75e-07 $l=2.5e-08 $layer=POLY_cond $X=5.415 $Y=1.202
+ $X2=5.44 $Y2=1.202
r57 13 19 6.557 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=5.73 $Y=1.18
+ $X2=5.895 $Y2=1.18
r58 13 22 0.397394 $w=2.88e-07 $l=1e-08 $layer=LI1_cond $X=5.73 $Y=1.18 $X2=5.72
+ $Y2=1.18
r59 10 20 19.9308 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.92 $Y=1.41
+ $X2=5.92 $Y2=1.202
r60 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.92 $Y=1.41
+ $X2=5.92 $Y2=1.985
r61 7 18 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.895 $Y=0.995
+ $X2=5.895 $Y2=1.202
r62 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.895 $Y=0.995
+ $X2=5.895 $Y2=0.56
r63 4 16 19.9308 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.44 $Y=1.41
+ $X2=5.44 $Y2=1.202
r64 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.44 $Y=1.41 $X2=5.44
+ $Y2=1.985
r65 1 15 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.415 $Y=0.995
+ $X2=5.415 $Y2=1.202
r66 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.415 $Y=0.995
+ $X2=5.415 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 39 41 44
+ 45 46 48 53 58 67 71 77 80 83 86 90
r108 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r109 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r110 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r111 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r112 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r113 75 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r114 75 87 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=4.83 $Y2=2.72
r115 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r116 72 86 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=4.86 $Y=2.72
+ $X2=4.727 $Y2=2.72
r117 72 74 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=4.86 $Y=2.72
+ $X2=6.21 $Y2=2.72
r118 71 89 5.26454 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=6.425 $Y=2.72
+ $X2=6.662 $Y2=2.72
r119 71 74 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.425 $Y=2.72
+ $X2=6.21 $Y2=2.72
r120 70 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r121 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r122 67 86 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=4.595 $Y=2.72
+ $X2=4.727 $Y2=2.72
r123 67 69 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.595 $Y=2.72
+ $X2=4.37 $Y2=2.72
r124 66 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r125 66 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r126 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r127 63 83 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.78 $Y=2.72
+ $X2=2.59 $Y2=2.72
r128 63 65 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.78 $Y=2.72
+ $X2=3.45 $Y2=2.72
r129 62 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r130 62 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r131 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r132 59 80 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.82 $Y=2.72
+ $X2=1.63 $Y2=2.72
r133 59 61 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.82 $Y=2.72
+ $X2=2.07 $Y2=2.72
r134 58 83 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.4 $Y=2.72 $X2=2.59
+ $Y2=2.72
r135 58 61 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.4 $Y=2.72
+ $X2=2.07 $Y2=2.72
r136 57 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r137 57 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r138 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r139 54 77 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.86 $Y=2.72
+ $X2=0.67 $Y2=2.72
r140 54 56 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.86 $Y=2.72
+ $X2=1.15 $Y2=2.72
r141 53 80 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.44 $Y=2.72
+ $X2=1.63 $Y2=2.72
r142 53 56 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.44 $Y=2.72
+ $X2=1.15 $Y2=2.72
r143 48 77 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.48 $Y=2.72
+ $X2=0.67 $Y2=2.72
r144 48 50 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.48 $Y=2.72
+ $X2=0.23 $Y2=2.72
r145 46 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r146 46 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r147 44 65 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=2.72
+ $X2=3.45 $Y2=2.72
r148 44 45 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.535 $Y=2.72
+ $X2=3.725 $Y2=2.72
r149 43 69 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.915 $Y=2.72
+ $X2=4.37 $Y2=2.72
r150 43 45 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.915 $Y=2.72
+ $X2=3.725 $Y2=2.72
r151 39 89 2.93215 $w=3.8e-07 $l=1.05924e-07 $layer=LI1_cond $X=6.615 $Y=2.635
+ $X2=6.662 $Y2=2.72
r152 39 41 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=6.615 $Y=2.635
+ $X2=6.615 $Y2=2
r153 35 86 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=4.727 $Y=2.635
+ $X2=4.727 $Y2=2.72
r154 35 37 11.9593 $w=2.63e-07 $l=2.75e-07 $layer=LI1_cond $X=4.727 $Y=2.635
+ $X2=4.727 $Y2=2.36
r155 31 45 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=2.635
+ $X2=3.725 $Y2=2.72
r156 31 33 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=3.725 $Y=2.635
+ $X2=3.725 $Y2=2.36
r157 27 83 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=2.635
+ $X2=2.59 $Y2=2.72
r158 27 29 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.59 $Y=2.635
+ $X2=2.59 $Y2=2.32
r159 23 80 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=2.635
+ $X2=1.63 $Y2=2.72
r160 23 25 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=1.63 $Y=2.635
+ $X2=1.63 $Y2=1.955
r161 19 77 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=2.635
+ $X2=0.67 $Y2=2.72
r162 19 21 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=0.67 $Y=2.635
+ $X2=0.67 $Y2=1.955
r163 6 41 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=6.49
+ $Y=1.485 $X2=6.64 $Y2=2
r164 5 37 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=4.575
+ $Y=1.485 $X2=4.725 $Y2=2.36
r165 4 33 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=3.6
+ $Y=1.485 $X2=3.75 $Y2=2.36
r166 3 29 600 $w=1.7e-07 $l=9.04599e-07 $layer=licon1_PDIFF $count=1 $X=2.47
+ $Y=1.485 $X2=2.615 $Y2=2.32
r167 2 25 300 $w=1.7e-07 $l=5.37634e-07 $layer=licon1_PDIFF $count=2 $X=1.51
+ $Y=1.485 $X2=1.655 $Y2=1.955
r168 1 21 300 $w=1.7e-07 $l=5.50591e-07 $layer=licon1_PDIFF $count=2 $X=0.52
+ $Y=1.485 $X2=0.695 $Y2=1.955
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_4%X 1 2 3 4 13 15 16 19 21 25 27 31 35 38 39
+ 40 43 45
c68 13 0 1.11396e-19 $X=0.645 $Y=0.72
r69 43 45 1.85214 $w=2.78e-07 $l=4.5e-08 $layer=LI1_cond $X=0.225 $Y=0.805
+ $X2=0.225 $Y2=0.85
r70 40 43 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.225 $Y=0.72
+ $X2=0.225 $Y2=0.805
r71 40 45 0.823174 $w=2.78e-07 $l=2e-08 $layer=LI1_cond $X=0.225 $Y=0.87
+ $X2=0.225 $Y2=0.85
r72 37 40 23.2547 $w=2.78e-07 $l=5.65e-07 $layer=LI1_cond $X=0.225 $Y=1.435
+ $X2=0.225 $Y2=0.87
r73 33 35 8.46412 $w=1.88e-07 $l=1.45e-07 $layer=LI1_cond $X=2.135 $Y=1.7
+ $X2=2.135 $Y2=1.845
r74 29 31 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.67 $Y=0.615
+ $X2=1.67 $Y2=0.42
r75 28 39 3.70371 $w=2.65e-07 $l=9e-08 $layer=LI1_cond $X=1.26 $Y=1.567 $X2=1.17
+ $Y2=1.567
r76 27 33 7.06018 $w=2.65e-07 $l=1.74138e-07 $layer=LI1_cond $X=2.04 $Y=1.567
+ $X2=2.135 $Y2=1.7
r77 27 28 33.921 $w=2.63e-07 $l=7.8e-07 $layer=LI1_cond $X=2.04 $Y=1.567
+ $X2=1.26 $Y2=1.567
r78 23 39 2.76582 $w=1.8e-07 $l=1.33e-07 $layer=LI1_cond $X=1.17 $Y=1.7 $X2=1.17
+ $Y2=1.567
r79 23 25 8.93434 $w=1.78e-07 $l=1.45e-07 $layer=LI1_cond $X=1.17 $Y=1.7
+ $X2=1.17 $Y2=1.845
r80 22 38 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0.71
+ $X2=0.73 $Y2=0.71
r81 21 29 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.585 $Y=0.71
+ $X2=1.67 $Y2=0.615
r82 21 22 44.9474 $w=1.88e-07 $l=7.7e-07 $layer=LI1_cond $X=1.585 $Y=0.71
+ $X2=0.815 $Y2=0.71
r83 17 38 1.54918 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.73 $Y=0.615
+ $X2=0.73 $Y2=0.71
r84 17 19 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.73 $Y=0.615
+ $X2=0.73 $Y2=0.42
r85 16 37 6.82321 $w=2.65e-07 $l=1.95141e-07 $layer=LI1_cond $X=0.365 $Y=1.567
+ $X2=0.225 $Y2=1.435
r86 15 39 3.70371 $w=2.65e-07 $l=9e-08 $layer=LI1_cond $X=1.08 $Y=1.567 $X2=1.17
+ $Y2=1.567
r87 15 16 31.0942 $w=2.63e-07 $l=7.15e-07 $layer=LI1_cond $X=1.08 $Y=1.567
+ $X2=0.365 $Y2=1.567
r88 14 40 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.365 $Y=0.72
+ $X2=0.225 $Y2=0.72
r89 13 38 4.92476 $w=1.8e-07 $l=8.9861e-08 $layer=LI1_cond $X=0.645 $Y=0.72
+ $X2=0.73 $Y2=0.71
r90 13 14 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.645 $Y=0.72
+ $X2=0.365 $Y2=0.72
r91 4 35 300 $w=1.7e-07 $l=4.2638e-07 $layer=licon1_PDIFF $count=2 $X=1.99
+ $Y=1.485 $X2=2.135 $Y2=1.845
r92 3 25 300 $w=1.7e-07 $l=4.2638e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.485 $X2=1.175 $Y2=1.845
r93 2 31 182 $w=1.7e-07 $l=2.59856e-07 $layer=licon1_NDIFF $count=1 $X=1.49
+ $Y=0.235 $X2=1.67 $Y2=0.42
r94 1 19 182 $w=1.7e-07 $l=2.59856e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.73 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_4%VGND 1 2 3 4 5 16 18 22 26 30 33 34 36 37
+ 38 40 45 61 62 68
r100 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r101 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r102 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.67
+ $Y2=0
r103 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r104 56 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r105 55 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r106 53 56 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=0 $X2=4.83
+ $Y2=0
r107 53 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r108 52 55 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=4.83
+ $Y2=0
r109 52 53 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r110 50 52 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.53
+ $Y2=0
r111 49 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r112 49 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r113 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r114 46 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.2
+ $Y2=0
r115 46 48 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.61
+ $Y2=0
r116 45 75 10.5525 $w=4.13e-07 $l=3.8e-07 $layer=LI1_cond $X=2.132 $Y=0
+ $X2=2.132 $Y2=0.38
r117 45 50 6.00275 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=2.132 $Y=0 $X2=2.34
+ $Y2=0
r118 45 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r119 45 48 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.925 $Y=0
+ $X2=1.61 $Y2=0
r120 44 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r121 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r122 41 65 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r123 41 43 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.69 $Y2=0
r124 40 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.2
+ $Y2=0
r125 40 43 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r126 38 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r127 38 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r128 36 58 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.065 $Y=0
+ $X2=5.75 $Y2=0
r129 36 37 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.065 $Y=0 $X2=6.16
+ $Y2=0
r130 35 61 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.255 $Y=0
+ $X2=6.67 $Y2=0
r131 35 37 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.255 $Y=0 $X2=6.16
+ $Y2=0
r132 33 55 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.98 $Y=0 $X2=4.83
+ $Y2=0
r133 33 34 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=4.98 $Y=0 $X2=5.137
+ $Y2=0
r134 32 58 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=5.295 $Y=0
+ $X2=5.75 $Y2=0
r135 32 34 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=5.295 $Y=0
+ $X2=5.137 $Y2=0
r136 28 37 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.16 $Y=0.085
+ $X2=6.16 $Y2=0
r137 28 30 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=6.16 $Y=0.085
+ $X2=6.16 $Y2=0.36
r138 24 34 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.137 $Y=0.085
+ $X2=5.137 $Y2=0
r139 24 26 10.061 $w=3.13e-07 $l=2.75e-07 $layer=LI1_cond $X=5.137 $Y=0.085
+ $X2=5.137 $Y2=0.36
r140 20 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.085 $X2=1.2
+ $Y2=0
r141 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0.36
r142 16 65 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r143 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r144 5 30 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=5.97
+ $Y=0.235 $X2=6.16 $Y2=0.36
r145 4 26 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=4.95
+ $Y=0.235 $X2=5.13 $Y2=0.36
r146 3 75 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=1.96
+ $Y=0.235 $X2=2.14 $Y2=0.38
r147 2 22 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.235 $X2=1.2 $Y2=0.36
r148 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_4%A_524_47# 1 2 3 4 13 17 18 19 20 23 25 29
+ 33
c70 20 0 6.40318e-20 $X=4.805 $Y=0.78
r71 27 29 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=6.615 $Y=0.695
+ $X2=6.615 $Y2=0.38
r72 26 33 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.845 $Y=0.78
+ $X2=5.655 $Y2=0.78
r73 25 27 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=6.425 $Y=0.78
+ $X2=6.615 $Y2=0.695
r74 25 26 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=6.425 $Y=0.78
+ $X2=5.845 $Y2=0.78
r75 21 33 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.655 $Y=0.695
+ $X2=5.655 $Y2=0.78
r76 21 23 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.655 $Y=0.695
+ $X2=5.655 $Y2=0.36
r77 19 33 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.465 $Y=0.78
+ $X2=5.655 $Y2=0.78
r78 19 20 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=5.465 $Y=0.78
+ $X2=4.805 $Y2=0.78
r79 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.64 $Y=0.695
+ $X2=4.805 $Y2=0.78
r80 17 32 2.82476 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=4.64 $Y=0.465
+ $X2=4.64 $Y2=0.36
r81 17 18 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=4.64 $Y=0.465
+ $X2=4.64 $Y2=0.695
r82 13 32 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=0.36
+ $X2=4.64 $Y2=0.36
r83 13 15 91.368 $w=2.08e-07 $l=1.73e-06 $layer=LI1_cond $X=4.475 $Y=0.36
+ $X2=2.745 $Y2=0.36
r84 4 29 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=6.45
+ $Y=0.235 $X2=6.64 $Y2=0.38
r85 3 23 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=5.49
+ $Y=0.235 $X2=5.68 $Y2=0.36
r86 2 32 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=4.475
+ $Y=0.235 $X2=4.64 $Y2=0.42
r87 1 15 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.62
+ $Y=0.235 $X2=2.745 $Y2=0.38
.ends

