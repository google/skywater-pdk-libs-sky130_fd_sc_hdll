* File: sky130_fd_sc_hdll__a211o_2.pex.spice
* Created: Wed Sep  2 08:15:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A211O_2%A_79_21# 1 2 3 10 12 13 15 16 18 19 21 25
+ 27 28 29 30 33 35 39 43 45 49
r102 48 49 1.98626 $w=3.64e-07 $l=1.5e-08 $layer=POLY_cond $X=0.95 $Y=1.202
+ $X2=0.965 $Y2=1.202
r103 47 48 60.25 $w=3.64e-07 $l=4.55e-07 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.95 $Y2=1.202
r104 46 47 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r105 41 43 2.88111 $w=3.78e-07 $l=9.5e-08 $layer=LI1_cond $X=3.745 $Y=1.66
+ $X2=3.745 $Y2=1.755
r106 37 39 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=3.745 $Y=0.695
+ $X2=3.745 $Y2=0.4
r107 36 45 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.855 $Y=0.785
+ $X2=2.665 $Y2=0.785
r108 35 37 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=3.555 $Y=0.785
+ $X2=3.745 $Y2=0.695
r109 35 36 43.1313 $w=1.78e-07 $l=7e-07 $layer=LI1_cond $X=3.555 $Y=0.785
+ $X2=2.855 $Y2=0.785
r110 31 45 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=2.665 $Y=0.695
+ $X2=2.665 $Y2=0.785
r111 31 33 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.665 $Y=0.695
+ $X2=2.665 $Y2=0.36
r112 29 41 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=3.555 $Y=1.575
+ $X2=3.745 $Y2=1.66
r113 29 30 143.529 $w=1.68e-07 $l=2.2e-06 $layer=LI1_cond $X=3.555 $Y=1.575
+ $X2=1.355 $Y2=1.575
r114 27 45 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.475 $Y=0.785
+ $X2=2.665 $Y2=0.785
r115 27 28 69.0101 $w=1.78e-07 $l=1.12e-06 $layer=LI1_cond $X=2.475 $Y=0.785
+ $X2=1.355 $Y2=0.785
r116 26 49 29.1319 $w=3.64e-07 $l=2.2e-07 $layer=POLY_cond $X=1.185 $Y=1.202
+ $X2=0.965 $Y2=1.202
r117 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.185
+ $Y=1.16 $X2=1.185 $Y2=1.16
r118 23 30 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=1.227 $Y=1.49
+ $X2=1.355 $Y2=1.575
r119 23 25 14.914 $w=2.53e-07 $l=3.3e-07 $layer=LI1_cond $X=1.227 $Y=1.49
+ $X2=1.227 $Y2=1.16
r120 22 28 7.08339 $w=1.8e-07 $l=1.67045e-07 $layer=LI1_cond $X=1.227 $Y=0.875
+ $X2=1.355 $Y2=0.785
r121 22 25 12.8802 $w=2.53e-07 $l=2.85e-07 $layer=LI1_cond $X=1.227 $Y=0.875
+ $X2=1.227 $Y2=1.16
r122 19 49 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r123 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r124 16 48 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.95 $Y=0.995
+ $X2=0.95 $Y2=1.202
r125 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.95 $Y=0.995
+ $X2=0.95 $Y2=0.56
r126 13 47 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r127 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r128 10 46 23.572 $w=1.5e-07 $l=2.02e-07 $layer=POLY_cond $X=0.47 $Y=1 $X2=0.47
+ $Y2=1.202
r129 10 12 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.47 $Y=1 $X2=0.47
+ $Y2=0.56
r130 3 43 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=3.625
+ $Y=1.485 $X2=3.77 $Y2=1.755
r131 2 39 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=3.585
+ $Y=0.235 $X2=3.77 $Y2=0.4
r132 1 33 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=2.5
+ $Y=0.235 $X2=2.69 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_2%A2 1 3 4 6 7 12
r33 12 13 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=2.005 $Y=1.202
+ $X2=2.03 $Y2=1.202
r34 10 12 34.4286 $w=3.64e-07 $l=2.6e-07 $layer=POLY_cond $X=1.745 $Y=1.202
+ $X2=2.005 $Y2=1.202
r35 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.745
+ $Y=1.16 $X2=1.745 $Y2=1.16
r36 4 13 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.03 $Y=0.995
+ $X2=2.03 $Y2=1.202
r37 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.03 $Y=0.995 $X2=2.03
+ $Y2=0.56
r38 1 12 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.005 $Y=1.41
+ $X2=2.005 $Y2=1.202
r39 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.005 $Y=1.41
+ $X2=2.005 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_2%A1 1 3 4 6 7 14
r30 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.485
+ $Y=1.16 $X2=2.485 $Y2=1.16
r31 7 14 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.52 $Y=1.16
+ $X2=2.485 $Y2=1.16
r32 4 10 47.4309 $w=3.07e-07 $l=2.81957e-07 $layer=POLY_cond $X=2.585 $Y=1.41
+ $X2=2.517 $Y2=1.16
r33 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.585 $Y=1.41
+ $X2=2.585 $Y2=1.985
r34 1 10 38.5336 $w=3.07e-07 $l=2.05925e-07 $layer=POLY_cond $X=2.425 $Y=0.995
+ $X2=2.517 $Y2=1.16
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.425 $Y=0.995
+ $X2=2.425 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_2%B1 1 3 4 6 7 14
r27 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.03
+ $Y=1.16 $X2=3.03 $Y2=1.16
r28 7 14 1.50319 $w=2.28e-07 $l=3e-08 $layer=LI1_cond $X=3.06 $Y=1.16 $X2=3.03
+ $Y2=1.16
r29 4 10 47.6478 $w=3.03e-07 $l=2.80624e-07 $layer=POLY_cond $X=3.125 $Y=1.41
+ $X2=3.06 $Y2=1.16
r30 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.125 $Y=1.41
+ $X2=3.125 $Y2=1.985
r31 1 10 38.5416 $w=3.03e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.97 $Y=0.995
+ $X2=3.06 $Y2=1.16
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.97 $Y=0.995 $X2=2.97
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_2%C1 1 3 4 6 7
r22 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.16 $X2=3.57 $Y2=1.16
r23 4 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.535 $Y=1.41
+ $X2=3.57 $Y2=1.16
r24 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.535 $Y=1.41
+ $X2=3.535 $Y2=1.985
r25 1 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.57 $Y2=1.16
r26 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.51 $Y=0.995 $X2=3.51
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_2%VPWR 1 2 3 10 12 16 20 24 27 28 29 39 40
+ 46
r53 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r54 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r55 37 40 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r56 36 39 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r57 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r58 34 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r59 34 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r60 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r61 31 46 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=1.227 $Y2=2.72
r62 31 33 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=2.07 $Y2=2.72
r63 29 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r64 29 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r65 27 33 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=2.72
+ $X2=2.07 $Y2=2.72
r66 27 28 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=2.155 $Y=2.72
+ $X2=2.292 $Y2=2.72
r67 26 36 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.43 $Y=2.72 $X2=2.53
+ $Y2=2.72
r68 26 28 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=2.43 $Y=2.72
+ $X2=2.292 $Y2=2.72
r69 22 28 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.292 $Y=2.635
+ $X2=2.292 $Y2=2.72
r70 22 24 11.734 $w=2.73e-07 $l=2.8e-07 $layer=LI1_cond $X=2.292 $Y=2.635
+ $X2=2.292 $Y2=2.355
r71 18 46 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.227 $Y=2.635
+ $X2=1.227 $Y2=2.72
r72 18 20 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=1.227 $Y=2.635
+ $X2=1.227 $Y2=2
r73 17 43 4.46799 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.192 $Y2=2.72
r74 16 46 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.1 $Y=2.72
+ $X2=1.227 $Y2=2.72
r75 16 17 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.1 $Y=2.72
+ $X2=0.385 $Y2=2.72
r76 12 15 26.5648 $w=2.93e-07 $l=6.8e-07 $layer=LI1_cond $X=0.237 $Y=1.655
+ $X2=0.237 $Y2=2.335
r77 10 43 3.00953 $w=2.95e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.237 $Y=2.635
+ $X2=0.192 $Y2=2.72
r78 10 15 11.7198 $w=2.93e-07 $l=3e-07 $layer=LI1_cond $X=0.237 $Y=2.635
+ $X2=0.237 $Y2=2.335
r79 3 24 600 $w=1.7e-07 $l=9.6933e-07 $layer=licon1_PDIFF $count=1 $X=2.095
+ $Y=1.485 $X2=2.305 $Y2=2.355
r80 2 20 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r81 1 15 400 $w=1.7e-07 $l=9.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.335
r82 1 12 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.655
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_2%X 1 2 7 10
r15 10 13 60.378 $w=2.28e-07 $l=1.205e-06 $layer=LI1_cond $X=0.72 $Y=0.42
+ $X2=0.72 $Y2=1.625
r16 7 13 29.3121 $w=2.28e-07 $l=5.85e-07 $layer=LI1_cond $X=0.72 $Y=2.21
+ $X2=0.72 $Y2=1.625
r17 2 13 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.625
r18 1 10 91 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_2%A_319_297# 1 2 9 14 16
r26 10 14 5.43773 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.935 $Y=1.93
+ $X2=1.745 $Y2=1.93
r27 9 16 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.715 $Y=1.93
+ $X2=2.88 $Y2=1.93
r28 9 10 48.0606 $w=1.78e-07 $l=7.8e-07 $layer=LI1_cond $X=2.715 $Y=1.93
+ $X2=1.935 $Y2=1.93
r29 2 16 300 $w=1.7e-07 $l=6.08933e-07 $layer=licon1_PDIFF $count=2 $X=2.675
+ $Y=1.485 $X2=2.88 $Y2=2
r30 1 14 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=1.595
+ $Y=1.485 $X2=1.72 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_2%VGND 1 2 3 10 12 16 19 20 21 36 37 45 51
r53 49 51 9.59153 $w=5.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.61 $Y=0.18
+ $X2=1.77 $Y2=0.18
r54 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r55 47 49 1.24121 $w=5.28e-07 $l=5.5e-08 $layer=LI1_cond $X=1.555 $Y=0.18
+ $X2=1.61 $Y2=0.18
r56 44 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r57 43 47 9.13984 $w=5.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1.15 $Y=0.18
+ $X2=1.555 $Y2=0.18
r58 43 45 9.25302 $w=5.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.15 $Y=0.18
+ $X2=1.005 $Y2=0.18
r59 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r60 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r61 34 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r62 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r63 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r64 31 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r65 30 33 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r66 30 51 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.77
+ $Y2=0
r67 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r68 27 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r69 26 45 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.005
+ $Y2=0
r70 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r71 24 40 4.46799 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.192
+ $Y2=0
r72 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.69
+ $Y2=0
r73 21 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r74 21 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r75 19 33 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.11 $Y=0 $X2=2.99
+ $Y2=0
r76 19 20 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=3.11 $Y=0 $X2=3.247
+ $Y2=0
r77 18 36 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.91
+ $Y2=0
r78 18 20 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.247
+ $Y2=0
r79 14 20 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=3.247 $Y=0.085
+ $X2=3.247 $Y2=0
r80 14 16 11.5244 $w=2.73e-07 $l=2.75e-07 $layer=LI1_cond $X=3.247 $Y=0.085
+ $X2=3.247 $Y2=0.36
r81 10 40 3.00953 $w=2.95e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.237 $Y=0.085
+ $X2=0.192 $Y2=0
r82 10 12 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.237 $Y=0.085
+ $X2=0.237 $Y2=0.38
r83 3 16 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=3.045
+ $Y=0.235 $X2=3.27 $Y2=0.36
r84 2 47 91 $w=1.7e-07 $l=5.89194e-07 $layer=licon1_NDIFF $count=2 $X=1.025
+ $Y=0.235 $X2=1.555 $Y2=0.36
r85 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

