* File: sky130_fd_sc_hdll__sdfbbp_1.pex.spice
* Created: Thu Aug 27 19:26:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%CLK 4 5 7 8 10 13 19 20 24 26
c41 13 0 2.71124e-20 $X=0.52 $Y=0.805
r42 24 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.24 $Y=1.235
+ $X2=0.24 $Y2=1.4
r43 24 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.24 $Y=1.235
+ $X2=0.24 $Y2=1.07
r44 19 20 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.26 $Y=1.19
+ $X2=0.26 $Y2=1.53
r45 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.235 $X2=0.24 $Y2=1.235
r46 11 13 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=0.3 $Y=0.805
+ $X2=0.52 $Y2=0.805
r47 8 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.805
r48 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.445
r49 5 15 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=0.495 $Y=1.665
+ $X2=0.3 $Y2=1.665
r50 5 7 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.74
+ $X2=0.495 $Y2=2.135
r51 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.3 $Y=1.59 $X2=0.3
+ $Y2=1.665
r52 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.3 $Y=1.59 $X2=0.3
+ $Y2=1.4
r53 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.3 $Y=0.88 $X2=0.3
+ $Y2=0.805
r54 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.3 $Y=0.88 $X2=0.3
+ $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_27_47# 1 2 8 9 11 14 16 18 19 21 23 24
+ 26 27 28 31 35 39 40 41 44 46 50 51 54 55 56 57 58 67 73 81 84
c256 51 0 1.42522e-19 $X=5.07 $Y=0.87
c257 44 0 1.70452e-19 $X=0.77 $Y=1.795
c258 41 0 5.65522e-20 $X=0.655 $Y=1.88
c259 27 0 1.11465e-19 $X=9.81 $Y=1.32
c260 24 0 3.92095e-19 $X=9.28 $Y=1.99
r261 83 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.195
+ $Y=1.74 $X2=9.195 $Y2=1.74
r262 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.44
+ $Y=1.74 $X2=5.44 $Y2=1.74
r263 72 73 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.235
+ $X2=0.99 $Y2=1.235
r264 67 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.26 $Y=1.87
+ $X2=9.26 $Y2=1.87
r265 65 81 6.36876 $w=3.78e-07 $l=2.1e-07 $layer=LI1_cond $X=5.23 $Y=1.765
+ $X2=5.44 $Y2=1.765
r266 65 89 3.48766 $w=3.78e-07 $l=1.15e-07 $layer=LI1_cond $X=5.23 $Y=1.765
+ $X2=5.115 $Y2=1.765
r267 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.23 $Y=1.87
+ $X2=5.23 $Y2=1.87
r268 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.74 $Y=1.87
+ $X2=0.74 $Y2=1.87
r269 58 64 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=1.87
+ $X2=5.23 $Y2=1.87
r270 57 67 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.115 $Y=1.87
+ $X2=9.26 $Y2=1.87
r271 57 58 4.6287 $w=1.4e-07 $l=3.74e-06 $layer=MET1_cond $X=9.115 $Y=1.87
+ $X2=5.375 $Y2=1.87
r272 56 60 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.885 $Y=1.87
+ $X2=0.74 $Y2=1.87
r273 55 64 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.085 $Y=1.87
+ $X2=5.23 $Y2=1.87
r274 55 56 5.19801 $w=1.4e-07 $l=4.2e-06 $layer=MET1_cond $X=5.085 $Y=1.87
+ $X2=0.885 $Y2=1.87
r275 51 75 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=5.07 $Y=0.87
+ $X2=4.94 $Y2=0.87
r276 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.07
+ $Y=0.87 $X2=5.07 $Y2=0.87
r277 48 89 2.9592 $w=2.6e-07 $l=1.9e-07 $layer=LI1_cond $X=5.115 $Y=1.575
+ $X2=5.115 $Y2=1.765
r278 48 50 31.2489 $w=2.58e-07 $l=7.05e-07 $layer=LI1_cond $X=5.115 $Y=1.575
+ $X2=5.115 $Y2=0.87
r279 47 72 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.8 $Y=1.235
+ $X2=0.965 $Y2=1.235
r280 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.8
+ $Y=1.235 $X2=0.8 $Y2=1.235
r281 44 61 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=1.795
+ $X2=0.77 $Y2=1.88
r282 44 46 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.77 $Y=1.795
+ $X2=0.77 $Y2=1.235
r283 43 46 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.77 $Y=0.805
+ $X2=0.77 $Y2=1.235
r284 42 54 3.4683 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.257 $Y2=1.88
r285 41 61 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.655 $Y=1.88
+ $X2=0.77 $Y2=1.88
r286 41 42 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.655 $Y=1.88
+ $X2=0.345 $Y2=1.88
r287 39 43 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.655 $Y=0.72
+ $X2=0.77 $Y2=0.805
r288 39 40 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.655 $Y=0.72
+ $X2=0.345 $Y2=0.72
r289 33 40 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.257 $Y=0.635
+ $X2=0.345 $Y2=0.72
r290 33 35 7.92208 $w=1.73e-07 $l=1.25e-07 $layer=LI1_cond $X=0.257 $Y=0.635
+ $X2=0.257 $Y2=0.51
r291 29 31 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=9.885 $Y=1.245
+ $X2=9.885 $Y2=0.415
r292 27 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.81 $Y=1.32
+ $X2=9.885 $Y2=1.245
r293 27 28 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.81 $Y=1.32
+ $X2=9.38 $Y2=1.32
r294 24 83 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=9.28 $Y=1.99
+ $X2=9.22 $Y2=1.74
r295 24 26 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=9.28 $Y=1.99
+ $X2=9.28 $Y2=2.275
r296 23 83 31.9848 $w=2.95e-07 $l=1.92678e-07 $layer=POLY_cond $X=9.28 $Y=1.575
+ $X2=9.22 $Y2=1.74
r297 22 28 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=9.28 $Y=1.395
+ $X2=9.38 $Y2=1.32
r298 22 23 59.6839 $w=2e-07 $l=1.8e-07 $layer=POLY_cond $X=9.28 $Y=1.395
+ $X2=9.28 $Y2=1.575
r299 19 80 46.5577 $w=3.26e-07 $l=2.64575e-07 $layer=POLY_cond $X=5.435 $Y=1.99
+ $X2=5.465 $Y2=1.74
r300 19 21 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.435 $Y=1.99
+ $X2=5.435 $Y2=2.275
r301 16 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.94 $Y=0.705
+ $X2=4.94 $Y2=0.87
r302 16 18 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.94 $Y=0.705
+ $X2=4.94 $Y2=0.415
r303 12 73 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=1.235
r304 12 14 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=0.445
r305 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.965 $Y=1.74
+ $X2=0.965 $Y2=2.135
r306 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.64 $X2=0.965
+ $Y2=1.74
r307 7 72 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=0.965 $Y=1.37
+ $X2=0.965 $Y2=1.235
r308 7 8 89.5258 $w=2e-07 $l=2.7e-07 $layer=POLY_cond $X=0.965 $Y=1.37 $X2=0.965
+ $Y2=1.64
r309 2 54 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r310 1 35 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%SCD 1 3 6 8 9 15
r39 15 16 3.31956 $w=3.63e-07 $l=2.5e-08 $layer=POLY_cond $X=1.955 $Y=1.532
+ $X2=1.98 $Y2=1.532
r40 13 15 36.5152 $w=3.63e-07 $l=2.75e-07 $layer=POLY_cond $X=1.68 $Y=1.532
+ $X2=1.955 $Y2=1.532
r41 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.49 $X2=1.68 $Y2=1.49
r42 8 9 12.5721 $w=2.73e-07 $l=3e-07 $layer=LI1_cond $X=1.627 $Y=1.19 $X2=1.627
+ $Y2=1.49
r43 4 16 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.98 $Y=1.325
+ $X2=1.98 $Y2=1.532
r44 4 6 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=1.98 $Y=1.325 $X2=1.98
+ $Y2=0.445
r45 1 15 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.955 $Y=1.74
+ $X2=1.955 $Y2=1.532
r46 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.955 $Y=1.74
+ $X2=1.955 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_453_315# 1 2 7 9 10 11 12 14 17 21 23
+ 25 26 27 28 29 45
c109 45 0 1.39584e-19 $X=4.045 $Y=0.93
c110 29 0 4.64297e-20 $X=3.105 $Y=1.66
c111 25 0 1.15331e-19 $X=3.725 $Y=0.71
c112 10 0 1.35433e-19 $X=2.895 $Y=1.65
r113 38 45 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=3.935 $Y=0.93
+ $X2=4.045 $Y2=0.93
r114 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.935
+ $Y=0.93 $X2=3.935 $Y2=0.93
r115 32 34 8.46025 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=1.74
+ $X2=3.105 $Y2=1.905
r116 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.045
+ $Y=1.74 $X2=3.045 $Y2=1.74
r117 29 32 2.88111 $w=3.18e-07 $l=8e-08 $layer=LI1_cond $X=3.105 $Y=1.66
+ $X2=3.105 $Y2=1.74
r118 27 37 9.00568 $w=2.92e-07 $l=2.03912e-07 $layer=LI1_cond $X=3.81 $Y=1.095
+ $X2=3.897 $Y2=0.93
r119 27 28 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.81 $Y=1.095
+ $X2=3.81 $Y2=1.575
r120 25 37 9.19178 $w=2.92e-07 $l=2.93666e-07 $layer=LI1_cond $X=3.725 $Y=0.71
+ $X2=3.897 $Y2=0.93
r121 25 26 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.725 $Y=0.71
+ $X2=3.325 $Y2=0.71
r122 24 29 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.265 $Y=1.66
+ $X2=3.105 $Y2=1.66
r123 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.725 $Y=1.66
+ $X2=3.81 $Y2=1.575
r124 23 24 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.725 $Y=1.66
+ $X2=3.265 $Y2=1.66
r125 19 26 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.225 $Y=0.625
+ $X2=3.325 $Y2=0.71
r126 19 21 8.59545 $w=1.98e-07 $l=1.55e-07 $layer=LI1_cond $X=3.225 $Y=0.625
+ $X2=3.225 $Y2=0.47
r127 17 34 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.18 $Y=2.3
+ $X2=3.18 $Y2=1.905
r128 12 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.045 $Y=0.765
+ $X2=4.045 $Y2=0.93
r129 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.045 $Y=0.765
+ $X2=4.045 $Y2=0.445
r130 10 33 18.9432 $w=2.85e-07 $l=9e-08 $layer=POLY_cond $X=3.037 $Y=1.65
+ $X2=3.037 $Y2=1.74
r131 10 11 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.895 $Y=1.65
+ $X2=2.465 $Y2=1.65
r132 7 11 27.2212 $w=1.5e-07 $l=1.3784e-07 $layer=POLY_cond $X=2.365 $Y=1.74
+ $X2=2.465 $Y2=1.65
r133 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.365 $Y=1.74
+ $X2=2.365 $Y2=2.135
r134 2 17 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=3.055
+ $Y=2.065 $X2=3.18 $Y2=2.3
r135 1 21 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.235 $X2=3.24 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%SCE 1 3 4 7 8 10 11 13 14 16 18 19 20 23
+ 28 29 30 31 38
c109 28 0 2.04036e-19 $X=2.095 $Y=0.887
c110 23 0 8.9001e-20 $X=2.4 $Y=0.93
c111 20 0 1.79188e-19 $X=3.49 $Y=1.912
c112 14 0 2.88088e-19 $X=3.86 $Y=1.91
c113 4 0 4.64297e-20 $X=3.39 $Y=0.81
r114 30 31 12.2447 $w=3.18e-07 $l=3.4e-07 $layer=LI1_cond $X=2.095 $Y=1.19
+ $X2=2.095 $Y2=1.53
r115 27 30 6.30242 $w=3.18e-07 $l=1.75e-07 $layer=LI1_cond $X=2.095 $Y=1.015
+ $X2=2.095 $Y2=1.19
r116 27 28 4.4274 $w=3e-07 $l=1.28e-07 $layer=LI1_cond $X=2.095 $Y=1.015
+ $X2=2.095 $Y2=0.887
r117 26 29 10.2897 $w=2.78e-07 $l=2.5e-07 $layer=LI1_cond $X=2.115 $Y=0.76
+ $X2=2.115 $Y2=0.51
r118 26 28 4.4274 $w=3e-07 $l=1.36635e-07 $layer=LI1_cond $X=2.115 $Y=0.76
+ $X2=2.095 $Y2=0.887
r119 24 38 49.7885 $w=3.6e-07 $l=1.85e-07 $layer=POLY_cond $X=2.4 $Y=0.915
+ $X2=2.585 $Y2=0.915
r120 24 35 9.61737 $w=3.6e-07 $l=6e-08 $layer=POLY_cond $X=2.4 $Y=0.915 $X2=2.34
+ $Y2=0.915
r121 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.4
+ $Y=0.93 $X2=2.4 $Y2=0.93
r122 21 28 2.0066 $w=2.5e-07 $l=1.61493e-07 $layer=LI1_cond $X=2.255 $Y=0.89
+ $X2=2.095 $Y2=0.887
r123 21 23 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=2.255 $Y=0.89
+ $X2=2.4 $Y2=0.89
r124 16 18 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.96 $Y=1.99
+ $X2=3.96 $Y2=2.275
r125 15 20 8.71579 $w=1.5e-07 $l=1.00995e-07 $layer=POLY_cond $X=3.59 $Y=1.91
+ $X2=3.49 $Y2=1.912
r126 14 16 27.2212 $w=1.5e-07 $l=1.34164e-07 $layer=POLY_cond $X=3.86 $Y=1.91
+ $X2=3.96 $Y2=1.99
r127 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.86 $Y=1.91
+ $X2=3.59 $Y2=1.91
r128 11 19 17.9196 $w=1.75e-07 $l=8.66025e-08 $layer=POLY_cond $X=3.515 $Y=0.735
+ $X2=3.49 $Y2=0.81
r129 11 13 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.515 $Y=0.735
+ $X2=3.515 $Y2=0.445
r130 8 20 16.6942 $w=1.9e-07 $l=7.8e-08 $layer=POLY_cond $X=3.49 $Y=1.99
+ $X2=3.49 $Y2=1.912
r131 8 10 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.49 $Y=1.99
+ $X2=3.49 $Y2=2.275
r132 7 20 16.6942 $w=1.9e-07 $l=7.7e-08 $layer=POLY_cond $X=3.49 $Y=1.835
+ $X2=3.49 $Y2=1.912
r133 6 19 17.9196 $w=1.75e-07 $l=7.5e-08 $layer=POLY_cond $X=3.49 $Y=0.885
+ $X2=3.49 $Y2=0.81
r134 6 7 314.998 $w=2e-07 $l=9.5e-07 $layer=POLY_cond $X=3.49 $Y=0.885 $X2=3.49
+ $Y2=1.835
r135 4 19 7.5188 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=3.39 $Y=0.81 $X2=3.49
+ $Y2=0.81
r136 4 38 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=3.39 $Y=0.81
+ $X2=2.585 $Y2=0.81
r137 1 35 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.34 $Y=0.735
+ $X2=2.34 $Y2=0.915
r138 1 3 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.34 $Y=0.735
+ $X2=2.34 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%D 2 3 5 8 10 11 16 19
r47 18 19 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=4.43 $Y=1.49
+ $X2=4.455 $Y2=1.49
r48 15 18 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=4.24 $Y=1.49 $X2=4.43
+ $Y2=1.49
r49 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.24
+ $Y=1.49 $X2=4.24 $Y2=1.49
r50 10 11 24.4894 $w=3.18e-07 $l=6.8e-07 $layer=LI1_cond $X=4.315 $Y=1.53
+ $X2=4.315 $Y2=2.21
r51 10 16 1.44055 $w=3.18e-07 $l=4e-08 $layer=LI1_cond $X=4.315 $Y=1.53
+ $X2=4.315 $Y2=1.49
r52 6 19 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.455 $Y=1.355
+ $X2=4.455 $Y2=1.49
r53 6 8 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=4.455 $Y=1.355
+ $X2=4.455 $Y2=0.445
r54 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=4.43 $Y=1.99 $X2=4.43
+ $Y2=2.275
r55 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.43 $Y=1.89 $X2=4.43
+ $Y2=1.99
r56 1 18 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=4.43 $Y=1.625 $X2=4.43
+ $Y2=1.49
r57 1 2 87.868 $w=2e-07 $l=2.65e-07 $layer=POLY_cond $X=4.43 $Y=1.625 $X2=4.43
+ $Y2=1.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_211_363# 1 2 8 9 11 12 13 16 19 20 22
+ 23 25 28 29 31 33 36 37 39 40 41 48 52 56 57 66
c230 52 0 1.11465e-19 $X=9.26 $Y=1.19
c231 39 0 9.29232e-20 $X=5.777 $Y=1.12
c232 31 0 1.21258e-19 $X=9.762 $Y=1.305
c233 29 0 1.7288e-19 $X=9.37 $Y=0.87
c234 8 0 4.36039e-20 $X=4.965 $Y=1.89
r235 56 59 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=5.615 $Y=0.93
+ $X2=5.615 $Y2=1.095
r236 56 58 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=5.615 $Y=0.93
+ $X2=5.615 $Y2=0.765
r237 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.64
+ $Y=0.93 $X2=5.64 $Y2=0.93
r238 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.26 $Y=1.19
+ $X2=9.26 $Y2=1.19
r239 48 50 0.0661242 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=5.74 $Y=0.85
+ $X2=5.74 $Y2=0.965
r240 48 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.74 $Y=0.85
+ $X2=5.74 $Y2=0.85
r241 44 70 60.0532 $w=2.03e-07 $l=1.11e-06 $layer=LI1_cond $X=1.217 $Y=0.85
+ $X2=1.217 $Y2=1.96
r242 44 66 18.3947 $w=2.03e-07 $l=3.4e-07 $layer=LI1_cond $X=1.217 $Y=0.85
+ $X2=1.217 $Y2=0.51
r243 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.235 $Y=0.85
+ $X2=1.235 $Y2=0.85
r244 40 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.115 $Y=1.19
+ $X2=9.26 $Y2=1.19
r245 40 41 3.99752 $w=1.4e-07 $l=3.23e-06 $layer=MET1_cond $X=9.115 $Y=1.19
+ $X2=5.885 $Y2=1.19
r246 39 41 0.0739737 $w=1.4e-07 $l=1.38651e-07 $layer=MET1_cond $X=5.777 $Y=1.12
+ $X2=5.885 $Y2=1.19
r247 39 50 0.110669 $w=2.15e-07 $l=1.55e-07 $layer=MET1_cond $X=5.777 $Y=1.12
+ $X2=5.777 $Y2=0.965
r248 37 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.38 $Y=0.85
+ $X2=1.235 $Y2=0.85
r249 36 48 0.0513368 $w=1.4e-07 $l=1.45e-07 $layer=MET1_cond $X=5.595 $Y=0.85
+ $X2=5.74 $Y2=0.85
r250 36 37 5.21657 $w=1.4e-07 $l=4.215e-06 $layer=MET1_cond $X=5.595 $Y=0.85
+ $X2=1.38 $Y2=0.85
r251 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.755
+ $Y=1.74 $X2=9.755 $Y2=1.74
r252 31 53 30.9313 $w=1.78e-07 $l=5.02e-07 $layer=LI1_cond $X=9.762 $Y=1.215
+ $X2=9.26 $Y2=1.215
r253 31 33 19.6593 $w=2.53e-07 $l=4.35e-07 $layer=LI1_cond $X=9.762 $Y=1.305
+ $X2=9.762 $Y2=1.74
r254 29 60 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=9.37 $Y=0.87
+ $X2=9.245 $Y2=0.87
r255 28 53 8.64332 $w=3.38e-07 $l=2.55e-07 $layer=LI1_cond $X=9.34 $Y=0.87
+ $X2=9.34 $Y2=1.125
r256 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.37
+ $Y=0.87 $X2=9.37 $Y2=0.87
r257 23 34 46.5577 $w=3.26e-07 $l=2.64575e-07 $layer=POLY_cond $X=9.75 $Y=1.99
+ $X2=9.78 $Y2=1.74
r258 23 25 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=9.75 $Y=1.99
+ $X2=9.75 $Y2=2.275
r259 20 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.245 $Y=0.705
+ $X2=9.245 $Y2=0.87
r260 20 22 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.245 $Y=0.705
+ $X2=9.245 $Y2=0.415
r261 19 59 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=5.555 $Y=1.245
+ $X2=5.555 $Y2=1.095
r262 16 58 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=5.53 $Y=0.415
+ $X2=5.53 $Y2=0.765
r263 12 19 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=5.455 $Y=1.32
+ $X2=5.555 $Y2=1.245
r264 12 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=5.455 $Y=1.32
+ $X2=5.065 $Y2=1.32
r265 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=4.965 $Y=1.99
+ $X2=4.965 $Y2=2.275
r266 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.965 $Y=1.89 $X2=4.965
+ $Y2=1.99
r267 7 13 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=4.965 $Y=1.395
+ $X2=5.065 $Y2=1.32
r268 7 8 164.131 $w=2e-07 $l=4.95e-07 $layer=POLY_cond $X=4.965 $Y=1.395
+ $X2=4.965 $Y2=1.89
r269 2 70 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.815 $X2=1.2 $Y2=1.96
r270 1 66 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_1197_21# 1 2 9 11 13 15 16 18 19 21 22
+ 26 28 30 31 32 35 41 45 55
c147 35 0 5.34811e-20 $X=6.17 $Y=1.74
c148 16 0 1.14486e-19 $X=8.46 $Y=1.57
c149 15 0 1.67562e-19 $X=8.46 $Y=1.47
r150 49 55 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=8.66 $Y=1.15
+ $X2=8.77 $Y2=1.15
r151 49 52 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=8.66 $Y=1.15 $X2=8.46
+ $Y2=1.15
r152 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.66
+ $Y=1.15 $X2=8.66 $Y2=1.15
r153 45 48 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=8.66 $Y=0.98
+ $X2=8.66 $Y2=1.15
r154 43 44 12.6207 $w=2.9e-07 $l=3e-07 $layer=LI1_cond $X=7.465 $Y=0.68
+ $X2=7.465 $Y2=0.98
r155 35 38 6.53051 $w=2.98e-07 $l=1.7e-07 $layer=LI1_cond $X=6.235 $Y=1.74
+ $X2=6.235 $Y2=1.91
r156 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.17
+ $Y=1.74 $X2=6.17 $Y2=1.74
r157 33 44 3.86198 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.655 $Y=0.98
+ $X2=7.465 $Y2=0.98
r158 32 45 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=8.445 $Y=0.98
+ $X2=8.66 $Y2=0.98
r159 32 33 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=8.445 $Y=0.98
+ $X2=7.655 $Y2=0.98
r160 30 44 5.64745 $w=2.9e-07 $l=1.00995e-07 $layer=LI1_cond $X=7.5 $Y=1.065
+ $X2=7.465 $Y2=0.98
r161 30 31 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=7.5 $Y=1.065
+ $X2=7.5 $Y2=1.785
r162 29 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.105 $Y=1.91
+ $X2=7.02 $Y2=1.91
r163 28 31 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.415 $Y=1.91
+ $X2=7.5 $Y2=1.785
r164 28 29 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=7.415 $Y=1.91
+ $X2=7.105 $Y2=1.91
r165 24 41 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.02 $Y=2.035
+ $X2=7.02 $Y2=1.91
r166 24 26 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.02 $Y=2.035
+ $X2=7.02 $Y2=2.21
r167 23 38 1.80669 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=6.385 $Y=1.91
+ $X2=6.235 $Y2=1.91
r168 22 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.935 $Y=1.91
+ $X2=7.02 $Y2=1.91
r169 22 23 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=6.935 $Y=1.91
+ $X2=6.385 $Y2=1.91
r170 19 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.77 $Y=0.985
+ $X2=8.77 $Y2=1.15
r171 19 21 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.77 $Y=0.985
+ $X2=8.77 $Y2=0.555
r172 16 18 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=8.46 $Y=1.57
+ $X2=8.46 $Y2=2.065
r173 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=8.46 $Y=1.47 $X2=8.46
+ $Y2=1.57
r174 14 52 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=8.46 $Y=1.315
+ $X2=8.46 $Y2=1.15
r175 14 15 51.3945 $w=2e-07 $l=1.55e-07 $layer=POLY_cond $X=8.46 $Y=1.315
+ $X2=8.46 $Y2=1.47
r176 11 36 46.2237 $w=3.35e-07 $l=2.89396e-07 $layer=POLY_cond $X=6.085 $Y=1.99
+ $X2=6.17 $Y2=1.74
r177 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.085 $Y=1.99
+ $X2=6.085 $Y2=2.275
r178 7 36 38.6365 $w=3.35e-07 $l=2.13014e-07 $layer=POLY_cond $X=6.06 $Y=1.575
+ $X2=6.17 $Y2=1.74
r179 7 9 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=6.06 $Y=1.575
+ $X2=6.06 $Y2=0.445
r180 2 41 600 $w=1.7e-07 $l=3.49142e-07 $layer=licon1_PDIFF $count=1 $X=6.755
+ $Y=2.065 $X2=7.02 $Y2=1.87
r181 2 26 600 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_PDIFF $count=1 $X=6.755
+ $Y=2.065 $X2=7.02 $Y2=2.21
r182 1 43 182 $w=1.7e-07 $l=5.08035e-07 $layer=licon1_NDIFF $count=1 $X=7.355
+ $Y=0.235 $X2=7.49 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%SET_B 2 3 5 8 11 12 14 17 19 20 22 23 25
+ 28 37 40
c130 37 0 1.51196e-19 $X=11.005 $Y=0.98
c131 20 0 1.59387e-19 $X=6.815 $Y=0.85
c132 19 0 5.20549e-20 $X=10.655 $Y=0.85
c133 11 0 1.07745e-19 $X=10.98 $Y=1.89
c134 3 0 5.34811e-20 $X=6.665 $Y=1.99
r135 36 37 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=10.98 $Y=0.98
+ $X2=11.005 $Y2=0.98
r136 33 36 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=10.83 $Y=0.98
+ $X2=10.98 $Y2=0.98
r137 28 31 37.7137 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.59 $Y=0.98
+ $X2=6.59 $Y2=1.145
r138 28 30 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.59 $Y=0.98
+ $X2=6.59 $Y2=0.815
r139 28 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.55
+ $Y=0.98 $X2=6.55 $Y2=0.98
r140 25 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0.85
+ $X2=6.67 $Y2=0.85
r141 23 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.83
+ $Y=0.98 $X2=10.83 $Y2=0.98
r142 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0.85
+ $X2=10.8 $Y2=0.85
r143 20 25 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.815 $Y=0.85
+ $X2=6.67 $Y2=0.85
r144 19 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=0.85
+ $X2=10.8 $Y2=0.85
r145 19 20 4.75247 $w=1.4e-07 $l=3.84e-06 $layer=MET1_cond $X=10.655 $Y=0.85
+ $X2=6.815 $Y2=0.85
r146 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.005 $Y=0.815
+ $X2=11.005 $Y2=0.98
r147 15 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=11.005 $Y=0.815
+ $X2=11.005 $Y2=0.445
r148 12 14 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=10.98 $Y=1.99
+ $X2=10.98 $Y2=2.275
r149 11 12 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=10.98 $Y=1.89 $X2=10.98
+ $Y2=1.99
r150 10 36 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=10.98 $Y=1.145
+ $X2=10.98 $Y2=0.98
r151 10 11 247.025 $w=2e-07 $l=7.45e-07 $layer=POLY_cond $X=10.98 $Y=1.145
+ $X2=10.98 $Y2=1.89
r152 8 30 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.69 $Y=0.445
+ $X2=6.69 $Y2=0.815
r153 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.665 $Y=1.99
+ $X2=6.665 $Y2=2.275
r154 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=6.665 $Y=1.89 $X2=6.665
+ $Y2=1.99
r155 2 31 247.025 $w=2e-07 $l=7.45e-07 $layer=POLY_cond $X=6.665 $Y=1.89
+ $X2=6.665 $Y2=1.145
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_1003_47# 1 2 7 9 12 14 18 23 25 26 31
c107 31 0 4.36039e-20 $X=6.215 $Y=1.3
c108 7 0 5.20549e-20 $X=7.255 $Y=1.57
r109 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.11
+ $Y=1.32 $X2=7.11 $Y2=1.32
r110 30 31 6.2444 $w=2.08e-07 $l=1.1e-07 $layer=LI1_cond $X=6.105 $Y=1.3
+ $X2=6.215 $Y2=1.3
r111 28 30 14.5238 $w=2.08e-07 $l=2.75e-07 $layer=LI1_cond $X=5.83 $Y=1.3
+ $X2=6.105 $Y2=1.3
r112 26 33 8.9562 $w=3.2e-07 $l=1.65e-07 $layer=LI1_cond $X=6.945 $Y=1.32
+ $X2=7.11 $Y2=1.32
r113 26 31 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.945 $Y=1.32
+ $X2=6.215 $Y2=1.32
r114 25 30 0.430812 $w=2.2e-07 $l=1.05e-07 $layer=LI1_cond $X=6.105 $Y=1.195
+ $X2=6.105 $Y2=1.3
r115 24 25 38.2402 $w=2.18e-07 $l=7.3e-07 $layer=LI1_cond $X=6.105 $Y=0.465
+ $X2=6.105 $Y2=1.195
r116 22 28 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.83 $Y=1.405
+ $X2=5.83 $Y2=1.3
r117 22 23 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=5.83 $Y=1.405
+ $X2=5.83 $Y2=2.25
r118 18 24 6.83662 $w=2e-07 $l=1.51987e-07 $layer=LI1_cond $X=5.995 $Y=0.365
+ $X2=6.105 $Y2=0.465
r119 18 20 40.4818 $w=1.98e-07 $l=7.3e-07 $layer=LI1_cond $X=5.995 $Y=0.365
+ $X2=5.265 $Y2=0.365
r120 14 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.745 $Y=2.335
+ $X2=5.83 $Y2=2.25
r121 14 16 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=5.745 $Y=2.335
+ $X2=5.2 $Y2=2.335
r122 10 34 38.7084 $w=3.43e-07 $l=2.14942e-07 $layer=POLY_cond $X=7.28 $Y=1.155
+ $X2=7.165 $Y2=1.32
r123 10 12 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.28 $Y=1.155 $X2=7.28
+ $Y2=0.555
r124 7 34 45.964 $w=3.43e-07 $l=2.91548e-07 $layer=POLY_cond $X=7.255 $Y=1.57
+ $X2=7.165 $Y2=1.32
r125 7 9 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=7.255 $Y=1.57
+ $X2=7.255 $Y2=2.065
r126 2 16 600 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=1 $X=5.055
+ $Y=2.065 $X2=5.2 $Y2=2.335
r127 1 20 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=5.015
+ $Y=0.235 $X2=5.265 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_1525_21# 1 2 9 11 13 14 16 19 21 22 23
+ 25 29 32 40 41 44 47 51 54 57
c155 54 0 6.44034e-20 $X=12 $Y=1.362
c156 32 0 2.82048e-19 $X=7.97 $Y=1.32
c157 25 0 1.4422e-19 $X=12.73 $Y=1.66
r158 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.215
+ $Y=1.32 $X2=12.215 $Y2=1.32
r159 54 56 31.7883 $w=3.26e-07 $l=2.15e-07 $layer=POLY_cond $X=12 $Y=1.362
+ $X2=12.215 $Y2=1.362
r160 53 54 11.8282 $w=3.26e-07 $l=8e-08 $layer=POLY_cond $X=11.92 $Y=1.362
+ $X2=12 $Y2=1.362
r161 50 51 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=7.7 $Y=1.362
+ $X2=7.725 $Y2=1.362
r162 48 57 11.2564 $w=2.13e-07 $l=2.1e-07 $layer=LI1_cond $X=12.237 $Y=1.53
+ $X2=12.237 $Y2=1.32
r163 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.25 $Y=1.53
+ $X2=12.25 $Y2=1.53
r164 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.8 $Y=1.53 $X2=8.8
+ $Y2=1.53
r165 41 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.945 $Y=1.53
+ $X2=8.8 $Y2=1.53
r166 40 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.105 $Y=1.53
+ $X2=12.25 $Y2=1.53
r167 40 41 3.91088 $w=1.4e-07 $l=3.16e-06 $layer=MET1_cond $X=12.105 $Y=1.53
+ $X2=8.945 $Y2=1.53
r168 39 48 2.41209 $w=2.13e-07 $l=4.5e-08 $layer=LI1_cond $X=12.237 $Y=1.575
+ $X2=12.237 $Y2=1.53
r169 38 57 21.1728 $w=2.13e-07 $l=3.95e-07 $layer=LI1_cond $X=12.237 $Y=0.925
+ $X2=12.237 $Y2=1.32
r170 36 44 31.9323 $w=2.38e-07 $l=6.65e-07 $layer=LI1_cond $X=8.135 $Y=1.535
+ $X2=8.8 $Y2=1.535
r171 35 36 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=7.97 $Y=1.535
+ $X2=8.135 $Y2=1.535
r172 33 51 32.3534 $w=3.65e-07 $l=2.45e-07 $layer=POLY_cond $X=7.97 $Y=1.362
+ $X2=7.725 $Y2=1.362
r173 32 35 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=7.97 $Y=1.32
+ $X2=7.97 $Y2=1.535
r174 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.97
+ $Y=1.32 $X2=7.97 $Y2=1.32
r175 27 29 18.0227 $w=1.98e-07 $l=3.25e-07 $layer=LI1_cond $X=12.715 $Y=0.755
+ $X2=12.715 $Y2=0.43
r176 23 39 6.93832 $w=1.7e-07 $l=1.44375e-07 $layer=LI1_cond $X=12.345 $Y=1.66
+ $X2=12.237 $Y2=1.575
r177 23 25 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=12.345 $Y=1.66
+ $X2=12.73 $Y2=1.66
r178 22 38 6.93832 $w=1.7e-07 $l=1.44375e-07 $layer=LI1_cond $X=12.345 $Y=0.84
+ $X2=12.237 $Y2=0.925
r179 21 27 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=12.615 $Y=0.84
+ $X2=12.715 $Y2=0.755
r180 21 22 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=12.615 $Y=0.84
+ $X2=12.345 $Y2=0.84
r181 17 54 20.933 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=12 $Y=1.155 $X2=12
+ $Y2=1.362
r182 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=12 $Y=1.155 $X2=12
+ $Y2=0.555
r183 14 53 16.6478 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=11.92 $Y=1.57
+ $X2=11.92 $Y2=1.362
r184 14 16 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=11.92 $Y=1.57
+ $X2=11.92 $Y2=2.065
r185 11 51 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.725 $Y=1.57
+ $X2=7.725 $Y2=1.362
r186 11 13 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=7.725 $Y=1.57
+ $X2=7.725 $Y2=2.065
r187 7 50 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.7 $Y=1.155
+ $X2=7.7 $Y2=1.362
r188 7 9 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.7 $Y=1.155 $X2=7.7
+ $Y2=0.555
r189 2 25 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=12.605
+ $Y=1.505 $X2=12.73 $Y2=1.66
r190 1 29 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=12.605
+ $Y=0.235 $X2=12.73 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_2058_21# 1 2 9 11 13 14 16 17 19 20 23
+ 25 26 28 29 31 34 36 37 41 44 45 48 50 53 54 57 58 60 63 67
c183 37 0 2.52352e-20 $X=14.435 $Y=1.612
c184 14 0 1.4422e-19 $X=13.5 $Y=1.41
c185 9 0 8.84721e-20 $X=10.365 $Y=0.445
r186 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.44
+ $Y=1.16 $X2=13.44 $Y2=1.16
r187 64 67 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=13.345 $Y=1.16
+ $X2=13.44 $Y2=1.16
r188 56 64 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.345 $Y=1.325
+ $X2=13.345 $Y2=1.16
r189 56 57 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=13.345 $Y=1.325
+ $X2=13.345 $Y2=1.915
r190 55 63 5.53942 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=11.915 $Y=2
+ $X2=11.822 $Y2=2
r191 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.26 $Y=2
+ $X2=13.345 $Y2=1.915
r192 54 55 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=13.26 $Y=2
+ $X2=11.915 $Y2=2
r193 53 63 1.03991 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=11.822 $Y=1.915
+ $X2=11.822 $Y2=2
r194 52 60 0.22998 $w=1.85e-07 $l=1.15521e-07 $layer=LI1_cond $X=11.822 $Y=0.815
+ $X2=11.75 $Y2=0.73
r195 52 53 65.9459 $w=1.83e-07 $l=1.1e-06 $layer=LI1_cond $X=11.822 $Y=0.815
+ $X2=11.822 $Y2=1.915
r196 51 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.36 $Y=2
+ $X2=11.275 $Y2=2
r197 50 63 5.53942 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=11.73 $Y=2
+ $X2=11.822 $Y2=2
r198 50 51 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=11.73 $Y=2 $X2=11.36
+ $Y2=2
r199 46 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.275 $Y=2.085
+ $X2=11.275 $Y2=2
r200 46 48 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=11.275 $Y=2.085
+ $X2=11.275 $Y2=2.21
r201 44 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.19 $Y=2
+ $X2=11.275 $Y2=2
r202 44 45 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=11.19 $Y=2 $X2=10.7
+ $Y2=2
r203 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.485
+ $Y=1.74 $X2=10.485 $Y2=1.74
r204 39 45 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=10.55 $Y=1.915
+ $X2=10.7 $Y2=2
r205 39 41 6.72258 $w=2.98e-07 $l=1.75e-07 $layer=LI1_cond $X=10.55 $Y=1.915
+ $X2=10.55 $Y2=1.74
r206 32 34 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=14.435 $Y=0.805
+ $X2=14.61 $Y2=0.805
r207 29 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.61 $Y=0.73
+ $X2=14.61 $Y2=0.805
r208 29 31 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=14.61 $Y=0.73
+ $X2=14.61 $Y2=0.445
r209 26 37 47.2549 $w=1.53e-07 $l=1.5e-07 $layer=POLY_cond $X=14.585 $Y=1.612
+ $X2=14.435 $Y2=1.612
r210 26 28 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=14.585 $Y=1.69
+ $X2=14.585 $Y2=2.085
r211 25 37 3.30671 $w=1.5e-07 $l=7.7e-08 $layer=POLY_cond $X=14.435 $Y=1.535
+ $X2=14.435 $Y2=1.612
r212 24 36 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=14.435 $Y=1.295
+ $X2=14.435 $Y2=1.16
r213 24 25 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=14.435 $Y=1.295
+ $X2=14.435 $Y2=1.535
r214 23 36 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=14.435 $Y=1.025
+ $X2=14.435 $Y2=1.16
r215 22 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.435 $Y=0.88
+ $X2=14.435 $Y2=0.805
r216 22 23 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=14.435 $Y=0.88
+ $X2=14.435 $Y2=1.025
r217 21 68 3.27186 $w=2.7e-07 $l=1.48e-07 $layer=POLY_cond $X=13.6 $Y=1.16
+ $X2=13.452 $Y2=1.16
r218 20 36 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=14.36 $Y=1.16
+ $X2=14.435 $Y2=1.16
r219 20 21 168.852 $w=2.7e-07 $l=7.6e-07 $layer=POLY_cond $X=14.36 $Y=1.16
+ $X2=13.6 $Y2=1.16
r220 17 68 38.8084 $w=2.75e-07 $l=1.98167e-07 $layer=POLY_cond $X=13.525
+ $Y=0.995 $X2=13.452 $Y2=1.16
r221 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.525 $Y=0.995
+ $X2=13.525 $Y2=0.56
r222 14 68 49.5676 $w=2.75e-07 $l=2.72947e-07 $layer=POLY_cond $X=13.5 $Y=1.41
+ $X2=13.452 $Y2=1.16
r223 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=13.5 $Y=1.41
+ $X2=13.5 $Y2=1.985
r224 11 42 45.964 $w=3.43e-07 $l=2.91548e-07 $layer=POLY_cond $X=10.39 $Y=1.99
+ $X2=10.48 $Y2=1.74
r225 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=10.39 $Y=1.99
+ $X2=10.39 $Y2=2.275
r226 7 42 38.7084 $w=3.43e-07 $l=2.14942e-07 $layer=POLY_cond $X=10.365 $Y=1.575
+ $X2=10.48 $Y2=1.74
r227 7 9 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=10.365 $Y=1.575
+ $X2=10.365 $Y2=0.445
r228 2 48 600 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=11.07
+ $Y=2.065 $X2=11.275 $Y2=2.21
r229 1 60 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=11.61
+ $Y=0.235 $X2=11.75 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_1864_47# 1 2 7 9 12 14 18 23 25 26 28
+ 30
c95 30 0 1.72149e-19 $X=11.425 $Y=1.24
c96 25 0 1.86429e-19 $X=10.145 $Y=2.25
r97 30 33 4.1907 $w=2.18e-07 $l=8e-08 $layer=LI1_cond $X=11.4 $Y=1.24 $X2=11.4
+ $Y2=1.32
r98 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.425
+ $Y=1.24 $X2=11.425 $Y2=1.24
r99 27 28 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.23 $Y=1.32
+ $X2=10.145 $Y2=1.32
r100 26 33 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=11.29 $Y=1.32
+ $X2=11.4 $Y2=1.32
r101 26 27 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=11.29 $Y=1.32
+ $X2=10.23 $Y2=1.32
r102 24 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.145 $Y=1.405
+ $X2=10.145 $Y2=1.32
r103 24 25 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=10.145 $Y=1.405
+ $X2=10.145 $Y2=2.25
r104 23 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.145 $Y=1.235
+ $X2=10.145 $Y2=1.32
r105 22 23 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=10.145 $Y=0.465
+ $X2=10.145 $Y2=1.235
r106 18 22 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=10.06 $Y=0.365
+ $X2=10.145 $Y2=0.465
r107 18 20 26.6182 $w=1.98e-07 $l=4.8e-07 $layer=LI1_cond $X=10.06 $Y=0.365
+ $X2=9.58 $Y2=0.365
r108 14 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.06 $Y=2.335
+ $X2=10.145 $Y2=2.25
r109 14 16 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=10.06 $Y=2.335
+ $X2=9.515 $Y2=2.335
r110 10 31 38.7299 $w=2.8e-07 $l=2.03101e-07 $layer=POLY_cond $X=11.535 $Y=1.075
+ $X2=11.45 $Y2=1.24
r111 10 12 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=11.535 $Y=1.075
+ $X2=11.535 $Y2=0.555
r112 7 31 62.9382 $w=2.8e-07 $l=3.58748e-07 $layer=POLY_cond $X=11.51 $Y=1.57
+ $X2=11.45 $Y2=1.24
r113 7 9 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=11.51 $Y=1.57
+ $X2=11.51 $Y2=2.065
r114 2 16 600 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=1 $X=9.37
+ $Y=2.065 $X2=9.515 $Y2=2.335
r115 1 20 182 $w=1.7e-07 $l=3.245e-07 $layer=licon1_NDIFF $count=1 $X=9.32
+ $Y=0.235 $X2=9.58 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%RESET_B 1 3 6 8 12
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.75
+ $Y=1.18 $X2=12.75 $Y2=1.18
r33 8 12 5.01062 $w=2.28e-07 $l=1e-07 $layer=LI1_cond $X=12.65 $Y=1.21 $X2=12.75
+ $Y2=1.21
r34 4 11 39.5463 $w=3.98e-07 $l=2.2798e-07 $layer=POLY_cond $X=12.99 $Y=1.015
+ $X2=12.84 $Y2=1.18
r35 4 6 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=12.99 $Y=1.015
+ $X2=12.99 $Y2=0.445
r36 1 11 44.909 $w=3.98e-07 $l=3.06186e-07 $layer=POLY_cond $X=12.965 $Y=1.43
+ $X2=12.84 $Y2=1.18
r37 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=12.965 $Y=1.43
+ $X2=12.965 $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_2845_47# 1 2 7 9 10 12 13 15 19 25 28
+ 29
c55 29 0 1.98844e-19 $X=14.417 $Y=1.16
r56 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.005
+ $Y=1.16 $X2=15.005 $Y2=1.16
r57 23 29 0.30096 $w=3.3e-07 $l=1.03e-07 $layer=LI1_cond $X=14.52 $Y=1.16
+ $X2=14.417 $Y2=1.16
r58 23 25 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=14.52 $Y=1.16
+ $X2=15.005 $Y2=1.16
r59 21 29 7.52254 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=14.417 $Y=1.325
+ $X2=14.417 $Y2=1.16
r60 21 28 21.6408 $w=2.03e-07 $l=4e-07 $layer=LI1_cond $X=14.417 $Y=1.325
+ $X2=14.417 $Y2=1.725
r61 17 29 7.52254 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=14.417 $Y=0.995
+ $X2=14.417 $Y2=1.16
r62 17 19 26.2395 $w=2.03e-07 $l=4.85e-07 $layer=LI1_cond $X=14.417 $Y=0.995
+ $X2=14.417 $Y2=0.51
r63 13 28 6.21614 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=14.392 $Y=1.852
+ $X2=14.392 $Y2=1.725
r64 13 15 2.62124 $w=2.53e-07 $l=5.8e-08 $layer=LI1_cond $X=14.392 $Y=1.852
+ $X2=14.392 $Y2=1.91
r65 10 26 38.532 $w=3.11e-07 $l=2.07123e-07 $layer=POLY_cond $X=15.135 $Y=0.995
+ $X2=15.04 $Y2=1.16
r66 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=15.135 $Y=0.995
+ $X2=15.135 $Y2=0.56
r67 7 26 47.2262 $w=3.11e-07 $l=2.82843e-07 $layer=POLY_cond $X=15.11 $Y=1.41
+ $X2=15.04 $Y2=1.16
r68 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.11 $Y=1.41
+ $X2=15.11 $Y2=1.985
r69 2 15 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=14.225
+ $Y=1.765 $X2=14.35 $Y2=1.91
r70 1 19 182 $w=1.7e-07 $l=3.51781e-07 $layer=licon1_NDIFF $count=1 $X=14.225
+ $Y=0.235 $X2=14.4 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%VPWR 1 2 3 4 5 6 7 8 9 30 32 36 40 44 48
+ 52 55 56 58 61 62 64 66 79 83 91 104 108 117 118 121 124 127 130 133 141 146
c212 118 0 4.74427e-19 $X=15.41 $Y=2.72
c213 79 0 1.633e-19 $X=6.205 $Y=2.72
c214 1 0 5.65522e-20 $X=0.585 $Y=1.815
r215 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.95 $Y=2.72
+ $X2=14.95 $Y2=2.72
r216 143 144 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r217 140 143 0.761141 $w=5.48e-07 $l=3.5e-08 $layer=LI1_cond $X=12.155 $Y=2.53
+ $X2=12.19 $Y2=2.53
r218 140 141 10.9193 $w=5.48e-07 $l=2.15e-07 $layer=LI1_cond $X=12.155 $Y=2.53
+ $X2=11.94 $Y2=2.53
r219 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r220 133 136 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=10.71 $Y=2.34
+ $X2=10.71 $Y2=2.72
r221 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r222 127 128 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r223 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r224 122 125 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r225 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r226 118 147 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.41 $Y=2.72
+ $X2=14.95 $Y2=2.72
r227 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.41 $Y=2.72
+ $X2=15.41 $Y2=2.72
r228 115 146 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=15.04 $Y=2.72
+ $X2=14.892 $Y2=2.72
r229 115 117 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=15.04 $Y=2.72
+ $X2=15.41 $Y2=2.72
r230 114 147 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=2.72
+ $X2=14.95 $Y2=2.72
r231 113 114 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.49 $Y=2.72
+ $X2=14.49 $Y2=2.72
r232 111 114 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.57 $Y=2.72
+ $X2=14.49 $Y2=2.72
r233 110 113 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=13.57 $Y=2.72
+ $X2=14.49 $Y2=2.72
r234 110 111 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.57 $Y=2.72
+ $X2=13.57 $Y2=2.72
r235 108 146 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=14.745 $Y=2.72
+ $X2=14.892 $Y2=2.72
r236 108 113 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=14.745 $Y=2.72
+ $X2=14.49 $Y2=2.72
r237 107 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=2.72
+ $X2=13.57 $Y2=2.72
r238 107 144 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.11 $Y=2.72
+ $X2=12.19 $Y2=2.72
r239 106 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r240 104 143 0.543672 $w=5.48e-07 $l=2.5e-08 $layer=LI1_cond $X=12.215 $Y=2.53
+ $X2=12.19 $Y2=2.53
r241 104 106 19.4635 $w=5.48e-07 $l=8.95e-07 $layer=LI1_cond $X=12.215 $Y=2.53
+ $X2=13.11 $Y2=2.53
r242 103 144 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=12.19 $Y2=2.72
r243 103 137 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=10.81 $Y2=2.72
r244 102 141 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=11.73 $Y=2.72
+ $X2=11.94 $Y2=2.72
r245 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r246 100 136 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.9 $Y=2.72
+ $X2=10.71 $Y2=2.72
r247 100 102 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=10.9 $Y=2.72
+ $X2=11.73 $Y2=2.72
r248 98 137 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=10.81 $Y2=2.72
r249 97 98 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r250 95 98 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=10.35 $Y2=2.72
r251 95 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.05 $Y2=2.72
r252 94 97 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=8.51 $Y=2.72
+ $X2=10.35 $Y2=2.72
r253 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r254 92 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.155 $Y=2.72
+ $X2=7.99 $Y2=2.72
r255 92 94 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.155 $Y=2.72
+ $X2=8.51 $Y2=2.72
r256 91 136 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.52 $Y=2.72
+ $X2=10.71 $Y2=2.72
r257 91 97 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=10.52 $Y=2.72
+ $X2=10.35 $Y2=2.72
r258 90 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r259 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r260 87 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r261 87 128 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r262 86 89 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r263 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r264 84 127 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.585 $Y=2.72
+ $X2=6.395 $Y2=2.72
r265 84 86 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.585 $Y=2.72
+ $X2=6.67 $Y2=2.72
r266 83 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.825 $Y=2.72
+ $X2=7.99 $Y2=2.72
r267 83 89 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=7.825 $Y=2.72
+ $X2=7.59 $Y2=2.72
r268 82 128 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=6.21 $Y2=2.72
r269 81 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r270 79 127 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.205 $Y=2.72
+ $X2=6.395 $Y2=2.72
r271 79 81 149.727 $w=1.68e-07 $l=2.295e-06 $layer=LI1_cond $X=6.205 $Y=2.72
+ $X2=3.91 $Y2=2.72
r272 78 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r273 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r274 75 78 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r275 75 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r276 74 77 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r277 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r278 72 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=2.72
+ $X2=1.72 $Y2=2.72
r279 72 74 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.885 $Y=2.72
+ $X2=2.07 $Y2=2.72
r280 66 121 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r281 64 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r282 62 66 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.515 $Y2=2.72
r283 62 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r284 61 110 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=13.43 $Y=2.72
+ $X2=13.57 $Y2=2.72
r285 60 61 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=13.265 $Y=2.53
+ $X2=13.43 $Y2=2.53
r286 58 106 0.97861 $w=5.48e-07 $l=4.5e-08 $layer=LI1_cond $X=13.155 $Y=2.53
+ $X2=13.11 $Y2=2.53
r287 58 60 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=13.155 $Y=2.53
+ $X2=13.265 $Y2=2.53
r288 55 77 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.51 $Y=2.72 $X2=3.45
+ $Y2=2.72
r289 55 56 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.51 $Y=2.72 $X2=3.7
+ $Y2=2.72
r290 54 81 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.89 $Y=2.72 $X2=3.91
+ $Y2=2.72
r291 54 56 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.89 $Y=2.72 $X2=3.7
+ $Y2=2.72
r292 50 146 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=14.892 $Y=2.635
+ $X2=14.892 $Y2=2.72
r293 50 52 27.1508 $w=2.93e-07 $l=6.95e-07 $layer=LI1_cond $X=14.892 $Y=2.635
+ $X2=14.892 $Y2=1.94
r294 46 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.99 $Y=2.635
+ $X2=7.99 $Y2=2.72
r295 46 48 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=7.99 $Y=2.635
+ $X2=7.99 $Y2=2
r296 42 127 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.395 $Y=2.635
+ $X2=6.395 $Y2=2.72
r297 42 44 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=6.395 $Y=2.635
+ $X2=6.395 $Y2=2.29
r298 38 56 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=2.635 $X2=3.7
+ $Y2=2.72
r299 38 40 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.7 $Y=2.635
+ $X2=3.7 $Y2=2.3
r300 34 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=2.635
+ $X2=1.72 $Y2=2.72
r301 34 36 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=1.72 $Y=2.635
+ $X2=1.72 $Y2=1.97
r302 33 121 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r303 32 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=2.72
+ $X2=1.72 $Y2=2.72
r304 32 33 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.555 $Y=2.72
+ $X2=0.895 $Y2=2.72
r305 28 121 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r306 28 30 12.5859 $w=3.78e-07 $l=4.15e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.22
r307 9 52 300 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=2 $X=14.675
+ $Y=1.765 $X2=14.875 $Y2=1.94
r308 8 60 600 $w=1.7e-07 $l=9.34117e-07 $layer=licon1_PDIFF $count=1 $X=13.055
+ $Y=1.505 $X2=13.265 $Y2=2.34
r309 7 140 600 $w=1.7e-07 $l=7.64068e-07 $layer=licon1_PDIFF $count=1 $X=12.01
+ $Y=1.645 $X2=12.155 $Y2=2.34
r310 6 133 600 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_PDIFF $count=1 $X=10.48
+ $Y=2.065 $X2=10.685 $Y2=2.34
r311 5 48 300 $w=1.7e-07 $l=4.33763e-07 $layer=licon1_PDIFF $count=2 $X=7.815
+ $Y=1.645 $X2=7.99 $Y2=2
r312 4 44 600 $w=1.7e-07 $l=3.07409e-07 $layer=licon1_PDIFF $count=1 $X=6.175
+ $Y=2.065 $X2=6.37 $Y2=2.29
r313 3 40 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=2.065 $X2=3.725 $Y2=2.3
r314 2 36 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=1.595
+ $Y=1.815 $X2=1.72 $Y2=1.97
r315 1 30 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.815 $X2=0.73 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_483_47# 1 2 3 4 16 18 19 24 26 29 30 33
+ 36 42
c119 36 0 4.95985e-20 $X=4.73 $Y=1.19
c120 30 0 1.15331e-19 $X=3.335 $Y=1.19
c121 26 0 4.64318e-20 $X=2.955 $Y=1.22
c122 16 0 1.60218e-19 $X=2.87 $Y=1.075
r123 37 46 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=4.73 $Y=1.19
+ $X2=4.73 $Y2=2.3
r124 37 42 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.73 $Y=1.19
+ $X2=4.73 $Y2=0.47
r125 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.73 $Y=1.19
+ $X2=4.73 $Y2=1.19
r126 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.19 $Y=1.19
+ $X2=3.19 $Y2=1.19
r127 30 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.335 $Y=1.19
+ $X2=3.19 $Y2=1.19
r128 29 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.585 $Y=1.19
+ $X2=4.73 $Y2=1.19
r129 29 30 1.54703 $w=1.4e-07 $l=1.25e-06 $layer=MET1_cond $X=4.585 $Y=1.19
+ $X2=3.335 $Y2=1.19
r130 27 28 11.4982 $w=2.26e-07 $l=2.13e-07 $layer=LI1_cond $X=2.657 $Y=1.22
+ $X2=2.87 $Y2=1.22
r131 26 33 9.33876 $w=2.88e-07 $l=2.35e-07 $layer=LI1_cond $X=2.955 $Y=1.22
+ $X2=3.19 $Y2=1.22
r132 26 28 4.20283 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.955 $Y=1.22
+ $X2=2.87 $Y2=1.22
r133 22 24 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=2.635 $Y=0.43
+ $X2=2.87 $Y2=0.43
r134 18 19 4.73279 $w=3.78e-07 $l=8.5e-08 $layer=LI1_cond $X=2.575 $Y=1.96
+ $X2=2.575 $Y2=1.875
r135 16 28 2.4068 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.87 $Y=1.075
+ $X2=2.87 $Y2=1.22
r136 15 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.87 $Y=0.595
+ $X2=2.87 $Y2=0.43
r137 15 16 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.87 $Y=0.595
+ $X2=2.87 $Y2=1.075
r138 13 27 1.0459 $w=2.15e-07 $l=1.45e-07 $layer=LI1_cond $X=2.657 $Y=1.365
+ $X2=2.657 $Y2=1.22
r139 13 19 27.337 $w=2.13e-07 $l=5.1e-07 $layer=LI1_cond $X=2.657 $Y=1.365
+ $X2=2.657 $Y2=1.875
r140 4 46 600 $w=1.7e-07 $l=3.23381e-07 $layer=licon1_PDIFF $count=1 $X=4.52
+ $Y=2.065 $X2=4.73 $Y2=2.3
r141 3 18 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=2.455
+ $Y=1.815 $X2=2.6 $Y2=1.96
r142 2 42 182 $w=1.7e-07 $l=3.19726e-07 $layer=licon1_NDIFF $count=1 $X=4.53
+ $Y=0.235 $X2=4.73 $Y2=0.47
r143 1 22 182 $w=1.7e-07 $l=3.02159e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.235 $X2=2.635 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%Q_N 1 2 11 12 13 14
c32 11 0 2.52352e-20 $X=13.83 $Y=1.815
r33 27 28 5.57099 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=13.915 $Y=0.55
+ $X2=13.915 $Y2=0.715
r34 13 14 13.2824 $w=2.93e-07 $l=3.4e-07 $layer=LI1_cond $X=13.967 $Y=0.85
+ $X2=13.967 $Y2=1.19
r35 13 28 5.27389 $w=2.93e-07 $l=1.35e-07 $layer=LI1_cond $X=13.967 $Y=0.85
+ $X2=13.967 $Y2=0.715
r36 12 27 1.15244 $w=3.98e-07 $l=4e-08 $layer=LI1_cond $X=13.915 $Y=0.51
+ $X2=13.915 $Y2=0.55
r37 9 14 7.14905 $w=2.93e-07 $l=1.83e-07 $layer=LI1_cond $X=13.967 $Y=1.373
+ $X2=13.967 $Y2=1.19
r38 9 11 16.6768 $w=3.26e-07 $l=4.67277e-07 $layer=LI1_cond $X=13.967 $Y=1.373
+ $X2=13.915 $Y2=1.815
r39 2 11 300 $w=1.7e-07 $l=4.33705e-07 $layer=licon1_PDIFF $count=2 $X=13.59
+ $Y=1.485 $X2=13.83 $Y2=1.815
r40 1 27 182 $w=1.7e-07 $l=4.14337e-07 $layer=licon1_NDIFF $count=1 $X=13.6
+ $Y=0.235 $X2=13.83 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%Q 1 2 10 11 12 13 14 15
r17 14 15 15.7703 $w=2.83e-07 $l=3.9e-07 $layer=LI1_cond $X=15.402 $Y=1.82
+ $X2=15.402 $Y2=2.21
r18 11 14 2.95187 $w=2.83e-07 $l=7.3e-08 $layer=LI1_cond $X=15.402 $Y=1.747
+ $X2=15.402 $Y2=1.82
r19 11 12 6.13081 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=15.402 $Y=1.747
+ $X2=15.402 $Y2=1.605
r20 10 12 38.2513 $w=2.33e-07 $l=7.8e-07 $layer=LI1_cond $X=15.427 $Y=0.825
+ $X2=15.427 $Y2=1.605
r21 9 13 6.99553 $w=2.83e-07 $l=1.73e-07 $layer=LI1_cond $X=15.402 $Y=0.683
+ $X2=15.402 $Y2=0.51
r22 9 10 6.13081 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=15.402 $Y=0.683
+ $X2=15.402 $Y2=0.825
r23 2 14 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=15.2
+ $Y=1.485 $X2=15.345 $Y2=1.82
r24 1 13 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=15.21
+ $Y=0.235 $X2=15.345 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%VGND 1 2 3 4 5 6 7 8 25 29 33 37 41 45 49
+ 52 53 55 56 57 59 61 67 79 93 97 107 108 112 118 121 131 134
c214 108 0 2.71124e-20 $X=15.41 $Y=0
c215 52 0 1.39584e-19 $X=6.385 $Y=0
c216 41 0 1.51196e-19 $X=10.635 $Y=0.36
c217 37 0 1.59387e-19 $X=6.47 $Y=0.36
r218 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.95 $Y=0
+ $X2=14.95 $Y2=0
r219 131 132 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r220 121 122 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r221 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r222 113 119 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.61 $Y2=0
r223 112 115 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.38
r224 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r225 108 135 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.41 $Y=0
+ $X2=14.95 $Y2=0
r226 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.41 $Y=0
+ $X2=15.41 $Y2=0
r227 105 134 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=15.04 $Y=0
+ $X2=14.895 $Y2=0
r228 105 107 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=15.04 $Y=0
+ $X2=15.41 $Y2=0
r229 104 135 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=0
+ $X2=14.95 $Y2=0
r230 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.49 $Y=0
+ $X2=14.49 $Y2=0
r231 101 104 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=14.49 $Y2=0
r232 101 132 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=13.11 $Y2=0
r233 100 103 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=13.57 $Y=0
+ $X2=14.49 $Y2=0
r234 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r235 98 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.43 $Y=0
+ $X2=13.265 $Y2=0
r236 98 100 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=13.43 $Y=0
+ $X2=13.57 $Y2=0
r237 97 134 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=14.75 $Y=0
+ $X2=14.895 $Y2=0
r238 97 103 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=14.75 $Y=0
+ $X2=14.49 $Y2=0
r239 96 132 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=13.11 $Y2=0
r240 95 96 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r241 93 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.1 $Y=0
+ $X2=13.265 $Y2=0
r242 93 95 149.401 $w=1.68e-07 $l=2.29e-06 $layer=LI1_cond $X=13.1 $Y=0
+ $X2=10.81 $Y2=0
r243 92 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=10.81 $Y2=0
r244 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r245 89 92 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=10.35 $Y2=0
r246 89 126 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=8.51 $Y2=0
r247 88 91 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=8.97 $Y=0
+ $X2=10.35 $Y2=0
r248 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r249 86 88 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.675 $Y=0 $X2=8.97
+ $Y2=0
r250 85 126 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.51 $Y2=0
r251 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r252 82 85 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=8.05 $Y2=0
r253 81 84 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.67 $Y=0 $X2=8.05
+ $Y2=0
r254 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r255 79 128 11.3748 $w=3.83e-07 $l=3.8e-07 $layer=LI1_cond $X=8.482 $Y=0
+ $X2=8.482 $Y2=0.38
r256 79 86 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=8.482 $Y=0
+ $X2=8.675 $Y2=0
r257 79 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r258 79 84 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=8.29 $Y=0 $X2=8.05
+ $Y2=0
r259 78 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r260 78 122 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=3.91 $Y2=0
r261 77 78 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r262 75 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.95 $Y=0
+ $X2=3.785 $Y2=0
r263 75 77 147.444 $w=1.68e-07 $l=2.26e-06 $layer=LI1_cond $X=3.95 $Y=0 $X2=6.21
+ $Y2=0
r264 74 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r265 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r266 71 74 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.45 $Y2=0
r267 71 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.61 $Y2=0
r268 70 73 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r269 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r270 68 118 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.805 $Y=0
+ $X2=1.68 $Y2=0
r271 68 70 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.805 $Y=0
+ $X2=2.07 $Y2=0
r272 67 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.62 $Y=0
+ $X2=3.785 $Y2=0
r273 67 73 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.62 $Y=0 $X2=3.45
+ $Y2=0
r274 61 112 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.705 $Y2=0
r275 59 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r276 57 61 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.515 $Y2=0
r277 57 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r278 55 91 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=10.41 $Y=0 $X2=10.35
+ $Y2=0
r279 55 56 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=10.41 $Y=0
+ $X2=10.565 $Y2=0
r280 54 95 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=10.72 $Y=0 $X2=10.81
+ $Y2=0
r281 54 56 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=10.72 $Y=0
+ $X2=10.565 $Y2=0
r282 52 77 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.385 $Y=0
+ $X2=6.21 $Y2=0
r283 52 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.385 $Y=0 $X2=6.47
+ $Y2=0
r284 51 81 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.555 $Y=0
+ $X2=6.67 $Y2=0
r285 51 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=0 $X2=6.47
+ $Y2=0
r286 47 134 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=14.895 $Y=0.085
+ $X2=14.895 $Y2=0
r287 47 49 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=14.895 $Y=0.085
+ $X2=14.895 $Y2=0.38
r288 43 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.265 $Y=0.085
+ $X2=13.265 $Y2=0
r289 43 45 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=13.265 $Y=0.085
+ $X2=13.265 $Y2=0.38
r290 39 56 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=10.565 $Y=0.085
+ $X2=10.565 $Y2=0
r291 39 41 10.2233 $w=3.08e-07 $l=2.75e-07 $layer=LI1_cond $X=10.565 $Y=0.085
+ $X2=10.565 $Y2=0.36
r292 35 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=0.085
+ $X2=6.47 $Y2=0
r293 35 37 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.47 $Y=0.085
+ $X2=6.47 $Y2=0.36
r294 31 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.785 $Y=0.085
+ $X2=3.785 $Y2=0
r295 31 33 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.785 $Y=0.085
+ $X2=3.785 $Y2=0.36
r296 27 118 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=0.085
+ $X2=1.68 $Y2=0
r297 27 29 17.7476 $w=2.48e-07 $l=3.85e-07 $layer=LI1_cond $X=1.68 $Y=0.085
+ $X2=1.68 $Y2=0.47
r298 26 112 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=0.705 $Y2=0
r299 25 118 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.555 $Y=0
+ $X2=1.68 $Y2=0
r300 25 26 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.555 $Y=0
+ $X2=0.895 $Y2=0
r301 8 49 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=14.685
+ $Y=0.235 $X2=14.875 $Y2=0.38
r302 7 45 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=13.065
+ $Y=0.235 $X2=13.265 $Y2=0.38
r303 6 41 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=10.44
+ $Y=0.235 $X2=10.635 $Y2=0.36
r304 5 128 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=8.33
+ $Y=0.235 $X2=8.455 $Y2=0.38
r305 4 37 182 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_NDIFF $count=1 $X=6.135
+ $Y=0.235 $X2=6.47 $Y2=0.36
r306 3 33 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=3.59
+ $Y=0.235 $X2=3.785 $Y2=0.36
r307 2 29 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.72 $Y2=0.47
r308 1 115 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_1353_47# 1 2 7 11 16
r23 14 16 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=6.94 $Y=0.36
+ $X2=7.105 $Y2=0.36
r24 9 11 7.10956 $w=1.93e-07 $l=1.25e-07 $layer=LI1_cond $X=7.947 $Y=0.425
+ $X2=7.947 $Y2=0.55
r25 7 9 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=7.85 $Y=0.34
+ $X2=7.947 $Y2=0.425
r26 7 16 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=7.85 $Y=0.34
+ $X2=7.105 $Y2=0.34
r27 2 11 182 $w=1.7e-07 $l=3.86814e-07 $layer=licon1_NDIFF $count=1 $X=7.775
+ $Y=0.235 $X2=7.935 $Y2=0.55
r28 1 14 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=6.765
+ $Y=0.235 $X2=6.94 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_2216_47# 1 2 7 10 12
r22 10 12 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=12.125 $Y=0.34
+ $X2=11.38 $Y2=0.34
r23 7 12 5.98033 $w=2.08e-07 $l=1.05e-07 $layer=LI1_cond $X=11.275 $Y=0.36
+ $X2=11.38 $Y2=0.36
r24 7 9 3.48571 $w=2.1e-07 $l=6e-08 $layer=LI1_cond $X=11.275 $Y=0.36 $X2=11.215
+ $Y2=0.36
r25 2 10 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=12.075
+ $Y=0.235 $X2=12.21 $Y2=0.42
r26 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=11.08
+ $Y=0.235 $X2=11.215 $Y2=0.38
.ends

