* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__mux2_2 A0 A1 S VGND VNB VPB VPWR X
X0 a_606_369# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X1 a_502_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_318_369# A1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X3 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 a_79_21# A0 a_606_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X5 VPWR a_280_21# a_318_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X6 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND S a_280_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR S a_280_21# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_79_21# A1 a_502_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_280_21# a_310_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_310_47# A0 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
