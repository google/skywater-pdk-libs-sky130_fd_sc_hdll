* File: sky130_fd_sc_hdll__a21oi_2.pex.spice
* Created: Thu Aug 27 18:53:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A21OI_2%A2 1 3 6 8 10 11 13 14 18 21 25
c76 18 0 2.26013e-19 $X=1.92 $Y=1.16
c77 11 0 4.91474e-21 $X=1.945 $Y=1.41
r78 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.4
+ $Y=1.16 $X2=0.4 $Y2=1.16
r79 21 31 1.19608 $w=5.48e-07 $l=5.5e-08 $layer=LI1_cond $X=0.42 $Y=1.53
+ $X2=0.42 $Y2=1.585
r80 21 25 8.04635 $w=5.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.42 $Y=1.53
+ $X2=0.42 $Y2=1.16
r81 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.92
+ $Y=1.16 $X2=1.92 $Y2=1.16
r82 16 18 10.2952 $w=3.73e-07 $l=3.35e-07 $layer=LI1_cond $X=1.942 $Y=1.495
+ $X2=1.942 $Y2=1.16
r83 15 31 7.39687 $w=1.8e-07 $l=2.75e-07 $layer=LI1_cond $X=0.695 $Y=1.585
+ $X2=0.42 $Y2=1.585
r84 14 16 7.97274 $w=1.8e-07 $l=2.27594e-07 $layer=LI1_cond $X=1.755 $Y=1.585
+ $X2=1.942 $Y2=1.495
r85 14 15 65.3131 $w=1.78e-07 $l=1.06e-06 $layer=LI1_cond $X=1.755 $Y=1.585
+ $X2=0.695 $Y2=1.585
r86 11 19 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=1.945 $Y=1.41
+ $X2=1.945 $Y2=1.16
r87 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.945 $Y=1.41
+ $X2=1.945 $Y2=1.985
r88 8 19 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.86 $Y=0.995
+ $X2=1.945 $Y2=1.16
r89 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.86 $Y=0.995
+ $X2=1.86 $Y2=0.56
r90 4 24 35.7103 $w=3.32e-07 $l=1.94165e-07 $layer=POLY_cond $X=0.54 $Y=1.015
+ $X2=0.425 $Y2=1.16
r91 4 6 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.54 $Y=1.015
+ $X2=0.54 $Y2=0.56
r92 1 24 46.3299 $w=3.32e-07 $l=2.91548e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.425 $Y2=1.16
r93 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_2%A1 1 3 4 6 7 9 10 12 13 19 20 23
r47 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.475 $Y=1.202
+ $X2=1.5 $Y2=1.202
r48 18 20 6.97632 $w=3.8e-07 $l=5.5e-08 $layer=POLY_cond $X=1.42 $Y=1.202
+ $X2=1.475 $Y2=1.202
r49 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.42
+ $Y=1.16 $X2=1.42 $Y2=1.16
r50 16 18 53.9079 $w=3.8e-07 $l=4.25e-07 $layer=POLY_cond $X=0.995 $Y=1.202
+ $X2=1.42 $Y2=1.202
r51 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.97 $Y=1.202
+ $X2=0.995 $Y2=1.202
r52 13 19 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.25 $Y=1.16
+ $X2=1.42 $Y2=1.16
r53 13 23 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.25 $Y=1.16 $X2=1.15
+ $Y2=1.16
r54 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.5 $Y=0.995
+ $X2=1.5 $Y2=1.202
r55 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.5 $Y=0.995 $X2=1.5
+ $Y2=0.56
r56 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.475 $Y=1.41
+ $X2=1.475 $Y2=1.202
r57 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.475 $Y=1.41
+ $X2=1.475 $Y2=1.985
r58 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.995 $Y=1.41
+ $X2=0.995 $Y2=1.202
r59 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.995 $Y=1.41
+ $X2=0.995 $Y2=1.985
r60 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.97 $Y=0.995
+ $X2=0.97 $Y2=1.202
r61 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.97 $Y=0.995 $X2=0.97
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_2%B1 3 5 7 10 12 14 15 20 21 25
r52 20 21 8.85098 $w=4.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.285 $Y=1.16
+ $X2=3.285 $Y2=1.53
r53 20 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.12
+ $Y=1.16 $X2=3.12 $Y2=1.16
r54 18 19 3.4233 $w=3.52e-07 $l=2.5e-08 $layer=POLY_cond $X=2.86 $Y=1.212
+ $X2=2.885 $Y2=1.212
r55 17 18 60.9347 $w=3.52e-07 $l=4.45e-07 $layer=POLY_cond $X=2.415 $Y=1.212
+ $X2=2.86 $Y2=1.212
r56 16 17 3.4233 $w=3.52e-07 $l=2.5e-08 $layer=POLY_cond $X=2.39 $Y=1.212
+ $X2=2.415 $Y2=1.212
r57 15 25 27.9249 $w=2.9e-07 $l=1.35e-07 $layer=POLY_cond $X=2.985 $Y=1.16
+ $X2=3.12 $Y2=1.16
r58 15 19 15.3312 $w=3.52e-07 $l=1.23288e-07 $layer=POLY_cond $X=2.985 $Y=1.16
+ $X2=2.885 $Y2=1.212
r59 12 19 18.4407 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=2.885 $Y=1.41
+ $X2=2.885 $Y2=1.212
r60 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.885 $Y=1.41
+ $X2=2.885 $Y2=1.985
r61 8 18 22.7654 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=2.86 $Y=1.015
+ $X2=2.86 $Y2=1.212
r62 8 10 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.86 $Y=1.015
+ $X2=2.86 $Y2=0.56
r63 5 17 18.4407 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=2.415 $Y=1.41
+ $X2=2.415 $Y2=1.212
r64 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.415 $Y=1.41
+ $X2=2.415 $Y2=1.985
r65 1 16 22.7654 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=2.39 $Y=1.015
+ $X2=2.39 $Y2=1.212
r66 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.39 $Y=1.015
+ $X2=2.39 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_2%A_27_297# 1 2 3 4 13 15 17 21 23 25 26 27
+ 28 31 36
c62 3 0 1.09571e-19 $X=2.035 $Y=1.485
r63 29 31 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=3.237 $Y=2.285
+ $X2=3.237 $Y2=1.96
r64 27 29 7.42255 $w=1.8e-07 $l=1.91792e-07 $layer=LI1_cond $X=3.085 $Y=2.375
+ $X2=3.237 $Y2=2.285
r65 27 28 45.596 $w=1.78e-07 $l=7.4e-07 $layer=LI1_cond $X=3.085 $Y=2.375
+ $X2=2.345 $Y2=2.375
r66 26 28 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.18 $Y=2.285
+ $X2=2.345 $Y2=2.375
r67 25 38 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=2.025 $X2=2.18
+ $Y2=1.94
r68 25 26 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.18 $Y=2.025
+ $X2=2.18 $Y2=2.285
r69 24 36 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.32 $Y=1.94
+ $X2=1.235 $Y2=1.98
r70 23 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=1.94
+ $X2=2.18 $Y2=1.94
r71 23 24 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.015 $Y=1.94
+ $X2=1.32 $Y2=1.94
r72 19 36 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.235 $Y=2.105
+ $X2=1.235 $Y2=1.98
r73 19 21 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.235 $Y=2.105
+ $X2=1.235 $Y2=2.3
r74 18 34 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=0.37 $Y=1.98 $X2=0.24
+ $Y2=1.98
r75 17 36 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=1.98 $X2=1.235
+ $Y2=1.98
r76 17 18 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=1.15 $Y=1.98
+ $X2=0.37 $Y2=1.98
r77 13 34 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=2.105
+ $X2=0.24 $Y2=1.98
r78 13 15 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=0.24 $Y=2.105
+ $X2=0.24 $Y2=2.3
r79 4 31 300 $w=1.7e-07 $l=5.84808e-07 $layer=licon1_PDIFF $count=2 $X=2.975
+ $Y=1.485 $X2=3.22 $Y2=1.96
r80 3 38 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=2.035
+ $Y=1.485 $X2=2.18 $Y2=2.02
r81 2 36 600 $w=1.7e-07 $l=5.24667e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.485 $X2=1.235 $Y2=1.94
r82 2 21 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.485 $X2=1.235 $Y2=2.3
r83 1 34 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=1.96
r84 1 15 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_2%VPWR 1 2 9 12 13 14 16 29 30 33
c55 2 0 1.16442e-19 $X=1.565 $Y=1.485
r56 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r57 33 36 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=0.73 $Y=2.36
+ $X2=0.73 $Y2=2.72
r58 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r59 27 30 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r60 26 29 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r61 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r62 24 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r63 24 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r64 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r65 21 36 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.92 $Y=2.72 $X2=0.73
+ $Y2=2.72
r66 21 23 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.92 $Y=2.72 $X2=1.61
+ $Y2=2.72
r67 16 36 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.54 $Y=2.72 $X2=0.73
+ $Y2=2.72
r68 16 18 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.54 $Y=2.72
+ $X2=0.23 $Y2=2.72
r69 14 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r70 14 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r71 12 23 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.625 $Y=2.72
+ $X2=1.61 $Y2=2.72
r72 12 13 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=2.72
+ $X2=1.71 $Y2=2.72
r73 11 26 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.795 $Y=2.72
+ $X2=2.07 $Y2=2.72
r74 11 13 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=2.72
+ $X2=1.71 $Y2=2.72
r75 7 13 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=2.635 $X2=1.71
+ $Y2=2.72
r76 7 9 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.71 $Y=2.635
+ $X2=1.71 $Y2=2.36
r77 2 9 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=1.565
+ $Y=1.485 $X2=1.71 $Y2=2.36
r78 1 33 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.485 $X2=0.755 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_2%Y 1 2 3 10 13 16 19 26 27 28 31
c48 27 0 4.91474e-21 $X=2.637 $Y=1.33
r49 28 31 3.24125 $w=3.18e-07 $l=9e-08 $layer=LI1_cond $X=2.705 $Y=0.51
+ $X2=2.705 $Y2=0.42
r50 24 28 3.78145 $w=3.18e-07 $l=1.05e-07 $layer=LI1_cond $X=2.705 $Y=0.615
+ $X2=2.705 $Y2=0.51
r51 24 26 2.49074 $w=3.87e-07 $l=1.14039e-07 $layer=LI1_cond $X=2.705 $Y=0.615
+ $X2=2.637 $Y2=0.7
r52 19 22 9.91976 $w=3.93e-07 $l=3.4e-07 $layer=LI1_cond $X=1.202 $Y=0.36
+ $X2=1.202 $Y2=0.7
r53 16 27 9.21954 $w=3.48e-07 $l=2.8e-07 $layer=LI1_cond $X=2.69 $Y=1.61
+ $X2=2.69 $Y2=1.33
r54 13 27 6.63479 $w=4.53e-07 $l=2.27e-07 $layer=LI1_cond $X=2.637 $Y=1.103
+ $X2=2.637 $Y2=1.33
r55 12 26 2.49074 $w=3.87e-07 $l=8.5e-08 $layer=LI1_cond $X=2.637 $Y=0.785
+ $X2=2.637 $Y2=0.7
r56 12 13 8.35941 $w=4.53e-07 $l=3.18e-07 $layer=LI1_cond $X=2.637 $Y=0.785
+ $X2=2.637 $Y2=1.103
r57 11 22 5.70203 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=1.4 $Y=0.7 $X2=1.202
+ $Y2=0.7
r58 10 26 4.42191 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=2.41 $Y=0.7
+ $X2=2.637 $Y2=0.7
r59 10 11 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=2.41 $Y=0.7 $X2=1.4
+ $Y2=0.7
r60 3 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.505
+ $Y=1.485 $X2=2.65 $Y2=1.61
r61 2 31 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=2.465
+ $Y=0.235 $X2=2.65 $Y2=0.42
r62 2 26 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=2.465
+ $Y=0.235 $X2=2.65 $Y2=0.76
r63 1 22 182 $w=1.7e-07 $l=5.51883e-07 $layer=licon1_NDIFF $count=1 $X=1.045
+ $Y=0.235 $X2=1.235 $Y2=0.7
r64 1 19 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=1.045
+ $Y=0.235 $X2=1.235 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_2%VGND 1 2 3 10 12 14 16 18 20 28 38 45
r48 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r49 38 41 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=2.1 $Y=0 $X2=2.1
+ $Y2=0.36
r50 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r51 32 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r52 32 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r53 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r54 29 38 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.29 $Y=0 $X2=2.1
+ $Y2=0
r55 29 31 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.29 $Y=0 $X2=2.99
+ $Y2=0
r56 28 44 4.49945 $w=1.7e-07 $l=2.92e-07 $layer=LI1_cond $X=3.095 $Y=0 $X2=3.387
+ $Y2=0
r57 28 31 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.095 $Y=0 $X2=2.99
+ $Y2=0
r58 27 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r59 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r60 24 27 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r61 23 26 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r62 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r63 21 34 4.4461 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.197
+ $Y2=0
r64 21 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.69
+ $Y2=0
r65 20 38 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.91 $Y=0 $X2=2.1
+ $Y2=0
r66 20 26 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.91 $Y=0 $X2=1.61
+ $Y2=0
r67 18 24 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r68 18 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r69 14 44 3.26672 $w=3.3e-07 $l=1.64085e-07 $layer=LI1_cond $X=3.26 $Y=0.085
+ $X2=3.387 $Y2=0
r70 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.26 $Y=0.085
+ $X2=3.26 $Y2=0.38
r71 10 34 3.03143 $w=2.95e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.247 $Y=0.085
+ $X2=0.197 $Y2=0
r72 10 12 10.7431 $w=2.93e-07 $l=2.75e-07 $layer=LI1_cond $X=0.247 $Y=0.085
+ $X2=0.247 $Y2=0.36
r73 3 16 91 $w=1.7e-07 $l=3.90832e-07 $layer=licon1_NDIFF $count=2 $X=2.935
+ $Y=0.235 $X2=3.26 $Y2=0.38
r74 2 41 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=1.935
+ $Y=0.235 $X2=2.125 $Y2=0.36
r75 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.36
.ends

