# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__dlrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dlrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 0.955000 1.765000 1.325000 ;
    END
  END D
  PIN GATE
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.435000 1.625000 ;
    END
  END GATE
  PIN Q
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.765000 0.255000 6.295000 0.495000 ;
        RECT 5.815000 2.255000 6.295000 2.465000 ;
        RECT 5.820000 0.495000 6.295000 0.885000 ;
        RECT 5.895000 1.495000 6.295000 2.255000 ;
        RECT 6.065000 0.885000 6.295000 1.495000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.890000 0.995000 5.385000 1.325000 ;
    END
  END RESET_B
  PIN VGND
    ANTENNADIFFAREA  0.564250 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.440000 0.085000 ;
        RECT 0.565000  0.085000 0.895000 0.465000 ;
        RECT 2.025000  0.085000 2.355000 0.445000 ;
        RECT 3.870000  0.085000 4.200000 0.610000 ;
        RECT 5.320000  0.085000 5.595000 0.625000 ;
        RECT 5.320000  0.625000 5.650000 0.825000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.131000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 6.440000 2.805000 ;
        RECT 0.565000 2.135000 0.895000 2.635000 ;
        RECT 2.055000 1.835000 2.325000 2.635000 ;
        RECT 4.050000 2.135000 4.635000 2.635000 ;
        RECT 5.345000 1.885000 5.675000 2.150000 ;
        RECT 5.345000 2.150000 5.645000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 1.795000 0.775000 1.965000 ;
      RECT 0.085000 1.965000 0.395000 2.465000 ;
      RECT 0.225000 0.280000 0.395000 0.635000 ;
      RECT 0.225000 0.635000 0.775000 0.805000 ;
      RECT 0.605000 0.805000 0.775000 1.070000 ;
      RECT 0.605000 1.070000 0.895000 1.400000 ;
      RECT 0.605000 1.400000 0.775000 1.795000 ;
      RECT 1.065000 0.280000 1.235000 1.685000 ;
      RECT 1.065000 1.685000 1.335000 2.465000 ;
      RECT 1.555000 1.495000 2.115000 1.665000 ;
      RECT 1.555000 1.665000 1.885000 2.465000 ;
      RECT 1.660000 0.345000 1.855000 0.615000 ;
      RECT 1.660000 0.615000 2.115000 0.765000 ;
      RECT 1.660000 0.765000 2.535000 0.785000 ;
      RECT 1.945000 0.785000 2.535000 1.095000 ;
      RECT 1.945000 1.095000 2.115000 1.495000 ;
      RECT 2.445000 1.265000 2.955000 1.685000 ;
      RECT 2.780000 0.735000 3.295000 1.095000 ;
      RECT 3.020000 2.165000 3.850000 2.385000 ;
      RECT 3.040000 0.280000 3.660000 0.565000 ;
      RECT 3.125000 1.095000 3.295000 1.575000 ;
      RECT 3.125000 1.575000 3.510000 1.995000 ;
      RECT 3.490000 0.565000 3.660000 0.995000 ;
      RECT 3.490000 0.995000 4.380000 1.165000 ;
      RECT 3.680000 1.165000 4.380000 1.325000 ;
      RECT 3.680000 1.325000 3.850000 2.165000 ;
      RECT 4.020000 1.535000 5.725000 1.705000 ;
      RECT 4.020000 1.705000 5.170000 1.865000 ;
      RECT 4.455000 0.255000 4.785000 0.825000 ;
      RECT 4.550000 0.825000 4.720000 1.535000 ;
      RECT 4.885000 1.865000 5.170000 2.465000 ;
      RECT 5.555000 1.055000 5.895000 1.325000 ;
      RECT 5.555000 1.325000 5.725000 1.535000 ;
    LAYER mcon ;
      RECT 0.605000 1.445000 0.775000 1.615000 ;
      RECT 1.115000 1.785000 1.285000 1.955000 ;
      RECT 2.725000 1.445000 2.895000 1.615000 ;
      RECT 3.280000 1.785000 3.450000 1.955000 ;
    LAYER met1 ;
      RECT 0.545000 1.415000 0.835000 1.460000 ;
      RECT 0.545000 1.460000 2.955000 1.600000 ;
      RECT 0.545000 1.600000 0.835000 1.645000 ;
      RECT 1.055000 1.755000 1.345000 1.800000 ;
      RECT 1.055000 1.800000 3.510000 1.940000 ;
      RECT 1.055000 1.940000 1.345000 1.985000 ;
      RECT 2.665000 1.415000 2.955000 1.460000 ;
      RECT 2.665000 1.600000 2.955000 1.645000 ;
      RECT 3.220000 1.755000 3.510000 1.800000 ;
      RECT 3.220000 1.940000 3.510000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlrtp_1
