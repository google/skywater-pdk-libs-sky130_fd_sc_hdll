* NGSPICE file created from sky130_fd_sc_hdll__o211a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 a_225_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=4.875e+11p pd=4.1e+06u as=4.4525e+11p ps=3.97e+06u
M1001 a_79_21# C1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=7.7e+11p pd=5.54e+06u as=1.07e+12p ps=8.14e+06u
M1002 VPWR B1 a_79_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_540_47# B1 a_225_47# VNB nshort w=650000u l=150000u
+  ad=3.64e+11p pd=2.42e+06u as=0p ps=0u
M1004 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1005 a_79_21# A2 a_315_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.45e+11p ps=2.69e+06u
M1006 a_79_21# C1 a_540_47# VNB nshort w=650000u l=150000u
+  ad=2.275e+11p pd=2e+06u as=0p ps=0u
M1007 a_315_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1009 VGND A1 a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

