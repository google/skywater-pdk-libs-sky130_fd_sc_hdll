* File: sky130_fd_sc_hdll__o32ai_1.pex.spice
* Created: Wed Sep  2 08:47:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O32AI_1%B1 1 3 4 6 7 8
r23 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r24 7 8 13.2318 $w=2.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.225 $Y=0.85
+ $X2=0.225 $Y2=1.16
r25 4 12 40.1292 $w=4.26e-07 $l=2.36525e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.352 $Y2=1.16
r26 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r27 1 12 44.7281 $w=4.26e-07 $l=3.13449e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.352 $Y2=1.16
r28 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_1%B2 1 3 4 6 7 16
r28 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.005
+ $Y=1.16 $X2=1.005 $Y2=1.16
r29 7 16 0.0964579 $w=6.18e-07 $l=5e-09 $layer=LI1_cond $X=1.15 $Y=1.305
+ $X2=1.155 $Y2=1.305
r30 7 11 2.79728 $w=6.18e-07 $l=1.45e-07 $layer=LI1_cond $X=1.15 $Y=1.305
+ $X2=1.005 $Y2=1.305
r31 4 10 38.5363 $w=3.15e-07 $l=1.96074e-07 $layer=POLY_cond $X=1.045 $Y=0.995
+ $X2=0.977 $Y2=1.16
r32 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.045 $Y=0.995
+ $X2=1.045 $Y2=0.56
r33 1 10 47.0331 $w=3.15e-07 $l=2.83725e-07 $layer=POLY_cond $X=0.905 $Y=1.41
+ $X2=0.977 $Y2=1.16
r34 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.905 $Y=1.41
+ $X2=0.905 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_1%A3 1 3 4 6 7 15
r26 7 15 0.964579 $w=6.18e-07 $l=5e-08 $layer=LI1_cond $X=1.565 $Y=1.305
+ $X2=1.615 $Y2=1.305
r27 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.565
+ $Y=1.16 $X2=1.565 $Y2=1.16
r28 4 10 49.9093 $w=2.71e-07 $l=2.7157e-07 $layer=POLY_cond $X=1.6 $Y=1.41
+ $X2=1.555 $Y2=1.16
r29 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.6 $Y=1.41 $X2=1.6
+ $Y2=1.985
r30 1 10 38.8824 $w=2.71e-07 $l=1.96914e-07 $layer=POLY_cond $X=1.485 $Y=0.995
+ $X2=1.555 $Y2=1.16
r31 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.485 $Y=0.995
+ $X2=1.485 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_1%A2 1 3 4 6 7 8 9 10
r31 9 10 13.5114 $w=2.88e-07 $l=3.4e-07 $layer=LI1_cond $X=2.06 $Y=1.87 $X2=2.06
+ $Y2=2.21
r32 8 9 13.5114 $w=2.88e-07 $l=3.4e-07 $layer=LI1_cond $X=2.06 $Y=1.53 $X2=2.06
+ $Y2=1.87
r33 7 8 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.06 $Y=1.16 $X2=2.06
+ $Y2=1.53
r34 7 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.12
+ $Y=1.16 $X2=2.12 $Y2=1.16
r35 4 16 38.7084 $w=3.43e-07 $l=2.14942e-07 $layer=POLY_cond $X=2.26 $Y=0.995
+ $X2=2.145 $Y2=1.16
r36 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.26 $Y=0.995 $X2=2.26
+ $Y2=0.56
r37 1 16 45.964 $w=3.43e-07 $l=2.91548e-07 $layer=POLY_cond $X=2.235 $Y=1.41
+ $X2=2.145 $Y2=1.16
r38 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.235 $Y=1.41
+ $X2=2.235 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_1%A1 1 3 4 6 7 11 15
r20 11 15 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.8 $Y=1.16 $X2=2.55
+ $Y2=1.16
r21 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.8
+ $Y=1.16 $X2=2.8 $Y2=1.16
r22 7 15 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=2.525 $Y=1.16
+ $X2=2.55 $Y2=1.16
r23 4 10 45.964 $w=3.43e-07 $l=2.91548e-07 $layer=POLY_cond $X=2.705 $Y=1.41
+ $X2=2.795 $Y2=1.16
r24 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.705 $Y=1.41
+ $X2=2.705 $Y2=1.985
r25 1 10 38.7084 $w=3.43e-07 $l=2.14942e-07 $layer=POLY_cond $X=2.68 $Y=0.995
+ $X2=2.795 $Y2=1.16
r26 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.68 $Y=0.995 $X2=2.68
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_1%VPWR 1 2 7 9 13 15 19 21 34
r34 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r35 28 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r36 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r37 25 28 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r38 24 27 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r39 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r40 22 30 4.22982 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.36 $Y=2.72 $X2=0.18
+ $Y2=2.72
r41 22 24 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.36 $Y=2.72
+ $X2=0.69 $Y2=2.72
r42 21 33 5.00668 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=2.785 $Y=2.72
+ $X2=3.002 $Y2=2.72
r43 21 27 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.785 $Y=2.72
+ $X2=2.53 $Y2=2.72
r44 19 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r45 19 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r46 15 18 22.3903 $w=3.48e-07 $l=6.8e-07 $layer=LI1_cond $X=2.96 $Y=1.66
+ $X2=2.96 $Y2=2.34
r47 13 33 2.93018 $w=3.5e-07 $l=1.03899e-07 $layer=LI1_cond $X=2.96 $Y=2.635
+ $X2=3.002 $Y2=2.72
r48 13 18 9.71345 $w=3.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.96 $Y=2.635
+ $X2=2.96 $Y2=2.34
r49 9 12 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.225 $Y=1.66
+ $X2=0.225 $Y2=2.34
r50 7 30 3.05487 $w=2.7e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.225 $Y=2.635
+ $X2=0.18 $Y2=2.72
r51 7 12 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.225 $Y=2.635
+ $X2=0.225 $Y2=2.34
r52 2 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.795
+ $Y=1.485 $X2=2.94 $Y2=2.34
r53 2 15 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.795
+ $Y=1.485 $X2=2.94 $Y2=1.66
r54 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r55 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_1%Y 1 2 11 13 15 16 30
r29 16 30 0.263841 $w=6.78e-07 $l=1.5e-08 $layer=LI1_cond $X=1.17 $Y=2.125
+ $X2=1.155 $Y2=2.125
r30 15 30 0.0879469 $w=6.78e-07 $l=5e-09 $layer=LI1_cond $X=1.15 $Y=2.125
+ $X2=1.155 $Y2=2.125
r31 15 27 0.175894 $w=6.78e-07 $l=1e-08 $layer=LI1_cond $X=1.15 $Y=2.125
+ $X2=1.14 $Y2=2.125
r32 13 24 2.30831 $w=6.8e-07 $l=1.1e-07 $layer=LI1_cond $X=0.64 $Y=2.125
+ $X2=0.75 $Y2=2.125
r33 13 27 6.15629 $w=6.78e-07 $l=3.5e-07 $layer=LI1_cond $X=0.79 $Y=2.125
+ $X2=1.14 $Y2=2.125
r34 13 24 0.703576 $w=6.78e-07 $l=4e-08 $layer=LI1_cond $X=0.79 $Y=2.125
+ $X2=0.75 $Y2=2.125
r35 8 13 36.6757 $w=3.08e-07 $l=9.6e-07 $layer=LI1_cond $X=0.64 $Y=0.825
+ $X2=0.64 $Y2=1.785
r36 8 11 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.64 $Y=0.74 $X2=0.73
+ $Y2=0.74
r37 2 27 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.995
+ $Y=1.485 $X2=1.14 $Y2=2
r38 1 11 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_1%A_27_47# 1 2 3 10 14 18
r31 23 24 11.0635 $w=3.73e-07 $l=3.6e-07 $layer=LI1_cond $X=1.252 $Y=0.38
+ $X2=1.252 $Y2=0.74
r32 16 18 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.47 $Y=0.655
+ $X2=2.47 $Y2=0.54
r33 15 24 5.38787 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=1.44 $Y=0.74
+ $X2=1.252 $Y2=0.74
r34 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.385 $Y=0.74
+ $X2=2.47 $Y2=0.655
r35 14 15 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=2.385 $Y=0.74
+ $X2=1.44 $Y2=0.74
r36 10 23 0.307318 $w=3.73e-07 $l=1e-08 $layer=LI1_cond $X=1.252 $Y=0.37
+ $X2=1.252 $Y2=0.38
r37 10 12 40.3355 $w=2.28e-07 $l=8.05e-07 $layer=LI1_cond $X=1.065 $Y=0.37
+ $X2=0.26 $Y2=0.37
r38 3 18 182 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.235 $X2=2.47 $Y2=0.54
r39 2 23 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.12
+ $Y=0.235 $X2=1.255 $Y2=0.38
r40 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_1%VGND 1 2 9 11 13 16 17 18 27 33
r38 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r39 30 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r40 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r41 27 32 5.08404 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.972
+ $Y2=0
r42 27 29 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.53
+ $Y2=0
r43 26 30 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r44 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r45 21 25 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r46 18 26 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r47 18 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r48 16 25 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.645 $Y=0 $X2=1.61
+ $Y2=0
r49 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.645 $Y=0 $X2=1.81
+ $Y2=0
r50 15 29 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=2.53
+ $Y2=0
r51 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=1.81
+ $Y2=0
r52 11 32 3.02572 $w=3.7e-07 $l=1.11781e-07 $layer=LI1_cond $X=2.91 $Y=0.085
+ $X2=2.972 $Y2=0
r53 11 13 9.1884 $w=3.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.91 $Y=0.085
+ $X2=2.91 $Y2=0.38
r54 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=0.085 $X2=1.81
+ $Y2=0
r55 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.81 $Y=0.085
+ $X2=1.81 $Y2=0.38
r56 2 13 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=2.755
+ $Y=0.235 $X2=2.91 $Y2=0.38
r57 1 9 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.235 $X2=1.81 $Y2=0.38
.ends

