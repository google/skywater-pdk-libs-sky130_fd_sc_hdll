# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nor4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.075000 1.075000 10.010000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.650000 1.075000 7.805000 1.285000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.445000 1.365000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.075000 1.395000 1.325000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  2.374000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.940000 1.415000 3.435000 1.705000 ;
        RECT 2.035000 0.255000 2.415000 0.725000 ;
        RECT 2.035000 0.725000 9.515000 0.905000 ;
        RECT 2.975000 0.255000 3.355000 0.725000 ;
        RECT 3.265000 0.905000 3.435000 1.415000 ;
        RECT 3.915000 0.255000 4.295000 0.725000 ;
        RECT 4.855000 0.255000 5.235000 0.725000 ;
        RECT 6.315000 0.255000 6.695000 0.725000 ;
        RECT 7.255000 0.255000 7.635000 0.725000 ;
        RECT 8.195000 0.255000 8.575000 0.725000 ;
        RECT 9.135000 0.255000 9.515000 0.725000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.085000  0.255000  0.445000 0.725000 ;
      RECT 0.085000  0.725000  0.835000 0.895000 ;
      RECT 0.085000  1.535000  0.835000 1.875000 ;
      RECT 0.085000  1.875000  3.825000 2.045000 ;
      RECT 0.085000  2.045000  0.365000 2.465000 ;
      RECT 0.535000  2.215000  0.915000 2.635000 ;
      RECT 0.665000  0.085000  0.835000 0.555000 ;
      RECT 0.665000  0.895000  0.835000 1.535000 ;
      RECT 1.005000  0.255000  1.385000 0.735000 ;
      RECT 1.005000  0.735000  1.735000 0.905000 ;
      RECT 1.005000  1.535000  1.735000 1.705000 ;
      RECT 1.565000  0.905000  1.735000 1.075000 ;
      RECT 1.565000  1.075000  3.095000 1.245000 ;
      RECT 1.565000  1.245000  1.735000 1.535000 ;
      RECT 1.615000  2.215000  3.825000 2.295000 ;
      RECT 1.615000  2.295000  5.695000 2.465000 ;
      RECT 1.695000  0.085000  1.865000 0.555000 ;
      RECT 2.635000  0.085000  2.805000 0.555000 ;
      RECT 3.575000  0.085000  3.745000 0.555000 ;
      RECT 3.655000  1.075000  5.405000 1.285000 ;
      RECT 3.655000  1.285000  3.825000 1.875000 ;
      RECT 4.045000  1.455000  7.595000 1.625000 ;
      RECT 4.045000  1.625000  4.255000 2.125000 ;
      RECT 4.475000  1.795000  4.725000 2.295000 ;
      RECT 4.515000  0.085000  4.685000 0.555000 ;
      RECT 4.945000  1.625000  5.195000 2.125000 ;
      RECT 5.415000  1.795000  5.695000 2.295000 ;
      RECT 5.455000  0.085000  6.145000 0.555000 ;
      RECT 5.880000  1.795000  6.185000 2.295000 ;
      RECT 5.880000  2.295000  8.065000 2.465000 ;
      RECT 6.405000  1.625000  6.655000 2.125000 ;
      RECT 6.875000  1.795000  7.125000 2.295000 ;
      RECT 6.915000  0.085000  7.085000 0.555000 ;
      RECT 7.345000  1.625000  7.595000 2.125000 ;
      RECT 7.815000  1.455000 10.010000 1.625000 ;
      RECT 7.815000  1.625000  8.065000 2.295000 ;
      RECT 7.855000  0.085000  8.025000 0.555000 ;
      RECT 8.285000  1.795000  8.535000 2.635000 ;
      RECT 8.755000  1.625000  9.005000 2.465000 ;
      RECT 8.795000  0.085000  8.965000 0.555000 ;
      RECT 9.225000  1.795000  9.475000 2.635000 ;
      RECT 9.695000  1.625000 10.010000 2.465000 ;
      RECT 9.735000  0.085000 10.010000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4bb_4
