* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__or2b_2 A B_N VGND VNB VPB VPWR X
X0 a_228_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR B_N a_27_53# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X2 VGND a_228_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_228_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 X a_228_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_318_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X6 a_27_53# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 X a_228_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VGND a_27_53# a_228_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_228_297# a_27_53# a_318_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
.ends
