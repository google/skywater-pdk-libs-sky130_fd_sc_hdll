* File: sky130_fd_sc_hdll__o221a_2.pex.spice
* Created: Thu Aug 27 19:20:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O221A_2%C1 1 3 4 6 7 8 9 18
r33 12 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r34 9 18 0.823174 $w=3.48e-07 $l=2.5e-08 $layer=LI1_cond $X=0.205 $Y=1.15
+ $X2=0.23 $Y2=1.15
r35 7 12 48.6364 $w=3.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.555 $Y=1.15
+ $X2=0.26 $Y2=1.15
r36 7 8 4.60329 $w=3.5e-07 $l=1.19164e-07 $layer=POLY_cond $X=0.555 $Y=1.15
+ $X2=0.655 $Y2=1.192
r37 4 8 36.1676 $w=1.65e-07 $l=2.29159e-07 $layer=POLY_cond $X=0.68 $Y=0.975
+ $X2=0.655 $Y2=1.192
r38 4 6 133.353 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=0.68 $Y=0.975
+ $X2=0.68 $Y2=0.56
r39 1 8 36.1676 $w=1.65e-07 $l=2.18e-07 $layer=POLY_cond $X=0.655 $Y=1.41
+ $X2=0.655 $Y2=1.192
r40 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.655 $Y=1.41
+ $X2=0.655 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_2%B1 1 3 4 6 7 14
r32 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.1
+ $Y=1.16 $X2=1.1 $Y2=1.16
r33 7 14 4.15909 $w=1.98e-07 $l=7.5e-08 $layer=LI1_cond $X=1.175 $Y=1.175
+ $X2=1.1 $Y2=1.175
r34 4 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=1.185 $Y=1.41
+ $X2=1.125 $Y2=1.16
r35 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.185 $Y=1.41
+ $X2=1.185 $Y2=1.985
r36 1 10 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.15 $Y=0.995
+ $X2=1.125 $Y2=1.16
r37 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.15 $Y=0.995 $X2=1.15
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_2%B2 1 3 4 6 7 8 18
r32 8 18 0.449004 $w=3.83e-07 $l=1.5e-08 $layer=LI1_cond $X=1.712 $Y=1.545
+ $X2=1.712 $Y2=1.53
r33 7 18 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=1.712 $Y=1.16
+ $X2=1.712 $Y2=1.53
r34 7 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.16 $X2=1.69 $Y2=1.16
r35 4 12 46.3664 $w=3.31e-07 $l=2.88097e-07 $layer=POLY_cond $X=1.61 $Y=1.41
+ $X2=1.692 $Y2=1.16
r36 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.61 $Y=1.41 $X2=1.61
+ $Y2=1.985
r37 1 12 38.6069 $w=3.31e-07 $l=2.11849e-07 $layer=POLY_cond $X=1.585 $Y=0.995
+ $X2=1.692 $Y2=1.16
r38 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.585 $Y=0.995
+ $X2=1.585 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_2%A2 1 3 4 6 7 8
r31 7 8 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.425 $Y=1.16
+ $X2=2.425 $Y2=1.53
r32 7 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.4 $Y=1.16
+ $X2=2.4 $Y2=1.16
r33 4 12 39.1188 $w=3.74e-07 $l=2.22486e-07 $layer=POLY_cond $X=2.61 $Y=0.995
+ $X2=2.475 $Y2=1.16
r34 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.61 $Y=0.995 $X2=2.61
+ $Y2=0.56
r35 1 12 45.2339 $w=3.74e-07 $l=3e-07 $layer=POLY_cond $X=2.585 $Y=1.41
+ $X2=2.475 $Y2=1.16
r36 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.585 $Y=1.41
+ $X2=2.585 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_2%A1 1 3 4 6 7 14
c32 1 0 1.87094e-19 $X=2.995 $Y=1.41
r33 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.03
+ $Y=1.16 $X2=3.03 $Y2=1.16
r34 7 14 10.8268 $w=2.08e-07 $l=2.05e-07 $layer=LI1_cond $X=3.235 $Y=1.18
+ $X2=3.03 $Y2=1.18
r35 4 10 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=3.08 $Y=0.995
+ $X2=3.055 $Y2=1.16
r36 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.08 $Y=0.995 $X2=3.08
+ $Y2=0.56
r37 1 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.995 $Y=1.41
+ $X2=3.055 $Y2=1.16
r38 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.995 $Y=1.41
+ $X2=2.995 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_2%A_38_47# 1 2 3 10 12 13 15 16 18 19 21 24
+ 28 30 31 32 35 37 38 41 42 43 45 51 54 55 59 65
c133 59 0 1.87094e-19 $X=3.71 $Y=1.16
r134 65 66 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.995 $Y=1.202
+ $X2=4.02 $Y2=1.202
r135 62 63 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.5 $Y=1.202
+ $X2=3.525 $Y2=1.202
r136 60 65 36.15 $w=3.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.71 $Y=1.202
+ $X2=3.995 $Y2=1.202
r137 60 63 23.4658 $w=3.8e-07 $l=1.85e-07 $layer=POLY_cond $X=3.71 $Y=1.202
+ $X2=3.525 $Y2=1.202
r138 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.71
+ $Y=1.16 $X2=3.71 $Y2=1.16
r139 56 59 5.54545 $w=2.08e-07 $l=1.05e-07 $layer=LI1_cond $X=3.605 $Y=1.18
+ $X2=3.71 $Y2=1.18
r140 53 55 8.87457 $w=5.88e-07 $l=1.05e-07 $layer=LI1_cond $X=2.35 $Y=2.17
+ $X2=2.455 $Y2=2.17
r141 53 54 19.9231 $w=5.88e-07 $l=6.5e-07 $layer=LI1_cond $X=2.35 $Y=2.17
+ $X2=1.7 $Y2=2.17
r142 44 56 0.430812 $w=2.2e-07 $l=1.05e-07 $layer=LI1_cond $X=3.605 $Y=1.285
+ $X2=3.605 $Y2=1.18
r143 44 45 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=3.605 $Y=1.285
+ $X2=3.605 $Y2=1.455
r144 42 45 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.495 $Y=1.54
+ $X2=3.605 $Y2=1.455
r145 42 43 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.495 $Y=1.54
+ $X2=2.965 $Y2=1.54
r146 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.88 $Y=1.625
+ $X2=2.965 $Y2=1.54
r147 40 41 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.88 $Y=1.625
+ $X2=2.88 $Y2=1.875
r148 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.795 $Y=1.96
+ $X2=2.88 $Y2=1.875
r149 38 55 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.795 $Y=1.96
+ $X2=2.455 $Y2=1.96
r150 37 54 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.35 $Y=1.96
+ $X2=1.7 $Y2=1.96
r151 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.265 $Y=1.875
+ $X2=1.35 $Y2=1.96
r152 34 35 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.265 $Y=1.67
+ $X2=1.265 $Y2=1.875
r153 33 51 2.07418 $w=2.25e-07 $l=5.45119e-07 $layer=LI1_cond $X=0.765 $Y=1.557
+ $X2=0.25 $Y2=1.495
r154 32 34 6.9898 $w=2.25e-07 $l=1.49579e-07 $layer=LI1_cond $X=1.18 $Y=1.557
+ $X2=1.265 $Y2=1.67
r155 32 33 21.2562 $w=2.23e-07 $l=4.15e-07 $layer=LI1_cond $X=1.18 $Y=1.557
+ $X2=0.765 $Y2=1.557
r156 31 51 4.35802 $w=2.75e-07 $l=4.29273e-07 $layer=LI1_cond $X=0.655 $Y=1.445
+ $X2=0.25 $Y2=1.495
r157 30 31 33.5256 $w=2.18e-07 $l=6.4e-07 $layer=LI1_cond $X=0.655 $Y=0.805
+ $X2=0.655 $Y2=1.445
r158 26 51 4.35802 $w=2.75e-07 $l=2.43926e-07 $layer=LI1_cond $X=0.415 $Y=1.67
+ $X2=0.25 $Y2=1.495
r159 26 28 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=0.415 $Y=1.67
+ $X2=0.415 $Y2=2.3
r160 22 30 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.335 $Y=0.72
+ $X2=0.655 $Y2=0.72
r161 22 24 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.335 $Y=0.635
+ $X2=0.335 $Y2=0.36
r162 19 66 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.02 $Y=0.995
+ $X2=4.02 $Y2=1.202
r163 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.02 $Y=0.995
+ $X2=4.02 $Y2=0.56
r164 16 65 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.995 $Y=1.41
+ $X2=3.995 $Y2=1.202
r165 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.995 $Y=1.41
+ $X2=3.995 $Y2=1.985
r166 13 63 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.525 $Y=1.41
+ $X2=3.525 $Y2=1.202
r167 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.525 $Y=1.41
+ $X2=3.525 $Y2=1.985
r168 10 62 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.5 $Y=0.995
+ $X2=3.5 $Y2=1.202
r169 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.5 $Y=0.995
+ $X2=3.5 $Y2=0.56
r170 3 53 150 $w=1.7e-07 $l=8.55132e-07 $layer=licon1_PDIFF $count=4 $X=1.7
+ $Y=1.485 $X2=2.35 $Y2=1.96
r171 2 51 400 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=0.23
+ $Y=1.485 $X2=0.415 $Y2=1.62
r172 2 28 400 $w=1.7e-07 $l=9.02773e-07 $layer=licon1_PDIFF $count=1 $X=0.23
+ $Y=1.485 $X2=0.415 $Y2=2.3
r173 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.19
+ $Y=0.235 $X2=0.335 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_2%VPWR 1 2 3 12 16 18 20 23 24 26 27 28 40
+ 46 50
r68 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r69 43 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r70 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r71 40 45 5.10308 $w=1.7e-07 $l=2.92e-07 $layer=LI1_cond $X=4.015 $Y=2.72
+ $X2=4.307 $Y2=2.72
r72 40 42 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.015 $Y=2.72
+ $X2=3.91 $Y2=2.72
r73 39 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r74 38 39 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r75 36 39 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r76 35 38 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r77 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r78 32 36 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r79 32 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r80 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r81 28 50 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=2.72
+ $X2=0.23 $Y2=2.72
r82 26 38 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.145 $Y=2.72
+ $X2=2.99 $Y2=2.72
r83 26 27 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.145 $Y=2.72
+ $X2=3.26 $Y2=2.72
r84 25 42 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.375 $Y=2.72
+ $X2=3.91 $Y2=2.72
r85 25 27 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.375 $Y=2.72
+ $X2=3.26 $Y2=2.72
r86 23 31 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.8 $Y=2.72 $X2=0.69
+ $Y2=2.72
r87 23 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.8 $Y=2.72
+ $X2=0.905 $Y2=2.72
r88 22 35 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.01 $Y=2.72
+ $X2=1.15 $Y2=2.72
r89 22 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.01 $Y=2.72
+ $X2=0.905 $Y2=2.72
r90 18 45 3.18069 $w=3.9e-07 $l=1.32868e-07 $layer=LI1_cond $X=4.21 $Y=2.635
+ $X2=4.307 $Y2=2.72
r91 18 20 9.89919 $w=3.88e-07 $l=3.35e-07 $layer=LI1_cond $X=4.21 $Y=2.635
+ $X2=4.21 $Y2=2.3
r92 14 27 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.26 $Y=2.635
+ $X2=3.26 $Y2=2.72
r93 14 16 33.8217 $w=2.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.26 $Y=2.635
+ $X2=3.26 $Y2=1.96
r94 10 24 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.905 $Y=2.635
+ $X2=0.905 $Y2=2.72
r95 10 12 32.7446 $w=2.08e-07 $l=6.2e-07 $layer=LI1_cond $X=0.905 $Y=2.635
+ $X2=0.905 $Y2=2.015
r96 3 20 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.085
+ $Y=1.485 $X2=4.23 $Y2=2.3
r97 2 16 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.085
+ $Y=1.485 $X2=3.23 $Y2=1.96
r98 1 12 300 $w=1.7e-07 $l=6.13433e-07 $layer=licon1_PDIFF $count=2 $X=0.745
+ $Y=1.485 $X2=0.925 $Y2=2.015
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_2%X 1 2 9 11 13 15 17 18 22 25 28
r46 25 28 0.185878 $w=3.08e-07 $l=5e-09 $layer=LI1_cond $X=4.335 $Y=1.875
+ $X2=4.335 $Y2=1.87
r47 22 25 2.69138 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.335 $Y=1.96
+ $X2=4.335 $Y2=1.875
r48 22 28 1.48702 $w=3.08e-07 $l=4e-08 $layer=LI1_cond $X=4.335 $Y=1.83
+ $X2=4.335 $Y2=1.87
r49 21 22 34.3874 $w=3.08e-07 $l=9.25e-07 $layer=LI1_cond $X=4.335 $Y=0.905
+ $X2=4.335 $Y2=1.83
r50 17 21 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=4.18 $Y=0.82
+ $X2=4.335 $Y2=0.905
r51 17 18 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.18 $Y=0.82
+ $X2=3.925 $Y2=0.82
r52 16 20 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.845 $Y=1.96
+ $X2=3.695 $Y2=1.96
r53 15 22 4.90781 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.18 $Y=1.96
+ $X2=4.335 $Y2=1.96
r54 15 16 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.18 $Y=1.96
+ $X2=3.845 $Y2=1.96
r55 11 20 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.695 $Y=2.045
+ $X2=3.695 $Y2=1.96
r56 11 13 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=3.695 $Y=2.045
+ $X2=3.695 $Y2=2.3
r57 7 18 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=3.735 $Y=0.735
+ $X2=3.925 $Y2=0.82
r58 7 9 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=3.735 $Y=0.735
+ $X2=3.735 $Y2=0.39
r59 2 20 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=3.615
+ $Y=1.485 $X2=3.76 $Y2=1.96
r60 2 13 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.615
+ $Y=1.485 $X2=3.76 $Y2=2.3
r61 1 9 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.575
+ $Y=0.235 $X2=3.76 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_2%A_151_47# 1 2 11
r17 8 11 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.89 $Y=0.38 $X2=1.83
+ $Y2=0.38
r18 2 11 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=1.66
+ $Y=0.235 $X2=1.83 $Y2=0.38
r19 1 8 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.755
+ $Y=0.235 $X2=0.89 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_2%A_245_47# 1 2 7 11 15 17
r36 13 15 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=2.795 $Y=0.735
+ $X2=2.795 $Y2=0.39
r37 11 13 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=2.605 $Y=0.82
+ $X2=2.795 $Y2=0.735
r38 11 17 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=2.605 $Y=0.82
+ $X2=1.57 $Y2=0.82
r39 7 17 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=1.44 $Y=0.775
+ $X2=1.57 $Y2=0.775
r40 7 9 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=1.44 $Y=0.775 $X2=1.36
+ $Y2=0.775
r41 2 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.685
+ $Y=0.235 $X2=2.82 $Y2=0.39
r42 1 9 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.225
+ $Y=0.235 $X2=1.36 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_2%VGND 1 2 3 12 16 20 23 24 26 27 28 29 30
+ 31 48 52
r63 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r64 45 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r65 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r66 42 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r67 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r68 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r69 39 52 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=0.23
+ $Y2=0
r70 38 39 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r71 34 38 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r72 34 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r73 31 52 0.00711354 $w=4.8e-07 $l=2.5e-08 $layer=MET1_cond $X=0.205 $Y=0
+ $X2=0.23 $Y2=0
r74 29 44 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.145 $Y=0 $X2=3.91
+ $Y2=0
r75 29 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.145 $Y=0 $X2=4.23
+ $Y2=0
r76 28 47 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=4.315 $Y=0 $X2=4.37
+ $Y2=0
r77 28 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.315 $Y=0 $X2=4.23
+ $Y2=0
r78 26 41 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.205 $Y=0 $X2=2.99
+ $Y2=0
r79 26 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.205 $Y=0 $X2=3.29
+ $Y2=0
r80 25 44 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.91
+ $Y2=0
r81 25 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.29
+ $Y2=0
r82 23 38 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.265 $Y=0 $X2=2.07
+ $Y2=0
r83 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.265 $Y=0 $X2=2.35
+ $Y2=0
r84 22 41 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.435 $Y=0 $X2=2.99
+ $Y2=0
r85 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=0 $X2=2.35
+ $Y2=0
r86 18 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.23 $Y=0.085
+ $X2=4.23 $Y2=0
r87 18 20 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.23 $Y=0.085
+ $X2=4.23 $Y2=0.39
r88 14 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.29 $Y=0.085
+ $X2=3.29 $Y2=0
r89 14 16 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.29 $Y=0.085
+ $X2=3.29 $Y2=0.39
r90 10 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.35 $Y=0.085
+ $X2=2.35 $Y2=0
r91 10 12 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.35 $Y=0.085
+ $X2=2.35 $Y2=0.39
r92 3 20 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.095
+ $Y=0.235 $X2=4.23 $Y2=0.39
r93 2 16 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.155
+ $Y=0.235 $X2=3.29 $Y2=0.39
r94 1 12 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.35 $Y2=0.39
.ends

