* File: sky130_fd_sc_hdll__o31ai_4.pxi.spice
* Created: Wed Sep  2 08:46:58 2020
* 
x_PM_SKY130_FD_SC_HDLL__O31AI_4%A1 N_A1_M1003_g N_A1_c_110_n N_A1_M1002_g
+ N_A1_M1014_g N_A1_c_111_n N_A1_M1006_g N_A1_M1015_g N_A1_c_112_n N_A1_M1013_g
+ N_A1_c_113_n N_A1_M1020_g N_A1_M1026_g A1 A1 A1 A1 N_A1_c_108_n A1 A1 A1
+ PM_SKY130_FD_SC_HDLL__O31AI_4%A1
x_PM_SKY130_FD_SC_HDLL__O31AI_4%A2 N_A2_M1008_g N_A2_c_198_n N_A2_M1001_g
+ N_A2_M1011_g N_A2_c_199_n N_A2_M1016_g N_A2_M1021_g N_A2_c_200_n N_A2_M1024_g
+ N_A2_c_201_n N_A2_M1031_g N_A2_M1029_g A2 A2 A2 A2 N_A2_c_197_n A2 A2 A2 A2
+ PM_SKY130_FD_SC_HDLL__O31AI_4%A2
x_PM_SKY130_FD_SC_HDLL__O31AI_4%A3 N_A3_M1000_g N_A3_c_292_n N_A3_M1005_g
+ N_A3_M1017_g N_A3_c_293_n N_A3_M1007_g N_A3_M1023_g N_A3_c_294_n N_A3_M1018_g
+ N_A3_c_295_n N_A3_M1028_g N_A3_M1027_g N_A3_c_288_n A3 A3 A3 A3 A3
+ N_A3_c_289_n N_A3_c_290_n A3 A3 A3 A3 A3 PM_SKY130_FD_SC_HDLL__O31AI_4%A3
x_PM_SKY130_FD_SC_HDLL__O31AI_4%B1 N_B1_M1004_g N_B1_c_363_n N_B1_M1010_g
+ N_B1_M1009_g N_B1_c_364_n N_B1_M1019_g N_B1_M1012_g N_B1_c_365_n N_B1_M1025_g
+ N_B1_M1022_g N_B1_c_366_n N_B1_M1030_g B1 B1 B1 N_B1_c_362_n B1 B1
+ PM_SKY130_FD_SC_HDLL__O31AI_4%B1
x_PM_SKY130_FD_SC_HDLL__O31AI_4%A_27_297# N_A_27_297#_M1002_s
+ N_A_27_297#_M1006_s N_A_27_297#_M1020_s N_A_27_297#_M1016_s
+ N_A_27_297#_M1031_s N_A_27_297#_c_428_n N_A_27_297#_c_429_n
+ N_A_27_297#_c_435_n N_A_27_297#_c_439_n N_A_27_297#_c_443_n
+ N_A_27_297#_c_447_n N_A_27_297#_c_448_n N_A_27_297#_c_458_n
+ N_A_27_297#_c_430_n N_A_27_297#_c_450_n N_A_27_297#_c_462_n
+ PM_SKY130_FD_SC_HDLL__O31AI_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__O31AI_4%VPWR N_VPWR_M1002_d N_VPWR_M1013_d
+ N_VPWR_M1010_s N_VPWR_M1025_s N_VPWR_c_511_n N_VPWR_c_512_n N_VPWR_c_513_n
+ N_VPWR_c_514_n N_VPWR_c_515_n N_VPWR_c_516_n N_VPWR_c_517_n N_VPWR_c_518_n
+ N_VPWR_c_519_n VPWR N_VPWR_c_520_n N_VPWR_c_510_n N_VPWR_c_522_n
+ N_VPWR_c_523_n PM_SKY130_FD_SC_HDLL__O31AI_4%VPWR
x_PM_SKY130_FD_SC_HDLL__O31AI_4%A_497_297# N_A_497_297#_M1001_d
+ N_A_497_297#_M1024_d N_A_497_297#_M1005_s N_A_497_297#_M1018_s
+ N_A_497_297#_c_623_n N_A_497_297#_c_636_n N_A_497_297#_c_624_n
+ N_A_497_297#_c_628_n N_A_497_297#_c_632_n N_A_497_297#_c_622_n
+ PM_SKY130_FD_SC_HDLL__O31AI_4%A_497_297#
x_PM_SKY130_FD_SC_HDLL__O31AI_4%Y N_Y_M1004_s N_Y_M1012_s N_Y_M1005_d
+ N_Y_M1007_d N_Y_M1028_d N_Y_M1019_d N_Y_M1030_d N_Y_c_722_n N_Y_c_690_n
+ N_Y_c_725_n N_Y_c_695_n Y Y Y Y Y Y Y Y Y Y Y N_Y_c_674_n Y Y Y Y Y
+ N_Y_c_675_n N_Y_c_676_n N_Y_c_677_n Y N_Y_c_678_n Y
+ PM_SKY130_FD_SC_HDLL__O31AI_4%Y
x_PM_SKY130_FD_SC_HDLL__O31AI_4%A_31_47# N_A_31_47#_M1003_d N_A_31_47#_M1014_d
+ N_A_31_47#_M1026_d N_A_31_47#_M1011_s N_A_31_47#_M1029_s N_A_31_47#_M1017_s
+ N_A_31_47#_M1027_s N_A_31_47#_M1009_d N_A_31_47#_M1022_d N_A_31_47#_c_753_n
+ N_A_31_47#_c_765_n N_A_31_47#_c_754_n N_A_31_47#_c_771_n N_A_31_47#_c_775_n
+ N_A_31_47#_c_779_n N_A_31_47#_c_788_n N_A_31_47#_c_792_n N_A_31_47#_c_796_n
+ N_A_31_47#_c_800_n N_A_31_47#_c_811_n N_A_31_47#_c_865_p N_A_31_47#_c_755_n
+ N_A_31_47#_c_824_n N_A_31_47#_c_869_p N_A_31_47#_c_756_n N_A_31_47#_c_757_n
+ N_A_31_47#_c_758_n N_A_31_47#_c_759_n N_A_31_47#_c_760_n N_A_31_47#_c_761_n
+ N_A_31_47#_c_762_n PM_SKY130_FD_SC_HDLL__O31AI_4%A_31_47#
x_PM_SKY130_FD_SC_HDLL__O31AI_4%VGND N_VGND_M1003_s N_VGND_M1015_s
+ N_VGND_M1008_d N_VGND_M1021_d N_VGND_M1000_d N_VGND_M1023_d N_VGND_c_903_n
+ N_VGND_c_904_n N_VGND_c_905_n N_VGND_c_906_n N_VGND_c_907_n N_VGND_c_908_n
+ N_VGND_c_909_n N_VGND_c_910_n N_VGND_c_911_n N_VGND_c_912_n N_VGND_c_913_n
+ N_VGND_c_914_n VGND N_VGND_c_915_n N_VGND_c_916_n N_VGND_c_917_n
+ N_VGND_c_918_n N_VGND_c_919_n N_VGND_c_920_n
+ PM_SKY130_FD_SC_HDLL__O31AI_4%VGND
cc_1 VNB N_A1_M1003_g 0.0248455f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_2 VNB N_A1_M1014_g 0.018541f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.56
cc_3 VNB N_A1_M1015_g 0.0190401f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.56
cc_4 VNB N_A1_M1026_g 0.0187919f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_5 VNB N_A1_c_108_n 0.0960913f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.217
cc_6 VNB A1 0.0144966f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.19
cc_7 VNB N_A2_M1008_g 0.0182928f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_8 VNB N_A2_M1011_g 0.018541f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.56
cc_9 VNB N_A2_M1021_g 0.0190401f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.56
cc_10 VNB N_A2_M1029_g 0.0187919f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_11 VNB A2 0.0058857f $X=-0.19 $Y=-0.24 $X2=1.68 $Y2=1.105
cc_12 VNB N_A2_c_197_n 0.0896153f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=1.217
cc_13 VNB N_A3_M1000_g 0.0245973f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_14 VNB N_A3_M1017_g 0.0239798f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.56
cc_15 VNB N_A3_M1023_g 0.020082f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.56
cc_16 VNB N_A3_M1027_g 0.0198226f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_17 VNB N_A3_c_288_n 0.0120068f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_18 VNB N_A3_c_289_n 0.030783f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_19 VNB N_A3_c_290_n 0.0899734f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.16
cc_20 VNB A3 0.00698319f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.24
cc_21 VNB N_B1_M1004_g 0.0177442f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_22 VNB N_B1_M1009_g 0.0184894f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.56
cc_23 VNB N_B1_M1012_g 0.0185367f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.56
cc_24 VNB N_B1_M1022_g 0.0249052f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.985
cc_25 VNB B1 0.0143034f $X=-0.19 $Y=-0.24 $X2=1.17 $Y2=1.105
cc_26 VNB N_B1_c_362_n 0.101665f $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=1.16
cc_27 VNB N_VPWR_c_510_n 0.364621f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.16
cc_28 VNB Y 0.00144061f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=1.217
cc_29 VNB N_A_31_47#_c_753_n 0.0188118f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_30 VNB N_A_31_47#_c_754_n 0.00983636f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_31_47#_c_755_n 0.001463f $X=-0.19 $Y=-0.24 $X2=0.745 $Y2=1.24
cc_32 VNB N_A_31_47#_c_756_n 0.0101084f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_31_47#_c_757_n 0.0186652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_31_47#_c_758_n 0.00146668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_31_47#_c_759_n 0.00356912f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_31_47#_c_760_n 0.00146668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_31_47#_c_761_n 0.00496288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_31_47#_c_762_n 0.00108591f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_903_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.985
cc_40 VNB N_VGND_c_904_n 0.0191455f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=1.025
cc_41 VNB N_VGND_c_905_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_42 VNB N_VGND_c_906_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_907_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.217
cc_44 VNB N_VGND_c_908_n 0.00530977f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_45 VNB N_VGND_c_909_n 0.0191455f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.16
cc_46 VNB N_VGND_c_910_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.16
cc_47 VNB N_VGND_c_911_n 0.0191455f $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=1.16
cc_48 VNB N_VGND_c_912_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=1.16
cc_49 VNB N_VGND_c_913_n 0.0165302f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.217
cc_50 VNB N_VGND_c_914_n 0.00708808f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.217
cc_51 VNB N_VGND_c_915_n 0.0623589f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_916_n 0.412442f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_917_n 0.0222518f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_918_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_919_n 0.0197062f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_920_n 0.01691f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VPB N_A1_c_110_n 0.0207821f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_58 VPB N_A1_c_111_n 0.0161549f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_59 VPB N_A1_c_112_n 0.0161549f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_60 VPB N_A1_c_113_n 0.0163866f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_61 VPB N_A1_c_108_n 0.0242435f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.217
cc_62 VPB A1 0.0166927f $X=-0.19 $Y=1.305 $X2=1.78 $Y2=1.19
cc_63 VPB N_A2_c_198_n 0.0163141f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_64 VPB N_A2_c_199_n 0.0161549f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_65 VPB N_A2_c_200_n 0.0161549f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_66 VPB N_A2_c_201_n 0.0198635f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_67 VPB A2 0.0179143f $X=-0.19 $Y=1.305 $X2=1.68 $Y2=1.105
cc_68 VPB N_A2_c_197_n 0.0236644f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=1.217
cc_69 VPB N_A3_c_292_n 0.0201091f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_70 VPB N_A3_c_293_n 0.0158911f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_71 VPB N_A3_c_294_n 0.0158911f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_72 VPB N_A3_c_295_n 0.015983f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_73 VPB N_A3_c_290_n 0.0286582f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.16
cc_74 VPB N_B1_c_363_n 0.0153951f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_75 VPB N_B1_c_364_n 0.0156918f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_76 VPB N_B1_c_365_n 0.0154218f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_77 VPB N_B1_c_366_n 0.0199377f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.56
cc_78 VPB N_B1_c_362_n 0.0282801f $X=-0.19 $Y=1.305 $X2=1.375 $Y2=1.16
cc_79 VPB N_A_27_297#_c_428_n 0.0131401f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=0.56
cc_80 VPB N_A_27_297#_c_429_n 0.0226427f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_27_297#_c_430_n 0.00471408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_511_n 0.00469739f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=0.56
cc_83 VPB N_VPWR_c_512_n 0.0206409f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_84 VPB N_VPWR_c_513_n 0.00469188f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.985
cc_85 VPB N_VPWR_c_514_n 4.04661e-19 $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.56
cc_86 VPB N_VPWR_c_515_n 4.04661e-19 $X=-0.19 $Y=1.305 $X2=1.17 $Y2=1.105
cc_87 VPB N_VPWR_c_516_n 0.116021f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_517_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_518_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.217
cc_90 VPB N_VPWR_c_519_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.217
cc_91 VPB N_VPWR_c_520_n 0.0190603f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.16
cc_92 VPB N_VPWR_c_510_n 0.0498316f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.16
cc_93 VPB N_VPWR_c_522_n 0.0230861f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.24
cc_94 VPB N_VPWR_c_523_n 0.00324032f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.24
cc_95 VPB N_A_497_297#_c_622_n 0.00738801f $X=-0.19 $Y=1.305 $X2=1.17 $Y2=1.105
cc_96 VPB Y 0.00182358f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.217
cc_97 VPB Y 0.00103485f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.217
cc_98 VPB Y 0.0326785f $X=-0.19 $Y=1.305 $X2=1.375 $Y2=1.217
cc_99 VPB N_Y_c_674_n 0.015166f $X=-0.19 $Y=1.305 $X2=0.745 $Y2=1.24
cc_100 VPB N_Y_c_675_n 0.00135271f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_Y_c_676_n 0.00378275f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_Y_c_677_n 0.00243899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_Y_c_678_n 0.0155574f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 N_A1_M1026_g N_A2_M1008_g 0.0162372f $X=1.95 $Y=0.56 $X2=0 $Y2=0
cc_105 N_A1_c_113_n N_A2_c_198_n 0.00992198f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_106 N_A1_c_108_n A2 0.00313533f $X=1.925 $Y=1.217 $X2=0 $Y2=0
cc_107 A1 A2 0.0269635f $X=1.78 $Y=1.19 $X2=0 $Y2=0
cc_108 N_A1_c_108_n N_A2_c_197_n 0.0162372f $X=1.925 $Y=1.217 $X2=0 $Y2=0
cc_109 A1 N_A2_c_197_n 3.07687e-19 $X=1.78 $Y=1.19 $X2=0 $Y2=0
cc_110 N_A1_c_110_n N_A_27_297#_c_428_n 8.12161e-19 $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_111 A1 N_A_27_297#_c_428_n 0.028375f $X=1.78 $Y=1.19 $X2=0 $Y2=0
cc_112 N_A1_c_110_n N_A_27_297#_c_429_n 0.00793864f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A1_c_111_n N_A_27_297#_c_429_n 6.16404e-19 $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A1_c_110_n N_A_27_297#_c_435_n 0.0144108f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A1_c_111_n N_A_27_297#_c_435_n 0.0110323f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A1_c_108_n N_A_27_297#_c_435_n 0.00125232f $X=1.925 $Y=1.217 $X2=0
+ $Y2=0
cc_117 A1 N_A_27_297#_c_435_n 0.0394639f $X=1.78 $Y=1.19 $X2=0 $Y2=0
cc_118 N_A1_c_110_n N_A_27_297#_c_439_n 6.53046e-19 $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A1_c_111_n N_A_27_297#_c_439_n 0.00985792f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A1_c_112_n N_A_27_297#_c_439_n 0.00793864f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A1_c_113_n N_A_27_297#_c_439_n 6.15975e-19 $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A1_c_112_n N_A_27_297#_c_443_n 0.0144108f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A1_c_113_n N_A_27_297#_c_443_n 0.0114971f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A1_c_108_n N_A_27_297#_c_443_n 0.00125645f $X=1.925 $Y=1.217 $X2=0
+ $Y2=0
cc_125 A1 N_A_27_297#_c_443_n 0.0383734f $X=1.78 $Y=1.19 $X2=0 $Y2=0
cc_126 N_A1_c_113_n N_A_27_297#_c_447_n 0.00553136f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A1_c_112_n N_A_27_297#_c_448_n 5.78464e-19 $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A1_c_113_n N_A_27_297#_c_448_n 0.00986416f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A1_c_111_n N_A_27_297#_c_450_n 0.00294943f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A1_c_112_n N_A_27_297#_c_450_n 8.12161e-19 $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A1_c_108_n N_A_27_297#_c_450_n 0.00132924f $X=1.925 $Y=1.217 $X2=0
+ $Y2=0
cc_132 A1 N_A_27_297#_c_450_n 0.0273952f $X=1.78 $Y=1.19 $X2=0 $Y2=0
cc_133 N_A1_c_110_n N_VPWR_c_511_n 0.00476657f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A1_c_111_n N_VPWR_c_511_n 0.00447692f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A1_c_111_n N_VPWR_c_512_n 0.00597712f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A1_c_112_n N_VPWR_c_512_n 0.00673617f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A1_c_112_n N_VPWR_c_513_n 0.00476657f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A1_c_113_n N_VPWR_c_513_n 0.00447307f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A1_c_113_n N_VPWR_c_516_n 0.00596194f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A1_c_110_n N_VPWR_c_510_n 0.0079958f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A1_c_111_n N_VPWR_c_510_n 0.0067049f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A1_c_112_n N_VPWR_c_510_n 0.00706625f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A1_c_113_n N_VPWR_c_510_n 0.00673919f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A1_c_110_n N_VPWR_c_522_n 0.00673617f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A1_M1003_g N_A_31_47#_c_753_n 0.00674948f $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_146 N_A1_M1014_g N_A_31_47#_c_753_n 5.42611e-19 $X=0.96 $Y=0.56 $X2=0 $Y2=0
cc_147 N_A1_M1003_g N_A_31_47#_c_765_n 0.0087374f $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_148 N_A1_M1014_g N_A_31_47#_c_765_n 0.0087374f $X=0.96 $Y=0.56 $X2=0 $Y2=0
cc_149 N_A1_c_108_n N_A_31_47#_c_765_n 0.00312059f $X=1.925 $Y=1.217 $X2=0 $Y2=0
cc_150 A1 N_A_31_47#_c_765_n 0.0369305f $X=1.78 $Y=1.19 $X2=0 $Y2=0
cc_151 N_A1_M1003_g N_A_31_47#_c_754_n 8.68782e-19 $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_152 A1 N_A_31_47#_c_754_n 0.0281907f $X=1.78 $Y=1.19 $X2=0 $Y2=0
cc_153 N_A1_M1003_g N_A_31_47#_c_771_n 5.22028e-19 $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_154 N_A1_M1014_g N_A_31_47#_c_771_n 0.00641183f $X=0.96 $Y=0.56 $X2=0 $Y2=0
cc_155 N_A1_M1015_g N_A_31_47#_c_771_n 0.00681792f $X=1.43 $Y=0.56 $X2=0 $Y2=0
cc_156 N_A1_M1026_g N_A_31_47#_c_771_n 5.31317e-19 $X=1.95 $Y=0.56 $X2=0 $Y2=0
cc_157 N_A1_M1015_g N_A_31_47#_c_775_n 0.00899636f $X=1.43 $Y=0.56 $X2=0 $Y2=0
cc_158 N_A1_M1026_g N_A_31_47#_c_775_n 0.00669407f $X=1.95 $Y=0.56 $X2=0 $Y2=0
cc_159 N_A1_c_108_n N_A_31_47#_c_775_n 0.00423509f $X=1.925 $Y=1.217 $X2=0 $Y2=0
cc_160 A1 N_A_31_47#_c_775_n 0.0360045f $X=1.78 $Y=1.19 $X2=0 $Y2=0
cc_161 N_A1_M1015_g N_A_31_47#_c_779_n 5.66697e-19 $X=1.43 $Y=0.56 $X2=0 $Y2=0
cc_162 N_A1_M1026_g N_A_31_47#_c_779_n 0.00843196f $X=1.95 $Y=0.56 $X2=0 $Y2=0
cc_163 N_A1_M1014_g N_A_31_47#_c_758_n 8.68782e-19 $X=0.96 $Y=0.56 $X2=0 $Y2=0
cc_164 N_A1_M1015_g N_A_31_47#_c_758_n 8.68782e-19 $X=1.43 $Y=0.56 $X2=0 $Y2=0
cc_165 N_A1_c_108_n N_A_31_47#_c_758_n 0.00323693f $X=1.925 $Y=1.217 $X2=0 $Y2=0
cc_166 A1 N_A_31_47#_c_758_n 0.0261364f $X=1.78 $Y=1.19 $X2=0 $Y2=0
cc_167 N_A1_M1026_g N_A_31_47#_c_759_n 0.00525283f $X=1.95 $Y=0.56 $X2=0 $Y2=0
cc_168 N_A1_M1003_g N_VGND_c_903_n 0.00376026f $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_169 N_A1_M1014_g N_VGND_c_903_n 0.00276126f $X=0.96 $Y=0.56 $X2=0 $Y2=0
cc_170 N_A1_M1014_g N_VGND_c_904_n 0.00422241f $X=0.96 $Y=0.56 $X2=0 $Y2=0
cc_171 N_A1_M1015_g N_VGND_c_904_n 0.00422241f $X=1.43 $Y=0.56 $X2=0 $Y2=0
cc_172 N_A1_M1015_g N_VGND_c_905_n 0.00382269f $X=1.43 $Y=0.56 $X2=0 $Y2=0
cc_173 N_A1_M1026_g N_VGND_c_905_n 0.00362873f $X=1.95 $Y=0.56 $X2=0 $Y2=0
cc_174 N_A1_M1026_g N_VGND_c_909_n 0.00395968f $X=1.95 $Y=0.56 $X2=0 $Y2=0
cc_175 N_A1_M1003_g N_VGND_c_916_n 0.00691918f $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_176 N_A1_M1014_g N_VGND_c_916_n 0.0059505f $X=0.96 $Y=0.56 $X2=0 $Y2=0
cc_177 N_A1_M1015_g N_VGND_c_916_n 0.00618861f $X=1.43 $Y=0.56 $X2=0 $Y2=0
cc_178 N_A1_M1026_g N_VGND_c_916_n 0.00581897f $X=1.95 $Y=0.56 $X2=0 $Y2=0
cc_179 N_A1_M1003_g N_VGND_c_917_n 0.00422241f $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_180 N_A2_M1029_g N_A3_M1000_g 0.0137836f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_181 A2 N_A3_c_288_n 0.00146591f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_182 N_A2_c_197_n N_A3_c_288_n 0.0137836f $X=3.805 $Y=1.217 $X2=0 $Y2=0
cc_183 A2 A3 0.0194357f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_184 N_A2_c_197_n A3 2.27279e-19 $X=3.805 $Y=1.217 $X2=0 $Y2=0
cc_185 N_A2_c_198_n N_A_27_297#_c_447_n 0.00378365f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_186 A2 N_A_27_297#_c_447_n 0.0125596f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_187 N_A2_c_198_n N_A_27_297#_c_448_n 0.00536381f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A2_c_199_n N_A_27_297#_c_448_n 5.32902e-19 $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A2_c_198_n N_A_27_297#_c_458_n 0.015794f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_190 N_A2_c_199_n N_A_27_297#_c_458_n 0.0101559f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_191 N_A2_c_200_n N_A_27_297#_c_430_n 0.0129706f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_192 N_A2_c_201_n N_A_27_297#_c_430_n 0.0115612f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A2_c_198_n N_A_27_297#_c_462_n 6.95719e-19 $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A2_c_199_n N_A_27_297#_c_462_n 0.00910731f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A2_c_200_n N_A_27_297#_c_462_n 0.00604378f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A2_c_201_n N_A_27_297#_c_462_n 9.68813e-19 $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A2_c_198_n N_VPWR_c_516_n 0.00429425f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A2_c_199_n N_VPWR_c_516_n 0.00430873f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A2_c_200_n N_VPWR_c_516_n 0.00430943f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_200 N_A2_c_201_n N_VPWR_c_516_n 0.00429453f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A2_c_198_n N_VPWR_c_510_n 0.00609019f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A2_c_199_n N_VPWR_c_510_n 0.00605584f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A2_c_200_n N_VPWR_c_510_n 0.0060559f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A2_c_201_n N_VPWR_c_510_n 0.00734734f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A2_c_201_n N_A_497_297#_c_623_n 0.00397427f $X=3.805 $Y=1.41 $X2=0
+ $Y2=0
cc_206 N_A2_c_198_n N_A_497_297#_c_624_n 0.00188234f $X=2.395 $Y=1.41 $X2=0
+ $Y2=0
cc_207 N_A2_c_199_n N_A_497_297#_c_624_n 0.00397606f $X=2.865 $Y=1.41 $X2=0
+ $Y2=0
cc_208 A2 N_A_497_297#_c_624_n 0.0142151f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_209 N_A2_c_197_n N_A_497_297#_c_624_n 9.26878e-19 $X=3.805 $Y=1.217 $X2=0
+ $Y2=0
cc_210 N_A2_c_199_n N_A_497_297#_c_628_n 0.0108069f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A2_c_200_n N_A_497_297#_c_628_n 0.0112356f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_212 A2 N_A_497_297#_c_628_n 0.0875041f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_213 N_A2_c_197_n N_A_497_297#_c_628_n 0.00138184f $X=3.805 $Y=1.217 $X2=0
+ $Y2=0
cc_214 N_A2_c_200_n N_A_497_297#_c_632_n 0.00527455f $X=3.335 $Y=1.41 $X2=0
+ $Y2=0
cc_215 N_A2_c_201_n N_A_497_297#_c_632_n 0.0217568f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A2_c_197_n N_A_497_297#_c_632_n 0.00128152f $X=3.805 $Y=1.217 $X2=0
+ $Y2=0
cc_217 N_A2_c_201_n N_Y_c_674_n 0.00617178f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A2_M1008_g N_A_31_47#_c_779_n 0.00674948f $X=2.37 $Y=0.56 $X2=0 $Y2=0
cc_219 N_A2_M1011_g N_A_31_47#_c_779_n 5.42233e-19 $X=2.84 $Y=0.56 $X2=0 $Y2=0
cc_220 N_A2_M1008_g N_A_31_47#_c_788_n 0.0087374f $X=2.37 $Y=0.56 $X2=0 $Y2=0
cc_221 N_A2_M1011_g N_A_31_47#_c_788_n 0.0087374f $X=2.84 $Y=0.56 $X2=0 $Y2=0
cc_222 A2 N_A_31_47#_c_788_n 0.0369305f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_223 N_A2_c_197_n N_A_31_47#_c_788_n 0.00312059f $X=3.805 $Y=1.217 $X2=0 $Y2=0
cc_224 N_A2_M1008_g N_A_31_47#_c_792_n 5.22028e-19 $X=2.37 $Y=0.56 $X2=0 $Y2=0
cc_225 N_A2_M1011_g N_A_31_47#_c_792_n 0.00641183f $X=2.84 $Y=0.56 $X2=0 $Y2=0
cc_226 N_A2_M1021_g N_A_31_47#_c_792_n 0.00681792f $X=3.31 $Y=0.56 $X2=0 $Y2=0
cc_227 N_A2_M1029_g N_A_31_47#_c_792_n 5.31317e-19 $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_228 N_A2_M1021_g N_A_31_47#_c_796_n 0.00899636f $X=3.31 $Y=0.56 $X2=0 $Y2=0
cc_229 N_A2_M1029_g N_A_31_47#_c_796_n 0.00626649f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_230 A2 N_A_31_47#_c_796_n 0.0370518f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_231 N_A2_c_197_n N_A_31_47#_c_796_n 0.00423509f $X=3.805 $Y=1.217 $X2=0 $Y2=0
cc_232 N_A2_M1021_g N_A_31_47#_c_800_n 5.66697e-19 $X=3.31 $Y=0.56 $X2=0 $Y2=0
cc_233 N_A2_M1029_g N_A_31_47#_c_800_n 0.00843196f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_234 N_A2_M1008_g N_A_31_47#_c_759_n 8.68782e-19 $X=2.37 $Y=0.56 $X2=0 $Y2=0
cc_235 A2 N_A_31_47#_c_759_n 0.0124322f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_236 N_A2_M1011_g N_A_31_47#_c_760_n 8.68782e-19 $X=2.84 $Y=0.56 $X2=0 $Y2=0
cc_237 N_A2_M1021_g N_A_31_47#_c_760_n 8.68782e-19 $X=3.31 $Y=0.56 $X2=0 $Y2=0
cc_238 A2 N_A_31_47#_c_760_n 0.0261364f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_239 N_A2_c_197_n N_A_31_47#_c_760_n 0.00323693f $X=3.805 $Y=1.217 $X2=0 $Y2=0
cc_240 N_A2_M1029_g N_A_31_47#_c_761_n 0.00239159f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_241 A2 N_A_31_47#_c_761_n 0.0125212f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_242 N_A2_M1008_g N_VGND_c_906_n 0.00376026f $X=2.37 $Y=0.56 $X2=0 $Y2=0
cc_243 N_A2_M1011_g N_VGND_c_906_n 0.00276126f $X=2.84 $Y=0.56 $X2=0 $Y2=0
cc_244 N_A2_M1021_g N_VGND_c_907_n 0.00382269f $X=3.31 $Y=0.56 $X2=0 $Y2=0
cc_245 N_A2_M1029_g N_VGND_c_907_n 0.00362873f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_246 N_A2_M1008_g N_VGND_c_909_n 0.00422241f $X=2.37 $Y=0.56 $X2=0 $Y2=0
cc_247 N_A2_M1011_g N_VGND_c_911_n 0.00422241f $X=2.84 $Y=0.56 $X2=0 $Y2=0
cc_248 N_A2_M1021_g N_VGND_c_911_n 0.00422241f $X=3.31 $Y=0.56 $X2=0 $Y2=0
cc_249 N_A2_M1008_g N_VGND_c_916_n 0.0059735f $X=2.37 $Y=0.56 $X2=0 $Y2=0
cc_250 N_A2_M1011_g N_VGND_c_916_n 0.0059505f $X=2.84 $Y=0.56 $X2=0 $Y2=0
cc_251 N_A2_M1021_g N_VGND_c_916_n 0.00618861f $X=3.31 $Y=0.56 $X2=0 $Y2=0
cc_252 N_A2_M1029_g N_VGND_c_916_n 0.00581897f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_253 N_A2_M1029_g N_VGND_c_919_n 0.00395968f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_254 N_A3_M1027_g N_B1_M1004_g 0.0217701f $X=6.295 $Y=0.56 $X2=0 $Y2=0
cc_255 N_A3_c_295_n N_B1_c_363_n 0.00959456f $X=6.27 $Y=1.41 $X2=0 $Y2=0
cc_256 N_A3_c_290_n N_B1_c_362_n 0.0217701f $X=6.27 $Y=1.217 $X2=0 $Y2=0
cc_257 A3 N_B1_c_362_n 0.00213713f $X=6.355 $Y=1.19 $X2=0 $Y2=0
cc_258 N_A3_c_292_n N_A_27_297#_c_430_n 0.00122868f $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A3_c_295_n N_VPWR_c_514_n 0.00127095f $X=6.27 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A3_c_292_n N_VPWR_c_516_n 0.00429453f $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A3_c_293_n N_VPWR_c_516_n 0.00429453f $X=5.33 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A3_c_294_n N_VPWR_c_516_n 0.00429453f $X=5.8 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A3_c_295_n N_VPWR_c_516_n 0.00672127f $X=6.27 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A3_c_292_n N_VPWR_c_510_n 0.00739666f $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A3_c_293_n N_VPWR_c_510_n 0.00606499f $X=5.33 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A3_c_294_n N_VPWR_c_510_n 0.00606499f $X=5.8 $Y=1.41 $X2=0 $Y2=0
cc_267 N_A3_c_295_n N_VPWR_c_510_n 0.0119297f $X=6.27 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A3_c_292_n N_A_497_297#_c_623_n 0.0265067f $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A3_c_293_n N_A_497_297#_c_636_n 0.0215684f $X=5.33 $Y=1.41 $X2=0 $Y2=0
cc_270 N_A3_c_294_n N_A_497_297#_c_636_n 0.0215684f $X=5.8 $Y=1.41 $X2=0 $Y2=0
cc_271 N_A3_c_295_n N_A_497_297#_c_636_n 0.00745123f $X=6.27 $Y=1.41 $X2=0 $Y2=0
cc_272 N_A3_M1027_g Y 8.70259e-19 $X=6.295 $Y=0.56 $X2=0 $Y2=0
cc_273 N_A3_c_290_n Y 8.72022e-19 $X=6.27 $Y=1.217 $X2=0 $Y2=0
cc_274 A3 Y 0.0179651f $X=6.355 $Y=1.19 $X2=0 $Y2=0
cc_275 N_A3_c_292_n N_Y_c_674_n 0.0131161f $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_276 N_A3_c_293_n N_Y_c_674_n 0.0127007f $X=5.33 $Y=1.41 $X2=0 $Y2=0
cc_277 N_A3_c_294_n N_Y_c_674_n 0.0127007f $X=5.8 $Y=1.41 $X2=0 $Y2=0
cc_278 N_A3_c_295_n N_Y_c_674_n 0.0178311f $X=6.27 $Y=1.41 $X2=0 $Y2=0
cc_279 N_A3_c_288_n N_Y_c_674_n 0.0141543f $X=4.325 $Y=1.16 $X2=0 $Y2=0
cc_280 N_A3_c_290_n N_Y_c_674_n 0.022637f $X=6.27 $Y=1.217 $X2=0 $Y2=0
cc_281 A3 N_Y_c_674_n 0.179429f $X=6.355 $Y=1.19 $X2=0 $Y2=0
cc_282 N_A3_M1000_g N_A_31_47#_c_800_n 0.0114904f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_283 N_A3_M1000_g N_A_31_47#_c_811_n 0.0105442f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_284 N_A3_M1017_g N_A_31_47#_c_811_n 0.0135834f $X=5.185 $Y=0.56 $X2=0 $Y2=0
cc_285 N_A3_c_289_n N_A_31_47#_c_811_n 0.0144f $X=4.76 $Y=1.16 $X2=0 $Y2=0
cc_286 N_A3_c_290_n N_A_31_47#_c_811_n 2.70619e-19 $X=6.27 $Y=1.217 $X2=0 $Y2=0
cc_287 A3 N_A_31_47#_c_811_n 0.0756647f $X=6.355 $Y=1.19 $X2=0 $Y2=0
cc_288 N_A3_M1023_g N_A_31_47#_c_755_n 0.0128768f $X=5.655 $Y=0.56 $X2=0 $Y2=0
cc_289 N_A3_M1027_g N_A_31_47#_c_755_n 0.0122836f $X=6.295 $Y=0.56 $X2=0 $Y2=0
cc_290 N_A3_c_290_n N_A_31_47#_c_755_n 0.00727706f $X=6.27 $Y=1.217 $X2=0 $Y2=0
cc_291 A3 N_A_31_47#_c_755_n 0.0690051f $X=6.355 $Y=1.19 $X2=0 $Y2=0
cc_292 N_A3_M1000_g N_A_31_47#_c_761_n 8.68782e-19 $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_293 A3 N_A_31_47#_c_761_n 0.00227082f $X=6.355 $Y=1.19 $X2=0 $Y2=0
cc_294 N_A3_c_290_n N_A_31_47#_c_762_n 0.00330072f $X=6.27 $Y=1.217 $X2=0 $Y2=0
cc_295 A3 N_A_31_47#_c_762_n 0.0129933f $X=6.355 $Y=1.19 $X2=0 $Y2=0
cc_296 N_A3_M1023_g N_VGND_c_908_n 0.00619024f $X=5.655 $Y=0.56 $X2=0 $Y2=0
cc_297 N_A3_M1027_g N_VGND_c_908_n 0.00701756f $X=6.295 $Y=0.56 $X2=0 $Y2=0
cc_298 N_A3_M1017_g N_VGND_c_913_n 0.00348405f $X=5.185 $Y=0.56 $X2=0 $Y2=0
cc_299 N_A3_M1023_g N_VGND_c_913_n 0.00436487f $X=5.655 $Y=0.56 $X2=0 $Y2=0
cc_300 N_A3_M1027_g N_VGND_c_915_n 0.00436487f $X=6.295 $Y=0.56 $X2=0 $Y2=0
cc_301 N_A3_M1000_g N_VGND_c_916_n 0.00726788f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_302 N_A3_M1017_g N_VGND_c_916_n 0.00426048f $X=5.185 $Y=0.56 $X2=0 $Y2=0
cc_303 N_A3_M1023_g N_VGND_c_916_n 0.00660368f $X=5.655 $Y=0.56 $X2=0 $Y2=0
cc_304 N_A3_M1027_g N_VGND_c_916_n 0.00650008f $X=6.295 $Y=0.56 $X2=0 $Y2=0
cc_305 N_A3_M1000_g N_VGND_c_919_n 0.00422241f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_306 N_A3_M1000_g N_VGND_c_920_n 0.0115201f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_307 N_A3_M1017_g N_VGND_c_920_n 0.0109061f $X=5.185 $Y=0.56 $X2=0 $Y2=0
cc_308 N_A3_M1023_g N_VGND_c_920_n 9.52286e-19 $X=5.655 $Y=0.56 $X2=0 $Y2=0
cc_309 N_B1_c_363_n N_VPWR_c_514_n 0.01571f $X=6.74 $Y=1.41 $X2=0 $Y2=0
cc_310 N_B1_c_364_n N_VPWR_c_514_n 0.0110779f $X=7.21 $Y=1.41 $X2=0 $Y2=0
cc_311 N_B1_c_365_n N_VPWR_c_514_n 6.04384e-19 $X=7.68 $Y=1.41 $X2=0 $Y2=0
cc_312 N_B1_c_364_n N_VPWR_c_515_n 6.40835e-19 $X=7.21 $Y=1.41 $X2=0 $Y2=0
cc_313 N_B1_c_365_n N_VPWR_c_515_n 0.014614f $X=7.68 $Y=1.41 $X2=0 $Y2=0
cc_314 N_B1_c_366_n N_VPWR_c_515_n 0.0128922f $X=8.15 $Y=1.41 $X2=0 $Y2=0
cc_315 N_B1_c_363_n N_VPWR_c_516_n 0.00427505f $X=6.74 $Y=1.41 $X2=0 $Y2=0
cc_316 N_B1_c_364_n N_VPWR_c_518_n 0.00622633f $X=7.21 $Y=1.41 $X2=0 $Y2=0
cc_317 N_B1_c_365_n N_VPWR_c_518_n 0.00427505f $X=7.68 $Y=1.41 $X2=0 $Y2=0
cc_318 N_B1_c_366_n N_VPWR_c_520_n 0.00622633f $X=8.15 $Y=1.41 $X2=0 $Y2=0
cc_319 N_B1_c_363_n N_VPWR_c_510_n 0.00735499f $X=6.74 $Y=1.41 $X2=0 $Y2=0
cc_320 N_B1_c_364_n N_VPWR_c_510_n 0.0104011f $X=7.21 $Y=1.41 $X2=0 $Y2=0
cc_321 N_B1_c_365_n N_VPWR_c_510_n 0.00732977f $X=7.68 $Y=1.41 $X2=0 $Y2=0
cc_322 N_B1_c_366_n N_VPWR_c_510_n 0.0115056f $X=8.15 $Y=1.41 $X2=0 $Y2=0
cc_323 N_B1_M1009_g N_Y_c_690_n 0.0112521f $X=7.185 $Y=0.56 $X2=0 $Y2=0
cc_324 N_B1_M1012_g N_Y_c_690_n 0.0106317f $X=7.655 $Y=0.56 $X2=0 $Y2=0
cc_325 N_B1_M1022_g N_Y_c_690_n 0.0037383f $X=8.125 $Y=0.56 $X2=0 $Y2=0
cc_326 B1 N_Y_c_690_n 0.0577744f $X=8.355 $Y=1.105 $X2=0 $Y2=0
cc_327 N_B1_c_362_n N_Y_c_690_n 0.00696439f $X=8.125 $Y=1.217 $X2=0 $Y2=0
cc_328 N_B1_M1004_g N_Y_c_695_n 0.00291048f $X=6.715 $Y=0.56 $X2=0 $Y2=0
cc_329 N_B1_M1004_g Y 0.00379829f $X=6.715 $Y=0.56 $X2=0 $Y2=0
cc_330 N_B1_c_363_n Y 0.00123141f $X=6.74 $Y=1.41 $X2=0 $Y2=0
cc_331 N_B1_M1009_g Y 0.00333472f $X=7.185 $Y=0.56 $X2=0 $Y2=0
cc_332 N_B1_c_364_n Y 8.20075e-19 $X=7.21 $Y=1.41 $X2=0 $Y2=0
cc_333 B1 Y 0.016985f $X=8.355 $Y=1.105 $X2=0 $Y2=0
cc_334 N_B1_c_362_n Y 0.0252277f $X=8.125 $Y=1.217 $X2=0 $Y2=0
cc_335 B1 Y 0.0139499f $X=8.355 $Y=1.105 $X2=0 $Y2=0
cc_336 N_B1_c_362_n Y 0.00409765f $X=8.125 $Y=1.217 $X2=0 $Y2=0
cc_337 N_B1_c_366_n Y 0.0114869f $X=8.15 $Y=1.41 $X2=0 $Y2=0
cc_338 N_B1_c_364_n N_Y_c_675_n 0.0184197f $X=7.21 $Y=1.41 $X2=0 $Y2=0
cc_339 B1 N_Y_c_675_n 0.0140845f $X=8.355 $Y=1.105 $X2=0 $Y2=0
cc_340 N_B1_c_362_n N_Y_c_675_n 0.00552408f $X=8.125 $Y=1.217 $X2=0 $Y2=0
cc_341 N_B1_c_363_n N_Y_c_676_n 0.0191608f $X=6.74 $Y=1.41 $X2=0 $Y2=0
cc_342 N_B1_c_362_n N_Y_c_676_n 0.00141271f $X=8.125 $Y=1.217 $X2=0 $Y2=0
cc_343 N_B1_c_365_n N_Y_c_677_n 0.0163251f $X=7.68 $Y=1.41 $X2=0 $Y2=0
cc_344 N_B1_c_366_n N_Y_c_677_n 0.0184695f $X=8.15 $Y=1.41 $X2=0 $Y2=0
cc_345 B1 N_Y_c_677_n 0.0563757f $X=8.355 $Y=1.105 $X2=0 $Y2=0
cc_346 N_B1_c_362_n N_Y_c_677_n 0.0103248f $X=8.125 $Y=1.217 $X2=0 $Y2=0
cc_347 B1 N_Y_c_678_n 0.0244039f $X=8.355 $Y=1.105 $X2=0 $Y2=0
cc_348 N_B1_c_362_n N_Y_c_678_n 5.73441e-19 $X=8.125 $Y=1.217 $X2=0 $Y2=0
cc_349 N_B1_M1004_g N_A_31_47#_c_824_n 0.014057f $X=6.715 $Y=0.56 $X2=0 $Y2=0
cc_350 N_B1_M1009_g N_A_31_47#_c_824_n 0.00923997f $X=7.185 $Y=0.56 $X2=0 $Y2=0
cc_351 N_B1_M1012_g N_A_31_47#_c_824_n 0.00931157f $X=7.655 $Y=0.56 $X2=0 $Y2=0
cc_352 N_B1_M1022_g N_A_31_47#_c_824_n 0.0108933f $X=8.125 $Y=0.56 $X2=0 $Y2=0
cc_353 B1 N_A_31_47#_c_824_n 0.00497946f $X=8.355 $Y=1.105 $X2=0 $Y2=0
cc_354 N_B1_c_362_n N_A_31_47#_c_824_n 0.00200338f $X=8.125 $Y=1.217 $X2=0 $Y2=0
cc_355 B1 N_A_31_47#_c_757_n 0.0237212f $X=8.355 $Y=1.105 $X2=0 $Y2=0
cc_356 N_B1_c_362_n N_A_31_47#_c_757_n 5.54902e-19 $X=8.125 $Y=1.217 $X2=0 $Y2=0
cc_357 N_B1_M1004_g N_VGND_c_915_n 0.00357877f $X=6.715 $Y=0.56 $X2=0 $Y2=0
cc_358 N_B1_M1009_g N_VGND_c_915_n 0.00357877f $X=7.185 $Y=0.56 $X2=0 $Y2=0
cc_359 N_B1_M1012_g N_VGND_c_915_n 0.00357877f $X=7.655 $Y=0.56 $X2=0 $Y2=0
cc_360 N_B1_M1022_g N_VGND_c_915_n 0.00357877f $X=8.125 $Y=0.56 $X2=0 $Y2=0
cc_361 N_B1_M1004_g N_VGND_c_916_n 0.00542415f $X=6.715 $Y=0.56 $X2=0 $Y2=0
cc_362 N_B1_M1009_g N_VGND_c_916_n 0.00548399f $X=7.185 $Y=0.56 $X2=0 $Y2=0
cc_363 N_B1_M1012_g N_VGND_c_916_n 0.00548399f $X=7.655 $Y=0.56 $X2=0 $Y2=0
cc_364 N_B1_M1022_g N_VGND_c_916_n 0.00642416f $X=8.125 $Y=0.56 $X2=0 $Y2=0
cc_365 N_A_27_297#_c_435_n N_VPWR_M1002_d 0.00336681f $X=1.005 $Y=1.745
+ $X2=-0.19 $Y2=1.305
cc_366 N_A_27_297#_c_443_n N_VPWR_M1013_d 0.00336681f $X=1.945 $Y=1.745 $X2=0
+ $Y2=0
cc_367 N_A_27_297#_c_429_n N_VPWR_c_511_n 0.0243541f $X=0.28 $Y=2.36 $X2=0 $Y2=0
cc_368 N_A_27_297#_c_435_n N_VPWR_c_511_n 0.0138732f $X=1.005 $Y=1.745 $X2=0
+ $Y2=0
cc_369 N_A_27_297#_c_439_n N_VPWR_c_511_n 0.029862f $X=1.22 $Y=2.36 $X2=0 $Y2=0
cc_370 N_A_27_297#_c_439_n N_VPWR_c_512_n 0.0223557f $X=1.22 $Y=2.36 $X2=0 $Y2=0
cc_371 N_A_27_297#_c_439_n N_VPWR_c_513_n 0.0244833f $X=1.22 $Y=2.36 $X2=0 $Y2=0
cc_372 N_A_27_297#_c_443_n N_VPWR_c_513_n 0.0138732f $X=1.945 $Y=1.745 $X2=0
+ $Y2=0
cc_373 N_A_27_297#_c_448_n N_VPWR_c_513_n 0.0308489f $X=2.135 $Y=2.205 $X2=0
+ $Y2=0
cc_374 N_A_27_297#_c_448_n N_VPWR_c_516_n 0.0224921f $X=2.135 $Y=2.205 $X2=0
+ $Y2=0
cc_375 N_A_27_297#_c_458_n N_VPWR_c_516_n 0.032562f $X=2.885 $Y=2.335 $X2=0
+ $Y2=0
cc_376 N_A_27_297#_c_430_n N_VPWR_c_516_n 0.0608402f $X=4.04 $Y=2.36 $X2=0 $Y2=0
cc_377 N_A_27_297#_c_462_n N_VPWR_c_516_n 0.0220286f $X=3.1 $Y=2.02 $X2=0 $Y2=0
cc_378 N_A_27_297#_M1002_s N_VPWR_c_510_n 0.00233913f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_379 N_A_27_297#_M1006_s N_VPWR_c_510_n 0.00231261f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_380 N_A_27_297#_M1020_s N_VPWR_c_510_n 0.00231261f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_381 N_A_27_297#_M1016_s N_VPWR_c_510_n 0.00231261f $X=2.955 $Y=1.485 $X2=0
+ $Y2=0
cc_382 N_A_27_297#_M1031_s N_VPWR_c_510_n 0.00233941f $X=3.895 $Y=1.485 $X2=0
+ $Y2=0
cc_383 N_A_27_297#_c_429_n N_VPWR_c_510_n 0.0134353f $X=0.28 $Y=2.36 $X2=0 $Y2=0
cc_384 N_A_27_297#_c_435_n N_VPWR_c_510_n 0.0128394f $X=1.005 $Y=1.745 $X2=0
+ $Y2=0
cc_385 N_A_27_297#_c_439_n N_VPWR_c_510_n 0.0140101f $X=1.22 $Y=2.36 $X2=0 $Y2=0
cc_386 N_A_27_297#_c_443_n N_VPWR_c_510_n 0.0128394f $X=1.945 $Y=1.745 $X2=0
+ $Y2=0
cc_387 N_A_27_297#_c_448_n N_VPWR_c_510_n 0.014078f $X=2.135 $Y=2.205 $X2=0
+ $Y2=0
cc_388 N_A_27_297#_c_458_n N_VPWR_c_510_n 0.0198173f $X=2.885 $Y=2.335 $X2=0
+ $Y2=0
cc_389 N_A_27_297#_c_430_n N_VPWR_c_510_n 0.0367241f $X=4.04 $Y=2.36 $X2=0 $Y2=0
cc_390 N_A_27_297#_c_462_n N_VPWR_c_510_n 0.0139179f $X=3.1 $Y=2.02 $X2=0 $Y2=0
cc_391 N_A_27_297#_c_429_n N_VPWR_c_522_n 0.0228244f $X=0.28 $Y=2.36 $X2=0 $Y2=0
cc_392 N_A_27_297#_c_458_n N_A_497_297#_M1001_d 0.0034842f $X=2.885 $Y=2.335
+ $X2=-0.19 $Y2=1.305
cc_393 N_A_27_297#_c_430_n N_A_497_297#_M1024_d 0.0035426f $X=4.04 $Y=2.36 $X2=0
+ $Y2=0
cc_394 N_A_27_297#_c_430_n N_A_497_297#_c_623_n 0.0182013f $X=4.04 $Y=2.36 $X2=0
+ $Y2=0
cc_395 N_A_27_297#_c_447_n N_A_497_297#_c_624_n 0.0193048f $X=2.135 $Y=1.895
+ $X2=0 $Y2=0
cc_396 N_A_27_297#_c_448_n N_A_497_297#_c_624_n 0.00853797f $X=2.135 $Y=2.205
+ $X2=0 $Y2=0
cc_397 N_A_27_297#_c_458_n N_A_497_297#_c_624_n 0.0129977f $X=2.885 $Y=2.335
+ $X2=0 $Y2=0
cc_398 N_A_27_297#_c_462_n N_A_497_297#_c_624_n 0.00746551f $X=3.1 $Y=2.02 $X2=0
+ $Y2=0
cc_399 N_A_27_297#_M1016_s N_A_497_297#_c_628_n 0.00341904f $X=2.955 $Y=1.485
+ $X2=0 $Y2=0
cc_400 N_A_27_297#_c_458_n N_A_497_297#_c_628_n 0.00366604f $X=2.885 $Y=2.335
+ $X2=0 $Y2=0
cc_401 N_A_27_297#_c_430_n N_A_497_297#_c_628_n 0.0052348f $X=4.04 $Y=2.36 $X2=0
+ $Y2=0
cc_402 N_A_27_297#_c_462_n N_A_497_297#_c_628_n 0.0205168f $X=3.1 $Y=2.02 $X2=0
+ $Y2=0
cc_403 N_A_27_297#_M1031_s N_A_497_297#_c_632_n 0.00980149f $X=3.895 $Y=1.485
+ $X2=0 $Y2=0
cc_404 N_A_27_297#_c_430_n N_A_497_297#_c_632_n 0.0506846f $X=4.04 $Y=2.36 $X2=0
+ $Y2=0
cc_405 N_A_27_297#_c_462_n N_A_497_297#_c_632_n 0.00676772f $X=3.1 $Y=2.02 $X2=0
+ $Y2=0
cc_406 N_A_27_297#_M1031_s N_A_497_297#_c_622_n 0.00941839f $X=3.895 $Y=1.485
+ $X2=0 $Y2=0
cc_407 N_A_27_297#_M1031_s N_Y_c_674_n 0.00276848f $X=3.895 $Y=1.485 $X2=0 $Y2=0
cc_408 N_VPWR_c_510_n N_A_497_297#_M1001_d 0.00232895f $X=8.51 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_409 N_VPWR_c_510_n N_A_497_297#_M1024_d 0.00232895f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_510_n N_A_497_297#_M1005_s 0.00231289f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_510_n N_A_497_297#_M1018_s 0.00231289f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_516_n N_A_497_297#_c_623_n 0.100707f $X=6.76 $Y=2.72 $X2=0 $Y2=0
cc_413 N_VPWR_c_510_n N_A_497_297#_c_623_n 0.0612129f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_510_n N_A_497_297#_c_632_n 0.00822431f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_415 N_VPWR_c_516_n N_A_497_297#_c_622_n 0.00398962f $X=6.76 $Y=2.72 $X2=0
+ $Y2=0
cc_416 N_VPWR_c_510_n N_Y_M1005_d 0.00262917f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_417 N_VPWR_c_510_n N_Y_M1007_d 0.00232895f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_418 N_VPWR_c_510_n N_Y_M1028_d 0.00647849f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_419 N_VPWR_c_510_n N_Y_M1019_d 0.00647849f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_420 N_VPWR_c_510_n N_Y_M1030_d 0.00430086f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_421 N_VPWR_c_514_n N_Y_c_722_n 0.0429267f $X=6.975 $Y=2.02 $X2=0 $Y2=0
cc_422 N_VPWR_c_516_n N_Y_c_722_n 0.0118139f $X=6.76 $Y=2.72 $X2=0 $Y2=0
cc_423 N_VPWR_c_510_n N_Y_c_722_n 0.00646998f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_424 N_VPWR_c_514_n N_Y_c_725_n 0.0351948f $X=6.975 $Y=2.02 $X2=0 $Y2=0
cc_425 N_VPWR_c_515_n N_Y_c_725_n 0.0429267f $X=7.915 $Y=2.02 $X2=0 $Y2=0
cc_426 N_VPWR_c_518_n N_Y_c_725_n 0.0118139f $X=7.7 $Y=2.72 $X2=0 $Y2=0
cc_427 N_VPWR_c_510_n N_Y_c_725_n 0.00646998f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_428 N_VPWR_c_515_n Y 0.0369515f $X=7.915 $Y=2.02 $X2=0 $Y2=0
cc_429 N_VPWR_c_520_n Y 0.0228703f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_430 N_VPWR_c_510_n Y 0.0124393f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_431 N_VPWR_M1010_s N_Y_c_675_n 7.64275e-19 $X=6.83 $Y=1.485 $X2=0 $Y2=0
cc_432 N_VPWR_M1010_s N_Y_c_676_n 0.00123197f $X=6.83 $Y=1.485 $X2=0 $Y2=0
cc_433 N_VPWR_c_514_n N_Y_c_676_n 0.0193265f $X=6.975 $Y=2.02 $X2=0 $Y2=0
cc_434 N_VPWR_M1025_s N_Y_c_677_n 0.00200765f $X=7.77 $Y=1.485 $X2=0 $Y2=0
cc_435 N_VPWR_c_515_n N_Y_c_677_n 0.0193613f $X=7.915 $Y=2.02 $X2=0 $Y2=0
cc_436 N_A_497_297#_c_623_n N_Y_M1005_d 0.0121702f $X=5.13 $Y=2.165 $X2=0 $Y2=0
cc_437 N_A_497_297#_c_622_n N_Y_M1005_d 0.00201952f $X=4.53 $Y=2.165 $X2=0 $Y2=0
cc_438 N_A_497_297#_c_636_n N_Y_M1007_d 0.00348699f $X=6.035 $Y=1.95 $X2=0 $Y2=0
cc_439 N_A_497_297#_c_636_n N_Y_c_722_n 0.038481f $X=6.035 $Y=1.95 $X2=0 $Y2=0
cc_440 N_A_497_297#_M1005_s N_Y_c_674_n 0.0018979f $X=4.95 $Y=1.485 $X2=0 $Y2=0
cc_441 N_A_497_297#_M1018_s N_Y_c_674_n 0.0018979f $X=5.89 $Y=1.485 $X2=0 $Y2=0
cc_442 N_A_497_297#_c_632_n N_Y_c_674_n 0.00883579f $X=4.005 $Y=1.815 $X2=0
+ $Y2=0
cc_443 N_A_497_297#_c_622_n N_Y_c_674_n 0.128693f $X=4.53 $Y=2.165 $X2=0 $Y2=0
cc_444 N_Y_c_690_n N_A_31_47#_M1009_d 0.00402197f $X=7.915 $Y=0.76 $X2=0 $Y2=0
cc_445 N_Y_M1004_s N_A_31_47#_c_824_n 0.00400271f $X=6.79 $Y=0.235 $X2=0 $Y2=0
cc_446 N_Y_M1012_s N_A_31_47#_c_824_n 0.00401579f $X=7.73 $Y=0.235 $X2=0 $Y2=0
cc_447 N_Y_c_690_n N_A_31_47#_c_824_n 0.0560055f $X=7.915 $Y=0.76 $X2=0 $Y2=0
cc_448 N_Y_c_695_n N_A_31_47#_c_824_n 0.0137702f $X=6.877 $Y=0.885 $X2=0 $Y2=0
cc_449 N_Y_c_690_n N_A_31_47#_c_757_n 0.0158916f $X=7.915 $Y=0.76 $X2=0 $Y2=0
cc_450 N_Y_M1004_s N_VGND_c_916_n 0.00256987f $X=6.79 $Y=0.235 $X2=0 $Y2=0
cc_451 N_Y_M1012_s N_VGND_c_916_n 0.00256987f $X=7.73 $Y=0.235 $X2=0 $Y2=0
cc_452 N_A_31_47#_c_765_n N_VGND_M1003_s 0.00435938f $X=1.005 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_453 N_A_31_47#_c_775_n N_VGND_M1015_s 0.00574199f $X=1.945 $Y=0.8 $X2=0 $Y2=0
cc_454 N_A_31_47#_c_788_n N_VGND_M1008_d 0.00435938f $X=2.885 $Y=0.8 $X2=0 $Y2=0
cc_455 N_A_31_47#_c_796_n N_VGND_M1021_d 0.00574199f $X=3.825 $Y=0.8 $X2=0 $Y2=0
cc_456 N_A_31_47#_c_811_n N_VGND_M1000_d 0.016993f $X=5.36 $Y=0.8 $X2=0 $Y2=0
cc_457 N_A_31_47#_c_755_n N_VGND_M1023_d 0.00815115f $X=6.42 $Y=0.8 $X2=0 $Y2=0
cc_458 N_A_31_47#_c_753_n N_VGND_c_903_n 0.0176569f $X=0.28 $Y=0.38 $X2=0 $Y2=0
cc_459 N_A_31_47#_c_765_n N_VGND_c_903_n 0.0126475f $X=1.005 $Y=0.8 $X2=0 $Y2=0
cc_460 N_A_31_47#_c_765_n N_VGND_c_904_n 0.0020257f $X=1.005 $Y=0.8 $X2=0 $Y2=0
cc_461 N_A_31_47#_c_771_n N_VGND_c_904_n 0.022318f $X=1.22 $Y=0.36 $X2=0 $Y2=0
cc_462 N_A_31_47#_c_775_n N_VGND_c_904_n 0.00271675f $X=1.945 $Y=0.8 $X2=0 $Y2=0
cc_463 N_A_31_47#_c_771_n N_VGND_c_905_n 0.0177507f $X=1.22 $Y=0.36 $X2=0 $Y2=0
cc_464 N_A_31_47#_c_775_n N_VGND_c_905_n 0.0131159f $X=1.945 $Y=0.8 $X2=0 $Y2=0
cc_465 N_A_31_47#_c_779_n N_VGND_c_905_n 0.0216501f $X=2.16 $Y=0.36 $X2=0 $Y2=0
cc_466 N_A_31_47#_c_779_n N_VGND_c_906_n 0.0177507f $X=2.16 $Y=0.36 $X2=0 $Y2=0
cc_467 N_A_31_47#_c_788_n N_VGND_c_906_n 0.0126475f $X=2.885 $Y=0.8 $X2=0 $Y2=0
cc_468 N_A_31_47#_c_792_n N_VGND_c_907_n 0.0177507f $X=3.1 $Y=0.36 $X2=0 $Y2=0
cc_469 N_A_31_47#_c_796_n N_VGND_c_907_n 0.0131159f $X=3.825 $Y=0.8 $X2=0 $Y2=0
cc_470 N_A_31_47#_c_800_n N_VGND_c_907_n 0.0216501f $X=4.04 $Y=0.36 $X2=0 $Y2=0
cc_471 N_A_31_47#_c_755_n N_VGND_c_908_n 0.02873f $X=6.42 $Y=0.8 $X2=0 $Y2=0
cc_472 N_A_31_47#_c_775_n N_VGND_c_909_n 0.00203275f $X=1.945 $Y=0.8 $X2=0 $Y2=0
cc_473 N_A_31_47#_c_779_n N_VGND_c_909_n 0.0222117f $X=2.16 $Y=0.36 $X2=0 $Y2=0
cc_474 N_A_31_47#_c_788_n N_VGND_c_909_n 0.00271675f $X=2.885 $Y=0.8 $X2=0 $Y2=0
cc_475 N_A_31_47#_c_788_n N_VGND_c_911_n 0.0020257f $X=2.885 $Y=0.8 $X2=0 $Y2=0
cc_476 N_A_31_47#_c_792_n N_VGND_c_911_n 0.022318f $X=3.1 $Y=0.36 $X2=0 $Y2=0
cc_477 N_A_31_47#_c_796_n N_VGND_c_911_n 0.00271675f $X=3.825 $Y=0.8 $X2=0 $Y2=0
cc_478 N_A_31_47#_c_811_n N_VGND_c_913_n 0.00270993f $X=5.36 $Y=0.8 $X2=0 $Y2=0
cc_479 N_A_31_47#_c_865_p N_VGND_c_913_n 0.00593095f $X=5.445 $Y=0.56 $X2=0
+ $Y2=0
cc_480 N_A_31_47#_c_755_n N_VGND_c_913_n 0.00293388f $X=6.42 $Y=0.8 $X2=0 $Y2=0
cc_481 N_A_31_47#_c_755_n N_VGND_c_915_n 0.00293388f $X=6.42 $Y=0.8 $X2=0 $Y2=0
cc_482 N_A_31_47#_c_824_n N_VGND_c_915_n 0.0959059f $X=8.3 $Y=0.365 $X2=0 $Y2=0
cc_483 N_A_31_47#_c_869_p N_VGND_c_915_n 0.0114055f $X=6.59 $Y=0.365 $X2=0 $Y2=0
cc_484 N_A_31_47#_c_756_n N_VGND_c_915_n 0.0200319f $X=8.442 $Y=0.475 $X2=0
+ $Y2=0
cc_485 N_A_31_47#_M1003_d N_VGND_c_916_n 0.00209319f $X=0.155 $Y=0.235 $X2=0
+ $Y2=0
cc_486 N_A_31_47#_M1014_d N_VGND_c_916_n 0.0025535f $X=1.035 $Y=0.235 $X2=0
+ $Y2=0
cc_487 N_A_31_47#_M1026_d N_VGND_c_916_n 0.00215201f $X=2.025 $Y=0.235 $X2=0
+ $Y2=0
cc_488 N_A_31_47#_M1011_s N_VGND_c_916_n 0.0025535f $X=2.915 $Y=0.235 $X2=0
+ $Y2=0
cc_489 N_A_31_47#_M1029_s N_VGND_c_916_n 0.00215201f $X=3.905 $Y=0.235 $X2=0
+ $Y2=0
cc_490 N_A_31_47#_M1017_s N_VGND_c_916_n 0.00339454f $X=5.26 $Y=0.235 $X2=0
+ $Y2=0
cc_491 N_A_31_47#_M1027_s N_VGND_c_916_n 0.00240924f $X=6.37 $Y=0.235 $X2=0
+ $Y2=0
cc_492 N_A_31_47#_M1009_d N_VGND_c_916_n 0.00255381f $X=7.26 $Y=0.235 $X2=0
+ $Y2=0
cc_493 N_A_31_47#_M1022_d N_VGND_c_916_n 0.00250318f $X=8.2 $Y=0.235 $X2=0 $Y2=0
cc_494 N_A_31_47#_c_753_n N_VGND_c_916_n 0.0133626f $X=0.28 $Y=0.38 $X2=0 $Y2=0
cc_495 N_A_31_47#_c_765_n N_VGND_c_916_n 0.009788f $X=1.005 $Y=0.8 $X2=0 $Y2=0
cc_496 N_A_31_47#_c_771_n N_VGND_c_916_n 0.0141185f $X=1.22 $Y=0.36 $X2=0 $Y2=0
cc_497 N_A_31_47#_c_775_n N_VGND_c_916_n 0.0100794f $X=1.945 $Y=0.8 $X2=0 $Y2=0
cc_498 N_A_31_47#_c_779_n N_VGND_c_916_n 0.0138899f $X=2.16 $Y=0.36 $X2=0 $Y2=0
cc_499 N_A_31_47#_c_788_n N_VGND_c_916_n 0.009788f $X=2.885 $Y=0.8 $X2=0 $Y2=0
cc_500 N_A_31_47#_c_792_n N_VGND_c_916_n 0.0141185f $X=3.1 $Y=0.36 $X2=0 $Y2=0
cc_501 N_A_31_47#_c_796_n N_VGND_c_916_n 0.0100794f $X=3.825 $Y=0.8 $X2=0 $Y2=0
cc_502 N_A_31_47#_c_800_n N_VGND_c_916_n 0.0138899f $X=4.04 $Y=0.36 $X2=0 $Y2=0
cc_503 N_A_31_47#_c_811_n N_VGND_c_916_n 0.0137173f $X=5.36 $Y=0.8 $X2=0 $Y2=0
cc_504 N_A_31_47#_c_865_p N_VGND_c_916_n 0.00590828f $X=5.445 $Y=0.56 $X2=0
+ $Y2=0
cc_505 N_A_31_47#_c_755_n N_VGND_c_916_n 0.0138213f $X=6.42 $Y=0.8 $X2=0 $Y2=0
cc_506 N_A_31_47#_c_824_n N_VGND_c_916_n 0.0610924f $X=8.3 $Y=0.365 $X2=0 $Y2=0
cc_507 N_A_31_47#_c_869_p N_VGND_c_916_n 0.0065339f $X=6.59 $Y=0.365 $X2=0 $Y2=0
cc_508 N_A_31_47#_c_756_n N_VGND_c_916_n 0.010954f $X=8.442 $Y=0.475 $X2=0 $Y2=0
cc_509 N_A_31_47#_c_753_n N_VGND_c_917_n 0.0227138f $X=0.28 $Y=0.38 $X2=0 $Y2=0
cc_510 N_A_31_47#_c_765_n N_VGND_c_917_n 0.00271675f $X=1.005 $Y=0.8 $X2=0 $Y2=0
cc_511 N_A_31_47#_c_796_n N_VGND_c_919_n 0.00203275f $X=3.825 $Y=0.8 $X2=0 $Y2=0
cc_512 N_A_31_47#_c_800_n N_VGND_c_919_n 0.0222117f $X=4.04 $Y=0.36 $X2=0 $Y2=0
cc_513 N_A_31_47#_c_811_n N_VGND_c_919_n 0.00301228f $X=5.36 $Y=0.8 $X2=0 $Y2=0
cc_514 N_A_31_47#_c_800_n N_VGND_c_920_n 0.0185147f $X=4.04 $Y=0.36 $X2=0 $Y2=0
cc_515 N_A_31_47#_c_811_n N_VGND_c_920_n 0.04936f $X=5.36 $Y=0.8 $X2=0 $Y2=0
cc_516 N_A_31_47#_c_865_p N_VGND_c_920_n 0.00960516f $X=5.445 $Y=0.56 $X2=0
+ $Y2=0
