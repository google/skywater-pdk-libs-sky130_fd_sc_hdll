* File: sky130_fd_sc_hdll__o22a_1.spice
* Created: Thu Aug 27 19:20:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o22a_1.pex.spice"
.subckt sky130_fd_sc_hdll__o22a_1  VNB VPB B1 B2 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_83_21#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.182 PD=1.82 PS=1.86 NRD=0 NRS=2.76 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_A_83_21#_M1008_d N_B1_M1008_g N_A_219_47#_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1009 N_A_219_47#_M1009_d N_B2_M1009_g N_A_83_21#_M1008_d VNB NSHORT L=0.15
+ W=0.65 AD=0.143 AS=0.08775 PD=1.09 PS=0.92 NRD=30.456 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_219_47#_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.143 PD=0.98 PS=1.09 NRD=10.152 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1004 N_A_219_47#_M1004_d N_A1_M1004_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.10725 PD=1.92 PS=0.98 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_A_83_21#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.355 AS=0.29 PD=1.71 PS=2.58 NRD=4.9053 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1005 A_299_297# N_B1_M1005_g N_VPWR_M1001_d VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.355 PD=1.29 PS=1.71 NRD=17.7103 NRS=9.8303 M=1 R=5.55556 SA=90001.1
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1003 N_A_83_21#_M1003_d N_B2_M1003_g A_299_297# VPB PHIGHVT L=0.18 W=1
+ AD=0.205 AS=0.145 PD=1.41 PS=1.29 NRD=0.9653 NRS=17.7103 M=1 R=5.55556
+ SA=90001.6 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1007 A_511_297# N_A2_M1007_g N_A_83_21#_M1003_d VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.205 PD=1.3 PS=1.41 NRD=18.6953 NRS=24.6053 M=1 R=5.55556 SA=90002.1
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g A_511_297# VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.15 PD=2.54 PS=1.3 NRD=0.9653 NRS=18.6953 M=1 R=5.55556 SA=90002.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hdll__o22a_1.pxi.spice"
*
.ends
*
*
