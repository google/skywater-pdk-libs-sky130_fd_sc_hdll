* File: sky130_fd_sc_hdll__inv_4.spice
* Created: Thu Aug 27 19:09:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__inv_4.pex.spice"
.subckt sky130_fd_sc_hdll__inv_4  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_Y_M1002_d N_A_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.2015 PD=0.97 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2 SB=75001.8
+ A=0.0975 P=1.6 MULT=1
MM1003 N_Y_M1002_d N_A_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.7 SB=75001.4
+ A=0.0975 P=1.6 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.2 SB=75000.9
+ A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1005_d N_A_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.32825 PD=0.97 PS=2.31 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.6 SB=75000.4
+ A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90001.8 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_Y_M1000_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.6
+ SB=90001.4 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1001_d N_A_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.1
+ SB=90000.9 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_Y_M1004_s VPB PHIGHVT L=0.18 W=1 AD=0.515
+ AS=0.145 PD=3.03 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.6
+ SB=90000.4 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hdll__inv_4.pxi.spice"
*
.ends
*
*
