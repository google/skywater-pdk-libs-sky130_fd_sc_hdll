# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a21o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.410000 0.365000 2.730000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.160000 0.750000 3.535000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.865000 0.995000 2.240000 1.410000 ;
    END
  END B1
  PIN VGND
    ANTENNADIFFAREA  0.854750 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  0.935000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  0.629500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.255000 0.825000 2.465000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.095000  1.665000 0.375000 2.635000 ;
      RECT 0.175000  0.085000 0.345000 0.555000 ;
      RECT 0.995000  0.655000 2.240000 0.825000 ;
      RECT 0.995000  0.825000 1.430000 1.690000 ;
      RECT 0.995000  1.690000 2.040000 1.920000 ;
      RECT 1.055000  2.220000 1.485000 2.635000 ;
      RECT 1.275000  0.085000 1.655000 0.445000 ;
      RECT 1.675000  1.920000 2.040000 2.465000 ;
      RECT 2.050000  0.255000 2.240000 0.655000 ;
      RECT 2.260000  1.670000 3.475000 1.935000 ;
      RECT 2.260000  1.935000 2.485000 2.465000 ;
      RECT 2.705000  2.125000 3.035000 2.635000 ;
      RECT 3.155000  0.085000 3.535000 0.565000 ;
      RECT 3.255000  1.935000 3.475000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21o_2
