* File: sky130_fd_sc_hdll__a21o_4.pxi.spice
* Created: Wed Sep  2 08:17:19 2020
* 
x_PM_SKY130_FD_SC_HDLL__A21O_4%A_84_21# N_A_84_21#_M1000_s N_A_84_21#_M1017_s
+ N_A_84_21#_M1011_s N_A_84_21#_c_76_n N_A_84_21#_M1002_g N_A_84_21#_c_84_n
+ N_A_84_21#_M1003_g N_A_84_21#_c_77_n N_A_84_21#_M1005_g N_A_84_21#_c_85_n
+ N_A_84_21#_M1012_g N_A_84_21#_c_78_n N_A_84_21#_M1008_g N_A_84_21#_c_86_n
+ N_A_84_21#_M1018_g N_A_84_21#_c_79_n N_A_84_21#_M1016_g N_A_84_21#_c_87_n
+ N_A_84_21#_M1019_g N_A_84_21#_c_80_n N_A_84_21#_c_81_n N_A_84_21#_c_92_p
+ N_A_84_21#_c_142_p N_A_84_21#_c_171_p N_A_84_21#_c_82_n N_A_84_21#_c_97_p
+ N_A_84_21#_c_117_p N_A_84_21#_c_83_n PM_SKY130_FD_SC_HDLL__A21O_4%A_84_21#
x_PM_SKY130_FD_SC_HDLL__A21O_4%B1 N_B1_c_201_n N_B1_M1000_g N_B1_c_205_n
+ N_B1_M1011_g N_B1_c_206_n N_B1_M1014_g N_B1_c_202_n N_B1_M1006_g B1
+ N_B1_c_204_n B1 PM_SKY130_FD_SC_HDLL__A21O_4%B1
x_PM_SKY130_FD_SC_HDLL__A21O_4%A2 N_A2_c_251_n N_A2_M1004_g N_A2_c_252_n
+ N_A2_M1007_g N_A2_c_253_n N_A2_M1010_g N_A2_c_254_n N_A2_M1013_g N_A2_c_255_n
+ N_A2_c_267_n N_A2_c_297_p A2 N_A2_c_256_n N_A2_c_257_n A2 N_A2_c_300_p
+ PM_SKY130_FD_SC_HDLL__A21O_4%A2
x_PM_SKY130_FD_SC_HDLL__A21O_4%A1 N_A1_c_335_n N_A1_M1017_g N_A1_c_339_n
+ N_A1_M1001_g N_A1_c_340_n N_A1_M1015_g N_A1_c_336_n N_A1_M1009_g A1
+ N_A1_c_338_n A1 PM_SKY130_FD_SC_HDLL__A21O_4%A1
x_PM_SKY130_FD_SC_HDLL__A21O_4%VPWR N_VPWR_M1003_d N_VPWR_M1012_d N_VPWR_M1019_d
+ N_VPWR_M1004_d N_VPWR_M1015_s N_VPWR_c_382_n N_VPWR_c_383_n N_VPWR_c_384_n
+ N_VPWR_c_385_n N_VPWR_c_386_n N_VPWR_c_387_n N_VPWR_c_388_n N_VPWR_c_389_n
+ N_VPWR_c_390_n VPWR N_VPWR_c_391_n N_VPWR_c_392_n N_VPWR_c_381_n
+ N_VPWR_c_394_n N_VPWR_c_395_n PM_SKY130_FD_SC_HDLL__A21O_4%VPWR
x_PM_SKY130_FD_SC_HDLL__A21O_4%X N_X_M1002_d N_X_M1008_d N_X_M1003_s N_X_M1018_s
+ N_X_c_508_n N_X_c_485_n N_X_c_486_n N_X_c_492_n N_X_c_496_n N_X_c_499_n X X
+ PM_SKY130_FD_SC_HDLL__A21O_4%X
x_PM_SKY130_FD_SC_HDLL__A21O_4%A_523_297# N_A_523_297#_M1011_d
+ N_A_523_297#_M1014_d N_A_523_297#_M1001_d N_A_523_297#_M1013_s
+ N_A_523_297#_c_534_n N_A_523_297#_c_535_n N_A_523_297#_c_575_n
+ N_A_523_297#_c_531_n N_A_523_297#_c_551_n N_A_523_297#_c_552_n
+ N_A_523_297#_c_584_n N_A_523_297#_c_556_n N_A_523_297#_c_532_n
+ N_A_523_297#_c_562_n N_A_523_297#_c_533_n
+ PM_SKY130_FD_SC_HDLL__A21O_4%A_523_297#
x_PM_SKY130_FD_SC_HDLL__A21O_4%VGND N_VGND_M1002_s N_VGND_M1005_s N_VGND_M1016_s
+ N_VGND_M1006_d N_VGND_M1010_d N_VGND_c_597_n N_VGND_c_598_n N_VGND_c_599_n
+ N_VGND_c_600_n N_VGND_c_601_n N_VGND_c_602_n N_VGND_c_603_n VGND
+ N_VGND_c_604_n N_VGND_c_605_n N_VGND_c_606_n N_VGND_c_607_n N_VGND_c_608_n
+ N_VGND_c_609_n PM_SKY130_FD_SC_HDLL__A21O_4%VGND
cc_1 VNB N_A_84_21#_c_76_n 0.0191599f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.995
cc_2 VNB N_A_84_21#_c_77_n 0.0169217f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=0.995
cc_3 VNB N_A_84_21#_c_78_n 0.0169495f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=0.995
cc_4 VNB N_A_84_21#_c_79_n 0.0197939f $X=-0.19 $Y=-0.24 $X2=1.935 $Y2=0.995
cc_5 VNB N_A_84_21#_c_80_n 0.00223883f $X=-0.19 $Y=-0.24 $X2=2.13 $Y2=1.16
cc_6 VNB N_A_84_21#_c_81_n 0.002509f $X=-0.19 $Y=-0.24 $X2=2.215 $Y2=0.995
cc_7 VNB N_A_84_21#_c_82_n 0.00202969f $X=-0.19 $Y=-0.24 $X2=3.21 $Y2=1.62
cc_8 VNB N_A_84_21#_c_83_n 0.0912528f $X=-0.19 $Y=-0.24 $X2=1.96 $Y2=1.202
cc_9 VNB N_B1_c_201_n 0.0202034f $X=-0.19 $Y=-0.24 $X2=3.025 $Y2=0.235
cc_10 VNB N_B1_c_202_n 0.0174882f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.995
cc_11 VNB B1 0.00406946f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.41
cc_12 VNB N_B1_c_204_n 0.0498307f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.985
cc_13 VNB N_A2_c_251_n 0.0213831f $X=-0.19 $Y=-0.24 $X2=3.025 $Y2=0.235
cc_14 VNB N_A2_c_252_n 0.0166832f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A2_c_253_n 0.0222254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A2_c_254_n 0.0316003f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.995
cc_17 VNB N_A2_c_255_n 5.56894e-19 $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.985
cc_18 VNB N_A2_c_256_n 0.00551268f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=0.56
cc_19 VNB N_A2_c_257_n 0.0153855f $X=-0.19 $Y=-0.24 $X2=1.935 $Y2=0.56
cc_20 VNB A2 4.09545e-19 $X=-0.19 $Y=-0.24 $X2=1.96 $Y2=1.985
cc_21 VNB N_A1_c_335_n 0.0172715f $X=-0.19 $Y=-0.24 $X2=3.025 $Y2=0.235
cc_22 VNB N_A1_c_336_n 0.0171772f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.995
cc_23 VNB A1 0.0024063f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.41
cc_24 VNB N_A1_c_338_n 0.0360975f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.985
cc_25 VNB N_VPWR_c_381_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.202
cc_26 VNB X 0.0193267f $X=-0.19 $Y=-0.24 $X2=1.96 $Y2=1.985
cc_27 VNB N_VGND_c_597_n 0.0108424f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=0.995
cc_28 VNB N_VGND_c_598_n 0.0119235f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=0.56
cc_29 VNB N_VGND_c_599_n 0.00227328f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=0.995
cc_30 VNB N_VGND_c_600_n 0.0157208f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=0.56
cc_31 VNB N_VGND_c_601_n 0.0331548f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=1.985
cc_32 VNB N_VGND_c_602_n 0.0164201f $X=-0.19 $Y=-0.24 $X2=1.935 $Y2=0.56
cc_33 VNB N_VGND_c_603_n 0.00507043f $X=-0.19 $Y=-0.24 $X2=1.935 $Y2=0.56
cc_34 VNB N_VGND_c_604_n 0.0136465f $X=-0.19 $Y=-0.24 $X2=1.96 $Y2=1.985
cc_35 VNB N_VGND_c_605_n 0.0440873f $X=-0.19 $Y=-0.24 $X2=3.21 $Y2=0.42
cc_36 VNB N_VGND_c_606_n 0.00546647f $X=-0.19 $Y=-0.24 $X2=4.62 $Y2=0.57
cc_37 VNB N_VGND_c_607_n 0.0191309f $X=-0.19 $Y=-0.24 $X2=1.26 $Y2=1.202
cc_38 VNB N_VGND_c_608_n 0.0191071f $X=-0.19 $Y=-0.24 $X2=1.935 $Y2=1.202
cc_39 VNB N_VGND_c_609_n 0.301236f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VPB N_A_84_21#_c_84_n 0.0185522f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.41
cc_41 VPB N_A_84_21#_c_85_n 0.0159888f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.41
cc_42 VPB N_A_84_21#_c_86_n 0.0162845f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=1.41
cc_43 VPB N_A_84_21#_c_87_n 0.0196726f $X=-0.19 $Y=1.305 $X2=1.96 $Y2=1.41
cc_44 VPB N_A_84_21#_c_80_n 0.00180214f $X=-0.19 $Y=1.305 $X2=2.13 $Y2=1.16
cc_45 VPB N_A_84_21#_c_82_n 0.00240585f $X=-0.19 $Y=1.305 $X2=3.21 $Y2=1.62
cc_46 VPB N_A_84_21#_c_83_n 0.0531128f $X=-0.19 $Y=1.305 $X2=1.96 $Y2=1.202
cc_47 VPB N_B1_c_205_n 0.0196006f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_B1_c_206_n 0.0164022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB B1 0.00744247f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.41
cc_50 VPB N_B1_c_204_n 0.0307902f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.985
cc_51 VPB N_A2_c_251_n 0.0254576f $X=-0.19 $Y=1.305 $X2=3.025 $Y2=0.235
cc_52 VPB N_A2_c_254_n 0.030702f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=0.995
cc_53 VPB N_A2_c_255_n 0.00173479f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.985
cc_54 VPB A2 0.00706632f $X=-0.19 $Y=1.305 $X2=1.96 $Y2=1.985
cc_55 VPB N_A1_c_339_n 0.0162056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A1_c_340_n 0.0159302f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A1_c_338_n 0.0195829f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.985
cc_58 VPB N_VPWR_c_382_n 0.0110369f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=0.995
cc_59 VPB N_VPWR_c_383_n 0.0243557f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=0.56
cc_60 VPB N_VPWR_c_384_n 3.38371e-19 $X=-0.19 $Y=1.305 $X2=1.455 $Y2=0.995
cc_61 VPB N_VPWR_c_385_n 0.018546f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=0.56
cc_62 VPB N_VPWR_c_386_n 0.00464386f $X=-0.19 $Y=1.305 $X2=1.935 $Y2=0.995
cc_63 VPB N_VPWR_c_387_n 0.00547137f $X=-0.19 $Y=1.305 $X2=1.96 $Y2=1.985
cc_64 VPB N_VPWR_c_388_n 0.0390762f $X=-0.19 $Y=1.305 $X2=1.26 $Y2=1.16
cc_65 VPB N_VPWR_c_389_n 0.00547137f $X=-0.19 $Y=1.305 $X2=1.99 $Y2=1.16
cc_66 VPB N_VPWR_c_390_n 0.0125866f $X=-0.19 $Y=1.305 $X2=2.215 $Y2=0.995
cc_67 VPB N_VPWR_c_391_n 0.0153876f $X=-0.19 $Y=1.305 $X2=3.21 $Y2=0.42
cc_68 VPB N_VPWR_c_392_n 0.0204162f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_69 VPB N_VPWR_c_381_n 0.0572424f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.202
cc_70 VPB N_VPWR_c_394_n 0.00503453f $X=-0.19 $Y=1.305 $X2=1.96 $Y2=1.202
cc_71 VPB N_VPWR_c_395_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB X 0.00958328f $X=-0.19 $Y=1.305 $X2=1.96 $Y2=1.985
cc_73 VPB N_A_523_297#_c_531_n 0.00333169f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.985
cc_74 VPB N_A_523_297#_c_532_n 0.0223011f $X=-0.19 $Y=1.305 $X2=1.99 $Y2=1.16
cc_75 VPB N_A_523_297#_c_533_n 0.0219742f $X=-0.19 $Y=1.305 $X2=2.3 $Y2=0.7
cc_76 N_A_84_21#_c_81_n N_B1_c_201_n 0.00468314f $X=2.215 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_77 N_A_84_21#_c_92_p N_B1_c_201_n 0.0153595f $X=3.125 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_78 N_A_84_21#_c_82_n N_B1_c_201_n 0.00341454f $X=3.21 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_79 N_A_84_21#_c_82_n N_B1_c_205_n 0.00603273f $X=3.21 $Y=1.62 $X2=0 $Y2=0
cc_80 N_A_84_21#_c_82_n N_B1_c_206_n 0.00364403f $X=3.21 $Y=1.62 $X2=0 $Y2=0
cc_81 N_A_84_21#_c_82_n N_B1_c_202_n 0.00341454f $X=3.21 $Y=1.62 $X2=0 $Y2=0
cc_82 N_A_84_21#_c_97_p N_B1_c_202_n 0.0146172f $X=4.485 $Y=0.755 $X2=0 $Y2=0
cc_83 N_A_84_21#_c_87_n B1 0.00264541f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_84_21#_c_80_n B1 0.0264328f $X=2.13 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_84_21#_c_92_p B1 0.0253655f $X=3.125 $Y=0.7 $X2=0 $Y2=0
cc_86 N_A_84_21#_c_82_n B1 0.0319957f $X=3.21 $Y=1.62 $X2=0 $Y2=0
cc_87 N_A_84_21#_c_83_n B1 0.0035725f $X=1.96 $Y=1.202 $X2=0 $Y2=0
cc_88 N_A_84_21#_c_80_n N_B1_c_204_n 0.00103082f $X=2.13 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A_84_21#_c_92_p N_B1_c_204_n 0.00435174f $X=3.125 $Y=0.7 $X2=0 $Y2=0
cc_90 N_A_84_21#_c_82_n N_B1_c_204_n 0.0259168f $X=3.21 $Y=1.62 $X2=0 $Y2=0
cc_91 N_A_84_21#_c_97_p N_B1_c_204_n 3.64185e-19 $X=4.485 $Y=0.755 $X2=0 $Y2=0
cc_92 N_A_84_21#_c_83_n N_B1_c_204_n 0.00622977f $X=1.96 $Y=1.202 $X2=0 $Y2=0
cc_93 N_A_84_21#_c_82_n N_A2_c_251_n 4.32833e-19 $X=3.21 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_94 N_A_84_21#_c_97_p N_A2_c_251_n 0.00376359f $X=4.485 $Y=0.755 $X2=-0.19
+ $Y2=-0.24
cc_95 N_A_84_21#_c_97_p N_A2_c_252_n 0.0118368f $X=4.485 $Y=0.755 $X2=0 $Y2=0
cc_96 N_A_84_21#_c_82_n N_A2_c_255_n 0.00424417f $X=3.21 $Y=1.62 $X2=0 $Y2=0
cc_97 N_A_84_21#_c_97_p N_A2_c_267_n 0.00269265f $X=4.485 $Y=0.755 $X2=0 $Y2=0
cc_98 N_A_84_21#_c_82_n N_A2_c_256_n 0.0102371f $X=3.21 $Y=1.62 $X2=0 $Y2=0
cc_99 N_A_84_21#_c_97_p N_A2_c_256_n 0.0283014f $X=4.485 $Y=0.755 $X2=0 $Y2=0
cc_100 N_A_84_21#_c_97_p N_A1_c_335_n 0.0112278f $X=4.485 $Y=0.755 $X2=-0.19
+ $Y2=-0.24
cc_101 N_A_84_21#_c_97_p A1 0.00848049f $X=4.485 $Y=0.755 $X2=0 $Y2=0
cc_102 N_A_84_21#_c_117_p A1 0.0208871f $X=4.62 $Y=0.57 $X2=0 $Y2=0
cc_103 N_A_84_21#_c_117_p N_A1_c_338_n 0.00444199f $X=4.62 $Y=0.57 $X2=0 $Y2=0
cc_104 N_A_84_21#_c_84_n N_VPWR_c_383_n 0.0132681f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A_84_21#_c_85_n N_VPWR_c_383_n 0.00127849f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_106 N_A_84_21#_c_84_n N_VPWR_c_384_n 0.00140714f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_107 N_A_84_21#_c_85_n N_VPWR_c_384_n 0.0160003f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A_84_21#_c_86_n N_VPWR_c_384_n 0.0127678f $X=1.48 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A_84_21#_c_87_n N_VPWR_c_384_n 0.00125009f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A_84_21#_c_86_n N_VPWR_c_385_n 0.00642146f $X=1.48 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A_84_21#_c_87_n N_VPWR_c_385_n 0.00686042f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A_84_21#_c_87_n N_VPWR_c_386_n 0.00348927f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_84_21#_c_80_n N_VPWR_c_386_n 0.0173684f $X=2.13 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_84_21#_c_83_n N_VPWR_c_386_n 0.00169403f $X=1.96 $Y=1.202 $X2=0 $Y2=0
cc_115 N_A_84_21#_c_84_n N_VPWR_c_391_n 0.00642146f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A_84_21#_c_85_n N_VPWR_c_391_n 0.00447018f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A_84_21#_M1011_s N_VPWR_c_381_n 0.00232895f $X=3.065 $Y=1.485 $X2=0
+ $Y2=0
cc_118 N_A_84_21#_c_84_n N_VPWR_c_381_n 0.0108125f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_84_21#_c_85_n N_VPWR_c_381_n 0.00774115f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_84_21#_c_86_n N_VPWR_c_381_n 0.0108125f $X=1.48 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_84_21#_c_87_n N_VPWR_c_381_n 0.0133008f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A_84_21#_c_76_n N_X_c_485_n 0.00884112f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_84_21#_c_77_n N_X_c_486_n 0.0100176f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A_84_21#_c_78_n N_X_c_486_n 0.0100176f $X=1.455 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_84_21#_c_79_n N_X_c_486_n 0.00302279f $X=1.935 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_84_21#_c_80_n N_X_c_486_n 0.0554287f $X=2.13 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A_84_21#_c_142_p N_X_c_486_n 0.0110614f $X=2.3 $Y=0.7 $X2=0 $Y2=0
cc_128 N_A_84_21#_c_83_n N_X_c_486_n 0.011212f $X=1.96 $Y=1.202 $X2=0 $Y2=0
cc_129 N_A_84_21#_c_85_n N_X_c_492_n 0.0140207f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_84_21#_c_86_n N_X_c_492_n 0.0155294f $X=1.48 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A_84_21#_c_80_n N_X_c_492_n 0.0348222f $X=2.13 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_84_21#_c_83_n N_X_c_492_n 0.00856313f $X=1.96 $Y=1.202 $X2=0 $Y2=0
cc_133 N_A_84_21#_c_87_n N_X_c_496_n 0.00210376f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_84_21#_c_80_n N_X_c_496_n 0.0128389f $X=2.13 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_84_21#_c_83_n N_X_c_496_n 0.00510469f $X=1.96 $Y=1.202 $X2=0 $Y2=0
cc_136 N_A_84_21#_c_87_n N_X_c_499_n 0.00495081f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A_84_21#_c_76_n X 0.00783436f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A_84_21#_c_84_n X 0.0217938f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_84_21#_c_77_n X 0.00485153f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_84_21#_c_85_n X 0.00392509f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_84_21#_c_80_n X 0.0271307f $X=2.13 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_84_21#_c_83_n X 0.0336972f $X=1.96 $Y=1.202 $X2=0 $Y2=0
cc_143 N_A_84_21#_c_82_n N_A_523_297#_c_534_n 0.0205562f $X=3.21 $Y=1.62 $X2=0
+ $Y2=0
cc_144 N_A_84_21#_M1011_s N_A_523_297#_c_535_n 0.00336374f $X=3.065 $Y=1.485
+ $X2=0 $Y2=0
cc_145 N_A_84_21#_c_82_n N_A_523_297#_c_535_n 0.0128008f $X=3.21 $Y=1.62 $X2=0
+ $Y2=0
cc_146 N_A_84_21#_c_82_n N_A_523_297#_c_531_n 0.0110013f $X=3.21 $Y=1.62 $X2=0
+ $Y2=0
cc_147 N_A_84_21#_c_97_p N_A_523_297#_c_531_n 0.00440519f $X=4.485 $Y=0.755
+ $X2=0 $Y2=0
cc_148 N_A_84_21#_c_81_n N_VGND_M1016_s 0.00301068f $X=2.215 $Y=0.995 $X2=0
+ $Y2=0
cc_149 N_A_84_21#_c_92_p N_VGND_M1016_s 0.0199211f $X=3.125 $Y=0.7 $X2=0 $Y2=0
cc_150 N_A_84_21#_c_142_p N_VGND_M1016_s 0.00507425f $X=2.3 $Y=0.7 $X2=0 $Y2=0
cc_151 N_A_84_21#_c_97_p N_VGND_M1006_d 0.00540394f $X=4.485 $Y=0.755 $X2=0
+ $Y2=0
cc_152 N_A_84_21#_c_76_n N_VGND_c_598_n 0.00905306f $X=0.495 $Y=0.995 $X2=0
+ $Y2=0
cc_153 N_A_84_21#_c_77_n N_VGND_c_598_n 0.00105862f $X=0.975 $Y=0.995 $X2=0
+ $Y2=0
cc_154 N_A_84_21#_c_97_p N_VGND_c_599_n 0.0133243f $X=4.485 $Y=0.755 $X2=0 $Y2=0
cc_155 N_A_84_21#_c_92_p N_VGND_c_602_n 0.00375101f $X=3.125 $Y=0.7 $X2=0 $Y2=0
cc_156 N_A_84_21#_c_171_p N_VGND_c_602_n 0.0118139f $X=3.21 $Y=0.42 $X2=0 $Y2=0
cc_157 N_A_84_21#_c_97_p N_VGND_c_602_n 0.00353953f $X=4.485 $Y=0.755 $X2=0
+ $Y2=0
cc_158 N_A_84_21#_c_76_n N_VGND_c_604_n 0.00350947f $X=0.495 $Y=0.995 $X2=0
+ $Y2=0
cc_159 N_A_84_21#_c_77_n N_VGND_c_604_n 0.0035176f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A_84_21#_c_97_p N_VGND_c_605_n 0.00822153f $X=4.485 $Y=0.755 $X2=0
+ $Y2=0
cc_161 N_A_84_21#_c_117_p N_VGND_c_605_n 0.00922285f $X=4.62 $Y=0.57 $X2=0 $Y2=0
cc_162 N_A_84_21#_c_76_n N_VGND_c_606_n 0.00106058f $X=0.495 $Y=0.995 $X2=0
+ $Y2=0
cc_163 N_A_84_21#_c_77_n N_VGND_c_606_n 0.00819243f $X=0.975 $Y=0.995 $X2=0
+ $Y2=0
cc_164 N_A_84_21#_c_78_n N_VGND_c_606_n 0.00939017f $X=1.455 $Y=0.995 $X2=0
+ $Y2=0
cc_165 N_A_84_21#_c_79_n N_VGND_c_606_n 0.00196005f $X=1.935 $Y=0.995 $X2=0
+ $Y2=0
cc_166 N_A_84_21#_c_78_n N_VGND_c_607_n 0.0035176f $X=1.455 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_84_21#_c_79_n N_VGND_c_607_n 0.00558173f $X=1.935 $Y=0.995 $X2=0
+ $Y2=0
cc_168 N_A_84_21#_c_79_n N_VGND_c_608_n 0.013604f $X=1.935 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_84_21#_c_80_n N_VGND_c_608_n 6.31205e-19 $X=2.13 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_84_21#_c_92_p N_VGND_c_608_n 0.0396902f $X=3.125 $Y=0.7 $X2=0 $Y2=0
cc_171 N_A_84_21#_c_142_p N_VGND_c_608_n 0.0141996f $X=2.3 $Y=0.7 $X2=0 $Y2=0
cc_172 N_A_84_21#_c_171_p N_VGND_c_608_n 0.0113729f $X=3.21 $Y=0.42 $X2=0 $Y2=0
cc_173 N_A_84_21#_c_83_n N_VGND_c_608_n 5.08643e-19 $X=1.96 $Y=1.202 $X2=0 $Y2=0
cc_174 N_A_84_21#_M1000_s N_VGND_c_609_n 0.00368335f $X=3.025 $Y=0.235 $X2=0
+ $Y2=0
cc_175 N_A_84_21#_M1017_s N_VGND_c_609_n 0.00481352f $X=4.435 $Y=0.235 $X2=0
+ $Y2=0
cc_176 N_A_84_21#_c_76_n N_VGND_c_609_n 0.00424411f $X=0.495 $Y=0.995 $X2=0
+ $Y2=0
cc_177 N_A_84_21#_c_77_n N_VGND_c_609_n 0.00424616f $X=0.975 $Y=0.995 $X2=0
+ $Y2=0
cc_178 N_A_84_21#_c_78_n N_VGND_c_609_n 0.00424616f $X=1.455 $Y=0.995 $X2=0
+ $Y2=0
cc_179 N_A_84_21#_c_79_n N_VGND_c_609_n 0.011515f $X=1.935 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_84_21#_c_92_p N_VGND_c_609_n 0.00884454f $X=3.125 $Y=0.7 $X2=0 $Y2=0
cc_181 N_A_84_21#_c_142_p N_VGND_c_609_n 8.9526e-19 $X=2.3 $Y=0.7 $X2=0 $Y2=0
cc_182 N_A_84_21#_c_171_p N_VGND_c_609_n 0.00646998f $X=3.21 $Y=0.42 $X2=0 $Y2=0
cc_183 N_A_84_21#_c_97_p N_VGND_c_609_n 0.0230737f $X=4.485 $Y=0.755 $X2=0 $Y2=0
cc_184 N_A_84_21#_c_117_p N_VGND_c_609_n 0.00967148f $X=4.62 $Y=0.57 $X2=0 $Y2=0
cc_185 N_A_84_21#_c_97_p A_801_47# 0.00534504f $X=4.485 $Y=0.755 $X2=-0.19
+ $Y2=-0.24
cc_186 N_B1_c_206_n N_A2_c_251_n 0.0200339f $X=3.445 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_187 N_B1_c_204_n N_A2_c_251_n 0.0260722f $X=3.445 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_188 N_B1_c_202_n N_A2_c_252_n 0.0235601f $X=3.47 $Y=0.995 $X2=0 $Y2=0
cc_189 N_B1_c_204_n N_A2_c_255_n 4.38741e-19 $X=3.445 $Y=1.202 $X2=0 $Y2=0
cc_190 N_B1_c_204_n N_A2_c_256_n 0.00256018f $X=3.445 $Y=1.202 $X2=0 $Y2=0
cc_191 N_B1_c_205_n N_VPWR_c_386_n 0.00786241f $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_192 B1 N_VPWR_c_386_n 6.92321e-19 $X=2.665 $Y=1.105 $X2=0 $Y2=0
cc_193 N_B1_c_206_n N_VPWR_c_387_n 0.00128781f $X=3.445 $Y=1.41 $X2=0 $Y2=0
cc_194 N_B1_c_205_n N_VPWR_c_388_n 0.00429453f $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_195 N_B1_c_206_n N_VPWR_c_388_n 0.00429453f $X=3.445 $Y=1.41 $X2=0 $Y2=0
cc_196 N_B1_c_205_n N_VPWR_c_381_n 0.00743756f $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_197 N_B1_c_206_n N_VPWR_c_381_n 0.00613207f $X=3.445 $Y=1.41 $X2=0 $Y2=0
cc_198 B1 N_A_523_297#_M1011_d 0.00372784f $X=2.665 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_199 B1 N_A_523_297#_c_534_n 0.0148026f $X=2.665 $Y=1.105 $X2=0 $Y2=0
cc_200 N_B1_c_204_n N_A_523_297#_c_534_n 6.95229e-19 $X=3.445 $Y=1.202 $X2=0
+ $Y2=0
cc_201 N_B1_c_205_n N_A_523_297#_c_535_n 0.0154468f $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_202 N_B1_c_206_n N_A_523_297#_c_535_n 0.0159634f $X=3.445 $Y=1.41 $X2=0 $Y2=0
cc_203 N_B1_c_206_n N_A_523_297#_c_531_n 5.67531e-19 $X=3.445 $Y=1.41 $X2=0
+ $Y2=0
cc_204 N_B1_c_202_n N_VGND_c_599_n 0.00178749f $X=3.47 $Y=0.995 $X2=0 $Y2=0
cc_205 N_B1_c_201_n N_VGND_c_602_n 0.00393283f $X=2.95 $Y=0.995 $X2=0 $Y2=0
cc_206 N_B1_c_202_n N_VGND_c_602_n 0.00430182f $X=3.47 $Y=0.995 $X2=0 $Y2=0
cc_207 N_B1_c_201_n N_VGND_c_608_n 0.00766662f $X=2.95 $Y=0.995 $X2=0 $Y2=0
cc_208 N_B1_c_202_n N_VGND_c_608_n 5.01938e-19 $X=3.47 $Y=0.995 $X2=0 $Y2=0
cc_209 N_B1_c_201_n N_VGND_c_609_n 0.00469688f $X=2.95 $Y=0.995 $X2=0 $Y2=0
cc_210 N_B1_c_202_n N_VGND_c_609_n 0.00601695f $X=3.47 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A2_c_252_n N_A1_c_335_n 0.0418594f $X=3.93 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_212 N_A2_c_251_n N_A1_c_339_n 0.0381051f $X=3.915 $Y=1.41 $X2=0 $Y2=0
cc_213 N_A2_c_255_n N_A1_c_339_n 0.00231141f $X=4.057 $Y=1.51 $X2=0 $Y2=0
cc_214 N_A2_c_267_n N_A1_c_339_n 0.0128971f $X=5.135 $Y=1.595 $X2=0 $Y2=0
cc_215 N_A2_c_254_n N_A1_c_340_n 0.0383927f $X=5.325 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A2_c_267_n N_A1_c_340_n 0.012329f $X=5.135 $Y=1.595 $X2=0 $Y2=0
cc_217 A2 N_A1_c_340_n 0.00225673f $X=5.18 $Y=1.445 $X2=0 $Y2=0
cc_218 N_A2_c_253_n N_A1_c_336_n 0.0307767f $X=5.3 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A2_c_251_n A1 2.47222e-19 $X=3.915 $Y=1.41 $X2=0 $Y2=0
cc_220 N_A2_c_254_n A1 0.00178471f $X=5.325 $Y=1.41 $X2=0 $Y2=0
cc_221 N_A2_c_267_n A1 0.0308222f $X=5.135 $Y=1.595 $X2=0 $Y2=0
cc_222 N_A2_c_256_n A1 0.0225433f $X=4.057 $Y=1.142 $X2=0 $Y2=0
cc_223 N_A2_c_257_n A1 0.0197242f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A2_c_251_n N_A1_c_338_n 0.0254638f $X=3.915 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A2_c_254_n N_A1_c_338_n 0.0307767f $X=5.325 $Y=1.41 $X2=0 $Y2=0
cc_226 N_A2_c_255_n N_A1_c_338_n 0.00318001f $X=4.057 $Y=1.51 $X2=0 $Y2=0
cc_227 N_A2_c_267_n N_A1_c_338_n 0.00618756f $X=5.135 $Y=1.595 $X2=0 $Y2=0
cc_228 N_A2_c_256_n N_A1_c_338_n 0.00186335f $X=4.057 $Y=1.142 $X2=0 $Y2=0
cc_229 N_A2_c_257_n N_A1_c_338_n 0.00117008f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_230 A2 N_A1_c_338_n 0.00278977f $X=5.18 $Y=1.445 $X2=0 $Y2=0
cc_231 N_A2_c_255_n N_VPWR_M1004_d 2.8034e-19 $X=4.057 $Y=1.51 $X2=0 $Y2=0
cc_232 N_A2_c_267_n N_VPWR_M1004_d 0.00212796f $X=5.135 $Y=1.595 $X2=0 $Y2=0
cc_233 N_A2_c_297_p N_VPWR_M1004_d 0.00116838f $X=4.17 $Y=1.595 $X2=0 $Y2=0
cc_234 N_A2_c_267_n N_VPWR_M1015_s 0.00644314f $X=5.135 $Y=1.595 $X2=0 $Y2=0
cc_235 A2 N_VPWR_M1015_s 3.02274e-19 $X=5.18 $Y=1.445 $X2=0 $Y2=0
cc_236 N_A2_c_300_p N_VPWR_M1015_s 4.58089e-19 $X=5.285 $Y=1.51 $X2=0 $Y2=0
cc_237 N_A2_c_251_n N_VPWR_c_387_n 0.0104236f $X=3.915 $Y=1.41 $X2=0 $Y2=0
cc_238 N_A2_c_251_n N_VPWR_c_388_n 0.0031857f $X=3.915 $Y=1.41 $X2=0 $Y2=0
cc_239 N_A2_c_254_n N_VPWR_c_389_n 0.0105364f $X=5.325 $Y=1.41 $X2=0 $Y2=0
cc_240 N_A2_c_254_n N_VPWR_c_392_n 0.00463375f $X=5.325 $Y=1.41 $X2=0 $Y2=0
cc_241 N_A2_c_251_n N_VPWR_c_381_n 0.0039001f $X=3.915 $Y=1.41 $X2=0 $Y2=0
cc_242 N_A2_c_254_n N_VPWR_c_381_n 0.00642292f $X=5.325 $Y=1.41 $X2=0 $Y2=0
cc_243 N_A2_c_267_n N_A_523_297#_M1001_d 0.00348955f $X=5.135 $Y=1.595 $X2=0
+ $Y2=0
cc_244 N_A2_c_251_n N_A_523_297#_c_535_n 0.00141217f $X=3.915 $Y=1.41 $X2=0
+ $Y2=0
cc_245 N_A2_c_251_n N_A_523_297#_c_531_n 0.00463826f $X=3.915 $Y=1.41 $X2=0
+ $Y2=0
cc_246 N_A2_c_255_n N_A_523_297#_c_531_n 0.00449863f $X=4.057 $Y=1.51 $X2=0
+ $Y2=0
cc_247 N_A2_c_297_p N_A_523_297#_c_531_n 0.0128305f $X=4.17 $Y=1.595 $X2=0 $Y2=0
cc_248 N_A2_c_256_n N_A_523_297#_c_531_n 0.00336061f $X=4.057 $Y=1.142 $X2=0
+ $Y2=0
cc_249 N_A2_c_251_n N_A_523_297#_c_551_n 0.0052858f $X=3.915 $Y=1.41 $X2=0 $Y2=0
cc_250 N_A2_c_251_n N_A_523_297#_c_552_n 0.0129464f $X=3.915 $Y=1.41 $X2=0 $Y2=0
cc_251 N_A2_c_267_n N_A_523_297#_c_552_n 0.0171783f $X=5.135 $Y=1.595 $X2=0
+ $Y2=0
cc_252 N_A2_c_297_p N_A_523_297#_c_552_n 0.0127265f $X=4.17 $Y=1.595 $X2=0 $Y2=0
cc_253 N_A2_c_256_n N_A_523_297#_c_552_n 0.00391327f $X=4.057 $Y=1.142 $X2=0
+ $Y2=0
cc_254 N_A2_c_254_n N_A_523_297#_c_556_n 0.0168236f $X=5.325 $Y=1.41 $X2=0 $Y2=0
cc_255 N_A2_c_267_n N_A_523_297#_c_556_n 0.0218994f $X=5.135 $Y=1.595 $X2=0
+ $Y2=0
cc_256 N_A2_c_257_n N_A_523_297#_c_556_n 0.00215221f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_257 N_A2_c_300_p N_A_523_297#_c_556_n 0.0164008f $X=5.285 $Y=1.51 $X2=0 $Y2=0
cc_258 N_A2_c_254_n N_A_523_297#_c_532_n 0.00761692f $X=5.325 $Y=1.41 $X2=0
+ $Y2=0
cc_259 A2 N_A_523_297#_c_532_n 0.0029503f $X=5.18 $Y=1.445 $X2=0 $Y2=0
cc_260 N_A2_c_267_n N_A_523_297#_c_562_n 0.0137194f $X=5.135 $Y=1.595 $X2=0
+ $Y2=0
cc_261 N_A2_c_254_n N_A_523_297#_c_533_n 0.0132625f $X=5.325 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A2_c_257_n N_A_523_297#_c_533_n 0.00240172f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_263 N_A2_c_252_n N_VGND_c_599_n 0.00921343f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A2_c_253_n N_VGND_c_601_n 0.0184132f $X=5.3 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A2_c_254_n N_VGND_c_601_n 0.00248023f $X=5.325 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A2_c_257_n N_VGND_c_601_n 0.0126389f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_267 N_A2_c_252_n N_VGND_c_605_n 0.00343403f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A2_c_253_n N_VGND_c_605_n 0.00585385f $X=5.3 $Y=0.995 $X2=0 $Y2=0
cc_269 N_A2_c_252_n N_VGND_c_609_n 0.00410952f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_270 N_A2_c_253_n N_VGND_c_609_n 0.0117951f $X=5.3 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A1_c_339_n N_VPWR_c_387_n 0.00658869f $X=4.385 $Y=1.41 $X2=0 $Y2=0
cc_272 N_A1_c_340_n N_VPWR_c_387_n 4.81844e-19 $X=4.855 $Y=1.41 $X2=0 $Y2=0
cc_273 N_A1_c_339_n N_VPWR_c_389_n 5.3082e-19 $X=4.385 $Y=1.41 $X2=0 $Y2=0
cc_274 N_A1_c_340_n N_VPWR_c_389_n 0.00935681f $X=4.855 $Y=1.41 $X2=0 $Y2=0
cc_275 N_A1_c_339_n N_VPWR_c_390_n 0.00463375f $X=4.385 $Y=1.41 $X2=0 $Y2=0
cc_276 N_A1_c_340_n N_VPWR_c_390_n 0.0031857f $X=4.855 $Y=1.41 $X2=0 $Y2=0
cc_277 N_A1_c_339_n N_VPWR_c_381_n 0.00530746f $X=4.385 $Y=1.41 $X2=0 $Y2=0
cc_278 N_A1_c_340_n N_VPWR_c_381_n 0.00382788f $X=4.855 $Y=1.41 $X2=0 $Y2=0
cc_279 N_A1_c_339_n N_A_523_297#_c_552_n 0.0115517f $X=4.385 $Y=1.41 $X2=0 $Y2=0
cc_280 N_A1_c_340_n N_A_523_297#_c_556_n 0.0111556f $X=4.855 $Y=1.41 $X2=0 $Y2=0
cc_281 N_A1_c_335_n N_VGND_c_599_n 0.00198574f $X=4.36 $Y=0.995 $X2=0 $Y2=0
cc_282 N_A1_c_335_n N_VGND_c_605_n 0.00430182f $X=4.36 $Y=0.995 $X2=0 $Y2=0
cc_283 N_A1_c_336_n N_VGND_c_605_n 0.00585385f $X=4.88 $Y=0.995 $X2=0 $Y2=0
cc_284 N_A1_c_335_n N_VGND_c_609_n 0.00626756f $X=4.36 $Y=0.995 $X2=0 $Y2=0
cc_285 N_A1_c_336_n N_VGND_c_609_n 0.0110915f $X=4.88 $Y=0.995 $X2=0 $Y2=0
cc_286 N_VPWR_c_381_n N_X_M1003_s 0.00737013f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_287 N_VPWR_c_381_n N_X_M1018_s 0.00522767f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_288 N_VPWR_c_383_n N_X_c_508_n 0.0146286f $X=0.28 $Y=2.02 $X2=0 $Y2=0
cc_289 N_VPWR_c_384_n N_X_c_508_n 0.0178565f $X=1.24 $Y=2.02 $X2=0 $Y2=0
cc_290 N_VPWR_c_391_n N_X_c_508_n 0.00405967f $X=1.025 $Y=2.72 $X2=0 $Y2=0
cc_291 N_VPWR_c_381_n N_X_c_508_n 0.00540609f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_292 N_VPWR_M1012_d N_X_c_492_n 0.00393627f $X=1.09 $Y=1.485 $X2=0 $Y2=0
cc_293 N_VPWR_c_384_n N_X_c_492_n 0.0200928f $X=1.24 $Y=2.02 $X2=0 $Y2=0
cc_294 N_VPWR_c_384_n N_X_c_499_n 0.0152212f $X=1.24 $Y=2.02 $X2=0 $Y2=0
cc_295 N_VPWR_c_385_n N_X_c_499_n 0.00531705f $X=2.065 $Y=2.72 $X2=0 $Y2=0
cc_296 N_VPWR_c_381_n N_X_c_499_n 0.00789534f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_297 N_VPWR_M1003_d X 0.0160803f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_298 N_VPWR_c_383_n X 0.0207391f $X=0.28 $Y=2.02 $X2=0 $Y2=0
cc_299 N_VPWR_c_381_n N_A_523_297#_M1011_d 0.00357188f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_300 N_VPWR_c_381_n N_A_523_297#_M1014_d 0.00260471f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_301 N_VPWR_c_381_n N_A_523_297#_M1001_d 0.00283933f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_302 N_VPWR_c_381_n N_A_523_297#_M1013_s 0.00387284f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_303 N_VPWR_c_386_n N_A_523_297#_c_534_n 0.026941f $X=2.2 $Y=1.68 $X2=0 $Y2=0
cc_304 N_VPWR_c_387_n N_A_523_297#_c_535_n 0.0141783f $X=4.15 $Y=2.36 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_388_n N_A_523_297#_c_535_n 0.053582f $X=3.935 $Y=2.72 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_381_n N_A_523_297#_c_535_n 0.0335752f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_386_n N_A_523_297#_c_575_n 0.00851268f $X=2.2 $Y=1.68 $X2=0
+ $Y2=0
cc_308 N_VPWR_c_388_n N_A_523_297#_c_575_n 0.0119545f $X=3.935 $Y=2.72 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_381_n N_A_523_297#_c_575_n 0.006547f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_310 N_VPWR_c_387_n N_A_523_297#_c_551_n 0.00146273f $X=4.15 $Y=2.36 $X2=0
+ $Y2=0
cc_311 N_VPWR_M1004_d N_A_523_297#_c_552_n 0.00401401f $X=4.005 $Y=1.485 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_387_n N_A_523_297#_c_552_n 0.0137903f $X=4.15 $Y=2.36 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_388_n N_A_523_297#_c_552_n 0.00204483f $X=3.935 $Y=2.72 $X2=0
+ $Y2=0
cc_314 N_VPWR_c_390_n N_A_523_297#_c_552_n 0.00275152f $X=4.875 $Y=2.72 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_381_n N_A_523_297#_c_552_n 0.0108873f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_316 N_VPWR_c_387_n N_A_523_297#_c_584_n 0.0116296f $X=4.15 $Y=2.36 $X2=0
+ $Y2=0
cc_317 N_VPWR_c_389_n N_A_523_297#_c_584_n 0.0141845f $X=5.09 $Y=2.36 $X2=0
+ $Y2=0
cc_318 N_VPWR_c_390_n N_A_523_297#_c_584_n 0.0117273f $X=4.875 $Y=2.72 $X2=0
+ $Y2=0
cc_319 N_VPWR_c_381_n N_A_523_297#_c_584_n 0.00645298f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_320 N_VPWR_M1015_s N_A_523_297#_c_556_n 0.0040301f $X=4.945 $Y=1.485 $X2=0
+ $Y2=0
cc_321 N_VPWR_c_389_n N_A_523_297#_c_556_n 0.0137903f $X=5.09 $Y=2.36 $X2=0
+ $Y2=0
cc_322 N_VPWR_c_390_n N_A_523_297#_c_556_n 0.00204483f $X=4.875 $Y=2.72 $X2=0
+ $Y2=0
cc_323 N_VPWR_c_392_n N_A_523_297#_c_556_n 0.00360937f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_324 N_VPWR_c_381_n N_A_523_297#_c_556_n 0.0123898f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_325 N_VPWR_c_389_n N_A_523_297#_c_533_n 0.00650951f $X=5.09 $Y=2.36 $X2=0
+ $Y2=0
cc_326 N_VPWR_c_392_n N_A_523_297#_c_533_n 0.015862f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_327 N_VPWR_c_381_n N_A_523_297#_c_533_n 0.0121599f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_328 N_X_c_485_n N_VGND_M1002_s 0.0108744f $X=0.68 $Y=0.7 $X2=-0.19 $Y2=-0.24
cc_329 X N_VGND_M1002_s 0.00485264f $X=0.145 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_330 N_X_c_486_n N_VGND_M1005_s 0.00435335f $X=1.72 $Y=0.7 $X2=0 $Y2=0
cc_331 N_X_c_485_n N_VGND_c_598_n 0.0200973f $X=0.68 $Y=0.7 $X2=0 $Y2=0
cc_332 N_X_c_485_n N_VGND_c_604_n 0.00399269f $X=0.68 $Y=0.7 $X2=0 $Y2=0
cc_333 N_X_c_486_n N_VGND_c_604_n 0.0057005f $X=1.72 $Y=0.7 $X2=0 $Y2=0
cc_334 N_X_c_486_n N_VGND_c_606_n 0.0196989f $X=1.72 $Y=0.7 $X2=0 $Y2=0
cc_335 N_X_c_486_n N_VGND_c_607_n 0.00768849f $X=1.72 $Y=0.7 $X2=0 $Y2=0
cc_336 N_X_M1002_d N_VGND_c_609_n 0.00375772f $X=0.57 $Y=0.235 $X2=0 $Y2=0
cc_337 N_X_M1008_d N_VGND_c_609_n 0.00375928f $X=1.53 $Y=0.235 $X2=0 $Y2=0
cc_338 N_X_c_485_n N_VGND_c_609_n 0.00811464f $X=0.68 $Y=0.7 $X2=0 $Y2=0
cc_339 N_X_c_486_n N_VGND_c_609_n 0.0241206f $X=1.72 $Y=0.7 $X2=0 $Y2=0
cc_340 N_A_523_297#_c_532_n N_VGND_c_601_n 0.00456504f $X=5.695 $Y=1.63 $X2=0
+ $Y2=0
cc_341 N_VGND_c_609_n A_801_47# 0.00341244f $X=5.75 $Y=0 $X2=-0.19 $Y2=-0.24
cc_342 N_VGND_c_609_n A_991_47# 0.0115413f $X=5.75 $Y=0 $X2=-0.19 $Y2=-0.24
