* File: sky130_fd_sc_hdll__einvp_1.spice
* Created: Wed Sep  2 08:31:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__einvp_1.pex.spice"
.subckt sky130_fd_sc_hdll__einvp_1  VNB VPB TE A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE	TE
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_TE_M1003_g N_A_27_47#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1005 A_204_47# N_TE_M1005_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.352625 AS=0.11785 PD=1.735 PS=1.18458 NRD=89.988 NRS=9.228 M=1 R=4.33333
+ SA=75000.5 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1002 N_Z_M1002_d N_A_M1002_g A_204_47# VNB NSHORT L=0.15 W=0.65 AD=0.208
+ AS=0.352625 PD=1.94 PS=1.735 NRD=8.304 NRS=89.988 M=1 R=4.33333 SA=75001.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_TE_M1001_g N_A_27_47#_M1001_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.250137 AS=0.1134 PD=1.12099 PS=1.38 NRD=7.0329 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90001.9 A=0.0756 P=1.2 MULT=1
MM1000 A_332_297# N_A_27_47#_M1000_g N_VPWR_M1001_d VPB PHIGHVT L=0.18 W=1
+ AD=0.2275 AS=0.595563 PD=1.455 PS=2.66901 NRD=33.9628 NRS=19.7 M=1 R=5.55556
+ SA=90000.9 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1004 N_Z_M1004_d N_A_M1004_g A_332_297# VPB PHIGHVT L=0.18 W=1 AD=0.28
+ AS=0.2275 PD=2.56 PS=1.455 NRD=2.9353 NRS=33.9628 M=1 R=5.55556 SA=90001.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.0397 P=9.49
pX7_noxref noxref_11 Z Z PROBETYPE=1
pX8_noxref noxref_12 Z Z PROBETYPE=1
*
.include "sky130_fd_sc_hdll__einvp_1.pxi.spice"
*
.ends
*
*
