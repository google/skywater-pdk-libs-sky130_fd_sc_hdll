* File: sky130_fd_sc_hdll__a221oi_1.pex.spice
* Created: Wed Sep  2 08:18:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A221OI_1%C1 1 3 4 6 7 12
c29 7 0 1.426e-19 $X=0.23 $Y=1.19
r30 12 13 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r31 10 12 32.4423 $w=3.64e-07 $l=2.45e-07 $layer=POLY_cond $X=0.25 $Y=1.202
+ $X2=0.495 $Y2=1.202
r32 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r33 4 13 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r34 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r35 1 12 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r36 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_1%B2 1 3 4 6 7 11 13
c26 1 0 2.70309e-19 $X=0.965 $Y=1.41
r27 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r28 7 11 10.0346 $w=2.08e-07 $l=1.9e-07 $layer=LI1_cond $X=0.75 $Y=1.18 $X2=0.94
+ $Y2=1.18
r29 7 13 2.64069 $w=2.08e-07 $l=5e-08 $layer=LI1_cond $X=0.75 $Y=1.18 $X2=0.7
+ $Y2=1.18
r30 4 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.05 $Y=0.995
+ $X2=0.965 $Y2=1.16
r31 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.05 $Y=0.995 $X2=1.05
+ $Y2=0.56
r32 1 10 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.16
r33 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_1%B1 1 3 4 6 7 8 14 21
r37 13 21 6.33766 $w=2.08e-07 $l=1.2e-07 $layer=LI1_cond $X=1.49 $Y=1.18
+ $X2=1.61 $Y2=1.18
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.49
+ $Y=1.16 $X2=1.49 $Y2=1.16
r39 8 14 2.64069 $w=2.08e-07 $l=5e-08 $layer=LI1_cond $X=1.62 $Y=1.18 $X2=1.67
+ $Y2=1.18
r40 8 21 0.528139 $w=2.08e-07 $l=1e-08 $layer=LI1_cond $X=1.62 $Y=1.18 $X2=1.61
+ $Y2=1.18
r41 7 14 8.94137 $w=2.88e-07 $l=2.25e-07 $layer=LI1_cond $X=1.67 $Y=0.85
+ $X2=1.67 $Y2=1.075
r42 4 12 47.0331 $w=3.15e-07 $l=2.83725e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.507 $Y2=1.16
r43 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r44 1 12 38.5363 $w=3.15e-07 $l=2.07918e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.507 $Y2=1.16
r45 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995 $X2=1.41
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_1%A1 1 3 4 6 7 8 13
c35 8 0 6.98876e-20 $X=2.07 $Y=0.85
r36 13 19 2.59521 $w=4.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.205 $Y=1.16
+ $X2=2.205 $Y2=1.075
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=1.16 $X2=2.26 $Y2=1.16
r38 8 19 7.1041 $w=3.63e-07 $l=2.25e-07 $layer=LI1_cond $X=2.167 $Y=0.85
+ $X2=2.167 $Y2=1.075
r39 7 13 0.785757 $w=4.38e-07 $l=3e-08 $layer=LI1_cond $X=2.205 $Y=1.19
+ $X2=2.205 $Y2=1.16
r40 4 12 38.8967 $w=3.59e-07 $l=2.18746e-07 $layer=POLY_cond $X=2.45 $Y=0.995
+ $X2=2.325 $Y2=1.16
r41 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.45 $Y=0.995 $X2=2.45
+ $Y2=0.56
r42 1 12 45.5371 $w=3.59e-07 $l=2.95804e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.325 $Y2=1.16
r43 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_1%A2 1 3 4 6 7 15
c31 1 0 6.98876e-20 $X=2.955 $Y=1.41
r32 7 15 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=1.16
+ $X2=2.955 $Y2=1.16
r33 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.87
+ $Y=1.16 $X2=2.87 $Y2=1.16
r34 4 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.98 $Y=0.995
+ $X2=2.895 $Y2=1.16
r35 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.98 $Y=0.995 $X2=2.98
+ $Y2=0.56
r36 1 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.955 $Y=1.41
+ $X2=2.895 $Y2=1.16
r37 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.955 $Y=1.41
+ $X2=2.955 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_1%Y 1 2 3 4 15 19 21 22 24 27 28 33 36 37
+ 38 39 40 41 42 43 49 50 52
c110 52 0 1.53436e-19 $X=3.355 $Y=0.85
r111 49 52 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=3.395 $Y=0.825
+ $X2=3.395 $Y2=0.85
r112 43 50 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.395 $Y=1.58
+ $X2=3.395 $Y2=1.495
r113 43 50 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=3.395 $Y=1.47
+ $X2=3.395 $Y2=1.495
r114 42 43 11.5244 $w=2.78e-07 $l=2.8e-07 $layer=LI1_cond $X=3.395 $Y=1.19
+ $X2=3.395 $Y2=1.47
r115 41 49 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.395 $Y=0.74
+ $X2=3.395 $Y2=0.825
r116 41 42 12.7592 $w=2.78e-07 $l=3.1e-07 $layer=LI1_cond $X=3.395 $Y=0.88
+ $X2=3.395 $Y2=1.19
r117 41 52 1.23476 $w=2.78e-07 $l=3e-08 $layer=LI1_cond $X=3.395 $Y=0.88
+ $X2=3.395 $Y2=0.85
r118 39 40 7.92208 $w=2.08e-07 $l=1.5e-07 $layer=LI1_cond $X=2.3 $Y=1.56
+ $X2=2.45 $Y2=1.56
r119 37 41 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.255 $Y=0.74
+ $X2=3.395 $Y2=0.74
r120 37 38 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.255 $Y=0.74
+ $X2=2.78 $Y2=0.74
r121 36 38 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.68 $Y=0.655
+ $X2=2.78 $Y2=0.74
r122 35 36 8.31818 $w=1.98e-07 $l=1.5e-07 $layer=LI1_cond $X=2.68 $Y=0.505
+ $X2=2.68 $Y2=0.655
r123 33 43 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.255 $Y=1.58
+ $X2=3.395 $Y2=1.58
r124 33 40 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=3.255 $Y=1.58
+ $X2=2.45 $Y2=1.58
r125 30 32 23.9708 $w=2.48e-07 $l=5.2e-07 $layer=LI1_cond $X=1.67 $Y=0.38
+ $X2=2.19 $Y2=0.38
r126 28 30 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.335 $Y=0.38
+ $X2=1.67 $Y2=0.38
r127 27 35 6.92652 $w=2.5e-07 $l=1.67705e-07 $layer=LI1_cond $X=2.58 $Y=0.38
+ $X2=2.68 $Y2=0.505
r128 27 32 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=2.58 $Y=0.38
+ $X2=2.19 $Y2=0.38
r129 25 28 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.25 $Y=0.505
+ $X2=1.335 $Y2=0.38
r130 25 26 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.25 $Y=0.505
+ $X2=1.25 $Y2=0.735
r131 24 39 127.545 $w=1.68e-07 $l=1.955e-06 $layer=LI1_cond $X=0.345 $Y=1.54
+ $X2=2.3 $Y2=1.54
r132 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.165 $Y=0.82
+ $X2=1.25 $Y2=0.735
r133 21 22 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.165 $Y=0.82
+ $X2=0.345 $Y2=0.82
r134 17 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.345 $Y2=1.54
r135 17 19 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.26 $Y2=1.65
r136 13 22 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.345 $Y2=0.82
r137 13 15 11.0909 $w=1.73e-07 $l=1.75e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.257 $Y2=0.56
r138 4 19 300 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.65
r139 3 32 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=2.065
+ $Y=0.235 $X2=2.19 $Y2=0.42
r140 2 30 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.42
r141 1 15 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_1%A_117_297# 1 2 9 12 13 15 17
c25 13 0 1.2771e-19 $X=1.56 $Y=2.36
r26 13 17 5.98033 $w=2.08e-07 $l=1.05e-07 $layer=LI1_cond $X=1.56 $Y=2.36
+ $X2=1.455 $Y2=2.36
r27 13 15 5.80952 $w=2.08e-07 $l=1.1e-07 $layer=LI1_cond $X=1.56 $Y=2.36
+ $X2=1.67 $Y2=2.36
r28 12 17 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.815 $Y=2.38
+ $X2=1.455 $Y2=2.38
r29 7 12 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=0.665 $Y=2.295
+ $X2=0.815 $Y2=2.38
r30 7 9 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=0.665 $Y=2.295
+ $X2=0.665 $Y2=1.96
r31 2 15 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
r32 1 9 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_1%A_211_297# 1 2 7 9 11 13 18 19
r29 16 18 5.59382 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.2 $Y=1.96 $X2=1.34
+ $Y2=1.96
r30 11 21 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=2.7 $Y=2.045 $X2=2.7
+ $Y2=1.94
r31 11 13 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=2.7 $Y=2.045
+ $X2=2.7 $Y2=2.3
r32 9 21 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.575 $Y=1.94 $X2=2.7
+ $Y2=1.94
r33 9 19 21.1255 $w=2.08e-07 $l=4e-07 $layer=LI1_cond $X=2.575 $Y=1.94 $X2=2.175
+ $Y2=1.94
r34 7 19 6.09095 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.05 $Y=1.92
+ $X2=2.175 $Y2=1.92
r35 7 18 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=2.05 $Y=1.92 $X2=1.34
+ $Y2=1.92
r36 2 21 600 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=1.485 $X2=2.66 $Y2=1.95
r37 2 13 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=1.485 $X2=2.66 $Y2=2.3
r38 1 16 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_1%VPWR 1 2 9 13 16 17 18 20 30 31 34
c50 2 0 1.53436e-19 $X=3.045 $Y=1.485
r51 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r52 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r53 28 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r54 28 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r55 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r56 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=2.72
+ $X2=2.19 $Y2=2.72
r57 25 27 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.355 $Y=2.72
+ $X2=2.99 $Y2=2.72
r58 20 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=2.19 $Y2=2.72
r59 20 22 117.107 $w=1.68e-07 $l=1.795e-06 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=0.23 $Y2=2.72
r60 18 35 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r61 18 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r62 16 27 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.045 $Y=2.72
+ $X2=2.99 $Y2=2.72
r63 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.045 $Y=2.72
+ $X2=3.21 $Y2=2.72
r64 15 30 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.375 $Y=2.72
+ $X2=3.45 $Y2=2.72
r65 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=2.72
+ $X2=3.21 $Y2=2.72
r66 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=2.635
+ $X2=3.21 $Y2=2.72
r67 11 13 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.21 $Y=2.635
+ $X2=3.21 $Y2=1.96
r68 7 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=2.635 $X2=2.19
+ $Y2=2.72
r69 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.19 $Y=2.635 $X2=2.19
+ $Y2=2.3
r70 2 13 300 $w=1.7e-07 $l=5.51362e-07 $layer=licon1_PDIFF $count=2 $X=3.045
+ $Y=1.485 $X2=3.21 $Y2=1.96
r71 1 9 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=2.065
+ $Y=1.485 $X2=2.19 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_1%VGND 1 2 9 13 16 17 18 20 33 34 37
r49 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r50 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r51 31 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r52 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r53 28 31 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r54 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r55 27 30 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r56 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r57 25 37 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r58 25 27 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.15
+ $Y2=0
r59 20 37 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r60 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r61 18 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r62 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r63 16 30 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=3.03 $Y=0 $X2=2.99
+ $Y2=0
r64 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.03 $Y=0 $X2=3.195
+ $Y2=0
r65 15 33 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.36 $Y=0 $X2=3.45
+ $Y2=0
r66 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.36 $Y=0 $X2=3.195
+ $Y2=0
r67 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.195 $Y=0.085
+ $X2=3.195 $Y2=0
r68 11 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.195 $Y=0.085
+ $X2=3.195 $Y2=0.4
r69 7 37 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r70 7 9 10.7662 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.44
r71 2 13 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.055
+ $Y=0.235 $X2=3.195 $Y2=0.4
r72 1 9 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.44
.ends

