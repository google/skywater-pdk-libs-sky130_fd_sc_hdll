* File: sky130_fd_sc_hdll__a31o_4.spice
* Created: Thu Aug 27 18:55:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a31o_4.pex.spice"
.subckt sky130_fd_sc_hdll__a31o_4  VNB VPB A3 A2 A1 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1016 N_VGND_M1016_d N_A3_M1016_g A_119_47# VNB NSHORT L=0.15 W=0.65 AD=0.2015
+ AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=19.38 M=1 R=4.33333 SA=75000.2 SB=75006
+ A=0.0975 P=1.6 MULT=1
MM1001 A_119_47# N_A2_M1001_g A_213_47# VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.08775 PD=0.97 PS=0.92 NRD=19.38 NRS=14.76 M=1 R=4.33333 SA=75000.7
+ SB=75005.5 A=0.0975 P=1.6 MULT=1
MM1005 A_213_47# N_A1_M1005_g N_A_297_47#_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=14.76 NRS=8.304 M=1 R=4.33333
+ SA=75001.1 SB=75005.1 A=0.0975 P=1.6 MULT=1
MM1017 A_401_47# N_A1_M1017_g N_A_297_47#_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=19.38 NRS=8.304 M=1 R=4.33333
+ SA=75001.6 SB=75004.6 A=0.0975 P=1.6 MULT=1
MM1014 A_495_47# N_A2_M1014_g A_401_47# VNB NSHORT L=0.15 W=0.65 AD=0.10725
+ AS=0.104 PD=0.98 PS=0.97 NRD=20.304 NRS=19.38 M=1 R=4.33333 SA=75002.1
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1019_d N_A3_M1019_g A_495_47# VNB NSHORT L=0.15 W=0.65 AD=0.1235
+ AS=0.10725 PD=1.03 PS=0.98 NRD=15.684 NRS=20.304 M=1 R=4.33333 SA=75002.6
+ SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1019_d N_B1_M1012_g N_A_297_47#_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.104 PD=1.03 PS=0.97 NRD=2.76 NRS=8.304 M=1 R=4.33333 SA=75003.1
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1021_d N_B1_M1021_g N_A_297_47#_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.28925 AS=0.104 PD=1.54 PS=0.97 NRD=23.076 NRS=0 M=1 R=4.33333 SA=75003.6
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1021_d N_A_297_47#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.28925 AS=0.104 PD=1.54 PS=0.97 NRD=23.076 NRS=0 M=1 R=4.33333 SA=75004.6
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A_297_47#_M1008_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75005.1
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1008_d N_A_297_47#_M1010_g N_X_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75005.6
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1023 N_VGND_M1023_d N_A_297_47#_M1023_g N_X_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.104 PD=1.82 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75006
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_27_297#_M1002_d N_A3_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.6 A=0.18 P=2.36 MULT=1
MM1000 N_A_27_297#_M1000_d N_A2_M1000_g N_VPWR_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1015 N_A_27_297#_M1000_d N_A1_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1022 N_A_27_297#_M1022_d N_A1_M1022_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1011 N_A_27_297#_M1022_d N_A2_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.175 PD=1.29 PS=1.35 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1007 N_A_27_297#_M1007_d N_A3_M1007_g N_VPWR_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=12.7853 NRS=12.7853 M=1 R=5.55556
+ SA=90002.6 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1009 N_A_27_297#_M1007_d N_B1_M1009_g N_A_297_47#_M1009_s VPB PHIGHVT L=0.18
+ W=1 AD=0.175 AS=0.145 PD=1.35 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1018 N_A_27_297#_M1018_d N_B1_M1018_g N_A_297_47#_M1009_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1003 N_X_M1003_d N_A_297_47#_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1006 N_X_M1003_d N_A_297_47#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1013 N_X_M1013_d N_A_297_47#_M1013_g N_VPWR_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1020 N_X_M1013_d N_A_297_47#_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX24_noxref VNB VPB NWDIODE A=11.6844 P=17.77
*
.include "sky130_fd_sc_hdll__a31o_4.pxi.spice"
*
.ends
*
*
