* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__isobufsrc_8 A SLEEP VGND VNB VPB VPWR X
X0 a_345_297# a_117_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 X SLEEP a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_117_297# a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_345_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 VPWR a_117_297# a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 VGND a_117_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_345_297# a_117_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_345_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 a_117_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND a_117_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 X SLEEP a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 VGND a_117_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND a_117_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_117_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 VPWR a_117_297# a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 X a_117_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 X a_117_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 X SLEEP a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 VPWR a_117_297# a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 a_345_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X26 X a_117_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 a_345_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 X a_117_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 X SLEEP a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X32 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 a_345_297# a_117_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X34 VGND A a_117_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 a_345_297# a_117_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
