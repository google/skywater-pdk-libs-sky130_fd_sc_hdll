* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
M1000 VPWR A a_614_297# VPB phighvt w=420000u l=180000u
+  ad=8.59325e+11p pd=7.99e+06u as=1.281e+11p ps=1.45e+06u
M1001 VGND C_N a_27_410# VNB nshort w=420000u l=150000u
+  ad=8.121e+11p pd=8.33e+06u as=1.302e+11p ps=1.46e+06u
M1002 a_336_413# a_216_93# VGND VNB nshort w=420000u l=150000u
+  ad=2.814e+11p pd=3.02e+06u as=0p ps=0u
M1003 a_216_93# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1004 VPWR a_336_413# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1005 X a_336_413# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_532_297# a_27_410# a_426_413# VPB phighvt w=420000u l=180000u
+  ad=9.66e+10p pd=1.3e+06u as=2.514e+11p ps=2.7e+06u
M1007 VGND A a_336_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_426_413# a_216_93# a_336_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1009 a_614_297# B a_532_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR C_N a_27_410# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1011 a_216_93# D_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
M1012 a_336_413# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_336_413# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1014 X a_336_413# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_27_410# a_336_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
