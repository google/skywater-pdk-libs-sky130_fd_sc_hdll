* File: sky130_fd_sc_hdll__xnor3_1.pex.spice
* Created: Thu Aug 27 19:29:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__XNOR3_1%A_83_21# 1 2 7 9 10 12 16 19 20 21 22 23
+ 25 27 29 30 32 34 36 38 39
c99 38 0 4.99043e-20 $X=0.635 $Y=1.33
r100 34 39 11.3723 $w=1.98e-07 $l=2e-07 $layer=LI1_cond $X=2.37 $Y=0.355
+ $X2=2.17 $Y2=0.355
r101 34 36 6.65455 $w=1.98e-07 $l=1.2e-07 $layer=LI1_cond $X=2.37 $Y=0.355
+ $X2=2.49 $Y2=0.355
r102 30 32 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=1.32 $Y=2.32
+ $X2=2.415 $Y2=2.32
r103 29 39 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=1.205 $Y=0.34
+ $X2=2.17 $Y2=0.34
r104 27 30 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.21 $Y=2.235
+ $X2=1.32 $Y2=2.32
r105 26 27 9.95292 $w=2.18e-07 $l=1.9e-07 $layer=LI1_cond $X=1.21 $Y=2.045
+ $X2=1.21 $Y2=2.235
r106 24 29 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.095 $Y=0.425
+ $X2=1.205 $Y2=0.34
r107 24 25 14.1436 $w=2.18e-07 $l=2.7e-07 $layer=LI1_cond $X=1.095 $Y=0.425
+ $X2=1.095 $Y2=0.695
r108 22 26 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.1 $Y=1.96
+ $X2=1.21 $Y2=2.045
r109 22 23 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.1 $Y=1.96
+ $X2=0.755 $Y2=1.96
r110 20 25 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.985 $Y=0.78
+ $X2=1.095 $Y2=0.695
r111 20 21 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.985 $Y=0.78
+ $X2=0.755 $Y2=0.78
r112 19 23 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.645 $Y=1.875
+ $X2=0.755 $Y2=1.96
r113 19 38 28.5492 $w=2.18e-07 $l=5.45e-07 $layer=LI1_cond $X=0.645 $Y=1.875
+ $X2=0.645 $Y2=1.33
r114 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.16 $X2=0.6 $Y2=1.16
r115 14 38 5.86323 $w=2.38e-07 $l=1.2e-07 $layer=LI1_cond $X=0.635 $Y=1.21
+ $X2=0.635 $Y2=1.33
r116 14 16 2.40092 $w=2.38e-07 $l=5e-08 $layer=LI1_cond $X=0.635 $Y=1.21
+ $X2=0.635 $Y2=1.16
r117 13 21 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=0.635 $Y=0.865
+ $X2=0.755 $Y2=0.78
r118 13 16 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=0.635 $Y=0.865
+ $X2=0.635 $Y2=1.16
r119 10 17 46.6797 $w=3.23e-07 $l=2.8592e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.592 $Y2=1.16
r120 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r121 7 17 38.5615 $w=3.23e-07 $l=2.09893e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.592 $Y2=1.16
r122 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=0.56
r123 2 32 600 $w=1.7e-07 $l=7.64068e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.625 $X2=2.415 $Y2=2.32
r124 1 36 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.345
+ $Y=0.245 $X2=2.49 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_1%C 1 3 7 8 10 11 13 15 18 19
c60 1 0 1.70967e-19 $X=1.055 $Y=0.995
r61 19 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.015
+ $Y=1.16 $X2=2.015 $Y2=1.16
r62 18 22 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=2.08 $Y=1.16
+ $X2=2.015 $Y2=1.16
r63 14 22 146.009 $w=3.3e-07 $l=8.35e-07 $layer=POLY_cond $X=1.18 $Y=1.16
+ $X2=2.015 $Y2=1.16
r64 14 15 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.18 $Y=1.16
+ $X2=1.08 $Y2=1.202
r65 11 18 39.7875 $w=2.42e-07 $l=1.9182e-07 $layer=POLY_cond $X=2.27 $Y=0.995
+ $X2=2.212 $Y2=1.16
r66 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.27 $Y=0.995
+ $X2=2.27 $Y2=0.565
r67 8 18 80.9439 $w=2.42e-07 $l=4.05685e-07 $layer=POLY_cond $X=2.18 $Y=1.55
+ $X2=2.212 $Y2=1.16
r68 8 10 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=2.18 $Y=1.55 $X2=2.18
+ $Y2=2.045
r69 4 15 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=1.08 $Y=1.41
+ $X2=1.08 $Y2=1.202
r70 4 7 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.08 $Y=1.41 $X2=1.08
+ $Y2=1.805
r71 1 15 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=1.08 $Y2=1.202
r72 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=1.055 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_1%A_226_93# 1 2 7 9 10 12 13 18 20 23 24 28
r70 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.16 $X2=2.69 $Y2=1.16
r71 25 28 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.585 $Y=1.16
+ $X2=2.69 $Y2=1.16
r72 22 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.585 $Y=1.325
+ $X2=2.585 $Y2=1.16
r73 22 23 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.585 $Y=1.325
+ $X2=2.585 $Y2=1.535
r74 21 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.545 $Y=1.62
+ $X2=1.46 $Y2=1.62
r75 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.5 $Y=1.62
+ $X2=2.585 $Y2=1.535
r76 20 21 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=2.5 $Y=1.62
+ $X2=1.545 $Y2=1.62
r77 16 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.46 $Y=1.535
+ $X2=1.46 $Y2=1.62
r78 16 18 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.46 $Y=1.535
+ $X2=1.46 $Y2=0.76
r79 13 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.375 $Y=1.62
+ $X2=1.46 $Y2=1.62
r80 13 15 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=1.375 $Y=1.62 $X2=1.315
+ $Y2=1.62
r81 10 29 38.578 $w=2.95e-07 $l=1.86145e-07 $layer=POLY_cond $X=2.76 $Y=0.995
+ $X2=2.715 $Y2=1.16
r82 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.76 $Y=0.995
+ $X2=2.76 $Y2=0.565
r83 7 29 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=2.715 $Y=1.41
+ $X2=2.715 $Y2=1.16
r84 7 9 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=2.715 $Y=1.41
+ $X2=2.715 $Y2=1.905
r85 2 15 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.17
+ $Y=1.485 $X2=1.315 $Y2=1.62
r86 1 18 182 $w=1.7e-07 $l=4.54148e-07 $layer=licon1_NDIFF $count=1 $X=1.13
+ $Y=0.465 $X2=1.46 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_1%A_783_297# 1 2 7 9 12 15 16 18 21 22 23 27
+ 35 37 38 39 40 47 49 50 55 57 60
c181 55 0 1.24749e-19 $X=7.24 $Y=1.11
c182 27 0 1.36535e-19 $X=4.22 $Y=1.58
r183 55 58 37.8858 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=7.262 $Y=1.11
+ $X2=7.262 $Y2=1.275
r184 55 57 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=7.262 $Y=1.11
+ $X2=7.262 $Y2=0.945
r185 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.24
+ $Y=1.11 $X2=7.24 $Y2=1.11
r186 50 56 11.8358 $w=2.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.17 $Y=0.85
+ $X2=7.17 $Y2=1.11
r187 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.12 $Y=0.85
+ $X2=7.12 $Y2=0.85
r188 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.64 $Y=0.85
+ $X2=5.64 $Y2=0.85
r189 42 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.16 $Y=0.85
+ $X2=4.16 $Y2=0.85
r190 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.785 $Y=0.85
+ $X2=5.64 $Y2=0.85
r191 39 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.975 $Y=0.85
+ $X2=7.12 $Y2=0.85
r192 39 40 1.47277 $w=1.4e-07 $l=1.19e-06 $layer=MET1_cond $X=6.975 $Y=0.85
+ $X2=5.785 $Y2=0.85
r193 38 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.305 $Y=0.85
+ $X2=4.16 $Y2=0.85
r194 37 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.495 $Y=0.85
+ $X2=5.64 $Y2=0.85
r195 37 38 1.47277 $w=1.4e-07 $l=1.19e-06 $layer=MET1_cond $X=5.495 $Y=0.85
+ $X2=4.305 $Y2=0.85
r196 35 47 7.65801 $w=2.08e-07 $l=1.45e-07 $layer=LI1_cond $X=5.62 $Y=0.995
+ $X2=5.62 $Y2=0.85
r197 31 35 6.28605 $w=2.73e-07 $l=1.5e-07 $layer=LI1_cond $X=5.47 $Y=1.132
+ $X2=5.62 $Y2=1.132
r198 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.47
+ $Y=1.16 $X2=5.47 $Y2=1.16
r199 28 60 28.0163 $w=2.88e-07 $l=7.05e-07 $layer=LI1_cond $X=4.22 $Y=1.445
+ $X2=4.22 $Y2=0.74
r200 27 28 0.275955 $w=2.9e-07 $l=1.35e-07 $layer=LI1_cond $X=4.22 $Y=1.58
+ $X2=4.22 $Y2=1.445
r201 25 27 6.82929 $w=2.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.06 $Y=1.58
+ $X2=4.22 $Y2=1.58
r202 22 32 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=5.73 $Y=1.16
+ $X2=5.47 $Y2=1.16
r203 22 23 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=5.73 $Y=1.16
+ $X2=5.83 $Y2=1.202
r204 21 57 131.747 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=7.345 $Y=0.535
+ $X2=7.345 $Y2=0.945
r205 16 18 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=7.32 $Y=1.57
+ $X2=7.32 $Y2=2.065
r206 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.32 $Y=1.47 $X2=7.32
+ $Y2=1.57
r207 15 58 64.6575 $w=2e-07 $l=1.95e-07 $layer=POLY_cond $X=7.32 $Y=1.47
+ $X2=7.32 $Y2=1.275
r208 10 23 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=5.855 $Y=0.995
+ $X2=5.83 $Y2=1.202
r209 10 12 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=5.855 $Y=0.995
+ $X2=5.855 $Y2=0.455
r210 7 23 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=5.83 $Y=1.41
+ $X2=5.83 $Y2=1.202
r211 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=5.83 $Y=1.41
+ $X2=5.83 $Y2=1.805
r212 2 25 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.915
+ $Y=1.485 $X2=4.06 $Y2=1.63
r213 1 60 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.145
+ $Y=0.235 $X2=4.28 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_1%B 1 3 6 8 9 13 16 18 19 22 24 25 28 31 33
+ 35 36 40 42 45
c136 42 0 1.94872e-19 $X=7.035 $Y=1.445
r137 38 42 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.845 $Y=1.53
+ $X2=7.12 $Y2=1.53
r138 38 40 3.92798 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=6.845 $Y=1.53
+ $X2=6.735 $Y2=1.53
r139 36 46 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=6.735 $Y=1.16
+ $X2=6.735 $Y2=1.325
r140 36 45 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=6.735 $Y=1.16
+ $X2=6.735 $Y2=0.995
r141 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.71
+ $Y=1.16 $X2=6.71 $Y2=1.16
r142 33 40 3.03526 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=6.735 $Y=1.445
+ $X2=6.735 $Y2=1.53
r143 33 35 14.9294 $w=2.18e-07 $l=2.85e-07 $layer=LI1_cond $X=6.735 $Y=1.445
+ $X2=6.735 $Y2=1.16
r144 31 32 29.1618 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=5.025 $Y=1.16
+ $X2=5.025 $Y2=1.085
r145 26 28 174.919 $w=1.8e-07 $l=4.5e-07 $layer=POLY_cond $X=6.755 $Y=2.415
+ $X2=6.755 $Y2=1.965
r146 25 28 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=6.755 $Y=1.57
+ $X2=6.755 $Y2=1.965
r147 24 25 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=6.755 $Y=1.47 $X2=6.755
+ $Y2=1.57
r148 24 46 48.0787 $w=2e-07 $l=1.45e-07 $layer=POLY_cond $X=6.755 $Y=1.47
+ $X2=6.755 $Y2=1.325
r149 22 45 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.65 $Y=0.565
+ $X2=6.65 $Y2=0.995
r150 18 26 27.2212 $w=1.5e-07 $l=1.67705e-07 $layer=POLY_cond $X=6.655 $Y=2.54
+ $X2=6.755 $Y2=2.415
r151 18 19 784.532 $w=1.5e-07 $l=1.53e-06 $layer=POLY_cond $X=6.655 $Y=2.54
+ $X2=5.125 $Y2=2.54
r152 16 32 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.05 $Y=0.565
+ $X2=5.05 $Y2=1.085
r153 11 19 27.2212 $w=1.5e-07 $l=1.36015e-07 $layer=POLY_cond $X=5.025 $Y=2.455
+ $X2=5.125 $Y2=2.54
r154 11 13 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=5.025 $Y=2.455
+ $X2=5.025 $Y2=1.905
r155 10 31 83.702 $w=2e-07 $l=2.5e-07 $layer=POLY_cond $X=5.025 $Y=1.41
+ $X2=5.025 $Y2=1.16
r156 10 13 192.411 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=5.025 $Y=1.41
+ $X2=5.025 $Y2=1.905
r157 8 31 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=4.925 $Y=1.16
+ $X2=5.025 $Y2=1.16
r158 8 9 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=4.925 $Y=1.16
+ $X2=4.145 $Y2=1.16
r159 4 9 21.6156 $w=2.33e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.07 $Y=1.085
+ $X2=4.145 $Y2=1.16
r160 4 6 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.07 $Y=1.085
+ $X2=4.07 $Y2=0.56
r161 1 4 50.6824 $w=2.33e-07 $l=3.43642e-07 $layer=POLY_cond $X=3.825 $Y=1.322
+ $X2=4.07 $Y2=1.085
r162 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.825 $Y=1.41
+ $X2=3.825 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_1%A 1 3 4 6 7 15
c38 1 0 1.94872e-19 $X=7.875 $Y=1.41
r39 11 15 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=7.77 $Y=1.2 $X2=8.04
+ $Y2=1.2
r40 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.77
+ $Y=1.16 $X2=7.77 $Y2=1.16
r41 7 15 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=8.045 $Y=1.2 $X2=8.04
+ $Y2=1.2
r42 4 10 38.532 $w=3.11e-07 $l=2.07123e-07 $layer=POLY_cond $X=7.9 $Y=0.995
+ $X2=7.805 $Y2=1.16
r43 4 6 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=7.9 $Y=0.995 $X2=7.9
+ $Y2=0.555
r44 1 10 47.2262 $w=3.11e-07 $l=2.82843e-07 $layer=POLY_cond $X=7.875 $Y=1.41
+ $X2=7.805 $Y2=1.16
r45 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.875 $Y=1.41
+ $X2=7.875 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_1%A_901_297# 1 2 3 4 13 15 16 18 21 23 27 28
+ 29 30 36 37 40 43 44
c130 30 0 1.41691e-19 $X=8.575 $Y=1.495
c131 13 0 3.96944e-20 $X=8.66 $Y=1.41
r132 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.63 $Y=0.51
+ $X2=7.63 $Y2=0.51
r133 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.67 $Y=0.51
+ $X2=4.67 $Y2=0.51
r134 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.815 $Y=0.51
+ $X2=4.67 $Y2=0.51
r135 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.485 $Y=0.51
+ $X2=7.63 $Y2=0.51
r136 36 37 3.30445 $w=1.4e-07 $l=2.67e-06 $layer=MET1_cond $X=7.485 $Y=0.51
+ $X2=4.815 $Y2=0.51
r137 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.635
+ $Y=1.16 $X2=8.635 $Y2=1.16
r138 32 34 17.9567 $w=2.31e-07 $l=3.4e-07 $layer=LI1_cond $X=8.63 $Y=0.82
+ $X2=8.63 $Y2=1.16
r139 31 44 8.94137 $w=2.88e-07 $l=2.25e-07 $layer=LI1_cond $X=7.66 $Y=0.735
+ $X2=7.66 $Y2=0.51
r140 29 34 9.58904 $w=2.31e-07 $l=1.90526e-07 $layer=LI1_cond $X=8.575 $Y=1.325
+ $X2=8.63 $Y2=1.16
r141 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.575 $Y=1.325
+ $X2=8.575 $Y2=1.495
r142 28 31 14.5133 $w=1.17e-07 $l=1.8262e-07 $layer=LI1_cond $X=7.805 $Y=0.82
+ $X2=7.66 $Y2=0.735
r143 27 32 2.5345 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=8.49 $Y=0.82 $X2=8.63
+ $Y2=0.82
r144 27 28 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=8.49 $Y=0.82
+ $X2=7.805 $Y2=0.82
r145 23 30 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=8.49 $Y=1.6
+ $X2=8.575 $Y2=1.495
r146 23 25 44.8918 $w=2.08e-07 $l=8.5e-07 $layer=LI1_cond $X=8.49 $Y=1.6
+ $X2=7.64 $Y2=1.6
r147 19 40 3.57235 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.63 $Y=0.595
+ $X2=4.63 $Y2=0.43
r148 19 21 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=4.63 $Y=0.595
+ $X2=4.63 $Y2=1.94
r149 16 35 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=8.685 $Y=0.995
+ $X2=8.66 $Y2=1.16
r150 16 18 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.685 $Y=0.995
+ $X2=8.685 $Y2=0.555
r151 13 35 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=8.66 $Y=1.41
+ $X2=8.66 $Y2=1.16
r152 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.66 $Y=1.41
+ $X2=8.66 $Y2=1.985
r153 4 25 600 $w=1.7e-07 $l=2.42178e-07 $layer=licon1_PDIFF $count=1 $X=7.41
+ $Y=1.645 $X2=7.64 $Y2=1.62
r154 3 21 600 $w=1.7e-07 $l=5.13712e-07 $layer=licon1_PDIFF $count=1 $X=4.505
+ $Y=1.485 $X2=4.63 $Y2=1.94
r155 2 44 182 $w=1.7e-07 $l=4.8775e-07 $layer=licon1_NDIFF $count=1 $X=7.42
+ $Y=0.235 $X2=7.64 $Y2=0.625
r156 1 40 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=4.665
+ $Y=0.245 $X2=4.79 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_1%X 1 2 9 11 13 16
r21 13 20 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=0.225 $Y=1.87
+ $X2=0.225 $Y2=2.3
r22 13 16 10.2897 $w=2.78e-07 $l=2.5e-07 $layer=LI1_cond $X=0.225 $Y=1.87
+ $X2=0.225 $Y2=1.62
r23 11 16 1.64635 $w=2.78e-07 $l=4e-08 $layer=LI1_cond $X=0.225 $Y=1.58
+ $X2=0.225 $Y2=1.62
r24 11 12 5.83872 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=0.225 $Y=1.58
+ $X2=0.225 $Y2=1.44
r25 9 12 39.0058 $w=2.58e-07 $l=8.8e-07 $layer=LI1_cond $X=0.215 $Y=0.56
+ $X2=0.215 $Y2=1.44
r26 2 20 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r27 2 16 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r28 1 9 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_1%VPWR 1 2 3 12 16 18 20 25 40 41 44 47 51
+ 55
c92 3 0 1.41691e-19 $X=7.965 $Y=1.485
r93 53 55 7.89897 $w=5.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.51 $Y=2.54
+ $X2=8.595 $Y2=2.54
r94 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r95 50 53 5.30337 $w=5.28e-07 $l=2.35e-07 $layer=LI1_cond $X=8.275 $Y=2.54
+ $X2=8.51 $Y2=2.54
r96 50 51 14.105 $w=5.28e-07 $l=3.6e-07 $layer=LI1_cond $X=8.275 $Y=2.54
+ $X2=7.915 $Y2=2.54
r97 47 48 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r98 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r99 41 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=8.51 $Y2=2.72
r100 40 55 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.97 $Y=2.72
+ $X2=8.595 $Y2=2.72
r101 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r102 37 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r103 36 51 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.59 $Y=2.72
+ $X2=7.915 $Y2=2.72
r104 36 37 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r105 34 37 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=7.59 $Y2=2.72
r106 34 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r107 33 36 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=7.59 $Y2=2.72
r108 33 34 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r109 31 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=3.59 $Y2=2.72
r110 31 33 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=3.91 $Y2=2.72
r111 29 48 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r112 29 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r113 28 29 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r114 26 44 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.92 $Y=2.72
+ $X2=0.727 $Y2=2.72
r115 26 28 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.92 $Y=2.72
+ $X2=1.15 $Y2=2.72
r116 25 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=2.72
+ $X2=3.59 $Y2=2.72
r117 25 28 148.422 $w=1.68e-07 $l=2.275e-06 $layer=LI1_cond $X=3.425 $Y=2.72
+ $X2=1.15 $Y2=2.72
r118 20 44 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.727 $Y2=2.72
r119 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.23 $Y2=2.72
r120 18 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r121 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r122 14 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.59 $Y=2.635
+ $X2=3.59 $Y2=2.72
r123 14 16 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.59 $Y=2.635
+ $X2=3.59 $Y2=2.32
r124 10 44 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.727 $Y=2.635
+ $X2=0.727 $Y2=2.72
r125 10 12 10.0278 $w=3.83e-07 $l=3.35e-07 $layer=LI1_cond $X=0.727 $Y=2.635
+ $X2=0.727 $Y2=2.3
r126 3 50 600 $w=1.7e-07 $l=1.01827e-06 $layer=licon1_PDIFF $count=1 $X=7.965
+ $Y=1.485 $X2=8.275 $Y2=2.36
r127 2 16 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.465
+ $Y=2.175 $X2=3.59 $Y2=2.32
r128 1 12 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.485 $X2=0.755 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_1%A_351_325# 1 2 3 4 13 17 22 24 25 28 29 30
+ 32 35 39 43 45 46 48
c153 29 0 1.36535e-19 $X=4.885 $Y=2.36
r154 46 47 17.602 $w=2.01e-07 $l=2.9e-07 $layer=LI1_cond $X=4.97 $Y=0.772
+ $X2=5.26 $Y2=0.772
r155 41 43 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.42 $Y=1.12
+ $X2=3.53 $Y2=1.12
r156 37 47 1.71937 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=5.26 $Y=0.655
+ $X2=5.26 $Y2=0.772
r157 37 39 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=5.26 $Y=0.655
+ $X2=5.26 $Y2=0.545
r158 33 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.055 $Y=2.36
+ $X2=4.97 $Y2=2.36
r159 33 35 131.786 $w=1.68e-07 $l=2.02e-06 $layer=LI1_cond $X=5.055 $Y=2.36
+ $X2=7.075 $Y2=2.36
r160 32 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.97 $Y=2.275
+ $X2=4.97 $Y2=2.36
r161 31 46 1.71937 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=4.97 $Y=0.89
+ $X2=4.97 $Y2=0.772
r162 31 32 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=4.97 $Y=0.89
+ $X2=4.97 $Y2=2.275
r163 29 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.885 $Y=2.36
+ $X2=4.97 $Y2=2.36
r164 29 30 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.885 $Y=2.36
+ $X2=4.36 $Y2=2.36
r165 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.275 $Y=2.275
+ $X2=4.36 $Y2=2.36
r166 27 28 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.275 $Y=2.065
+ $X2=4.275 $Y2=2.275
r167 26 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=1.98
+ $X2=3.53 $Y2=1.98
r168 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.19 $Y=1.98
+ $X2=4.275 $Y2=2.065
r169 25 26 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=4.19 $Y=1.98
+ $X2=3.615 $Y2=1.98
r170 24 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.53 $Y=1.895
+ $X2=3.53 $Y2=1.98
r171 23 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.53 $Y=1.205
+ $X2=3.53 $Y2=1.12
r172 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.53 $Y=1.205
+ $X2=3.53 $Y2=1.895
r173 22 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=1.035
+ $X2=3.42 $Y2=1.12
r174 21 22 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.42 $Y=0.455
+ $X2=3.42 $Y2=1.035
r175 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.335 $Y=0.37
+ $X2=3.42 $Y2=0.455
r176 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.335 $Y=0.37
+ $X2=3.04 $Y2=0.37
r177 13 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.445 $Y=1.98
+ $X2=3.53 $Y2=1.98
r178 13 15 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=3.445 $Y=1.98
+ $X2=1.945 $Y2=1.98
r179 4 35 600 $w=1.7e-07 $l=8.21995e-07 $layer=licon1_PDIFF $count=1 $X=6.845
+ $Y=1.645 $X2=7.075 $Y2=2.36
r180 3 15 600 $w=1.7e-07 $l=4.39858e-07 $layer=licon1_PDIFF $count=1 $X=1.755
+ $Y=1.625 $X2=1.945 $Y2=1.98
r181 2 39 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=5.125
+ $Y=0.245 $X2=5.26 $Y2=0.545
r182 1 19 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=2.835
+ $Y=0.245 $X2=3.04 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_1%A_375_49# 1 2 3 4 13 16 17 19 21 24 26 27
+ 29 34 35 36 37 40 43
c136 29 0 1.24749e-19 $X=6.92 $Y=0.38
r137 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.64 $Y=1.53
+ $X2=5.64 $Y2=1.53
r138 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.19 $Y=1.53
+ $X2=3.19 $Y2=1.53
r139 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.335 $Y=1.53
+ $X2=3.19 $Y2=1.53
r140 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.495 $Y=1.53
+ $X2=5.64 $Y2=1.53
r141 36 37 2.67326 $w=1.4e-07 $l=2.16e-06 $layer=MET1_cond $X=5.495 $Y=1.53
+ $X2=3.335 $Y2=1.53
r142 32 34 10.6148 $w=2.78e-07 $l=2.15e-07 $layer=LI1_cond $X=2.01 $Y=0.765
+ $X2=2.225 $Y2=0.765
r143 27 35 11.5258 $w=2.08e-07 $l=2.1e-07 $layer=LI1_cond $X=6.835 $Y=0.36
+ $X2=6.625 $Y2=0.36
r144 27 29 4.48918 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=6.835 $Y=0.36
+ $X2=6.92 $Y2=0.36
r145 26 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.115 $Y=0.34
+ $X2=6.625 $Y2=0.34
r146 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.03 $Y=0.425
+ $X2=6.115 $Y2=0.34
r147 23 24 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.03 $Y=0.425
+ $X2=6.03 $Y2=1.445
r148 22 44 6.03523 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=5.7 $Y=1.53
+ $X2=5.492 $Y2=1.53
r149 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.945 $Y=1.53
+ $X2=6.03 $Y2=1.445
r150 21 22 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.945 $Y=1.53
+ $X2=5.7 $Y2=1.53
r151 17 44 2.46632 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.492 $Y=1.615
+ $X2=5.492 $Y2=1.53
r152 17 19 0.138849 $w=4.13e-07 $l=5e-09 $layer=LI1_cond $X=5.492 $Y=1.615
+ $X2=5.492 $Y2=1.62
r153 16 40 8.59825 $w=3.35e-07 $l=1.55997e-07 $layer=LI1_cond $X=3.08 $Y=1.375
+ $X2=3.082 $Y2=1.53
r154 15 16 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.08 $Y=0.795
+ $X2=3.08 $Y2=1.375
r155 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.995 $Y=0.71
+ $X2=3.08 $Y2=0.795
r156 13 34 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.995 $Y=0.71
+ $X2=2.225 $Y2=0.71
r157 4 19 300 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_PDIFF $count=2 $X=5.115
+ $Y=1.485 $X2=5.46 $Y2=1.62
r158 3 40 600 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=2.805
+ $Y=1.485 $X2=3.055 $Y2=1.61
r159 2 29 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=6.725
+ $Y=0.245 $X2=6.92 $Y2=0.38
r160 1 32 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.875
+ $Y=0.245 $X2=2.01 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_1%A_1184_297# 1 2 3 4 15 18 23 26 29 31 36
r66 34 36 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=8.895 $Y=0.42
+ $X2=9.025 $Y2=0.42
r67 28 29 17.0922 $w=2.28e-07 $l=3.25e-07 $layer=LI1_cond $X=8.9 $Y=1.99
+ $X2=8.575 $Y2=1.99
r68 26 31 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.025 $Y=1.875
+ $X2=9.025 $Y2=1.99
r69 25 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.025 $Y=0.585
+ $X2=9.025 $Y2=0.42
r70 25 26 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=9.025 $Y=0.585
+ $X2=9.025 $Y2=1.875
r71 21 31 3.15669 $w=2.28e-07 $l=6.3e-08 $layer=LI1_cond $X=8.962 $Y=1.99
+ $X2=9.025 $Y2=1.99
r72 21 28 3.10659 $w=2.28e-07 $l=6.2e-08 $layer=LI1_cond $X=8.962 $Y=1.99
+ $X2=8.9 $Y2=1.99
r73 21 23 7.61784 $w=2.93e-07 $l=1.95e-07 $layer=LI1_cond $X=8.962 $Y=2.105
+ $X2=8.962 $Y2=2.3
r74 20 29 134.07 $w=1.68e-07 $l=2.055e-06 $layer=LI1_cond $X=6.52 $Y=2.02
+ $X2=8.575 $Y2=2.02
r75 18 20 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.455 $Y=2.02
+ $X2=6.52 $Y2=2.02
r76 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.37 $Y=1.935
+ $X2=6.455 $Y2=2.02
r77 13 15 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=6.37 $Y=1.935
+ $X2=6.37 $Y2=0.76
r78 4 28 600 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=1 $X=8.75
+ $Y=1.485 $X2=8.9 $Y2=1.96
r79 4 23 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=8.75
+ $Y=1.485 $X2=8.9 $Y2=2.3
r80 3 20 600 $w=1.7e-07 $l=8.25227e-07 $layer=licon1_PDIFF $count=1 $X=5.92
+ $Y=1.485 $X2=6.52 $Y2=2.02
r81 2 34 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=8.76
+ $Y=0.235 $X2=8.895 $Y2=0.42
r82 1 15 182 $w=1.7e-07 $l=7.01302e-07 $layer=licon1_NDIFF $count=1 $X=5.93
+ $Y=0.245 $X2=6.37 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_1%VGND 1 2 3 12 16 20 23 24 25 27 39 45 46
+ 49 52
c104 46 0 1.70967e-19 $X=8.97 $Y=0
c105 20 0 3.96944e-20 $X=8.285 $Y=0.4
r106 52 53 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r107 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r108 46 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=8.05
+ $Y2=0
r109 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r110 43 52 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=8.51 $Y=0 $X2=8.28
+ $Y2=0
r111 43 45 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=8.51 $Y=0 $X2=8.97
+ $Y2=0
r112 42 53 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=3.91 $Y=0 $X2=8.05
+ $Y2=0
r113 41 42 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r114 39 52 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=8.05 $Y=0 $X2=8.28
+ $Y2=0
r115 39 41 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=8.05 $Y=0 $X2=3.91
+ $Y2=0
r116 38 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r117 37 38 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r118 35 38 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r119 35 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r120 34 37 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r121 34 35 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r122 32 49 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.665
+ $Y2=0
r123 32 34 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=0
+ $X2=1.15 $Y2=0
r124 27 49 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.665
+ $Y2=0
r125 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r126 25 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r127 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r128 23 37 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.675 $Y=0
+ $X2=3.45 $Y2=0
r129 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=0 $X2=3.76
+ $Y2=0
r130 22 41 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.845 $Y=0 $X2=3.91
+ $Y2=0
r131 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.845 $Y=0 $X2=3.76
+ $Y2=0
r132 18 52 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.28 $Y=0.085
+ $X2=8.28 $Y2=0
r133 18 20 8.19054 $w=4.58e-07 $l=3.15e-07 $layer=LI1_cond $X=8.28 $Y=0.085
+ $X2=8.28 $Y2=0.4
r134 14 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.76 $Y=0.085
+ $X2=3.76 $Y2=0
r135 14 16 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.76 $Y=0.085
+ $X2=3.76 $Y2=0.36
r136 10 49 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=0.085
+ $X2=0.665 $Y2=0
r137 10 12 10.5641 $w=2.98e-07 $l=2.75e-07 $layer=LI1_cond $X=0.665 $Y=0.085
+ $X2=0.665 $Y2=0.36
r138 3 20 182 $w=1.7e-07 $l=3.83732e-07 $layer=licon1_NDIFF $count=1 $X=7.975
+ $Y=0.235 $X2=8.285 $Y2=0.4
r139 2 16 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=3.605
+ $Y=0.235 $X2=3.76 $Y2=0.36
r140 1 12 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.73 $Y2=0.36
.ends

