* File: sky130_fd_sc_hdll__clkmux2_4.pxi.spice
* Created: Thu Aug 27 19:03:37 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_4%A_79_199# N_A_79_199#_M1005_d
+ N_A_79_199#_M1013_d N_A_79_199#_c_97_n N_A_79_199#_M1000_g N_A_79_199#_M1003_g
+ N_A_79_199#_M1008_g N_A_79_199#_c_98_n N_A_79_199#_M1004_g N_A_79_199#_c_99_n
+ N_A_79_199#_M1010_g N_A_79_199#_M1011_g N_A_79_199#_M1014_g
+ N_A_79_199#_c_100_n N_A_79_199#_M1015_g N_A_79_199#_c_93_n N_A_79_199#_c_94_n
+ N_A_79_199#_c_187_p N_A_79_199#_c_95_n N_A_79_199#_c_125_p N_A_79_199#_c_108_p
+ N_A_79_199#_c_119_p N_A_79_199#_c_114_p N_A_79_199#_c_96_n
+ PM_SKY130_FD_SC_HDLL__CLKMUX2_4%A_79_199#
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_4%S N_S_c_222_n N_S_M1012_g N_S_M1016_g
+ N_S_c_224_n N_S_M1006_g N_S_M1002_g N_S_c_230_n N_S_c_248_n N_S_c_296_p
+ N_S_c_231_n N_S_c_271_p N_S_c_288_p N_S_c_226_n N_S_c_227_n S S
+ PM_SKY130_FD_SC_HDLL__CLKMUX2_4%S
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_4%A1 N_A1_M1005_g N_A1_c_318_n N_A1_M1007_g
+ N_A1_c_319_n N_A1_c_320_n N_A1_c_335_n N_A1_c_337_n A1 A1
+ PM_SKY130_FD_SC_HDLL__CLKMUX2_4%A1
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_4%A0 N_A0_c_390_n N_A0_M1013_g N_A0_c_391_n
+ N_A0_c_392_n N_A0_M1009_g N_A0_c_387_n A0 N_A0_c_388_n N_A0_c_389_n
+ PM_SKY130_FD_SC_HDLL__CLKMUX2_4%A0
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_4%A_925_21# N_A_925_21#_M1002_d
+ N_A_925_21#_M1006_d N_A_925_21#_M1001_g N_A_925_21#_c_437_n
+ N_A_925_21#_c_446_n N_A_925_21#_M1017_g N_A_925_21#_c_438_n
+ N_A_925_21#_c_439_n N_A_925_21#_c_440_n N_A_925_21#_c_441_n
+ N_A_925_21#_c_442_n N_A_925_21#_c_447_n N_A_925_21#_c_443_n
+ N_A_925_21#_c_444_n PM_SKY130_FD_SC_HDLL__CLKMUX2_4%A_925_21#
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_4%VPWR N_VPWR_M1000_d N_VPWR_M1004_d
+ N_VPWR_M1015_d N_VPWR_M1017_d N_VPWR_c_505_n N_VPWR_c_506_n N_VPWR_c_507_n
+ N_VPWR_c_508_n N_VPWR_c_509_n N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_512_n
+ VPWR N_VPWR_c_513_n N_VPWR_c_514_n N_VPWR_c_504_n N_VPWR_c_516_n
+ N_VPWR_c_517_n PM_SKY130_FD_SC_HDLL__CLKMUX2_4%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_4%X N_X_M1003_d N_X_M1011_d N_X_M1000_s
+ N_X_M1010_s N_X_c_574_n N_X_c_576_n N_X_c_570_n N_X_c_581_n N_X_c_572_n
+ N_X_c_585_n N_X_c_586_n N_X_c_588_n N_X_c_573_n X X X
+ PM_SKY130_FD_SC_HDLL__CLKMUX2_4%X
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_4%VGND N_VGND_M1003_s N_VGND_M1008_s
+ N_VGND_M1014_s N_VGND_M1001_d N_VGND_c_626_n N_VGND_c_627_n N_VGND_c_628_n
+ N_VGND_c_629_n VGND N_VGND_c_630_n N_VGND_c_631_n N_VGND_c_632_n
+ N_VGND_c_633_n N_VGND_c_634_n N_VGND_c_635_n N_VGND_c_636_n
+ PM_SKY130_FD_SC_HDLL__CLKMUX2_4%VGND
cc_1 VNB N_A_79_199#_M1003_g 0.0323163f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.495
cc_2 VNB N_A_79_199#_M1008_g 0.0238495f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.495
cc_3 VNB N_A_79_199#_M1011_g 0.0229096f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=0.495
cc_4 VNB N_A_79_199#_M1014_g 0.0241174f $X=-0.19 $Y=-0.24 $X2=1.87 $Y2=0.495
cc_5 VNB N_A_79_199#_c_93_n 0.00195867f $X=-0.19 $Y=-0.24 $X2=2 $Y2=1.16
cc_6 VNB N_A_79_199#_c_94_n 0.0180054f $X=-0.19 $Y=-0.24 $X2=2.815 $Y2=0.74
cc_7 VNB N_A_79_199#_c_95_n 0.00510464f $X=-0.19 $Y=-0.24 $X2=2.905 $Y2=1.955
cc_8 VNB N_A_79_199#_c_96_n 0.0967082f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_9 VNB N_S_c_222_n 0.0252932f $X=-0.19 $Y=-0.24 $X2=3.115 $Y2=0.235
cc_10 VNB N_S_M1016_g 0.0317183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_S_c_224_n 0.0209544f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_12 VNB N_S_M1002_g 0.0335245f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_S_c_226_n 5.74134e-19 $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_14 VNB N_S_c_227_n 0.0037048f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A1_M1005_g 0.0226218f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A1_c_318_n 0.0236121f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A1_c_319_n 0.0049634f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_18 VNB N_A1_c_320_n 0.0364624f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.495
cc_19 VNB A1 0.00997405f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.495
cc_20 VNB N_A0_M1009_g 0.0254644f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_21 VNB N_A0_c_387_n 0.00955013f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.495
cc_22 VNB N_A0_c_388_n 0.028761f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.495
cc_23 VNB N_A0_c_389_n 0.00455985f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.495
cc_24 VNB N_A_925_21#_M1001_g 0.02497f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_25 VNB N_A_925_21#_c_437_n 0.0070328f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.495
cc_26 VNB N_A_925_21#_c_438_n 5.32232e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_27 VNB N_A_925_21#_c_439_n 0.0308747f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_28 VNB N_A_925_21#_c_440_n 0.00551271f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_29 VNB N_A_925_21#_c_441_n 8.46441e-19 $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_30 VNB N_A_925_21#_c_442_n 0.0158392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_925_21#_c_443_n 0.0211382f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_32 VNB N_A_925_21#_c_444_n 0.0166335f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_33 VNB N_VPWR_c_504_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.202
cc_34 VNB N_X_c_570_n 0.00481412f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_35 VNB X 0.0014592f $X=-0.19 $Y=-0.24 $X2=2 $Y2=1.16
cc_36 VNB N_VGND_c_626_n 0.0124957f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_627_n 0.00458818f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.495
cc_38 VNB N_VGND_c_628_n 0.00397623f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_39 VNB N_VGND_c_629_n 0.00290835f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_40 VNB N_VGND_c_630_n 0.0177162f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_631_n 0.0156469f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_42 VNB N_VGND_c_632_n 0.0702689f $X=-0.19 $Y=-0.24 $X2=2 $Y2=1.16
cc_43 VNB N_VGND_c_633_n 0.0249556f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_634_n 0.304888f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=2.04
cc_45 VNB N_VGND_c_635_n 0.00480536f $X=-0.19 $Y=-0.24 $X2=2.902 $Y2=0.54
cc_46 VNB N_VGND_c_636_n 0.00564938f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=1.202
cc_47 VPB N_A_79_199#_c_97_n 0.0210619f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_48 VPB N_A_79_199#_c_98_n 0.0162324f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_49 VPB N_A_79_199#_c_99_n 0.015932f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_50 VPB N_A_79_199#_c_100_n 0.0174332f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_51 VPB N_A_79_199#_c_93_n 7.30825e-19 $X=-0.19 $Y=1.305 $X2=2 $Y2=1.16
cc_52 VPB N_A_79_199#_c_95_n 0.00428087f $X=-0.19 $Y=1.305 $X2=2.905 $Y2=1.955
cc_53 VPB N_A_79_199#_c_96_n 0.0557501f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_54 VPB N_S_c_222_n 0.0321847f $X=-0.19 $Y=1.305 $X2=3.115 $Y2=0.235
cc_55 VPB N_S_c_224_n 0.0330042f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_56 VPB N_S_c_230_n 0.0014488f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=0.495
cc_57 VPB N_S_c_231_n 6.63611e-19 $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_58 VPB N_S_c_226_n 6.16925e-19 $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_59 VPB N_S_c_227_n 0.00199981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB S 0.00455426f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_61 VPB N_A1_c_318_n 0.0304527f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A1_c_319_n 0.00280765f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.995
cc_63 VPB A1 0.00558813f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=0.495
cc_64 VPB N_A0_c_390_n 0.0205128f $X=-0.19 $Y=1.305 $X2=3.115 $Y2=0.235
cc_65 VPB N_A0_c_391_n 0.0406981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A0_c_392_n 0.00979353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A0_c_387_n 8.40892e-19 $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.495
cc_68 VPB N_A0_c_389_n 0.0023903f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=0.495
cc_69 VPB N_A_925_21#_c_437_n 0.00378234f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.495
cc_70 VPB N_A_925_21#_c_446_n 0.0224682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_925_21#_c_447_n 0.0267191f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_72 VPB N_A_925_21#_c_443_n 0.0225129f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_73 VPB N_VPWR_c_505_n 0.0114791f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_506_n 0.00466634f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=0.495
cc_75 VPB N_VPWR_c_507_n 0.00449767f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_76 VPB N_VPWR_c_508_n 0.0186115f $X=-0.19 $Y=1.305 $X2=1.45 $Y2=0.495
cc_77 VPB N_VPWR_c_509_n 0.00522692f $X=-0.19 $Y=1.305 $X2=1.87 $Y2=0.495
cc_78 VPB N_VPWR_c_510_n 0.00497347f $X=-0.19 $Y=1.305 $X2=2 $Y2=0.825
cc_79 VPB N_VPWR_c_511_n 0.062713f $X=-0.19 $Y=1.305 $X2=2 $Y2=1.16
cc_80 VPB N_VPWR_c_512_n 0.00439107f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_513_n 0.017949f $X=-0.19 $Y=1.305 $X2=2.905 $Y2=0.825
cc_82 VPB N_VPWR_c_514_n 0.0232568f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_83 VPB N_VPWR_c_504_n 0.0519448f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.202
cc_84 VPB N_VPWR_c_516_n 0.00458379f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_85 VPB N_VPWR_c_517_n 0.00525664f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_X_c_572_n 0.0020094f $X=-0.19 $Y=1.305 $X2=1.87 $Y2=0.495
cc_87 VPB N_X_c_573_n 0.00153266f $X=-0.19 $Y=1.305 $X2=2 $Y2=1.16
cc_88 N_A_79_199#_c_100_n N_S_c_222_n 0.0152157f $X=1.905 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_89 N_A_79_199#_c_93_n N_S_c_222_n 0.0010611f $X=2 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_90 N_A_79_199#_c_94_n N_S_c_222_n 0.00185825f $X=2.815 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_91 N_A_79_199#_c_95_n N_S_c_222_n 0.00377629f $X=2.905 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_92 N_A_79_199#_c_108_p N_S_c_222_n 6.79013e-19 $X=2.99 $Y=2.04 $X2=-0.19
+ $Y2=-0.24
cc_93 N_A_79_199#_c_96_n N_S_c_222_n 0.0236603f $X=1.905 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_94 N_A_79_199#_M1014_g N_S_M1016_g 0.0136976f $X=1.87 $Y=0.495 $X2=0 $Y2=0
cc_95 N_A_79_199#_c_93_n N_S_M1016_g 0.00297788f $X=2 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_79_199#_c_94_n N_S_M1016_g 0.0132761f $X=2.815 $Y=0.74 $X2=0 $Y2=0
cc_97 N_A_79_199#_c_95_n N_S_M1016_g 0.00349105f $X=2.905 $Y=1.955 $X2=0 $Y2=0
cc_98 N_A_79_199#_c_114_p N_S_M1016_g 0.007128f $X=2.902 $Y=0.54 $X2=0 $Y2=0
cc_99 N_A_79_199#_c_100_n N_S_c_230_n 6.36201e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A_79_199#_c_96_n N_S_c_230_n 4.77161e-19 $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_101 N_A_79_199#_M1013_d N_S_c_248_n 0.02385f $X=3.19 $Y=1.545 $X2=0 $Y2=0
cc_102 N_A_79_199#_c_108_p N_S_c_248_n 0.0100943f $X=2.99 $Y=2.04 $X2=0 $Y2=0
cc_103 N_A_79_199#_c_119_p N_S_c_248_n 0.0768599f $X=4.05 $Y=2.04 $X2=0 $Y2=0
cc_104 N_A_79_199#_c_93_n N_S_c_227_n 0.0151538f $X=2 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_79_199#_c_94_n N_S_c_227_n 0.0210402f $X=2.815 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A_79_199#_c_95_n N_S_c_227_n 0.0573306f $X=2.905 $Y=1.955 $X2=0 $Y2=0
cc_107 N_A_79_199#_c_96_n N_S_c_227_n 0.00131225f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_108 N_A_79_199#_c_95_n N_A1_M1005_g 2.48191e-19 $X=2.905 $Y=1.955 $X2=0 $Y2=0
cc_109 N_A_79_199#_c_125_p N_A1_M1005_g 0.0166772f $X=3.415 $Y=0.455 $X2=0 $Y2=0
cc_110 N_A_79_199#_c_114_p N_A1_M1005_g 0.0113941f $X=2.902 $Y=0.54 $X2=0 $Y2=0
cc_111 N_A_79_199#_c_119_p N_A1_c_318_n 0.00495514f $X=4.05 $Y=2.04 $X2=0 $Y2=0
cc_112 N_A_79_199#_M1013_d N_A1_c_319_n 0.00263273f $X=3.19 $Y=1.545 $X2=0 $Y2=0
cc_113 N_A_79_199#_c_95_n N_A1_c_319_n 0.053476f $X=2.905 $Y=1.955 $X2=0 $Y2=0
cc_114 N_A_79_199#_c_125_p N_A1_c_319_n 0.0126222f $X=3.415 $Y=0.455 $X2=0 $Y2=0
cc_115 N_A_79_199#_c_114_p N_A1_c_319_n 0.00119858f $X=2.902 $Y=0.54 $X2=0 $Y2=0
cc_116 N_A_79_199#_c_95_n N_A1_c_320_n 0.00712155f $X=2.905 $Y=1.955 $X2=0 $Y2=0
cc_117 N_A_79_199#_c_125_p N_A1_c_320_n 0.00418341f $X=3.415 $Y=0.455 $X2=0
+ $Y2=0
cc_118 N_A_79_199#_M1013_d N_A1_c_335_n 0.0262928f $X=3.19 $Y=1.545 $X2=0 $Y2=0
cc_119 N_A_79_199#_c_119_p N_A1_c_335_n 0.0639496f $X=4.05 $Y=2.04 $X2=0 $Y2=0
cc_120 N_A_79_199#_M1013_d N_A1_c_337_n 9.09665e-19 $X=3.19 $Y=1.545 $X2=0 $Y2=0
cc_121 N_A_79_199#_c_119_p N_A1_c_337_n 0.00891696f $X=4.05 $Y=2.04 $X2=0 $Y2=0
cc_122 N_A_79_199#_c_95_n N_A0_c_390_n 0.00328666f $X=2.905 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_123 N_A_79_199#_c_119_p N_A0_c_390_n 0.0138346f $X=4.05 $Y=2.04 $X2=-0.19
+ $Y2=-0.24
cc_124 N_A_79_199#_c_119_p N_A0_c_391_n 0.00104228f $X=4.05 $Y=2.04 $X2=0 $Y2=0
cc_125 N_A_79_199#_c_95_n N_A0_c_392_n 0.00173321f $X=2.905 $Y=1.955 $X2=0 $Y2=0
cc_126 N_A_79_199#_c_125_p N_A0_M1009_g 0.00342458f $X=3.415 $Y=0.455 $X2=0
+ $Y2=0
cc_127 N_A_79_199#_c_114_p N_A0_M1009_g 8.26503e-19 $X=2.902 $Y=0.54 $X2=0 $Y2=0
cc_128 N_A_79_199#_c_125_p N_A0_c_389_n 0.0299622f $X=3.415 $Y=0.455 $X2=0 $Y2=0
cc_129 N_A_79_199#_c_97_n N_VPWR_c_506_n 0.00354318f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_130 N_A_79_199#_c_98_n N_VPWR_c_507_n 0.0017219f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A_79_199#_c_99_n N_VPWR_c_507_n 0.00288097f $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_132 N_A_79_199#_c_96_n N_VPWR_c_507_n 0.00554477f $X=1.905 $Y=1.202 $X2=0
+ $Y2=0
cc_133 N_A_79_199#_c_99_n N_VPWR_c_508_n 0.00628074f $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_134 N_A_79_199#_c_100_n N_VPWR_c_508_n 0.00673617f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_135 N_A_79_199#_c_100_n N_VPWR_c_509_n 0.00333241f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_136 N_A_79_199#_c_93_n N_VPWR_c_509_n 0.00473648f $X=2 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_79_199#_c_94_n N_VPWR_c_509_n 0.00586099f $X=2.815 $Y=0.74 $X2=0
+ $Y2=0
cc_138 N_A_79_199#_c_96_n N_VPWR_c_509_n 0.0020312f $X=1.905 $Y=1.202 $X2=0
+ $Y2=0
cc_139 N_A_79_199#_c_97_n N_VPWR_c_513_n 0.00673617f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_140 N_A_79_199#_c_98_n N_VPWR_c_513_n 0.00673617f $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_141 N_A_79_199#_M1013_d N_VPWR_c_504_n 0.00817943f $X=3.19 $Y=1.545 $X2=0
+ $Y2=0
cc_142 N_A_79_199#_c_97_n N_VPWR_c_504_n 0.0126298f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_79_199#_c_98_n N_VPWR_c_504_n 0.0117184f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_79_199#_c_99_n N_VPWR_c_504_n 0.0106841f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_79_199#_c_100_n N_VPWR_c_504_n 0.0120575f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_146 N_A_79_199#_c_97_n N_X_c_574_n 0.00275587f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_79_199#_c_98_n N_X_c_574_n 0.00194755f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_79_199#_c_97_n N_X_c_576_n 0.00902937f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_79_199#_c_98_n N_X_c_576_n 0.00861078f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_79_199#_M1003_g N_X_c_570_n 0.0070553f $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_151 N_A_79_199#_M1008_g N_X_c_570_n 0.00401395f $X=0.93 $Y=0.495 $X2=0 $Y2=0
cc_152 N_A_79_199#_c_96_n N_X_c_570_n 0.00859968f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_153 N_A_79_199#_c_96_n N_X_c_581_n 0.0533f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_154 N_A_79_199#_c_97_n N_X_c_572_n 0.00206704f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_79_199#_c_98_n N_X_c_572_n 0.00108107f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_79_199#_c_96_n N_X_c_572_n 0.00549618f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_157 N_A_79_199#_c_96_n N_X_c_585_n 0.0246193f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_158 N_A_79_199#_c_93_n N_X_c_586_n 0.0198056f $X=2 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A_79_199#_c_96_n N_X_c_586_n 0.0154879f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_160 N_A_79_199#_c_99_n N_X_c_588_n 0.00226869f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A_79_199#_c_100_n N_X_c_588_n 0.00286667f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_79_199#_c_96_n N_X_c_588_n 0.00176607f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_163 N_A_79_199#_c_98_n N_X_c_573_n 5.02384e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_79_199#_c_99_n N_X_c_573_n 0.00245897f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A_79_199#_c_100_n N_X_c_573_n 0.0021314f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_79_199#_c_96_n N_X_c_573_n 0.00532378f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_167 N_A_79_199#_M1008_g X 0.00112312f $X=0.93 $Y=0.495 $X2=0 $Y2=0
cc_168 N_A_79_199#_M1011_g X 0.0154249f $X=1.45 $Y=0.495 $X2=0 $Y2=0
cc_169 N_A_79_199#_M1014_g X 0.00218271f $X=1.87 $Y=0.495 $X2=0 $Y2=0
cc_170 N_A_79_199#_c_93_n X 0.0174378f $X=2 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_79_199#_c_187_p X 0.00995765f $X=2.085 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A_79_199#_c_96_n X 0.00677505f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_173 N_A_79_199#_c_99_n X 0.0103556f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_79_199#_c_100_n X 0.00862367f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_79_199#_c_95_n A_523_309# 0.00524208f $X=2.905 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_176 N_A_79_199#_c_108_p A_523_309# 0.00299062f $X=2.99 $Y=2.04 $X2=-0.19
+ $Y2=-0.24
cc_177 N_A_79_199#_c_94_n N_VGND_M1014_s 0.00213207f $X=2.815 $Y=0.74 $X2=0
+ $Y2=0
cc_178 N_A_79_199#_c_187_p N_VGND_M1014_s 8.75693e-19 $X=2.085 $Y=0.74 $X2=0
+ $Y2=0
cc_179 N_A_79_199#_M1003_g N_VGND_c_627_n 0.0045924f $X=0.51 $Y=0.495 $X2=0
+ $Y2=0
cc_180 N_A_79_199#_M1008_g N_VGND_c_628_n 0.00193867f $X=0.93 $Y=0.495 $X2=0
+ $Y2=0
cc_181 N_A_79_199#_M1011_g N_VGND_c_628_n 0.00314364f $X=1.45 $Y=0.495 $X2=0
+ $Y2=0
cc_182 N_A_79_199#_c_96_n N_VGND_c_628_n 0.00413946f $X=1.905 $Y=1.202 $X2=0
+ $Y2=0
cc_183 N_A_79_199#_M1011_g N_VGND_c_629_n 6.08654e-19 $X=1.45 $Y=0.495 $X2=0
+ $Y2=0
cc_184 N_A_79_199#_M1014_g N_VGND_c_629_n 0.00757456f $X=1.87 $Y=0.495 $X2=0
+ $Y2=0
cc_185 N_A_79_199#_c_94_n N_VGND_c_629_n 0.014523f $X=2.815 $Y=0.74 $X2=0 $Y2=0
cc_186 N_A_79_199#_c_187_p N_VGND_c_629_n 0.00929542f $X=2.085 $Y=0.74 $X2=0
+ $Y2=0
cc_187 N_A_79_199#_c_114_p N_VGND_c_629_n 0.00829663f $X=2.902 $Y=0.54 $X2=0
+ $Y2=0
cc_188 N_A_79_199#_c_96_n N_VGND_c_629_n 5.28291e-19 $X=1.905 $Y=1.202 $X2=0
+ $Y2=0
cc_189 N_A_79_199#_M1003_g N_VGND_c_630_n 0.00585385f $X=0.51 $Y=0.495 $X2=0
+ $Y2=0
cc_190 N_A_79_199#_M1008_g N_VGND_c_630_n 0.00585385f $X=0.93 $Y=0.495 $X2=0
+ $Y2=0
cc_191 N_A_79_199#_M1011_g N_VGND_c_631_n 0.00510997f $X=1.45 $Y=0.495 $X2=0
+ $Y2=0
cc_192 N_A_79_199#_M1014_g N_VGND_c_631_n 0.0046653f $X=1.87 $Y=0.495 $X2=0
+ $Y2=0
cc_193 N_A_79_199#_c_94_n N_VGND_c_632_n 0.00916117f $X=2.815 $Y=0.74 $X2=0
+ $Y2=0
cc_194 N_A_79_199#_c_125_p N_VGND_c_632_n 0.0319877f $X=3.415 $Y=0.455 $X2=0
+ $Y2=0
cc_195 N_A_79_199#_c_114_p N_VGND_c_632_n 0.0102622f $X=2.902 $Y=0.54 $X2=0
+ $Y2=0
cc_196 N_A_79_199#_M1005_d N_VGND_c_634_n 0.00824573f $X=3.115 $Y=0.235 $X2=0
+ $Y2=0
cc_197 N_A_79_199#_M1003_g N_VGND_c_634_n 0.0116294f $X=0.51 $Y=0.495 $X2=0
+ $Y2=0
cc_198 N_A_79_199#_M1008_g N_VGND_c_634_n 0.0109403f $X=0.93 $Y=0.495 $X2=0
+ $Y2=0
cc_199 N_A_79_199#_M1011_g N_VGND_c_634_n 0.00917818f $X=1.45 $Y=0.495 $X2=0
+ $Y2=0
cc_200 N_A_79_199#_M1014_g N_VGND_c_634_n 0.00796766f $X=1.87 $Y=0.495 $X2=0
+ $Y2=0
cc_201 N_A_79_199#_c_94_n N_VGND_c_634_n 0.0151571f $X=2.815 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A_79_199#_c_187_p N_VGND_c_634_n 8.0899e-19 $X=2.085 $Y=0.74 $X2=0
+ $Y2=0
cc_203 N_A_79_199#_c_125_p N_VGND_c_634_n 0.0187496f $X=3.415 $Y=0.455 $X2=0
+ $Y2=0
cc_204 N_A_79_199#_c_114_p N_VGND_c_634_n 0.00662435f $X=2.902 $Y=0.54 $X2=0
+ $Y2=0
cc_205 N_A_79_199#_c_114_p A_525_47# 0.00646906f $X=2.902 $Y=0.54 $X2=-0.19
+ $Y2=-0.24
cc_206 N_S_M1016_g N_A1_M1005_g 0.0169272f $X=2.55 $Y=0.445 $X2=0 $Y2=0
cc_207 N_S_c_248_n N_A1_c_318_n 0.0140173f $X=4.625 $Y=2.38 $X2=0 $Y2=0
cc_208 N_S_c_231_n N_A1_c_318_n 3.3557e-19 $X=4.71 $Y=1.63 $X2=0 $Y2=0
cc_209 N_S_c_222_n N_A1_c_320_n 0.0169272f $X=2.525 $Y=1.47 $X2=0 $Y2=0
cc_210 N_S_c_227_n N_A1_c_320_n 2.91356e-19 $X=2.48 $Y=1.16 $X2=0 $Y2=0
cc_211 N_S_c_248_n N_A1_c_335_n 0.00421347f $X=4.625 $Y=2.38 $X2=0 $Y2=0
cc_212 N_S_c_231_n A1 0.0117446f $X=4.71 $Y=1.63 $X2=0 $Y2=0
cc_213 N_S_c_222_n N_A0_c_390_n 0.031348f $X=2.525 $Y=1.47 $X2=-0.19 $Y2=-0.24
cc_214 N_S_c_248_n N_A0_c_390_n 0.0134713f $X=4.625 $Y=2.38 $X2=-0.19 $Y2=-0.24
cc_215 N_S_c_222_n N_A0_c_392_n 0.00442896f $X=2.525 $Y=1.47 $X2=0 $Y2=0
cc_216 N_S_M1002_g N_A_925_21#_M1001_g 0.0166525f $X=5.32 $Y=0.495 $X2=0 $Y2=0
cc_217 N_S_c_224_n N_A_925_21#_c_437_n 0.00791167f $X=5.295 $Y=1.47 $X2=0 $Y2=0
cc_218 N_S_c_226_n N_A_925_21#_c_437_n 0.00114571f $X=5.27 $Y=1.22 $X2=0 $Y2=0
cc_219 N_S_c_224_n N_A_925_21#_c_446_n 0.0253237f $X=5.295 $Y=1.47 $X2=0 $Y2=0
cc_220 N_S_c_248_n N_A_925_21#_c_446_n 0.00665392f $X=4.625 $Y=2.38 $X2=0 $Y2=0
cc_221 N_S_c_231_n N_A_925_21#_c_446_n 0.00936369f $X=4.71 $Y=1.63 $X2=0 $Y2=0
cc_222 N_S_c_271_p N_A_925_21#_c_446_n 0.0169742f $X=4.71 $Y=2.295 $X2=0 $Y2=0
cc_223 N_S_c_226_n N_A_925_21#_c_446_n 9.61528e-19 $X=5.27 $Y=1.22 $X2=0 $Y2=0
cc_224 S N_A_925_21#_c_446_n 0.00468862f $X=5.185 $Y=1.445 $X2=0 $Y2=0
cc_225 N_S_c_224_n N_A_925_21#_c_438_n 4.2108e-19 $X=5.295 $Y=1.47 $X2=0 $Y2=0
cc_226 N_S_M1002_g N_A_925_21#_c_438_n 0.00105012f $X=5.32 $Y=0.495 $X2=0 $Y2=0
cc_227 N_S_c_231_n N_A_925_21#_c_438_n 0.00529971f $X=4.71 $Y=1.63 $X2=0 $Y2=0
cc_228 N_S_c_226_n N_A_925_21#_c_438_n 0.00549551f $X=5.27 $Y=1.22 $X2=0 $Y2=0
cc_229 S N_A_925_21#_c_438_n 0.00442941f $X=5.185 $Y=1.445 $X2=0 $Y2=0
cc_230 N_S_c_224_n N_A_925_21#_c_439_n 0.0078874f $X=5.295 $Y=1.47 $X2=0 $Y2=0
cc_231 N_S_M1002_g N_A_925_21#_c_439_n 0.00773768f $X=5.32 $Y=0.495 $X2=0 $Y2=0
cc_232 N_S_c_226_n N_A_925_21#_c_439_n 4.28614e-19 $X=5.27 $Y=1.22 $X2=0 $Y2=0
cc_233 S N_A_925_21#_c_439_n 0.00155646f $X=5.185 $Y=1.445 $X2=0 $Y2=0
cc_234 N_S_c_224_n N_A_925_21#_c_440_n 0.00210123f $X=5.295 $Y=1.47 $X2=0 $Y2=0
cc_235 N_S_M1002_g N_A_925_21#_c_440_n 0.0151946f $X=5.32 $Y=0.495 $X2=0 $Y2=0
cc_236 N_S_c_226_n N_A_925_21#_c_440_n 0.0131349f $X=5.27 $Y=1.22 $X2=0 $Y2=0
cc_237 S N_A_925_21#_c_440_n 0.00986081f $X=5.185 $Y=1.445 $X2=0 $Y2=0
cc_238 N_S_c_224_n N_A_925_21#_c_447_n 0.00747341f $X=5.295 $Y=1.47 $X2=0 $Y2=0
cc_239 N_S_c_288_p N_A_925_21#_c_447_n 6.43652e-19 $X=5.28 $Y=1.44 $X2=0 $Y2=0
cc_240 N_S_c_224_n N_A_925_21#_c_443_n 0.0171101f $X=5.295 $Y=1.47 $X2=0 $Y2=0
cc_241 N_S_M1002_g N_A_925_21#_c_443_n 0.00462428f $X=5.32 $Y=0.495 $X2=0 $Y2=0
cc_242 N_S_c_288_p N_A_925_21#_c_443_n 0.0123401f $X=5.28 $Y=1.44 $X2=0 $Y2=0
cc_243 N_S_c_226_n N_A_925_21#_c_443_n 0.0228671f $X=5.27 $Y=1.22 $X2=0 $Y2=0
cc_244 S N_VPWR_M1017_d 0.00577639f $X=5.185 $Y=1.445 $X2=0 $Y2=0
cc_245 N_S_c_222_n N_VPWR_c_509_n 0.0105378f $X=2.525 $Y=1.47 $X2=0 $Y2=0
cc_246 N_S_c_230_n N_VPWR_c_509_n 0.0589849f $X=2.55 $Y=2.295 $X2=0 $Y2=0
cc_247 N_S_c_296_p N_VPWR_c_509_n 0.0138248f $X=2.65 $Y=2.38 $X2=0 $Y2=0
cc_248 N_S_c_224_n N_VPWR_c_510_n 0.00324489f $X=5.295 $Y=1.47 $X2=0 $Y2=0
cc_249 N_S_c_248_n N_VPWR_c_510_n 0.0136491f $X=4.625 $Y=2.38 $X2=0 $Y2=0
cc_250 N_S_c_271_p N_VPWR_c_510_n 0.0330344f $X=4.71 $Y=2.295 $X2=0 $Y2=0
cc_251 S N_VPWR_c_510_n 0.0129774f $X=5.185 $Y=1.445 $X2=0 $Y2=0
cc_252 N_S_c_222_n N_VPWR_c_511_n 0.00451973f $X=2.525 $Y=1.47 $X2=0 $Y2=0
cc_253 N_S_c_248_n N_VPWR_c_511_n 0.127436f $X=4.625 $Y=2.38 $X2=0 $Y2=0
cc_254 N_S_c_296_p N_VPWR_c_511_n 0.0124588f $X=2.65 $Y=2.38 $X2=0 $Y2=0
cc_255 N_S_c_224_n N_VPWR_c_514_n 0.00673617f $X=5.295 $Y=1.47 $X2=0 $Y2=0
cc_256 N_S_c_222_n N_VPWR_c_504_n 0.00727617f $X=2.525 $Y=1.47 $X2=0 $Y2=0
cc_257 N_S_c_224_n N_VPWR_c_504_n 0.0130085f $X=5.295 $Y=1.47 $X2=0 $Y2=0
cc_258 N_S_c_248_n N_VPWR_c_504_n 0.07773f $X=4.625 $Y=2.38 $X2=0 $Y2=0
cc_259 N_S_c_296_p N_VPWR_c_504_n 0.00693792f $X=2.65 $Y=2.38 $X2=0 $Y2=0
cc_260 N_S_c_248_n A_523_309# 0.0100148f $X=4.625 $Y=2.38 $X2=-0.19 $Y2=-0.24
cc_261 N_S_c_248_n A_875_309# 0.00646556f $X=4.625 $Y=2.38 $X2=-0.19 $Y2=-0.24
cc_262 N_S_M1016_g N_VGND_c_629_n 0.00567875f $X=2.55 $Y=0.445 $X2=0 $Y2=0
cc_263 N_S_M1016_g N_VGND_c_632_n 0.00428022f $X=2.55 $Y=0.445 $X2=0 $Y2=0
cc_264 N_S_M1002_g N_VGND_c_632_n 0.00646436f $X=5.32 $Y=0.495 $X2=0 $Y2=0
cc_265 N_S_M1002_g N_VGND_c_633_n 0.00433717f $X=5.32 $Y=0.495 $X2=0 $Y2=0
cc_266 N_S_M1016_g N_VGND_c_634_n 0.006683f $X=2.55 $Y=0.445 $X2=0 $Y2=0
cc_267 N_S_M1002_g N_VGND_c_634_n 0.00761805f $X=5.32 $Y=0.495 $X2=0 $Y2=0
cc_268 N_A1_c_319_n N_A0_c_390_n 0.00408958f $X=3.245 $Y=0.975 $X2=-0.19
+ $Y2=-0.24
cc_269 N_A1_c_337_n N_A0_c_390_n 0.00649431f $X=3.33 $Y=1.7 $X2=-0.19 $Y2=-0.24
cc_270 N_A1_c_318_n N_A0_c_391_n 0.00277644f $X=4.285 $Y=1.47 $X2=0 $Y2=0
cc_271 N_A1_c_319_n N_A0_c_391_n 0.0101853f $X=3.245 $Y=0.975 $X2=0 $Y2=0
cc_272 N_A1_c_335_n N_A0_c_391_n 0.016411f $X=4.165 $Y=1.7 $X2=0 $Y2=0
cc_273 A1 N_A0_c_391_n 0.00120799f $X=4.285 $Y=0.765 $X2=0 $Y2=0
cc_274 N_A1_c_319_n N_A0_c_392_n 0.00201932f $X=3.245 $Y=0.975 $X2=0 $Y2=0
cc_275 N_A1_c_320_n N_A0_c_392_n 0.0292599f $X=3.245 $Y=0.975 $X2=0 $Y2=0
cc_276 N_A1_M1005_g N_A0_M1009_g 0.0140866f $X=3.04 $Y=0.445 $X2=0 $Y2=0
cc_277 N_A1_c_319_n N_A0_M1009_g 2.42785e-19 $X=3.245 $Y=0.975 $X2=0 $Y2=0
cc_278 A1 N_A0_M1009_g 0.00248702f $X=4.285 $Y=0.765 $X2=0 $Y2=0
cc_279 N_A1_c_318_n N_A0_c_387_n 0.00936614f $X=4.285 $Y=1.47 $X2=0 $Y2=0
cc_280 A1 N_A0_c_387_n 2.12428e-19 $X=4.285 $Y=0.765 $X2=0 $Y2=0
cc_281 N_A1_c_318_n N_A0_c_388_n 0.00503691f $X=4.285 $Y=1.47 $X2=0 $Y2=0
cc_282 N_A1_c_319_n N_A0_c_388_n 0.00486025f $X=3.245 $Y=0.975 $X2=0 $Y2=0
cc_283 N_A1_c_320_n N_A0_c_388_n 0.0169793f $X=3.245 $Y=0.975 $X2=0 $Y2=0
cc_284 N_A1_c_335_n N_A0_c_388_n 2.70133e-19 $X=4.165 $Y=1.7 $X2=0 $Y2=0
cc_285 A1 N_A0_c_388_n 0.00144026f $X=4.285 $Y=0.765 $X2=0 $Y2=0
cc_286 N_A1_M1005_g N_A0_c_389_n 0.00121146f $X=3.04 $Y=0.445 $X2=0 $Y2=0
cc_287 N_A1_c_318_n N_A0_c_389_n 0.00240846f $X=4.285 $Y=1.47 $X2=0 $Y2=0
cc_288 N_A1_c_319_n N_A0_c_389_n 0.0256133f $X=3.245 $Y=0.975 $X2=0 $Y2=0
cc_289 N_A1_c_320_n N_A0_c_389_n 9.69032e-19 $X=3.245 $Y=0.975 $X2=0 $Y2=0
cc_290 N_A1_c_335_n N_A0_c_389_n 0.0231818f $X=4.165 $Y=1.7 $X2=0 $Y2=0
cc_291 A1 N_A0_c_389_n 0.0929962f $X=4.285 $Y=0.765 $X2=0 $Y2=0
cc_292 A1 N_A_925_21#_M1001_g 0.0260542f $X=4.285 $Y=0.765 $X2=0 $Y2=0
cc_293 N_A1_c_318_n N_A_925_21#_c_446_n 0.0556404f $X=4.285 $Y=1.47 $X2=0 $Y2=0
cc_294 N_A1_c_335_n N_A_925_21#_c_446_n 6.59428e-19 $X=4.165 $Y=1.7 $X2=0 $Y2=0
cc_295 A1 N_A_925_21#_c_446_n 5.7392e-19 $X=4.285 $Y=0.765 $X2=0 $Y2=0
cc_296 A1 N_A_925_21#_c_438_n 0.0179199f $X=4.285 $Y=0.765 $X2=0 $Y2=0
cc_297 N_A1_c_318_n N_A_925_21#_c_439_n 0.0213383f $X=4.285 $Y=1.47 $X2=0 $Y2=0
cc_298 A1 N_A_925_21#_c_441_n 0.0105375f $X=4.285 $Y=0.765 $X2=0 $Y2=0
cc_299 N_A1_c_318_n N_VPWR_c_511_n 0.00429453f $X=4.285 $Y=1.47 $X2=0 $Y2=0
cc_300 N_A1_c_318_n N_VPWR_c_504_n 0.0073872f $X=4.285 $Y=1.47 $X2=0 $Y2=0
cc_301 N_A1_c_335_n A_875_309# 0.0019065f $X=4.165 $Y=1.7 $X2=-0.19 $Y2=-0.24
cc_302 A1 A_875_309# 5.87758e-19 $X=4.285 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_303 N_A1_M1005_g N_VGND_c_632_n 0.00357842f $X=3.04 $Y=0.445 $X2=0 $Y2=0
cc_304 A1 N_VGND_c_632_n 0.041242f $X=4.285 $Y=0.765 $X2=0 $Y2=0
cc_305 N_A1_M1005_g N_VGND_c_634_n 0.00598057f $X=3.04 $Y=0.445 $X2=0 $Y2=0
cc_306 A1 N_VGND_c_634_n 0.0110914f $X=4.285 $Y=0.765 $X2=0 $Y2=0
cc_307 A1 A_754_47# 0.0167608f $X=4.285 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_308 N_A0_c_390_n N_VPWR_c_511_n 0.00429453f $X=3.1 $Y=1.47 $X2=0 $Y2=0
cc_309 N_A0_c_390_n N_VPWR_c_504_n 0.00770108f $X=3.1 $Y=1.47 $X2=0 $Y2=0
cc_310 N_A0_M1009_g N_VGND_c_632_n 0.00435091f $X=3.695 $Y=0.445 $X2=0 $Y2=0
cc_311 N_A0_c_389_n N_VGND_c_632_n 0.0205158f $X=3.755 $Y=0.98 $X2=0 $Y2=0
cc_312 N_A0_M1009_g N_VGND_c_634_n 0.00904666f $X=3.695 $Y=0.445 $X2=0 $Y2=0
cc_313 N_A0_c_389_n N_VGND_c_634_n 0.0119866f $X=3.755 $Y=0.98 $X2=0 $Y2=0
cc_314 N_A0_c_389_n A_754_47# 0.00656391f $X=3.755 $Y=0.98 $X2=-0.19 $Y2=-0.24
cc_315 N_A_925_21#_c_446_n N_VPWR_c_510_n 0.00744201f $X=4.725 $Y=1.47 $X2=0
+ $Y2=0
cc_316 N_A_925_21#_c_446_n N_VPWR_c_511_n 0.00459563f $X=4.725 $Y=1.47 $X2=0
+ $Y2=0
cc_317 N_A_925_21#_c_447_n N_VPWR_c_514_n 0.0259839f $X=5.53 $Y=2 $X2=0 $Y2=0
cc_318 N_A_925_21#_M1006_d N_VPWR_c_504_n 0.00233913f $X=5.385 $Y=1.545 $X2=0
+ $Y2=0
cc_319 N_A_925_21#_c_446_n N_VPWR_c_504_n 0.00704825f $X=4.725 $Y=1.47 $X2=0
+ $Y2=0
cc_320 N_A_925_21#_c_447_n N_VPWR_c_504_n 0.0151509f $X=5.53 $Y=2 $X2=0 $Y2=0
cc_321 N_A_925_21#_c_440_n N_VGND_M1001_d 0.00234003f $X=5.415 $Y=0.78 $X2=0
+ $Y2=0
cc_322 N_A_925_21#_M1001_g N_VGND_c_632_n 0.023697f $X=4.7 $Y=0.445 $X2=0 $Y2=0
cc_323 N_A_925_21#_c_439_n N_VGND_c_632_n 6.87788e-19 $X=4.79 $Y=1.02 $X2=0
+ $Y2=0
cc_324 N_A_925_21#_c_440_n N_VGND_c_632_n 0.0210008f $X=5.415 $Y=0.78 $X2=0
+ $Y2=0
cc_325 N_A_925_21#_c_441_n N_VGND_c_632_n 0.0115145f $X=4.875 $Y=0.78 $X2=0
+ $Y2=0
cc_326 N_A_925_21#_c_440_n N_VGND_c_633_n 0.00345018f $X=5.415 $Y=0.78 $X2=0
+ $Y2=0
cc_327 N_A_925_21#_c_442_n N_VGND_c_633_n 0.0157596f $X=5.53 $Y=0.455 $X2=0
+ $Y2=0
cc_328 N_A_925_21#_c_444_n N_VGND_c_633_n 0.00189167f $X=5.59 $Y=0.78 $X2=0
+ $Y2=0
cc_329 N_A_925_21#_M1002_d N_VGND_c_634_n 0.00218371f $X=5.395 $Y=0.235 $X2=0
+ $Y2=0
cc_330 N_A_925_21#_M1001_g N_VGND_c_634_n 0.00251647f $X=4.7 $Y=0.445 $X2=0
+ $Y2=0
cc_331 N_A_925_21#_c_440_n N_VGND_c_634_n 0.00766116f $X=5.415 $Y=0.78 $X2=0
+ $Y2=0
cc_332 N_A_925_21#_c_441_n N_VGND_c_634_n 7.21038e-19 $X=4.875 $Y=0.78 $X2=0
+ $Y2=0
cc_333 N_A_925_21#_c_442_n N_VGND_c_634_n 0.0093388f $X=5.53 $Y=0.455 $X2=0
+ $Y2=0
cc_334 N_A_925_21#_c_444_n N_VGND_c_634_n 0.00302259f $X=5.59 $Y=0.78 $X2=0
+ $Y2=0
cc_335 N_VPWR_c_504_n N_X_M1000_s 0.00231261f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_336 N_VPWR_c_504_n N_X_M1010_s 0.00231261f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_337 N_VPWR_c_513_n N_X_c_576_n 0.0189467f $X=1.065 $Y=2.72 $X2=0 $Y2=0
cc_338 N_VPWR_c_504_n N_X_c_576_n 0.0123027f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_339 N_VPWR_c_507_n N_X_c_581_n 0.0165498f $X=1.2 $Y=1.66 $X2=0 $Y2=0
cc_340 N_VPWR_c_508_n X 0.0209921f $X=2.005 $Y=2.72 $X2=0 $Y2=0
cc_341 N_VPWR_c_504_n X 0.0133313f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_342 N_VPWR_c_504_n A_523_309# 0.00317215f $X=5.75 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_343 N_VPWR_c_504_n A_875_309# 0.00208801f $X=5.75 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_344 N_X_c_581_n N_VGND_c_628_n 0.0100833f $X=1.475 $Y=1.195 $X2=0 $Y2=0
cc_345 X N_VGND_c_628_n 0.0299439f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_346 N_X_c_570_n N_VGND_c_630_n 0.0145891f $X=0.72 $Y=0.49 $X2=0 $Y2=0
cc_347 X N_VGND_c_631_n 0.0165462f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_348 N_X_M1003_d N_VGND_c_634_n 0.00258466f $X=0.585 $Y=0.235 $X2=0 $Y2=0
cc_349 N_X_M1011_d N_VGND_c_634_n 0.00393857f $X=1.525 $Y=0.235 $X2=0 $Y2=0
cc_350 N_X_c_570_n N_VGND_c_634_n 0.00993603f $X=0.72 $Y=0.49 $X2=0 $Y2=0
cc_351 X N_VGND_c_634_n 0.0100971f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_352 N_VGND_c_634_n A_525_47# 0.0034784f $X=5.75 $Y=0 $X2=-0.19 $Y2=-0.24
cc_353 N_VGND_c_634_n A_754_47# 0.0188707f $X=5.75 $Y=0 $X2=-0.19 $Y2=-0.24
