* File: sky130_fd_sc_hdll__clkbuf_16.pxi.spice
* Created: Wed Sep  2 08:25:19 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKBUF_16%A N_A_c_150_n N_A_M1013_g N_A_M1006_g
+ N_A_c_151_n N_A_M1014_g N_A_M1007_g N_A_c_152_n N_A_M1030_g N_A_M1011_g
+ N_A_c_153_n N_A_M1034_g N_A_M1023_g A A N_A_c_149_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_16%A
x_PM_SKY130_FD_SC_HDLL__CLKBUF_16%A_118_297# N_A_118_297#_M1006_d
+ N_A_118_297#_M1011_d N_A_118_297#_M1013_d N_A_118_297#_M1030_d
+ N_A_118_297#_M1000_g N_A_118_297#_c_228_n N_A_118_297#_M1003_g
+ N_A_118_297#_M1001_g N_A_118_297#_c_229_n N_A_118_297#_M1004_g
+ N_A_118_297#_M1002_g N_A_118_297#_c_230_n N_A_118_297#_M1008_g
+ N_A_118_297#_M1005_g N_A_118_297#_c_231_n N_A_118_297#_M1009_g
+ N_A_118_297#_M1012_g N_A_118_297#_c_232_n N_A_118_297#_M1010_g
+ N_A_118_297#_M1017_g N_A_118_297#_c_233_n N_A_118_297#_M1015_g
+ N_A_118_297#_M1019_g N_A_118_297#_c_234_n N_A_118_297#_M1016_g
+ N_A_118_297#_M1020_g N_A_118_297#_c_235_n N_A_118_297#_M1018_g
+ N_A_118_297#_M1021_g N_A_118_297#_c_236_n N_A_118_297#_M1022_g
+ N_A_118_297#_M1024_g N_A_118_297#_c_237_n N_A_118_297#_M1025_g
+ N_A_118_297#_M1027_g N_A_118_297#_c_238_n N_A_118_297#_M1026_g
+ N_A_118_297#_M1032_g N_A_118_297#_c_239_n N_A_118_297#_M1028_g
+ N_A_118_297#_M1033_g N_A_118_297#_c_240_n N_A_118_297#_M1029_g
+ N_A_118_297#_M1036_g N_A_118_297#_c_241_n N_A_118_297#_M1031_g
+ N_A_118_297#_M1037_g N_A_118_297#_c_242_n N_A_118_297#_M1035_g
+ N_A_118_297#_c_243_n N_A_118_297#_M1038_g N_A_118_297#_M1039_g
+ N_A_118_297#_c_224_n N_A_118_297#_c_244_n N_A_118_297#_c_257_n
+ N_A_118_297#_c_225_n N_A_118_297#_c_245_n N_A_118_297#_c_226_n
+ N_A_118_297#_c_265_n N_A_118_297#_c_267_n N_A_118_297#_c_227_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_16%A_118_297#
x_PM_SKY130_FD_SC_HDLL__CLKBUF_16%VPWR N_VPWR_M1013_s N_VPWR_M1014_s
+ N_VPWR_M1034_s N_VPWR_M1004_s N_VPWR_M1009_s N_VPWR_M1015_s N_VPWR_M1018_s
+ N_VPWR_M1025_s N_VPWR_M1028_s N_VPWR_M1031_s N_VPWR_M1038_s N_VPWR_c_486_n
+ N_VPWR_c_487_n N_VPWR_c_488_n N_VPWR_c_489_n N_VPWR_c_490_n N_VPWR_c_491_n
+ N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_494_n N_VPWR_c_495_n N_VPWR_c_496_n
+ N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_500_n N_VPWR_c_501_n
+ N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n N_VPWR_c_506_n
+ N_VPWR_c_507_n N_VPWR_c_508_n N_VPWR_c_509_n N_VPWR_c_510_n N_VPWR_c_511_n
+ N_VPWR_c_512_n N_VPWR_c_513_n N_VPWR_c_514_n VPWR N_VPWR_c_515_n
+ N_VPWR_c_516_n N_VPWR_c_517_n N_VPWR_c_485_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_16%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKBUF_16%X N_X_M1000_s N_X_M1002_s N_X_M1012_s
+ N_X_M1019_s N_X_M1021_s N_X_M1027_s N_X_M1033_s N_X_M1037_s N_X_M1003_d
+ N_X_M1008_d N_X_M1010_d N_X_M1016_d N_X_M1022_d N_X_M1026_d N_X_M1029_d
+ N_X_M1035_d N_X_c_631_n N_X_c_632_n N_X_c_633_n N_X_c_664_n N_X_c_634_n
+ N_X_c_635_n N_X_c_674_n N_X_c_636_n N_X_c_637_n N_X_c_684_n N_X_c_638_n
+ N_X_c_639_n N_X_c_695_n N_X_c_640_n N_X_c_641_n N_X_c_705_n N_X_c_642_n
+ N_X_c_643_n N_X_c_644_n N_X_c_645_n N_X_c_777_n N_X_c_646_n N_X_c_724_n
+ N_X_c_647_n N_X_c_728_n N_X_c_648_n N_X_c_732_n N_X_c_649_n N_X_c_737_n
+ N_X_c_650_n N_X_c_741_n N_X_c_651_n N_X_c_745_n N_X_c_652_n X X X N_X_c_756_n
+ X PM_SKY130_FD_SC_HDLL__CLKBUF_16%X
x_PM_SKY130_FD_SC_HDLL__CLKBUF_16%VGND N_VGND_M1006_s N_VGND_M1007_s
+ N_VGND_M1023_s N_VGND_M1001_d N_VGND_M1005_d N_VGND_M1017_d N_VGND_M1020_d
+ N_VGND_M1024_d N_VGND_M1032_d N_VGND_M1036_d N_VGND_M1039_d N_VGND_c_851_n
+ N_VGND_c_852_n N_VGND_c_853_n N_VGND_c_854_n N_VGND_c_855_n N_VGND_c_856_n
+ N_VGND_c_857_n N_VGND_c_858_n N_VGND_c_859_n N_VGND_c_860_n N_VGND_c_861_n
+ N_VGND_c_862_n N_VGND_c_863_n N_VGND_c_864_n N_VGND_c_865_n N_VGND_c_866_n
+ N_VGND_c_867_n N_VGND_c_868_n N_VGND_c_869_n N_VGND_c_870_n N_VGND_c_871_n
+ N_VGND_c_872_n N_VGND_c_873_n N_VGND_c_874_n N_VGND_c_875_n N_VGND_c_876_n
+ N_VGND_c_877_n N_VGND_c_878_n N_VGND_c_879_n VGND N_VGND_c_880_n
+ N_VGND_c_881_n N_VGND_c_882_n N_VGND_c_883_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_16%VGND
cc_1 VNB N_A_M1006_g 0.0301185f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.445
cc_2 VNB N_A_M1007_g 0.0244402f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=0.445
cc_3 VNB N_A_M1011_g 0.0244401f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=0.445
cc_4 VNB N_A_M1023_g 0.0241662f $X=-0.19 $Y=-0.24 $X2=1.965 $Y2=0.445
cc_5 VNB A 0.023702f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_6 VNB N_A_c_149_n 0.125209f $X=-0.19 $Y=-0.24 $X2=1.965 $Y2=1.155
cc_7 VNB N_A_118_297#_M1000_g 0.0268891f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.41
cc_8 VNB N_A_118_297#_M1001_g 0.0258077f $X=-0.19 $Y=-0.24 $X2=1.94 $Y2=1.41
cc_9 VNB N_A_118_297#_M1002_g 0.0258075f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_10 VNB N_A_118_297#_M1005_g 0.0258077f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_118_297#_M1012_g 0.0258075f $X=-0.19 $Y=-0.24 $X2=1.94 $Y2=1.155
cc_12 VNB N_A_118_297#_M1017_g 0.0258057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_118_297#_M1019_g 0.0254848f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_118_297#_M1020_g 0.0257277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_118_297#_M1021_g 0.0257274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_118_297#_M1024_g 0.0258076f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_118_297#_M1027_g 0.0258074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_118_297#_M1032_g 0.0258076f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_118_297#_M1033_g 0.0258074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_118_297#_M1036_g 0.0258078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_118_297#_M1037_g 0.0261948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_118_297#_M1039_g 0.033665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_118_297#_c_224_n 0.00481185f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_118_297#_c_225_n 0.00524031f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_118_297#_c_226_n 0.00429043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_118_297#_c_227_n 0.349639f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_485_n 0.421552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_X_c_631_n 0.0017582f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_X_c_632_n 0.00733625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_X_c_633_n 0.00426583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_X_c_634_n 0.00149815f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_X_c_635_n 0.00733625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_X_c_636_n 0.00140668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_X_c_637_n 0.00603057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_X_c_638_n 7.61769e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_X_c_639_n 0.00708778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_X_c_640_n 0.00148721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_X_c_641_n 0.00739565f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_X_c_642_n 0.00148721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_X_c_643_n 0.00739565f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_X_c_644_n 0.00202124f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_X_c_645_n 0.00148721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_X_c_646_n 0.0015723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_X_c_647_n 0.0018976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_X_c_648_n 0.0018976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_X_c_649_n 0.0024696f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_X_c_650_n 0.0018976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_X_c_651_n 0.0018976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_X_c_652_n 0.0018976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB X 0.0329822f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_851_n 0.0107531f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_52 VNB N_VGND_c_852_n 0.0196988f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_853_n 0.0199238f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.155
cc_54 VNB N_VGND_c_854_n 0.00523594f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=1.155
cc_55 VNB N_VGND_c_855_n 0.0199238f $X=-0.19 $Y=-0.24 $X2=1.965 $Y2=1.155
cc_56 VNB N_VGND_c_856_n 0.00522139f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_857_n 0.00523594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_858_n 0.00523594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_859_n 0.00511236f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_860_n 0.00515183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_861_n 0.00518f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_862_n 0.00518f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_863_n 0.00523594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_864_n 0.0109745f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_865_n 0.0184458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_866_n 0.0190904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_867_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_868_n 0.0182806f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_869_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_870_n 0.0182806f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_871_n 0.0046855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_872_n 0.0183422f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_873_n 0.0046855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_874_n 0.0185624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_875_n 0.00478165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_876_n 0.0185624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_877_n 0.00478165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_878_n 0.0185258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_879_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_880_n 0.0182774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_881_n 0.00497572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_882_n 0.00500104f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_883_n 0.465174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VPB N_A_c_150_n 0.0211429f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_85 VPB N_A_c_151_n 0.0163977f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.41
cc_86 VPB N_A_c_152_n 0.0163977f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.41
cc_87 VPB N_A_c_153_n 0.0165782f $X=-0.19 $Y=1.305 $X2=1.94 $Y2=1.41
cc_88 VPB A 0.00127249f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_89 VPB N_A_c_149_n 0.0494902f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=1.155
cc_90 VPB N_A_118_297#_c_228_n 0.0166021f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.985
cc_91 VPB N_A_118_297#_c_229_n 0.0164285f $X=-0.19 $Y=1.305 $X2=1.94 $Y2=1.985
cc_92 VPB N_A_118_297#_c_230_n 0.0164285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_118_297#_c_231_n 0.0164285f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.155
cc_94 VPB N_A_118_297#_c_232_n 0.0164285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_118_297#_c_233_n 0.0164285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_118_297#_c_234_n 0.0164285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_118_297#_c_235_n 0.0163875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_118_297#_c_236_n 0.0163875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_118_297#_c_237_n 0.0164285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_118_297#_c_238_n 0.0164285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_118_297#_c_239_n 0.0164285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_118_297#_c_240_n 0.0164269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_118_297#_c_241_n 0.0164158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_118_297#_c_242_n 0.0157624f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_118_297#_c_243_n 0.0193677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_118_297#_c_244_n 0.00139844f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_118_297#_c_245_n 0.00140153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_118_297#_c_226_n 0.00459688f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_118_297#_c_227_n 0.209766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_486_n 0.0108797f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_111 VPB N_VPWR_c_487_n 0.0309762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_488_n 0.0199257f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.155
cc_113 VPB N_VPWR_c_489_n 0.00522213f $X=-0.19 $Y=1.305 $X2=1.485 $Y2=1.155
cc_114 VPB N_VPWR_c_490_n 0.0199013f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=1.155
cc_115 VPB N_VPWR_c_491_n 0.00504594f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_492_n 0.00504594f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_493_n 0.00504594f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_494_n 0.00504594f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_495_n 0.00496467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_496_n 0.00496485f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_497_n 0.00496485f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_498_n 0.00501892f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_499_n 0.0103988f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_500_n 0.0281929f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_501_n 0.0199172f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_502_n 0.00502323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_503_n 0.0199172f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_504_n 0.00502323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_505_n 0.0199172f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_506_n 0.00502323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_507_n 0.0199172f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_508_n 0.00473193f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_509_n 0.0203974f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_510_n 0.00473193f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_511_n 0.0203974f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_512_n 0.00473193f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_513_n 0.0203974f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_514_n 0.00499086f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_515_n 0.0204288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_516_n 0.00497514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_517_n 0.00508796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_485_n 0.0439962f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB X 0.0198539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 N_A_M1023_g N_A_118_297#_M1000_g 0.0220223f $X=1.965 $Y=0.445 $X2=0 $Y2=0
cc_145 N_A_c_153_n N_A_118_297#_c_228_n 0.0221268f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_M1006_g N_A_118_297#_c_224_n 0.00434374f $X=0.525 $Y=0.445 $X2=0
+ $Y2=0
cc_147 N_A_M1007_g N_A_118_297#_c_224_n 0.00875058f $X=1.005 $Y=0.445 $X2=0
+ $Y2=0
cc_148 A N_A_118_297#_c_224_n 0.0195449f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_149 N_A_c_149_n N_A_118_297#_c_224_n 0.0184072f $X=1.965 $Y=1.155 $X2=0 $Y2=0
cc_150 N_A_c_150_n N_A_118_297#_c_244_n 0.00336448f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_c_151_n N_A_118_297#_c_244_n 0.00339176f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_c_149_n N_A_118_297#_c_244_n 0.0124529f $X=1.965 $Y=1.155 $X2=0 $Y2=0
cc_153 N_A_c_149_n N_A_118_297#_c_257_n 0.0686685f $X=1.965 $Y=1.155 $X2=0 $Y2=0
cc_154 N_A_M1011_g N_A_118_297#_c_225_n 0.00680043f $X=1.485 $Y=0.445 $X2=0
+ $Y2=0
cc_155 N_A_M1023_g N_A_118_297#_c_225_n 0.00813566f $X=1.965 $Y=0.445 $X2=0
+ $Y2=0
cc_156 N_A_c_149_n N_A_118_297#_c_225_n 0.0186314f $X=1.965 $Y=1.155 $X2=0 $Y2=0
cc_157 N_A_c_152_n N_A_118_297#_c_245_n 0.00320023f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_c_153_n N_A_118_297#_c_245_n 0.00325155f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_c_149_n N_A_118_297#_c_245_n 0.0102852f $X=1.965 $Y=1.155 $X2=0 $Y2=0
cc_160 N_A_c_149_n N_A_118_297#_c_226_n 0.027109f $X=1.965 $Y=1.155 $X2=0 $Y2=0
cc_161 A N_A_118_297#_c_265_n 0.0161665f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_162 N_A_c_149_n N_A_118_297#_c_265_n 0.0100412f $X=1.965 $Y=1.155 $X2=0 $Y2=0
cc_163 N_A_c_149_n N_A_118_297#_c_267_n 0.00588528f $X=1.965 $Y=1.155 $X2=0
+ $Y2=0
cc_164 N_A_c_149_n N_A_118_297#_c_227_n 0.0220223f $X=1.965 $Y=1.155 $X2=0 $Y2=0
cc_165 N_A_c_150_n N_VPWR_c_487_n 0.00484201f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_166 A N_VPWR_c_487_n 0.0102593f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_167 N_A_c_149_n N_VPWR_c_487_n 0.00616128f $X=1.965 $Y=1.155 $X2=0 $Y2=0
cc_168 N_A_c_150_n N_VPWR_c_488_n 0.00702461f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_c_151_n N_VPWR_c_488_n 0.00702461f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_c_151_n N_VPWR_c_489_n 0.00303578f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_c_152_n N_VPWR_c_489_n 0.00303578f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A_c_149_n N_VPWR_c_489_n 0.00269579f $X=1.965 $Y=1.155 $X2=0 $Y2=0
cc_173 N_A_c_152_n N_VPWR_c_490_n 0.00702461f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_c_153_n N_VPWR_c_490_n 0.00702461f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_c_153_n N_VPWR_c_491_n 0.00303578f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A_c_150_n N_VPWR_c_485_n 0.0133506f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A_c_151_n N_VPWR_c_485_n 0.0124599f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A_c_152_n N_VPWR_c_485_n 0.0125388f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_c_153_n N_VPWR_c_485_n 0.0125621f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_M1006_g N_VGND_c_852_n 0.00683213f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_181 A N_VGND_c_852_n 0.0266668f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_182 N_A_c_149_n N_VGND_c_852_n 0.00159897f $X=1.965 $Y=1.155 $X2=0 $Y2=0
cc_183 N_A_M1006_g N_VGND_c_853_n 0.00585385f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_184 N_A_M1007_g N_VGND_c_853_n 0.00585385f $X=1.005 $Y=0.445 $X2=0 $Y2=0
cc_185 N_A_M1007_g N_VGND_c_854_n 0.00320795f $X=1.005 $Y=0.445 $X2=0 $Y2=0
cc_186 N_A_M1011_g N_VGND_c_854_n 0.0048757f $X=1.485 $Y=0.445 $X2=0 $Y2=0
cc_187 N_A_c_149_n N_VGND_c_854_n 0.00390083f $X=1.965 $Y=1.155 $X2=0 $Y2=0
cc_188 N_A_M1011_g N_VGND_c_855_n 0.00585385f $X=1.485 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A_M1023_g N_VGND_c_855_n 0.00585385f $X=1.965 $Y=0.445 $X2=0 $Y2=0
cc_190 N_A_M1023_g N_VGND_c_856_n 0.00313954f $X=1.965 $Y=0.445 $X2=0 $Y2=0
cc_191 N_A_M1006_g N_VGND_c_883_n 0.0117978f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_192 N_A_M1007_g N_VGND_c_883_n 0.0109017f $X=1.005 $Y=0.445 $X2=0 $Y2=0
cc_193 N_A_M1011_g N_VGND_c_883_n 0.0110272f $X=1.485 $Y=0.445 $X2=0 $Y2=0
cc_194 N_A_M1023_g N_VGND_c_883_n 0.0107987f $X=1.965 $Y=0.445 $X2=0 $Y2=0
cc_195 A N_VGND_c_883_n 0.00161553f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_196 N_A_118_297#_c_244_n N_VPWR_c_488_n 0.0151021f $X=0.74 $Y=1.96 $X2=0
+ $Y2=0
cc_197 N_A_118_297#_c_257_n N_VPWR_c_489_n 0.00759905f $X=1.58 $Y=1.2 $X2=0
+ $Y2=0
cc_198 N_A_118_297#_c_245_n N_VPWR_c_490_n 0.0148098f $X=1.7 $Y=1.92 $X2=0 $Y2=0
cc_199 N_A_118_297#_c_228_n N_VPWR_c_491_n 0.00303578f $X=2.42 $Y=1.41 $X2=0
+ $Y2=0
cc_200 N_A_118_297#_c_226_n N_VPWR_c_491_n 0.00850896f $X=8.305 $Y=1.16 $X2=0
+ $Y2=0
cc_201 N_A_118_297#_c_229_n N_VPWR_c_492_n 0.00398486f $X=2.9 $Y=1.41 $X2=0
+ $Y2=0
cc_202 N_A_118_297#_c_230_n N_VPWR_c_492_n 0.00398486f $X=3.38 $Y=1.41 $X2=0
+ $Y2=0
cc_203 N_A_118_297#_c_231_n N_VPWR_c_493_n 0.00398486f $X=3.86 $Y=1.41 $X2=0
+ $Y2=0
cc_204 N_A_118_297#_c_232_n N_VPWR_c_493_n 0.00398486f $X=4.34 $Y=1.41 $X2=0
+ $Y2=0
cc_205 N_A_118_297#_c_233_n N_VPWR_c_494_n 0.00398486f $X=4.82 $Y=1.41 $X2=0
+ $Y2=0
cc_206 N_A_118_297#_c_234_n N_VPWR_c_494_n 0.00398486f $X=5.3 $Y=1.41 $X2=0
+ $Y2=0
cc_207 N_A_118_297#_c_235_n N_VPWR_c_495_n 0.0039448f $X=5.78 $Y=1.41 $X2=0
+ $Y2=0
cc_208 N_A_118_297#_c_236_n N_VPWR_c_495_n 0.00386731f $X=6.255 $Y=1.41 $X2=0
+ $Y2=0
cc_209 N_A_118_297#_c_237_n N_VPWR_c_496_n 0.00392752f $X=6.735 $Y=1.41 $X2=0
+ $Y2=0
cc_210 N_A_118_297#_c_238_n N_VPWR_c_496_n 0.00388876f $X=7.215 $Y=1.41 $X2=0
+ $Y2=0
cc_211 N_A_118_297#_c_239_n N_VPWR_c_497_n 0.00392752f $X=7.695 $Y=1.41 $X2=0
+ $Y2=0
cc_212 N_A_118_297#_c_240_n N_VPWR_c_497_n 0.00388876f $X=8.175 $Y=1.41 $X2=0
+ $Y2=0
cc_213 N_A_118_297#_c_241_n N_VPWR_c_498_n 0.00393961f $X=8.655 $Y=1.41 $X2=0
+ $Y2=0
cc_214 N_A_118_297#_c_242_n N_VPWR_c_498_n 0.00397892f $X=9.135 $Y=1.41 $X2=0
+ $Y2=0
cc_215 N_A_118_297#_c_227_n N_VPWR_c_498_n 7.89682e-19 $X=9.615 $Y=1.18 $X2=0
+ $Y2=0
cc_216 N_A_118_297#_c_243_n N_VPWR_c_500_n 0.00866749f $X=9.615 $Y=1.41 $X2=0
+ $Y2=0
cc_217 N_A_118_297#_c_228_n N_VPWR_c_501_n 0.00709843f $X=2.42 $Y=1.41 $X2=0
+ $Y2=0
cc_218 N_A_118_297#_c_229_n N_VPWR_c_501_n 0.00709843f $X=2.9 $Y=1.41 $X2=0
+ $Y2=0
cc_219 N_A_118_297#_c_230_n N_VPWR_c_503_n 0.00709843f $X=3.38 $Y=1.41 $X2=0
+ $Y2=0
cc_220 N_A_118_297#_c_231_n N_VPWR_c_503_n 0.00709843f $X=3.86 $Y=1.41 $X2=0
+ $Y2=0
cc_221 N_A_118_297#_c_232_n N_VPWR_c_505_n 0.00709843f $X=4.34 $Y=1.41 $X2=0
+ $Y2=0
cc_222 N_A_118_297#_c_233_n N_VPWR_c_505_n 0.00709843f $X=4.82 $Y=1.41 $X2=0
+ $Y2=0
cc_223 N_A_118_297#_c_234_n N_VPWR_c_507_n 0.00709843f $X=5.3 $Y=1.41 $X2=0
+ $Y2=0
cc_224 N_A_118_297#_c_235_n N_VPWR_c_507_n 0.00709843f $X=5.78 $Y=1.41 $X2=0
+ $Y2=0
cc_225 N_A_118_297#_c_236_n N_VPWR_c_509_n 0.00709843f $X=6.255 $Y=1.41 $X2=0
+ $Y2=0
cc_226 N_A_118_297#_c_237_n N_VPWR_c_509_n 0.00709843f $X=6.735 $Y=1.41 $X2=0
+ $Y2=0
cc_227 N_A_118_297#_c_238_n N_VPWR_c_511_n 0.00709843f $X=7.215 $Y=1.41 $X2=0
+ $Y2=0
cc_228 N_A_118_297#_c_239_n N_VPWR_c_511_n 0.00709843f $X=7.695 $Y=1.41 $X2=0
+ $Y2=0
cc_229 N_A_118_297#_c_240_n N_VPWR_c_513_n 0.00709843f $X=8.175 $Y=1.41 $X2=0
+ $Y2=0
cc_230 N_A_118_297#_c_241_n N_VPWR_c_513_n 0.00709843f $X=8.655 $Y=1.41 $X2=0
+ $Y2=0
cc_231 N_A_118_297#_c_242_n N_VPWR_c_515_n 0.00702461f $X=9.135 $Y=1.41 $X2=0
+ $Y2=0
cc_232 N_A_118_297#_c_243_n N_VPWR_c_515_n 0.00688861f $X=9.615 $Y=1.41 $X2=0
+ $Y2=0
cc_233 N_A_118_297#_M1013_d N_VPWR_c_485_n 0.00430227f $X=0.59 $Y=1.485 $X2=0
+ $Y2=0
cc_234 N_A_118_297#_M1030_d N_VPWR_c_485_n 0.00421554f $X=1.55 $Y=1.485 $X2=0
+ $Y2=0
cc_235 N_A_118_297#_c_228_n N_VPWR_c_485_n 0.0125397f $X=2.42 $Y=1.41 $X2=0
+ $Y2=0
cc_236 N_A_118_297#_c_229_n N_VPWR_c_485_n 0.0125948f $X=2.9 $Y=1.41 $X2=0 $Y2=0
cc_237 N_A_118_297#_c_230_n N_VPWR_c_485_n 0.0125948f $X=3.38 $Y=1.41 $X2=0
+ $Y2=0
cc_238 N_A_118_297#_c_231_n N_VPWR_c_485_n 0.0125948f $X=3.86 $Y=1.41 $X2=0
+ $Y2=0
cc_239 N_A_118_297#_c_232_n N_VPWR_c_485_n 0.0125948f $X=4.34 $Y=1.41 $X2=0
+ $Y2=0
cc_240 N_A_118_297#_c_233_n N_VPWR_c_485_n 0.0125948f $X=4.82 $Y=1.41 $X2=0
+ $Y2=0
cc_241 N_A_118_297#_c_234_n N_VPWR_c_485_n 0.0125948f $X=5.3 $Y=1.41 $X2=0 $Y2=0
cc_242 N_A_118_297#_c_235_n N_VPWR_c_485_n 0.0125817f $X=5.78 $Y=1.41 $X2=0
+ $Y2=0
cc_243 N_A_118_297#_c_236_n N_VPWR_c_485_n 0.0126045f $X=6.255 $Y=1.41 $X2=0
+ $Y2=0
cc_244 N_A_118_297#_c_237_n N_VPWR_c_485_n 0.0126062f $X=6.735 $Y=1.41 $X2=0
+ $Y2=0
cc_245 N_A_118_297#_c_238_n N_VPWR_c_485_n 0.0126177f $X=7.215 $Y=1.41 $X2=0
+ $Y2=0
cc_246 N_A_118_297#_c_239_n N_VPWR_c_485_n 0.0126062f $X=7.695 $Y=1.41 $X2=0
+ $Y2=0
cc_247 N_A_118_297#_c_240_n N_VPWR_c_485_n 0.0126177f $X=8.175 $Y=1.41 $X2=0
+ $Y2=0
cc_248 N_A_118_297#_c_241_n N_VPWR_c_485_n 0.0126062f $X=8.655 $Y=1.41 $X2=0
+ $Y2=0
cc_249 N_A_118_297#_c_242_n N_VPWR_c_485_n 0.0126172f $X=9.135 $Y=1.41 $X2=0
+ $Y2=0
cc_250 N_A_118_297#_c_243_n N_VPWR_c_485_n 0.0132896f $X=9.615 $Y=1.41 $X2=0
+ $Y2=0
cc_251 N_A_118_297#_c_244_n N_VPWR_c_485_n 0.00935836f $X=0.74 $Y=1.96 $X2=0
+ $Y2=0
cc_252 N_A_118_297#_c_245_n N_VPWR_c_485_n 0.00952853f $X=1.7 $Y=1.92 $X2=0
+ $Y2=0
cc_253 N_A_118_297#_M1000_g N_X_c_631_n 0.00377354f $X=2.395 $Y=0.445 $X2=0
+ $Y2=0
cc_254 N_A_118_297#_M1001_g N_X_c_631_n 0.00228345f $X=2.875 $Y=0.445 $X2=0
+ $Y2=0
cc_255 N_A_118_297#_M1001_g N_X_c_632_n 0.0124132f $X=2.875 $Y=0.445 $X2=0 $Y2=0
cc_256 N_A_118_297#_M1002_g N_X_c_632_n 0.0128559f $X=3.355 $Y=0.445 $X2=0 $Y2=0
cc_257 N_A_118_297#_c_226_n N_X_c_632_n 0.0503195f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_258 N_A_118_297#_c_227_n N_X_c_632_n 0.00400618f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_259 N_A_118_297#_M1000_g N_X_c_633_n 0.00545572f $X=2.395 $Y=0.445 $X2=0
+ $Y2=0
cc_260 N_A_118_297#_c_226_n N_X_c_633_n 0.021367f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A_118_297#_c_227_n N_X_c_633_n 0.00415703f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_262 N_A_118_297#_c_229_n N_X_c_664_n 0.017751f $X=2.9 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A_118_297#_c_230_n N_X_c_664_n 0.017751f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A_118_297#_c_226_n N_X_c_664_n 0.0450774f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_265 N_A_118_297#_c_227_n N_X_c_664_n 0.00670724f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_266 N_A_118_297#_M1002_g N_X_c_634_n 0.00519179f $X=3.355 $Y=0.445 $X2=0
+ $Y2=0
cc_267 N_A_118_297#_M1005_g N_X_c_634_n 0.00228345f $X=3.835 $Y=0.445 $X2=0
+ $Y2=0
cc_268 N_A_118_297#_M1005_g N_X_c_635_n 0.0128559f $X=3.835 $Y=0.445 $X2=0 $Y2=0
cc_269 N_A_118_297#_M1012_g N_X_c_635_n 0.0128559f $X=4.315 $Y=0.445 $X2=0 $Y2=0
cc_270 N_A_118_297#_c_226_n N_X_c_635_n 0.0503195f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_271 N_A_118_297#_c_227_n N_X_c_635_n 0.00400618f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_272 N_A_118_297#_c_231_n N_X_c_674_n 0.017751f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_273 N_A_118_297#_c_232_n N_X_c_674_n 0.017751f $X=4.34 $Y=1.41 $X2=0 $Y2=0
cc_274 N_A_118_297#_c_226_n N_X_c_674_n 0.0450774f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_275 N_A_118_297#_c_227_n N_X_c_674_n 0.00670724f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_276 N_A_118_297#_M1012_g N_X_c_636_n 0.00519179f $X=4.315 $Y=0.445 $X2=0
+ $Y2=0
cc_277 N_A_118_297#_M1017_g N_X_c_636_n 0.00130218f $X=4.795 $Y=0.445 $X2=0
+ $Y2=0
cc_278 N_A_118_297#_M1017_g N_X_c_637_n 0.0128559f $X=4.795 $Y=0.445 $X2=0 $Y2=0
cc_279 N_A_118_297#_M1019_g N_X_c_637_n 0.0102303f $X=5.275 $Y=0.445 $X2=0 $Y2=0
cc_280 N_A_118_297#_c_226_n N_X_c_637_n 0.0455574f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_281 N_A_118_297#_c_227_n N_X_c_637_n 0.00400618f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_282 N_A_118_297#_c_233_n N_X_c_684_n 0.017751f $X=4.82 $Y=1.41 $X2=0 $Y2=0
cc_283 N_A_118_297#_c_234_n N_X_c_684_n 0.017751f $X=5.3 $Y=1.41 $X2=0 $Y2=0
cc_284 N_A_118_297#_c_226_n N_X_c_684_n 0.0450774f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_285 N_A_118_297#_c_227_n N_X_c_684_n 0.00670724f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_286 N_A_118_297#_M1017_g N_X_c_638_n 5.07314e-19 $X=4.795 $Y=0.445 $X2=0
+ $Y2=0
cc_287 N_A_118_297#_M1019_g N_X_c_638_n 0.00667092f $X=5.275 $Y=0.445 $X2=0
+ $Y2=0
cc_288 N_A_118_297#_M1020_g N_X_c_638_n 0.00237691f $X=5.755 $Y=0.445 $X2=0
+ $Y2=0
cc_289 N_A_118_297#_M1020_g N_X_c_639_n 0.0128288f $X=5.755 $Y=0.445 $X2=0 $Y2=0
cc_290 N_A_118_297#_M1021_g N_X_c_639_n 0.0128288f $X=6.23 $Y=0.445 $X2=0 $Y2=0
cc_291 N_A_118_297#_c_226_n N_X_c_639_n 0.0492155f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_292 N_A_118_297#_c_227_n N_X_c_639_n 0.00387264f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_293 N_A_118_297#_c_235_n N_X_c_695_n 0.0177094f $X=5.78 $Y=1.41 $X2=0 $Y2=0
cc_294 N_A_118_297#_c_236_n N_X_c_695_n 0.0177094f $X=6.255 $Y=1.41 $X2=0 $Y2=0
cc_295 N_A_118_297#_c_226_n N_X_c_695_n 0.0443468f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_296 N_A_118_297#_c_227_n N_X_c_695_n 0.00659124f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_297 N_A_118_297#_M1021_g N_X_c_640_n 0.0021663f $X=6.23 $Y=0.445 $X2=0 $Y2=0
cc_298 N_A_118_297#_M1024_g N_X_c_640_n 0.0022534f $X=6.71 $Y=0.445 $X2=0 $Y2=0
cc_299 N_A_118_297#_M1024_g N_X_c_641_n 0.0128559f $X=6.71 $Y=0.445 $X2=0 $Y2=0
cc_300 N_A_118_297#_M1027_g N_X_c_641_n 0.0128559f $X=7.19 $Y=0.445 $X2=0 $Y2=0
cc_301 N_A_118_297#_c_226_n N_X_c_641_n 0.0503195f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_302 N_A_118_297#_c_227_n N_X_c_641_n 0.00400618f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_303 N_A_118_297#_c_237_n N_X_c_705_n 0.017751f $X=6.735 $Y=1.41 $X2=0 $Y2=0
cc_304 N_A_118_297#_c_238_n N_X_c_705_n 0.017751f $X=7.215 $Y=1.41 $X2=0 $Y2=0
cc_305 N_A_118_297#_c_226_n N_X_c_705_n 0.0450774f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_306 N_A_118_297#_c_227_n N_X_c_705_n 0.00670724f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_307 N_A_118_297#_M1027_g N_X_c_642_n 0.0021663f $X=7.19 $Y=0.445 $X2=0 $Y2=0
cc_308 N_A_118_297#_M1032_g N_X_c_642_n 0.0022534f $X=7.67 $Y=0.445 $X2=0 $Y2=0
cc_309 N_A_118_297#_M1032_g N_X_c_643_n 0.0128559f $X=7.67 $Y=0.445 $X2=0 $Y2=0
cc_310 N_A_118_297#_M1033_g N_X_c_643_n 0.0128559f $X=8.15 $Y=0.445 $X2=0 $Y2=0
cc_311 N_A_118_297#_c_226_n N_X_c_643_n 0.0503195f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_312 N_A_118_297#_c_227_n N_X_c_643_n 0.00400618f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_313 N_A_118_297#_c_239_n N_X_c_644_n 0.017751f $X=7.695 $Y=1.41 $X2=0 $Y2=0
cc_314 N_A_118_297#_c_240_n N_X_c_644_n 0.017751f $X=8.175 $Y=1.41 $X2=0 $Y2=0
cc_315 N_A_118_297#_M1036_g N_X_c_644_n 0.0147462f $X=8.63 $Y=0.445 $X2=0 $Y2=0
cc_316 N_A_118_297#_c_226_n N_X_c_644_n 0.0454078f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_317 N_A_118_297#_c_227_n N_X_c_644_n 0.00670724f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_318 N_A_118_297#_M1033_g N_X_c_645_n 0.0021663f $X=8.15 $Y=0.445 $X2=0 $Y2=0
cc_319 N_A_118_297#_M1036_g N_X_c_645_n 0.0022534f $X=8.63 $Y=0.445 $X2=0 $Y2=0
cc_320 N_A_118_297#_M1037_g N_X_c_646_n 0.00525012f $X=9.11 $Y=0.445 $X2=0 $Y2=0
cc_321 N_A_118_297#_M1039_g N_X_c_646_n 0.00525012f $X=9.64 $Y=0.445 $X2=0 $Y2=0
cc_322 N_A_118_297#_c_226_n N_X_c_724_n 0.0177415f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_323 N_A_118_297#_c_227_n N_X_c_724_n 0.00635512f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_324 N_A_118_297#_c_226_n N_X_c_647_n 0.021367f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_325 N_A_118_297#_c_227_n N_X_c_647_n 0.00415703f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_326 N_A_118_297#_c_226_n N_X_c_728_n 0.0177415f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_327 N_A_118_297#_c_227_n N_X_c_728_n 0.00635512f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_328 N_A_118_297#_c_226_n N_X_c_648_n 0.021367f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A_118_297#_c_227_n N_X_c_648_n 0.00415703f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_330 N_A_118_297#_c_226_n N_X_c_732_n 0.0177415f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_331 N_A_118_297#_c_227_n N_X_c_732_n 0.00635512f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_332 N_A_118_297#_M1019_g N_X_c_649_n 0.00240228f $X=5.275 $Y=0.445 $X2=0
+ $Y2=0
cc_333 N_A_118_297#_c_226_n N_X_c_649_n 0.0266872f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_334 N_A_118_297#_c_227_n N_X_c_649_n 0.00415703f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_335 N_A_118_297#_c_226_n N_X_c_737_n 0.0177415f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A_118_297#_c_227_n N_X_c_737_n 0.00635512f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_337 N_A_118_297#_c_226_n N_X_c_650_n 0.021367f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_338 N_A_118_297#_c_227_n N_X_c_650_n 0.00415703f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_339 N_A_118_297#_c_226_n N_X_c_741_n 0.0177415f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_340 N_A_118_297#_c_227_n N_X_c_741_n 0.00635512f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_341 N_A_118_297#_c_226_n N_X_c_651_n 0.021367f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_342 N_A_118_297#_c_227_n N_X_c_651_n 0.00415703f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_343 N_A_118_297#_c_226_n N_X_c_745_n 0.0177415f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_344 N_A_118_297#_c_227_n N_X_c_745_n 0.00635512f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_345 N_A_118_297#_c_226_n N_X_c_652_n 0.021367f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_346 N_A_118_297#_c_227_n N_X_c_652_n 0.00415703f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_347 N_A_118_297#_c_241_n X 0.0207323f $X=8.655 $Y=1.41 $X2=0 $Y2=0
cc_348 N_A_118_297#_M1037_g X 0.0130265f $X=9.11 $Y=0.445 $X2=0 $Y2=0
cc_349 N_A_118_297#_c_242_n X 0.0194145f $X=9.135 $Y=1.41 $X2=0 $Y2=0
cc_350 N_A_118_297#_c_243_n X 0.0214176f $X=9.615 $Y=1.41 $X2=0 $Y2=0
cc_351 N_A_118_297#_M1039_g X 0.014443f $X=9.64 $Y=0.445 $X2=0 $Y2=0
cc_352 N_A_118_297#_c_226_n X 0.0349671f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_353 N_A_118_297#_c_227_n X 0.0905049f $X=9.615 $Y=1.18 $X2=0 $Y2=0
cc_354 N_A_118_297#_c_243_n N_X_c_756_n 0.0157494f $X=9.615 $Y=1.41 $X2=0 $Y2=0
cc_355 N_A_118_297#_c_224_n N_VGND_c_853_n 0.0152148f $X=0.74 $Y=0.445 $X2=0
+ $Y2=0
cc_356 N_A_118_297#_c_257_n N_VGND_c_854_n 0.00863012f $X=1.58 $Y=1.2 $X2=0
+ $Y2=0
cc_357 N_A_118_297#_c_225_n N_VGND_c_855_n 0.0152148f $X=1.7 $Y=0.445 $X2=0
+ $Y2=0
cc_358 N_A_118_297#_M1000_g N_VGND_c_856_n 0.00313954f $X=2.395 $Y=0.445 $X2=0
+ $Y2=0
cc_359 N_A_118_297#_c_226_n N_VGND_c_856_n 0.0091835f $X=8.305 $Y=1.16 $X2=0
+ $Y2=0
cc_360 N_A_118_297#_M1001_g N_VGND_c_857_n 0.00484691f $X=2.875 $Y=0.445 $X2=0
+ $Y2=0
cc_361 N_A_118_297#_M1002_g N_VGND_c_857_n 0.00313102f $X=3.355 $Y=0.445 $X2=0
+ $Y2=0
cc_362 N_A_118_297#_M1005_g N_VGND_c_858_n 0.00484691f $X=3.835 $Y=0.445 $X2=0
+ $Y2=0
cc_363 N_A_118_297#_M1012_g N_VGND_c_858_n 0.00313102f $X=4.315 $Y=0.445 $X2=0
+ $Y2=0
cc_364 N_A_118_297#_M1017_g N_VGND_c_859_n 0.0048031f $X=4.795 $Y=0.445 $X2=0
+ $Y2=0
cc_365 N_A_118_297#_M1019_g N_VGND_c_859_n 0.00302263f $X=5.275 $Y=0.445 $X2=0
+ $Y2=0
cc_366 N_A_118_297#_M1020_g N_VGND_c_860_n 0.00479609f $X=5.755 $Y=0.445 $X2=0
+ $Y2=0
cc_367 N_A_118_297#_M1021_g N_VGND_c_860_n 0.00304452f $X=6.23 $Y=0.445 $X2=0
+ $Y2=0
cc_368 N_A_118_297#_M1024_g N_VGND_c_861_n 0.00486187f $X=6.71 $Y=0.445 $X2=0
+ $Y2=0
cc_369 N_A_118_297#_M1027_g N_VGND_c_861_n 0.00305844f $X=7.19 $Y=0.445 $X2=0
+ $Y2=0
cc_370 N_A_118_297#_M1032_g N_VGND_c_862_n 0.00486187f $X=7.67 $Y=0.445 $X2=0
+ $Y2=0
cc_371 N_A_118_297#_M1033_g N_VGND_c_862_n 0.00305844f $X=8.15 $Y=0.445 $X2=0
+ $Y2=0
cc_372 N_A_118_297#_M1036_g N_VGND_c_863_n 0.00489124f $X=8.63 $Y=0.445 $X2=0
+ $Y2=0
cc_373 N_A_118_297#_M1037_g N_VGND_c_863_n 0.00313102f $X=9.11 $Y=0.445 $X2=0
+ $Y2=0
cc_374 N_A_118_297#_c_227_n N_VGND_c_863_n 7.1871e-19 $X=9.615 $Y=1.18 $X2=0
+ $Y2=0
cc_375 N_A_118_297#_M1039_g N_VGND_c_865_n 0.00488085f $X=9.64 $Y=0.445 $X2=0
+ $Y2=0
cc_376 N_A_118_297#_M1000_g N_VGND_c_866_n 0.00585385f $X=2.395 $Y=0.445 $X2=0
+ $Y2=0
cc_377 N_A_118_297#_M1001_g N_VGND_c_866_n 0.00439206f $X=2.875 $Y=0.445 $X2=0
+ $Y2=0
cc_378 N_A_118_297#_M1002_g N_VGND_c_868_n 0.00439206f $X=3.355 $Y=0.445 $X2=0
+ $Y2=0
cc_379 N_A_118_297#_M1005_g N_VGND_c_868_n 0.00439206f $X=3.835 $Y=0.445 $X2=0
+ $Y2=0
cc_380 N_A_118_297#_M1012_g N_VGND_c_870_n 0.00439206f $X=4.315 $Y=0.445 $X2=0
+ $Y2=0
cc_381 N_A_118_297#_M1017_g N_VGND_c_870_n 0.00439206f $X=4.795 $Y=0.445 $X2=0
+ $Y2=0
cc_382 N_A_118_297#_M1019_g N_VGND_c_872_n 0.00438144f $X=5.275 $Y=0.445 $X2=0
+ $Y2=0
cc_383 N_A_118_297#_M1020_g N_VGND_c_872_n 0.00439206f $X=5.755 $Y=0.445 $X2=0
+ $Y2=0
cc_384 N_A_118_297#_M1021_g N_VGND_c_874_n 0.00439206f $X=6.23 $Y=0.445 $X2=0
+ $Y2=0
cc_385 N_A_118_297#_M1024_g N_VGND_c_874_n 0.00439206f $X=6.71 $Y=0.445 $X2=0
+ $Y2=0
cc_386 N_A_118_297#_M1027_g N_VGND_c_876_n 0.00439206f $X=7.19 $Y=0.445 $X2=0
+ $Y2=0
cc_387 N_A_118_297#_M1032_g N_VGND_c_876_n 0.00439206f $X=7.67 $Y=0.445 $X2=0
+ $Y2=0
cc_388 N_A_118_297#_M1033_g N_VGND_c_878_n 0.00439206f $X=8.15 $Y=0.445 $X2=0
+ $Y2=0
cc_389 N_A_118_297#_M1036_g N_VGND_c_878_n 0.00439206f $X=8.63 $Y=0.445 $X2=0
+ $Y2=0
cc_390 N_A_118_297#_M1037_g N_VGND_c_880_n 0.00439071f $X=9.11 $Y=0.445 $X2=0
+ $Y2=0
cc_391 N_A_118_297#_M1039_g N_VGND_c_880_n 0.00439071f $X=9.64 $Y=0.445 $X2=0
+ $Y2=0
cc_392 N_A_118_297#_M1006_d N_VGND_c_883_n 0.00549964f $X=0.6 $Y=0.235 $X2=0
+ $Y2=0
cc_393 N_A_118_297#_M1011_d N_VGND_c_883_n 0.00549964f $X=1.56 $Y=0.235 $X2=0
+ $Y2=0
cc_394 N_A_118_297#_M1000_g N_VGND_c_883_n 0.0107987f $X=2.395 $Y=0.445 $X2=0
+ $Y2=0
cc_395 N_A_118_297#_M1001_g N_VGND_c_883_n 0.00628867f $X=2.875 $Y=0.445 $X2=0
+ $Y2=0
cc_396 N_A_118_297#_M1002_g N_VGND_c_883_n 0.00616322f $X=3.355 $Y=0.445 $X2=0
+ $Y2=0
cc_397 N_A_118_297#_M1005_g N_VGND_c_883_n 0.00628867f $X=3.835 $Y=0.445 $X2=0
+ $Y2=0
cc_398 N_A_118_297#_M1012_g N_VGND_c_883_n 0.00616322f $X=4.315 $Y=0.445 $X2=0
+ $Y2=0
cc_399 N_A_118_297#_M1017_g N_VGND_c_883_n 0.00628867f $X=4.795 $Y=0.445 $X2=0
+ $Y2=0
cc_400 N_A_118_297#_M1019_g N_VGND_c_883_n 0.00612682f $X=5.275 $Y=0.445 $X2=0
+ $Y2=0
cc_401 N_A_118_297#_M1020_g N_VGND_c_883_n 0.00627675f $X=5.755 $Y=0.445 $X2=0
+ $Y2=0
cc_402 N_A_118_297#_M1021_g N_VGND_c_883_n 0.00617638f $X=6.23 $Y=0.445 $X2=0
+ $Y2=0
cc_403 N_A_118_297#_M1024_g N_VGND_c_883_n 0.00628867f $X=6.71 $Y=0.445 $X2=0
+ $Y2=0
cc_404 N_A_118_297#_M1027_g N_VGND_c_883_n 0.00618831f $X=7.19 $Y=0.445 $X2=0
+ $Y2=0
cc_405 N_A_118_297#_M1032_g N_VGND_c_883_n 0.00628867f $X=7.67 $Y=0.445 $X2=0
+ $Y2=0
cc_406 N_A_118_297#_M1033_g N_VGND_c_883_n 0.00618831f $X=8.15 $Y=0.445 $X2=0
+ $Y2=0
cc_407 N_A_118_297#_M1036_g N_VGND_c_883_n 0.00628867f $X=8.63 $Y=0.445 $X2=0
+ $Y2=0
cc_408 N_A_118_297#_M1037_g N_VGND_c_883_n 0.00627824f $X=9.11 $Y=0.445 $X2=0
+ $Y2=0
cc_409 N_A_118_297#_M1039_g N_VGND_c_883_n 0.00709099f $X=9.64 $Y=0.445 $X2=0
+ $Y2=0
cc_410 N_A_118_297#_c_224_n N_VGND_c_883_n 0.00950576f $X=0.74 $Y=0.445 $X2=0
+ $Y2=0
cc_411 N_A_118_297#_c_225_n N_VGND_c_883_n 0.00950576f $X=1.7 $Y=0.445 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_485_n N_X_M1003_d 0.00386843f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_413 N_VPWR_c_485_n N_X_M1008_d 0.00386843f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_414 N_VPWR_c_485_n N_X_M1010_d 0.00386843f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_415 N_VPWR_c_485_n N_X_M1016_d 0.00386843f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_416 N_VPWR_c_485_n N_X_M1022_d 0.00386843f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_417 N_VPWR_c_485_n N_X_M1026_d 0.00386843f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_418 N_VPWR_c_485_n N_X_M1029_d 0.00386843f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_419 N_VPWR_c_485_n N_X_M1035_d 0.00313952f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_420 N_VPWR_M1004_s N_X_c_664_n 0.00357164f $X=2.99 $Y=1.485 $X2=0 $Y2=0
cc_421 N_VPWR_c_492_n N_X_c_664_n 0.0154924f $X=3.14 $Y=2.22 $X2=0 $Y2=0
cc_422 N_VPWR_M1009_s N_X_c_674_n 0.00357164f $X=3.95 $Y=1.485 $X2=0 $Y2=0
cc_423 N_VPWR_c_493_n N_X_c_674_n 0.0154924f $X=4.1 $Y=2.22 $X2=0 $Y2=0
cc_424 N_VPWR_M1015_s N_X_c_684_n 0.00357164f $X=4.91 $Y=1.485 $X2=0 $Y2=0
cc_425 N_VPWR_c_494_n N_X_c_684_n 0.0154924f $X=5.06 $Y=2.22 $X2=0 $Y2=0
cc_426 N_VPWR_M1018_s N_X_c_695_n 0.00347562f $X=5.87 $Y=1.485 $X2=0 $Y2=0
cc_427 N_VPWR_c_495_n N_X_c_695_n 0.0150759f $X=6.02 $Y=2.22 $X2=0 $Y2=0
cc_428 N_VPWR_M1025_s N_X_c_705_n 0.00357164f $X=6.825 $Y=1.485 $X2=0 $Y2=0
cc_429 N_VPWR_c_496_n N_X_c_705_n 0.0154924f $X=6.975 $Y=2.22 $X2=0 $Y2=0
cc_430 N_VPWR_M1028_s N_X_c_644_n 0.00357164f $X=7.785 $Y=1.485 $X2=0 $Y2=0
cc_431 N_VPWR_c_497_n N_X_c_644_n 0.0154924f $X=7.935 $Y=2.22 $X2=0 $Y2=0
cc_432 N_VPWR_c_513_n N_X_c_777_n 0.0156448f $X=8.77 $Y=2.717 $X2=0 $Y2=0
cc_433 N_VPWR_c_485_n N_X_c_777_n 0.00987681f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_434 N_VPWR_c_501_n N_X_c_724_n 0.0156448f $X=3.01 $Y=2.717 $X2=0 $Y2=0
cc_435 N_VPWR_c_485_n N_X_c_724_n 0.00987681f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_436 N_VPWR_c_503_n N_X_c_728_n 0.0156448f $X=3.97 $Y=2.717 $X2=0 $Y2=0
cc_437 N_VPWR_c_485_n N_X_c_728_n 0.00987681f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_438 N_VPWR_c_505_n N_X_c_732_n 0.0156448f $X=4.93 $Y=2.717 $X2=0 $Y2=0
cc_439 N_VPWR_c_485_n N_X_c_732_n 0.00987681f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_440 N_VPWR_c_507_n N_X_c_737_n 0.0156448f $X=5.89 $Y=2.717 $X2=0 $Y2=0
cc_441 N_VPWR_c_485_n N_X_c_737_n 0.00987681f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_442 N_VPWR_c_509_n N_X_c_741_n 0.0156448f $X=6.85 $Y=2.717 $X2=0 $Y2=0
cc_443 N_VPWR_c_485_n N_X_c_741_n 0.00987681f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_444 N_VPWR_c_511_n N_X_c_745_n 0.0156448f $X=7.81 $Y=2.717 $X2=0 $Y2=0
cc_445 N_VPWR_c_485_n N_X_c_745_n 0.00987681f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_446 N_VPWR_M1031_s X 0.00213384f $X=8.745 $Y=1.485 $X2=0 $Y2=0
cc_447 N_VPWR_M1038_s X 0.00359002f $X=9.705 $Y=1.485 $X2=0 $Y2=0
cc_448 N_VPWR_c_498_n X 0.0157372f $X=8.895 $Y=2.22 $X2=0 $Y2=0
cc_449 N_VPWR_c_500_n X 0.023778f $X=9.855 $Y=2.22 $X2=0 $Y2=0
cc_450 N_VPWR_c_515_n N_X_c_756_n 0.0164721f $X=9.755 $Y=2.72 $X2=0 $Y2=0
cc_451 N_VPWR_c_485_n N_X_c_756_n 0.0110241f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_452 N_X_c_632_n N_VGND_c_857_n 0.0185136f $X=3.49 $Y=0.82 $X2=0 $Y2=0
cc_453 N_X_c_635_n N_VGND_c_858_n 0.0185136f $X=4.45 $Y=0.82 $X2=0 $Y2=0
cc_454 N_X_c_637_n N_VGND_c_859_n 0.0179867f $X=5.345 $Y=0.82 $X2=0 $Y2=0
cc_455 N_X_c_639_n N_VGND_c_860_n 0.0177638f $X=6.355 $Y=0.82 $X2=0 $Y2=0
cc_456 N_X_c_641_n N_VGND_c_861_n 0.0181624f $X=7.315 $Y=0.82 $X2=0 $Y2=0
cc_457 N_X_c_643_n N_VGND_c_862_n 0.0181624f $X=8.275 $Y=0.82 $X2=0 $Y2=0
cc_458 X N_VGND_c_863_n 0.0207327f $X=9.375 $Y=0.765 $X2=0 $Y2=0
cc_459 X N_VGND_c_865_n 0.0243436f $X=9.375 $Y=0.765 $X2=0 $Y2=0
cc_460 N_X_c_631_n N_VGND_c_866_n 0.0141875f $X=2.66 $Y=0.445 $X2=0 $Y2=0
cc_461 N_X_c_632_n N_VGND_c_866_n 0.00299761f $X=3.49 $Y=0.82 $X2=0 $Y2=0
cc_462 N_X_c_632_n N_VGND_c_868_n 0.00299761f $X=3.49 $Y=0.82 $X2=0 $Y2=0
cc_463 N_X_c_634_n N_VGND_c_868_n 0.0141875f $X=3.62 $Y=0.445 $X2=0 $Y2=0
cc_464 N_X_c_635_n N_VGND_c_868_n 0.00299761f $X=4.45 $Y=0.82 $X2=0 $Y2=0
cc_465 N_X_c_635_n N_VGND_c_870_n 0.00299761f $X=4.45 $Y=0.82 $X2=0 $Y2=0
cc_466 N_X_c_636_n N_VGND_c_870_n 0.0141875f $X=4.58 $Y=0.445 $X2=0 $Y2=0
cc_467 N_X_c_637_n N_VGND_c_870_n 0.00299761f $X=5.345 $Y=0.82 $X2=0 $Y2=0
cc_468 N_X_c_637_n N_VGND_c_872_n 0.00226107f $X=5.345 $Y=0.82 $X2=0 $Y2=0
cc_469 N_X_c_638_n N_VGND_c_872_n 0.0163978f $X=5.54 $Y=0.445 $X2=0 $Y2=0
cc_470 N_X_c_639_n N_VGND_c_872_n 0.00299761f $X=6.355 $Y=0.82 $X2=0 $Y2=0
cc_471 N_X_c_639_n N_VGND_c_874_n 0.00299761f $X=6.355 $Y=0.82 $X2=0 $Y2=0
cc_472 N_X_c_640_n N_VGND_c_874_n 0.0143045f $X=6.495 $Y=0.445 $X2=0 $Y2=0
cc_473 N_X_c_641_n N_VGND_c_874_n 0.00314713f $X=7.315 $Y=0.82 $X2=0 $Y2=0
cc_474 N_X_c_641_n N_VGND_c_876_n 0.00299761f $X=7.315 $Y=0.82 $X2=0 $Y2=0
cc_475 N_X_c_642_n N_VGND_c_876_n 0.0143045f $X=7.455 $Y=0.445 $X2=0 $Y2=0
cc_476 N_X_c_643_n N_VGND_c_876_n 0.00314713f $X=8.275 $Y=0.82 $X2=0 $Y2=0
cc_477 N_X_c_643_n N_VGND_c_878_n 0.00299761f $X=8.275 $Y=0.82 $X2=0 $Y2=0
cc_478 N_X_c_644_n N_VGND_c_878_n 0.00307254f $X=8.275 $Y=1.615 $X2=0 $Y2=0
cc_479 N_X_c_645_n N_VGND_c_878_n 0.0143045f $X=8.415 $Y=0.445 $X2=0 $Y2=0
cc_480 N_X_c_646_n N_VGND_c_880_n 0.0156284f $X=9.375 $Y=0.445 $X2=0 $Y2=0
cc_481 X N_VGND_c_880_n 0.00665978f $X=9.375 $Y=0.765 $X2=0 $Y2=0
cc_482 N_X_M1000_s N_VGND_c_883_n 0.00482172f $X=2.47 $Y=0.235 $X2=0 $Y2=0
cc_483 N_X_M1002_s N_VGND_c_883_n 0.00300326f $X=3.43 $Y=0.235 $X2=0 $Y2=0
cc_484 N_X_M1012_s N_VGND_c_883_n 0.00300326f $X=4.39 $Y=0.235 $X2=0 $Y2=0
cc_485 N_X_M1019_s N_VGND_c_883_n 0.00270667f $X=5.35 $Y=0.235 $X2=0 $Y2=0
cc_486 N_X_M1021_s N_VGND_c_883_n 0.00300326f $X=6.305 $Y=0.235 $X2=0 $Y2=0
cc_487 N_X_M1027_s N_VGND_c_883_n 0.00300326f $X=7.265 $Y=0.235 $X2=0 $Y2=0
cc_488 N_X_M1033_s N_VGND_c_883_n 0.00300326f $X=8.225 $Y=0.235 $X2=0 $Y2=0
cc_489 N_X_M1037_s N_VGND_c_883_n 0.00365899f $X=9.185 $Y=0.235 $X2=0 $Y2=0
cc_490 N_X_c_631_n N_VGND_c_883_n 0.00979224f $X=2.66 $Y=0.445 $X2=0 $Y2=0
cc_491 N_X_c_632_n N_VGND_c_883_n 0.0109571f $X=3.49 $Y=0.82 $X2=0 $Y2=0
cc_492 N_X_c_634_n N_VGND_c_883_n 0.00979224f $X=3.62 $Y=0.445 $X2=0 $Y2=0
cc_493 N_X_c_635_n N_VGND_c_883_n 0.0109571f $X=4.45 $Y=0.82 $X2=0 $Y2=0
cc_494 N_X_c_636_n N_VGND_c_883_n 0.00979224f $X=4.58 $Y=0.445 $X2=0 $Y2=0
cc_495 N_X_c_637_n N_VGND_c_883_n 0.00961597f $X=5.345 $Y=0.82 $X2=0 $Y2=0
cc_496 N_X_c_638_n N_VGND_c_883_n 0.0122303f $X=5.54 $Y=0.445 $X2=0 $Y2=0
cc_497 N_X_c_639_n N_VGND_c_883_n 0.010901f $X=6.355 $Y=0.82 $X2=0 $Y2=0
cc_498 N_X_c_640_n N_VGND_c_883_n 0.00979224f $X=6.495 $Y=0.445 $X2=0 $Y2=0
cc_499 N_X_c_641_n N_VGND_c_883_n 0.0111819f $X=7.315 $Y=0.82 $X2=0 $Y2=0
cc_500 N_X_c_642_n N_VGND_c_883_n 0.00979224f $X=7.455 $Y=0.445 $X2=0 $Y2=0
cc_501 N_X_c_643_n N_VGND_c_883_n 0.0111819f $X=8.275 $Y=0.82 $X2=0 $Y2=0
cc_502 N_X_c_644_n N_VGND_c_883_n 0.00510452f $X=8.275 $Y=1.615 $X2=0 $Y2=0
cc_503 N_X_c_645_n N_VGND_c_883_n 0.00979224f $X=8.415 $Y=0.445 $X2=0 $Y2=0
cc_504 N_X_c_646_n N_VGND_c_883_n 0.00981584f $X=9.375 $Y=0.445 $X2=0 $Y2=0
cc_505 X N_VGND_c_883_n 0.0132278f $X=9.375 $Y=0.765 $X2=0 $Y2=0
