* File: sky130_fd_sc_hdll__a21o_8.pxi.spice
* Created: Thu Aug 27 18:53:09 2020
* 
x_PM_SKY130_FD_SC_HDLL__A21O_8%A2 N_A2_c_112_n N_A2_M1011_g N_A2_c_113_n
+ N_A2_M1000_g N_A2_c_114_n N_A2_M1014_g N_A2_c_115_n N_A2_M1017_g N_A2_c_121_n
+ N_A2_c_122_n N_A2_c_163_p N_A2_c_116_n N_A2_c_117_n N_A2_c_118_n A2
+ PM_SKY130_FD_SC_HDLL__A21O_8%A2
x_PM_SKY130_FD_SC_HDLL__A21O_8%A1 N_A1_c_204_n N_A1_M1003_g N_A1_c_200_n
+ N_A1_M1008_g N_A1_c_201_n N_A1_M1004_g N_A1_c_205_n N_A1_M1024_g A1
+ N_A1_c_202_n N_A1_c_203_n PM_SKY130_FD_SC_HDLL__A21O_8%A1
x_PM_SKY130_FD_SC_HDLL__A21O_8%B1 N_B1_c_256_n N_B1_M1009_g N_B1_c_252_n
+ N_B1_M1016_g N_B1_c_253_n N_B1_M1023_g N_B1_c_257_n N_B1_M1012_g B1
+ N_B1_c_255_n PM_SKY130_FD_SC_HDLL__A21O_8%B1
x_PM_SKY130_FD_SC_HDLL__A21O_8%A_213_47# N_A_213_47#_M1008_d N_A_213_47#_M1016_d
+ N_A_213_47#_M1009_s N_A_213_47#_c_319_n N_A_213_47#_M1005_g
+ N_A_213_47#_c_306_n N_A_213_47#_M1001_g N_A_213_47#_c_307_n
+ N_A_213_47#_M1002_g N_A_213_47#_c_320_n N_A_213_47#_M1007_g
+ N_A_213_47#_c_321_n N_A_213_47#_M1013_g N_A_213_47#_c_308_n
+ N_A_213_47#_M1006_g N_A_213_47#_c_309_n N_A_213_47#_M1010_g
+ N_A_213_47#_c_322_n N_A_213_47#_M1015_g N_A_213_47#_c_323_n
+ N_A_213_47#_M1018_g N_A_213_47#_c_310_n N_A_213_47#_M1019_g
+ N_A_213_47#_c_311_n N_A_213_47#_M1020_g N_A_213_47#_c_324_n
+ N_A_213_47#_M1021_g N_A_213_47#_c_325_n N_A_213_47#_M1025_g
+ N_A_213_47#_c_312_n N_A_213_47#_M1022_g N_A_213_47#_c_313_n
+ N_A_213_47#_M1026_g N_A_213_47#_c_326_n N_A_213_47#_M1027_g
+ N_A_213_47#_c_329_n N_A_213_47#_c_331_n N_A_213_47#_c_314_n
+ N_A_213_47#_c_336_n N_A_213_47#_c_315_n N_A_213_47#_c_358_n
+ N_A_213_47#_c_316_n N_A_213_47#_c_317_n N_A_213_47#_c_414_p
+ N_A_213_47#_c_365_n N_A_213_47#_c_366_n N_A_213_47#_c_318_n
+ PM_SKY130_FD_SC_HDLL__A21O_8%A_213_47#
x_PM_SKY130_FD_SC_HDLL__A21O_8%A_27_297# N_A_27_297#_M1011_s N_A_27_297#_M1003_d
+ N_A_27_297#_M1017_s N_A_27_297#_M1012_d N_A_27_297#_c_521_n
+ N_A_27_297#_c_522_n N_A_27_297#_c_532_n N_A_27_297#_c_536_n
+ N_A_27_297#_c_539_n N_A_27_297#_c_523_n N_A_27_297#_c_524_n
+ N_A_27_297#_c_541_n N_A_27_297#_c_525_n N_A_27_297#_c_526_n
+ N_A_27_297#_c_544_n N_A_27_297#_c_547_n PM_SKY130_FD_SC_HDLL__A21O_8%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A21O_8%VPWR N_VPWR_M1011_d N_VPWR_M1024_s N_VPWR_M1005_s
+ N_VPWR_M1007_s N_VPWR_M1015_s N_VPWR_M1021_s N_VPWR_M1027_s N_VPWR_c_593_n
+ N_VPWR_c_594_n N_VPWR_c_595_n N_VPWR_c_596_n N_VPWR_c_597_n N_VPWR_c_598_n
+ N_VPWR_c_599_n N_VPWR_c_600_n N_VPWR_c_601_n N_VPWR_c_602_n N_VPWR_c_603_n
+ N_VPWR_c_604_n N_VPWR_c_605_n N_VPWR_c_606_n N_VPWR_c_607_n N_VPWR_c_608_n
+ N_VPWR_c_609_n N_VPWR_c_610_n VPWR N_VPWR_c_611_n N_VPWR_c_612_n
+ N_VPWR_c_592_n N_VPWR_c_614_n N_VPWR_c_615_n PM_SKY130_FD_SC_HDLL__A21O_8%VPWR
x_PM_SKY130_FD_SC_HDLL__A21O_8%X N_X_M1001_d N_X_M1006_d N_X_M1019_d N_X_M1022_d
+ N_X_M1005_d N_X_M1013_d N_X_M1018_d N_X_M1025_d N_X_c_724_n N_X_c_797_n
+ N_X_c_716_n N_X_c_717_n N_X_c_734_n N_X_c_738_n N_X_c_742_n N_X_c_801_n
+ N_X_c_718_n N_X_c_750_n N_X_c_754_n N_X_c_805_n N_X_c_719_n N_X_c_761_n
+ N_X_c_764_n N_X_c_720_n N_X_c_810_n N_X_c_770_n N_X_c_721_n N_X_c_776_n
+ N_X_c_722_n N_X_c_782_n X PM_SKY130_FD_SC_HDLL__A21O_8%X
x_PM_SKY130_FD_SC_HDLL__A21O_8%VGND N_VGND_M1000_s N_VGND_M1014_s N_VGND_M1023_s
+ N_VGND_M1002_s N_VGND_M1010_s N_VGND_M1020_s N_VGND_M1026_s N_VGND_c_843_n
+ N_VGND_c_844_n N_VGND_c_845_n N_VGND_c_846_n N_VGND_c_847_n N_VGND_c_848_n
+ N_VGND_c_849_n N_VGND_c_850_n N_VGND_c_851_n N_VGND_c_852_n N_VGND_c_853_n
+ N_VGND_c_854_n N_VGND_c_855_n N_VGND_c_856_n N_VGND_c_857_n VGND
+ N_VGND_c_858_n N_VGND_c_859_n N_VGND_c_860_n N_VGND_c_861_n N_VGND_c_862_n
+ N_VGND_c_863_n PM_SKY130_FD_SC_HDLL__A21O_8%VGND
cc_1 VNB N_A2_c_112_n 0.0293869f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_A2_c_113_n 0.0211848f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.995
cc_3 VNB N_A2_c_114_n 0.017665f $X=-0.19 $Y=-0.24 $X2=1.82 $Y2=0.995
cc_4 VNB N_A2_c_115_n 0.0197856f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_5 VNB N_A2_c_116_n 2.55318e-19 $X=-0.19 $Y=-0.24 $X2=1.79 $Y2=1.46
cc_6 VNB N_A2_c_117_n 0.0199748f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.172
cc_7 VNB N_A2_c_118_n 0.00458328f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_8 VNB N_A1_c_200_n 0.0161331f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.995
cc_9 VNB N_A1_c_201_n 0.0161021f $X=-0.19 $Y=-0.24 $X2=1.82 $Y2=0.995
cc_10 VNB N_A1_c_202_n 0.00291039f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.172
cc_11 VNB N_A1_c_203_n 0.035465f $X=-0.19 $Y=-0.24 $X2=1.79 $Y2=1.172
cc_12 VNB N_B1_c_252_n 0.0170767f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.995
cc_13 VNB N_B1_c_253_n 0.0201851f $X=-0.19 $Y=-0.24 $X2=1.82 $Y2=0.995
cc_14 VNB B1 0.00256212f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.29
cc_15 VNB N_B1_c_255_n 0.0540894f $X=-0.19 $Y=-0.24 $X2=1.79 $Y2=1.46
cc_16 VNB N_A_213_47#_c_306_n 0.0191654f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.29
cc_17 VNB N_A_213_47#_c_307_n 0.0169283f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.545
cc_18 VNB N_A_213_47#_c_308_n 0.0169331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_213_47#_c_309_n 0.0169331f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_20 VNB N_A_213_47#_c_310_n 0.0169331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_213_47#_c_311_n 0.0169059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_213_47#_c_312_n 0.0159577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_213_47#_c_313_n 0.0214454f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_213_47#_c_314_n 0.00115748f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_213_47#_c_315_n 0.00103672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_213_47#_c_316_n 0.00339889f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_213_47#_c_317_n 0.00399351f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_213_47#_c_318_n 0.169466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_592_n 0.326667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB X 0.00235317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_843_n 0.0138449f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.172
cc_32 VNB N_VGND_c_844_n 0.0297009f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_33 VNB N_VGND_c_845_n 0.00501005f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_34 VNB N_VGND_c_846_n 0.00413904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_847_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_848_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_849_n 0.0329153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_850_n 0.0172699f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_851_n 0.00515784f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_852_n 0.0165909f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_853_n 0.00515784f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_854_n 0.0165909f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_855_n 0.00515784f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_856_n 0.0172686f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_857_n 0.00480536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_858_n 0.0384028f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_859_n 0.0131219f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_860_n 0.385252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_861_n 0.00631346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_862_n 0.0159607f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_863_n 0.0229593f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VPB N_A2_c_112_n 0.0332672f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_53 VPB N_A2_c_115_n 0.0243889f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_54 VPB N_A2_c_121_n 0.00148131f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.46
cc_55 VPB N_A2_c_122_n 0.0102624f $X=-0.19 $Y=1.305 $X2=1.705 $Y2=1.545
cc_56 VPB N_A2_c_116_n 0.00148131f $X=-0.19 $Y=1.305 $X2=1.79 $Y2=1.46
cc_57 VPB N_A1_c_204_n 0.016105f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_58 VPB N_A1_c_205_n 0.016105f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_59 VPB N_A1_c_203_n 0.0195118f $X=-0.19 $Y=1.305 $X2=1.79 $Y2=1.172
cc_60 VPB N_B1_c_256_n 0.0161061f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_61 VPB N_B1_c_257_n 0.0195953f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_62 VPB B1 0.00260515f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.29
cc_63 VPB N_B1_c_255_n 0.0295495f $X=-0.19 $Y=1.305 $X2=1.79 $Y2=1.46
cc_64 VPB N_A_213_47#_c_319_n 0.0197254f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_65 VPB N_A_213_47#_c_320_n 0.0157197f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.172
cc_66 VPB N_A_213_47#_c_321_n 0.0157197f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.172
cc_67 VPB N_A_213_47#_c_322_n 0.0157197f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_68 VPB N_A_213_47#_c_323_n 0.0157197f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_213_47#_c_324_n 0.015696f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_213_47#_c_325_n 0.0153999f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_213_47#_c_326_n 0.0199368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_213_47#_c_315_n 9.30672e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_213_47#_c_318_n 0.102536f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_297#_c_521_n 0.0153465f $X=-0.19 $Y=1.305 $X2=1.705 $Y2=1.545
cc_75 VPB N_A_27_297#_c_522_n 0.0194072f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.172
cc_76 VPB N_A_27_297#_c_523_n 0.00407295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_297#_c_524_n 0.0019327f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.172
cc_78 VPB N_A_27_297#_c_525_n 0.00645964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_27_297#_c_526_n 0.00717518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_593_n 0.00466368f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_81 VPB N_VPWR_c_594_n 0.0167297f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_82 VPB N_VPWR_c_595_n 0.0046582f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_83 VPB N_VPWR_c_596_n 0.00462153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_597_n 3.40287e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_598_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_599_n 3.38822e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_600_n 0.0510468f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_601_n 0.0404498f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_602_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_603_n 0.0167344f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_604_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_605_n 0.0147329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_606_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_607_n 0.0147329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_608_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_609_n 0.0164162f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_610_n 0.00593688f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_611_n 0.0172595f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_612_n 0.0115308f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_592_n 0.0623934f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_614_n 0.00516022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_615_n 0.00515985f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_X_c_716_n 0.00180924f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.172
cc_104 VPB N_X_c_717_n 0.00215492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_X_c_718_n 0.00180924f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_X_c_719_n 0.00224041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_X_c_720_n 0.00230295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_X_c_721_n 0.00162501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_X_c_722_n 0.00162501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB X 0.00275881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 N_A2_c_112_n N_A1_c_204_n 0.0364735f $X=0.495 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_112 N_A2_c_121_n N_A1_c_204_n 0.00101315f $X=0.61 $Y=1.46 $X2=-0.19 $Y2=-0.24
cc_113 N_A2_c_122_n N_A1_c_204_n 0.0118662f $X=1.705 $Y=1.545 $X2=-0.19
+ $Y2=-0.24
cc_114 N_A2_c_113_n N_A1_c_200_n 0.0418602f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A2_c_114_n N_A1_c_201_n 0.0440841f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A2_c_115_n N_A1_c_205_n 0.0364735f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A2_c_122_n N_A1_c_205_n 0.0118662f $X=1.705 $Y=1.545 $X2=0 $Y2=0
cc_118 N_A2_c_116_n N_A1_c_205_n 0.00101315f $X=1.79 $Y=1.46 $X2=0 $Y2=0
cc_119 N_A2_c_112_n N_A1_c_202_n 2.66334e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A2_c_115_n N_A1_c_202_n 2.67076e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A2_c_122_n N_A1_c_202_n 0.0477309f $X=1.705 $Y=1.545 $X2=0 $Y2=0
cc_122 N_A2_c_117_n N_A1_c_202_n 0.0205474f $X=0.525 $Y=1.172 $X2=0 $Y2=0
cc_123 N_A2_c_118_n N_A1_c_202_n 0.0196709f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A2_c_112_n N_A1_c_203_n 0.0260406f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A2_c_115_n N_A1_c_203_n 0.0259586f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A2_c_121_n N_A1_c_203_n 0.0024835f $X=0.61 $Y=1.46 $X2=0 $Y2=0
cc_127 N_A2_c_122_n N_A1_c_203_n 0.0081936f $X=1.705 $Y=1.545 $X2=0 $Y2=0
cc_128 N_A2_c_116_n N_A1_c_203_n 0.00250084f $X=1.79 $Y=1.46 $X2=0 $Y2=0
cc_129 N_A2_c_117_n N_A1_c_203_n 8.47697e-19 $X=0.525 $Y=1.172 $X2=0 $Y2=0
cc_130 N_A2_c_118_n N_A1_c_203_n 7.65384e-19 $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A2_c_115_n N_B1_c_256_n 0.00914847f $X=1.905 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_132 N_A2_c_114_n N_B1_c_252_n 0.0223862f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A2_c_115_n N_B1_c_255_n 0.02115f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A2_c_116_n N_B1_c_255_n 3.96194e-19 $X=1.79 $Y=1.46 $X2=0 $Y2=0
cc_135 N_A2_c_118_n N_B1_c_255_n 0.00207728f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A2_c_113_n N_A_213_47#_c_329_n 0.00116223f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A2_c_114_n N_A_213_47#_c_329_n 0.00153389f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A2_c_114_n N_A_213_47#_c_331_n 0.0142266f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A2_c_115_n N_A_213_47#_c_331_n 0.00318656f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A2_c_122_n N_A_213_47#_c_331_n 0.00493675f $X=1.705 $Y=1.545 $X2=0
+ $Y2=0
cc_141 N_A2_c_118_n N_A_213_47#_c_331_n 0.0211231f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A2_c_113_n N_A_213_47#_c_314_n 6.08286e-19 $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A2_c_114_n N_A_213_47#_c_336_n 8.26073e-19 $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A2_c_114_n N_A_213_47#_c_315_n 4.98365e-19 $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A2_c_115_n N_A_213_47#_c_315_n 0.00110089f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A2_c_116_n N_A_213_47#_c_315_n 0.00434447f $X=1.79 $Y=1.46 $X2=0 $Y2=0
cc_147 N_A2_c_118_n N_A_213_47#_c_315_n 0.00960727f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A2_c_122_n N_A_27_297#_M1003_d 0.00187091f $X=1.705 $Y=1.545 $X2=0
+ $Y2=0
cc_149 N_A2_c_112_n N_A_27_297#_c_521_n 0.00128062f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A2_c_163_p N_A_27_297#_c_521_n 0.00812827f $X=0.695 $Y=1.545 $X2=0
+ $Y2=0
cc_151 N_A2_c_117_n N_A_27_297#_c_521_n 0.022168f $X=0.525 $Y=1.172 $X2=0 $Y2=0
cc_152 N_A2_c_112_n N_A_27_297#_c_522_n 0.00681523f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A2_c_112_n N_A_27_297#_c_532_n 0.0121086f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A2_c_122_n N_A_27_297#_c_532_n 0.0197085f $X=1.705 $Y=1.545 $X2=0 $Y2=0
cc_155 N_A2_c_163_p N_A_27_297#_c_532_n 0.00871932f $X=0.695 $Y=1.545 $X2=0
+ $Y2=0
cc_156 N_A2_c_117_n N_A_27_297#_c_532_n 0.00280628f $X=0.525 $Y=1.172 $X2=0
+ $Y2=0
cc_157 N_A2_c_115_n N_A_27_297#_c_536_n 0.0121086f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A2_c_122_n N_A_27_297#_c_536_n 0.0280721f $X=1.705 $Y=1.545 $X2=0 $Y2=0
cc_159 N_A2_c_118_n N_A_27_297#_c_536_n 0.00285382f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A2_c_115_n N_A_27_297#_c_539_n 0.00486243f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A2_c_122_n N_A_27_297#_c_523_n 0.00811046f $X=1.705 $Y=1.545 $X2=0
+ $Y2=0
cc_162 N_A2_c_115_n N_A_27_297#_c_541_n 0.00195885f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A2_c_112_n N_A_27_297#_c_526_n 7.83256e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A2_c_117_n N_A_27_297#_c_526_n 0.00134292f $X=0.525 $Y=1.172 $X2=0
+ $Y2=0
cc_165 N_A2_c_112_n N_A_27_297#_c_544_n 5.15302e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A2_c_115_n N_A_27_297#_c_544_n 5.15302e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A2_c_122_n N_A_27_297#_c_544_n 0.0172506f $X=1.705 $Y=1.545 $X2=0 $Y2=0
cc_168 N_A2_c_115_n N_A_27_297#_c_547_n 8.09873e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A2_c_118_n N_A_27_297#_c_547_n 0.00146178f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A2_c_122_n N_VPWR_M1011_d 0.00130005f $X=1.705 $Y=1.545 $X2=-0.19
+ $Y2=-0.24
cc_171 N_A2_c_163_p N_VPWR_M1011_d 5.84953e-19 $X=0.695 $Y=1.545 $X2=-0.19
+ $Y2=-0.24
cc_172 N_A2_c_122_n N_VPWR_M1024_s 0.00186483f $X=1.705 $Y=1.545 $X2=0 $Y2=0
cc_173 N_A2_c_112_n N_VPWR_c_593_n 0.00309049f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A2_c_115_n N_VPWR_c_595_n 0.00309049f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A2_c_115_n N_VPWR_c_601_n 0.00518316f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A2_c_112_n N_VPWR_c_611_n 0.00519834f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A2_c_112_n N_VPWR_c_592_n 0.00767899f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A2_c_115_n N_VPWR_c_592_n 0.00680185f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A2_c_112_n N_VGND_c_844_n 0.00474596f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A2_c_113_n N_VGND_c_844_n 0.0176088f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A2_c_117_n N_VGND_c_844_n 0.0243306f $X=0.525 $Y=1.172 $X2=0 $Y2=0
cc_182 N_A2_c_114_n N_VGND_c_845_n 0.00475459f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A2_c_113_n N_VGND_c_858_n 0.0046653f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A2_c_114_n N_VGND_c_858_n 0.00430895f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A2_c_113_n N_VGND_c_860_n 0.00796999f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A2_c_114_n N_VGND_c_860_n 0.00623871f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A1_c_200_n N_A_213_47#_c_329_n 0.00712196f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A1_c_201_n N_A_213_47#_c_329_n 0.00761603f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A1_c_201_n N_A_213_47#_c_331_n 0.00910922f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A1_c_202_n N_A_213_47#_c_331_n 0.0102215f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A1_c_200_n N_A_213_47#_c_314_n 0.0040234f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A1_c_201_n N_A_213_47#_c_314_n 9.7745e-19 $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A1_c_202_n N_A_213_47#_c_314_n 0.0211043f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A1_c_203_n N_A_213_47#_c_314_n 0.00224326f $X=1.41 $Y=1.202 $X2=0 $Y2=0
cc_195 N_A1_c_204_n N_A_27_297#_c_522_n 5.15302e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A1_c_204_n N_A_27_297#_c_532_n 0.0108454f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A1_c_205_n N_A_27_297#_c_536_n 0.0108454f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A1_c_205_n N_A_27_297#_c_539_n 4.72751e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A1_c_204_n N_A_27_297#_c_544_n 0.00769006f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_200 N_A1_c_205_n N_A_27_297#_c_544_n 0.00769006f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A1_c_204_n N_VPWR_c_593_n 0.00173895f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A1_c_204_n N_VPWR_c_594_n 0.00519834f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A1_c_205_n N_VPWR_c_594_n 0.00519834f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A1_c_205_n N_VPWR_c_595_n 0.00173895f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A1_c_204_n N_VPWR_c_592_n 0.00676756f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A1_c_205_n N_VPWR_c_592_n 0.00676756f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A1_c_200_n N_VGND_c_844_n 0.00302624f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A1_c_200_n N_VGND_c_858_n 0.00542163f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A1_c_201_n N_VGND_c_858_n 0.00418572f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A1_c_200_n N_VGND_c_860_n 0.00970348f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A1_c_201_n N_VGND_c_860_n 0.00578774f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_212 B1 N_A_213_47#_c_319_n 0.00228471f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_213 N_B1_c_252_n N_A_213_47#_c_331_n 0.0139202f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_214 N_B1_c_252_n N_A_213_47#_c_336_n 0.00640026f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_215 N_B1_c_256_n N_A_213_47#_c_315_n 0.00506273f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_216 N_B1_c_252_n N_A_213_47#_c_315_n 0.00314306f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_217 N_B1_c_253_n N_A_213_47#_c_315_n 0.00279934f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B1_c_257_n N_A_213_47#_c_315_n 0.0046097f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_219 B1 N_A_213_47#_c_315_n 0.0421322f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_220 N_B1_c_255_n N_A_213_47#_c_315_n 0.0299017f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_221 N_B1_c_253_n N_A_213_47#_c_358_n 0.0172949f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_222 B1 N_A_213_47#_c_358_n 0.0235839f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_223 N_B1_c_255_n N_A_213_47#_c_358_n 0.00728832f $X=2.845 $Y=1.202 $X2=0
+ $Y2=0
cc_224 N_B1_c_253_n N_A_213_47#_c_316_n 0.00222925f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_225 N_B1_c_255_n N_A_213_47#_c_316_n 7.80627e-19 $X=2.845 $Y=1.202 $X2=0
+ $Y2=0
cc_226 B1 N_A_213_47#_c_317_n 0.0103841f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_227 N_B1_c_255_n N_A_213_47#_c_317_n 0.00164768f $X=2.845 $Y=1.202 $X2=0
+ $Y2=0
cc_228 N_B1_c_252_n N_A_213_47#_c_365_n 5.73461e-19 $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_229 N_B1_c_256_n N_A_213_47#_c_366_n 0.0037767f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_230 N_B1_c_255_n N_A_213_47#_c_366_n 9.13766e-19 $X=2.845 $Y=1.202 $X2=0
+ $Y2=0
cc_231 B1 N_A_213_47#_c_318_n 0.00275109f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_232 N_B1_c_255_n N_A_213_47#_c_318_n 0.00576975f $X=2.845 $Y=1.202 $X2=0
+ $Y2=0
cc_233 B1 N_A_27_297#_M1012_d 0.00431235f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_234 N_B1_c_256_n N_A_27_297#_c_523_n 2.03034e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_235 N_B1_c_256_n N_A_27_297#_c_524_n 0.0137768f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_236 N_B1_c_257_n N_A_27_297#_c_524_n 0.0134429f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_237 N_B1_c_256_n N_A_27_297#_c_525_n 4.38946e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_238 N_B1_c_257_n N_A_27_297#_c_525_n 0.00878804f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_239 B1 N_A_27_297#_c_525_n 0.0194936f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_240 N_B1_c_255_n N_A_27_297#_c_525_n 9.68667e-19 $X=2.845 $Y=1.202 $X2=0
+ $Y2=0
cc_241 N_B1_c_257_n N_VPWR_c_596_n 0.00677716f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_242 B1 N_VPWR_c_596_n 0.00633255f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_243 N_B1_c_256_n N_VPWR_c_601_n 0.00429453f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_244 N_B1_c_257_n N_VPWR_c_601_n 0.00429425f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_245 N_B1_c_256_n N_VPWR_c_592_n 0.00609021f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_246 N_B1_c_257_n N_VPWR_c_592_n 0.00734732f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_247 N_B1_c_252_n N_VGND_c_845_n 0.00338986f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_248 N_B1_c_252_n N_VGND_c_860_n 0.00604629f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_249 N_B1_c_253_n N_VGND_c_860_n 0.00701283f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_250 N_B1_c_252_n N_VGND_c_862_n 0.00417768f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_251 N_B1_c_253_n N_VGND_c_862_n 0.00430895f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_252 N_B1_c_253_n N_VGND_c_863_n 0.00353715f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A_213_47#_c_331_n N_A_27_297#_c_523_n 0.00791064f $X=2.445 $Y=0.78
+ $X2=0 $Y2=0
cc_254 N_A_213_47#_c_315_n N_A_27_297#_c_523_n 0.0131458f $X=2.61 $Y=1.62 $X2=0
+ $Y2=0
cc_255 N_A_213_47#_M1009_s N_A_27_297#_c_524_n 0.00344383f $X=2.465 $Y=1.485
+ $X2=0 $Y2=0
cc_256 N_A_213_47#_c_366_n N_A_27_297#_c_524_n 0.0147165f $X=2.61 $Y=1.96 $X2=0
+ $Y2=0
cc_257 N_A_213_47#_c_315_n N_A_27_297#_c_525_n 2.79839e-19 $X=2.61 $Y=1.62 $X2=0
+ $Y2=0
cc_258 N_A_213_47#_c_319_n N_VPWR_c_596_n 0.00349953f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_259 N_A_213_47#_c_358_n N_VPWR_c_596_n 0.00248426f $X=3.565 $Y=0.78 $X2=0
+ $Y2=0
cc_260 N_A_213_47#_c_317_n N_VPWR_c_596_n 0.0110476f $X=3.735 $Y=1.155 $X2=0
+ $Y2=0
cc_261 N_A_213_47#_c_319_n N_VPWR_c_597_n 6.17091e-19 $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_262 N_A_213_47#_c_320_n N_VPWR_c_597_n 0.0128989f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_263 N_A_213_47#_c_321_n N_VPWR_c_597_n 0.0128391f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_264 N_A_213_47#_c_322_n N_VPWR_c_597_n 6.06824e-19 $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_265 N_A_213_47#_c_321_n N_VPWR_c_598_n 6.06824e-19 $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_266 N_A_213_47#_c_322_n N_VPWR_c_598_n 0.0128391f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_267 N_A_213_47#_c_323_n N_VPWR_c_598_n 0.0128391f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_268 N_A_213_47#_c_324_n N_VPWR_c_598_n 6.06824e-19 $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_269 N_A_213_47#_c_323_n N_VPWR_c_599_n 6.06824e-19 $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_270 N_A_213_47#_c_324_n N_VPWR_c_599_n 0.0128391f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_271 N_A_213_47#_c_325_n N_VPWR_c_599_n 0.0128792f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_272 N_A_213_47#_c_326_n N_VPWR_c_599_n 6.1369e-19 $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_273 N_A_213_47#_c_326_n N_VPWR_c_600_n 0.00457324f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_274 N_A_213_47#_c_318_n N_VPWR_c_600_n 0.00217332f $X=7.1 $Y=1.202 $X2=0
+ $Y2=0
cc_275 N_A_213_47#_c_319_n N_VPWR_c_603_n 0.00702461f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_276 N_A_213_47#_c_320_n N_VPWR_c_603_n 0.00622633f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_277 N_A_213_47#_c_321_n N_VPWR_c_605_n 0.00622633f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_278 N_A_213_47#_c_322_n N_VPWR_c_605_n 0.00622633f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_279 N_A_213_47#_c_323_n N_VPWR_c_607_n 0.00622633f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_280 N_A_213_47#_c_324_n N_VPWR_c_607_n 0.00622633f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_281 N_A_213_47#_c_325_n N_VPWR_c_609_n 0.00622633f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_282 N_A_213_47#_c_326_n N_VPWR_c_609_n 0.00700684f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_283 N_A_213_47#_M1009_s N_VPWR_c_592_n 0.00232895f $X=2.465 $Y=1.485 $X2=0
+ $Y2=0
cc_284 N_A_213_47#_c_319_n N_VPWR_c_592_n 0.0136664f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_285 N_A_213_47#_c_320_n N_VPWR_c_592_n 0.0104011f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_286 N_A_213_47#_c_321_n N_VPWR_c_592_n 0.0104011f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_287 N_A_213_47#_c_322_n N_VPWR_c_592_n 0.0104011f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_288 N_A_213_47#_c_323_n N_VPWR_c_592_n 0.0104011f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_289 N_A_213_47#_c_324_n N_VPWR_c_592_n 0.0104011f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_290 N_A_213_47#_c_325_n N_VPWR_c_592_n 0.0104011f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_291 N_A_213_47#_c_326_n N_VPWR_c_592_n 0.013396f $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_292 N_A_213_47#_c_306_n N_X_c_724_n 0.0106602f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_293 N_A_213_47#_c_307_n N_X_c_724_n 0.00639957f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_294 N_A_213_47#_c_308_n N_X_c_724_n 5.17822e-19 $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_295 N_A_213_47#_c_320_n N_X_c_716_n 0.0150944f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_296 N_A_213_47#_c_321_n N_X_c_716_n 0.0151703f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_297 N_A_213_47#_c_414_p N_X_c_716_n 0.0477325f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_298 N_A_213_47#_c_318_n N_X_c_716_n 0.00798413f $X=7.1 $Y=1.202 $X2=0 $Y2=0
cc_299 N_A_213_47#_c_319_n N_X_c_717_n 0.0013234f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_300 N_A_213_47#_c_414_p N_X_c_717_n 0.0222834f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_301 N_A_213_47#_c_318_n N_X_c_717_n 0.00743165f $X=7.1 $Y=1.202 $X2=0 $Y2=0
cc_302 N_A_213_47#_c_307_n N_X_c_734_n 0.00893375f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_303 N_A_213_47#_c_308_n N_X_c_734_n 0.00893375f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_304 N_A_213_47#_c_414_p N_X_c_734_n 0.0391608f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_305 N_A_213_47#_c_318_n N_X_c_734_n 0.00446519f $X=7.1 $Y=1.202 $X2=0 $Y2=0
cc_306 N_A_213_47#_c_306_n N_X_c_738_n 0.00227599f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_307 N_A_213_47#_c_307_n N_X_c_738_n 8.68219e-19 $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_308 N_A_213_47#_c_414_p N_X_c_738_n 0.0211425f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_309 N_A_213_47#_c_318_n N_X_c_738_n 0.00218937f $X=7.1 $Y=1.202 $X2=0 $Y2=0
cc_310 N_A_213_47#_c_307_n N_X_c_742_n 5.17822e-19 $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_311 N_A_213_47#_c_308_n N_X_c_742_n 0.00639957f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_312 N_A_213_47#_c_309_n N_X_c_742_n 0.00639957f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_313 N_A_213_47#_c_310_n N_X_c_742_n 5.17822e-19 $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_314 N_A_213_47#_c_322_n N_X_c_718_n 0.0151703f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_315 N_A_213_47#_c_323_n N_X_c_718_n 0.0151703f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_316 N_A_213_47#_c_414_p N_X_c_718_n 0.0477325f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_317 N_A_213_47#_c_318_n N_X_c_718_n 0.00798413f $X=7.1 $Y=1.202 $X2=0 $Y2=0
cc_318 N_A_213_47#_c_309_n N_X_c_750_n 0.00893375f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_319 N_A_213_47#_c_310_n N_X_c_750_n 0.00893375f $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_320 N_A_213_47#_c_414_p N_X_c_750_n 0.0391608f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_321 N_A_213_47#_c_318_n N_X_c_750_n 0.00446519f $X=7.1 $Y=1.202 $X2=0 $Y2=0
cc_322 N_A_213_47#_c_309_n N_X_c_754_n 5.17822e-19 $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_323 N_A_213_47#_c_310_n N_X_c_754_n 0.00639957f $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_324 N_A_213_47#_c_311_n N_X_c_754_n 0.00639957f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_325 N_A_213_47#_c_312_n N_X_c_754_n 5.17822e-19 $X=6.68 $Y=0.995 $X2=0 $Y2=0
cc_326 N_A_213_47#_c_324_n N_X_c_719_n 0.0169197f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_327 N_A_213_47#_c_414_p N_X_c_719_n 0.00348096f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_328 N_A_213_47#_c_318_n N_X_c_719_n 0.00836679f $X=7.1 $Y=1.202 $X2=0 $Y2=0
cc_329 N_A_213_47#_c_311_n N_X_c_761_n 0.0101833f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_330 N_A_213_47#_c_414_p N_X_c_761_n 0.00135861f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_331 N_A_213_47#_c_318_n N_X_c_761_n 0.00531719f $X=7.1 $Y=1.202 $X2=0 $Y2=0
cc_332 N_A_213_47#_c_311_n N_X_c_764_n 5.17822e-19 $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_333 N_A_213_47#_c_312_n N_X_c_764_n 0.00639957f $X=6.68 $Y=0.995 $X2=0 $Y2=0
cc_334 N_A_213_47#_c_313_n N_X_c_764_n 0.00506666f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_335 N_A_213_47#_c_325_n N_X_c_720_n 0.013198f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_336 N_A_213_47#_c_326_n N_X_c_720_n 3.7313e-19 $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_337 N_A_213_47#_c_318_n N_X_c_720_n 0.00763541f $X=7.1 $Y=1.202 $X2=0 $Y2=0
cc_338 N_A_213_47#_c_308_n N_X_c_770_n 8.68219e-19 $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_339 N_A_213_47#_c_309_n N_X_c_770_n 8.68219e-19 $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_340 N_A_213_47#_c_414_p N_X_c_770_n 0.0211425f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_341 N_A_213_47#_c_318_n N_X_c_770_n 0.00218937f $X=7.1 $Y=1.202 $X2=0 $Y2=0
cc_342 N_A_213_47#_c_414_p N_X_c_721_n 0.0222834f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_343 N_A_213_47#_c_318_n N_X_c_721_n 0.00743165f $X=7.1 $Y=1.202 $X2=0 $Y2=0
cc_344 N_A_213_47#_c_310_n N_X_c_776_n 8.68219e-19 $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_345 N_A_213_47#_c_311_n N_X_c_776_n 8.68219e-19 $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_346 N_A_213_47#_c_414_p N_X_c_776_n 0.0211425f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_347 N_A_213_47#_c_318_n N_X_c_776_n 0.00218937f $X=7.1 $Y=1.202 $X2=0 $Y2=0
cc_348 N_A_213_47#_c_414_p N_X_c_722_n 0.0222834f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_349 N_A_213_47#_c_318_n N_X_c_722_n 0.00743165f $X=7.1 $Y=1.202 $X2=0 $Y2=0
cc_350 N_A_213_47#_c_312_n N_X_c_782_n 0.00785862f $X=6.68 $Y=0.995 $X2=0 $Y2=0
cc_351 N_A_213_47#_c_313_n N_X_c_782_n 0.00328757f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_352 N_A_213_47#_c_318_n N_X_c_782_n 0.0027324f $X=7.1 $Y=1.202 $X2=0 $Y2=0
cc_353 N_A_213_47#_c_311_n X 0.00252921f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_354 N_A_213_47#_c_324_n X 6.96836e-19 $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_355 N_A_213_47#_c_325_n X 0.00143298f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_356 N_A_213_47#_c_312_n X 0.00310338f $X=6.68 $Y=0.995 $X2=0 $Y2=0
cc_357 N_A_213_47#_c_313_n X 0.00200553f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_358 N_A_213_47#_c_326_n X 7.22019e-19 $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_359 N_A_213_47#_c_414_p X 0.00913163f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_360 N_A_213_47#_c_318_n X 0.0384257f $X=7.1 $Y=1.202 $X2=0 $Y2=0
cc_361 N_A_213_47#_c_331_n N_VGND_M1014_s 0.00924222f $X=2.445 $Y=0.78 $X2=0
+ $Y2=0
cc_362 N_A_213_47#_c_358_n N_VGND_M1023_s 0.0301698f $X=3.565 $Y=0.78 $X2=0
+ $Y2=0
cc_363 N_A_213_47#_c_329_n N_VGND_c_844_n 0.0124356f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_364 N_A_213_47#_c_314_n N_VGND_c_844_n 0.00693247f $X=1.365 $Y=0.78 $X2=0
+ $Y2=0
cc_365 N_A_213_47#_c_331_n N_VGND_c_845_n 0.0247398f $X=2.445 $Y=0.78 $X2=0
+ $Y2=0
cc_366 N_A_213_47#_c_307_n N_VGND_c_846_n 0.00166738f $X=4.28 $Y=0.995 $X2=0
+ $Y2=0
cc_367 N_A_213_47#_c_308_n N_VGND_c_846_n 0.00166854f $X=4.8 $Y=0.995 $X2=0
+ $Y2=0
cc_368 N_A_213_47#_c_309_n N_VGND_c_847_n 0.00166854f $X=5.22 $Y=0.995 $X2=0
+ $Y2=0
cc_369 N_A_213_47#_c_310_n N_VGND_c_847_n 0.00166854f $X=5.74 $Y=0.995 $X2=0
+ $Y2=0
cc_370 N_A_213_47#_c_311_n N_VGND_c_848_n 0.00166854f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_371 N_A_213_47#_c_312_n N_VGND_c_848_n 0.00166854f $X=6.68 $Y=0.995 $X2=0
+ $Y2=0
cc_372 N_A_213_47#_c_313_n N_VGND_c_849_n 0.00372903f $X=7.1 $Y=0.995 $X2=0
+ $Y2=0
cc_373 N_A_213_47#_c_318_n N_VGND_c_849_n 0.00171941f $X=7.1 $Y=1.202 $X2=0
+ $Y2=0
cc_374 N_A_213_47#_c_306_n N_VGND_c_850_n 0.00541359f $X=3.86 $Y=0.995 $X2=0
+ $Y2=0
cc_375 N_A_213_47#_c_307_n N_VGND_c_850_n 0.00420025f $X=4.28 $Y=0.995 $X2=0
+ $Y2=0
cc_376 N_A_213_47#_c_308_n N_VGND_c_852_n 0.00420025f $X=4.8 $Y=0.995 $X2=0
+ $Y2=0
cc_377 N_A_213_47#_c_309_n N_VGND_c_852_n 0.00420025f $X=5.22 $Y=0.995 $X2=0
+ $Y2=0
cc_378 N_A_213_47#_c_310_n N_VGND_c_854_n 0.00420025f $X=5.74 $Y=0.995 $X2=0
+ $Y2=0
cc_379 N_A_213_47#_c_311_n N_VGND_c_854_n 0.00420025f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_380 N_A_213_47#_c_312_n N_VGND_c_856_n 0.00419913f $X=6.68 $Y=0.995 $X2=0
+ $Y2=0
cc_381 N_A_213_47#_c_313_n N_VGND_c_856_n 0.00541359f $X=7.1 $Y=0.995 $X2=0
+ $Y2=0
cc_382 N_A_213_47#_c_329_n N_VGND_c_858_n 0.0166744f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_383 N_A_213_47#_c_331_n N_VGND_c_858_n 0.00789631f $X=2.445 $Y=0.78 $X2=0
+ $Y2=0
cc_384 N_A_213_47#_M1008_d N_VGND_c_860_n 0.00216035f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_385 N_A_213_47#_M1016_d N_VGND_c_860_n 0.00215201f $X=2.475 $Y=0.235 $X2=0
+ $Y2=0
cc_386 N_A_213_47#_c_306_n N_VGND_c_860_n 0.0109518f $X=3.86 $Y=0.995 $X2=0
+ $Y2=0
cc_387 N_A_213_47#_c_307_n N_VGND_c_860_n 0.0058995f $X=4.28 $Y=0.995 $X2=0
+ $Y2=0
cc_388 N_A_213_47#_c_308_n N_VGND_c_860_n 0.0058995f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_389 N_A_213_47#_c_309_n N_VGND_c_860_n 0.0058995f $X=5.22 $Y=0.995 $X2=0
+ $Y2=0
cc_390 N_A_213_47#_c_310_n N_VGND_c_860_n 0.0058995f $X=5.74 $Y=0.995 $X2=0
+ $Y2=0
cc_391 N_A_213_47#_c_311_n N_VGND_c_860_n 0.0058995f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_392 N_A_213_47#_c_312_n N_VGND_c_860_n 0.00589754f $X=6.68 $Y=0.995 $X2=0
+ $Y2=0
cc_393 N_A_213_47#_c_313_n N_VGND_c_860_n 0.0106244f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_394 N_A_213_47#_c_329_n N_VGND_c_860_n 0.0120611f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_395 N_A_213_47#_c_331_n N_VGND_c_860_n 0.0201864f $X=2.445 $Y=0.78 $X2=0
+ $Y2=0
cc_396 N_A_213_47#_c_336_n N_VGND_c_860_n 0.0112677f $X=2.61 $Y=0.42 $X2=0 $Y2=0
cc_397 N_A_213_47#_c_358_n N_VGND_c_860_n 0.00740747f $X=3.565 $Y=0.78 $X2=0
+ $Y2=0
cc_398 N_A_213_47#_c_331_n N_VGND_c_862_n 0.00224243f $X=2.445 $Y=0.78 $X2=0
+ $Y2=0
cc_399 N_A_213_47#_c_336_n N_VGND_c_862_n 0.0169239f $X=2.61 $Y=0.42 $X2=0 $Y2=0
cc_400 N_A_213_47#_c_358_n N_VGND_c_862_n 0.00243213f $X=3.565 $Y=0.78 $X2=0
+ $Y2=0
cc_401 N_A_213_47#_c_306_n N_VGND_c_863_n 0.00853918f $X=3.86 $Y=0.995 $X2=0
+ $Y2=0
cc_402 N_A_213_47#_c_358_n N_VGND_c_863_n 0.0614132f $X=3.565 $Y=0.78 $X2=0
+ $Y2=0
cc_403 N_A_213_47#_c_331_n A_131_47# 0.00554514f $X=2.445 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_404 N_A_27_297#_c_532_n N_VPWR_M1011_d 0.00368875f $X=1.035 $Y=1.885
+ $X2=-0.19 $Y2=1.305
cc_405 N_A_27_297#_c_536_n N_VPWR_M1024_s 0.00368875f $X=1.975 $Y=1.885 $X2=0
+ $Y2=0
cc_406 N_A_27_297#_c_532_n N_VPWR_c_593_n 0.0138616f $X=1.035 $Y=1.885 $X2=0
+ $Y2=0
cc_407 N_A_27_297#_c_532_n N_VPWR_c_594_n 0.00209157f $X=1.035 $Y=1.885 $X2=0
+ $Y2=0
cc_408 N_A_27_297#_c_536_n N_VPWR_c_594_n 0.00209157f $X=1.975 $Y=1.885 $X2=0
+ $Y2=0
cc_409 N_A_27_297#_c_544_n N_VPWR_c_594_n 0.0189225f $X=1.2 $Y=1.885 $X2=0 $Y2=0
cc_410 N_A_27_297#_c_536_n N_VPWR_c_595_n 0.0138616f $X=1.975 $Y=1.885 $X2=0
+ $Y2=0
cc_411 N_A_27_297#_c_524_n N_VPWR_c_596_n 0.0113145f $X=2.915 $Y=2.38 $X2=0
+ $Y2=0
cc_412 N_A_27_297#_c_525_n N_VPWR_c_596_n 0.0318764f $X=3.08 $Y=1.87 $X2=0 $Y2=0
cc_413 N_A_27_297#_c_536_n N_VPWR_c_601_n 0.00209157f $X=1.975 $Y=1.885 $X2=0
+ $Y2=0
cc_414 N_A_27_297#_c_524_n N_VPWR_c_601_n 0.0575925f $X=2.915 $Y=2.38 $X2=0
+ $Y2=0
cc_415 N_A_27_297#_c_541_n N_VPWR_c_601_n 0.0173953f $X=2.275 $Y=2.38 $X2=0
+ $Y2=0
cc_416 N_A_27_297#_c_522_n N_VPWR_c_611_n 0.0210576f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_417 N_A_27_297#_c_532_n N_VPWR_c_611_n 0.00209157f $X=1.035 $Y=1.885 $X2=0
+ $Y2=0
cc_418 N_A_27_297#_M1011_s N_VPWR_c_592_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_419 N_A_27_297#_M1003_d N_VPWR_c_592_n 0.00231261f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_420 N_A_27_297#_M1017_s N_VPWR_c_592_n 0.00231262f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_421 N_A_27_297#_M1012_d N_VPWR_c_592_n 0.00217517f $X=2.935 $Y=1.485 $X2=0
+ $Y2=0
cc_422 N_A_27_297#_c_522_n N_VPWR_c_592_n 0.0124606f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_423 N_A_27_297#_c_532_n N_VPWR_c_592_n 0.00811004f $X=1.035 $Y=1.885 $X2=0
+ $Y2=0
cc_424 N_A_27_297#_c_536_n N_VPWR_c_592_n 0.00811004f $X=1.975 $Y=1.885 $X2=0
+ $Y2=0
cc_425 N_A_27_297#_c_524_n N_VPWR_c_592_n 0.0347586f $X=2.915 $Y=2.38 $X2=0
+ $Y2=0
cc_426 N_A_27_297#_c_541_n N_VPWR_c_592_n 0.0113829f $X=2.275 $Y=2.38 $X2=0
+ $Y2=0
cc_427 N_A_27_297#_c_544_n N_VPWR_c_592_n 0.0123059f $X=1.2 $Y=1.885 $X2=0 $Y2=0
cc_428 N_VPWR_c_592_n N_X_M1005_d 0.00300692f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_429 N_VPWR_c_592_n N_X_M1013_d 0.00300692f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_430 N_VPWR_c_592_n N_X_M1018_d 0.00300692f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_431 N_VPWR_c_592_n N_X_M1025_d 0.00300692f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_432 N_VPWR_c_603_n N_X_c_797_n 0.0156407f $X=4.375 $Y=2.72 $X2=0 $Y2=0
cc_433 N_VPWR_c_592_n N_X_c_797_n 0.0103212f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_434 N_VPWR_M1007_s N_X_c_716_n 0.00187091f $X=4.395 $Y=1.485 $X2=0 $Y2=0
cc_435 N_VPWR_c_597_n N_X_c_716_n 0.0171295f $X=4.54 $Y=1.87 $X2=0 $Y2=0
cc_436 N_VPWR_c_605_n N_X_c_801_n 0.0156407f $X=5.315 $Y=2.72 $X2=0 $Y2=0
cc_437 N_VPWR_c_592_n N_X_c_801_n 0.0103212f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_438 N_VPWR_M1015_s N_X_c_718_n 0.00187091f $X=5.335 $Y=1.485 $X2=0 $Y2=0
cc_439 N_VPWR_c_598_n N_X_c_718_n 0.0171295f $X=5.48 $Y=1.87 $X2=0 $Y2=0
cc_440 N_VPWR_c_607_n N_X_c_805_n 0.0156407f $X=6.255 $Y=2.72 $X2=0 $Y2=0
cc_441 N_VPWR_c_592_n N_X_c_805_n 0.0103212f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_442 N_VPWR_M1021_s N_X_c_719_n 0.00187091f $X=6.275 $Y=1.485 $X2=0 $Y2=0
cc_443 N_VPWR_c_599_n N_X_c_719_n 0.0171295f $X=6.42 $Y=1.87 $X2=0 $Y2=0
cc_444 N_VPWR_c_600_n N_X_c_720_n 0.00802397f $X=7.36 $Y=1.63 $X2=0 $Y2=0
cc_445 N_VPWR_c_609_n N_X_c_810_n 0.0156407f $X=7.215 $Y=2.72 $X2=0 $Y2=0
cc_446 N_VPWR_c_592_n N_X_c_810_n 0.0103212f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_447 N_VPWR_c_600_n N_VGND_c_849_n 0.0103464f $X=7.36 $Y=1.63 $X2=0 $Y2=0
cc_448 N_X_c_734_n N_VGND_M1002_s 0.00500678f $X=4.845 $Y=0.78 $X2=0 $Y2=0
cc_449 N_X_c_750_n N_VGND_M1010_s 0.00500678f $X=5.785 $Y=0.78 $X2=0 $Y2=0
cc_450 N_X_c_761_n N_VGND_M1020_s 0.00625323f $X=6.545 $Y=0.78 $X2=0 $Y2=0
cc_451 X N_VGND_M1020_s 2.58287e-19 $X=6.585 $Y=1.105 $X2=0 $Y2=0
cc_452 N_X_c_734_n N_VGND_c_846_n 0.0198794f $X=4.845 $Y=0.78 $X2=0 $Y2=0
cc_453 N_X_c_750_n N_VGND_c_847_n 0.0198794f $X=5.785 $Y=0.78 $X2=0 $Y2=0
cc_454 N_X_c_761_n N_VGND_c_848_n 0.019613f $X=6.545 $Y=0.78 $X2=0 $Y2=0
cc_455 N_X_c_782_n N_VGND_c_848_n 2.57371e-19 $X=6.8 $Y=0.78 $X2=0 $Y2=0
cc_456 X N_VGND_c_849_n 7.9475e-19 $X=6.585 $Y=1.105 $X2=0 $Y2=0
cc_457 N_X_c_724_n N_VGND_c_850_n 0.018787f $X=4.07 $Y=0.36 $X2=0 $Y2=0
cc_458 N_X_c_734_n N_VGND_c_850_n 0.00211912f $X=4.845 $Y=0.78 $X2=0 $Y2=0
cc_459 N_X_c_734_n N_VGND_c_852_n 0.00211912f $X=4.845 $Y=0.78 $X2=0 $Y2=0
cc_460 N_X_c_742_n N_VGND_c_852_n 0.018787f $X=5.01 $Y=0.36 $X2=0 $Y2=0
cc_461 N_X_c_750_n N_VGND_c_852_n 0.00211912f $X=5.785 $Y=0.78 $X2=0 $Y2=0
cc_462 N_X_c_750_n N_VGND_c_854_n 0.00211912f $X=5.785 $Y=0.78 $X2=0 $Y2=0
cc_463 N_X_c_754_n N_VGND_c_854_n 0.018787f $X=5.95 $Y=0.36 $X2=0 $Y2=0
cc_464 N_X_c_761_n N_VGND_c_854_n 0.00211912f $X=6.545 $Y=0.78 $X2=0 $Y2=0
cc_465 N_X_c_764_n N_VGND_c_856_n 0.018802f $X=6.89 $Y=0.36 $X2=0 $Y2=0
cc_466 N_X_c_782_n N_VGND_c_856_n 0.00229847f $X=6.8 $Y=0.78 $X2=0 $Y2=0
cc_467 N_X_M1001_d N_VGND_c_860_n 0.00215201f $X=3.935 $Y=0.235 $X2=0 $Y2=0
cc_468 N_X_M1006_d N_VGND_c_860_n 0.00215201f $X=4.875 $Y=0.235 $X2=0 $Y2=0
cc_469 N_X_M1019_d N_VGND_c_860_n 0.00215201f $X=5.815 $Y=0.235 $X2=0 $Y2=0
cc_470 N_X_M1022_d N_VGND_c_860_n 0.00215201f $X=6.755 $Y=0.235 $X2=0 $Y2=0
cc_471 N_X_c_724_n N_VGND_c_860_n 0.0121864f $X=4.07 $Y=0.36 $X2=0 $Y2=0
cc_472 N_X_c_734_n N_VGND_c_860_n 0.00897448f $X=4.845 $Y=0.78 $X2=0 $Y2=0
cc_473 N_X_c_742_n N_VGND_c_860_n 0.0121864f $X=5.01 $Y=0.36 $X2=0 $Y2=0
cc_474 N_X_c_750_n N_VGND_c_860_n 0.00897448f $X=5.785 $Y=0.78 $X2=0 $Y2=0
cc_475 N_X_c_754_n N_VGND_c_860_n 0.0121864f $X=5.95 $Y=0.36 $X2=0 $Y2=0
cc_476 N_X_c_761_n N_VGND_c_860_n 0.00498522f $X=6.545 $Y=0.78 $X2=0 $Y2=0
cc_477 N_X_c_764_n N_VGND_c_860_n 0.0121937f $X=6.89 $Y=0.36 $X2=0 $Y2=0
cc_478 N_X_c_782_n N_VGND_c_860_n 0.00427984f $X=6.8 $Y=0.78 $X2=0 $Y2=0
cc_479 N_VGND_c_860_n A_297_47# 0.0111139f $X=7.59 $Y=0 $X2=-0.19 $Y2=-0.24
cc_480 N_VGND_c_860_n A_131_47# 0.00318778f $X=7.59 $Y=0 $X2=-0.19 $Y2=-0.24
