* File: sky130_fd_sc_hdll__nand2b_2.pxi.spice
* Created: Wed Sep  2 08:37:19 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND2B_2%A_N N_A_N_c_51_n N_A_N_M1009_g N_A_N_c_52_n
+ N_A_N_M1006_g A_N A_N PM_SKY130_FD_SC_HDLL__NAND2B_2%A_N
x_PM_SKY130_FD_SC_HDLL__NAND2B_2%A_27_93# N_A_27_93#_M1009_s N_A_27_93#_M1006_s
+ N_A_27_93#_c_82_n N_A_27_93#_M1001_g N_A_27_93#_M1000_g N_A_27_93#_c_83_n
+ N_A_27_93#_M1007_g N_A_27_93#_M1002_g N_A_27_93#_c_78_n N_A_27_93#_c_93_n
+ N_A_27_93#_c_79_n N_A_27_93#_c_80_n N_A_27_93#_c_86_n N_A_27_93#_c_81_n
+ PM_SKY130_FD_SC_HDLL__NAND2B_2%A_27_93#
x_PM_SKY130_FD_SC_HDLL__NAND2B_2%B N_B_c_140_n N_B_M1004_g N_B_M1003_g
+ N_B_c_141_n N_B_M1008_g N_B_M1005_g B B B N_B_c_139_n B
+ PM_SKY130_FD_SC_HDLL__NAND2B_2%B
x_PM_SKY130_FD_SC_HDLL__NAND2B_2%VPWR N_VPWR_M1006_d N_VPWR_M1007_d
+ N_VPWR_M1008_d N_VPWR_c_188_n N_VPWR_c_189_n N_VPWR_c_190_n N_VPWR_c_191_n
+ N_VPWR_c_192_n N_VPWR_c_193_n VPWR N_VPWR_c_194_n N_VPWR_c_195_n
+ N_VPWR_c_187_n PM_SKY130_FD_SC_HDLL__NAND2B_2%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND2B_2%Y N_Y_M1000_s N_Y_M1001_s N_Y_M1004_s
+ N_Y_c_233_n N_Y_c_234_n N_Y_c_246_n N_Y_c_237_n Y Y Y Y N_Y_c_231_n Y
+ PM_SKY130_FD_SC_HDLL__NAND2B_2%Y
x_PM_SKY130_FD_SC_HDLL__NAND2B_2%VGND N_VGND_M1009_d N_VGND_M1003_s
+ N_VGND_c_275_n N_VGND_c_276_n N_VGND_c_277_n N_VGND_c_278_n VGND
+ N_VGND_c_279_n N_VGND_c_280_n N_VGND_c_281_n N_VGND_c_282_n
+ PM_SKY130_FD_SC_HDLL__NAND2B_2%VGND
x_PM_SKY130_FD_SC_HDLL__NAND2B_2%A_215_47# N_A_215_47#_M1000_d
+ N_A_215_47#_M1002_d N_A_215_47#_M1005_d N_A_215_47#_c_319_n
+ N_A_215_47#_c_327_n N_A_215_47#_c_320_n N_A_215_47#_c_321_n
+ N_A_215_47#_c_322_n PM_SKY130_FD_SC_HDLL__NAND2B_2%A_215_47#
cc_1 VNB N_A_N_c_51_n 0.0242977f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_N_c_52_n 0.0275905f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_3 VNB A_N 0.00546266f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_4 VNB N_A_27_93#_M1000_g 0.0232023f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.16
cc_5 VNB N_A_27_93#_M1002_g 0.017197f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_93#_c_78_n 0.0213871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_93#_c_79_n 0.00340013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_93#_c_80_n 0.0123578f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_93#_c_81_n 0.0725464f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B_M1003_g 0.0180965f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.695
cc_11 VNB N_B_M1005_g 0.0244194f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB B 0.0161406f $X=-0.19 $Y=-0.24 $X2=0.745 $Y2=1.16
cc_13 VNB B 0.00141012f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_B_c_139_n 0.0449304f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VPWR_c_187_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_275_n 0.0127513f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=1.16
cc_17 VNB N_VGND_c_276_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_277_n 0.0405294f $X=-0.19 $Y=-0.24 $X2=0.745 $Y2=1.16
cc_19 VNB N_VGND_c_278_n 0.00323881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_279_n 0.0197486f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_280_n 0.0181414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_281_n 0.203025f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_282_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_215_47#_c_319_n 0.00303415f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.16
cc_25 VNB N_A_215_47#_c_320_n 0.00681087f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_26 VNB N_A_215_47#_c_321_n 0.0142118f $X=-0.19 $Y=-0.24 $X2=0.745 $Y2=1.16
cc_27 VNB N_A_215_47#_c_322_n 0.0172779f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VPB N_A_N_c_52_n 0.0331179f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_29 VPB A_N 0.00127365f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_30 VPB N_A_27_93#_c_82_n 0.0193086f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_31 VPB N_A_27_93#_c_83_n 0.017309f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.16
cc_32 VPB N_A_27_93#_c_78_n 0.00899582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A_27_93#_c_79_n 0.00132417f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_27_93#_c_86_n 0.0153447f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_27_93#_c_81_n 0.0128857f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_B_c_140_n 0.0177189f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_37 VPB N_B_c_141_n 0.0192593f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB B 0.0158653f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_B_c_139_n 0.014484f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_188_n 0.0235272f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.16
cc_41 VPB N_VPWR_c_189_n 0.00588144f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_190_n 0.0119842f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_191_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_192_n 0.0225792f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_193_n 0.00718421f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_194_n 0.0196192f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_195_n 0.0270701f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_187_n 0.0633335f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_Y_c_231_n 0.00351661f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 N_A_N_c_52_n N_A_27_93#_c_82_n 0.0164156f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_51 N_A_N_c_52_n N_A_27_93#_M1000_g 3.59662e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_52 N_A_N_c_51_n N_A_27_93#_c_78_n 0.0161951f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_53 N_A_N_c_52_n N_A_27_93#_c_78_n 0.00310122f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_54 A_N N_A_27_93#_c_78_n 0.0245673f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_55 N_A_N_c_52_n N_A_27_93#_c_93_n 0.0187674f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_56 A_N N_A_27_93#_c_93_n 0.0272949f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_57 N_A_N_c_52_n N_A_27_93#_c_79_n 0.00123604f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_58 A_N N_A_27_93#_c_79_n 0.0253713f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_59 N_A_N_c_52_n N_A_27_93#_c_86_n 0.0037072f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_60 N_A_N_c_52_n N_A_27_93#_c_81_n 0.0224545f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_61 A_N N_A_27_93#_c_81_n 0.00222183f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_62 N_A_N_c_52_n N_VPWR_c_188_n 0.00392799f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_63 N_A_N_c_52_n N_VPWR_c_195_n 0.00393512f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_64 N_A_N_c_52_n N_VPWR_c_187_n 0.00500987f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_65 N_A_N_c_51_n N_VGND_c_275_n 0.00505361f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_66 N_A_N_c_52_n N_VGND_c_275_n 0.00290622f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_67 A_N N_VGND_c_275_n 0.0113158f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_68 N_A_N_c_51_n N_VGND_c_279_n 0.00510437f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_69 N_A_N_c_51_n N_VGND_c_281_n 0.00512902f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_70 N_A_27_93#_c_83_n N_B_c_140_n 0.024863f $X=1.565 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_71 N_A_27_93#_M1002_g N_B_M1003_g 0.0132767f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_72 N_A_27_93#_c_81_n B 0.00169515f $X=1.565 $Y=1.217 $X2=0 $Y2=0
cc_73 N_A_27_93#_c_81_n N_B_c_139_n 0.0213215f $X=1.565 $Y=1.217 $X2=0 $Y2=0
cc_74 N_A_27_93#_c_93_n N_VPWR_M1006_d 0.00604907f $X=1.02 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_75 N_A_27_93#_c_82_n N_VPWR_c_188_n 0.00752789f $X=1.035 $Y=1.41 $X2=0 $Y2=0
cc_76 N_A_27_93#_c_93_n N_VPWR_c_188_n 0.0196888f $X=1.02 $Y=1.58 $X2=0 $Y2=0
cc_77 N_A_27_93#_c_83_n N_VPWR_c_189_n 0.00689826f $X=1.565 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A_27_93#_c_82_n N_VPWR_c_192_n 0.00702461f $X=1.035 $Y=1.41 $X2=0 $Y2=0
cc_79 N_A_27_93#_c_83_n N_VPWR_c_192_n 0.00523619f $X=1.565 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A_27_93#_c_82_n N_VPWR_c_187_n 0.0139371f $X=1.035 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_27_93#_c_83_n N_VPWR_c_187_n 0.00750777f $X=1.565 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A_27_93#_c_93_n N_Y_M1001_s 0.00193341f $X=1.02 $Y=1.58 $X2=0 $Y2=0
cc_83 N_A_27_93#_c_81_n N_Y_c_233_n 0.00337255f $X=1.565 $Y=1.217 $X2=0 $Y2=0
cc_84 N_A_27_93#_c_83_n N_Y_c_234_n 0.0102419f $X=1.565 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A_27_93#_c_93_n N_Y_c_234_n 6.71458e-19 $X=1.02 $Y=1.58 $X2=0 $Y2=0
cc_86 N_A_27_93#_c_81_n N_Y_c_234_n 0.00765408f $X=1.565 $Y=1.217 $X2=0 $Y2=0
cc_87 N_A_27_93#_c_83_n N_Y_c_237_n 7.80904e-19 $X=1.565 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A_27_93#_c_82_n N_Y_c_231_n 3.84971e-19 $X=1.035 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A_27_93#_M1000_g N_Y_c_231_n 0.0181396f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_90 N_A_27_93#_c_83_n N_Y_c_231_n 0.0136191f $X=1.565 $Y=1.41 $X2=0 $Y2=0
cc_91 N_A_27_93#_M1002_g N_Y_c_231_n 0.00702384f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_92 N_A_27_93#_c_79_n N_Y_c_231_n 0.0263774f $X=1.105 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_27_93#_c_81_n N_Y_c_231_n 0.0260976f $X=1.565 $Y=1.217 $X2=0 $Y2=0
cc_94 N_A_27_93#_M1000_g N_VGND_c_275_n 0.0077417f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_95 N_A_27_93#_M1000_g N_VGND_c_277_n 0.00357877f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_96 N_A_27_93#_M1002_g N_VGND_c_277_n 0.00357877f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_97 N_A_27_93#_c_80_n N_VGND_c_279_n 0.00593412f $X=0.26 $Y=0.675 $X2=0 $Y2=0
cc_98 N_A_27_93#_M1000_g N_VGND_c_281_n 0.00655123f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_99 N_A_27_93#_M1002_g N_VGND_c_281_n 0.00525237f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_100 N_A_27_93#_c_80_n N_VGND_c_281_n 0.00761143f $X=0.26 $Y=0.675 $X2=0 $Y2=0
cc_101 N_A_27_93#_M1000_g N_A_215_47#_c_319_n 0.0124471f $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_102 N_A_27_93#_M1002_g N_A_215_47#_c_319_n 0.0124471f $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_103 N_A_27_93#_c_79_n N_A_215_47#_c_319_n 0.00579922f $X=1.105 $Y=1.16 $X2=0
+ $Y2=0
cc_104 N_A_27_93#_c_81_n N_A_215_47#_c_319_n 0.00404198f $X=1.565 $Y=1.217 $X2=0
+ $Y2=0
cc_105 B N_VPWR_M1008_d 0.00699604f $X=2.915 $Y=1.445 $X2=0 $Y2=0
cc_106 N_B_c_140_n N_VPWR_c_189_n 0.00560707f $X=2.215 $Y=1.41 $X2=0 $Y2=0
cc_107 N_B_c_141_n N_VPWR_c_191_n 0.00697547f $X=2.695 $Y=1.41 $X2=0 $Y2=0
cc_108 B N_VPWR_c_191_n 0.00206711f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_109 B N_VPWR_c_191_n 0.00921873f $X=2.915 $Y=1.445 $X2=0 $Y2=0
cc_110 N_B_c_140_n N_VPWR_c_194_n 0.00514793f $X=2.215 $Y=1.41 $X2=0 $Y2=0
cc_111 N_B_c_141_n N_VPWR_c_194_n 0.00688798f $X=2.695 $Y=1.41 $X2=0 $Y2=0
cc_112 N_B_c_140_n N_VPWR_c_187_n 0.00716634f $X=2.215 $Y=1.41 $X2=0 $Y2=0
cc_113 N_B_c_141_n N_VPWR_c_187_n 0.0131773f $X=2.695 $Y=1.41 $X2=0 $Y2=0
cc_114 N_B_c_140_n N_Y_c_233_n 0.0135455f $X=2.215 $Y=1.41 $X2=0 $Y2=0
cc_115 B N_Y_c_233_n 0.00432305f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_116 N_B_c_141_n N_Y_c_246_n 0.00973393f $X=2.695 $Y=1.41 $X2=0 $Y2=0
cc_117 B N_Y_c_246_n 0.0149129f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_118 B N_Y_c_246_n 0.00779671f $X=2.915 $Y=1.445 $X2=0 $Y2=0
cc_119 N_B_c_139_n N_Y_c_246_n 0.00596949f $X=2.695 $Y=1.217 $X2=0 $Y2=0
cc_120 N_B_c_140_n N_Y_c_237_n 0.00780325f $X=2.215 $Y=1.41 $X2=0 $Y2=0
cc_121 N_B_c_141_n N_Y_c_237_n 0.00755651f $X=2.695 $Y=1.41 $X2=0 $Y2=0
cc_122 B N_Y_c_237_n 0.00101442f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_123 N_B_c_140_n N_Y_c_231_n 0.00491505f $X=2.215 $Y=1.41 $X2=0 $Y2=0
cc_124 N_B_M1003_g N_Y_c_231_n 6.76644e-19 $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_125 B N_Y_c_231_n 0.0103076f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_126 N_B_c_139_n N_Y_c_231_n 0.00304806f $X=2.695 $Y=1.217 $X2=0 $Y2=0
cc_127 N_B_M1003_g N_VGND_c_276_n 0.00369356f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_128 N_B_M1005_g N_VGND_c_276_n 0.00276126f $X=2.72 $Y=0.56 $X2=0 $Y2=0
cc_129 N_B_M1003_g N_VGND_c_277_n 0.00418507f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_130 N_B_M1005_g N_VGND_c_280_n 0.00420025f $X=2.72 $Y=0.56 $X2=0 $Y2=0
cc_131 N_B_M1003_g N_VGND_c_281_n 0.00594321f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_132 N_B_M1005_g N_VGND_c_281_n 0.00676597f $X=2.72 $Y=0.56 $X2=0 $Y2=0
cc_133 N_B_M1003_g N_A_215_47#_c_327_n 0.00271016f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_134 N_B_M1003_g N_A_215_47#_c_320_n 0.00498742f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_135 N_B_M1005_g N_A_215_47#_c_320_n 4.68334e-19 $X=2.72 $Y=0.56 $X2=0 $Y2=0
cc_136 B N_A_215_47#_c_320_n 0.0076014f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_137 N_B_c_139_n N_A_215_47#_c_320_n 0.00169611f $X=2.695 $Y=1.217 $X2=0 $Y2=0
cc_138 N_B_M1003_g N_A_215_47#_c_321_n 0.00967151f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_139 N_B_M1005_g N_A_215_47#_c_321_n 0.0109805f $X=2.72 $Y=0.56 $X2=0 $Y2=0
cc_140 B N_A_215_47#_c_321_n 0.0693881f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_141 N_B_c_139_n N_A_215_47#_c_321_n 0.00321256f $X=2.695 $Y=1.217 $X2=0 $Y2=0
cc_142 N_B_M1003_g N_A_215_47#_c_322_n 5.17586e-19 $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_143 N_B_M1005_g N_A_215_47#_c_322_n 0.00620156f $X=2.72 $Y=0.56 $X2=0 $Y2=0
cc_144 N_VPWR_c_187_n N_Y_M1001_s 0.00315011f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_145 N_VPWR_c_187_n N_Y_M1004_s 0.00239291f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_146 N_VPWR_M1007_d N_Y_c_233_n 0.0120611f $X=1.655 $Y=1.485 $X2=0 $Y2=0
cc_147 N_VPWR_c_189_n N_Y_c_233_n 0.0220603f $X=1.92 $Y=2.34 $X2=0 $Y2=0
cc_148 N_VPWR_c_194_n N_Y_c_233_n 0.00237402f $X=2.845 $Y=2.72 $X2=0 $Y2=0
cc_149 N_VPWR_c_187_n N_Y_c_233_n 0.00533331f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_150 N_VPWR_M1007_d N_Y_c_234_n 8.8477e-19 $X=1.655 $Y=1.485 $X2=0 $Y2=0
cc_151 N_VPWR_c_189_n N_Y_c_234_n 0.00504736f $X=1.92 $Y=2.34 $X2=0 $Y2=0
cc_152 N_VPWR_c_192_n N_Y_c_234_n 0.023283f $X=1.725 $Y=2.72 $X2=0 $Y2=0
cc_153 N_VPWR_c_187_n N_Y_c_234_n 0.0193719f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_154 N_VPWR_c_191_n N_Y_c_237_n 0.0374578f $X=2.93 $Y=2 $X2=0 $Y2=0
cc_155 N_VPWR_c_194_n N_Y_c_237_n 0.0189613f $X=2.845 $Y=2.72 $X2=0 $Y2=0
cc_156 N_VPWR_c_187_n N_Y_c_237_n 0.0123549f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_157 N_VPWR_M1007_d N_Y_c_231_n 0.00483788f $X=1.655 $Y=1.485 $X2=0 $Y2=0
cc_158 N_Y_M1000_s N_VGND_c_281_n 0.00216833f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_159 N_Y_M1000_s N_A_215_47#_c_319_n 0.00305226f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_160 N_Y_c_231_n N_A_215_47#_c_319_n 0.016329f $X=1.62 $Y=0.72 $X2=0 $Y2=0
cc_161 N_Y_c_231_n N_A_215_47#_c_320_n 0.00880289f $X=1.62 $Y=0.72 $X2=0 $Y2=0
cc_162 N_VGND_c_281_n N_A_215_47#_M1000_d 0.00209344f $X=2.99 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_163 N_VGND_c_281_n N_A_215_47#_M1002_d 0.00215206f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_164 N_VGND_c_281_n N_A_215_47#_M1005_d 0.00209319f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_165 N_VGND_c_275_n N_A_215_47#_c_319_n 0.0127155f $X=0.68 $Y=0.61 $X2=0 $Y2=0
cc_166 N_VGND_c_277_n N_A_215_47#_c_319_n 0.0521531f $X=2.425 $Y=0 $X2=0 $Y2=0
cc_167 N_VGND_c_281_n N_A_215_47#_c_319_n 0.0329109f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_168 N_VGND_c_276_n N_A_215_47#_c_327_n 0.0135136f $X=2.51 $Y=0.36 $X2=0 $Y2=0
cc_169 N_VGND_c_277_n N_A_215_47#_c_327_n 0.0152108f $X=2.425 $Y=0 $X2=0 $Y2=0
cc_170 N_VGND_c_281_n N_A_215_47#_c_327_n 0.00940698f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_171 N_VGND_c_276_n N_A_215_47#_c_320_n 0.003527f $X=2.51 $Y=0.36 $X2=0 $Y2=0
cc_172 N_VGND_M1003_s N_A_215_47#_c_321_n 0.00249128f $X=2.325 $Y=0.235 $X2=0
+ $Y2=0
cc_173 N_VGND_c_276_n N_A_215_47#_c_321_n 0.0127545f $X=2.51 $Y=0.36 $X2=0 $Y2=0
cc_174 N_VGND_c_277_n N_A_215_47#_c_321_n 0.00287272f $X=2.425 $Y=0 $X2=0 $Y2=0
cc_175 N_VGND_c_280_n N_A_215_47#_c_321_n 0.00214238f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_176 N_VGND_c_281_n N_A_215_47#_c_321_n 0.0100688f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_177 N_VGND_c_280_n N_A_215_47#_c_322_n 0.0209752f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_178 N_VGND_c_281_n N_A_215_47#_c_322_n 0.0124119f $X=2.99 $Y=0 $X2=0 $Y2=0
