* File: sky130_fd_sc_hdll__o32ai_4.pxi.spice
* Created: Thu Aug 27 19:23:00 2020
* 
x_PM_SKY130_FD_SC_HDLL__O32AI_4%B2 N_B2_c_136_n N_B2_M1002_g N_B2_M1004_g
+ N_B2_c_137_n N_B2_M1016_g N_B2_M1026_g N_B2_c_138_n N_B2_M1025_g N_B2_M1027_g
+ N_B2_c_139_n N_B2_M1036_g N_B2_M1038_g B2 B2 B2 N_B2_c_134_n N_B2_c_135_n B2
+ PM_SKY130_FD_SC_HDLL__O32AI_4%B2
x_PM_SKY130_FD_SC_HDLL__O32AI_4%B1 N_B1_M1005_g N_B1_c_209_n N_B1_M1000_g
+ N_B1_M1024_g N_B1_c_210_n N_B1_M1007_g N_B1_M1028_g N_B1_c_211_n N_B1_M1022_g
+ N_B1_c_212_n N_B1_M1034_g N_B1_M1039_g B1 B1 B1 N_B1_c_207_n N_B1_c_208_n B1
+ B1 B1 PM_SKY130_FD_SC_HDLL__O32AI_4%B1
x_PM_SKY130_FD_SC_HDLL__O32AI_4%A3 N_A3_M1012_g N_A3_M1013_g N_A3_c_279_n
+ N_A3_M1011_g N_A3_M1017_g N_A3_c_280_n N_A3_M1021_g N_A3_c_281_n N_A3_M1029_g
+ N_A3_M1031_g N_A3_c_282_n N_A3_M1037_g N_A3_c_275_n A3 A3 A3 A3 N_A3_c_277_n
+ N_A3_c_278_n A3 A3 A3 A3 PM_SKY130_FD_SC_HDLL__O32AI_4%A3
x_PM_SKY130_FD_SC_HDLL__O32AI_4%A2 N_A2_M1006_g N_A2_c_364_n N_A2_M1001_g
+ N_A2_M1009_g N_A2_c_365_n N_A2_M1008_g N_A2_M1019_g N_A2_c_366_n N_A2_M1014_g
+ N_A2_c_367_n N_A2_M1018_g N_A2_M1033_g A2 A2 A2 N_A2_c_362_n N_A2_c_363_n A2
+ A2 A2 PM_SKY130_FD_SC_HDLL__O32AI_4%A2
x_PM_SKY130_FD_SC_HDLL__O32AI_4%A1 N_A1_M1015_g N_A1_c_443_n N_A1_M1003_g
+ N_A1_M1020_g N_A1_c_444_n N_A1_M1010_g N_A1_M1032_g N_A1_c_445_n N_A1_M1023_g
+ N_A1_c_438_n N_A1_c_439_n N_A1_M1035_g N_A1_c_448_n N_A1_M1030_g A1 A1 A1 A1
+ N_A1_c_442_n A1 A1 A1 PM_SKY130_FD_SC_HDLL__O32AI_4%A1
x_PM_SKY130_FD_SC_HDLL__O32AI_4%A_27_297# N_A_27_297#_M1002_d
+ N_A_27_297#_M1016_d N_A_27_297#_M1036_d N_A_27_297#_M1007_d
+ N_A_27_297#_M1034_d N_A_27_297#_c_513_n N_A_27_297#_c_514_n
+ N_A_27_297#_c_519_n N_A_27_297#_c_534_p N_A_27_297#_c_521_n
+ N_A_27_297#_c_552_p N_A_27_297#_c_525_n N_A_27_297#_c_523_n
+ N_A_27_297#_c_559_p N_A_27_297#_c_527_n N_A_27_297#_c_515_n
+ N_A_27_297#_c_516_n N_A_27_297#_c_569_p N_A_27_297#_c_543_p
+ PM_SKY130_FD_SC_HDLL__O32AI_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__O32AI_4%Y N_Y_M1004_s N_Y_M1027_s N_Y_M1005_s
+ N_Y_M1028_s N_Y_M1002_s N_Y_M1025_s N_Y_M1011_d N_Y_M1029_d N_Y_c_590_n
+ N_Y_c_601_n N_Y_c_605_n N_Y_c_591_n N_Y_c_592_n N_Y_c_594_n N_Y_c_640_n
+ N_Y_c_609_n N_Y_c_614_n N_Y_c_702_p N_Y_c_672_n N_Y_c_644_n N_Y_c_649_n Y
+ PM_SKY130_FD_SC_HDLL__O32AI_4%Y
x_PM_SKY130_FD_SC_HDLL__O32AI_4%VPWR N_VPWR_M1000_s N_VPWR_M1022_s
+ N_VPWR_M1003_s N_VPWR_M1010_s N_VPWR_M1030_s N_VPWR_c_720_n N_VPWR_c_721_n
+ N_VPWR_c_722_n N_VPWR_c_723_n N_VPWR_c_724_n N_VPWR_c_725_n N_VPWR_c_726_n
+ N_VPWR_c_727_n N_VPWR_c_728_n N_VPWR_c_729_n VPWR N_VPWR_c_730_n
+ N_VPWR_c_731_n N_VPWR_c_732_n N_VPWR_c_733_n N_VPWR_c_734_n N_VPWR_c_719_n
+ PM_SKY130_FD_SC_HDLL__O32AI_4%VPWR
x_PM_SKY130_FD_SC_HDLL__O32AI_4%A_886_297# N_A_886_297#_M1011_s
+ N_A_886_297#_M1021_s N_A_886_297#_M1037_s N_A_886_297#_M1008_s
+ N_A_886_297#_M1018_s N_A_886_297#_c_868_n N_A_886_297#_c_869_n
+ N_A_886_297#_c_872_n N_A_886_297#_c_891_n N_A_886_297#_c_874_n
+ N_A_886_297#_c_897_n N_A_886_297#_c_876_n N_A_886_297#_c_927_p
+ N_A_886_297#_c_878_n N_A_886_297#_c_870_n N_A_886_297#_c_871_n
+ N_A_886_297#_c_917_n N_A_886_297#_c_919_n N_A_886_297#_c_921_n
+ PM_SKY130_FD_SC_HDLL__O32AI_4%A_886_297#
x_PM_SKY130_FD_SC_HDLL__O32AI_4%A_1352_297# N_A_1352_297#_M1001_d
+ N_A_1352_297#_M1014_d N_A_1352_297#_M1003_d N_A_1352_297#_M1023_d
+ N_A_1352_297#_c_940_n N_A_1352_297#_c_938_n N_A_1352_297#_c_956_n
+ N_A_1352_297#_c_959_n N_A_1352_297#_c_963_n N_A_1352_297#_c_966_n
+ N_A_1352_297#_c_939_n N_A_1352_297#_c_950_n N_A_1352_297#_c_968_n
+ PM_SKY130_FD_SC_HDLL__O32AI_4%A_1352_297#
x_PM_SKY130_FD_SC_HDLL__O32AI_4%A_27_47# N_A_27_47#_M1004_d N_A_27_47#_M1026_d
+ N_A_27_47#_M1038_d N_A_27_47#_M1024_d N_A_27_47#_M1039_d N_A_27_47#_M1013_d
+ N_A_27_47#_M1031_d N_A_27_47#_M1009_d N_A_27_47#_M1033_d N_A_27_47#_M1020_d
+ N_A_27_47#_M1035_d N_A_27_47#_c_1004_n N_A_27_47#_c_1005_n N_A_27_47#_c_1022_n
+ N_A_27_47#_c_1033_n N_A_27_47#_c_1006_n N_A_27_47#_c_1007_n
+ N_A_27_47#_c_1041_n N_A_27_47#_c_1008_n N_A_27_47#_c_1056_n
+ N_A_27_47#_c_1009_n N_A_27_47#_c_1077_n N_A_27_47#_c_1010_n
+ N_A_27_47#_c_1011_n N_A_27_47#_c_1012_n N_A_27_47#_c_1013_n
+ N_A_27_47#_c_1014_n N_A_27_47#_c_1015_n N_A_27_47#_c_1016_n
+ N_A_27_47#_c_1017_n N_A_27_47#_c_1018_n PM_SKY130_FD_SC_HDLL__O32AI_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__O32AI_4%VGND N_VGND_M1012_s N_VGND_M1017_s
+ N_VGND_M1006_s N_VGND_M1019_s N_VGND_M1015_s N_VGND_M1032_s N_VGND_c_1176_n
+ N_VGND_c_1177_n N_VGND_c_1178_n N_VGND_c_1179_n N_VGND_c_1180_n
+ N_VGND_c_1181_n N_VGND_c_1182_n N_VGND_c_1183_n N_VGND_c_1184_n
+ N_VGND_c_1185_n N_VGND_c_1186_n N_VGND_c_1187_n N_VGND_c_1188_n
+ N_VGND_c_1189_n N_VGND_c_1190_n N_VGND_c_1191_n N_VGND_c_1192_n
+ N_VGND_c_1193_n VGND N_VGND_c_1194_n N_VGND_c_1195_n
+ PM_SKY130_FD_SC_HDLL__O32AI_4%VGND
cc_1 VNB N_B2_M1004_g 0.0234929f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_2 VNB N_B2_M1026_g 0.0178489f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_3 VNB N_B2_M1027_g 0.0178244f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_4 VNB N_B2_M1038_g 0.0176682f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_5 VNB N_B2_c_134_n 0.00806404f $X=-0.19 $Y=-0.24 $X2=1.67 $Y2=1.16
cc_6 VNB N_B2_c_135_n 0.093221f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.212
cc_7 VNB N_B1_M1005_g 0.0176684f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_8 VNB N_B1_M1024_g 0.0178246f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_9 VNB N_B1_M1028_g 0.0183265f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_10 VNB N_B1_M1039_g 0.0182733f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_11 VNB N_B1_c_207_n 0.00242518f $X=-0.19 $Y=-0.24 $X2=1.67 $Y2=1.16
cc_12 VNB N_B1_c_208_n 0.0705577f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.212
cc_13 VNB N_A3_M1012_g 0.0175554f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_14 VNB N_A3_M1013_g 0.0178447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A3_M1017_g 0.019236f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A3_M1031_g 0.0220017f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_17 VNB N_A3_c_275_n 0.00897557f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_18 VNB A3 0.00140887f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A3_c_277_n 0.0130289f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.212
cc_20 VNB N_A3_c_278_n 0.0768683f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A2_M1006_g 0.0206103f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_22 VNB N_A2_M1009_g 0.0178447f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_23 VNB N_A2_M1019_g 0.0183223f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_24 VNB N_A2_M1033_g 0.0240946f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_25 VNB N_A2_c_362_n 0.00411926f $X=-0.19 $Y=-0.24 $X2=1.67 $Y2=1.16
cc_26 VNB N_A2_c_363_n 0.0808208f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.212
cc_27 VNB N_A1_M1015_g 0.023617f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_28 VNB N_A1_M1020_g 0.0178447f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_29 VNB N_A1_M1032_g 0.0182764f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_30 VNB N_A1_c_438_n 0.0139169f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_31 VNB N_A1_c_439_n 0.057597f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_32 VNB N_A1_M1035_g 0.0240303f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_33 VNB A1 0.00988511f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A1_c_442_n 0.0292002f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.175
cc_35 VNB N_Y_c_590_n 0.00825728f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.015
cc_36 VNB N_Y_c_591_n 0.00744161f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.212
cc_37 VNB N_Y_c_592_n 0.00852537f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.212
cc_38 VNB N_VPWR_c_719_n 0.459507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_27_47#_c_1004_n 0.00922242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_27_47#_c_1005_n 0.0184553f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_41 VNB N_A_27_47#_c_1006_n 0.00370005f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.212
cc_42 VNB N_A_27_47#_c_1007_n 0.00247521f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.212
cc_43 VNB N_A_27_47#_c_1008_n 0.00247521f $X=-0.19 $Y=-0.24 $X2=1.165 $Y2=1.175
cc_44 VNB N_A_27_47#_c_1009_n 0.00450643f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_27_47#_c_1010_n 0.0123645f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_27_47#_c_1011_n 0.0191373f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_27_47#_c_1012_n 0.00252813f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_27_47#_c_1013_n 0.00357456f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_27_47#_c_1014_n 0.0132745f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_27_47#_c_1015_n 0.00252813f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_27_47#_c_1016_n 0.00289984f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_27_47#_c_1017_n 0.011017f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_27_47#_c_1018_n 0.00252813f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1176_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_1177_n 0.00563047f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.015
cc_56 VNB N_VGND_c_1178_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_57 VNB N_VGND_c_1179_n 0.00469188f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1180_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_59 VNB N_VGND_c_1181_n 0.00493975f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.212
cc_60 VNB N_VGND_c_1182_n 0.102171f $X=-0.19 $Y=-0.24 $X2=1.67 $Y2=1.212
cc_61 VNB N_VGND_c_1183_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=1.67 $Y2=1.16
cc_62 VNB N_VGND_c_1184_n 0.0192031f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.212
cc_63 VNB N_VGND_c_1185_n 0.006319f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.212
cc_64 VNB N_VGND_c_1186_n 0.0278283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1187_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1188_n 0.0192031f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1189_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.175
cc_68 VNB N_VGND_c_1190_n 0.0319176f $X=-0.19 $Y=-0.24 $X2=1.165 $Y2=1.175
cc_69 VNB N_VGND_c_1191_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=1.67 $Y2=1.175
cc_70 VNB N_VGND_c_1192_n 0.0192031f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1193_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1194_n 0.0189951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1195_n 0.506619f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VPB N_B2_c_136_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_75 VPB N_B2_c_137_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_76 VPB N_B2_c_138_n 0.016261f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_77 VPB N_B2_c_139_n 0.0165318f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_78 VPB N_B2_c_135_n 0.0577082f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.212
cc_79 VPB N_B1_c_209_n 0.0160813f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_80 VPB N_B1_c_210_n 0.0160897f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_81 VPB N_B1_c_211_n 0.0158129f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_82 VPB N_B1_c_212_n 0.0209165f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_83 VPB N_B1_c_208_n 0.0491191f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.212
cc_84 VPB N_A3_c_279_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_85 VPB N_A3_c_280_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_86 VPB N_A3_c_281_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_87 VPB N_A3_c_282_n 0.016445f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.56
cc_88 VPB N_A3_c_275_n 0.00397253f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_89 VPB N_A3_c_277_n 0.00809277f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.212
cc_90 VPB N_A3_c_278_n 0.0502939f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A2_c_364_n 0.016445f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_92 VPB N_A2_c_365_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_93 VPB N_A2_c_366_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_94 VPB N_A2_c_367_n 0.0210879f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_95 VPB N_A2_c_363_n 0.0493915f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.212
cc_96 VPB N_A1_c_443_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_97 VPB N_A1_c_444_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_98 VPB N_A1_c_445_n 0.0166236f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_99 VPB N_A1_c_438_n 0.00825307f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_100 VPB N_A1_c_439_n 0.0360716f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_101 VPB N_A1_c_448_n 0.0214479f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A1_c_442_n 0.0166586f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.175
cc_103 VPB N_A_27_297#_c_513_n 0.00922995f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_104 VPB N_A_27_297#_c_514_n 0.0291185f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.015
cc_105 VPB N_A_27_297#_c_515_n 0.00184995f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.212
cc_106 VPB N_A_27_297#_c_516_n 0.00435684f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.212
cc_107 VPB N_Y_c_591_n 0.00336294f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.212
cc_108 VPB N_Y_c_594_n 0.0108306f $X=-0.19 $Y=1.305 $X2=1.67 $Y2=1.16
cc_109 VPB N_VPWR_c_720_n 4.04661e-19 $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.015
cc_110 VPB N_VPWR_c_721_n 4.04661e-19 $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_111 VPB N_VPWR_c_722_n 0.0114084f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.56
cc_112 VPB N_VPWR_c_723_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_113 VPB N_VPWR_c_724_n 0.0106521f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_725_n 0.0425695f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_726_n 0.113361f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.212
cc_116 VPB N_VPWR_c_727_n 0.00477947f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.212
cc_117 VPB N_VPWR_c_728_n 0.0206409f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.212
cc_118 VPB N_VPWR_c_729_n 0.00324069f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.212
cc_119 VPB N_VPWR_c_730_n 0.0563727f $X=-0.19 $Y=1.305 $X2=1.67 $Y2=1.16
cc_120 VPB N_VPWR_c_731_n 0.0127061f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.175
cc_121 VPB N_VPWR_c_732_n 0.0221761f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_733_n 0.00503156f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_734_n 0.00503156f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_719_n 0.0624475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_886_297#_c_868_n 0.00218721f $X=-0.19 $Y=1.305 $X2=1.435
+ $Y2=1.985
cc_126 VPB N_A_886_297#_c_869_n 0.0040066f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.015
cc_127 VPB N_A_886_297#_c_870_n 0.00218721f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.212
cc_128 VPB N_A_886_297#_c_871_n 0.00410007f $X=-0.19 $Y=1.305 $X2=1.435
+ $Y2=1.212
cc_129 VPB N_A_1352_297#_c_938_n 0.0132401f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_130 N_B2_M1038_g N_B1_M1005_g 0.0207012f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_131 N_B2_c_139_n N_B1_c_209_n 0.0324142f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_132 N_B2_c_135_n N_B1_c_208_n 0.0207012f $X=1.905 $Y=1.212 $X2=0 $Y2=0
cc_133 N_B2_c_134_n N_A_27_297#_c_514_n 0.0153565f $X=1.67 $Y=1.16 $X2=0 $Y2=0
cc_134 N_B2_c_135_n N_A_27_297#_c_514_n 0.00537148f $X=1.905 $Y=1.212 $X2=0
+ $Y2=0
cc_135 N_B2_c_136_n N_A_27_297#_c_519_n 0.0135433f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_136 N_B2_c_137_n N_A_27_297#_c_519_n 0.0122129f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_137 N_B2_c_138_n N_A_27_297#_c_521_n 0.0114822f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_138 N_B2_c_139_n N_A_27_297#_c_521_n 0.0130207f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_139 N_B2_c_139_n N_A_27_297#_c_523_n 0.0014328f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_140 N_B2_M1004_g N_Y_c_590_n 0.00607102f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_141 N_B2_M1026_g N_Y_c_590_n 0.0112895f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_142 N_B2_M1027_g N_Y_c_590_n 0.0112895f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_143 N_B2_M1038_g N_Y_c_590_n 0.0127785f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_144 N_B2_c_134_n N_Y_c_590_n 0.0970482f $X=1.67 $Y=1.16 $X2=0 $Y2=0
cc_145 N_B2_c_135_n N_Y_c_590_n 0.00994084f $X=1.905 $Y=1.212 $X2=0 $Y2=0
cc_146 N_B2_c_137_n N_Y_c_601_n 0.0113777f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_147 N_B2_c_138_n N_Y_c_601_n 0.00844992f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_148 N_B2_c_134_n N_Y_c_601_n 0.0285071f $X=1.67 $Y=1.16 $X2=0 $Y2=0
cc_149 N_B2_c_135_n N_Y_c_601_n 0.00623548f $X=1.905 $Y=1.212 $X2=0 $Y2=0
cc_150 N_B2_c_139_n N_Y_c_605_n 0.0120917f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_151 N_B2_c_139_n N_Y_c_591_n 0.00205706f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_152 N_B2_M1038_g N_Y_c_591_n 0.00958372f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_153 N_B2_c_134_n N_Y_c_591_n 0.0130702f $X=1.67 $Y=1.16 $X2=0 $Y2=0
cc_154 N_B2_c_136_n N_Y_c_609_n 0.0106394f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_155 N_B2_c_137_n N_Y_c_609_n 0.00689028f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_156 N_B2_c_138_n N_Y_c_609_n 5.03725e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_157 N_B2_c_134_n N_Y_c_609_n 0.0201192f $X=1.67 $Y=1.16 $X2=0 $Y2=0
cc_158 N_B2_c_135_n N_Y_c_609_n 0.00639631f $X=1.905 $Y=1.212 $X2=0 $Y2=0
cc_159 N_B2_c_138_n N_Y_c_614_n 0.002228f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_160 N_B2_c_139_n N_Y_c_614_n 0.00122806f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_161 N_B2_c_134_n N_Y_c_614_n 0.0201184f $X=1.67 $Y=1.16 $X2=0 $Y2=0
cc_162 N_B2_c_135_n N_Y_c_614_n 0.00639631f $X=1.905 $Y=1.212 $X2=0 $Y2=0
cc_163 N_B2_c_137_n Y 5.39594e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_164 N_B2_c_138_n Y 0.00814852f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_165 N_B2_c_139_n Y 0.00707207f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_166 N_B2_c_139_n N_VPWR_c_720_n 0.00123447f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_167 N_B2_c_136_n N_VPWR_c_730_n 0.00429453f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_168 N_B2_c_137_n N_VPWR_c_730_n 0.00429453f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_169 N_B2_c_138_n N_VPWR_c_730_n 0.00429453f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_170 N_B2_c_139_n N_VPWR_c_730_n 0.00429453f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_171 N_B2_c_136_n N_VPWR_c_719_n 0.00697643f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_172 N_B2_c_137_n N_VPWR_c_719_n 0.00606499f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_173 N_B2_c_138_n N_VPWR_c_719_n 0.00606499f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_174 N_B2_c_139_n N_VPWR_c_719_n 0.00616881f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_175 N_B2_M1004_g N_A_27_47#_c_1005_n 0.00497296f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_176 N_B2_c_134_n N_A_27_47#_c_1005_n 0.0190063f $X=1.67 $Y=1.16 $X2=0 $Y2=0
cc_177 N_B2_c_135_n N_A_27_47#_c_1005_n 0.00569691f $X=1.905 $Y=1.212 $X2=0
+ $Y2=0
cc_178 N_B2_M1004_g N_A_27_47#_c_1022_n 0.0100644f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_179 N_B2_M1026_g N_A_27_47#_c_1022_n 0.00915601f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_180 N_B2_M1027_g N_A_27_47#_c_1022_n 0.00915601f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_181 N_B2_M1038_g N_A_27_47#_c_1022_n 0.00915601f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_182 N_B2_c_134_n N_A_27_47#_c_1022_n 0.00349337f $X=1.67 $Y=1.16 $X2=0 $Y2=0
cc_183 N_B2_c_135_n N_A_27_47#_c_1022_n 0.00160484f $X=1.905 $Y=1.212 $X2=0
+ $Y2=0
cc_184 N_B2_M1004_g N_VGND_c_1182_n 0.00357877f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_185 N_B2_M1026_g N_VGND_c_1182_n 0.00357877f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_186 N_B2_M1027_g N_VGND_c_1182_n 0.00357877f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_187 N_B2_M1038_g N_VGND_c_1182_n 0.00357877f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_188 N_B2_M1004_g N_VGND_c_1195_n 0.00635588f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_189 N_B2_M1026_g N_VGND_c_1195_n 0.00548399f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_190 N_B2_M1027_g N_VGND_c_1195_n 0.00548399f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_191 N_B2_M1038_g N_VGND_c_1195_n 0.00542082f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_192 N_B1_M1039_g N_A3_M1012_g 0.0144883f $X=3.825 $Y=0.56 $X2=0 $Y2=0
cc_193 N_B1_c_207_n N_A3_c_275_n 8.49417e-19 $X=3.565 $Y=1.16 $X2=0 $Y2=0
cc_194 N_B1_c_208_n N_A3_c_275_n 0.0144883f $X=3.8 $Y=1.212 $X2=0 $Y2=0
cc_195 N_B1_c_207_n A3 0.0140536f $X=3.565 $Y=1.16 $X2=0 $Y2=0
cc_196 N_B1_c_208_n A3 2.32892e-19 $X=3.8 $Y=1.212 $X2=0 $Y2=0
cc_197 N_B1_c_209_n N_A_27_297#_c_521_n 0.00127104f $X=2.39 $Y=1.41 $X2=0 $Y2=0
cc_198 N_B1_c_209_n N_A_27_297#_c_525_n 0.0124008f $X=2.39 $Y=1.41 $X2=0 $Y2=0
cc_199 N_B1_c_210_n N_A_27_297#_c_525_n 0.011553f $X=2.86 $Y=1.41 $X2=0 $Y2=0
cc_200 N_B1_c_211_n N_A_27_297#_c_527_n 0.0110194f $X=3.33 $Y=1.41 $X2=0 $Y2=0
cc_201 N_B1_c_212_n N_A_27_297#_c_527_n 0.0115961f $X=3.8 $Y=1.41 $X2=0 $Y2=0
cc_202 N_B1_c_212_n N_A_27_297#_c_516_n 0.0049102f $X=3.8 $Y=1.41 $X2=0 $Y2=0
cc_203 N_B1_M1005_g N_Y_c_591_n 0.00936751f $X=2.365 $Y=0.56 $X2=0 $Y2=0
cc_204 N_B1_c_209_n N_Y_c_591_n 0.00204392f $X=2.39 $Y=1.41 $X2=0 $Y2=0
cc_205 N_B1_c_207_n N_Y_c_591_n 0.0158867f $X=3.565 $Y=1.16 $X2=0 $Y2=0
cc_206 N_B1_M1005_g N_Y_c_592_n 0.0123401f $X=2.365 $Y=0.56 $X2=0 $Y2=0
cc_207 N_B1_M1024_g N_Y_c_592_n 0.0112895f $X=2.835 $Y=0.56 $X2=0 $Y2=0
cc_208 N_B1_M1028_g N_Y_c_592_n 0.011285f $X=3.305 $Y=0.56 $X2=0 $Y2=0
cc_209 N_B1_M1039_g N_Y_c_592_n 2.03781e-19 $X=3.825 $Y=0.56 $X2=0 $Y2=0
cc_210 N_B1_c_207_n N_Y_c_592_n 0.0975986f $X=3.565 $Y=1.16 $X2=0 $Y2=0
cc_211 N_B1_c_208_n N_Y_c_592_n 0.0111243f $X=3.8 $Y=1.212 $X2=0 $Y2=0
cc_212 N_B1_c_209_n N_Y_c_594_n 0.0134413f $X=2.39 $Y=1.41 $X2=0 $Y2=0
cc_213 N_B1_c_210_n N_Y_c_594_n 0.0122688f $X=2.86 $Y=1.41 $X2=0 $Y2=0
cc_214 N_B1_c_211_n N_Y_c_594_n 0.0122688f $X=3.33 $Y=1.41 $X2=0 $Y2=0
cc_215 N_B1_c_212_n N_Y_c_594_n 0.0142686f $X=3.8 $Y=1.41 $X2=0 $Y2=0
cc_216 N_B1_c_207_n N_Y_c_594_n 0.0763672f $X=3.565 $Y=1.16 $X2=0 $Y2=0
cc_217 N_B1_c_208_n N_Y_c_594_n 0.0184849f $X=3.8 $Y=1.212 $X2=0 $Y2=0
cc_218 N_B1_c_209_n Y 9.18366e-19 $X=2.39 $Y=1.41 $X2=0 $Y2=0
cc_219 N_B1_c_209_n N_VPWR_c_720_n 0.0116502f $X=2.39 $Y=1.41 $X2=0 $Y2=0
cc_220 N_B1_c_210_n N_VPWR_c_720_n 0.00799817f $X=2.86 $Y=1.41 $X2=0 $Y2=0
cc_221 N_B1_c_211_n N_VPWR_c_720_n 5.90726e-19 $X=3.33 $Y=1.41 $X2=0 $Y2=0
cc_222 N_B1_c_210_n N_VPWR_c_721_n 6.47527e-19 $X=2.86 $Y=1.41 $X2=0 $Y2=0
cc_223 N_B1_c_211_n N_VPWR_c_721_n 0.0108702f $X=3.33 $Y=1.41 $X2=0 $Y2=0
cc_224 N_B1_c_212_n N_VPWR_c_721_n 0.00935472f $X=3.8 $Y=1.41 $X2=0 $Y2=0
cc_225 N_B1_c_212_n N_VPWR_c_726_n 0.00464801f $X=3.8 $Y=1.41 $X2=0 $Y2=0
cc_226 N_B1_c_209_n N_VPWR_c_730_n 0.00319306f $X=2.39 $Y=1.41 $X2=0 $Y2=0
cc_227 N_B1_c_210_n N_VPWR_c_731_n 0.00464801f $X=2.86 $Y=1.41 $X2=0 $Y2=0
cc_228 N_B1_c_211_n N_VPWR_c_731_n 0.00319306f $X=3.33 $Y=1.41 $X2=0 $Y2=0
cc_229 N_B1_c_209_n N_VPWR_c_719_n 0.00396435f $X=2.39 $Y=1.41 $X2=0 $Y2=0
cc_230 N_B1_c_210_n N_VPWR_c_719_n 0.00539343f $X=2.86 $Y=1.41 $X2=0 $Y2=0
cc_231 N_B1_c_211_n N_VPWR_c_719_n 0.00390143f $X=3.33 $Y=1.41 $X2=0 $Y2=0
cc_232 N_B1_c_212_n N_VPWR_c_719_n 0.0067251f $X=3.8 $Y=1.41 $X2=0 $Y2=0
cc_233 N_B1_M1005_g N_A_27_47#_c_1022_n 0.00915601f $X=2.365 $Y=0.56 $X2=0 $Y2=0
cc_234 N_B1_M1024_g N_A_27_47#_c_1022_n 0.00915601f $X=2.835 $Y=0.56 $X2=0 $Y2=0
cc_235 N_B1_M1028_g N_A_27_47#_c_1022_n 0.00947663f $X=3.305 $Y=0.56 $X2=0 $Y2=0
cc_236 N_B1_M1039_g N_A_27_47#_c_1022_n 0.0114382f $X=3.825 $Y=0.56 $X2=0 $Y2=0
cc_237 N_B1_c_207_n N_A_27_47#_c_1022_n 0.00449518f $X=3.565 $Y=1.16 $X2=0 $Y2=0
cc_238 N_B1_M1005_g N_VGND_c_1182_n 0.00357877f $X=2.365 $Y=0.56 $X2=0 $Y2=0
cc_239 N_B1_M1024_g N_VGND_c_1182_n 0.00357877f $X=2.835 $Y=0.56 $X2=0 $Y2=0
cc_240 N_B1_M1028_g N_VGND_c_1182_n 0.00357877f $X=3.305 $Y=0.56 $X2=0 $Y2=0
cc_241 N_B1_M1039_g N_VGND_c_1182_n 0.00357877f $X=3.825 $Y=0.56 $X2=0 $Y2=0
cc_242 N_B1_M1005_g N_VGND_c_1195_n 0.00542082f $X=2.365 $Y=0.56 $X2=0 $Y2=0
cc_243 N_B1_M1024_g N_VGND_c_1195_n 0.00548399f $X=2.835 $Y=0.56 $X2=0 $Y2=0
cc_244 N_B1_M1028_g N_VGND_c_1195_n 0.00560377f $X=3.305 $Y=0.56 $X2=0 $Y2=0
cc_245 N_B1_M1039_g N_VGND_c_1195_n 0.005504f $X=3.825 $Y=0.56 $X2=0 $Y2=0
cc_246 N_A3_M1031_g N_A2_M1006_g 0.00469042f $X=5.815 $Y=0.56 $X2=0 $Y2=0
cc_247 N_A3_c_282_n N_A2_c_364_n 0.0229948f $X=6.2 $Y=1.41 $X2=0 $Y2=0
cc_248 A3 N_A2_c_362_n 0.00733776f $X=5.675 $Y=1.105 $X2=0 $Y2=0
cc_249 N_A3_c_278_n N_A2_c_362_n 0.00234519f $X=5.815 $Y=1.212 $X2=0 $Y2=0
cc_250 N_A3_c_278_n N_A2_c_363_n 0.0214954f $X=5.815 $Y=1.212 $X2=0 $Y2=0
cc_251 N_A3_c_279_n N_Y_c_594_n 0.0133775f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_252 N_A3_c_275_n N_Y_c_594_n 0.0128941f $X=4.32 $Y=1.16 $X2=0 $Y2=0
cc_253 A3 N_Y_c_594_n 0.0383986f $X=5.675 $Y=1.105 $X2=0 $Y2=0
cc_254 N_A3_c_280_n N_Y_c_640_n 0.0113777f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_255 N_A3_c_281_n N_Y_c_640_n 0.00844992f $X=5.73 $Y=1.41 $X2=0 $Y2=0
cc_256 A3 N_Y_c_640_n 0.0285071f $X=5.675 $Y=1.105 $X2=0 $Y2=0
cc_257 N_A3_c_278_n N_Y_c_640_n 0.00565948f $X=5.815 $Y=1.212 $X2=0 $Y2=0
cc_258 N_A3_c_279_n N_Y_c_644_n 0.0112633f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A3_c_280_n N_Y_c_644_n 0.00689028f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A3_c_281_n N_Y_c_644_n 5.04446e-19 $X=5.73 $Y=1.41 $X2=0 $Y2=0
cc_261 A3 N_Y_c_644_n 0.0170249f $X=5.675 $Y=1.105 $X2=0 $Y2=0
cc_262 N_A3_c_278_n N_Y_c_644_n 0.00644066f $X=5.815 $Y=1.212 $X2=0 $Y2=0
cc_263 N_A3_c_280_n N_Y_c_649_n 5.398e-19 $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A3_c_281_n N_Y_c_649_n 0.0103765f $X=5.73 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A3_c_282_n N_Y_c_649_n 0.00986171f $X=6.2 $Y=1.41 $X2=0 $Y2=0
cc_266 A3 N_Y_c_649_n 0.0125766f $X=5.675 $Y=1.105 $X2=0 $Y2=0
cc_267 N_A3_c_278_n N_Y_c_649_n 0.00643186f $X=5.815 $Y=1.212 $X2=0 $Y2=0
cc_268 N_A3_c_279_n N_VPWR_c_726_n 0.00429453f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A3_c_280_n N_VPWR_c_726_n 0.00429453f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_270 N_A3_c_281_n N_VPWR_c_726_n 0.00429453f $X=5.73 $Y=1.41 $X2=0 $Y2=0
cc_271 N_A3_c_282_n N_VPWR_c_726_n 0.00429453f $X=6.2 $Y=1.41 $X2=0 $Y2=0
cc_272 N_A3_c_279_n N_VPWR_c_719_n 0.00734734f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_273 N_A3_c_280_n N_VPWR_c_719_n 0.00606499f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_274 N_A3_c_281_n N_VPWR_c_719_n 0.00606499f $X=5.73 $Y=1.41 $X2=0 $Y2=0
cc_275 N_A3_c_282_n N_VPWR_c_719_n 0.00609021f $X=6.2 $Y=1.41 $X2=0 $Y2=0
cc_276 N_A3_c_279_n N_A_886_297#_c_872_n 0.0122129f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_277 N_A3_c_280_n N_A_886_297#_c_872_n 0.0122129f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_278 N_A3_c_281_n N_A_886_297#_c_874_n 0.0115355f $X=5.73 $Y=1.41 $X2=0 $Y2=0
cc_279 N_A3_c_282_n N_A_886_297#_c_874_n 0.0151209f $X=6.2 $Y=1.41 $X2=0 $Y2=0
cc_280 N_A3_c_282_n N_A_1352_297#_c_939_n 0.00107778f $X=6.2 $Y=1.41 $X2=0 $Y2=0
cc_281 N_A3_M1012_g N_A_27_47#_c_1033_n 0.00271016f $X=4.245 $Y=0.56 $X2=0 $Y2=0
cc_282 N_A3_M1012_g N_A_27_47#_c_1006_n 0.00547261f $X=4.245 $Y=0.56 $X2=0 $Y2=0
cc_283 N_A3_M1013_g N_A_27_47#_c_1006_n 5.3593e-19 $X=4.715 $Y=0.56 $X2=0 $Y2=0
cc_284 A3 N_A_27_47#_c_1006_n 0.00230247f $X=5.675 $Y=1.105 $X2=0 $Y2=0
cc_285 N_A3_M1012_g N_A_27_47#_c_1007_n 0.00879805f $X=4.245 $Y=0.56 $X2=0 $Y2=0
cc_286 N_A3_M1013_g N_A_27_47#_c_1007_n 0.00874287f $X=4.715 $Y=0.56 $X2=0 $Y2=0
cc_287 A3 N_A_27_47#_c_1007_n 0.0395004f $X=5.675 $Y=1.105 $X2=0 $Y2=0
cc_288 N_A3_c_277_n N_A_27_47#_c_1007_n 0.00328139f $X=4.64 $Y=1.16 $X2=0 $Y2=0
cc_289 N_A3_M1012_g N_A_27_47#_c_1041_n 5.82865e-19 $X=4.245 $Y=0.56 $X2=0 $Y2=0
cc_290 N_A3_M1013_g N_A_27_47#_c_1041_n 0.00678142f $X=4.715 $Y=0.56 $X2=0 $Y2=0
cc_291 N_A3_M1017_g N_A_27_47#_c_1041_n 0.00785018f $X=5.185 $Y=0.56 $X2=0 $Y2=0
cc_292 N_A3_M1031_g N_A_27_47#_c_1041_n 9.07158e-19 $X=5.815 $Y=0.56 $X2=0 $Y2=0
cc_293 N_A3_M1013_g N_A_27_47#_c_1012_n 0.00113905f $X=4.715 $Y=0.56 $X2=0 $Y2=0
cc_294 N_A3_M1017_g N_A_27_47#_c_1012_n 0.00113905f $X=5.185 $Y=0.56 $X2=0 $Y2=0
cc_295 A3 N_A_27_47#_c_1012_n 0.0306019f $X=5.675 $Y=1.105 $X2=0 $Y2=0
cc_296 N_A3_c_278_n N_A_27_47#_c_1012_n 0.00342373f $X=5.815 $Y=1.212 $X2=0
+ $Y2=0
cc_297 N_A3_M1017_g N_A_27_47#_c_1013_n 0.00951792f $X=5.185 $Y=0.56 $X2=0 $Y2=0
cc_298 N_A3_M1031_g N_A_27_47#_c_1013_n 0.0115541f $X=5.815 $Y=0.56 $X2=0 $Y2=0
cc_299 A3 N_A_27_47#_c_1013_n 0.0603122f $X=5.675 $Y=1.105 $X2=0 $Y2=0
cc_300 N_A3_c_278_n N_A_27_47#_c_1013_n 0.0226407f $X=5.815 $Y=1.212 $X2=0 $Y2=0
cc_301 N_A3_M1012_g N_VGND_c_1176_n 0.00375751f $X=4.245 $Y=0.56 $X2=0 $Y2=0
cc_302 N_A3_M1013_g N_VGND_c_1176_n 0.00276126f $X=4.715 $Y=0.56 $X2=0 $Y2=0
cc_303 N_A3_M1017_g N_VGND_c_1177_n 0.00620702f $X=5.185 $Y=0.56 $X2=0 $Y2=0
cc_304 N_A3_M1031_g N_VGND_c_1177_n 0.00524095f $X=5.815 $Y=0.56 $X2=0 $Y2=0
cc_305 N_A3_M1012_g N_VGND_c_1182_n 0.00422898f $X=4.245 $Y=0.56 $X2=0 $Y2=0
cc_306 N_A3_M1013_g N_VGND_c_1184_n 0.00424416f $X=4.715 $Y=0.56 $X2=0 $Y2=0
cc_307 N_A3_M1017_g N_VGND_c_1184_n 0.00424416f $X=5.185 $Y=0.56 $X2=0 $Y2=0
cc_308 N_A3_M1031_g N_VGND_c_1186_n 0.00439206f $X=5.815 $Y=0.56 $X2=0 $Y2=0
cc_309 N_A3_M1012_g N_VGND_c_1195_n 0.00602209f $X=4.245 $Y=0.56 $X2=0 $Y2=0
cc_310 N_A3_M1013_g N_VGND_c_1195_n 0.00599001f $X=4.715 $Y=0.56 $X2=0 $Y2=0
cc_311 N_A3_M1017_g N_VGND_c_1195_n 0.00650836f $X=5.185 $Y=0.56 $X2=0 $Y2=0
cc_312 N_A3_M1031_g N_VGND_c_1195_n 0.00717549f $X=5.815 $Y=0.56 $X2=0 $Y2=0
cc_313 N_A2_c_364_n N_Y_c_649_n 9.91702e-19 $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_314 N_A2_c_367_n N_VPWR_c_722_n 0.00228307f $X=8.08 $Y=1.41 $X2=0 $Y2=0
cc_315 N_A2_c_364_n N_VPWR_c_726_n 0.00429453f $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_316 N_A2_c_365_n N_VPWR_c_726_n 0.00429453f $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_317 N_A2_c_366_n N_VPWR_c_726_n 0.00429453f $X=7.61 $Y=1.41 $X2=0 $Y2=0
cc_318 N_A2_c_367_n N_VPWR_c_726_n 0.00429453f $X=8.08 $Y=1.41 $X2=0 $Y2=0
cc_319 N_A2_c_364_n N_VPWR_c_719_n 0.00609021f $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_320 N_A2_c_365_n N_VPWR_c_719_n 0.00606499f $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_321 N_A2_c_366_n N_VPWR_c_719_n 0.00606499f $X=7.61 $Y=1.41 $X2=0 $Y2=0
cc_322 N_A2_c_367_n N_VPWR_c_719_n 0.00734734f $X=8.08 $Y=1.41 $X2=0 $Y2=0
cc_323 N_A2_c_364_n N_A_886_297#_c_876_n 0.0135433f $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_324 N_A2_c_365_n N_A_886_297#_c_876_n 0.0122129f $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_325 N_A2_c_366_n N_A_886_297#_c_878_n 0.0115355f $X=7.61 $Y=1.41 $X2=0 $Y2=0
cc_326 N_A2_c_367_n N_A_886_297#_c_878_n 0.0122129f $X=8.08 $Y=1.41 $X2=0 $Y2=0
cc_327 N_A2_c_365_n N_A_1352_297#_c_940_n 0.0113777f $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_328 N_A2_c_366_n N_A_1352_297#_c_940_n 0.00844992f $X=7.61 $Y=1.41 $X2=0
+ $Y2=0
cc_329 N_A2_c_362_n N_A_1352_297#_c_940_n 0.0285071f $X=7.845 $Y=1.16 $X2=0
+ $Y2=0
cc_330 N_A2_c_363_n N_A_1352_297#_c_940_n 0.00623548f $X=8.08 $Y=1.212 $X2=0
+ $Y2=0
cc_331 N_A2_c_367_n N_A_1352_297#_c_938_n 0.0151858f $X=8.08 $Y=1.41 $X2=0 $Y2=0
cc_332 N_A2_c_364_n N_A_1352_297#_c_939_n 0.0129876f $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_333 N_A2_c_365_n N_A_1352_297#_c_939_n 0.00689028f $X=7.14 $Y=1.41 $X2=0
+ $Y2=0
cc_334 N_A2_c_366_n N_A_1352_297#_c_939_n 5.03725e-19 $X=7.61 $Y=1.41 $X2=0
+ $Y2=0
cc_335 N_A2_c_362_n N_A_1352_297#_c_939_n 0.0201192f $X=7.845 $Y=1.16 $X2=0
+ $Y2=0
cc_336 N_A2_c_363_n N_A_1352_297#_c_939_n 0.00639631f $X=8.08 $Y=1.212 $X2=0
+ $Y2=0
cc_337 N_A2_c_365_n N_A_1352_297#_c_950_n 5.398e-19 $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_338 N_A2_c_366_n N_A_1352_297#_c_950_n 0.0103765f $X=7.61 $Y=1.41 $X2=0 $Y2=0
cc_339 N_A2_c_367_n N_A_1352_297#_c_950_n 0.0113799f $X=8.08 $Y=1.41 $X2=0 $Y2=0
cc_340 N_A2_c_362_n N_A_1352_297#_c_950_n 0.0201192f $X=7.845 $Y=1.16 $X2=0
+ $Y2=0
cc_341 N_A2_c_363_n N_A_1352_297#_c_950_n 0.00617453f $X=8.08 $Y=1.212 $X2=0
+ $Y2=0
cc_342 N_A2_M1006_g N_A_27_47#_c_1008_n 0.00990019f $X=6.645 $Y=0.56 $X2=0 $Y2=0
cc_343 N_A2_M1009_g N_A_27_47#_c_1008_n 0.00879805f $X=7.115 $Y=0.56 $X2=0 $Y2=0
cc_344 N_A2_c_363_n N_A_27_47#_c_1008_n 0.00328139f $X=8.08 $Y=1.212 $X2=0 $Y2=0
cc_345 N_A2_M1006_g N_A_27_47#_c_1056_n 5.86828e-19 $X=6.645 $Y=0.56 $X2=0 $Y2=0
cc_346 N_A2_M1009_g N_A_27_47#_c_1056_n 0.00683102f $X=7.115 $Y=0.56 $X2=0 $Y2=0
cc_347 N_A2_M1019_g N_A_27_47#_c_1056_n 0.00718011f $X=7.585 $Y=0.56 $X2=0 $Y2=0
cc_348 N_A2_M1033_g N_A_27_47#_c_1056_n 5.92369e-19 $X=8.105 $Y=0.56 $X2=0 $Y2=0
cc_349 N_A2_M1006_g N_A_27_47#_c_1014_n 0.00718522f $X=6.645 $Y=0.56 $X2=0 $Y2=0
cc_350 N_A2_M1009_g N_A_27_47#_c_1014_n 5.88234e-19 $X=7.115 $Y=0.56 $X2=0 $Y2=0
cc_351 N_A2_c_362_n N_A_27_47#_c_1014_n 0.0459421f $X=7.845 $Y=1.16 $X2=0 $Y2=0
cc_352 N_A2_M1009_g N_A_27_47#_c_1015_n 0.00113905f $X=7.115 $Y=0.56 $X2=0 $Y2=0
cc_353 N_A2_M1019_g N_A_27_47#_c_1015_n 0.00113905f $X=7.585 $Y=0.56 $X2=0 $Y2=0
cc_354 N_A2_c_362_n N_A_27_47#_c_1015_n 0.0306019f $X=7.845 $Y=1.16 $X2=0 $Y2=0
cc_355 N_A2_c_363_n N_A_27_47#_c_1015_n 0.00340841f $X=8.08 $Y=1.212 $X2=0 $Y2=0
cc_356 N_A2_M1019_g N_A_27_47#_c_1016_n 0.00905701f $X=7.585 $Y=0.56 $X2=0 $Y2=0
cc_357 N_A2_M1033_g N_A_27_47#_c_1016_n 0.00722392f $X=8.105 $Y=0.56 $X2=0 $Y2=0
cc_358 N_A2_c_362_n N_A_27_47#_c_1016_n 0.0335381f $X=7.845 $Y=1.16 $X2=0 $Y2=0
cc_359 N_A2_c_363_n N_A_27_47#_c_1016_n 0.00445332f $X=8.08 $Y=1.212 $X2=0 $Y2=0
cc_360 N_A2_M1019_g N_A_27_47#_c_1017_n 6.31595e-19 $X=7.585 $Y=0.56 $X2=0 $Y2=0
cc_361 N_A2_M1033_g N_A_27_47#_c_1017_n 0.0128668f $X=8.105 $Y=0.56 $X2=0 $Y2=0
cc_362 N_A2_M1006_g N_VGND_c_1178_n 0.00384711f $X=6.645 $Y=0.56 $X2=0 $Y2=0
cc_363 N_A2_M1009_g N_VGND_c_1178_n 0.00276126f $X=7.115 $Y=0.56 $X2=0 $Y2=0
cc_364 N_A2_M1019_g N_VGND_c_1179_n 0.00382269f $X=7.585 $Y=0.56 $X2=0 $Y2=0
cc_365 N_A2_M1033_g N_VGND_c_1179_n 0.00364096f $X=8.105 $Y=0.56 $X2=0 $Y2=0
cc_366 N_A2_M1006_g N_VGND_c_1186_n 0.00433784f $X=6.645 $Y=0.56 $X2=0 $Y2=0
cc_367 N_A2_M1009_g N_VGND_c_1188_n 0.00424416f $X=7.115 $Y=0.56 $X2=0 $Y2=0
cc_368 N_A2_M1019_g N_VGND_c_1188_n 0.00424416f $X=7.585 $Y=0.56 $X2=0 $Y2=0
cc_369 N_A2_M1033_g N_VGND_c_1190_n 0.00395831f $X=8.105 $Y=0.56 $X2=0 $Y2=0
cc_370 N_A2_M1006_g N_VGND_c_1195_n 0.00685134f $X=6.645 $Y=0.56 $X2=0 $Y2=0
cc_371 N_A2_M1009_g N_VGND_c_1195_n 0.00599001f $X=7.115 $Y=0.56 $X2=0 $Y2=0
cc_372 N_A2_M1019_g N_VGND_c_1195_n 0.00622812f $X=7.585 $Y=0.56 $X2=0 $Y2=0
cc_373 N_A2_M1033_g N_VGND_c_1195_n 0.00714991f $X=8.105 $Y=0.56 $X2=0 $Y2=0
cc_374 N_A1_c_443_n N_VPWR_c_722_n 0.00673063f $X=9.07 $Y=1.41 $X2=0 $Y2=0
cc_375 N_A1_c_444_n N_VPWR_c_723_n 0.0052072f $X=9.54 $Y=1.41 $X2=0 $Y2=0
cc_376 N_A1_c_445_n N_VPWR_c_723_n 0.004751f $X=10.01 $Y=1.41 $X2=0 $Y2=0
cc_377 N_A1_c_448_n N_VPWR_c_725_n 0.00917994f $X=10.525 $Y=1.41 $X2=0 $Y2=0
cc_378 A1 N_VPWR_c_725_n 0.0166705f $X=10.72 $Y=1.105 $X2=0 $Y2=0
cc_379 N_A1_c_442_n N_VPWR_c_725_n 0.00353507f $X=10.525 $Y=1.212 $X2=0 $Y2=0
cc_380 N_A1_c_443_n N_VPWR_c_728_n 0.00597712f $X=9.07 $Y=1.41 $X2=0 $Y2=0
cc_381 N_A1_c_444_n N_VPWR_c_728_n 0.00673617f $X=9.54 $Y=1.41 $X2=0 $Y2=0
cc_382 N_A1_c_445_n N_VPWR_c_732_n 0.00597712f $X=10.01 $Y=1.41 $X2=0 $Y2=0
cc_383 N_A1_c_448_n N_VPWR_c_732_n 0.00702461f $X=10.525 $Y=1.41 $X2=0 $Y2=0
cc_384 N_A1_c_443_n N_VPWR_c_719_n 0.0112769f $X=9.07 $Y=1.41 $X2=0 $Y2=0
cc_385 N_A1_c_444_n N_VPWR_c_719_n 0.0118438f $X=9.54 $Y=1.41 $X2=0 $Y2=0
cc_386 N_A1_c_445_n N_VPWR_c_719_n 0.0101051f $X=10.01 $Y=1.41 $X2=0 $Y2=0
cc_387 N_A1_c_448_n N_VPWR_c_719_n 0.0135496f $X=10.525 $Y=1.41 $X2=0 $Y2=0
cc_388 N_A1_c_443_n N_A_1352_297#_c_938_n 0.0135615f $X=9.07 $Y=1.41 $X2=0 $Y2=0
cc_389 N_A1_c_443_n N_A_1352_297#_c_956_n 0.0178402f $X=9.07 $Y=1.41 $X2=0 $Y2=0
cc_390 N_A1_c_444_n N_A_1352_297#_c_956_n 0.0106251f $X=9.54 $Y=1.41 $X2=0 $Y2=0
cc_391 N_A1_c_445_n N_A_1352_297#_c_956_n 6.24674e-19 $X=10.01 $Y=1.41 $X2=0
+ $Y2=0
cc_392 N_A1_c_444_n N_A_1352_297#_c_959_n 0.0141085f $X=9.54 $Y=1.41 $X2=0 $Y2=0
cc_393 N_A1_c_445_n N_A_1352_297#_c_959_n 0.010322f $X=10.01 $Y=1.41 $X2=0 $Y2=0
cc_394 N_A1_c_439_n N_A_1352_297#_c_959_n 0.00623548f $X=10.11 $Y=1.16 $X2=0
+ $Y2=0
cc_395 A1 N_A_1352_297#_c_959_n 0.0285071f $X=10.72 $Y=1.105 $X2=0 $Y2=0
cc_396 N_A1_c_445_n N_A_1352_297#_c_963_n 0.00225158f $X=10.01 $Y=1.41 $X2=0
+ $Y2=0
cc_397 N_A1_c_438_n N_A_1352_297#_c_963_n 0.00707949f $X=10.425 $Y=1.16 $X2=0
+ $Y2=0
cc_398 A1 N_A_1352_297#_c_963_n 0.0213064f $X=10.72 $Y=1.105 $X2=0 $Y2=0
cc_399 N_A1_c_444_n N_A_1352_297#_c_966_n 6.48386e-19 $X=9.54 $Y=1.41 $X2=0
+ $Y2=0
cc_400 N_A1_c_445_n N_A_1352_297#_c_966_n 0.0130707f $X=10.01 $Y=1.41 $X2=0
+ $Y2=0
cc_401 N_A1_c_443_n N_A_1352_297#_c_968_n 0.00225158f $X=9.07 $Y=1.41 $X2=0
+ $Y2=0
cc_402 N_A1_c_444_n N_A_1352_297#_c_968_n 6.2e-19 $X=9.54 $Y=1.41 $X2=0 $Y2=0
cc_403 N_A1_c_439_n N_A_1352_297#_c_968_n 0.00642534f $X=10.11 $Y=1.16 $X2=0
+ $Y2=0
cc_404 A1 N_A_1352_297#_c_968_n 0.020318f $X=10.72 $Y=1.105 $X2=0 $Y2=0
cc_405 N_A1_M1015_g N_A_27_47#_c_1009_n 0.0161317f $X=9.045 $Y=0.56 $X2=0 $Y2=0
cc_406 N_A1_M1020_g N_A_27_47#_c_1009_n 0.00879805f $X=9.515 $Y=0.56 $X2=0 $Y2=0
cc_407 N_A1_c_439_n N_A_27_47#_c_1009_n 0.00328139f $X=10.11 $Y=1.16 $X2=0 $Y2=0
cc_408 A1 N_A_27_47#_c_1009_n 0.0334263f $X=10.72 $Y=1.105 $X2=0 $Y2=0
cc_409 N_A1_M1015_g N_A_27_47#_c_1077_n 9.20069e-19 $X=9.045 $Y=0.56 $X2=0 $Y2=0
cc_410 N_A1_M1020_g N_A_27_47#_c_1077_n 0.00697449f $X=9.515 $Y=0.56 $X2=0 $Y2=0
cc_411 N_A1_M1032_g N_A_27_47#_c_1077_n 0.00732269f $X=9.985 $Y=0.56 $X2=0 $Y2=0
cc_412 N_A1_M1035_g N_A_27_47#_c_1077_n 6.02058e-19 $X=10.5 $Y=0.56 $X2=0 $Y2=0
cc_413 N_A1_M1032_g N_A_27_47#_c_1010_n 0.00903265f $X=9.985 $Y=0.56 $X2=0 $Y2=0
cc_414 N_A1_c_438_n N_A_27_47#_c_1010_n 0.00433613f $X=10.425 $Y=1.16 $X2=0
+ $Y2=0
cc_415 N_A1_M1035_g N_A_27_47#_c_1010_n 0.0103146f $X=10.5 $Y=0.56 $X2=0 $Y2=0
cc_416 A1 N_A_27_47#_c_1010_n 0.073856f $X=10.72 $Y=1.105 $X2=0 $Y2=0
cc_417 N_A1_c_442_n N_A_27_47#_c_1010_n 0.006417f $X=10.525 $Y=1.212 $X2=0 $Y2=0
cc_418 N_A1_M1032_g N_A_27_47#_c_1011_n 6.5576e-19 $X=9.985 $Y=0.56 $X2=0 $Y2=0
cc_419 N_A1_M1035_g N_A_27_47#_c_1011_n 0.00698027f $X=10.5 $Y=0.56 $X2=0 $Y2=0
cc_420 N_A1_M1015_g N_A_27_47#_c_1017_n 0.0152198f $X=9.045 $Y=0.56 $X2=0 $Y2=0
cc_421 N_A1_M1020_g N_A_27_47#_c_1018_n 0.00113905f $X=9.515 $Y=0.56 $X2=0 $Y2=0
cc_422 N_A1_M1032_g N_A_27_47#_c_1018_n 0.00113905f $X=9.985 $Y=0.56 $X2=0 $Y2=0
cc_423 N_A1_c_439_n N_A_27_47#_c_1018_n 0.00340841f $X=10.11 $Y=1.16 $X2=0 $Y2=0
cc_424 A1 N_A_27_47#_c_1018_n 0.0306019f $X=10.72 $Y=1.105 $X2=0 $Y2=0
cc_425 N_A1_M1015_g N_VGND_c_1180_n 0.00433891f $X=9.045 $Y=0.56 $X2=0 $Y2=0
cc_426 N_A1_M1020_g N_VGND_c_1180_n 0.00276126f $X=9.515 $Y=0.56 $X2=0 $Y2=0
cc_427 N_A1_M1032_g N_VGND_c_1181_n 0.00544034f $X=9.985 $Y=0.56 $X2=0 $Y2=0
cc_428 N_A1_M1035_g N_VGND_c_1181_n 0.00289099f $X=10.5 $Y=0.56 $X2=0 $Y2=0
cc_429 N_A1_M1015_g N_VGND_c_1190_n 0.00439206f $X=9.045 $Y=0.56 $X2=0 $Y2=0
cc_430 N_A1_M1020_g N_VGND_c_1192_n 0.00424416f $X=9.515 $Y=0.56 $X2=0 $Y2=0
cc_431 N_A1_M1032_g N_VGND_c_1192_n 0.00424416f $X=9.985 $Y=0.56 $X2=0 $Y2=0
cc_432 N_A1_M1035_g N_VGND_c_1194_n 0.00424416f $X=10.5 $Y=0.56 $X2=0 $Y2=0
cc_433 N_A1_M1015_g N_VGND_c_1195_n 0.00758272f $X=9.045 $Y=0.56 $X2=0 $Y2=0
cc_434 N_A1_M1020_g N_VGND_c_1195_n 0.00599001f $X=9.515 $Y=0.56 $X2=0 $Y2=0
cc_435 N_A1_M1032_g N_VGND_c_1195_n 0.00627058f $X=9.985 $Y=0.56 $X2=0 $Y2=0
cc_436 N_A1_M1035_g N_VGND_c_1195_n 0.00698226f $X=10.5 $Y=0.56 $X2=0 $Y2=0
cc_437 N_A_27_297#_c_519_n N_Y_M1002_s 0.00354696f $X=1.115 $Y=2.36 $X2=0 $Y2=0
cc_438 N_A_27_297#_c_521_n N_Y_M1025_s 0.00354696f $X=2.07 $Y=2.36 $X2=0 $Y2=0
cc_439 N_A_27_297#_M1016_d N_Y_c_601_n 0.00342641f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_440 N_A_27_297#_c_519_n N_Y_c_601_n 0.0039635f $X=1.115 $Y=2.36 $X2=0 $Y2=0
cc_441 N_A_27_297#_c_534_p N_Y_c_601_n 0.0135833f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_442 N_A_27_297#_c_521_n N_Y_c_601_n 0.00273065f $X=2.07 $Y=2.36 $X2=0 $Y2=0
cc_443 N_A_27_297#_c_521_n N_Y_c_605_n 0.00359503f $X=2.07 $Y=2.36 $X2=0 $Y2=0
cc_444 N_A_27_297#_M1007_d N_Y_c_594_n 0.00344767f $X=2.95 $Y=1.485 $X2=0 $Y2=0
cc_445 N_A_27_297#_M1034_d N_Y_c_594_n 0.00720894f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_446 N_A_27_297#_c_525_n N_Y_c_594_n 0.0373684f $X=3.01 $Y=1.92 $X2=0 $Y2=0
cc_447 N_A_27_297#_c_523_n N_Y_c_594_n 3.67789e-19 $X=2.24 $Y=1.92 $X2=0 $Y2=0
cc_448 N_A_27_297#_c_527_n N_Y_c_594_n 0.0373345f $X=3.95 $Y=1.92 $X2=0 $Y2=0
cc_449 N_A_27_297#_c_515_n N_Y_c_594_n 0.0203373f $X=4.075 $Y=2.005 $X2=0 $Y2=0
cc_450 N_A_27_297#_c_543_p N_Y_c_594_n 0.0136738f $X=3.095 $Y=1.92 $X2=0 $Y2=0
cc_451 N_A_27_297#_c_514_n N_Y_c_609_n 0.0460215f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_452 N_A_27_297#_c_519_n N_Y_c_609_n 0.0198628f $X=1.115 $Y=2.36 $X2=0 $Y2=0
cc_453 N_A_27_297#_c_534_p N_Y_c_609_n 0.0153021f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_454 N_A_27_297#_M1036_d N_Y_c_672_n 0.00210464f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_455 N_A_27_297#_c_521_n N_Y_c_672_n 4.54881e-19 $X=2.07 $Y=2.36 $X2=0 $Y2=0
cc_456 N_A_27_297#_c_523_n N_Y_c_672_n 0.0147478f $X=2.24 $Y=1.92 $X2=0 $Y2=0
cc_457 N_A_27_297#_c_534_p Y 0.0187207f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_458 N_A_27_297#_c_521_n Y 0.0209463f $X=2.07 $Y=2.36 $X2=0 $Y2=0
cc_459 N_A_27_297#_c_552_p Y 0.00488151f $X=2.155 $Y=2.17 $X2=0 $Y2=0
cc_460 N_A_27_297#_c_523_n Y 0.011653f $X=2.24 $Y=1.92 $X2=0 $Y2=0
cc_461 N_A_27_297#_c_525_n N_VPWR_M1000_s 0.00350529f $X=3.01 $Y=1.92 $X2=-0.19
+ $Y2=1.305
cc_462 N_A_27_297#_c_527_n N_VPWR_M1022_s 0.00350529f $X=3.95 $Y=1.92 $X2=0
+ $Y2=0
cc_463 N_A_27_297#_c_521_n N_VPWR_c_720_n 0.0175144f $X=2.07 $Y=2.36 $X2=0 $Y2=0
cc_464 N_A_27_297#_c_552_p N_VPWR_c_720_n 0.00593609f $X=2.155 $Y=2.17 $X2=0
+ $Y2=0
cc_465 N_A_27_297#_c_525_n N_VPWR_c_720_n 0.0200892f $X=3.01 $Y=1.92 $X2=0 $Y2=0
cc_466 N_A_27_297#_c_559_p N_VPWR_c_720_n 0.0153021f $X=3.095 $Y=2.26 $X2=0
+ $Y2=0
cc_467 N_A_27_297#_c_559_p N_VPWR_c_721_n 0.0186638f $X=3.095 $Y=2.26 $X2=0
+ $Y2=0
cc_468 N_A_27_297#_c_527_n N_VPWR_c_721_n 0.0200892f $X=3.95 $Y=1.92 $X2=0 $Y2=0
cc_469 N_A_27_297#_c_516_n N_VPWR_c_721_n 0.0182679f $X=4.035 $Y=2.26 $X2=0
+ $Y2=0
cc_470 N_A_27_297#_c_527_n N_VPWR_c_726_n 0.00265246f $X=3.95 $Y=1.92 $X2=0
+ $Y2=0
cc_471 N_A_27_297#_c_516_n N_VPWR_c_726_n 0.017395f $X=4.035 $Y=2.26 $X2=0 $Y2=0
cc_472 N_A_27_297#_c_513_n N_VPWR_c_730_n 0.0179936f $X=0.217 $Y=2.255 $X2=0
+ $Y2=0
cc_473 N_A_27_297#_c_519_n N_VPWR_c_730_n 0.0419729f $X=1.115 $Y=2.36 $X2=0
+ $Y2=0
cc_474 N_A_27_297#_c_521_n N_VPWR_c_730_n 0.0549103f $X=2.07 $Y=2.36 $X2=0 $Y2=0
cc_475 N_A_27_297#_c_525_n N_VPWR_c_730_n 0.00196845f $X=3.01 $Y=1.92 $X2=0
+ $Y2=0
cc_476 N_A_27_297#_c_569_p N_VPWR_c_730_n 0.0118886f $X=1.2 $Y=2.34 $X2=0 $Y2=0
cc_477 N_A_27_297#_c_525_n N_VPWR_c_731_n 0.00265246f $X=3.01 $Y=1.92 $X2=0
+ $Y2=0
cc_478 N_A_27_297#_c_559_p N_VPWR_c_731_n 0.00929594f $X=3.095 $Y=2.26 $X2=0
+ $Y2=0
cc_479 N_A_27_297#_c_527_n N_VPWR_c_731_n 0.00196845f $X=3.95 $Y=1.92 $X2=0
+ $Y2=0
cc_480 N_A_27_297#_M1002_d N_VPWR_c_719_n 0.00217523f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_481 N_A_27_297#_M1016_d N_VPWR_c_719_n 0.00231272f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_482 N_A_27_297#_M1036_d N_VPWR_c_719_n 0.00273854f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_483 N_A_27_297#_M1007_d N_VPWR_c_719_n 0.00290587f $X=2.95 $Y=1.485 $X2=0
+ $Y2=0
cc_484 N_A_27_297#_M1034_d N_VPWR_c_719_n 0.00246452f $X=3.89 $Y=1.485 $X2=0
+ $Y2=0
cc_485 N_A_27_297#_c_513_n N_VPWR_c_719_n 0.0098205f $X=0.217 $Y=2.255 $X2=0
+ $Y2=0
cc_486 N_A_27_297#_c_519_n N_VPWR_c_719_n 0.0270046f $X=1.115 $Y=2.36 $X2=0
+ $Y2=0
cc_487 N_A_27_297#_c_521_n N_VPWR_c_719_n 0.0341783f $X=2.07 $Y=2.36 $X2=0 $Y2=0
cc_488 N_A_27_297#_c_525_n N_VPWR_c_719_n 0.0104808f $X=3.01 $Y=1.92 $X2=0 $Y2=0
cc_489 N_A_27_297#_c_559_p N_VPWR_c_719_n 0.00631544f $X=3.095 $Y=2.26 $X2=0
+ $Y2=0
cc_490 N_A_27_297#_c_527_n N_VPWR_c_719_n 0.0104808f $X=3.95 $Y=1.92 $X2=0 $Y2=0
cc_491 N_A_27_297#_c_516_n N_VPWR_c_719_n 0.00953181f $X=4.035 $Y=2.26 $X2=0
+ $Y2=0
cc_492 N_A_27_297#_c_569_p N_VPWR_c_719_n 0.00653405f $X=1.2 $Y=2.34 $X2=0 $Y2=0
cc_493 N_A_27_297#_c_516_n N_A_886_297#_c_868_n 0.0168365f $X=4.035 $Y=2.26
+ $X2=0 $Y2=0
cc_494 N_A_27_297#_c_515_n N_A_886_297#_c_869_n 0.0136296f $X=4.075 $Y=2.005
+ $X2=0 $Y2=0
cc_495 N_A_27_297#_c_516_n N_A_886_297#_c_869_n 0.0183843f $X=4.035 $Y=2.26
+ $X2=0 $Y2=0
cc_496 N_A_27_297#_c_514_n N_A_27_47#_c_1005_n 7.42972e-19 $X=0.26 $Y=1.66 $X2=0
+ $Y2=0
cc_497 N_Y_c_594_n N_VPWR_M1000_s 0.00351601f $X=4.86 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_498 N_Y_c_594_n N_VPWR_M1022_s 0.00351601f $X=4.86 $Y=1.58 $X2=0 $Y2=0
cc_499 N_Y_M1002_s N_VPWR_c_719_n 0.00232895f $X=0.585 $Y=1.485 $X2=0 $Y2=0
cc_500 N_Y_M1025_s N_VPWR_c_719_n 0.00232895f $X=1.525 $Y=1.485 $X2=0 $Y2=0
cc_501 N_Y_M1011_d N_VPWR_c_719_n 0.00232895f $X=4.88 $Y=1.485 $X2=0 $Y2=0
cc_502 N_Y_M1029_d N_VPWR_c_719_n 0.00232895f $X=5.82 $Y=1.485 $X2=0 $Y2=0
cc_503 N_Y_c_594_n N_A_886_297#_M1011_s 0.00504403f $X=4.86 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_504 N_Y_c_640_n N_A_886_297#_M1021_s 0.00342641f $X=5.75 $Y=1.58 $X2=0 $Y2=0
cc_505 N_Y_c_594_n N_A_886_297#_c_869_n 0.0201714f $X=4.86 $Y=1.58 $X2=0 $Y2=0
cc_506 N_Y_c_644_n N_A_886_297#_c_869_n 0.0155816f $X=5.025 $Y=1.66 $X2=0 $Y2=0
cc_507 N_Y_M1011_d N_A_886_297#_c_872_n 0.00354696f $X=4.88 $Y=1.485 $X2=0 $Y2=0
cc_508 N_Y_c_594_n N_A_886_297#_c_872_n 0.0039635f $X=4.86 $Y=1.58 $X2=0 $Y2=0
cc_509 N_Y_c_640_n N_A_886_297#_c_872_n 0.0039635f $X=5.75 $Y=1.58 $X2=0 $Y2=0
cc_510 N_Y_c_644_n N_A_886_297#_c_872_n 0.0162509f $X=5.025 $Y=1.66 $X2=0 $Y2=0
cc_511 N_Y_c_640_n N_A_886_297#_c_891_n 0.0135833f $X=5.75 $Y=1.58 $X2=0 $Y2=0
cc_512 N_Y_c_644_n N_A_886_297#_c_891_n 0.0151355f $X=5.025 $Y=1.66 $X2=0 $Y2=0
cc_513 N_Y_c_649_n N_A_886_297#_c_891_n 0.0186638f $X=5.965 $Y=1.66 $X2=0 $Y2=0
cc_514 N_Y_M1029_d N_A_886_297#_c_874_n 0.00354696f $X=5.82 $Y=1.485 $X2=0 $Y2=0
cc_515 N_Y_c_640_n N_A_886_297#_c_874_n 0.00273065f $X=5.75 $Y=1.58 $X2=0 $Y2=0
cc_516 N_Y_c_649_n N_A_886_297#_c_874_n 0.0198628f $X=5.965 $Y=1.66 $X2=0 $Y2=0
cc_517 N_Y_c_649_n N_A_886_297#_c_897_n 0.0153021f $X=5.965 $Y=1.66 $X2=0 $Y2=0
cc_518 N_Y_c_649_n N_A_1352_297#_c_939_n 0.0102243f $X=5.965 $Y=1.66 $X2=0 $Y2=0
cc_519 N_Y_c_590_n N_A_27_47#_M1026_d 0.0022437f $X=2.055 $Y=0.78 $X2=0 $Y2=0
cc_520 N_Y_c_702_p N_A_27_47#_M1038_d 0.00191657f $X=2.145 $Y=0.78 $X2=0 $Y2=0
cc_521 N_Y_c_592_n N_A_27_47#_M1024_d 0.0022437f $X=3.565 $Y=0.74 $X2=0 $Y2=0
cc_522 N_Y_c_590_n N_A_27_47#_c_1005_n 0.0200858f $X=2.055 $Y=0.78 $X2=0 $Y2=0
cc_523 N_Y_M1004_s N_A_27_47#_c_1022_n 0.00410554f $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_524 N_Y_M1027_s N_A_27_47#_c_1022_n 0.00410554f $X=1.535 $Y=0.235 $X2=0 $Y2=0
cc_525 N_Y_M1005_s N_A_27_47#_c_1022_n 0.00410554f $X=2.44 $Y=0.235 $X2=0 $Y2=0
cc_526 N_Y_M1028_s N_A_27_47#_c_1022_n 0.00519908f $X=3.38 $Y=0.235 $X2=0 $Y2=0
cc_527 N_Y_c_590_n N_A_27_47#_c_1022_n 0.0726287f $X=2.055 $Y=0.78 $X2=0 $Y2=0
cc_528 N_Y_c_592_n N_A_27_47#_c_1022_n 0.071066f $X=3.565 $Y=0.74 $X2=0 $Y2=0
cc_529 N_Y_c_702_p N_A_27_47#_c_1022_n 0.0121347f $X=2.145 $Y=0.78 $X2=0 $Y2=0
cc_530 N_Y_c_592_n N_A_27_47#_c_1006_n 0.00140356f $X=3.565 $Y=0.74 $X2=0 $Y2=0
cc_531 N_Y_c_594_n N_A_27_47#_c_1006_n 0.00745598f $X=4.86 $Y=1.58 $X2=0 $Y2=0
cc_532 N_Y_c_649_n N_A_27_47#_c_1014_n 0.00441221f $X=5.965 $Y=1.66 $X2=0 $Y2=0
cc_533 N_Y_M1004_s N_VGND_c_1195_n 0.00256987f $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_534 N_Y_M1027_s N_VGND_c_1195_n 0.00256987f $X=1.535 $Y=0.235 $X2=0 $Y2=0
cc_535 N_Y_M1005_s N_VGND_c_1195_n 0.00256987f $X=2.44 $Y=0.235 $X2=0 $Y2=0
cc_536 N_Y_M1028_s N_VGND_c_1195_n 0.00297142f $X=3.38 $Y=0.235 $X2=0 $Y2=0
cc_537 N_VPWR_c_719_n N_A_886_297#_M1011_s 0.00217523f $X=10.81 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_538 N_VPWR_c_719_n N_A_886_297#_M1021_s 0.00231272f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_719_n N_A_886_297#_M1037_s 0.00231272f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_719_n N_A_886_297#_M1008_s 0.00231272f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_719_n N_A_886_297#_M1018_s 0.00217523f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_542 N_VPWR_c_726_n N_A_886_297#_c_868_n 0.017537f $X=8.67 $Y=2.72 $X2=0 $Y2=0
cc_543 N_VPWR_c_719_n N_A_886_297#_c_868_n 0.00960883f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_544 N_VPWR_c_726_n N_A_886_297#_c_872_n 0.0419729f $X=8.67 $Y=2.72 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_719_n N_A_886_297#_c_872_n 0.0270046f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_726_n N_A_886_297#_c_874_n 0.0419729f $X=8.67 $Y=2.72 $X2=0
+ $Y2=0
cc_547 N_VPWR_c_719_n N_A_886_297#_c_874_n 0.0270046f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_548 N_VPWR_c_726_n N_A_886_297#_c_876_n 0.0419729f $X=8.67 $Y=2.72 $X2=0
+ $Y2=0
cc_549 N_VPWR_c_719_n N_A_886_297#_c_876_n 0.0270046f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_550 N_VPWR_c_726_n N_A_886_297#_c_878_n 0.0419729f $X=8.67 $Y=2.72 $X2=0
+ $Y2=0
cc_551 N_VPWR_c_719_n N_A_886_297#_c_878_n 0.0270046f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_552 N_VPWR_c_722_n N_A_886_297#_c_870_n 0.0168365f $X=8.835 $Y=2 $X2=0 $Y2=0
cc_553 N_VPWR_c_726_n N_A_886_297#_c_870_n 0.017537f $X=8.67 $Y=2.72 $X2=0 $Y2=0
cc_554 N_VPWR_c_719_n N_A_886_297#_c_870_n 0.00960883f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_555 N_VPWR_c_722_n N_A_886_297#_c_871_n 0.0309728f $X=8.835 $Y=2 $X2=0 $Y2=0
cc_556 N_VPWR_c_726_n N_A_886_297#_c_917_n 0.0118886f $X=8.67 $Y=2.72 $X2=0
+ $Y2=0
cc_557 N_VPWR_c_719_n N_A_886_297#_c_917_n 0.00653405f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_726_n N_A_886_297#_c_919_n 0.0118886f $X=8.67 $Y=2.72 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_719_n N_A_886_297#_c_919_n 0.00653405f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_560 N_VPWR_c_726_n N_A_886_297#_c_921_n 0.0118886f $X=8.67 $Y=2.72 $X2=0
+ $Y2=0
cc_561 N_VPWR_c_719_n N_A_886_297#_c_921_n 0.00653405f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_562 N_VPWR_c_719_n N_A_1352_297#_M1001_d 0.00232895f $X=10.81 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_563 N_VPWR_c_719_n N_A_1352_297#_M1014_d 0.00232895f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_564 N_VPWR_c_719_n N_A_1352_297#_M1003_d 0.00231261f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_565 N_VPWR_c_719_n N_A_1352_297#_M1023_d 0.00354185f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_566 N_VPWR_M1003_s N_A_1352_297#_c_938_n 0.00726124f $X=8.71 $Y=1.485 $X2=0
+ $Y2=0
cc_567 N_VPWR_c_722_n N_A_1352_297#_c_938_n 0.0202979f $X=8.835 $Y=2 $X2=0 $Y2=0
cc_568 N_VPWR_c_722_n N_A_1352_297#_c_956_n 0.0483931f $X=8.835 $Y=2 $X2=0 $Y2=0
cc_569 N_VPWR_c_723_n N_A_1352_297#_c_956_n 0.0385613f $X=9.775 $Y=2 $X2=0 $Y2=0
cc_570 N_VPWR_c_728_n N_A_1352_297#_c_956_n 0.0223557f $X=9.69 $Y=2.72 $X2=0
+ $Y2=0
cc_571 N_VPWR_c_719_n N_A_1352_297#_c_956_n 0.0140101f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_572 N_VPWR_M1010_s N_A_1352_297#_c_959_n 0.00342641f $X=9.63 $Y=1.485 $X2=0
+ $Y2=0
cc_573 N_VPWR_c_723_n N_A_1352_297#_c_959_n 0.0136682f $X=9.775 $Y=2 $X2=0 $Y2=0
cc_574 N_VPWR_c_723_n N_A_1352_297#_c_966_n 0.0470327f $X=9.775 $Y=2 $X2=0 $Y2=0
cc_575 N_VPWR_c_732_n N_A_1352_297#_c_966_n 0.0233349f $X=10.675 $Y=2.72 $X2=0
+ $Y2=0
cc_576 N_VPWR_c_719_n N_A_1352_297#_c_966_n 0.0141694f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_577 N_A_886_297#_c_876_n N_A_1352_297#_M1001_d 0.00354696f $X=7.29 $Y=2.36
+ $X2=-0.19 $Y2=1.305
cc_578 N_A_886_297#_c_878_n N_A_1352_297#_M1014_d 0.00354696f $X=8.23 $Y=2.36
+ $X2=0 $Y2=0
cc_579 N_A_886_297#_M1008_s N_A_1352_297#_c_940_n 0.00342641f $X=7.23 $Y=1.485
+ $X2=0 $Y2=0
cc_580 N_A_886_297#_c_876_n N_A_1352_297#_c_940_n 0.0039635f $X=7.29 $Y=2.36
+ $X2=0 $Y2=0
cc_581 N_A_886_297#_c_927_p N_A_1352_297#_c_940_n 0.0135833f $X=7.375 $Y=2 $X2=0
+ $Y2=0
cc_582 N_A_886_297#_c_878_n N_A_1352_297#_c_940_n 0.00273065f $X=8.23 $Y=2.36
+ $X2=0 $Y2=0
cc_583 N_A_886_297#_M1018_s N_A_1352_297#_c_938_n 0.00726124f $X=8.17 $Y=1.485
+ $X2=0 $Y2=0
cc_584 N_A_886_297#_c_878_n N_A_1352_297#_c_938_n 0.0039635f $X=8.23 $Y=2.36
+ $X2=0 $Y2=0
cc_585 N_A_886_297#_c_871_n N_A_1352_297#_c_938_n 0.0201715f $X=8.315 $Y=2 $X2=0
+ $Y2=0
cc_586 N_A_886_297#_c_897_n N_A_1352_297#_c_939_n 0.0186638f $X=6.435 $Y=2 $X2=0
+ $Y2=0
cc_587 N_A_886_297#_c_876_n N_A_1352_297#_c_939_n 0.0198628f $X=7.29 $Y=2.36
+ $X2=0 $Y2=0
cc_588 N_A_886_297#_c_927_p N_A_1352_297#_c_939_n 0.0153021f $X=7.375 $Y=2 $X2=0
+ $Y2=0
cc_589 N_A_886_297#_c_927_p N_A_1352_297#_c_950_n 0.0186638f $X=7.375 $Y=2 $X2=0
+ $Y2=0
cc_590 N_A_886_297#_c_878_n N_A_1352_297#_c_950_n 0.0198628f $X=8.23 $Y=2.36
+ $X2=0 $Y2=0
cc_591 N_A_886_297#_c_871_n N_A_1352_297#_c_950_n 0.0157482f $X=8.315 $Y=2 $X2=0
+ $Y2=0
cc_592 N_A_1352_297#_c_938_n N_A_27_47#_c_1016_n 0.0323114f $X=9.09 $Y=1.58
+ $X2=0 $Y2=0
cc_593 N_A_27_47#_c_1007_n N_VGND_M1012_s 0.00259473f $X=4.76 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_594 N_A_27_47#_c_1013_n N_VGND_M1017_s 0.00532376f $X=5.91 $Y=0.58 $X2=0
+ $Y2=0
cc_595 N_A_27_47#_c_1008_n N_VGND_M1006_s 0.00259473f $X=7.16 $Y=0.82 $X2=0
+ $Y2=0
cc_596 N_A_27_47#_c_1016_n N_VGND_M1019_s 0.00357604f $X=8.1 $Y=0.58 $X2=0 $Y2=0
cc_597 N_A_27_47#_c_1009_n N_VGND_M1015_s 0.00259473f $X=9.56 $Y=0.82 $X2=0
+ $Y2=0
cc_598 N_A_27_47#_c_1010_n N_VGND_M1032_s 0.00312516f $X=10.545 $Y=0.82 $X2=0
+ $Y2=0
cc_599 N_A_27_47#_c_1033_n N_VGND_c_1176_n 0.0135136f $X=4.075 $Y=0.465 $X2=0
+ $Y2=0
cc_600 N_A_27_47#_c_1006_n N_VGND_c_1176_n 0.00471242f $X=4.075 $Y=0.735 $X2=0
+ $Y2=0
cc_601 N_A_27_47#_c_1007_n N_VGND_c_1176_n 0.0115453f $X=4.76 $Y=0.82 $X2=0
+ $Y2=0
cc_602 N_A_27_47#_c_1041_n N_VGND_c_1177_n 0.0186586f $X=4.975 $Y=0.38 $X2=0
+ $Y2=0
cc_603 N_A_27_47#_c_1013_n N_VGND_c_1177_n 0.0229481f $X=5.91 $Y=0.58 $X2=0
+ $Y2=0
cc_604 N_A_27_47#_c_1008_n N_VGND_c_1178_n 0.0115453f $X=7.16 $Y=0.82 $X2=0
+ $Y2=0
cc_605 N_A_27_47#_c_1014_n N_VGND_c_1178_n 0.0173695f $X=6.58 $Y=0.58 $X2=0
+ $Y2=0
cc_606 N_A_27_47#_c_1056_n N_VGND_c_1179_n 0.0177507f $X=7.375 $Y=0.38 $X2=0
+ $Y2=0
cc_607 N_A_27_47#_c_1016_n N_VGND_c_1179_n 0.0119729f $X=8.1 $Y=0.58 $X2=0 $Y2=0
cc_608 N_A_27_47#_c_1017_n N_VGND_c_1179_n 0.0227149f $X=8.84 $Y=0.58 $X2=0
+ $Y2=0
cc_609 N_A_27_47#_c_1009_n N_VGND_c_1180_n 0.0115453f $X=9.56 $Y=0.82 $X2=0
+ $Y2=0
cc_610 N_A_27_47#_c_1017_n N_VGND_c_1180_n 0.0129622f $X=8.84 $Y=0.58 $X2=0
+ $Y2=0
cc_611 N_A_27_47#_c_1077_n N_VGND_c_1181_n 0.0180625f $X=9.775 $Y=0.38 $X2=0
+ $Y2=0
cc_612 N_A_27_47#_c_1010_n N_VGND_c_1181_n 0.0147523f $X=10.545 $Y=0.82 $X2=0
+ $Y2=0
cc_613 N_A_27_47#_c_1004_n N_VGND_c_1182_n 0.0179343f $X=0.217 $Y=0.465 $X2=0
+ $Y2=0
cc_614 N_A_27_47#_c_1022_n N_VGND_c_1182_n 0.202979f $X=3.95 $Y=0.36 $X2=0 $Y2=0
cc_615 N_A_27_47#_c_1033_n N_VGND_c_1182_n 0.0152108f $X=4.075 $Y=0.465 $X2=0
+ $Y2=0
cc_616 N_A_27_47#_c_1007_n N_VGND_c_1182_n 0.00260082f $X=4.76 $Y=0.82 $X2=0
+ $Y2=0
cc_617 N_A_27_47#_c_1007_n N_VGND_c_1184_n 0.00193763f $X=4.76 $Y=0.82 $X2=0
+ $Y2=0
cc_618 N_A_27_47#_c_1041_n N_VGND_c_1184_n 0.0223596f $X=4.975 $Y=0.38 $X2=0
+ $Y2=0
cc_619 N_A_27_47#_c_1013_n N_VGND_c_1184_n 0.00260082f $X=5.91 $Y=0.58 $X2=0
+ $Y2=0
cc_620 N_A_27_47#_c_1008_n N_VGND_c_1186_n 0.00286294f $X=7.16 $Y=0.82 $X2=0
+ $Y2=0
cc_621 N_A_27_47#_c_1013_n N_VGND_c_1186_n 0.00248202f $X=5.91 $Y=0.58 $X2=0
+ $Y2=0
cc_622 N_A_27_47#_c_1014_n N_VGND_c_1186_n 0.0433668f $X=6.58 $Y=0.58 $X2=0
+ $Y2=0
cc_623 N_A_27_47#_c_1008_n N_VGND_c_1188_n 0.00193763f $X=7.16 $Y=0.82 $X2=0
+ $Y2=0
cc_624 N_A_27_47#_c_1056_n N_VGND_c_1188_n 0.0223596f $X=7.375 $Y=0.38 $X2=0
+ $Y2=0
cc_625 N_A_27_47#_c_1016_n N_VGND_c_1188_n 0.00260082f $X=8.1 $Y=0.58 $X2=0
+ $Y2=0
cc_626 N_A_27_47#_c_1009_n N_VGND_c_1190_n 0.00445989f $X=9.56 $Y=0.82 $X2=0
+ $Y2=0
cc_627 N_A_27_47#_c_1016_n N_VGND_c_1190_n 0.00194552f $X=8.1 $Y=0.58 $X2=0
+ $Y2=0
cc_628 N_A_27_47#_c_1017_n N_VGND_c_1190_n 0.0493628f $X=8.84 $Y=0.58 $X2=0
+ $Y2=0
cc_629 N_A_27_47#_c_1009_n N_VGND_c_1192_n 0.00193763f $X=9.56 $Y=0.82 $X2=0
+ $Y2=0
cc_630 N_A_27_47#_c_1077_n N_VGND_c_1192_n 0.0223596f $X=9.775 $Y=0.38 $X2=0
+ $Y2=0
cc_631 N_A_27_47#_c_1010_n N_VGND_c_1192_n 0.00260082f $X=10.545 $Y=0.82 $X2=0
+ $Y2=0
cc_632 N_A_27_47#_c_1010_n N_VGND_c_1194_n 0.00193763f $X=10.545 $Y=0.82 $X2=0
+ $Y2=0
cc_633 N_A_27_47#_c_1011_n N_VGND_c_1194_n 0.0244796f $X=10.76 $Y=0.38 $X2=0
+ $Y2=0
cc_634 N_A_27_47#_M1004_d N_VGND_c_1195_n 0.00250318f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_635 N_A_27_47#_M1026_d N_VGND_c_1195_n 0.00255381f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_636 N_A_27_47#_M1038_d N_VGND_c_1195_n 0.00227273f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_637 N_A_27_47#_M1024_d N_VGND_c_1195_n 0.00255381f $X=2.91 $Y=0.235 $X2=0
+ $Y2=0
cc_638 N_A_27_47#_M1039_d N_VGND_c_1195_n 0.00215206f $X=3.9 $Y=0.235 $X2=0
+ $Y2=0
cc_639 N_A_27_47#_M1013_d N_VGND_c_1195_n 0.0025535f $X=4.79 $Y=0.235 $X2=0
+ $Y2=0
cc_640 N_A_27_47#_M1031_d N_VGND_c_1195_n 0.00559598f $X=5.89 $Y=0.235 $X2=0
+ $Y2=0
cc_641 N_A_27_47#_M1009_d N_VGND_c_1195_n 0.0025535f $X=7.19 $Y=0.235 $X2=0
+ $Y2=0
cc_642 N_A_27_47#_M1033_d N_VGND_c_1195_n 0.00707417f $X=8.18 $Y=0.235 $X2=0
+ $Y2=0
cc_643 N_A_27_47#_M1020_d N_VGND_c_1195_n 0.0025535f $X=9.59 $Y=0.235 $X2=0
+ $Y2=0
cc_644 N_A_27_47#_M1035_d N_VGND_c_1195_n 0.00250309f $X=10.575 $Y=0.235 $X2=0
+ $Y2=0
cc_645 N_A_27_47#_c_1004_n N_VGND_c_1195_n 0.00980895f $X=0.217 $Y=0.465 $X2=0
+ $Y2=0
cc_646 N_A_27_47#_c_1022_n N_VGND_c_1195_n 0.128846f $X=3.95 $Y=0.36 $X2=0 $Y2=0
cc_647 N_A_27_47#_c_1033_n N_VGND_c_1195_n 0.00940698f $X=4.075 $Y=0.465 $X2=0
+ $Y2=0
cc_648 N_A_27_47#_c_1007_n N_VGND_c_1195_n 0.00964063f $X=4.76 $Y=0.82 $X2=0
+ $Y2=0
cc_649 N_A_27_47#_c_1041_n N_VGND_c_1195_n 0.0141302f $X=4.975 $Y=0.38 $X2=0
+ $Y2=0
cc_650 N_A_27_47#_c_1008_n N_VGND_c_1195_n 0.0100655f $X=7.16 $Y=0.82 $X2=0
+ $Y2=0
cc_651 N_A_27_47#_c_1056_n N_VGND_c_1195_n 0.0141302f $X=7.375 $Y=0.38 $X2=0
+ $Y2=0
cc_652 N_A_27_47#_c_1009_n N_VGND_c_1195_n 0.0136855f $X=9.56 $Y=0.82 $X2=0
+ $Y2=0
cc_653 N_A_27_47#_c_1077_n N_VGND_c_1195_n 0.0141302f $X=9.775 $Y=0.38 $X2=0
+ $Y2=0
cc_654 N_A_27_47#_c_1010_n N_VGND_c_1195_n 0.00985487f $X=10.545 $Y=0.82 $X2=0
+ $Y2=0
cc_655 N_A_27_47#_c_1011_n N_VGND_c_1195_n 0.0143352f $X=10.76 $Y=0.38 $X2=0
+ $Y2=0
cc_656 N_A_27_47#_c_1013_n N_VGND_c_1195_n 0.0114569f $X=5.91 $Y=0.58 $X2=0
+ $Y2=0
cc_657 N_A_27_47#_c_1014_n N_VGND_c_1195_n 0.02564f $X=6.58 $Y=0.58 $X2=0 $Y2=0
cc_658 N_A_27_47#_c_1016_n N_VGND_c_1195_n 0.00993102f $X=8.1 $Y=0.58 $X2=0
+ $Y2=0
cc_659 N_A_27_47#_c_1017_n N_VGND_c_1195_n 0.0280109f $X=8.84 $Y=0.58 $X2=0
+ $Y2=0
