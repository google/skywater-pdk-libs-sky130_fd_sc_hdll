* NGSPICE file created from sky130_fd_sc_hdll__or4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
M1000 X a_335_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=1.20363e+12p ps=1.058e+07u
M1001 a_425_297# a_224_297# a_335_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.5e+11p pd=2.7e+06u as=2.7e+11p ps=2.54e+06u
M1002 VGND A a_335_297# VNB nshort w=650000u l=150000u
+  ad=1.2044e+12p pd=1.129e+07u as=4.355e+11p ps=3.94e+06u
M1003 VPWR A a_625_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1004 a_224_297# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1005 a_335_297# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_335_297# VGND VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=0p ps=0u
M1007 VPWR a_335_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND C_N a_27_410# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1009 a_625_297# B a_531_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1010 a_531_297# a_27_410# a_425_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_335_297# a_224_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_27_410# a_335_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_335_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR C_N a_27_410# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1015 X a_335_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_335_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_224_297# D_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1018 VPWR a_335_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_335_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

