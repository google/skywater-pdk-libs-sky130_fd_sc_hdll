* File: sky130_fd_sc_hdll__and3_4.spice
* Created: Wed Sep  2 08:22:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and3_4.pex.spice"
.subckt sky130_fd_sc_hdll__and3_4  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 A_185_47# N_A_M1002_g N_A_85_297#_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.160875 AS=0.19825 PD=1.145 PS=1.91 NRD=35.532 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1006 A_314_47# N_B_M1006_g A_185_47# VNB NSHORT L=0.15 W=0.65 AD=0.06825
+ AS=0.160875 PD=0.86 PS=1.145 NRD=9.228 NRS=35.532 M=1 R=4.33333 SA=75000.9
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_C_M1007_g A_314_47# VNB NSHORT L=0.15 W=0.65 AD=0.154375
+ AS=0.06825 PD=1.125 PS=0.86 NRD=27.684 NRS=9.228 M=1 R=4.33333 SA=75001.2
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1003_d N_A_85_297#_M1003_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.154375 PD=0.98 PS=1.125 NRD=9.228 NRS=8.304 M=1 R=4.33333
+ SA=75001.9 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1008 N_X_M1003_d N_A_85_297#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75002.3
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1011 N_X_M1011_d N_A_85_297#_M1011_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.10725 PD=1.03 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75002.8
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1012 N_X_M1011_d N_A_85_297#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.18525 PD=1.03 PS=1.87 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75003.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1013 N_VPWR_M1013_d N_A_M1013_g N_A_85_297#_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.2325 AS=0.31 PD=1.465 PS=2.62 NRD=24.6053 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.3 A=0.18 P=2.36 MULT=1
MM1001 N_A_85_297#_M1001_d N_B_M1001_g N_VPWR_M1013_d VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.2325 PD=1.3 PS=1.465 NRD=1.9503 NRS=11.8003 M=1 R=5.55556
+ SA=90000.9 SB=90002.7 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_C_M1009_g N_A_85_297#_M1001_d VPB PHIGHVT L=0.18 W=1
+ AD=0.1875 AS=0.15 PD=1.375 PS=1.3 NRD=8.8453 NRS=1.9503 M=1 R=5.55556
+ SA=90001.3 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1000 N_X_M1000_d N_A_85_297#_M1000_g N_VPWR_M1009_d VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.1875 PD=1.3 PS=1.375 NRD=1.9503 NRS=9.8303 M=1 R=5.55556
+ SA=90001.9 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1004 N_X_M1000_d N_A_85_297#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.4
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1005 N_X_M1005_d N_A_85_297#_M1005_g N_VPWR_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.9
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1010 N_X_M1005_d N_A_85_297#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90003.3
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
pX15_noxref noxref_12 C C PROBETYPE=1
*
.include "sky130_fd_sc_hdll__and3_4.pxi.spice"
*
.ends
*
*
