* File: sky130_fd_sc_hdll__clkinv_2.pxi.spice
* Created: Thu Aug 27 19:02:46 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKINV_2%A N_A_c_41_n N_A_M1001_g N_A_c_42_n N_A_M1002_g
+ N_A_M1000_g N_A_c_36_n N_A_c_37_n N_A_c_44_n N_A_M1004_g N_A_M1003_g
+ N_A_c_39_n A A A A A PM_SKY130_FD_SC_HDLL__CLKINV_2%A
x_PM_SKY130_FD_SC_HDLL__CLKINV_2%Y N_Y_M1000_s N_Y_M1001_d N_Y_M1002_d
+ N_Y_c_124_p N_Y_c_90_n N_Y_c_91_n N_Y_c_120_p N_Y_c_87_n Y Y Y N_Y_c_89_n Y
+ PM_SKY130_FD_SC_HDLL__CLKINV_2%Y
x_PM_SKY130_FD_SC_HDLL__CLKINV_2%VPWR N_VPWR_M1001_s N_VPWR_M1004_s
+ N_VPWR_c_136_n N_VPWR_c_137_n N_VPWR_c_138_n VPWR N_VPWR_c_139_n
+ N_VPWR_c_135_n N_VPWR_c_141_n N_VPWR_c_142_n
+ PM_SKY130_FD_SC_HDLL__CLKINV_2%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKINV_2%VGND N_VGND_M1000_d N_VGND_M1003_d
+ N_VGND_c_162_n N_VGND_c_163_n VGND N_VGND_c_164_n N_VGND_c_165_n
+ N_VGND_c_166_n N_VGND_c_167_n N_VGND_c_168_n N_VGND_c_169_n
+ PM_SKY130_FD_SC_HDLL__CLKINV_2%VGND
cc_1 VNB N_A_M1000_g 0.0430151f $X=-0.19 $Y=-0.24 $X2=1.04 $Y2=0.445
cc_2 VNB N_A_c_36_n 0.0183225f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=1.16
cc_3 VNB N_A_c_37_n 0.0811477f $X=-0.19 $Y=-0.24 $X2=1.115 $Y2=1.16
cc_4 VNB N_A_M1003_g 0.0365712f $X=-0.19 $Y=-0.24 $X2=1.52 $Y2=0.445
cc_5 VNB N_A_c_39_n 0.0141158f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=1.217
cc_6 VNB A 0.0140604f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.19
cc_7 VNB N_Y_c_87_n 0.00219255f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.105
cc_8 VNB Y 0.0238967f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_Y_c_89_n 0.0245153f $X=-0.19 $Y=-0.24 $X2=1.04 $Y2=1.212
cc_10 VNB N_VPWR_c_135_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_VGND_c_162_n 0.0211888f $X=-0.19 $Y=-0.24 $X2=1.04 $Y2=0.445
cc_12 VNB N_VGND_c_163_n 0.0157142f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=1.41
cc_13 VNB N_VGND_c_164_n 0.0199636f $X=-0.19 $Y=-0.24 $X2=1.52 $Y2=0.445
cc_14 VNB N_VGND_c_165_n 0.0158182f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.105
cc_15 VNB N_VGND_c_166_n 0.013929f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.16
cc_16 VNB N_VGND_c_167_n 0.16655f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.212
cc_17 VNB N_VGND_c_168_n 0.00661087f $X=-0.19 $Y=-0.24 $X2=1.05 $Y2=1.212
cc_18 VNB N_VGND_c_169_n 0.00577191f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.177
cc_19 VPB N_A_c_41_n 0.0205439f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.41
cc_20 VPB N_A_c_42_n 0.0162776f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.41
cc_21 VPB N_A_c_37_n 0.0223263f $X=-0.19 $Y=1.305 $X2=1.115 $Y2=1.16
cc_22 VPB N_A_c_44_n 0.019664f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=1.41
cc_23 VPB N_A_c_39_n 0.00766741f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=1.217
cc_24 VPB N_Y_c_90_n 0.00201747f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=1.985
cc_25 VPB N_Y_c_91_n 0.00853539f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=1.985
cc_26 VPB Y 0.00837634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB Y 0.0227786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB N_VPWR_c_136_n 0.00522213f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=1.16
cc_29 VPB N_VPWR_c_137_n 0.0204001f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=1.41
cc_30 VPB N_VPWR_c_138_n 0.00520816f $X=-0.19 $Y=1.305 $X2=1.52 $Y2=0.445
cc_31 VPB N_VPWR_c_139_n 0.016145f $X=-0.19 $Y=1.305 $X2=1.06 $Y2=1.105
cc_32 VPB N_VPWR_c_135_n 0.0598401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_141_n 0.0249217f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.212
cc_34 VPB N_VPWR_c_142_n 0.00487897f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.212
cc_35 N_A_c_41_n N_Y_c_90_n 0.0187135f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_36 N_A_c_42_n N_Y_c_90_n 0.0176117f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_37 N_A_c_37_n N_Y_c_90_n 0.00769645f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_38 A N_Y_c_90_n 0.0496881f $X=1.15 $Y=1.19 $X2=0 $Y2=0
cc_39 N_A_c_37_n N_Y_c_91_n 0.00589614f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_40 A N_Y_c_91_n 0.0209563f $X=1.15 $Y=1.19 $X2=0 $Y2=0
cc_41 N_A_M1000_g N_Y_c_87_n 0.00197368f $X=1.04 $Y=0.445 $X2=0 $Y2=0
cc_42 N_A_M1003_g N_Y_c_87_n 0.00454178f $X=1.52 $Y=0.445 $X2=0 $Y2=0
cc_43 N_A_c_42_n Y 2.39795e-19 $X=1 $Y=1.41 $X2=0 $Y2=0
cc_44 N_A_M1000_g Y 6.78834e-19 $X=1.04 $Y=0.445 $X2=0 $Y2=0
cc_45 N_A_c_37_n Y 5.69444e-19 $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_46 N_A_c_44_n Y 0.00224713f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_47 N_A_M1003_g Y 0.00630543f $X=1.52 $Y=0.445 $X2=0 $Y2=0
cc_48 N_A_c_39_n Y 0.0195369f $X=1.495 $Y=1.217 $X2=0 $Y2=0
cc_49 A Y 0.0174542f $X=1.15 $Y=1.19 $X2=0 $Y2=0
cc_50 N_A_c_37_n Y 0.00730986f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_51 N_A_c_44_n Y 0.0204201f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_52 N_A_c_39_n Y 3.54423e-19 $X=1.495 $Y=1.217 $X2=0 $Y2=0
cc_53 A Y 0.0184556f $X=1.15 $Y=1.19 $X2=0 $Y2=0
cc_54 N_A_M1000_g N_Y_c_89_n 0.00573988f $X=1.04 $Y=0.445 $X2=0 $Y2=0
cc_55 N_A_c_36_n N_Y_c_89_n 0.00347009f $X=1.395 $Y=1.16 $X2=0 $Y2=0
cc_56 N_A_M1003_g N_Y_c_89_n 0.0132947f $X=1.52 $Y=0.445 $X2=0 $Y2=0
cc_57 A N_Y_c_89_n 0.0153343f $X=1.15 $Y=1.19 $X2=0 $Y2=0
cc_58 N_A_c_41_n N_VPWR_c_136_n 0.00303578f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_59 N_A_c_42_n N_VPWR_c_136_n 0.00303578f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_60 N_A_c_42_n N_VPWR_c_137_n 0.00702461f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_61 N_A_c_44_n N_VPWR_c_137_n 0.00702461f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_62 N_A_c_44_n N_VPWR_c_138_n 0.00479709f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_63 N_A_c_41_n N_VPWR_c_135_n 0.0134823f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_64 N_A_c_42_n N_VPWR_c_135_n 0.0125774f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_65 N_A_c_44_n N_VPWR_c_135_n 0.0136509f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_66 N_A_c_41_n N_VPWR_c_141_n 0.00702461f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_67 N_A_M1000_g N_VGND_c_162_n 0.00515421f $X=1.04 $Y=0.445 $X2=0 $Y2=0
cc_68 N_A_c_37_n N_VGND_c_162_n 0.00703816f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_69 A N_VGND_c_162_n 0.0130871f $X=1.15 $Y=1.19 $X2=0 $Y2=0
cc_70 N_A_M1000_g N_VGND_c_163_n 6.45214e-19 $X=1.04 $Y=0.445 $X2=0 $Y2=0
cc_71 N_A_M1003_g N_VGND_c_163_n 0.0120485f $X=1.52 $Y=0.445 $X2=0 $Y2=0
cc_72 N_A_M1000_g N_VGND_c_165_n 0.00585385f $X=1.04 $Y=0.445 $X2=0 $Y2=0
cc_73 N_A_M1003_g N_VGND_c_165_n 0.00218133f $X=1.52 $Y=0.445 $X2=0 $Y2=0
cc_74 N_A_M1000_g N_VGND_c_167_n 0.0122475f $X=1.04 $Y=0.445 $X2=0 $Y2=0
cc_75 N_A_M1003_g N_VGND_c_167_n 0.00303238f $X=1.52 $Y=0.445 $X2=0 $Y2=0
cc_76 N_Y_c_90_n N_VPWR_M1001_s 0.00197722f $X=1.11 $Y=1.545 $X2=-0.19 $Y2=-0.24
cc_77 Y N_VPWR_M1004_s 0.00310571f $X=1.52 $Y=1.445 $X2=0 $Y2=0
cc_78 N_Y_c_90_n N_VPWR_c_136_n 0.0151327f $X=1.11 $Y=1.545 $X2=0 $Y2=0
cc_79 N_Y_c_120_p N_VPWR_c_137_n 0.0135664f $X=1.24 $Y=1.83 $X2=0 $Y2=0
cc_80 Y N_VPWR_c_138_n 0.0195651f $X=1.52 $Y=1.445 $X2=0 $Y2=0
cc_81 N_Y_M1001_d N_VPWR_c_135_n 0.00295932f $X=0.155 $Y=1.485 $X2=0 $Y2=0
cc_82 N_Y_M1002_d N_VPWR_c_135_n 0.00452262f $X=1.09 $Y=1.485 $X2=0 $Y2=0
cc_83 N_Y_c_124_p N_VPWR_c_135_n 0.00960102f $X=0.28 $Y=1.83 $X2=0 $Y2=0
cc_84 N_Y_c_120_p N_VPWR_c_135_n 0.00979076f $X=1.24 $Y=1.83 $X2=0 $Y2=0
cc_85 N_Y_c_124_p N_VPWR_c_141_n 0.0138754f $X=0.28 $Y=1.83 $X2=0 $Y2=0
cc_86 N_Y_c_87_n N_VGND_c_163_n 0.0209587f $X=1.255 $Y=0.445 $X2=0 $Y2=0
cc_87 N_Y_c_89_n N_VGND_c_163_n 0.0270926f $X=1.837 $Y=0.895 $X2=0 $Y2=0
cc_88 N_Y_c_87_n N_VGND_c_165_n 0.0118258f $X=1.255 $Y=0.445 $X2=0 $Y2=0
cc_89 N_Y_c_89_n N_VGND_c_165_n 0.00247477f $X=1.837 $Y=0.895 $X2=0 $Y2=0
cc_90 N_Y_c_89_n N_VGND_c_166_n 0.00387867f $X=1.837 $Y=0.895 $X2=0 $Y2=0
cc_91 N_Y_M1000_s N_VGND_c_167_n 0.00349695f $X=1.115 $Y=0.235 $X2=0 $Y2=0
cc_92 N_Y_c_87_n N_VGND_c_167_n 0.00838499f $X=1.255 $Y=0.445 $X2=0 $Y2=0
cc_93 N_Y_c_89_n N_VGND_c_167_n 0.0123932f $X=1.837 $Y=0.895 $X2=0 $Y2=0
