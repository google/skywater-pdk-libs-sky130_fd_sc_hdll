* File: sky130_fd_sc_hdll__nand4bb_1.pex.spice
* Created: Wed Sep  2 08:39:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_1%B_N 3 5 6 8 9 10 14 16
c33 16 0 7.02603e-20 $X=0.562 $Y=0.995
c34 9 0 6.28491e-20 $X=0.695 $Y=1.19
r35 14 17 37.7183 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.562 $Y=1.16
+ $X2=0.562 $Y2=1.325
r36 14 16 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.562 $Y=1.16
+ $X2=0.562 $Y2=0.995
r37 9 10 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.627 $Y=1.16
+ $X2=0.627 $Y2=1.53
r38 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.595
+ $Y=1.16 $X2=0.595 $Y2=1.16
r39 6 8 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r40 5 6 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.89 $X2=0.495
+ $Y2=1.99
r41 5 17 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.495 $Y=1.89
+ $X2=0.495 $Y2=1.325
r42 3 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.47 $Y=0.675
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_1%D 1 3 4 6 7
r35 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.16
+ $Y=1.16 $X2=1.16 $Y2=1.16
r36 4 10 46.2237 $w=3.35e-07 $l=2.89396e-07 $layer=POLY_cond $X=1.04 $Y=1.41
+ $X2=1.125 $Y2=1.16
r37 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.04 $Y=1.41 $X2=1.04
+ $Y2=1.985
r38 1 10 38.6365 $w=3.35e-07 $l=2.13014e-07 $layer=POLY_cond $X=1.015 $Y=0.995
+ $X2=1.125 $Y2=1.16
r39 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.015 $Y=0.995
+ $X2=1.015 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_1%C 1 3 4 6 7 8
c34 7 0 6.28491e-20 $X=1.59 $Y=0.765
r35 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.675
+ $Y=1.16 $X2=1.675 $Y2=1.16
r36 7 8 13.4814 $w=2.63e-07 $l=3.1e-07 $layer=LI1_cond $X=1.627 $Y=0.85
+ $X2=1.627 $Y2=1.16
r37 4 12 49.9093 $w=2.71e-07 $l=2.7157e-07 $layer=POLY_cond $X=1.62 $Y=1.41
+ $X2=1.665 $Y2=1.16
r38 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.62 $Y=1.41 $X2=1.62
+ $Y2=1.985
r39 1 12 38.8824 $w=2.71e-07 $l=1.96914e-07 $layer=POLY_cond $X=1.595 $Y=0.995
+ $X2=1.665 $Y2=1.16
r40 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.595 $Y=0.995
+ $X2=1.595 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_1%A_27_93# 1 2 7 9 10 12 15 18 19 20 23 27
+ 32 33
c85 20 0 7.02603e-20 $X=1.22 $Y=0.46
r86 32 33 12.0264 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=0.255 $Y=2.34
+ $X2=0.255 $Y2=2.065
r87 30 33 73.5169 $w=1.73e-07 $l=1.16e-06 $layer=LI1_cond $X=0.172 $Y=0.905
+ $X2=0.172 $Y2=2.065
r88 29 30 5.92518 $w=3.38e-07 $l=9.5e-08 $layer=LI1_cond $X=0.255 $Y=0.81
+ $X2=0.255 $Y2=0.905
r89 27 29 6.77908 $w=3.38e-07 $l=2e-07 $layer=LI1_cond $X=0.255 $Y=0.61
+ $X2=0.255 $Y2=0.81
r90 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.155
+ $Y=1.16 $X2=2.155 $Y2=1.16
r91 21 23 27.8891 $w=2.48e-07 $l=6.05e-07 $layer=LI1_cond $X=2.115 $Y=0.555
+ $X2=2.115 $Y2=1.16
r92 19 21 6.98266 $w=1.9e-07 $l=1.65831e-07 $layer=LI1_cond $X=1.99 $Y=0.46
+ $X2=2.115 $Y2=0.555
r93 19 20 44.9474 $w=1.88e-07 $l=7.7e-07 $layer=LI1_cond $X=1.99 $Y=0.46
+ $X2=1.22 $Y2=0.46
r94 17 20 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.135 $Y=0.555
+ $X2=1.22 $Y2=0.46
r95 17 18 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.135 $Y=0.555
+ $X2=1.135 $Y2=0.715
r96 16 29 4.14298 $w=1.9e-07 $l=1.7e-07 $layer=LI1_cond $X=0.425 $Y=0.81
+ $X2=0.255 $Y2=0.81
r97 15 18 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.05 $Y=0.81
+ $X2=1.135 $Y2=0.715
r98 15 16 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=1.05 $Y=0.81
+ $X2=0.425 $Y2=0.81
r99 10 24 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.12 $Y=1.41
+ $X2=2.155 $Y2=1.16
r100 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.12 $Y=1.41
+ $X2=2.12 $Y2=1.985
r101 7 24 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.095 $Y=0.995
+ $X2=2.155 $Y2=1.16
r102 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.095 $Y=0.995
+ $X2=2.095 $Y2=0.56
r103 2 32 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.34
r104 1 27 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_1%A_500_21# 1 2 7 9 10 12 15 18 19 22 25
+ 29 31 33
r68 32 33 3.35655 $w=3.59e-07 $l=2.5e-08 $layer=POLY_cond $X=2.575 $Y=1.202
+ $X2=2.6 $Y2=1.202
r69 27 29 3.77524 $w=2.88e-07 $l=9.5e-08 $layer=LI1_cond $X=3.875 $Y=0.4
+ $X2=3.97 $Y2=0.4
r70 25 31 3.80849 $w=2.42e-07 $l=1.15888e-07 $layer=LI1_cond $X=3.97 $Y=1.835
+ $X2=3.897 $Y2=1.92
r71 24 29 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.97 $Y=0.545
+ $X2=3.97 $Y2=0.4
r72 24 25 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=3.97 $Y=0.545
+ $X2=3.97 $Y2=1.835
r73 20 31 3.80849 $w=2.42e-07 $l=8.5e-08 $layer=LI1_cond $X=3.897 $Y=2.005
+ $X2=3.897 $Y2=1.92
r74 20 22 10.7927 $w=3.13e-07 $l=2.95e-07 $layer=LI1_cond $X=3.897 $Y=2.005
+ $X2=3.897 $Y2=2.3
r75 18 31 2.64776 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=3.74 $Y=1.92
+ $X2=3.897 $Y2=1.92
r76 18 19 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.74 $Y=1.92
+ $X2=3.125 $Y2=1.92
r77 16 33 44.9777 $w=3.59e-07 $l=3.35e-07 $layer=POLY_cond $X=2.935 $Y=1.202
+ $X2=2.6 $Y2=1.202
r78 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.935
+ $Y=1.16 $X2=2.935 $Y2=1.16
r79 13 19 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=2.987 $Y=1.835
+ $X2=3.125 $Y2=1.92
r80 13 15 28.2872 $w=2.73e-07 $l=6.75e-07 $layer=LI1_cond $X=2.987 $Y=1.835
+ $X2=2.987 $Y2=1.16
r81 10 33 18.9031 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.6 $Y=1.41 $X2=2.6
+ $Y2=1.202
r82 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.6 $Y=1.41 $X2=2.6
+ $Y2=1.985
r83 7 32 23.2387 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.575 $Y=0.995
+ $X2=2.575 $Y2=1.202
r84 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.575 $Y=0.995
+ $X2=2.575 $Y2=0.56
r85 2 22 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=3.68
+ $Y=2.065 $X2=3.825 $Y2=2.3
r86 1 27 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=3.64
+ $Y=0.235 $X2=3.875 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_1%A_N 3 6 7 9 10 11 12 17
r37 17 20 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.65 $Y=1.155
+ $X2=3.65 $Y2=1.32
r38 17 19 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.65 $Y=1.155
+ $X2=3.65 $Y2=0.99
r39 11 12 10.5406 $w=4.08e-07 $l=3.75e-07 $layer=LI1_cond $X=3.505 $Y=1.155
+ $X2=3.505 $Y2=1.53
r40 11 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.625
+ $Y=1.155 $X2=3.625 $Y2=1.155
r41 10 11 8.57305 $w=4.08e-07 $l=3.05e-07 $layer=LI1_cond $X=3.505 $Y=0.85
+ $X2=3.505 $Y2=1.155
r42 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.59 $Y=1.99 $X2=3.59
+ $Y2=2.275
r43 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.59 $Y=1.89 $X2=3.59
+ $Y2=1.99
r44 6 20 188.999 $w=2e-07 $l=5.7e-07 $layer=POLY_cond $X=3.59 $Y=1.89 $X2=3.59
+ $Y2=1.32
r45 3 19 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.565 $Y=0.445
+ $X2=3.565 $Y2=0.99
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_1%VPWR 1 2 3 14 18 21 22 23 35 36 39 44 47
r61 46 47 10.3517 $w=6.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=2.49
+ $X2=3.52 $Y2=2.49
r62 42 46 6.92966 $w=6.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.99 $Y=2.49
+ $X2=3.355 $Y2=2.49
r63 42 44 11.7756 $w=6.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.99 $Y=2.49
+ $X2=2.75 $Y2=2.49
r64 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r65 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r66 36 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=2.99 $Y2=2.72
r67 35 47 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=3.52 $Y2=2.72
r68 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r69 32 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r70 31 44 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=2.75 $Y2=2.72
r71 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r72 28 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r73 28 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r74 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r75 25 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=2.72
+ $X2=0.81 $Y2=2.72
r76 25 27 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.975 $Y=2.72
+ $X2=1.61 $Y2=2.72
r77 23 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r78 21 27 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=2.72
+ $X2=1.61 $Y2=2.72
r79 21 22 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=1.695 $Y=2.72
+ $X2=1.855 $Y2=2.72
r80 20 31 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.015 $Y=2.72
+ $X2=2.53 $Y2=2.72
r81 20 22 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=2.015 $Y=2.72
+ $X2=1.855 $Y2=2.72
r82 16 22 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=2.635
+ $X2=1.855 $Y2=2.72
r83 16 18 22.8688 $w=3.18e-07 $l=6.35e-07 $layer=LI1_cond $X=1.855 $Y=2.635
+ $X2=1.855 $Y2=2
r84 12 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=2.635
+ $X2=0.81 $Y2=2.72
r85 12 14 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.81 $Y=2.635
+ $X2=0.81 $Y2=2
r86 3 46 300 $w=1.7e-07 $l=1.14e-06 $layer=licon1_PDIFF $count=2 $X=2.69
+ $Y=1.485 $X2=3.355 $Y2=2.34
r87 2 18 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=1.71
+ $Y=1.485 $X2=1.86 $Y2=2
r88 1 14 300 $w=1.7e-07 $l=2.40312e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=2.065 $X2=0.795 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_1%Y 1 2 3 10 12 14 18 22 23 24 25 35 41 48
r47 53 54 8.95361 $w=4.88e-07 $l=3.45e-07 $layer=LI1_cond $X=2.435 $Y=1.66
+ $X2=2.435 $Y2=2.005
r48 51 53 1.95278 $w=4.88e-07 $l=8e-08 $layer=LI1_cond $X=2.435 $Y=1.58
+ $X2=2.435 $Y2=1.66
r49 48 49 3.24739 $w=4.88e-07 $l=3.5e-08 $layer=LI1_cond $X=2.435 $Y=1.53
+ $X2=2.435 $Y2=1.495
r50 35 46 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.545 $Y=0.85
+ $X2=2.545 $Y2=0.825
r51 25 51 0.610244 $w=4.88e-07 $l=2.5e-08 $layer=LI1_cond $X=2.435 $Y=1.555
+ $X2=2.435 $Y2=1.58
r52 25 48 0.610244 $w=4.88e-07 $l=2.5e-08 $layer=LI1_cond $X=2.435 $Y=1.555
+ $X2=2.435 $Y2=1.53
r53 25 49 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.545 $Y=1.47
+ $X2=2.545 $Y2=1.495
r54 24 25 11.9513 $w=2.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.545 $Y=1.19
+ $X2=2.545 $Y2=1.47
r55 23 46 4.1624 $w=5.88e-07 $l=3e-08 $layer=LI1_cond $X=2.705 $Y=0.795
+ $X2=2.705 $Y2=0.825
r56 23 24 13.2318 $w=2.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.545 $Y=0.88
+ $X2=2.545 $Y2=1.19
r57 23 35 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=2.545 $Y=0.88
+ $X2=2.545 $Y2=0.85
r58 22 23 5.77767 $w=5.88e-07 $l=2.85e-07 $layer=LI1_cond $X=2.705 $Y=0.51
+ $X2=2.705 $Y2=0.795
r59 22 41 2.63543 $w=5.88e-07 $l=1.3e-07 $layer=LI1_cond $X=2.705 $Y=0.51
+ $X2=2.705 $Y2=0.38
r60 18 54 9.89919 $w=3.88e-07 $l=3.35e-07 $layer=LI1_cond $X=2.385 $Y=2.34
+ $X2=2.385 $Y2=2.005
r61 15 21 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=1.58
+ $X2=1.32 $Y2=1.58
r62 14 51 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=2.19 $Y=1.58
+ $X2=2.435 $Y2=1.58
r63 14 15 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.19 $Y=1.58
+ $X2=1.485 $Y2=1.58
r64 10 21 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.32 $Y=1.665 $X2=1.32
+ $Y2=1.58
r65 10 12 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.32 $Y=1.665
+ $X2=1.32 $Y2=2.34
r66 3 53 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.21
+ $Y=1.485 $X2=2.355 $Y2=1.66
r67 3 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.21
+ $Y=1.485 $X2=2.355 $Y2=2.34
r68 2 21 400 $w=1.7e-07 $l=2.63344e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=1.485 $X2=1.32 $Y2=1.66
r69 2 12 400 $w=1.7e-07 $l=9.45238e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=1.485 $X2=1.32 $Y2=2.34
r70 1 41 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=2.65
+ $Y=0.235 $X2=2.835 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_1%VGND 1 2 11 15 17 19 29 30 33 36
r50 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r51 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r52 30 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=3.45
+ $Y2=0
r53 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r54 27 36 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.54 $Y=0 $X2=3.365
+ $Y2=0
r55 27 29 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.54 $Y=0 $X2=3.91
+ $Y2=0
r56 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r57 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r58 23 26 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r59 23 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r60 22 25 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r61 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r62 20 33 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.762
+ $Y2=0
r63 20 22 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=1.15
+ $Y2=0
r64 19 36 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.19 $Y=0 $X2=3.365
+ $Y2=0
r65 19 25 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.19 $Y=0 $X2=2.99
+ $Y2=0
r66 17 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r67 13 36 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.365 $Y=0.085
+ $X2=3.365 $Y2=0
r68 13 15 9.71345 $w=3.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.365 $Y=0.085
+ $X2=3.365 $Y2=0.38
r69 9 33 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.762 $Y=0.085
+ $X2=0.762 $Y2=0
r70 9 11 14.4668 $w=2.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.762 $Y=0.085
+ $X2=0.762 $Y2=0.38
r71 2 15 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.23
+ $Y=0.235 $X2=3.355 $Y2=0.38
r72 1 11 182 $w=1.7e-07 $l=2.89396e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.465 $X2=0.795 $Y2=0.38
.ends

