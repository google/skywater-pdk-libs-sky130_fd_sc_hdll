* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
X0 X a_197_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VPWR a_197_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 VGND a_197_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND A2 a_635_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_197_21# a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 a_27_297# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_635_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_197_21# A2 a_823_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VPWR A1 a_823_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 X a_197_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 X a_197_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 a_823_297# A2 a_197_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 VPWR a_197_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 a_635_47# a_27_297# a_197_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 X a_197_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_635_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR a_27_297# a_197_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_27_297# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_823_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 VGND A1 a_635_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VGND a_197_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_197_21# a_27_297# a_635_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
