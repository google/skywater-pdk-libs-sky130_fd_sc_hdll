* NGSPICE file created from sky130_fd_sc_hdll__isobufsrc_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__isobufsrc_2 A SLEEP VGND VNB VPB VPWR X
M1000 VPWR SLEEP a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=4.034e+11p pd=3.96e+06u as=8.5e+11p ps=7.7e+06u
M1001 VGND A a_271_21# VNB nshort w=420000u l=150000u
+  ad=6.5345e+11p pd=6.97e+06u as=1.092e+11p ps=1.36e+06u
M1002 a_27_297# a_271_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1003 X a_271_21# a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=4.81e+11p pd=4.08e+06u as=0p ps=0u
M1005 VGND a_271_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A a_271_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1007 a_27_297# SLEEP VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_271_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND SLEEP X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

