# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__sdfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.755000 1.355000 3.125000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.960000 0.305000 10.440000 0.825000 ;
        RECT  9.980000 1.505000 10.440000 2.465000 ;
        RECT 10.220000 0.825000 10.440000 1.505000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.615000 0.265000 11.870000 2.325000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 1.055000 4.345000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.860000 0.615000 3.535000 0.785000 ;
        RECT 1.860000 0.785000 2.030000 1.685000 ;
        RECT 3.315000 0.785000 3.535000 1.115000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.150000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.860000 0.805000 ;
      RECT  0.175000  1.795000  0.895000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  0.515000  2.135000  0.895000 2.635000 ;
      RECT  0.665000  0.805000  0.860000 0.970000 ;
      RECT  0.665000  0.970000  0.895000 1.795000 ;
      RECT  1.115000  0.345000  1.285000 2.465000 ;
      RECT  1.520000  0.255000  1.905000 0.445000 ;
      RECT  1.520000  0.445000  1.690000 1.860000 ;
      RECT  1.520000  1.860000  3.530000 2.075000 ;
      RECT  1.520000  2.075000  1.805000 2.445000 ;
      RECT  1.975000  2.245000  2.355000 2.635000 ;
      RECT  2.145000  0.085000  2.475000 0.445000 ;
      RECT  2.250000  0.955000  2.695000 1.125000 ;
      RECT  2.250000  1.125000  2.420000 1.860000 ;
      RECT  2.875000  2.245000  3.870000 2.415000 ;
      RECT  3.050000  0.275000  3.875000 0.445000 ;
      RECT  3.335000  1.355000  3.555000 1.685000 ;
      RECT  3.335000  1.685000  3.530000 1.860000 ;
      RECT  3.700000  1.825000  4.685000 1.995000 ;
      RECT  3.700000  1.995000  3.870000 2.245000 ;
      RECT  3.705000  0.445000  3.875000 0.715000 ;
      RECT  3.705000  0.715000  4.685000 0.885000 ;
      RECT  4.090000  2.165000  4.260000 2.635000 ;
      RECT  4.095000  0.085000  4.295000 0.545000 ;
      RECT  4.515000  0.365000  4.865000 0.535000 ;
      RECT  4.515000  0.535000  4.685000 0.715000 ;
      RECT  4.515000  0.885000  4.685000 1.825000 ;
      RECT  4.515000  1.995000  4.685000 2.070000 ;
      RECT  4.515000  2.070000  4.800000 2.440000 ;
      RECT  4.855000  0.705000  5.485000 1.035000 ;
      RECT  4.855000  1.035000  5.145000 1.905000 ;
      RECT  4.995000  2.190000  6.215000 2.360000 ;
      RECT  5.085000  0.365000  5.875000 0.535000 ;
      RECT  5.335000  1.655000  5.825000 2.010000 ;
      RECT  5.705000  0.535000  5.875000 1.315000 ;
      RECT  5.705000  1.315000  6.555000 1.485000 ;
      RECT  5.995000  1.485000  6.555000 1.575000 ;
      RECT  5.995000  1.575000  6.215000 2.190000 ;
      RECT  6.095000  0.765000  6.945000 1.065000 ;
      RECT  6.095000  1.065000  6.265000 1.095000 ;
      RECT  6.175000  0.085000  6.545000 0.585000 ;
      RECT  6.385000  1.245000  6.555000 1.315000 ;
      RECT  6.385000  1.835000  6.555000 2.635000 ;
      RECT  6.725000  0.365000  7.235000 0.535000 ;
      RECT  6.725000  0.535000  6.945000 0.765000 ;
      RECT  6.725000  1.065000  6.945000 2.135000 ;
      RECT  6.725000  2.135000  7.025000 2.465000 ;
      RECT  7.115000  0.705000  7.715000 1.035000 ;
      RECT  7.115000  1.245000  7.355000 1.965000 ;
      RECT  7.250000  2.165000  8.285000 2.335000 ;
      RECT  7.515000  0.365000  8.155000 0.535000 ;
      RECT  7.525000  1.035000  7.715000 1.575000 ;
      RECT  7.525000  1.575000  7.895000 1.905000 ;
      RECT  7.935000  0.535000  8.155000 0.995000 ;
      RECT  7.935000  0.995000  9.045000 1.325000 ;
      RECT  7.935000  1.325000  8.285000 1.405000 ;
      RECT  8.115000  1.405000  8.285000 2.165000 ;
      RECT  8.380000  0.085000  8.800000 0.615000 ;
      RECT  8.485000  1.575000  9.400000 1.905000 ;
      RECT  8.515000  2.135000  8.820000 2.635000 ;
      RECT  9.070000  0.300000  9.400000 0.825000 ;
      RECT  9.110000  1.905000  9.400000 2.455000 ;
      RECT  9.215000  0.825000  9.400000 0.995000 ;
      RECT  9.215000  0.995000 10.050000 1.325000 ;
      RECT  9.215000  1.325000  9.400000 1.575000 ;
      RECT  9.620000  0.085000  9.790000 0.695000 ;
      RECT  9.620000  1.625000  9.790000 2.635000 ;
      RECT 10.610000  0.345000 10.860000 0.995000 ;
      RECT 10.610000  0.995000 11.440000 1.325000 ;
      RECT 10.610000  1.325000 10.860000 2.425000 ;
      RECT 11.065000  0.085000 11.395000 0.805000 ;
      RECT 11.090000  1.495000 11.395000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.695000  1.785000  0.865000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.115000  0.425000  1.285000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  0.765000  5.375000 0.935000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.615000  1.785000  5.785000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.175000  1.785000  7.345000 1.955000 ;
      RECT  7.185000  0.765000  7.355000 0.935000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
    LAYER met1 ;
      RECT 0.635000 1.755000 0.925000 1.800000 ;
      RECT 0.635000 1.800000 7.405000 1.940000 ;
      RECT 0.635000 1.940000 0.925000 1.985000 ;
      RECT 1.005000 0.395000 1.345000 0.440000 ;
      RECT 1.005000 0.440000 5.285000 0.580000 ;
      RECT 1.005000 0.580000 1.345000 0.625000 ;
      RECT 5.145000 0.580000 5.285000 0.735000 ;
      RECT 5.145000 0.735000 5.435000 0.780000 ;
      RECT 5.145000 0.780000 7.415000 0.920000 ;
      RECT 5.145000 0.920000 5.435000 0.965000 ;
      RECT 5.555000 1.755000 5.845000 1.800000 ;
      RECT 5.555000 1.940000 5.845000 1.985000 ;
      RECT 7.115000 1.755000 7.405000 1.800000 ;
      RECT 7.115000 1.940000 7.405000 1.985000 ;
      RECT 7.125000 0.735000 7.415000 0.780000 ;
      RECT 7.125000 0.920000 7.415000 0.965000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfxbp_1
END LIBRARY
