# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__muxb16to1_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__muxb16to1_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  51.98000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D[0]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.395000 1.055000 1.785000 1.325000 ;
    END
  END D[0]
  PIN D[1]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.095000 1.055000 12.485000 1.325000 ;
    END
  END D[1]
  PIN D[2]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.275000 1.055000 14.665000 1.325000 ;
    END
  END D[2]
  PIN D[3]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 23.975000 1.055000 25.365000 1.325000 ;
    END
  END D[3]
  PIN D[4]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 26.615000 1.055000 28.005000 1.325000 ;
    END
  END D[4]
  PIN D[5]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 37.315000 1.055000 38.705000 1.325000 ;
    END
  END D[5]
  PIN D[6]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 39.495000 1.055000 40.885000 1.325000 ;
    END
  END D[6]
  PIN D[7]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 50.195000 1.055000 51.585000 1.325000 ;
    END
  END D[7]
  PIN D[8]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.395000 4.115000 1.785000 4.385000 ;
    END
  END D[8]
  PIN D[9]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.095000 4.115000 12.485000 4.385000 ;
    END
  END D[9]
  PIN D[10]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.275000 4.115000 14.665000 4.385000 ;
    END
  END D[10]
  PIN D[11]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 23.975000 4.115000 25.365000 4.385000 ;
    END
  END D[11]
  PIN D[12]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 26.615000 4.115000 28.005000 4.385000 ;
    END
  END D[12]
  PIN D[13]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 37.315000 4.115000 38.705000 4.385000 ;
    END
  END D[13]
  PIN D[14]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 39.495000 4.115000 40.885000 4.385000 ;
    END
  END D[14]
  PIN D[15]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 50.195000 4.115000 51.585000 4.385000 ;
    END
  END D[15]
  PIN S[0]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.760000 0.995000 6.355000 1.325000 ;
    END
  END S[0]
  PIN S[1]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.525000 0.995000 7.120000 1.325000 ;
    END
  END S[1]
  PIN S[2]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.640000 0.995000 19.235000 1.325000 ;
    END
  END S[2]
  PIN S[3]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.405000 0.995000 20.000000 1.325000 ;
    END
  END S[3]
  PIN S[4]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 31.980000 0.995000 32.575000 1.325000 ;
    END
  END S[4]
  PIN S[5]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 32.745000 0.995000 33.340000 1.325000 ;
    END
  END S[5]
  PIN S[6]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 44.860000 0.995000 45.455000 1.325000 ;
    END
  END S[6]
  PIN S[7]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 45.625000 0.995000 46.220000 1.325000 ;
    END
  END S[7]
  PIN S[8]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.760000 4.115000 6.355000 4.445000 ;
    END
  END S[8]
  PIN S[9]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.525000 4.115000 7.120000 4.445000 ;
    END
  END S[9]
  PIN S[10]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.640000 4.115000 19.235000 4.445000 ;
    END
  END S[10]
  PIN S[11]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.405000 4.115000 20.000000 4.445000 ;
    END
  END S[11]
  PIN S[12]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 31.980000 4.115000 32.575000 4.445000 ;
    END
  END S[12]
  PIN S[13]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 32.745000 4.115000 33.340000 4.445000 ;
    END
  END S[13]
  PIN S[14]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 44.860000 4.115000 45.455000 4.445000 ;
    END
  END S[14]
  PIN S[15]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 45.625000 4.115000 46.220000 4.445000 ;
    END
  END S[15]
  PIN VNB
    ANTENNADIFFAREA  0.089250 ;
    PORT
      LAYER li1 ;
        RECT 25.845000 0.265000 26.135000 0.810000 ;
    END
    PORT
      LAYER li1 ;
        RECT 25.845000 4.630000 26.135000 5.175000 ;
    END
  END VNB
  PIN VPB
    ANTENNADIFFAREA  0.297500 ;
    PORT
      LAYER li1 ;
        RECT 25.845000 1.470000 26.135000 2.455000 ;
        RECT 25.845000 2.985000 26.135000 3.970000 ;
    END
  END VPB
  PIN Z
    ANTENNADIFFAREA  12.10240 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865000 0.595000 3.195000 0.885000 ;
        RECT 2.865000 4.555000 3.195000 4.845000 ;
        RECT 2.965000 0.885000 3.195000 1.065000 ;
        RECT 2.965000 1.065000 4.235000 1.365000 ;
        RECT 2.965000 1.365000 3.295000 4.075000 ;
        RECT 2.965000 4.075000 4.235000 4.375000 ;
        RECT 2.965000 4.375000 3.195000 4.555000 ;
        RECT 3.705000 0.595000 4.035000 1.065000 ;
        RECT 3.705000 4.375000 4.035000 4.845000 ;
        RECT 3.905000 1.365000 4.235000 4.075000 ;
      LAYER mcon ;
        RECT 3.045000 1.785000 3.215000 1.955000 ;
        RECT 3.045000 3.485000 3.215000 3.655000 ;
        RECT 3.985000 1.785000 4.155000 1.955000 ;
        RECT 3.985000 3.485000 4.155000 3.655000 ;
    END
    PORT
      LAYER met1 ;
        RECT  2.985000 1.755000  3.275000 1.800000 ;
        RECT  2.985000 1.800000 48.995000 1.940000 ;
        RECT  2.985000 1.940000  3.275000 1.985000 ;
        RECT  2.985000 3.455000  3.275000 3.500000 ;
        RECT  2.985000 3.500000 48.995000 3.640000 ;
        RECT  2.985000 3.640000  3.275000 3.685000 ;
        RECT  3.925000 1.755000  4.215000 1.800000 ;
        RECT  3.925000 1.940000  4.215000 1.985000 ;
        RECT  3.925000 3.455000  4.215000 3.500000 ;
        RECT  3.925000 3.640000  4.215000 3.685000 ;
        RECT  8.665000 1.755000  8.955000 1.800000 ;
        RECT  8.665000 1.940000  8.955000 1.985000 ;
        RECT  8.665000 3.455000  8.955000 3.500000 ;
        RECT  8.665000 3.640000  8.955000 3.685000 ;
        RECT  9.605000 1.755000  9.895000 1.800000 ;
        RECT  9.605000 1.940000  9.895000 1.985000 ;
        RECT  9.605000 3.455000  9.895000 3.500000 ;
        RECT  9.605000 3.640000  9.895000 3.685000 ;
        RECT 15.865000 1.755000 16.155000 1.800000 ;
        RECT 15.865000 1.940000 16.155000 1.985000 ;
        RECT 15.865000 3.455000 16.155000 3.500000 ;
        RECT 15.865000 3.640000 16.155000 3.685000 ;
        RECT 16.805000 1.755000 17.095000 1.800000 ;
        RECT 16.805000 1.940000 17.095000 1.985000 ;
        RECT 16.805000 3.455000 17.095000 3.500000 ;
        RECT 16.805000 3.640000 17.095000 3.685000 ;
        RECT 21.545000 1.755000 21.835000 1.800000 ;
        RECT 21.545000 1.940000 21.835000 1.985000 ;
        RECT 21.545000 3.455000 21.835000 3.500000 ;
        RECT 21.545000 3.640000 21.835000 3.685000 ;
        RECT 22.485000 1.755000 22.775000 1.800000 ;
        RECT 22.485000 1.940000 22.775000 1.985000 ;
        RECT 22.485000 3.455000 22.775000 3.500000 ;
        RECT 22.485000 3.640000 22.775000 3.685000 ;
        RECT 29.205000 1.755000 29.495000 1.800000 ;
        RECT 29.205000 1.940000 29.495000 1.985000 ;
        RECT 29.205000 3.455000 29.495000 3.500000 ;
        RECT 29.205000 3.640000 29.495000 3.685000 ;
        RECT 30.145000 1.755000 30.435000 1.800000 ;
        RECT 30.145000 1.940000 30.435000 1.985000 ;
        RECT 30.145000 3.455000 30.435000 3.500000 ;
        RECT 30.145000 3.640000 30.435000 3.685000 ;
        RECT 34.885000 1.755000 35.175000 1.800000 ;
        RECT 34.885000 1.940000 35.175000 1.985000 ;
        RECT 34.885000 3.455000 35.175000 3.500000 ;
        RECT 34.885000 3.640000 35.175000 3.685000 ;
        RECT 35.825000 1.755000 36.115000 1.800000 ;
        RECT 35.825000 1.940000 36.115000 1.985000 ;
        RECT 35.825000 3.455000 36.115000 3.500000 ;
        RECT 35.825000 3.640000 36.115000 3.685000 ;
        RECT 42.085000 1.755000 42.375000 1.800000 ;
        RECT 42.085000 1.940000 42.375000 1.985000 ;
        RECT 42.085000 3.455000 42.375000 3.500000 ;
        RECT 42.085000 3.640000 42.375000 3.685000 ;
        RECT 43.025000 1.755000 43.315000 1.800000 ;
        RECT 43.025000 1.940000 43.315000 1.985000 ;
        RECT 43.025000 3.455000 43.315000 3.500000 ;
        RECT 43.025000 3.640000 43.315000 3.685000 ;
        RECT 47.765000 1.755000 48.055000 1.800000 ;
        RECT 47.765000 1.940000 48.055000 1.985000 ;
        RECT 47.765000 3.455000 48.055000 3.500000 ;
        RECT 47.765000 3.640000 48.055000 3.685000 ;
        RECT 48.705000 1.755000 48.995000 1.800000 ;
        RECT 48.705000 1.940000 48.995000 1.985000 ;
        RECT 48.705000 3.455000 48.995000 3.500000 ;
        RECT 48.705000 3.640000 48.995000 3.685000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 51.980000 0.085000 ;
        RECT  0.145000  0.085000  0.395000 0.885000 ;
        RECT  1.065000  0.085000  1.335000 0.545000 ;
        RECT  2.005000  0.085000  2.255000 0.545000 ;
        RECT  4.960000  0.085000  5.250000 0.610000 ;
        RECT  5.880000  0.085000  6.170000 0.610000 ;
        RECT  6.710000  0.085000  7.000000 0.610000 ;
        RECT  7.630000  0.085000  7.920000 0.610000 ;
        RECT 10.625000  0.085000 10.875000 0.545000 ;
        RECT 11.545000  0.085000 11.815000 0.545000 ;
        RECT 12.485000  0.085000 12.735000 0.885000 ;
        RECT 13.025000  0.085000 13.275000 0.885000 ;
        RECT 13.945000  0.085000 14.215000 0.545000 ;
        RECT 14.885000  0.085000 15.135000 0.545000 ;
        RECT 17.840000  0.085000 18.130000 0.610000 ;
        RECT 18.760000  0.085000 19.050000 0.610000 ;
        RECT 19.590000  0.085000 19.880000 0.610000 ;
        RECT 20.510000  0.085000 20.800000 0.610000 ;
        RECT 23.505000  0.085000 23.755000 0.545000 ;
        RECT 24.425000  0.085000 24.695000 0.545000 ;
        RECT 25.365000  0.085000 25.615000 0.885000 ;
        RECT 26.365000  0.085000 26.615000 0.885000 ;
        RECT 27.285000  0.085000 27.555000 0.545000 ;
        RECT 28.225000  0.085000 28.475000 0.545000 ;
        RECT 31.180000  0.085000 31.470000 0.610000 ;
        RECT 32.100000  0.085000 32.390000 0.610000 ;
        RECT 32.930000  0.085000 33.220000 0.610000 ;
        RECT 33.850000  0.085000 34.140000 0.610000 ;
        RECT 36.845000  0.085000 37.095000 0.545000 ;
        RECT 37.765000  0.085000 38.035000 0.545000 ;
        RECT 38.705000  0.085000 38.955000 0.885000 ;
        RECT 39.245000  0.085000 39.495000 0.885000 ;
        RECT 40.165000  0.085000 40.435000 0.545000 ;
        RECT 41.105000  0.085000 41.355000 0.545000 ;
        RECT 44.060000  0.085000 44.350000 0.610000 ;
        RECT 44.980000  0.085000 45.270000 0.610000 ;
        RECT 45.810000  0.085000 46.100000 0.610000 ;
        RECT 46.730000  0.085000 47.020000 0.610000 ;
        RECT 49.725000  0.085000 49.975000 0.545000 ;
        RECT 50.645000  0.085000 50.915000 0.545000 ;
        RECT 51.585000  0.085000 51.835000 0.885000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
        RECT 10.725000 -0.085000 10.895000 0.085000 ;
        RECT 11.185000 -0.085000 11.355000 0.085000 ;
        RECT 11.645000 -0.085000 11.815000 0.085000 ;
        RECT 12.105000 -0.085000 12.275000 0.085000 ;
        RECT 12.565000 -0.085000 12.735000 0.085000 ;
        RECT 13.025000 -0.085000 13.195000 0.085000 ;
        RECT 13.485000 -0.085000 13.655000 0.085000 ;
        RECT 13.945000 -0.085000 14.115000 0.085000 ;
        RECT 14.405000 -0.085000 14.575000 0.085000 ;
        RECT 14.865000 -0.085000 15.035000 0.085000 ;
        RECT 15.325000 -0.085000 15.495000 0.085000 ;
        RECT 15.785000 -0.085000 15.955000 0.085000 ;
        RECT 16.245000 -0.085000 16.415000 0.085000 ;
        RECT 16.705000 -0.085000 16.875000 0.085000 ;
        RECT 17.165000 -0.085000 17.335000 0.085000 ;
        RECT 17.625000 -0.085000 17.795000 0.085000 ;
        RECT 18.085000 -0.085000 18.255000 0.085000 ;
        RECT 18.545000 -0.085000 18.715000 0.085000 ;
        RECT 19.005000 -0.085000 19.175000 0.085000 ;
        RECT 19.465000 -0.085000 19.635000 0.085000 ;
        RECT 19.925000 -0.085000 20.095000 0.085000 ;
        RECT 20.385000 -0.085000 20.555000 0.085000 ;
        RECT 20.845000 -0.085000 21.015000 0.085000 ;
        RECT 21.305000 -0.085000 21.475000 0.085000 ;
        RECT 21.765000 -0.085000 21.935000 0.085000 ;
        RECT 22.225000 -0.085000 22.395000 0.085000 ;
        RECT 22.685000 -0.085000 22.855000 0.085000 ;
        RECT 23.145000 -0.085000 23.315000 0.085000 ;
        RECT 23.605000 -0.085000 23.775000 0.085000 ;
        RECT 24.065000 -0.085000 24.235000 0.085000 ;
        RECT 24.525000 -0.085000 24.695000 0.085000 ;
        RECT 24.985000 -0.085000 25.155000 0.085000 ;
        RECT 25.445000 -0.085000 25.615000 0.085000 ;
        RECT 25.905000 -0.085000 26.075000 0.085000 ;
        RECT 26.365000 -0.085000 26.535000 0.085000 ;
        RECT 26.825000 -0.085000 26.995000 0.085000 ;
        RECT 27.285000 -0.085000 27.455000 0.085000 ;
        RECT 27.745000 -0.085000 27.915000 0.085000 ;
        RECT 28.205000 -0.085000 28.375000 0.085000 ;
        RECT 28.665000 -0.085000 28.835000 0.085000 ;
        RECT 29.125000 -0.085000 29.295000 0.085000 ;
        RECT 29.585000 -0.085000 29.755000 0.085000 ;
        RECT 30.045000 -0.085000 30.215000 0.085000 ;
        RECT 30.505000 -0.085000 30.675000 0.085000 ;
        RECT 30.965000 -0.085000 31.135000 0.085000 ;
        RECT 31.425000 -0.085000 31.595000 0.085000 ;
        RECT 31.885000 -0.085000 32.055000 0.085000 ;
        RECT 32.345000 -0.085000 32.515000 0.085000 ;
        RECT 32.805000 -0.085000 32.975000 0.085000 ;
        RECT 33.265000 -0.085000 33.435000 0.085000 ;
        RECT 33.725000 -0.085000 33.895000 0.085000 ;
        RECT 34.185000 -0.085000 34.355000 0.085000 ;
        RECT 34.645000 -0.085000 34.815000 0.085000 ;
        RECT 35.105000 -0.085000 35.275000 0.085000 ;
        RECT 35.565000 -0.085000 35.735000 0.085000 ;
        RECT 36.025000 -0.085000 36.195000 0.085000 ;
        RECT 36.485000 -0.085000 36.655000 0.085000 ;
        RECT 36.945000 -0.085000 37.115000 0.085000 ;
        RECT 37.405000 -0.085000 37.575000 0.085000 ;
        RECT 37.865000 -0.085000 38.035000 0.085000 ;
        RECT 38.325000 -0.085000 38.495000 0.085000 ;
        RECT 38.785000 -0.085000 38.955000 0.085000 ;
        RECT 39.245000 -0.085000 39.415000 0.085000 ;
        RECT 39.705000 -0.085000 39.875000 0.085000 ;
        RECT 40.165000 -0.085000 40.335000 0.085000 ;
        RECT 40.625000 -0.085000 40.795000 0.085000 ;
        RECT 41.085000 -0.085000 41.255000 0.085000 ;
        RECT 41.545000 -0.085000 41.715000 0.085000 ;
        RECT 42.005000 -0.085000 42.175000 0.085000 ;
        RECT 42.465000 -0.085000 42.635000 0.085000 ;
        RECT 42.925000 -0.085000 43.095000 0.085000 ;
        RECT 43.385000 -0.085000 43.555000 0.085000 ;
        RECT 43.845000 -0.085000 44.015000 0.085000 ;
        RECT 44.305000 -0.085000 44.475000 0.085000 ;
        RECT 44.765000 -0.085000 44.935000 0.085000 ;
        RECT 45.225000 -0.085000 45.395000 0.085000 ;
        RECT 45.685000 -0.085000 45.855000 0.085000 ;
        RECT 46.145000 -0.085000 46.315000 0.085000 ;
        RECT 46.605000 -0.085000 46.775000 0.085000 ;
        RECT 47.065000 -0.085000 47.235000 0.085000 ;
        RECT 47.525000 -0.085000 47.695000 0.085000 ;
        RECT 47.985000 -0.085000 48.155000 0.085000 ;
        RECT 48.445000 -0.085000 48.615000 0.085000 ;
        RECT 48.905000 -0.085000 49.075000 0.085000 ;
        RECT 49.365000 -0.085000 49.535000 0.085000 ;
        RECT 49.825000 -0.085000 49.995000 0.085000 ;
        RECT 50.285000 -0.085000 50.455000 0.085000 ;
        RECT 50.745000 -0.085000 50.915000 0.085000 ;
        RECT 51.205000 -0.085000 51.375000 0.085000 ;
        RECT 51.665000 -0.085000 51.835000 0.085000 ;
    END
    PORT
      LAYER li1 ;
        RECT  0.000000 5.355000 51.980000 5.525000 ;
        RECT  0.145000 4.555000  0.395000 5.355000 ;
        RECT  1.065000 4.895000  1.335000 5.355000 ;
        RECT  2.005000 4.895000  2.255000 5.355000 ;
        RECT  4.960000 4.830000  5.250000 5.355000 ;
        RECT  5.880000 4.830000  6.170000 5.355000 ;
        RECT  6.710000 4.830000  7.000000 5.355000 ;
        RECT  7.630000 4.830000  7.920000 5.355000 ;
        RECT 10.625000 4.895000 10.875000 5.355000 ;
        RECT 11.545000 4.895000 11.815000 5.355000 ;
        RECT 12.485000 4.555000 12.735000 5.355000 ;
        RECT 13.025000 4.555000 13.275000 5.355000 ;
        RECT 13.945000 4.895000 14.215000 5.355000 ;
        RECT 14.885000 4.895000 15.135000 5.355000 ;
        RECT 17.840000 4.830000 18.130000 5.355000 ;
        RECT 18.760000 4.830000 19.050000 5.355000 ;
        RECT 19.590000 4.830000 19.880000 5.355000 ;
        RECT 20.510000 4.830000 20.800000 5.355000 ;
        RECT 23.505000 4.895000 23.755000 5.355000 ;
        RECT 24.425000 4.895000 24.695000 5.355000 ;
        RECT 25.365000 4.555000 25.615000 5.355000 ;
        RECT 26.365000 4.555000 26.615000 5.355000 ;
        RECT 27.285000 4.895000 27.555000 5.355000 ;
        RECT 28.225000 4.895000 28.475000 5.355000 ;
        RECT 31.180000 4.830000 31.470000 5.355000 ;
        RECT 32.100000 4.830000 32.390000 5.355000 ;
        RECT 32.930000 4.830000 33.220000 5.355000 ;
        RECT 33.850000 4.830000 34.140000 5.355000 ;
        RECT 36.845000 4.895000 37.095000 5.355000 ;
        RECT 37.765000 4.895000 38.035000 5.355000 ;
        RECT 38.705000 4.555000 38.955000 5.355000 ;
        RECT 39.245000 4.555000 39.495000 5.355000 ;
        RECT 40.165000 4.895000 40.435000 5.355000 ;
        RECT 41.105000 4.895000 41.355000 5.355000 ;
        RECT 44.060000 4.830000 44.350000 5.355000 ;
        RECT 44.980000 4.830000 45.270000 5.355000 ;
        RECT 45.810000 4.830000 46.100000 5.355000 ;
        RECT 46.730000 4.830000 47.020000 5.355000 ;
        RECT 49.725000 4.895000 49.975000 5.355000 ;
        RECT 50.645000 4.895000 50.915000 5.355000 ;
        RECT 51.585000 4.555000 51.835000 5.355000 ;
      LAYER mcon ;
        RECT  0.145000 5.355000  0.315000 5.525000 ;
        RECT  0.605000 5.355000  0.775000 5.525000 ;
        RECT  1.065000 5.355000  1.235000 5.525000 ;
        RECT  1.525000 5.355000  1.695000 5.525000 ;
        RECT  1.985000 5.355000  2.155000 5.525000 ;
        RECT  2.445000 5.355000  2.615000 5.525000 ;
        RECT  2.905000 5.355000  3.075000 5.525000 ;
        RECT  3.365000 5.355000  3.535000 5.525000 ;
        RECT  3.825000 5.355000  3.995000 5.525000 ;
        RECT  4.285000 5.355000  4.455000 5.525000 ;
        RECT  4.745000 5.355000  4.915000 5.525000 ;
        RECT  5.205000 5.355000  5.375000 5.525000 ;
        RECT  5.665000 5.355000  5.835000 5.525000 ;
        RECT  6.125000 5.355000  6.295000 5.525000 ;
        RECT  6.585000 5.355000  6.755000 5.525000 ;
        RECT  7.045000 5.355000  7.215000 5.525000 ;
        RECT  7.505000 5.355000  7.675000 5.525000 ;
        RECT  7.965000 5.355000  8.135000 5.525000 ;
        RECT  8.425000 5.355000  8.595000 5.525000 ;
        RECT  8.885000 5.355000  9.055000 5.525000 ;
        RECT  9.345000 5.355000  9.515000 5.525000 ;
        RECT  9.805000 5.355000  9.975000 5.525000 ;
        RECT 10.265000 5.355000 10.435000 5.525000 ;
        RECT 10.725000 5.355000 10.895000 5.525000 ;
        RECT 11.185000 5.355000 11.355000 5.525000 ;
        RECT 11.645000 5.355000 11.815000 5.525000 ;
        RECT 12.105000 5.355000 12.275000 5.525000 ;
        RECT 12.565000 5.355000 12.735000 5.525000 ;
        RECT 13.025000 5.355000 13.195000 5.525000 ;
        RECT 13.485000 5.355000 13.655000 5.525000 ;
        RECT 13.945000 5.355000 14.115000 5.525000 ;
        RECT 14.405000 5.355000 14.575000 5.525000 ;
        RECT 14.865000 5.355000 15.035000 5.525000 ;
        RECT 15.325000 5.355000 15.495000 5.525000 ;
        RECT 15.785000 5.355000 15.955000 5.525000 ;
        RECT 16.245000 5.355000 16.415000 5.525000 ;
        RECT 16.705000 5.355000 16.875000 5.525000 ;
        RECT 17.165000 5.355000 17.335000 5.525000 ;
        RECT 17.625000 5.355000 17.795000 5.525000 ;
        RECT 18.085000 5.355000 18.255000 5.525000 ;
        RECT 18.545000 5.355000 18.715000 5.525000 ;
        RECT 19.005000 5.355000 19.175000 5.525000 ;
        RECT 19.465000 5.355000 19.635000 5.525000 ;
        RECT 19.925000 5.355000 20.095000 5.525000 ;
        RECT 20.385000 5.355000 20.555000 5.525000 ;
        RECT 20.845000 5.355000 21.015000 5.525000 ;
        RECT 21.305000 5.355000 21.475000 5.525000 ;
        RECT 21.765000 5.355000 21.935000 5.525000 ;
        RECT 22.225000 5.355000 22.395000 5.525000 ;
        RECT 22.685000 5.355000 22.855000 5.525000 ;
        RECT 23.145000 5.355000 23.315000 5.525000 ;
        RECT 23.605000 5.355000 23.775000 5.525000 ;
        RECT 24.065000 5.355000 24.235000 5.525000 ;
        RECT 24.525000 5.355000 24.695000 5.525000 ;
        RECT 24.985000 5.355000 25.155000 5.525000 ;
        RECT 25.445000 5.355000 25.615000 5.525000 ;
        RECT 25.905000 5.355000 26.075000 5.525000 ;
        RECT 26.365000 5.355000 26.535000 5.525000 ;
        RECT 26.825000 5.355000 26.995000 5.525000 ;
        RECT 27.285000 5.355000 27.455000 5.525000 ;
        RECT 27.745000 5.355000 27.915000 5.525000 ;
        RECT 28.205000 5.355000 28.375000 5.525000 ;
        RECT 28.665000 5.355000 28.835000 5.525000 ;
        RECT 29.125000 5.355000 29.295000 5.525000 ;
        RECT 29.585000 5.355000 29.755000 5.525000 ;
        RECT 30.045000 5.355000 30.215000 5.525000 ;
        RECT 30.505000 5.355000 30.675000 5.525000 ;
        RECT 30.965000 5.355000 31.135000 5.525000 ;
        RECT 31.425000 5.355000 31.595000 5.525000 ;
        RECT 31.885000 5.355000 32.055000 5.525000 ;
        RECT 32.345000 5.355000 32.515000 5.525000 ;
        RECT 32.805000 5.355000 32.975000 5.525000 ;
        RECT 33.265000 5.355000 33.435000 5.525000 ;
        RECT 33.725000 5.355000 33.895000 5.525000 ;
        RECT 34.185000 5.355000 34.355000 5.525000 ;
        RECT 34.645000 5.355000 34.815000 5.525000 ;
        RECT 35.105000 5.355000 35.275000 5.525000 ;
        RECT 35.565000 5.355000 35.735000 5.525000 ;
        RECT 36.025000 5.355000 36.195000 5.525000 ;
        RECT 36.485000 5.355000 36.655000 5.525000 ;
        RECT 36.945000 5.355000 37.115000 5.525000 ;
        RECT 37.405000 5.355000 37.575000 5.525000 ;
        RECT 37.865000 5.355000 38.035000 5.525000 ;
        RECT 38.325000 5.355000 38.495000 5.525000 ;
        RECT 38.785000 5.355000 38.955000 5.525000 ;
        RECT 39.245000 5.355000 39.415000 5.525000 ;
        RECT 39.705000 5.355000 39.875000 5.525000 ;
        RECT 40.165000 5.355000 40.335000 5.525000 ;
        RECT 40.625000 5.355000 40.795000 5.525000 ;
        RECT 41.085000 5.355000 41.255000 5.525000 ;
        RECT 41.545000 5.355000 41.715000 5.525000 ;
        RECT 42.005000 5.355000 42.175000 5.525000 ;
        RECT 42.465000 5.355000 42.635000 5.525000 ;
        RECT 42.925000 5.355000 43.095000 5.525000 ;
        RECT 43.385000 5.355000 43.555000 5.525000 ;
        RECT 43.845000 5.355000 44.015000 5.525000 ;
        RECT 44.305000 5.355000 44.475000 5.525000 ;
        RECT 44.765000 5.355000 44.935000 5.525000 ;
        RECT 45.225000 5.355000 45.395000 5.525000 ;
        RECT 45.685000 5.355000 45.855000 5.525000 ;
        RECT 46.145000 5.355000 46.315000 5.525000 ;
        RECT 46.605000 5.355000 46.775000 5.525000 ;
        RECT 47.065000 5.355000 47.235000 5.525000 ;
        RECT 47.525000 5.355000 47.695000 5.525000 ;
        RECT 47.985000 5.355000 48.155000 5.525000 ;
        RECT 48.445000 5.355000 48.615000 5.525000 ;
        RECT 48.905000 5.355000 49.075000 5.525000 ;
        RECT 49.365000 5.355000 49.535000 5.525000 ;
        RECT 49.825000 5.355000 49.995000 5.525000 ;
        RECT 50.285000 5.355000 50.455000 5.525000 ;
        RECT 50.745000 5.355000 50.915000 5.525000 ;
        RECT 51.205000 5.355000 51.375000 5.525000 ;
        RECT 51.665000 5.355000 51.835000 5.525000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 51.980000 0.240000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 51.980000 5.680000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 2.795000 2.805000 ;
        RECT 0.125000 1.495000 0.395000 2.635000 ;
        RECT 0.125000 2.805000 0.395000 3.945000 ;
        RECT 1.065000 1.835000 1.335000 2.635000 ;
        RECT 1.065000 2.805000 1.335000 3.605000 ;
        RECT 2.005000 1.835000 2.275000 2.635000 ;
        RECT 2.005000 2.805000 2.275000 3.605000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
    END
    PORT
      LAYER li1 ;
        RECT 10.085000 2.635000 15.675000 2.805000 ;
        RECT 10.605000 1.835000 10.875000 2.635000 ;
        RECT 10.605000 2.805000 10.875000 3.605000 ;
        RECT 11.545000 1.835000 11.815000 2.635000 ;
        RECT 11.545000 2.805000 11.815000 3.605000 ;
        RECT 12.485000 1.495000 12.755000 2.635000 ;
        RECT 12.485000 2.805000 12.755000 3.945000 ;
        RECT 13.005000 1.495000 13.275000 2.635000 ;
        RECT 13.005000 2.805000 13.275000 3.945000 ;
        RECT 13.945000 1.835000 14.215000 2.635000 ;
        RECT 13.945000 2.805000 14.215000 3.605000 ;
        RECT 14.885000 1.835000 15.155000 2.635000 ;
        RECT 14.885000 2.805000 15.155000 3.605000 ;
      LAYER mcon ;
        RECT 10.265000 2.635000 10.435000 2.805000 ;
        RECT 10.725000 2.635000 10.895000 2.805000 ;
        RECT 11.185000 2.635000 11.355000 2.805000 ;
        RECT 11.645000 2.635000 11.815000 2.805000 ;
        RECT 12.105000 2.635000 12.275000 2.805000 ;
        RECT 12.565000 2.635000 12.735000 2.805000 ;
        RECT 13.025000 2.635000 13.195000 2.805000 ;
        RECT 13.485000 2.635000 13.655000 2.805000 ;
        RECT 13.945000 2.635000 14.115000 2.805000 ;
        RECT 14.405000 2.635000 14.575000 2.805000 ;
        RECT 14.865000 2.635000 15.035000 2.805000 ;
        RECT 15.325000 2.635000 15.495000 2.805000 ;
    END
    PORT
      LAYER li1 ;
        RECT 22.965000 2.635000 29.015000 2.805000 ;
        RECT 23.485000 1.835000 23.755000 2.635000 ;
        RECT 23.485000 2.805000 23.755000 3.605000 ;
        RECT 24.425000 1.835000 24.695000 2.635000 ;
        RECT 24.425000 2.805000 24.695000 3.605000 ;
        RECT 25.365000 1.495000 25.635000 2.635000 ;
        RECT 25.365000 2.805000 25.635000 3.945000 ;
        RECT 26.345000 1.495000 26.615000 2.635000 ;
        RECT 26.345000 2.805000 26.615000 3.945000 ;
        RECT 27.285000 1.835000 27.555000 2.635000 ;
        RECT 27.285000 2.805000 27.555000 3.605000 ;
        RECT 28.225000 1.835000 28.495000 2.635000 ;
        RECT 28.225000 2.805000 28.495000 3.605000 ;
      LAYER mcon ;
        RECT 23.145000 2.635000 23.315000 2.805000 ;
        RECT 23.605000 2.635000 23.775000 2.805000 ;
        RECT 24.065000 2.635000 24.235000 2.805000 ;
        RECT 24.525000 2.635000 24.695000 2.805000 ;
        RECT 24.985000 2.635000 25.155000 2.805000 ;
        RECT 25.445000 2.635000 25.615000 2.805000 ;
        RECT 25.905000 2.635000 26.075000 2.805000 ;
        RECT 26.365000 2.635000 26.535000 2.805000 ;
        RECT 26.825000 2.635000 26.995000 2.805000 ;
        RECT 27.285000 2.635000 27.455000 2.805000 ;
        RECT 27.745000 2.635000 27.915000 2.805000 ;
        RECT 28.205000 2.635000 28.375000 2.805000 ;
        RECT 28.665000 2.635000 28.835000 2.805000 ;
    END
    PORT
      LAYER li1 ;
        RECT 36.305000 2.635000 41.895000 2.805000 ;
        RECT 36.825000 1.835000 37.095000 2.635000 ;
        RECT 36.825000 2.805000 37.095000 3.605000 ;
        RECT 37.765000 1.835000 38.035000 2.635000 ;
        RECT 37.765000 2.805000 38.035000 3.605000 ;
        RECT 38.705000 1.495000 38.975000 2.635000 ;
        RECT 38.705000 2.805000 38.975000 3.945000 ;
        RECT 39.225000 1.495000 39.495000 2.635000 ;
        RECT 39.225000 2.805000 39.495000 3.945000 ;
        RECT 40.165000 1.835000 40.435000 2.635000 ;
        RECT 40.165000 2.805000 40.435000 3.605000 ;
        RECT 41.105000 1.835000 41.375000 2.635000 ;
        RECT 41.105000 2.805000 41.375000 3.605000 ;
      LAYER mcon ;
        RECT 36.485000 2.635000 36.655000 2.805000 ;
        RECT 36.945000 2.635000 37.115000 2.805000 ;
        RECT 37.405000 2.635000 37.575000 2.805000 ;
        RECT 37.865000 2.635000 38.035000 2.805000 ;
        RECT 38.325000 2.635000 38.495000 2.805000 ;
        RECT 38.785000 2.635000 38.955000 2.805000 ;
        RECT 39.245000 2.635000 39.415000 2.805000 ;
        RECT 39.705000 2.635000 39.875000 2.805000 ;
        RECT 40.165000 2.635000 40.335000 2.805000 ;
        RECT 40.625000 2.635000 40.795000 2.805000 ;
        RECT 41.085000 2.635000 41.255000 2.805000 ;
        RECT 41.545000 2.635000 41.715000 2.805000 ;
    END
    PORT
      LAYER li1 ;
        RECT 49.185000 2.635000 51.980000 2.805000 ;
        RECT 49.705000 1.835000 49.975000 2.635000 ;
        RECT 49.705000 2.805000 49.975000 3.605000 ;
        RECT 50.645000 1.835000 50.915000 2.635000 ;
        RECT 50.645000 2.805000 50.915000 3.605000 ;
        RECT 51.585000 1.495000 51.855000 2.635000 ;
        RECT 51.585000 2.805000 51.855000 3.945000 ;
      LAYER mcon ;
        RECT 49.365000 2.635000 49.535000 2.805000 ;
        RECT 49.825000 2.635000 49.995000 2.805000 ;
        RECT 50.285000 2.635000 50.455000 2.805000 ;
        RECT 50.745000 2.635000 50.915000 2.805000 ;
        RECT 51.205000 2.635000 51.375000 2.805000 ;
        RECT 51.665000 2.635000 51.835000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 51.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.565000 0.255000  0.895000 0.715000 ;
      RECT  0.565000 0.715000  2.695000 0.885000 ;
      RECT  0.565000 1.495000  2.795000 1.665000 ;
      RECT  0.565000 1.665000  0.895000 2.465000 ;
      RECT  0.565000 2.975000  0.895000 3.775000 ;
      RECT  0.565000 3.775000  2.795000 3.945000 ;
      RECT  0.565000 4.555000  2.695000 4.725000 ;
      RECT  0.565000 4.725000  0.895000 5.185000 ;
      RECT  1.505000 0.255000  1.835000 0.715000 ;
      RECT  1.505000 1.665000  1.835000 2.465000 ;
      RECT  1.505000 2.975000  1.835000 3.775000 ;
      RECT  1.505000 4.725000  1.835000 5.185000 ;
      RECT  2.425000 0.255000  4.455000 0.425000 ;
      RECT  2.425000 0.425000  2.695000 0.715000 ;
      RECT  2.425000 4.725000  2.695000 5.015000 ;
      RECT  2.425000 5.015000  4.455000 5.185000 ;
      RECT  2.495000 1.665000  2.795000 2.465000 ;
      RECT  2.495000 2.975000  2.795000 3.775000 ;
      RECT  3.365000 0.425000  3.535000 0.770000 ;
      RECT  3.365000 4.670000  3.535000 5.015000 ;
      RECT  3.465000 1.535000  3.735000 2.465000 ;
      RECT  3.465000 2.975000  3.735000 3.905000 ;
      RECT  4.205000 0.425000  4.455000 0.770000 ;
      RECT  4.205000 4.670000  4.455000 5.015000 ;
      RECT  4.405000 1.065000  5.590000 1.395000 ;
      RECT  4.405000 1.565000  4.705000 2.465000 ;
      RECT  4.405000 2.635000  8.475000 2.805000 ;
      RECT  4.405000 2.975000  4.705000 3.875000 ;
      RECT  4.405000 4.045000  5.590000 4.375000 ;
      RECT  4.950000 1.605000  5.225000 2.635000 ;
      RECT  4.950000 2.805000  5.225000 3.835000 ;
      RECT  5.420000 0.280000  5.670000 0.825000 ;
      RECT  5.420000 0.825000  5.590000 1.065000 ;
      RECT  5.420000 1.395000  5.590000 1.605000 ;
      RECT  5.420000 1.605000  5.750000 2.465000 ;
      RECT  5.420000 2.975000  5.750000 3.835000 ;
      RECT  5.420000 3.835000  5.590000 4.045000 ;
      RECT  5.420000 4.375000  5.590000 4.615000 ;
      RECT  5.420000 4.615000  5.670000 5.160000 ;
      RECT  5.920000 1.605000  6.220000 2.635000 ;
      RECT  5.920000 2.805000  6.220000 3.835000 ;
      RECT  6.660000 1.605000  6.960000 2.635000 ;
      RECT  6.660000 2.805000  6.960000 3.835000 ;
      RECT  7.130000 1.605000  7.460000 2.465000 ;
      RECT  7.130000 2.975000  7.460000 3.835000 ;
      RECT  7.210000 0.280000  7.460000 0.825000 ;
      RECT  7.210000 4.615000  7.460000 5.160000 ;
      RECT  7.290000 0.825000  7.460000 1.065000 ;
      RECT  7.290000 1.065000  8.475000 1.395000 ;
      RECT  7.290000 1.395000  7.460000 1.605000 ;
      RECT  7.290000 3.835000  7.460000 4.045000 ;
      RECT  7.290000 4.045000  8.475000 4.375000 ;
      RECT  7.290000 4.375000  7.460000 4.615000 ;
      RECT  7.655000 1.605000  7.930000 2.635000 ;
      RECT  7.655000 2.805000  7.930000 3.835000 ;
      RECT  8.175000 1.565000  8.475000 2.465000 ;
      RECT  8.175000 2.975000  8.475000 3.875000 ;
      RECT  8.425000 0.255000 10.455000 0.425000 ;
      RECT  8.425000 0.425000  8.675000 0.770000 ;
      RECT  8.425000 4.670000  8.675000 5.015000 ;
      RECT  8.425000 5.015000 10.455000 5.185000 ;
      RECT  8.645000 1.065000  9.915000 1.365000 ;
      RECT  8.645000 1.365000  8.975000 4.075000 ;
      RECT  8.645000 4.075000  9.915000 4.375000 ;
      RECT  8.845000 0.595000  9.175000 1.065000 ;
      RECT  8.845000 4.375000  9.175000 4.845000 ;
      RECT  9.145000 1.535000  9.415000 2.465000 ;
      RECT  9.145000 2.975000  9.415000 3.905000 ;
      RECT  9.345000 0.425000  9.515000 0.770000 ;
      RECT  9.345000 4.670000  9.515000 5.015000 ;
      RECT  9.585000 1.365000  9.915000 4.075000 ;
      RECT  9.685000 0.595000 10.015000 0.885000 ;
      RECT  9.685000 0.885000  9.915000 1.065000 ;
      RECT  9.685000 4.375000  9.915000 4.555000 ;
      RECT  9.685000 4.555000 10.015000 4.845000 ;
      RECT 10.085000 1.495000 12.315000 1.665000 ;
      RECT 10.085000 1.665000 10.385000 2.465000 ;
      RECT 10.085000 2.975000 10.385000 3.775000 ;
      RECT 10.085000 3.775000 12.315000 3.945000 ;
      RECT 10.185000 0.425000 10.455000 0.715000 ;
      RECT 10.185000 0.715000 12.315000 0.885000 ;
      RECT 10.185000 4.555000 12.315000 4.725000 ;
      RECT 10.185000 4.725000 10.455000 5.015000 ;
      RECT 11.045000 0.255000 11.375000 0.715000 ;
      RECT 11.045000 1.665000 11.375000 2.465000 ;
      RECT 11.045000 2.975000 11.375000 3.775000 ;
      RECT 11.045000 4.725000 11.375000 5.185000 ;
      RECT 11.985000 0.255000 12.315000 0.715000 ;
      RECT 11.985000 1.665000 12.315000 2.465000 ;
      RECT 11.985000 2.975000 12.315000 3.775000 ;
      RECT 11.985000 4.725000 12.315000 5.185000 ;
      RECT 13.445000 0.255000 13.775000 0.715000 ;
      RECT 13.445000 0.715000 15.575000 0.885000 ;
      RECT 13.445000 1.495000 15.675000 1.665000 ;
      RECT 13.445000 1.665000 13.775000 2.465000 ;
      RECT 13.445000 2.975000 13.775000 3.775000 ;
      RECT 13.445000 3.775000 15.675000 3.945000 ;
      RECT 13.445000 4.555000 15.575000 4.725000 ;
      RECT 13.445000 4.725000 13.775000 5.185000 ;
      RECT 14.385000 0.255000 14.715000 0.715000 ;
      RECT 14.385000 1.665000 14.715000 2.465000 ;
      RECT 14.385000 2.975000 14.715000 3.775000 ;
      RECT 14.385000 4.725000 14.715000 5.185000 ;
      RECT 15.305000 0.255000 17.335000 0.425000 ;
      RECT 15.305000 0.425000 15.575000 0.715000 ;
      RECT 15.305000 4.725000 15.575000 5.015000 ;
      RECT 15.305000 5.015000 17.335000 5.185000 ;
      RECT 15.375000 1.665000 15.675000 2.465000 ;
      RECT 15.375000 2.975000 15.675000 3.775000 ;
      RECT 15.745000 0.595000 16.075000 0.885000 ;
      RECT 15.745000 4.555000 16.075000 4.845000 ;
      RECT 15.845000 0.885000 16.075000 1.065000 ;
      RECT 15.845000 1.065000 17.115000 1.365000 ;
      RECT 15.845000 1.365000 16.175000 4.075000 ;
      RECT 15.845000 4.075000 17.115000 4.375000 ;
      RECT 15.845000 4.375000 16.075000 4.555000 ;
      RECT 16.245000 0.425000 16.415000 0.770000 ;
      RECT 16.245000 4.670000 16.415000 5.015000 ;
      RECT 16.345000 1.535000 16.615000 2.465000 ;
      RECT 16.345000 2.975000 16.615000 3.905000 ;
      RECT 16.585000 0.595000 16.915000 1.065000 ;
      RECT 16.585000 4.375000 16.915000 4.845000 ;
      RECT 16.785000 1.365000 17.115000 4.075000 ;
      RECT 17.085000 0.425000 17.335000 0.770000 ;
      RECT 17.085000 4.670000 17.335000 5.015000 ;
      RECT 17.285000 1.065000 18.470000 1.395000 ;
      RECT 17.285000 1.565000 17.585000 2.465000 ;
      RECT 17.285000 2.635000 21.355000 2.805000 ;
      RECT 17.285000 2.975000 17.585000 3.875000 ;
      RECT 17.285000 4.045000 18.470000 4.375000 ;
      RECT 17.830000 1.605000 18.105000 2.635000 ;
      RECT 17.830000 2.805000 18.105000 3.835000 ;
      RECT 18.300000 0.280000 18.550000 0.825000 ;
      RECT 18.300000 0.825000 18.470000 1.065000 ;
      RECT 18.300000 1.395000 18.470000 1.605000 ;
      RECT 18.300000 1.605000 18.630000 2.465000 ;
      RECT 18.300000 2.975000 18.630000 3.835000 ;
      RECT 18.300000 3.835000 18.470000 4.045000 ;
      RECT 18.300000 4.375000 18.470000 4.615000 ;
      RECT 18.300000 4.615000 18.550000 5.160000 ;
      RECT 18.800000 1.605000 19.100000 2.635000 ;
      RECT 18.800000 2.805000 19.100000 3.835000 ;
      RECT 19.540000 1.605000 19.840000 2.635000 ;
      RECT 19.540000 2.805000 19.840000 3.835000 ;
      RECT 20.010000 1.605000 20.340000 2.465000 ;
      RECT 20.010000 2.975000 20.340000 3.835000 ;
      RECT 20.090000 0.280000 20.340000 0.825000 ;
      RECT 20.090000 4.615000 20.340000 5.160000 ;
      RECT 20.170000 0.825000 20.340000 1.065000 ;
      RECT 20.170000 1.065000 21.355000 1.395000 ;
      RECT 20.170000 1.395000 20.340000 1.605000 ;
      RECT 20.170000 3.835000 20.340000 4.045000 ;
      RECT 20.170000 4.045000 21.355000 4.375000 ;
      RECT 20.170000 4.375000 20.340000 4.615000 ;
      RECT 20.535000 1.605000 20.810000 2.635000 ;
      RECT 20.535000 2.805000 20.810000 3.835000 ;
      RECT 21.055000 1.565000 21.355000 2.465000 ;
      RECT 21.055000 2.975000 21.355000 3.875000 ;
      RECT 21.305000 0.255000 23.335000 0.425000 ;
      RECT 21.305000 0.425000 21.555000 0.770000 ;
      RECT 21.305000 4.670000 21.555000 5.015000 ;
      RECT 21.305000 5.015000 23.335000 5.185000 ;
      RECT 21.525000 1.065000 22.795000 1.365000 ;
      RECT 21.525000 1.365000 21.855000 4.075000 ;
      RECT 21.525000 4.075000 22.795000 4.375000 ;
      RECT 21.725000 0.595000 22.055000 1.065000 ;
      RECT 21.725000 4.375000 22.055000 4.845000 ;
      RECT 22.025000 1.535000 22.295000 2.465000 ;
      RECT 22.025000 2.975000 22.295000 3.905000 ;
      RECT 22.225000 0.425000 22.395000 0.770000 ;
      RECT 22.225000 4.670000 22.395000 5.015000 ;
      RECT 22.465000 1.365000 22.795000 4.075000 ;
      RECT 22.565000 0.595000 22.895000 0.885000 ;
      RECT 22.565000 0.885000 22.795000 1.065000 ;
      RECT 22.565000 4.375000 22.795000 4.555000 ;
      RECT 22.565000 4.555000 22.895000 4.845000 ;
      RECT 22.965000 1.495000 25.195000 1.665000 ;
      RECT 22.965000 1.665000 23.265000 2.465000 ;
      RECT 22.965000 2.975000 23.265000 3.775000 ;
      RECT 22.965000 3.775000 25.195000 3.945000 ;
      RECT 23.065000 0.425000 23.335000 0.715000 ;
      RECT 23.065000 0.715000 25.195000 0.885000 ;
      RECT 23.065000 4.555000 25.195000 4.725000 ;
      RECT 23.065000 4.725000 23.335000 5.015000 ;
      RECT 23.925000 0.255000 24.255000 0.715000 ;
      RECT 23.925000 1.665000 24.255000 2.465000 ;
      RECT 23.925000 2.975000 24.255000 3.775000 ;
      RECT 23.925000 4.725000 24.255000 5.185000 ;
      RECT 24.865000 0.255000 25.195000 0.715000 ;
      RECT 24.865000 1.665000 25.195000 2.465000 ;
      RECT 24.865000 2.975000 25.195000 3.775000 ;
      RECT 24.865000 4.725000 25.195000 5.185000 ;
      RECT 26.785000 0.255000 27.115000 0.715000 ;
      RECT 26.785000 0.715000 28.915000 0.885000 ;
      RECT 26.785000 1.495000 29.015000 1.665000 ;
      RECT 26.785000 1.665000 27.115000 2.465000 ;
      RECT 26.785000 2.975000 27.115000 3.775000 ;
      RECT 26.785000 3.775000 29.015000 3.945000 ;
      RECT 26.785000 4.555000 28.915000 4.725000 ;
      RECT 26.785000 4.725000 27.115000 5.185000 ;
      RECT 27.725000 0.255000 28.055000 0.715000 ;
      RECT 27.725000 1.665000 28.055000 2.465000 ;
      RECT 27.725000 2.975000 28.055000 3.775000 ;
      RECT 27.725000 4.725000 28.055000 5.185000 ;
      RECT 28.645000 0.255000 30.675000 0.425000 ;
      RECT 28.645000 0.425000 28.915000 0.715000 ;
      RECT 28.645000 4.725000 28.915000 5.015000 ;
      RECT 28.645000 5.015000 30.675000 5.185000 ;
      RECT 28.715000 1.665000 29.015000 2.465000 ;
      RECT 28.715000 2.975000 29.015000 3.775000 ;
      RECT 29.085000 0.595000 29.415000 0.885000 ;
      RECT 29.085000 4.555000 29.415000 4.845000 ;
      RECT 29.185000 0.885000 29.415000 1.065000 ;
      RECT 29.185000 1.065000 30.455000 1.365000 ;
      RECT 29.185000 1.365000 29.515000 4.075000 ;
      RECT 29.185000 4.075000 30.455000 4.375000 ;
      RECT 29.185000 4.375000 29.415000 4.555000 ;
      RECT 29.585000 0.425000 29.755000 0.770000 ;
      RECT 29.585000 4.670000 29.755000 5.015000 ;
      RECT 29.685000 1.535000 29.955000 2.465000 ;
      RECT 29.685000 2.975000 29.955000 3.905000 ;
      RECT 29.925000 0.595000 30.255000 1.065000 ;
      RECT 29.925000 4.375000 30.255000 4.845000 ;
      RECT 30.125000 1.365000 30.455000 4.075000 ;
      RECT 30.425000 0.425000 30.675000 0.770000 ;
      RECT 30.425000 4.670000 30.675000 5.015000 ;
      RECT 30.625000 1.065000 31.810000 1.395000 ;
      RECT 30.625000 1.565000 30.925000 2.465000 ;
      RECT 30.625000 2.635000 34.695000 2.805000 ;
      RECT 30.625000 2.975000 30.925000 3.875000 ;
      RECT 30.625000 4.045000 31.810000 4.375000 ;
      RECT 31.170000 1.605000 31.445000 2.635000 ;
      RECT 31.170000 2.805000 31.445000 3.835000 ;
      RECT 31.640000 0.280000 31.890000 0.825000 ;
      RECT 31.640000 0.825000 31.810000 1.065000 ;
      RECT 31.640000 1.395000 31.810000 1.605000 ;
      RECT 31.640000 1.605000 31.970000 2.465000 ;
      RECT 31.640000 2.975000 31.970000 3.835000 ;
      RECT 31.640000 3.835000 31.810000 4.045000 ;
      RECT 31.640000 4.375000 31.810000 4.615000 ;
      RECT 31.640000 4.615000 31.890000 5.160000 ;
      RECT 32.140000 1.605000 32.440000 2.635000 ;
      RECT 32.140000 2.805000 32.440000 3.835000 ;
      RECT 32.880000 1.605000 33.180000 2.635000 ;
      RECT 32.880000 2.805000 33.180000 3.835000 ;
      RECT 33.350000 1.605000 33.680000 2.465000 ;
      RECT 33.350000 2.975000 33.680000 3.835000 ;
      RECT 33.430000 0.280000 33.680000 0.825000 ;
      RECT 33.430000 4.615000 33.680000 5.160000 ;
      RECT 33.510000 0.825000 33.680000 1.065000 ;
      RECT 33.510000 1.065000 34.695000 1.395000 ;
      RECT 33.510000 1.395000 33.680000 1.605000 ;
      RECT 33.510000 3.835000 33.680000 4.045000 ;
      RECT 33.510000 4.045000 34.695000 4.375000 ;
      RECT 33.510000 4.375000 33.680000 4.615000 ;
      RECT 33.875000 1.605000 34.150000 2.635000 ;
      RECT 33.875000 2.805000 34.150000 3.835000 ;
      RECT 34.395000 1.565000 34.695000 2.465000 ;
      RECT 34.395000 2.975000 34.695000 3.875000 ;
      RECT 34.645000 0.255000 36.675000 0.425000 ;
      RECT 34.645000 0.425000 34.895000 0.770000 ;
      RECT 34.645000 4.670000 34.895000 5.015000 ;
      RECT 34.645000 5.015000 36.675000 5.185000 ;
      RECT 34.865000 1.065000 36.135000 1.365000 ;
      RECT 34.865000 1.365000 35.195000 4.075000 ;
      RECT 34.865000 4.075000 36.135000 4.375000 ;
      RECT 35.065000 0.595000 35.395000 1.065000 ;
      RECT 35.065000 4.375000 35.395000 4.845000 ;
      RECT 35.365000 1.535000 35.635000 2.465000 ;
      RECT 35.365000 2.975000 35.635000 3.905000 ;
      RECT 35.565000 0.425000 35.735000 0.770000 ;
      RECT 35.565000 4.670000 35.735000 5.015000 ;
      RECT 35.805000 1.365000 36.135000 4.075000 ;
      RECT 35.905000 0.595000 36.235000 0.885000 ;
      RECT 35.905000 0.885000 36.135000 1.065000 ;
      RECT 35.905000 4.375000 36.135000 4.555000 ;
      RECT 35.905000 4.555000 36.235000 4.845000 ;
      RECT 36.305000 1.495000 38.535000 1.665000 ;
      RECT 36.305000 1.665000 36.605000 2.465000 ;
      RECT 36.305000 2.975000 36.605000 3.775000 ;
      RECT 36.305000 3.775000 38.535000 3.945000 ;
      RECT 36.405000 0.425000 36.675000 0.715000 ;
      RECT 36.405000 0.715000 38.535000 0.885000 ;
      RECT 36.405000 4.555000 38.535000 4.725000 ;
      RECT 36.405000 4.725000 36.675000 5.015000 ;
      RECT 37.265000 0.255000 37.595000 0.715000 ;
      RECT 37.265000 1.665000 37.595000 2.465000 ;
      RECT 37.265000 2.975000 37.595000 3.775000 ;
      RECT 37.265000 4.725000 37.595000 5.185000 ;
      RECT 38.205000 0.255000 38.535000 0.715000 ;
      RECT 38.205000 1.665000 38.535000 2.465000 ;
      RECT 38.205000 2.975000 38.535000 3.775000 ;
      RECT 38.205000 4.725000 38.535000 5.185000 ;
      RECT 39.665000 0.255000 39.995000 0.715000 ;
      RECT 39.665000 0.715000 41.795000 0.885000 ;
      RECT 39.665000 1.495000 41.895000 1.665000 ;
      RECT 39.665000 1.665000 39.995000 2.465000 ;
      RECT 39.665000 2.975000 39.995000 3.775000 ;
      RECT 39.665000 3.775000 41.895000 3.945000 ;
      RECT 39.665000 4.555000 41.795000 4.725000 ;
      RECT 39.665000 4.725000 39.995000 5.185000 ;
      RECT 40.605000 0.255000 40.935000 0.715000 ;
      RECT 40.605000 1.665000 40.935000 2.465000 ;
      RECT 40.605000 2.975000 40.935000 3.775000 ;
      RECT 40.605000 4.725000 40.935000 5.185000 ;
      RECT 41.525000 0.255000 43.555000 0.425000 ;
      RECT 41.525000 0.425000 41.795000 0.715000 ;
      RECT 41.525000 4.725000 41.795000 5.015000 ;
      RECT 41.525000 5.015000 43.555000 5.185000 ;
      RECT 41.595000 1.665000 41.895000 2.465000 ;
      RECT 41.595000 2.975000 41.895000 3.775000 ;
      RECT 41.965000 0.595000 42.295000 0.885000 ;
      RECT 41.965000 4.555000 42.295000 4.845000 ;
      RECT 42.065000 0.885000 42.295000 1.065000 ;
      RECT 42.065000 1.065000 43.335000 1.365000 ;
      RECT 42.065000 1.365000 42.395000 4.075000 ;
      RECT 42.065000 4.075000 43.335000 4.375000 ;
      RECT 42.065000 4.375000 42.295000 4.555000 ;
      RECT 42.465000 0.425000 42.635000 0.770000 ;
      RECT 42.465000 4.670000 42.635000 5.015000 ;
      RECT 42.565000 1.535000 42.835000 2.465000 ;
      RECT 42.565000 2.975000 42.835000 3.905000 ;
      RECT 42.805000 0.595000 43.135000 1.065000 ;
      RECT 42.805000 4.375000 43.135000 4.845000 ;
      RECT 43.005000 1.365000 43.335000 4.075000 ;
      RECT 43.305000 0.425000 43.555000 0.770000 ;
      RECT 43.305000 4.670000 43.555000 5.015000 ;
      RECT 43.505000 1.065000 44.690000 1.395000 ;
      RECT 43.505000 1.565000 43.805000 2.465000 ;
      RECT 43.505000 2.635000 47.575000 2.805000 ;
      RECT 43.505000 2.975000 43.805000 3.875000 ;
      RECT 43.505000 4.045000 44.690000 4.375000 ;
      RECT 44.050000 1.605000 44.325000 2.635000 ;
      RECT 44.050000 2.805000 44.325000 3.835000 ;
      RECT 44.520000 0.280000 44.770000 0.825000 ;
      RECT 44.520000 0.825000 44.690000 1.065000 ;
      RECT 44.520000 1.395000 44.690000 1.605000 ;
      RECT 44.520000 1.605000 44.850000 2.465000 ;
      RECT 44.520000 2.975000 44.850000 3.835000 ;
      RECT 44.520000 3.835000 44.690000 4.045000 ;
      RECT 44.520000 4.375000 44.690000 4.615000 ;
      RECT 44.520000 4.615000 44.770000 5.160000 ;
      RECT 45.020000 1.605000 45.320000 2.635000 ;
      RECT 45.020000 2.805000 45.320000 3.835000 ;
      RECT 45.760000 1.605000 46.060000 2.635000 ;
      RECT 45.760000 2.805000 46.060000 3.835000 ;
      RECT 46.230000 1.605000 46.560000 2.465000 ;
      RECT 46.230000 2.975000 46.560000 3.835000 ;
      RECT 46.310000 0.280000 46.560000 0.825000 ;
      RECT 46.310000 4.615000 46.560000 5.160000 ;
      RECT 46.390000 0.825000 46.560000 1.065000 ;
      RECT 46.390000 1.065000 47.575000 1.395000 ;
      RECT 46.390000 1.395000 46.560000 1.605000 ;
      RECT 46.390000 3.835000 46.560000 4.045000 ;
      RECT 46.390000 4.045000 47.575000 4.375000 ;
      RECT 46.390000 4.375000 46.560000 4.615000 ;
      RECT 46.755000 1.605000 47.030000 2.635000 ;
      RECT 46.755000 2.805000 47.030000 3.835000 ;
      RECT 47.275000 1.565000 47.575000 2.465000 ;
      RECT 47.275000 2.975000 47.575000 3.875000 ;
      RECT 47.525000 0.255000 49.555000 0.425000 ;
      RECT 47.525000 0.425000 47.775000 0.770000 ;
      RECT 47.525000 4.670000 47.775000 5.015000 ;
      RECT 47.525000 5.015000 49.555000 5.185000 ;
      RECT 47.745000 1.065000 49.015000 1.365000 ;
      RECT 47.745000 1.365000 48.075000 4.075000 ;
      RECT 47.745000 4.075000 49.015000 4.375000 ;
      RECT 47.945000 0.595000 48.275000 1.065000 ;
      RECT 47.945000 4.375000 48.275000 4.845000 ;
      RECT 48.245000 1.535000 48.515000 2.465000 ;
      RECT 48.245000 2.975000 48.515000 3.905000 ;
      RECT 48.445000 0.425000 48.615000 0.770000 ;
      RECT 48.445000 4.670000 48.615000 5.015000 ;
      RECT 48.685000 1.365000 49.015000 4.075000 ;
      RECT 48.785000 0.595000 49.115000 0.885000 ;
      RECT 48.785000 0.885000 49.015000 1.065000 ;
      RECT 48.785000 4.375000 49.015000 4.555000 ;
      RECT 48.785000 4.555000 49.115000 4.845000 ;
      RECT 49.185000 1.495000 51.415000 1.665000 ;
      RECT 49.185000 1.665000 49.485000 2.465000 ;
      RECT 49.185000 2.975000 49.485000 3.775000 ;
      RECT 49.185000 3.775000 51.415000 3.945000 ;
      RECT 49.285000 0.425000 49.555000 0.715000 ;
      RECT 49.285000 0.715000 51.415000 0.885000 ;
      RECT 49.285000 4.555000 51.415000 4.725000 ;
      RECT 49.285000 4.725000 49.555000 5.015000 ;
      RECT 50.145000 0.255000 50.475000 0.715000 ;
      RECT 50.145000 1.665000 50.475000 2.465000 ;
      RECT 50.145000 2.975000 50.475000 3.775000 ;
      RECT 50.145000 4.725000 50.475000 5.185000 ;
      RECT 51.085000 0.255000 51.415000 0.715000 ;
      RECT 51.085000 1.665000 51.415000 2.465000 ;
      RECT 51.085000 2.975000 51.415000 3.775000 ;
      RECT 51.085000 4.725000 51.415000 5.185000 ;
    LAYER mcon ;
      RECT  0.645000 2.140000  0.815000 2.310000 ;
      RECT  0.645000 3.130000  0.815000 3.300000 ;
      RECT  1.585000 2.140000  1.755000 2.310000 ;
      RECT  1.585000 3.130000  1.755000 3.300000 ;
      RECT  2.565000 2.140000  2.735000 2.310000 ;
      RECT  2.565000 3.130000  2.735000 3.300000 ;
      RECT  3.515000 2.140000  3.685000 2.310000 ;
      RECT  3.515000 3.130000  3.685000 3.300000 ;
      RECT  4.465000 2.140000  4.635000 2.310000 ;
      RECT  4.465000 3.130000  4.635000 3.300000 ;
      RECT  4.745000 2.635000  4.915000 2.805000 ;
      RECT  5.205000 2.635000  5.375000 2.805000 ;
      RECT  5.665000 2.635000  5.835000 2.805000 ;
      RECT  6.125000 2.635000  6.295000 2.805000 ;
      RECT  6.585000 2.635000  6.755000 2.805000 ;
      RECT  7.045000 2.635000  7.215000 2.805000 ;
      RECT  7.505000 2.635000  7.675000 2.805000 ;
      RECT  7.965000 2.635000  8.135000 2.805000 ;
      RECT  8.245000 2.140000  8.415000 2.310000 ;
      RECT  8.245000 3.130000  8.415000 3.300000 ;
      RECT  8.725000 1.785000  8.895000 1.955000 ;
      RECT  8.725000 3.485000  8.895000 3.655000 ;
      RECT  9.195000 2.140000  9.365000 2.310000 ;
      RECT  9.195000 3.130000  9.365000 3.300000 ;
      RECT  9.665000 1.785000  9.835000 1.955000 ;
      RECT  9.665000 3.485000  9.835000 3.655000 ;
      RECT 10.145000 2.140000 10.315000 2.310000 ;
      RECT 10.145000 3.130000 10.315000 3.300000 ;
      RECT 11.125000 2.140000 11.295000 2.310000 ;
      RECT 11.125000 3.130000 11.295000 3.300000 ;
      RECT 12.065000 2.140000 12.235000 2.310000 ;
      RECT 12.065000 3.130000 12.235000 3.300000 ;
      RECT 13.525000 2.140000 13.695000 2.310000 ;
      RECT 13.525000 3.130000 13.695000 3.300000 ;
      RECT 14.465000 2.140000 14.635000 2.310000 ;
      RECT 14.465000 3.130000 14.635000 3.300000 ;
      RECT 15.445000 2.140000 15.615000 2.310000 ;
      RECT 15.445000 3.130000 15.615000 3.300000 ;
      RECT 15.925000 1.785000 16.095000 1.955000 ;
      RECT 15.925000 3.485000 16.095000 3.655000 ;
      RECT 16.395000 2.140000 16.565000 2.310000 ;
      RECT 16.395000 3.130000 16.565000 3.300000 ;
      RECT 16.865000 1.785000 17.035000 1.955000 ;
      RECT 16.865000 3.485000 17.035000 3.655000 ;
      RECT 17.345000 2.140000 17.515000 2.310000 ;
      RECT 17.345000 3.130000 17.515000 3.300000 ;
      RECT 17.625000 2.635000 17.795000 2.805000 ;
      RECT 18.085000 2.635000 18.255000 2.805000 ;
      RECT 18.545000 2.635000 18.715000 2.805000 ;
      RECT 19.005000 2.635000 19.175000 2.805000 ;
      RECT 19.465000 2.635000 19.635000 2.805000 ;
      RECT 19.925000 2.635000 20.095000 2.805000 ;
      RECT 20.385000 2.635000 20.555000 2.805000 ;
      RECT 20.845000 2.635000 21.015000 2.805000 ;
      RECT 21.125000 2.140000 21.295000 2.310000 ;
      RECT 21.125000 3.130000 21.295000 3.300000 ;
      RECT 21.605000 1.785000 21.775000 1.955000 ;
      RECT 21.605000 3.485000 21.775000 3.655000 ;
      RECT 22.075000 2.140000 22.245000 2.310000 ;
      RECT 22.075000 3.130000 22.245000 3.300000 ;
      RECT 22.545000 1.785000 22.715000 1.955000 ;
      RECT 22.545000 3.485000 22.715000 3.655000 ;
      RECT 23.025000 2.140000 23.195000 2.310000 ;
      RECT 23.025000 3.130000 23.195000 3.300000 ;
      RECT 24.005000 2.140000 24.175000 2.310000 ;
      RECT 24.005000 3.130000 24.175000 3.300000 ;
      RECT 24.945000 2.140000 25.115000 2.310000 ;
      RECT 24.945000 3.130000 25.115000 3.300000 ;
      RECT 26.865000 2.140000 27.035000 2.310000 ;
      RECT 26.865000 3.130000 27.035000 3.300000 ;
      RECT 27.805000 2.140000 27.975000 2.310000 ;
      RECT 27.805000 3.130000 27.975000 3.300000 ;
      RECT 28.785000 2.140000 28.955000 2.310000 ;
      RECT 28.785000 3.130000 28.955000 3.300000 ;
      RECT 29.265000 1.785000 29.435000 1.955000 ;
      RECT 29.265000 3.485000 29.435000 3.655000 ;
      RECT 29.735000 2.140000 29.905000 2.310000 ;
      RECT 29.735000 3.130000 29.905000 3.300000 ;
      RECT 30.205000 1.785000 30.375000 1.955000 ;
      RECT 30.205000 3.485000 30.375000 3.655000 ;
      RECT 30.685000 2.140000 30.855000 2.310000 ;
      RECT 30.685000 3.130000 30.855000 3.300000 ;
      RECT 30.965000 2.635000 31.135000 2.805000 ;
      RECT 31.425000 2.635000 31.595000 2.805000 ;
      RECT 31.885000 2.635000 32.055000 2.805000 ;
      RECT 32.345000 2.635000 32.515000 2.805000 ;
      RECT 32.805000 2.635000 32.975000 2.805000 ;
      RECT 33.265000 2.635000 33.435000 2.805000 ;
      RECT 33.725000 2.635000 33.895000 2.805000 ;
      RECT 34.185000 2.635000 34.355000 2.805000 ;
      RECT 34.465000 2.140000 34.635000 2.310000 ;
      RECT 34.465000 3.130000 34.635000 3.300000 ;
      RECT 34.945000 1.785000 35.115000 1.955000 ;
      RECT 34.945000 3.485000 35.115000 3.655000 ;
      RECT 35.415000 2.140000 35.585000 2.310000 ;
      RECT 35.415000 3.130000 35.585000 3.300000 ;
      RECT 35.885000 1.785000 36.055000 1.955000 ;
      RECT 35.885000 3.485000 36.055000 3.655000 ;
      RECT 36.365000 2.140000 36.535000 2.310000 ;
      RECT 36.365000 3.130000 36.535000 3.300000 ;
      RECT 37.345000 2.140000 37.515000 2.310000 ;
      RECT 37.345000 3.130000 37.515000 3.300000 ;
      RECT 38.285000 2.140000 38.455000 2.310000 ;
      RECT 38.285000 3.130000 38.455000 3.300000 ;
      RECT 39.745000 2.140000 39.915000 2.310000 ;
      RECT 39.745000 3.130000 39.915000 3.300000 ;
      RECT 40.685000 2.140000 40.855000 2.310000 ;
      RECT 40.685000 3.130000 40.855000 3.300000 ;
      RECT 41.665000 2.140000 41.835000 2.310000 ;
      RECT 41.665000 3.130000 41.835000 3.300000 ;
      RECT 42.145000 1.785000 42.315000 1.955000 ;
      RECT 42.145000 3.485000 42.315000 3.655000 ;
      RECT 42.615000 2.140000 42.785000 2.310000 ;
      RECT 42.615000 3.130000 42.785000 3.300000 ;
      RECT 43.085000 1.785000 43.255000 1.955000 ;
      RECT 43.085000 3.485000 43.255000 3.655000 ;
      RECT 43.565000 2.140000 43.735000 2.310000 ;
      RECT 43.565000 3.130000 43.735000 3.300000 ;
      RECT 43.845000 2.635000 44.015000 2.805000 ;
      RECT 44.305000 2.635000 44.475000 2.805000 ;
      RECT 44.765000 2.635000 44.935000 2.805000 ;
      RECT 45.225000 2.635000 45.395000 2.805000 ;
      RECT 45.685000 2.635000 45.855000 2.805000 ;
      RECT 46.145000 2.635000 46.315000 2.805000 ;
      RECT 46.605000 2.635000 46.775000 2.805000 ;
      RECT 47.065000 2.635000 47.235000 2.805000 ;
      RECT 47.345000 2.140000 47.515000 2.310000 ;
      RECT 47.345000 3.130000 47.515000 3.300000 ;
      RECT 47.825000 1.785000 47.995000 1.955000 ;
      RECT 47.825000 3.485000 47.995000 3.655000 ;
      RECT 48.295000 2.140000 48.465000 2.310000 ;
      RECT 48.295000 3.130000 48.465000 3.300000 ;
      RECT 48.765000 1.785000 48.935000 1.955000 ;
      RECT 48.765000 3.485000 48.935000 3.655000 ;
      RECT 49.245000 2.140000 49.415000 2.310000 ;
      RECT 49.245000 3.130000 49.415000 3.300000 ;
      RECT 50.225000 2.140000 50.395000 2.310000 ;
      RECT 50.225000 3.130000 50.395000 3.300000 ;
      RECT 51.165000 2.140000 51.335000 2.310000 ;
      RECT 51.165000 3.130000 51.335000 3.300000 ;
    LAYER met1 ;
      RECT  0.585000 2.110000  0.875000 2.155000 ;
      RECT  0.585000 2.155000  4.695000 2.295000 ;
      RECT  0.585000 2.295000  0.875000 2.340000 ;
      RECT  0.585000 3.100000  0.875000 3.145000 ;
      RECT  0.585000 3.145000  4.695000 3.285000 ;
      RECT  0.585000 3.285000  0.875000 3.330000 ;
      RECT  1.525000 2.110000  1.815000 2.155000 ;
      RECT  1.525000 2.295000  1.815000 2.340000 ;
      RECT  1.525000 3.100000  1.815000 3.145000 ;
      RECT  1.525000 3.285000  1.815000 3.330000 ;
      RECT  2.505000 2.110000  2.795000 2.155000 ;
      RECT  2.505000 2.295000  2.795000 2.340000 ;
      RECT  2.505000 3.100000  2.795000 3.145000 ;
      RECT  2.505000 3.285000  2.795000 3.330000 ;
      RECT  3.455000 2.110000  3.745000 2.155000 ;
      RECT  3.455000 2.295000  3.745000 2.340000 ;
      RECT  3.455000 3.100000  3.745000 3.145000 ;
      RECT  3.455000 3.285000  3.745000 3.330000 ;
      RECT  4.405000 2.110000  4.695000 2.155000 ;
      RECT  4.405000 2.295000  4.695000 2.340000 ;
      RECT  4.405000 3.100000  4.695000 3.145000 ;
      RECT  4.405000 3.285000  4.695000 3.330000 ;
      RECT  8.185000 2.110000  8.475000 2.155000 ;
      RECT  8.185000 2.155000 12.295000 2.295000 ;
      RECT  8.185000 2.295000  8.475000 2.340000 ;
      RECT  8.185000 3.100000  8.475000 3.145000 ;
      RECT  8.185000 3.145000 12.295000 3.285000 ;
      RECT  8.185000 3.285000  8.475000 3.330000 ;
      RECT  9.135000 2.110000  9.425000 2.155000 ;
      RECT  9.135000 2.295000  9.425000 2.340000 ;
      RECT  9.135000 3.100000  9.425000 3.145000 ;
      RECT  9.135000 3.285000  9.425000 3.330000 ;
      RECT 10.085000 2.110000 10.375000 2.155000 ;
      RECT 10.085000 2.295000 10.375000 2.340000 ;
      RECT 10.085000 3.100000 10.375000 3.145000 ;
      RECT 10.085000 3.285000 10.375000 3.330000 ;
      RECT 11.065000 2.110000 11.355000 2.155000 ;
      RECT 11.065000 2.295000 11.355000 2.340000 ;
      RECT 11.065000 3.100000 11.355000 3.145000 ;
      RECT 11.065000 3.285000 11.355000 3.330000 ;
      RECT 12.005000 2.110000 12.295000 2.155000 ;
      RECT 12.005000 2.295000 12.295000 2.340000 ;
      RECT 12.005000 3.100000 12.295000 3.145000 ;
      RECT 12.005000 3.285000 12.295000 3.330000 ;
      RECT 13.465000 2.110000 13.755000 2.155000 ;
      RECT 13.465000 2.155000 17.575000 2.295000 ;
      RECT 13.465000 2.295000 13.755000 2.340000 ;
      RECT 13.465000 3.100000 13.755000 3.145000 ;
      RECT 13.465000 3.145000 17.575000 3.285000 ;
      RECT 13.465000 3.285000 13.755000 3.330000 ;
      RECT 14.405000 2.110000 14.695000 2.155000 ;
      RECT 14.405000 2.295000 14.695000 2.340000 ;
      RECT 14.405000 3.100000 14.695000 3.145000 ;
      RECT 14.405000 3.285000 14.695000 3.330000 ;
      RECT 15.385000 2.110000 15.675000 2.155000 ;
      RECT 15.385000 2.295000 15.675000 2.340000 ;
      RECT 15.385000 3.100000 15.675000 3.145000 ;
      RECT 15.385000 3.285000 15.675000 3.330000 ;
      RECT 16.335000 2.110000 16.625000 2.155000 ;
      RECT 16.335000 2.295000 16.625000 2.340000 ;
      RECT 16.335000 3.100000 16.625000 3.145000 ;
      RECT 16.335000 3.285000 16.625000 3.330000 ;
      RECT 17.285000 2.110000 17.575000 2.155000 ;
      RECT 17.285000 2.295000 17.575000 2.340000 ;
      RECT 17.285000 3.100000 17.575000 3.145000 ;
      RECT 17.285000 3.285000 17.575000 3.330000 ;
      RECT 21.065000 2.110000 21.355000 2.155000 ;
      RECT 21.065000 2.155000 25.175000 2.295000 ;
      RECT 21.065000 2.295000 21.355000 2.340000 ;
      RECT 21.065000 3.100000 21.355000 3.145000 ;
      RECT 21.065000 3.145000 25.175000 3.285000 ;
      RECT 21.065000 3.285000 21.355000 3.330000 ;
      RECT 22.015000 2.110000 22.305000 2.155000 ;
      RECT 22.015000 2.295000 22.305000 2.340000 ;
      RECT 22.015000 3.100000 22.305000 3.145000 ;
      RECT 22.015000 3.285000 22.305000 3.330000 ;
      RECT 22.965000 2.110000 23.255000 2.155000 ;
      RECT 22.965000 2.295000 23.255000 2.340000 ;
      RECT 22.965000 3.100000 23.255000 3.145000 ;
      RECT 22.965000 3.285000 23.255000 3.330000 ;
      RECT 23.945000 2.110000 24.235000 2.155000 ;
      RECT 23.945000 2.295000 24.235000 2.340000 ;
      RECT 23.945000 3.100000 24.235000 3.145000 ;
      RECT 23.945000 3.285000 24.235000 3.330000 ;
      RECT 24.885000 2.110000 25.175000 2.155000 ;
      RECT 24.885000 2.295000 25.175000 2.340000 ;
      RECT 24.885000 3.100000 25.175000 3.145000 ;
      RECT 24.885000 3.285000 25.175000 3.330000 ;
      RECT 26.805000 2.110000 27.095000 2.155000 ;
      RECT 26.805000 2.155000 30.915000 2.295000 ;
      RECT 26.805000 2.295000 27.095000 2.340000 ;
      RECT 26.805000 3.100000 27.095000 3.145000 ;
      RECT 26.805000 3.145000 30.915000 3.285000 ;
      RECT 26.805000 3.285000 27.095000 3.330000 ;
      RECT 27.745000 2.110000 28.035000 2.155000 ;
      RECT 27.745000 2.295000 28.035000 2.340000 ;
      RECT 27.745000 3.100000 28.035000 3.145000 ;
      RECT 27.745000 3.285000 28.035000 3.330000 ;
      RECT 28.725000 2.110000 29.015000 2.155000 ;
      RECT 28.725000 2.295000 29.015000 2.340000 ;
      RECT 28.725000 3.100000 29.015000 3.145000 ;
      RECT 28.725000 3.285000 29.015000 3.330000 ;
      RECT 29.675000 2.110000 29.965000 2.155000 ;
      RECT 29.675000 2.295000 29.965000 2.340000 ;
      RECT 29.675000 3.100000 29.965000 3.145000 ;
      RECT 29.675000 3.285000 29.965000 3.330000 ;
      RECT 30.625000 2.110000 30.915000 2.155000 ;
      RECT 30.625000 2.295000 30.915000 2.340000 ;
      RECT 30.625000 3.100000 30.915000 3.145000 ;
      RECT 30.625000 3.285000 30.915000 3.330000 ;
      RECT 34.405000 2.110000 34.695000 2.155000 ;
      RECT 34.405000 2.155000 38.515000 2.295000 ;
      RECT 34.405000 2.295000 34.695000 2.340000 ;
      RECT 34.405000 3.100000 34.695000 3.145000 ;
      RECT 34.405000 3.145000 38.515000 3.285000 ;
      RECT 34.405000 3.285000 34.695000 3.330000 ;
      RECT 35.355000 2.110000 35.645000 2.155000 ;
      RECT 35.355000 2.295000 35.645000 2.340000 ;
      RECT 35.355000 3.100000 35.645000 3.145000 ;
      RECT 35.355000 3.285000 35.645000 3.330000 ;
      RECT 36.305000 2.110000 36.595000 2.155000 ;
      RECT 36.305000 2.295000 36.595000 2.340000 ;
      RECT 36.305000 3.100000 36.595000 3.145000 ;
      RECT 36.305000 3.285000 36.595000 3.330000 ;
      RECT 37.285000 2.110000 37.575000 2.155000 ;
      RECT 37.285000 2.295000 37.575000 2.340000 ;
      RECT 37.285000 3.100000 37.575000 3.145000 ;
      RECT 37.285000 3.285000 37.575000 3.330000 ;
      RECT 38.225000 2.110000 38.515000 2.155000 ;
      RECT 38.225000 2.295000 38.515000 2.340000 ;
      RECT 38.225000 3.100000 38.515000 3.145000 ;
      RECT 38.225000 3.285000 38.515000 3.330000 ;
      RECT 39.685000 2.110000 39.975000 2.155000 ;
      RECT 39.685000 2.155000 43.795000 2.295000 ;
      RECT 39.685000 2.295000 39.975000 2.340000 ;
      RECT 39.685000 3.100000 39.975000 3.145000 ;
      RECT 39.685000 3.145000 43.795000 3.285000 ;
      RECT 39.685000 3.285000 39.975000 3.330000 ;
      RECT 40.625000 2.110000 40.915000 2.155000 ;
      RECT 40.625000 2.295000 40.915000 2.340000 ;
      RECT 40.625000 3.100000 40.915000 3.145000 ;
      RECT 40.625000 3.285000 40.915000 3.330000 ;
      RECT 41.605000 2.110000 41.895000 2.155000 ;
      RECT 41.605000 2.295000 41.895000 2.340000 ;
      RECT 41.605000 3.100000 41.895000 3.145000 ;
      RECT 41.605000 3.285000 41.895000 3.330000 ;
      RECT 42.555000 2.110000 42.845000 2.155000 ;
      RECT 42.555000 2.295000 42.845000 2.340000 ;
      RECT 42.555000 3.100000 42.845000 3.145000 ;
      RECT 42.555000 3.285000 42.845000 3.330000 ;
      RECT 43.505000 2.110000 43.795000 2.155000 ;
      RECT 43.505000 2.295000 43.795000 2.340000 ;
      RECT 43.505000 3.100000 43.795000 3.145000 ;
      RECT 43.505000 3.285000 43.795000 3.330000 ;
      RECT 47.285000 2.110000 47.575000 2.155000 ;
      RECT 47.285000 2.155000 51.395000 2.295000 ;
      RECT 47.285000 2.295000 47.575000 2.340000 ;
      RECT 47.285000 3.100000 47.575000 3.145000 ;
      RECT 47.285000 3.145000 51.395000 3.285000 ;
      RECT 47.285000 3.285000 47.575000 3.330000 ;
      RECT 48.235000 2.110000 48.525000 2.155000 ;
      RECT 48.235000 2.295000 48.525000 2.340000 ;
      RECT 48.235000 3.100000 48.525000 3.145000 ;
      RECT 48.235000 3.285000 48.525000 3.330000 ;
      RECT 49.185000 2.110000 49.475000 2.155000 ;
      RECT 49.185000 2.295000 49.475000 2.340000 ;
      RECT 49.185000 3.100000 49.475000 3.145000 ;
      RECT 49.185000 3.285000 49.475000 3.330000 ;
      RECT 50.165000 2.110000 50.455000 2.155000 ;
      RECT 50.165000 2.295000 50.455000 2.340000 ;
      RECT 50.165000 3.100000 50.455000 3.145000 ;
      RECT 50.165000 3.285000 50.455000 3.330000 ;
      RECT 51.105000 2.110000 51.395000 2.155000 ;
      RECT 51.105000 2.295000 51.395000 2.340000 ;
      RECT 51.105000 3.100000 51.395000 3.145000 ;
      RECT 51.105000 3.285000 51.395000 3.330000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb16to1_4
END LIBRARY
