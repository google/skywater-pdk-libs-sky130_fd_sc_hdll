# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__sdlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdlclkp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.745000 1.075000 5.035000 1.120000 ;
        RECT 4.745000 1.120000 6.230000 1.260000 ;
        RECT 4.745000 1.260000 5.035000 1.305000 ;
        RECT 5.940000 1.075000 6.230000 1.120000 ;
        RECT 5.940000 1.260000 6.230000 1.305000 ;
    END
  END CLK
  PIN GATE
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 0.955000 1.235000 1.955000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.480250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.985000 0.255000 7.235000 2.465000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.330000 1.665000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.615000 ;
      RECT 0.085000  0.615000 1.295000 0.785000 ;
      RECT 0.085000  1.835000 0.345000 2.635000 ;
      RECT 0.515000  0.085000 0.895000 0.445000 ;
      RECT 0.515000  0.785000 0.685000 2.125000 ;
      RECT 0.515000  2.125000 1.280000 2.465000 ;
      RECT 1.115000  0.255000 1.295000 0.615000 ;
      RECT 1.465000  0.255000 2.645000 0.535000 ;
      RECT 1.465000  0.705000 1.800000 1.205000 ;
      RECT 1.465000  1.205000 1.960000 1.955000 ;
      RECT 1.610000  2.125000 2.300000 2.465000 ;
      RECT 1.970000  0.705000 2.305000 1.035000 ;
      RECT 2.130000  1.205000 3.205000 1.375000 ;
      RECT 2.130000  1.375000 2.300000 2.125000 ;
      RECT 2.470000  1.575000 2.665000 1.635000 ;
      RECT 2.470000  1.635000 3.545000 1.905000 ;
      RECT 2.475000  0.535000 2.645000 0.995000 ;
      RECT 2.475000  0.995000 3.205000 1.205000 ;
      RECT 2.520000  2.075000 3.105000 2.635000 ;
      RECT 2.910000  0.085000 3.080000 0.825000 ;
      RECT 3.325000  1.905000 3.545000 1.915000 ;
      RECT 3.325000  1.915000 5.735000 2.085000 ;
      RECT 3.325000  2.085000 3.545000 2.465000 ;
      RECT 3.375000  0.255000 3.545000 1.635000 ;
      RECT 3.735000  0.255000 4.065000 0.935000 ;
      RECT 3.735000  0.935000 3.905000 1.575000 ;
      RECT 3.735000  1.575000 4.145000 1.745000 ;
      RECT 3.885000  2.255000 5.735000 2.635000 ;
      RECT 4.075000  1.105000 4.550000 1.275000 ;
      RECT 4.285000  0.085000 4.615000 0.445000 ;
      RECT 4.365000  1.275000 4.550000 1.495000 ;
      RECT 4.365000  1.495000 5.215000 1.745000 ;
      RECT 4.380000  0.615000 5.215000 0.785000 ;
      RECT 4.380000  0.785000 4.550000 1.105000 ;
      RECT 4.745000  0.995000 5.060000 1.325000 ;
      RECT 4.965000  0.255000 5.215000 0.615000 ;
      RECT 5.385000  0.995000 5.735000 1.915000 ;
      RECT 5.535000  0.255000 5.705000 0.615000 ;
      RECT 5.535000  0.615000 6.815000 0.785000 ;
      RECT 5.955000  0.995000 6.395000 1.325000 ;
      RECT 5.955000  1.495000 6.815000 2.085000 ;
      RECT 5.955000  2.085000 6.125000 2.465000 ;
      RECT 6.325000  0.085000 6.685000 0.445000 ;
      RECT 6.385000  2.255000 6.715000 2.635000 ;
      RECT 6.645000  0.785000 6.815000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.625000  1.445000 1.795000 1.615000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.135000  0.765000 2.305000 0.935000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.800000  0.765000 3.970000 0.935000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.365000  1.445000 4.535000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 4.805000  1.105000 4.975000 1.275000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.000000  1.105000 6.170000 1.275000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
    LAYER met1 ;
      RECT 1.565000 1.415000 1.855000 1.460000 ;
      RECT 1.565000 1.460000 4.595000 1.600000 ;
      RECT 1.565000 1.600000 1.855000 1.645000 ;
      RECT 2.075000 0.735000 2.365000 0.780000 ;
      RECT 2.075000 0.780000 4.030000 0.920000 ;
      RECT 2.075000 0.920000 2.365000 0.965000 ;
      RECT 3.740000 0.735000 4.030000 0.780000 ;
      RECT 3.740000 0.920000 4.030000 0.965000 ;
      RECT 4.305000 1.415000 4.595000 1.460000 ;
      RECT 4.305000 1.600000 4.595000 1.645000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdlclkp_1
