* NGSPICE file created from sky130_fd_sc_hdll__xor2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__xor2_1 A B VGND VNB VPB VPWR X
M1000 VPWR A a_125_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.6e+11p pd=5.12e+06u as=3e+11p ps=2.6e+06u
M1001 X a_35_297# a_315_297# VPB phighvt w=1e+06u l=180000u
+  ad=4.5e+11p pd=2.9e+06u as=5.7e+11p ps=5.14e+06u
M1002 a_35_297# B VGND VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=7.28e+11p ps=6.14e+06u
M1003 VGND A a_35_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_35_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=5.46e+11p ps=2.98e+06u
M1005 VPWR B a_315_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_125_297# B a_35_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1007 a_317_47# A VGND VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=0p ps=0u
M1008 X B a_317_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_315_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

