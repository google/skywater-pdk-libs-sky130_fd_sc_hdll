* File: sky130_fd_sc_hdll__o2bb2a_2.pex.spice
* Created: Wed Sep  2 08:46:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_2%A_84_21# 1 2 7 9 10 12 13 15 16 18 21 25
+ 26 27 31 34 37 40 41 42 48
c118 16 0 1.10934e-19 $X=0.99 $Y=1.41
r119 47 48 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r120 46 47 57.504 $w=3.73e-07 $l=4.45e-07 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.965 $Y2=1.202
r121 45 46 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r122 42 44 0.699809 $w=5.23e-07 $l=3e-08 $layer=LI1_cond $X=3.132 $Y=1.97
+ $X2=3.132 $Y2=2
r123 40 41 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=2.905 $Y=1.075
+ $X2=2.905 $Y2=1.245
r124 39 40 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.895 $Y=0.69
+ $X2=2.895 $Y2=1.075
r125 37 39 10.7341 $w=2.43e-07 $l=2.05e-07 $layer=LI1_cond $X=2.857 $Y=0.485
+ $X2=2.857 $Y2=0.69
r126 31 42 17.0847 $w=5.23e-07 $l=5.73324e-07 $layer=LI1_cond $X=2.915 $Y=1.495
+ $X2=3.132 $Y2=1.97
r127 31 41 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.915 $Y=1.495
+ $X2=2.915 $Y2=1.245
r128 26 42 7.43996 $w=1.7e-07 $l=3.02e-07 $layer=LI1_cond $X=2.83 $Y=1.97
+ $X2=3.132 $Y2=1.97
r129 26 27 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=2.83 $Y=1.97
+ $X2=1.37 $Y2=1.97
r130 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.285 $Y=1.885
+ $X2=1.37 $Y2=1.97
r131 24 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=1.615
+ $X2=1.285 $Y2=1.53
r132 24 25 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.285 $Y=1.615
+ $X2=1.285 $Y2=1.885
r133 22 48 2.58445 $w=3.73e-07 $l=2e-08 $layer=POLY_cond $X=1.01 $Y=1.202
+ $X2=0.99 $Y2=1.202
r134 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.01
+ $Y=1.16 $X2=1.01 $Y2=1.16
r135 19 34 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.035 $Y=1.53
+ $X2=1.285 $Y2=1.53
r136 19 21 14.9294 $w=2.18e-07 $l=2.85e-07 $layer=LI1_cond $X=1.035 $Y=1.445
+ $X2=1.035 $Y2=1.16
r137 16 48 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.99 $Y=1.41
+ $X2=0.99 $Y2=1.202
r138 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.99 $Y=1.41
+ $X2=0.99 $Y2=1.985
r139 13 47 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.965 $Y=0.995
+ $X2=0.965 $Y2=1.202
r140 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.965 $Y=0.995
+ $X2=0.965 $Y2=0.56
r141 10 46 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.52 $Y=1.41
+ $X2=0.52 $Y2=1.202
r142 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.52 $Y=1.41
+ $X2=0.52 $Y2=1.985
r143 7 45 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=0.995
+ $X2=0.495 $Y2=1.202
r144 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.495 $Y=0.995
+ $X2=0.495 $Y2=0.56
r145 2 44 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=3.125
+ $Y=1.845 $X2=3.27 $Y2=2
r146 1 37 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=2.695
+ $Y=0.235 $X2=2.82 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_2%A1_N 3 6 7 9 10 13 19
c42 10 0 1.59802e-19 $X=1.525 $Y=1.095
c43 3 0 1.1853e-19 $X=1.49 $Y=0.445
r44 13 16 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.575 $Y=1.16
+ $X2=1.575 $Y2=1.325
r45 13 15 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.575 $Y=1.16
+ $X2=1.575 $Y2=0.995
r46 13 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.55
+ $Y=1.16 $X2=1.55 $Y2=1.16
r47 10 19 3.32727 $w=1.98e-07 $l=6e-08 $layer=LI1_cond $X=1.61 $Y=1.175 $X2=1.55
+ $Y2=1.175
r48 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.515 $Y=1.77
+ $X2=1.515 $Y2=2.165
r49 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.515 $Y=1.67 $X2=1.515
+ $Y2=1.77
r50 6 16 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=1.515 $Y=1.67
+ $X2=1.515 $Y2=1.325
r51 3 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.49 $Y=0.445
+ $X2=1.49 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_2%A2_N 3 5 6 8 9 12 14 17
c43 12 0 1.59802e-19 $X=2.09 $Y=0.935
r44 13 17 13.2609 $w=4.14e-07 $l=4.5e-07 $layer=LI1_cond $X=2.09 $Y=0.74
+ $X2=1.64 $Y2=0.74
r45 12 15 37.7413 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=0.935
+ $X2=2.11 $Y2=1.1
r46 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=0.935
+ $X2=2.11 $Y2=0.77
r47 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.09
+ $Y=0.935 $X2=2.09 $Y2=0.935
r48 9 17 5.98801 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.64 $Y=0.51 $X2=1.64
+ $Y2=0.74
r49 6 8 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.125 $Y=1.77
+ $X2=2.125 $Y2=2.165
r50 5 6 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.125 $Y=1.67 $X2=2.125
+ $Y2=1.77
r51 5 15 188.999 $w=2e-07 $l=5.7e-07 $layer=POLY_cond $X=2.125 $Y=1.67 $X2=2.125
+ $Y2=1.1
r52 3 14 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=2.02 $Y=0.445
+ $X2=2.02 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_2%A_321_369# 1 2 7 9 12 14 15 16 20 27 29
c69 20 0 1.1853e-19 $X=2.395 $Y=0.48
c70 16 0 1.10934e-19 $X=2.395 $Y=1.605
r71 27 29 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=2.527 $Y=1.52
+ $X2=2.527 $Y2=1.355
r72 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.575
+ $Y=1.52 $X2=2.575 $Y2=1.52
r73 24 29 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=2.48 $Y=0.565
+ $X2=2.48 $Y2=1.355
r74 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.395 $Y=0.48
+ $X2=2.48 $Y2=0.565
r75 20 22 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.395 $Y=0.48
+ $X2=2.27 $Y2=0.48
r76 16 27 3.69652 $w=2.63e-07 $l=8.5e-08 $layer=LI1_cond $X=2.527 $Y=1.605
+ $X2=2.527 $Y2=1.52
r77 16 18 29.8588 $w=2.18e-07 $l=5.7e-07 $layer=LI1_cond $X=2.395 $Y=1.605
+ $X2=1.825 $Y2=1.605
r78 14 28 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.935 $Y=1.52
+ $X2=2.575 $Y2=1.52
r79 14 15 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=2.935 $Y=1.52
+ $X2=3.035 $Y2=1.562
r80 10 15 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=3.06 $Y=1.355
+ $X2=3.035 $Y2=1.562
r81 10 12 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=3.06 $Y=1.355
+ $X2=3.06 $Y2=0.445
r82 7 15 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=3.035 $Y=1.77
+ $X2=3.035 $Y2=1.562
r83 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.035 $Y=1.77
+ $X2=3.035 $Y2=2.165
r84 2 18 600 $w=1.7e-07 $l=3.09354e-07 $layer=licon1_PDIFF $count=1 $X=1.605
+ $Y=1.845 $X2=1.825 $Y2=1.63
r85 1 22 182 $w=1.7e-07 $l=3.2078e-07 $layer=licon1_NDIFF $count=1 $X=2.095
+ $Y=0.235 $X2=2.27 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_2%B2 2 3 5 8 12 13 14 18 22 26 28
r51 18 20 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.525 $Y=1.16
+ $X2=3.525 $Y2=0.995
r52 14 28 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=3.825 $Y=2.21
+ $X2=3.825 $Y2=2.23
r53 14 26 12.8783 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=3.825 $Y=2.21
+ $X2=3.825 $Y2=1.915
r54 13 22 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=3.46 $Y=1.2 $X2=3.44
+ $Y2=1.2
r55 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.5
+ $Y=1.16 $X2=3.5 $Y2=1.16
r56 12 13 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=3.655 $Y=1.2
+ $X2=3.46 $Y2=1.2
r57 10 12 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.74 $Y=1.325
+ $X2=3.655 $Y2=1.2
r58 10 26 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.74 $Y=1.325
+ $X2=3.74 $Y2=1.915
r59 8 20 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.55 $Y=0.445
+ $X2=3.55 $Y2=0.995
r60 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.525 $Y=1.77
+ $X2=3.525 $Y2=2.165
r61 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.525 $Y=1.67 $X2=3.525
+ $Y2=1.77
r62 1 18 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.525 $Y=1.325
+ $X2=3.525 $Y2=1.16
r63 1 2 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=3.525 $Y=1.325
+ $X2=3.525 $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_2%B1 3 6 7 9 10 11 18 25
r30 16 18 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.05 $Y=1.16
+ $X2=4.215 $Y2=1.16
r31 14 16 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=4.025 $Y=1.16
+ $X2=4.05 $Y2=1.16
r32 11 25 0.128611 $w=4.63e-07 $l=5e-09 $layer=LI1_cond $X=4.232 $Y=1.53
+ $X2=4.232 $Y2=1.525
r33 10 25 9.38857 $w=4.63e-07 $l=3.65e-07 $layer=LI1_cond $X=4.232 $Y=1.16
+ $X2=4.232 $Y2=1.525
r34 10 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.215
+ $Y=1.16 $X2=4.215 $Y2=1.16
r35 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=4.05 $Y=1.77 $X2=4.05
+ $Y2=2.165
r36 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.05 $Y=1.67 $X2=4.05
+ $Y2=1.77
r37 5 16 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.05 $Y=1.325 $X2=4.05
+ $Y2=1.16
r38 5 6 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=4.05 $Y=1.325 $X2=4.05
+ $Y2=1.67
r39 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.025 $Y=0.995
+ $X2=4.025 $Y2=1.16
r40 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.025 $Y=0.995
+ $X2=4.025 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_2%VPWR 1 2 3 4 13 15 21 23 25 27 29 34 39
+ 51 54 62 66
r62 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r63 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r64 48 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r65 46 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r66 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r67 43 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r68 43 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r69 42 45 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r70 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r71 40 42 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.765 $Y=2.72
+ $X2=2.99 $Y2=2.72
r72 39 61 4.58008 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=4.165 $Y=2.72
+ $X2=4.382 $Y2=2.72
r73 39 45 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.165 $Y=2.72
+ $X2=3.91 $Y2=2.72
r74 38 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r75 38 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r76 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r77 35 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.39 $Y=2.72 $X2=1.2
+ $Y2=2.72
r78 35 37 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.39 $Y=2.72
+ $X2=2.07 $Y2=2.72
r79 34 40 5.85399 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=2.562 $Y=2.72
+ $X2=2.765 $Y2=2.72
r80 34 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r81 34 54 11.3822 $w=4.03e-07 $l=4e-07 $layer=LI1_cond $X=2.562 $Y=2.72
+ $X2=2.562 $Y2=2.32
r82 34 37 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.36 $Y=2.72
+ $X2=2.07 $Y2=2.72
r83 33 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r84 33 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r85 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r86 30 48 4.06635 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=2.72
+ $X2=0.182 $Y2=2.72
r87 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=2.72
+ $X2=0.69 $Y2=2.72
r88 29 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.01 $Y=2.72 $X2=1.2
+ $Y2=2.72
r89 29 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.01 $Y=2.72 $X2=0.69
+ $Y2=2.72
r90 27 66 0.00284542 $w=4.8e-07 $l=1e-08 $layer=MET1_cond $X=0.22 $Y=2.72
+ $X2=0.23 $Y2=2.72
r91 23 61 3.06042 $w=3.15e-07 $l=1.11018e-07 $layer=LI1_cond $X=4.322 $Y=2.635
+ $X2=4.382 $Y2=2.72
r92 23 25 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=4.322 $Y=2.635
+ $X2=4.322 $Y2=2
r93 19 51 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.72
r94 19 21 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.32
r95 15 18 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.237 $Y=1.62
+ $X2=0.237 $Y2=2.3
r96 13 48 3.11087 $w=2.55e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.237 $Y=2.635
+ $X2=0.182 $Y2=2.72
r97 13 18 15.1399 $w=2.53e-07 $l=3.35e-07 $layer=LI1_cond $X=0.237 $Y=2.635
+ $X2=0.237 $Y2=2.3
r98 4 25 300 $w=1.7e-07 $l=2.19203e-07 $layer=licon1_PDIFF $count=2 $X=4.14
+ $Y=1.845 $X2=4.295 $Y2=2
r99 3 54 600 $w=1.7e-07 $l=6.25999e-07 $layer=licon1_PDIFF $count=1 $X=2.215
+ $Y=1.845 $X2=2.565 $Y2=2.32
r100 2 21 600 $w=1.7e-07 $l=9.04599e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.485 $X2=1.225 $Y2=2.32
r101 1 18 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r102 1 15 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_2%X 1 2 10 13 14 15 18
r30 15 18 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=0.687 $Y=2.21
+ $X2=0.687 $Y2=1.96
r31 13 18 0.491205 $w=3.03e-07 $l=1.3e-08 $layer=LI1_cond $X=0.687 $Y=1.947
+ $X2=0.687 $Y2=1.96
r32 13 14 6.65738 $w=3.03e-07 $l=1.52e-07 $layer=LI1_cond $X=0.687 $Y=1.947
+ $X2=0.687 $Y2=1.795
r33 12 14 50.8123 $w=2.18e-07 $l=9.7e-07 $layer=LI1_cond $X=0.645 $Y=0.825
+ $X2=0.645 $Y2=1.795
r34 10 12 15.7188 $w=3.83e-07 $l=4.55e-07 $layer=LI1_cond $X=0.727 $Y=0.37
+ $X2=0.727 $Y2=0.825
r35 2 18 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.61
+ $Y=1.485 $X2=0.755 $Y2=1.96
r36 1 10 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.235 $X2=0.755 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_2%VGND 1 2 3 10 12 14 18 22 25 26 27 37 38
+ 44 49
r58 45 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.23
+ $Y2=0
r59 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r60 41 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r61 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r62 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r63 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r64 32 35 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=3.45
+ $Y2=0
r65 32 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r66 31 34 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=3.45
+ $Y2=0
r67 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r68 29 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.22
+ $Y2=0
r69 29 31 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.61
+ $Y2=0
r70 27 49 0.00284542 $w=4.8e-07 $l=1e-08 $layer=MET1_cond $X=0.22 $Y=0 $X2=0.23
+ $Y2=0
r71 25 34 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.675 $Y=0 $X2=3.45
+ $Y2=0
r72 25 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=0 $X2=3.76
+ $Y2=0
r73 24 37 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.845 $Y=0 $X2=4.37
+ $Y2=0
r74 24 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.845 $Y=0 $X2=3.76
+ $Y2=0
r75 20 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.76 $Y=0.085
+ $X2=3.76 $Y2=0
r76 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.76 $Y=0.085
+ $X2=3.76 $Y2=0.39
r77 16 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r78 16 18 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.525
r79 15 41 4.06635 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r80 14 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.22
+ $Y2=0
r81 14 15 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=0 $X2=0.365
+ $Y2=0
r82 10 41 3.11087 $w=2.55e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.237 $Y=0.085
+ $X2=0.182 $Y2=0
r83 10 12 12.8802 $w=2.53e-07 $l=2.85e-07 $layer=LI1_cond $X=0.237 $Y=0.085
+ $X2=0.237 $Y2=0.37
r84 3 22 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.625
+ $Y=0.235 $X2=3.76 $Y2=0.39
r85 2 18 182 $w=1.7e-07 $l=3.69188e-07 $layer=licon1_NDIFF $count=1 $X=1.04
+ $Y=0.235 $X2=1.22 $Y2=0.525
r86 1 12 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_2%A_627_47# 1 2 9 11 12 15
r31 13 15 8.56945 $w=3.88e-07 $l=2.9e-07 $layer=LI1_cond $X=4.21 $Y=0.725
+ $X2=4.21 $Y2=0.435
r32 11 13 8.0953 $w=1.8e-07 $l=2.35743e-07 $layer=LI1_cond $X=4.015 $Y=0.815
+ $X2=4.21 $Y2=0.725
r33 11 12 35.7374 $w=1.78e-07 $l=5.8e-07 $layer=LI1_cond $X=4.015 $Y=0.815
+ $X2=3.435 $Y2=0.815
r34 7 12 6.94918 $w=1.8e-07 $l=1.53542e-07 $layer=LI1_cond $X=3.32 $Y=0.725
+ $X2=3.435 $Y2=0.815
r35 7 9 12.0255 $w=2.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.32 $Y=0.725 $X2=3.32
+ $Y2=0.485
r36 2 15 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=4.1
+ $Y=0.235 $X2=4.24 $Y2=0.435
r37 1 9 182 $w=1.7e-07 $l=3.18198e-07 $layer=licon1_NDIFF $count=1 $X=3.135
+ $Y=0.235 $X2=3.29 $Y2=0.485
.ends

