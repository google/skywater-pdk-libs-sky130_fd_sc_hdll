* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hdll__muxb4to1_1 D[3] D[2] D[1] D[0] S[3] S[2] S[1] S[0] VGND VNB VPB VPWR Z
*.PININFO D[3]:I D[2]:I D[1]:I D[0]:I S[3]:I S[2]:I S[1]:I S[0]:I
*.PININFO VGND:I VNB:I VPB:I VPWR:I Z:O
MMNA00 Z S[0] VNB nshort m=1 w=0.52 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 net87 D[0] VNB nshort m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 SB0 S[0] VNB nshort m=1 w=0.52 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI30 Z S[2] VNB nshort m=1 w=0.52 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI29 net51 D[2] VNB nshort m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI28 SB2 S[2] VNB nshort m=1 w=0.52 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI27 SB3 S[3] VNB nshort m=1 w=0.52 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI26 net63 D[3] VNB nshort m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Z S[3] VNB nshort m=1 w=0.52 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI13 Z S[1] VNB nshort m=1 w=0.52 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI12 net75 D[1] VNB nshort m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI11 SB1 S[1] VNB nshort m=1 w=0.52 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI35 net99 SB2 VPB phighvt m=1 w=0.82 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI34 SB2 S[2] VPB phighvt m=1 w=1.0 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR D[0] VPB phighvt m=1 w=1.0 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 net135 SB0 VPB phighvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 SB3 S[3] VPB phighvt m=1 w=1.0 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net111 SB3 VPB phighvt m=1 w=0.82 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI31 VPWR D[3] VPB phighvt m=1 w=1.0 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 SB0 S[0] VPB phighvt m=1 w=1.0 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI15 net123 SB1 VPB phighvt m=1 w=0.82 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI16 VPWR D[1] VPB phighvt m=1 w=1.0 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI14 SB1 S[1] VPB phighvt m=1 w=1.0 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI36 VPWR D[2] VPB phighvt m=1 w=1.0 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_hdll__muxb4to1_1
