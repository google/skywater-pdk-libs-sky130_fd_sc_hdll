* File: sky130_fd_sc_hdll__sedfxbp_2.pxi.spice
* Created: Thu Aug 27 19:28:39 2020
* 
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%CLK N_CLK_c_298_n N_CLK_c_302_n N_CLK_c_303_n
+ N_CLK_M1007_g N_CLK_c_299_n N_CLK_M1037_g CLK
+ PM_SKY130_FD_SC_HDLL__SEDFXBP_2%CLK
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_27_47# N_A_27_47#_M1037_s N_A_27_47#_M1007_s
+ N_A_27_47#_c_348_n N_A_27_47#_c_349_n N_A_27_47#_M1041_g N_A_27_47#_M1001_g
+ N_A_27_47#_M1013_g N_A_27_47#_c_350_n N_A_27_47#_M1032_g N_A_27_47#_c_351_n
+ N_A_27_47#_c_352_n N_A_27_47#_M1003_g N_A_27_47#_c_337_n N_A_27_47#_M1021_g
+ N_A_27_47#_c_597_p N_A_27_47#_c_339_n N_A_27_47#_c_340_n N_A_27_47#_c_354_n
+ N_A_27_47#_c_490_p N_A_27_47#_c_341_n N_A_27_47#_c_342_n N_A_27_47#_c_343_n
+ N_A_27_47#_c_344_n N_A_27_47#_c_357_n N_A_27_47#_c_358_n N_A_27_47#_c_359_n
+ N_A_27_47#_c_360_n N_A_27_47#_c_361_n N_A_27_47#_c_362_n N_A_27_47#_c_363_n
+ N_A_27_47#_c_345_n N_A_27_47#_c_346_n N_A_27_47#_c_347_n
+ PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%D N_D_c_616_n N_D_c_621_n N_D_M1023_g
+ N_D_M1043_g D N_D_c_619_n PM_SKY130_FD_SC_HDLL__SEDFXBP_2%D
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_455_324# N_A_455_324#_M1034_s
+ N_A_455_324#_M1006_s N_A_455_324#_c_669_n N_A_455_324#_M1029_g
+ N_A_455_324#_c_670_n N_A_455_324#_c_671_n N_A_455_324#_M1035_g
+ N_A_455_324#_c_672_n N_A_455_324#_c_664_n N_A_455_324#_c_665_n
+ N_A_455_324#_c_666_n N_A_455_324#_c_667_n N_A_455_324#_c_674_n
+ N_A_455_324#_c_668_n PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_455_324#
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%DE N_DE_M1045_g N_DE_c_762_n N_DE_c_763_n
+ N_DE_c_769_n N_DE_M1006_g N_DE_M1034_g N_DE_c_770_n N_DE_c_771_n N_DE_M1025_g
+ N_DE_c_765_n N_DE_c_772_n N_DE_c_773_n DE N_DE_c_766_n DE
+ PM_SKY130_FD_SC_HDLL__SEDFXBP_2%DE
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_851_264# N_A_851_264#_M1018_s
+ N_A_851_264#_M1005_s N_A_851_264#_c_869_n N_A_851_264#_M1026_g
+ N_A_851_264#_M1009_g N_A_851_264#_c_852_n N_A_851_264#_c_872_n
+ N_A_851_264#_M1039_g N_A_851_264#_M1004_g N_A_851_264#_c_854_n
+ N_A_851_264#_c_855_n N_A_851_264#_M1011_g N_A_851_264#_M1017_g
+ N_A_851_264#_c_857_n N_A_851_264#_c_858_n N_A_851_264#_M1020_g
+ N_A_851_264#_M1033_g N_A_851_264#_c_860_n N_A_851_264#_c_861_n
+ N_A_851_264#_c_862_n N_A_851_264#_c_876_n N_A_851_264#_c_863_n
+ N_A_851_264#_c_864_n N_A_851_264#_c_865_n N_A_851_264#_c_866_n
+ N_A_851_264#_c_867_n N_A_851_264#_c_1063_p N_A_851_264#_c_868_n
+ PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_851_264#
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_955_21# N_A_955_21#_M1015_s
+ N_A_955_21#_M1022_s N_A_955_21#_c_1083_n N_A_955_21#_M1019_g
+ N_A_955_21#_c_1084_n N_A_955_21#_c_1085_n N_A_955_21#_c_1086_n
+ N_A_955_21#_c_1087_n N_A_955_21#_M1014_g N_A_955_21#_c_1088_n
+ N_A_955_21#_c_1089_n N_A_955_21#_c_1090_n N_A_955_21#_c_1091_n
+ N_A_955_21#_c_1096_n N_A_955_21#_c_1092_n N_A_955_21#_c_1098_n
+ N_A_955_21#_c_1093_n PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_955_21#
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%SCD N_SCD_c_1201_n N_SCD_M1036_g N_SCD_M1038_g
+ SCD PM_SKY130_FD_SC_HDLL__SEDFXBP_2%SCD
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%SCE N_SCE_c_1248_n N_SCE_M1030_g
+ N_SCE_c_1241_n N_SCE_c_1250_n N_SCE_M1022_g N_SCE_M1015_g N_SCE_c_1243_n
+ N_SCE_c_1244_n N_SCE_M1024_g N_SCE_c_1251_n SCE N_SCE_c_1247_n SCE
+ PM_SKY130_FD_SC_HDLL__SEDFXBP_2%SCE
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_211_363# N_A_211_363#_M1001_d
+ N_A_211_363#_M1041_d N_A_211_363#_c_1342_n N_A_211_363#_c_1343_n
+ N_A_211_363#_M1027_g N_A_211_363#_c_1333_n N_A_211_363#_M1042_g
+ N_A_211_363#_c_1335_n N_A_211_363#_M1012_g N_A_211_363#_c_1345_n
+ N_A_211_363#_M1046_g N_A_211_363#_c_1336_n N_A_211_363#_c_1337_n
+ N_A_211_363#_c_1346_n N_A_211_363#_c_1347_n N_A_211_363#_c_1348_n
+ N_A_211_363#_c_1349_n N_A_211_363#_c_1397_n N_A_211_363#_c_1338_n
+ N_A_211_363#_c_1339_n N_A_211_363#_c_1340_n N_A_211_363#_c_1341_n
+ PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_211_363#
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_1787_159# N_A_1787_159#_M1047_d
+ N_A_1787_159#_M1000_d N_A_1787_159#_c_1547_n N_A_1787_159#_c_1559_n
+ N_A_1787_159#_M1028_g N_A_1787_159#_M1040_g N_A_1787_159#_c_1560_n
+ N_A_1787_159#_c_1561_n N_A_1787_159#_M1002_g N_A_1787_159#_M1010_g
+ N_A_1787_159#_c_1550_n N_A_1787_159#_c_1551_n N_A_1787_159#_c_1552_n
+ N_A_1787_159#_c_1553_n N_A_1787_159#_c_1564_n N_A_1787_159#_c_1554_n
+ N_A_1787_159#_c_1555_n N_A_1787_159#_c_1556_n N_A_1787_159#_c_1557_n
+ PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_1787_159#
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_1611_413# N_A_1611_413#_M1013_d
+ N_A_1611_413#_M1027_d N_A_1611_413#_c_1672_n N_A_1611_413#_c_1679_n
+ N_A_1611_413#_M1000_g N_A_1611_413#_M1047_g N_A_1611_413#_c_1673_n
+ N_A_1611_413#_c_1674_n N_A_1611_413#_c_1675_n N_A_1611_413#_c_1676_n
+ N_A_1611_413#_c_1686_n N_A_1611_413#_c_1691_n N_A_1611_413#_c_1677_n
+ N_A_1611_413#_c_1682_n N_A_1611_413#_c_1678_n
+ PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_1611_413#
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_2266_413# N_A_2266_413#_M1012_d
+ N_A_2266_413#_M1003_d N_A_2266_413#_c_1788_n N_A_2266_413#_M1018_g
+ N_A_2266_413#_c_1789_n N_A_2266_413#_M1005_g N_A_2266_413#_c_1782_n
+ N_A_2266_413#_c_1783_n N_A_2266_413#_c_1784_n N_A_2266_413#_M1031_g
+ N_A_2266_413#_c_1792_n N_A_2266_413#_M1008_g N_A_2266_413#_c_1793_n
+ N_A_2266_413#_M1016_g N_A_2266_413#_c_1785_n N_A_2266_413#_M1044_g
+ N_A_2266_413#_c_1786_n N_A_2266_413#_c_1801_n N_A_2266_413#_c_1805_n
+ N_A_2266_413#_c_1795_n N_A_2266_413#_c_1796_n N_A_2266_413#_c_1787_n
+ N_A_2266_413#_c_1798_n N_A_2266_413#_c_1799_n N_A_2266_413#_c_1800_n
+ PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_2266_413#
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%VPWR N_VPWR_M1007_d N_VPWR_M1029_d
+ N_VPWR_M1006_d N_VPWR_M1022_d N_VPWR_M1028_d N_VPWR_M1002_s N_VPWR_M1039_d
+ N_VPWR_M1020_d N_VPWR_M1005_d N_VPWR_M1016_d N_VPWR_c_1918_n N_VPWR_c_1919_n
+ N_VPWR_c_1920_n N_VPWR_c_1921_n N_VPWR_c_1922_n N_VPWR_c_1923_n
+ N_VPWR_c_1924_n N_VPWR_c_1925_n N_VPWR_c_1926_n N_VPWR_c_1927_n
+ N_VPWR_c_1928_n N_VPWR_c_1929_n N_VPWR_c_1930_n N_VPWR_c_1931_n
+ N_VPWR_c_1932_n N_VPWR_c_1933_n N_VPWR_c_1934_n N_VPWR_c_1935_n VPWR
+ N_VPWR_c_1936_n N_VPWR_c_1937_n N_VPWR_c_1938_n N_VPWR_c_1939_n
+ N_VPWR_c_1940_n N_VPWR_c_1941_n N_VPWR_c_1917_n N_VPWR_c_1943_n
+ N_VPWR_c_1944_n N_VPWR_c_1945_n N_VPWR_c_1946_n N_VPWR_c_1947_n
+ N_VPWR_c_1948_n N_VPWR_c_1949_n PM_SKY130_FD_SC_HDLL__SEDFXBP_2%VPWR
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_319_47# N_A_319_47#_M1043_s
+ N_A_319_47#_M1009_d N_A_319_47#_M1023_s N_A_319_47#_M1026_d
+ N_A_319_47#_c_2152_n N_A_319_47#_c_2145_n N_A_319_47#_c_2154_n
+ N_A_319_47#_c_2146_n N_A_319_47#_c_2147_n N_A_319_47#_c_2148_n
+ N_A_319_47#_c_2176_n N_A_319_47#_c_2149_n N_A_319_47#_c_2150_n
+ N_A_319_47#_c_2151_n PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_319_47#
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_985_47# N_A_985_47#_M1019_d
+ N_A_985_47#_M1024_d N_A_985_47#_M1030_d N_A_985_47#_M1014_d
+ N_A_985_47#_c_2269_n N_A_985_47#_c_2270_n N_A_985_47#_c_2260_n
+ N_A_985_47#_c_2282_n N_A_985_47#_c_2346_n N_A_985_47#_c_2261_n
+ N_A_985_47#_c_2271_n N_A_985_47#_c_2262_n N_A_985_47#_c_2263_n
+ N_A_985_47#_c_2286_n N_A_985_47#_c_2264_n N_A_985_47#_c_2265_n
+ N_A_985_47#_c_2266_n N_A_985_47#_c_2267_n N_A_985_47#_c_2320_n
+ N_A_985_47#_c_2268_n PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_985_47#
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%Q_N N_Q_N_M1017_s N_Q_N_M1011_s N_Q_N_c_2398_n
+ N_Q_N_c_2396_n Q_N PM_SKY130_FD_SC_HDLL__SEDFXBP_2%Q_N
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%Q N_Q_M1031_s N_Q_M1008_s Q N_Q_c_2426_n
+ PM_SKY130_FD_SC_HDLL__SEDFXBP_2%Q
x_PM_SKY130_FD_SC_HDLL__SEDFXBP_2%VGND N_VGND_M1037_d N_VGND_M1045_d
+ N_VGND_M1034_d N_VGND_M1015_d N_VGND_M1040_d N_VGND_M1010_s N_VGND_M1004_d
+ N_VGND_M1033_d N_VGND_M1018_d N_VGND_M1044_d N_VGND_c_2446_n N_VGND_c_2447_n
+ N_VGND_c_2448_n N_VGND_c_2449_n N_VGND_c_2450_n N_VGND_c_2451_n
+ N_VGND_c_2452_n N_VGND_c_2453_n N_VGND_c_2454_n N_VGND_c_2455_n
+ N_VGND_c_2456_n N_VGND_c_2457_n N_VGND_c_2458_n N_VGND_c_2459_n
+ N_VGND_c_2460_n N_VGND_c_2461_n VGND N_VGND_c_2462_n N_VGND_c_2463_n
+ N_VGND_c_2464_n N_VGND_c_2465_n N_VGND_c_2466_n N_VGND_c_2467_n
+ N_VGND_c_2468_n N_VGND_c_2469_n N_VGND_c_2470_n N_VGND_c_2471_n
+ N_VGND_c_2472_n N_VGND_c_2473_n N_VGND_c_2474_n N_VGND_c_2475_n
+ N_VGND_c_2476_n PM_SKY130_FD_SC_HDLL__SEDFXBP_2%VGND
cc_1 VNB N_CLK_c_298_n 0.0607903f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.325
cc_2 VNB N_CLK_c_299_n 0.0173562f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_3 VNB CLK 0.0188452f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_27_47#_M1001_g 0.0407387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_27_47#_M1013_g 0.0226463f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_c_337_n 0.0172417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_M1021_g 0.0473175f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_339_n 0.00353743f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_340_n 0.00651432f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_341_n 0.00717927f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_342_n 0.00381138f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_343_n 0.0337321f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_344_n 0.00481323f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_345_n 0.0272085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_346_n 0.00998637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_347_n 0.00232986f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_D_c_616_n 0.0138173f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.59
cc_18 VNB N_D_M1043_g 0.0309027f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_19 VNB D 0.00799811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_D_c_619_n 0.0194093f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_21 VNB N_A_455_324#_M1035_g 0.022764f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_455_324#_c_664_n 0.00785922f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_455_324#_c_665_n 0.00185686f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_455_324#_c_666_n 0.00358193f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_455_324#_c_667_n 0.0343111f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_455_324#_c_668_n 0.00239244f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_DE_M1045_g 0.021472f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.74
cc_28 VNB N_DE_c_762_n 0.0423212f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_29 VNB N_DE_c_763_n 0.0199457f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_30 VNB N_DE_M1034_g 0.0240367f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_DE_c_765_n 0.00610496f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_DE_c_766_n 0.0393836f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB DE 0.00860916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_851_264#_M1009_g 0.0497249f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_851_264#_c_852_n 0.00428343f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_36 VNB N_A_851_264#_M1004_g 0.0320214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_851_264#_c_854_n 0.0139483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_851_264#_c_855_n 0.010325f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_851_264#_M1017_g 0.0194597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_851_264#_c_857_n 0.00981196f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_851_264#_c_858_n 0.0154134f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_851_264#_M1033_g 0.0216027f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_851_264#_c_860_n 0.0346803f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_851_264#_c_861_n 0.0105805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_851_264#_c_862_n 0.0039678f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_851_264#_c_863_n 0.0320138f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_851_264#_c_864_n 0.00234899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_851_264#_c_865_n 0.0518632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_851_264#_c_866_n 0.00529256f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_851_264#_c_867_n 0.0137497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_851_264#_c_868_n 0.00964094f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_955_21#_c_1083_n 0.0196804f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_53 VNB N_A_955_21#_c_1084_n 0.0481338f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_955_21#_c_1085_n 0.00817921f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.665
cc_55 VNB N_A_955_21#_c_1086_n 0.0171161f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_56 VNB N_A_955_21#_c_1087_n 0.0126951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_955_21#_c_1088_n 0.0105942f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_58 VNB N_A_955_21#_c_1089_n 0.0348285f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_955_21#_c_1090_n 0.00278382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_955_21#_c_1091_n 0.00492913f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_955_21#_c_1092_n 0.00242064f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_955_21#_c_1093_n 0.00209066f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_SCD_c_1201_n 0.00932499f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.325
cc_64 VNB N_SCD_M1038_g 0.0270642f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_65 VNB SCD 0.00977457f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_66 VNB N_SCE_c_1241_n 0.00789916f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_67 VNB N_SCE_M1015_g 0.0230411f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_SCE_c_1243_n 0.0624009f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_69 VNB N_SCE_c_1244_n 0.011117f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_SCE_M1024_g 0.0325532f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_71 VNB SCE 0.00613801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_SCE_c_1247_n 0.0500998f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_211_363#_c_1333_n 0.0156862f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_211_363#_M1042_g 0.0445483f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_75 VNB N_A_211_363#_c_1335_n 0.0190887f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_211_363#_c_1336_n 0.00834745f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_211_363#_c_1337_n 0.0351046f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_211_363#_c_1338_n 0.00914674f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_211_363#_c_1339_n 0.00271227f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_211_363#_c_1340_n 0.0180788f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_211_363#_c_1341_n 0.0128135f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_1787_159#_c_1547_n 0.0152162f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_83 VNB N_A_1787_159#_M1040_g 0.0207384f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1787_159#_M1010_g 0.0293639f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_1787_159#_c_1550_n 0.0249115f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_1787_159#_c_1551_n 0.00801699f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_1787_159#_c_1552_n 0.00935939f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_1787_159#_c_1553_n 0.00632297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_1787_159#_c_1554_n 0.0048611f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_1787_159#_c_1555_n 0.0179853f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_1787_159#_c_1556_n 0.00296193f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_A_1787_159#_c_1557_n 0.0348905f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_A_1611_413#_c_1672_n 0.0123393f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_94 VNB N_A_1611_413#_c_1673_n 0.0186444f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_95 VNB N_A_1611_413#_c_1674_n 0.0155462f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_96 VNB N_A_1611_413#_c_1675_n 0.00937366f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_97 VNB N_A_1611_413#_c_1676_n 0.0013343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_A_1611_413#_c_1677_n 0.0120473f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_A_1611_413#_c_1678_n 0.00183626f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_A_2266_413#_M1018_g 0.0347962f $X=-0.19 $Y=-0.24 $X2=0.495
+ $Y2=1.665
cc_101 VNB N_A_2266_413#_c_1782_n 0.0160411f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_102 VNB N_A_2266_413#_c_1783_n 0.0127576f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_103 VNB N_A_2266_413#_c_1784_n 0.0174548f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_A_2266_413#_c_1785_n 0.0224588f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_A_2266_413#_c_1786_n 0.0446091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_A_2266_413#_c_1787_n 0.00885691f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VPWR_c_1917_n 0.687231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_A_319_47#_c_2145_n 0.0139975f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_A_319_47#_c_2146_n 0.00299149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_A_319_47#_c_2147_n 0.00512225f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_A_319_47#_c_2148_n 0.00419923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_A_319_47#_c_2149_n 0.00440827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_A_319_47#_c_2150_n 0.0031955f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_A_319_47#_c_2151_n 0.00404434f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_A_985_47#_c_2260_n 3.20364e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_A_985_47#_c_2261_n 0.00225385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_A_985_47#_c_2262_n 0.0127253f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_A_985_47#_c_2263_n 0.00860855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_A_985_47#_c_2264_n 0.00551087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_A_985_47#_c_2265_n 7.96116e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_A_985_47#_c_2266_n 3.04222e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_A_985_47#_c_2267_n 0.00804403f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_A_985_47#_c_2268_n 0.00374428f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_Q_N_c_2396_n 0.00144373f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_125 VNB N_Q_c_2426_n 0.00103515f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2446_n 0.00487083f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2447_n 0.0165213f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2448_n 4.14276e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2449_n 0.00698291f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2450_n 0.00312457f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2451_n 0.00532105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2452_n 0.0096851f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2453_n 0.0176082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2454_n 0.00925922f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2455_n 0.0342122f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2456_n 0.023337f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2457_n 0.00526448f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2458_n 0.0212244f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2459_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2460_n 0.0207574f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2461_n 0.00500104f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2462_n 0.0154125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2463_n 0.04097f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2464_n 0.0688491f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2465_n 0.0632245f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2466_n 0.0526425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2467_n 0.0289267f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2468_n 0.0142356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2469_n 0.767424f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2470_n 0.0085923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2471_n 0.00597653f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2472_n 0.00503538f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2473_n 0.00332923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2474_n 0.00626777f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2475_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2476_n 0.00451684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_157 VPB N_CLK_c_298_n 0.00482568f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_158 VPB N_CLK_c_302_n 0.0148284f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.59
cc_159 VPB N_CLK_c_303_n 0.0462588f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.74
cc_160 VPB CLK 0.017793f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_161 VPB N_A_27_47#_c_348_n 0.0181622f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_162 VPB N_A_27_47#_c_349_n 0.0252424f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_163 VPB N_A_27_47#_c_350_n 0.0523214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_27_47#_c_351_n 0.0155789f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_27_47#_c_352_n 0.0223707f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_27_47#_c_337_n 0.0236548f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_27_47#_c_354_n 0.0019617f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_27_47#_c_341_n 0.00381244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_27_47#_c_344_n 0.00305108f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_27_47#_c_357_n 0.0035907f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_27_47#_c_358_n 0.0363003f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_27_47#_c_359_n 0.00167529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_27_47#_c_360_n 0.0139626f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_27_47#_c_361_n 0.00104792f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_27_47#_c_362_n 0.00810591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_27_47#_c_363_n 0.00485115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_27_47#_c_345_n 0.0122883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_27_47#_c_346_n 0.0226921f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_27_47#_c_347_n 0.00668639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_D_c_616_n 0.0418959f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.59
cc_181 VPB N_D_c_621_n 0.0191809f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.74
cc_182 VPB D 0.0062301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_455_324#_c_669_n 0.0182034f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_184 VPB N_A_455_324#_c_670_n 0.00981795f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_455_324#_c_671_n 0.0100724f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.665
cc_186 VPB N_A_455_324#_c_672_n 0.00766443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_455_324#_c_665_n 0.00615652f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_455_324#_c_674_n 0.0411589f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_DE_c_763_n 0.0115068f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_190 VPB N_DE_c_769_n 0.0196068f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_191 VPB N_DE_c_770_n 0.0203478f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_192 VPB N_DE_c_771_n 0.0168391f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_DE_c_772_n 0.0145969f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_DE_c_773_n 0.0186843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB DE 0.00252241f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_A_851_264#_c_869_n 0.0578051f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_197 VPB N_A_851_264#_M1009_g 8.38539e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_A_851_264#_c_852_n 0.0345155f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.16
cc_199 VPB N_A_851_264#_c_872_n 0.0241801f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_200 VPB N_A_851_264#_c_855_n 0.0227078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_A_851_264#_c_858_n 0.0288671f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_A_851_264#_c_862_n 0.0151347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_A_851_264#_c_876_n 0.00672509f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_A_851_264#_c_867_n 6.92652e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_A_955_21#_c_1087_n 0.0437816f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_A_955_21#_c_1091_n 0.00606327f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_A_955_21#_c_1096_n 0.00533522f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_A_955_21#_c_1092_n 0.00164978f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_A_955_21#_c_1098_n 0.0117193f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_SCD_c_1201_n 0.0408369f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_211 VPB SCD 0.00359136f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_212 VPB N_SCE_c_1248_n 0.0197112f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_213 VPB N_SCE_c_1241_n 0.0295713f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_214 VPB N_SCE_c_1250_n 0.0203812f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_215 VPB N_SCE_c_1251_n 0.0221203f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB SCE 0.00360919f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_SCE_c_1247_n 0.0402931f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_A_211_363#_c_1342_n 0.0247149f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_219 VPB N_A_211_363#_c_1343_n 0.0247192f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_220 VPB N_A_211_363#_c_1333_n 0.0149739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_A_211_363#_c_1345_n 0.0534851f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_A_211_363#_c_1346_n 0.0410924f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_A_211_363#_c_1347_n 0.00567492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_A_211_363#_c_1348_n 0.0216005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_A_211_363#_c_1349_n 0.00120291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_A_211_363#_c_1338_n 0.00694839f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_A_211_363#_c_1339_n 0.00152248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_A_211_363#_c_1340_n 0.0145882f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_A_211_363#_c_1341_n 0.00996908f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB N_A_1787_159#_c_1547_n 0.0337045f $X=-0.19 $Y=1.305 $X2=0.52
+ $Y2=0.445
cc_231 VPB N_A_1787_159#_c_1559_n 0.0249303f $X=-0.19 $Y=1.305 $X2=0.31
+ $Y2=1.665
cc_232 VPB N_A_1787_159#_c_1560_n 0.03542f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_233 VPB N_A_1787_159#_c_1561_n 0.0276825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_A_1787_159#_c_1551_n 0.00992693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_A_1787_159#_c_1552_n 0.00154645f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_A_1787_159#_c_1564_n 0.0156409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_A_1787_159#_c_1554_n 0.00366659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_A_1611_413#_c_1679_n 0.0213145f $X=-0.19 $Y=1.305 $X2=0.31
+ $Y2=1.665
cc_239 VPB N_A_1611_413#_c_1675_n 0.0189038f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_240 VPB N_A_1611_413#_c_1676_n 0.0207029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 VPB N_A_1611_413#_c_1682_n 0.00398435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_242 VPB N_A_1611_413#_c_1678_n 0.00937022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_243 VPB N_A_2266_413#_c_1788_n 0.0387442f $X=-0.19 $Y=1.305 $X2=0.52
+ $Y2=0.445
cc_244 VPB N_A_2266_413#_c_1789_n 0.0194331f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_245 VPB N_A_2266_413#_c_1782_n 0.011803f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_246 VPB N_A_2266_413#_c_1783_n 0.0252249f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_247 VPB N_A_2266_413#_c_1792_n 0.0164032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_248 VPB N_A_2266_413#_c_1793_n 0.0202373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_249 VPB N_A_2266_413#_c_1786_n 0.0235016f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_250 VPB N_A_2266_413#_c_1795_n 0.00756022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_251 VPB N_A_2266_413#_c_1796_n 0.00270536f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_252 VPB N_A_2266_413#_c_1787_n 0.00515957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_253 VPB N_A_2266_413#_c_1798_n 0.0033711f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_254 VPB N_A_2266_413#_c_1799_n 0.0427106f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_255 VPB N_A_2266_413#_c_1800_n 0.00417984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1918_n 0.00126291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1919_n 0.00853665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1920_n 0.007127f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1921_n 0.00571282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1922_n 0.0696924f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1923_n 0.00506553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1924_n 0.00900651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1925_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1926_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1927_n 0.0196453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1928_n 0.01027f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1929_n 0.0475361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1930_n 0.0209492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1931_n 0.00372488f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1932_n 0.0204002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1933_n 0.00555304f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1934_n 0.0211826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1935_n 0.00497514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1936_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1937_n 0.0397223f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1938_n 0.0727682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1939_n 0.0530696f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1940_n 0.0317155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1941_n 0.0142356f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_1917_n 0.0912717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_281 VPB N_VPWR_c_1943_n 0.0054556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_282 VPB N_VPWR_c_1944_n 0.00580385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_283 VPB N_VPWR_c_1945_n 0.00660741f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_284 VPB N_VPWR_c_1946_n 0.00449095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_285 VPB N_VPWR_c_1947_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_286 VPB N_VPWR_c_1948_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_287 VPB N_VPWR_c_1949_n 0.00449427f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_288 VPB N_A_319_47#_c_2152_n 0.00774922f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_289 VPB N_A_319_47#_c_2145_n 0.00993433f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_290 VPB N_A_319_47#_c_2154_n 0.00168019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_291 VPB N_A_319_47#_c_2146_n 0.00408201f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_292 VPB N_A_985_47#_c_2269_n 0.00307437f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.16
cc_293 VPB N_A_985_47#_c_2270_n 0.00414607f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_294 VPB N_A_985_47#_c_2271_n 0.00411328f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_295 VPB N_A_985_47#_c_2262_n 0.00951926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_296 VPB N_A_985_47#_c_2264_n 0.00658861f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_297 N_CLK_c_302_n N_A_27_47#_c_348_n 0.00267643f $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_298 N_CLK_c_303_n N_A_27_47#_c_348_n 0.0066814f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_299 CLK N_A_27_47#_c_348_n 8.10055e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_300 N_CLK_c_303_n N_A_27_47#_c_349_n 0.0193458f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_301 N_CLK_c_298_n N_A_27_47#_M1001_g 0.00195891f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_302 N_CLK_c_299_n N_A_27_47#_M1001_g 0.0154156f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_303 N_CLK_c_298_n N_A_27_47#_c_339_n 0.0107746f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_304 N_CLK_c_299_n N_A_27_47#_c_339_n 0.00644237f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_305 CLK N_A_27_47#_c_339_n 0.00774265f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_306 N_CLK_c_298_n N_A_27_47#_c_340_n 0.00622672f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_307 CLK N_A_27_47#_c_340_n 0.0144574f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_308 N_CLK_c_303_n N_A_27_47#_c_354_n 0.0170291f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_309 CLK N_A_27_47#_c_354_n 0.00769886f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_310 N_CLK_c_298_n N_A_27_47#_c_341_n 0.00280606f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_311 N_CLK_c_302_n N_A_27_47#_c_341_n 4.49617e-19 $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_312 N_CLK_c_303_n N_A_27_47#_c_341_n 0.00442243f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_313 CLK N_A_27_47#_c_341_n 0.0421632f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_314 N_CLK_c_298_n N_A_27_47#_c_357_n 2.46885e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_315 N_CLK_c_303_n N_A_27_47#_c_357_n 0.00784199f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_316 CLK N_A_27_47#_c_357_n 0.0153591f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_317 N_CLK_c_303_n N_A_27_47#_c_359_n 0.00102492f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_318 N_CLK_c_298_n N_A_27_47#_c_345_n 0.0130772f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_319 CLK N_A_27_47#_c_345_n 0.00184152f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_320 N_CLK_c_303_n N_VPWR_c_1918_n 0.0125197f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_321 N_CLK_c_303_n N_VPWR_c_1936_n 0.00304525f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_322 N_CLK_c_303_n N_VPWR_c_1917_n 0.00454898f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_323 N_CLK_c_298_n N_VGND_c_2462_n 6.28829e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_324 N_CLK_c_299_n N_VGND_c_2462_n 0.00198377f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_325 N_CLK_c_299_n N_VGND_c_2469_n 0.00367064f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_326 N_CLK_c_299_n N_VGND_c_2470_n 0.0142867f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_327 N_A_27_47#_c_348_n N_D_c_616_n 0.00409608f $X=0.965 $Y=1.64 $X2=0 $Y2=0
cc_328 N_A_27_47#_c_358_n N_D_c_616_n 0.00191722f $X=8.285 $Y=1.87 $X2=0 $Y2=0
cc_329 N_A_27_47#_c_358_n N_D_c_621_n 0.00555057f $X=8.285 $Y=1.87 $X2=0 $Y2=0
cc_330 N_A_27_47#_c_358_n D 0.00999475f $X=8.285 $Y=1.87 $X2=0 $Y2=0
cc_331 N_A_27_47#_M1001_g N_D_c_619_n 0.00409608f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_332 N_A_27_47#_c_358_n N_A_455_324#_c_669_n 0.00424473f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_333 N_A_27_47#_c_358_n N_A_455_324#_c_670_n 0.00790328f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_334 N_A_27_47#_c_358_n N_A_455_324#_c_672_n 0.0224406f $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_358_n N_A_455_324#_c_665_n 0.00660521f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_336 N_A_27_47#_c_358_n N_DE_c_769_n 0.00475911f $X=8.285 $Y=1.87 $X2=0 $Y2=0
cc_337 N_A_27_47#_c_358_n N_DE_c_770_n 0.00347671f $X=8.285 $Y=1.87 $X2=0 $Y2=0
cc_338 N_A_27_47#_c_358_n N_DE_c_771_n 0.00684461f $X=8.285 $Y=1.87 $X2=0 $Y2=0
cc_339 N_A_27_47#_c_358_n N_DE_c_772_n 2.07787e-19 $X=8.285 $Y=1.87 $X2=0 $Y2=0
cc_340 N_A_27_47#_c_358_n N_DE_c_773_n 3.29055e-19 $X=8.285 $Y=1.87 $X2=0 $Y2=0
cc_341 N_A_27_47#_c_358_n N_A_851_264#_c_869_n 0.00648269f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_342 N_A_27_47#_c_337_n N_A_851_264#_c_852_n 0.0110221f $X=11.92 $Y=1.32 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_M1021_g N_A_851_264#_M1004_g 0.0320946f $X=11.995 $Y=0.415
+ $X2=0 $Y2=0
cc_344 N_A_27_47#_M1021_g N_A_851_264#_c_861_n 0.0110221f $X=11.995 $Y=0.415
+ $X2=0 $Y2=0
cc_345 N_A_27_47#_c_358_n N_A_851_264#_c_876_n 0.00953293f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_346 N_A_27_47#_c_337_n N_A_851_264#_c_865_n 2.99626e-19 $X=11.92 $Y=1.32
+ $X2=0 $Y2=0
cc_347 N_A_27_47#_M1021_g N_A_851_264#_c_865_n 0.00914271f $X=11.995 $Y=0.415
+ $X2=0 $Y2=0
cc_348 N_A_27_47#_c_342_n N_A_851_264#_c_865_n 0.030906f $X=8.285 $Y=0.845 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_343_n N_A_851_264#_c_865_n 0.00164034f $X=8.065 $Y=0.87
+ $X2=0 $Y2=0
cc_350 N_A_27_47#_c_346_n N_A_851_264#_c_865_n 8.58822e-19 $X=11.235 $Y=1.32
+ $X2=0 $Y2=0
cc_351 N_A_27_47#_c_347_n N_A_851_264#_c_865_n 0.00657388f $X=11.21 $Y=1.41
+ $X2=0 $Y2=0
cc_352 N_A_27_47#_c_358_n N_A_955_21#_c_1087_n 0.00278526f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_353 N_A_27_47#_c_358_n N_A_955_21#_c_1091_n 0.00420532f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_354 N_A_27_47#_c_358_n N_A_955_21#_c_1096_n 0.0424464f $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_358_n N_A_955_21#_c_1092_n 0.00628866f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_356 N_A_27_47#_c_358_n N_A_955_21#_c_1098_n 0.0222884f $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_358_n N_SCD_c_1201_n 0.0038756f $X=8.285 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_358 N_A_27_47#_c_358_n SCD 0.00346426f $X=8.285 $Y=1.87 $X2=0 $Y2=0
cc_359 N_A_27_47#_c_358_n N_SCE_c_1248_n 0.00459204f $X=8.285 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_360 N_A_27_47#_c_358_n N_SCE_c_1241_n 0.00181115f $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_358_n N_SCE_c_1250_n 9.20215e-19 $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_c_358_n SCE 0.00649921f $X=8.285 $Y=1.87 $X2=0 $Y2=0
cc_363 N_A_27_47#_c_358_n N_SCE_c_1247_n 2.07787e-19 $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_358_n N_A_211_363#_M1041_d 0.00143359f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_365 N_A_27_47#_c_350_n N_A_211_363#_c_1342_n 0.0168071f $X=8.47 $Y=1.99 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_344_n N_A_211_363#_c_1342_n 7.27568e-19 $X=8.37 $Y=1.655
+ $X2=0 $Y2=0
cc_367 N_A_27_47#_c_358_n N_A_211_363#_c_1342_n 0.00322923f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_368 N_A_27_47#_c_362_n N_A_211_363#_c_1342_n 0.00242228f $X=8.43 $Y=1.87
+ $X2=0 $Y2=0
cc_369 N_A_27_47#_c_350_n N_A_211_363#_c_1343_n 0.00983697f $X=8.47 $Y=1.99
+ $X2=0 $Y2=0
cc_370 N_A_27_47#_c_358_n N_A_211_363#_c_1343_n 0.00394649f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_371 N_A_27_47#_c_350_n N_A_211_363#_c_1333_n 0.021571f $X=8.47 $Y=1.99 $X2=0
+ $Y2=0
cc_372 N_A_27_47#_c_344_n N_A_211_363#_c_1333_n 0.0124116f $X=8.37 $Y=1.655
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_362_n N_A_211_363#_c_1333_n 0.00177023f $X=8.43 $Y=1.87
+ $X2=0 $Y2=0
cc_374 N_A_27_47#_M1013_g N_A_211_363#_M1042_g 0.0144482f $X=8.075 $Y=0.415
+ $X2=0 $Y2=0
cc_375 N_A_27_47#_c_342_n N_A_211_363#_M1042_g 0.00159135f $X=8.285 $Y=0.845
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_c_343_n N_A_211_363#_M1042_g 0.0129656f $X=8.065 $Y=0.87 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_c_344_n N_A_211_363#_M1042_g 0.00498229f $X=8.37 $Y=1.655
+ $X2=0 $Y2=0
cc_378 N_A_27_47#_M1021_g N_A_211_363#_c_1335_n 0.0136144f $X=11.995 $Y=0.415
+ $X2=0 $Y2=0
cc_379 N_A_27_47#_c_351_n N_A_211_363#_c_1345_n 0.0185582f $X=11.24 $Y=1.89
+ $X2=0 $Y2=0
cc_380 N_A_27_47#_c_352_n N_A_211_363#_c_1345_n 0.0115366f $X=11.24 $Y=1.99
+ $X2=0 $Y2=0
cc_381 N_A_27_47#_c_337_n N_A_211_363#_c_1345_n 0.0254956f $X=11.92 $Y=1.32
+ $X2=0 $Y2=0
cc_382 N_A_27_47#_c_347_n N_A_211_363#_c_1345_n 8.74813e-19 $X=11.21 $Y=1.41
+ $X2=0 $Y2=0
cc_383 N_A_27_47#_M1021_g N_A_211_363#_c_1336_n 0.00817915f $X=11.995 $Y=0.415
+ $X2=0 $Y2=0
cc_384 N_A_27_47#_c_346_n N_A_211_363#_c_1336_n 9.61914e-19 $X=11.235 $Y=1.32
+ $X2=0 $Y2=0
cc_385 N_A_27_47#_M1021_g N_A_211_363#_c_1337_n 0.0125766f $X=11.995 $Y=0.415
+ $X2=0 $Y2=0
cc_386 N_A_27_47#_c_346_n N_A_211_363#_c_1337_n 0.0237533f $X=11.235 $Y=1.32
+ $X2=0 $Y2=0
cc_387 N_A_27_47#_c_347_n N_A_211_363#_c_1337_n 9.45568e-19 $X=11.21 $Y=1.41
+ $X2=0 $Y2=0
cc_388 N_A_27_47#_c_358_n N_A_211_363#_c_1346_n 0.514674f $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_c_348_n N_A_211_363#_c_1347_n 0.00667151f $X=0.965 $Y=1.64
+ $X2=0 $Y2=0
cc_390 N_A_27_47#_c_349_n N_A_211_363#_c_1347_n 5.76646e-19 $X=0.965 $Y=1.74
+ $X2=0 $Y2=0
cc_391 N_A_27_47#_c_341_n N_A_211_363#_c_1347_n 0.00696231f $X=0.81 $Y=1.235
+ $X2=0 $Y2=0
cc_392 N_A_27_47#_c_358_n N_A_211_363#_c_1347_n 0.0309287f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_393 N_A_27_47#_c_350_n N_A_211_363#_c_1348_n 0.00216832f $X=8.47 $Y=1.99
+ $X2=0 $Y2=0
cc_394 N_A_27_47#_c_337_n N_A_211_363#_c_1348_n 0.00218822f $X=11.92 $Y=1.32
+ $X2=0 $Y2=0
cc_395 N_A_27_47#_c_342_n N_A_211_363#_c_1348_n 0.00220528f $X=8.285 $Y=0.845
+ $X2=0 $Y2=0
cc_396 N_A_27_47#_c_344_n N_A_211_363#_c_1348_n 0.0124914f $X=8.37 $Y=1.655
+ $X2=0 $Y2=0
cc_397 N_A_27_47#_c_358_n N_A_211_363#_c_1348_n 0.00995021f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_398 N_A_27_47#_c_360_n N_A_211_363#_c_1348_n 0.196783f $X=11.075 $Y=1.87
+ $X2=0 $Y2=0
cc_399 N_A_27_47#_c_361_n N_A_211_363#_c_1348_n 0.0298939f $X=8.625 $Y=1.87
+ $X2=0 $Y2=0
cc_400 N_A_27_47#_c_362_n N_A_211_363#_c_1348_n 0.00803098f $X=8.43 $Y=1.87
+ $X2=0 $Y2=0
cc_401 N_A_27_47#_c_363_n N_A_211_363#_c_1348_n 0.0303318f $X=11.245 $Y=1.87
+ $X2=0 $Y2=0
cc_402 N_A_27_47#_c_346_n N_A_211_363#_c_1348_n 0.00376297f $X=11.235 $Y=1.32
+ $X2=0 $Y2=0
cc_403 N_A_27_47#_c_347_n N_A_211_363#_c_1348_n 0.0173469f $X=11.21 $Y=1.41
+ $X2=0 $Y2=0
cc_404 N_A_27_47#_c_342_n N_A_211_363#_c_1349_n 0.0013998f $X=8.285 $Y=0.845
+ $X2=0 $Y2=0
cc_405 N_A_27_47#_c_344_n N_A_211_363#_c_1349_n 0.0026225f $X=8.37 $Y=1.655
+ $X2=0 $Y2=0
cc_406 N_A_27_47#_c_358_n N_A_211_363#_c_1349_n 0.0312586f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_407 N_A_27_47#_c_347_n N_A_211_363#_c_1397_n 6.55244e-19 $X=11.21 $Y=1.41
+ $X2=0 $Y2=0
cc_408 N_A_27_47#_c_351_n N_A_211_363#_c_1338_n 0.00138907f $X=11.24 $Y=1.89
+ $X2=0 $Y2=0
cc_409 N_A_27_47#_c_352_n N_A_211_363#_c_1338_n 6.84267e-19 $X=11.24 $Y=1.99
+ $X2=0 $Y2=0
cc_410 N_A_27_47#_c_337_n N_A_211_363#_c_1338_n 0.0204748f $X=11.92 $Y=1.32
+ $X2=0 $Y2=0
cc_411 N_A_27_47#_c_363_n N_A_211_363#_c_1338_n 0.00833156f $X=11.245 $Y=1.87
+ $X2=0 $Y2=0
cc_412 N_A_27_47#_c_346_n N_A_211_363#_c_1338_n 0.00355741f $X=11.235 $Y=1.32
+ $X2=0 $Y2=0
cc_413 N_A_27_47#_c_347_n N_A_211_363#_c_1338_n 0.0524851f $X=11.21 $Y=1.41
+ $X2=0 $Y2=0
cc_414 N_A_27_47#_c_350_n N_A_211_363#_c_1339_n 3.56164e-19 $X=8.47 $Y=1.99
+ $X2=0 $Y2=0
cc_415 N_A_27_47#_c_342_n N_A_211_363#_c_1339_n 0.0150461f $X=8.285 $Y=0.845
+ $X2=0 $Y2=0
cc_416 N_A_27_47#_c_343_n N_A_211_363#_c_1339_n 0.0014811f $X=8.065 $Y=0.87
+ $X2=0 $Y2=0
cc_417 N_A_27_47#_c_344_n N_A_211_363#_c_1339_n 0.0374134f $X=8.37 $Y=1.655
+ $X2=0 $Y2=0
cc_418 N_A_27_47#_c_358_n N_A_211_363#_c_1339_n 0.00512466f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_419 N_A_27_47#_c_362_n N_A_211_363#_c_1339_n 0.0054038f $X=8.43 $Y=1.87 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_c_342_n N_A_211_363#_c_1340_n 0.00120953f $X=8.285 $Y=0.845
+ $X2=0 $Y2=0
cc_421 N_A_27_47#_c_343_n N_A_211_363#_c_1340_n 0.0243754f $X=8.065 $Y=0.87
+ $X2=0 $Y2=0
cc_422 N_A_27_47#_c_344_n N_A_211_363#_c_1340_n 0.00284165f $X=8.37 $Y=1.655
+ $X2=0 $Y2=0
cc_423 N_A_27_47#_c_358_n N_A_211_363#_c_1340_n 5.87167e-19 $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_424 N_A_27_47#_c_349_n N_A_211_363#_c_1341_n 0.00679553f $X=0.965 $Y=1.74
+ $X2=0 $Y2=0
cc_425 N_A_27_47#_M1001_g N_A_211_363#_c_1341_n 0.0179095f $X=0.99 $Y=0.445
+ $X2=0 $Y2=0
cc_426 N_A_27_47#_c_339_n N_A_211_363#_c_1341_n 0.0105335f $X=0.665 $Y=0.72
+ $X2=0 $Y2=0
cc_427 N_A_27_47#_c_490_p N_A_211_363#_c_1341_n 0.00861371f $X=0.78 $Y=1.795
+ $X2=0 $Y2=0
cc_428 N_A_27_47#_c_341_n N_A_211_363#_c_1341_n 0.0573128f $X=0.81 $Y=1.235
+ $X2=0 $Y2=0
cc_429 N_A_27_47#_c_358_n N_A_211_363#_c_1341_n 0.0127022f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_430 N_A_27_47#_c_359_n N_A_211_363#_c_1341_n 0.00258866f $X=0.915 $Y=1.87
+ $X2=0 $Y2=0
cc_431 N_A_27_47#_c_350_n N_A_1787_159#_c_1547_n 0.0209375f $X=8.47 $Y=1.99
+ $X2=0 $Y2=0
cc_432 N_A_27_47#_c_344_n N_A_1787_159#_c_1547_n 0.00160354f $X=8.37 $Y=1.655
+ $X2=0 $Y2=0
cc_433 N_A_27_47#_c_360_n N_A_1787_159#_c_1547_n 6.76291e-19 $X=11.075 $Y=1.87
+ $X2=0 $Y2=0
cc_434 N_A_27_47#_c_362_n N_A_1787_159#_c_1547_n 0.00193479f $X=8.43 $Y=1.87
+ $X2=0 $Y2=0
cc_435 N_A_27_47#_c_350_n N_A_1787_159#_c_1559_n 0.0233814f $X=8.47 $Y=1.99
+ $X2=0 $Y2=0
cc_436 N_A_27_47#_c_360_n N_A_1787_159#_c_1559_n 6.48115e-19 $X=11.075 $Y=1.87
+ $X2=0 $Y2=0
cc_437 N_A_27_47#_c_351_n N_A_1787_159#_c_1560_n 0.008386f $X=11.24 $Y=1.89
+ $X2=0 $Y2=0
cc_438 N_A_27_47#_c_360_n N_A_1787_159#_c_1560_n 0.00459776f $X=11.075 $Y=1.87
+ $X2=0 $Y2=0
cc_439 N_A_27_47#_c_363_n N_A_1787_159#_c_1560_n 6.96835e-19 $X=11.245 $Y=1.87
+ $X2=0 $Y2=0
cc_440 N_A_27_47#_c_347_n N_A_1787_159#_c_1560_n 0.00631585f $X=11.21 $Y=1.41
+ $X2=0 $Y2=0
cc_441 N_A_27_47#_c_352_n N_A_1787_159#_c_1561_n 0.0336123f $X=11.24 $Y=1.99
+ $X2=0 $Y2=0
cc_442 N_A_27_47#_c_360_n N_A_1787_159#_c_1561_n 0.00472081f $X=11.075 $Y=1.87
+ $X2=0 $Y2=0
cc_443 N_A_27_47#_c_363_n N_A_1787_159#_c_1561_n 6.96835e-19 $X=11.245 $Y=1.87
+ $X2=0 $Y2=0
cc_444 N_A_27_47#_c_346_n N_A_1787_159#_c_1551_n 0.0192899f $X=11.235 $Y=1.32
+ $X2=0 $Y2=0
cc_445 N_A_27_47#_c_347_n N_A_1787_159#_c_1551_n 0.00204249f $X=11.21 $Y=1.41
+ $X2=0 $Y2=0
cc_446 N_A_27_47#_c_360_n N_A_1787_159#_c_1564_n 0.0292026f $X=11.075 $Y=1.87
+ $X2=0 $Y2=0
cc_447 N_A_27_47#_c_346_n N_A_1787_159#_c_1554_n 4.77663e-19 $X=11.235 $Y=1.32
+ $X2=0 $Y2=0
cc_448 N_A_27_47#_c_347_n N_A_1787_159#_c_1554_n 0.00497295f $X=11.21 $Y=1.41
+ $X2=0 $Y2=0
cc_449 N_A_27_47#_c_360_n N_A_1611_413#_c_1679_n 0.00297942f $X=11.075 $Y=1.87
+ $X2=0 $Y2=0
cc_450 N_A_27_47#_c_360_n N_A_1611_413#_c_1675_n 2.40114e-19 $X=11.075 $Y=1.87
+ $X2=0 $Y2=0
cc_451 N_A_27_47#_c_350_n N_A_1611_413#_c_1686_n 0.011692f $X=8.47 $Y=1.99 $X2=0
+ $Y2=0
cc_452 N_A_27_47#_c_358_n N_A_1611_413#_c_1686_n 0.00635946f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_453 N_A_27_47#_c_360_n N_A_1611_413#_c_1686_n 0.00551164f $X=11.075 $Y=1.87
+ $X2=0 $Y2=0
cc_454 N_A_27_47#_c_361_n N_A_1611_413#_c_1686_n 0.00137467f $X=8.625 $Y=1.87
+ $X2=0 $Y2=0
cc_455 N_A_27_47#_c_362_n N_A_1611_413#_c_1686_n 0.0312078f $X=8.43 $Y=1.87
+ $X2=0 $Y2=0
cc_456 N_A_27_47#_M1013_g N_A_1611_413#_c_1691_n 0.00355834f $X=8.075 $Y=0.415
+ $X2=0 $Y2=0
cc_457 N_A_27_47#_c_342_n N_A_1611_413#_c_1691_n 0.0205671f $X=8.285 $Y=0.845
+ $X2=0 $Y2=0
cc_458 N_A_27_47#_c_343_n N_A_1611_413#_c_1691_n 0.00269571f $X=8.065 $Y=0.87
+ $X2=0 $Y2=0
cc_459 N_A_27_47#_c_342_n N_A_1611_413#_c_1677_n 0.0124197f $X=8.285 $Y=0.845
+ $X2=0 $Y2=0
cc_460 N_A_27_47#_c_344_n N_A_1611_413#_c_1677_n 0.0208376f $X=8.37 $Y=1.655
+ $X2=0 $Y2=0
cc_461 N_A_27_47#_c_350_n N_A_1611_413#_c_1682_n 0.00170495f $X=8.47 $Y=1.99
+ $X2=0 $Y2=0
cc_462 N_A_27_47#_c_344_n N_A_1611_413#_c_1682_n 0.00189525f $X=8.37 $Y=1.655
+ $X2=0 $Y2=0
cc_463 N_A_27_47#_c_360_n N_A_1611_413#_c_1682_n 0.0158254f $X=11.075 $Y=1.87
+ $X2=0 $Y2=0
cc_464 N_A_27_47#_c_361_n N_A_1611_413#_c_1682_n 4.1916e-19 $X=8.625 $Y=1.87
+ $X2=0 $Y2=0
cc_465 N_A_27_47#_c_362_n N_A_1611_413#_c_1682_n 0.0259876f $X=8.43 $Y=1.87
+ $X2=0 $Y2=0
cc_466 N_A_27_47#_c_350_n N_A_1611_413#_c_1678_n 5.89706e-19 $X=8.47 $Y=1.99
+ $X2=0 $Y2=0
cc_467 N_A_27_47#_c_344_n N_A_1611_413#_c_1678_n 0.0121159f $X=8.37 $Y=1.655
+ $X2=0 $Y2=0
cc_468 N_A_27_47#_c_360_n N_A_1611_413#_c_1678_n 0.00326146f $X=11.075 $Y=1.87
+ $X2=0 $Y2=0
cc_469 N_A_27_47#_c_362_n N_A_1611_413#_c_1678_n 0.00725124f $X=8.43 $Y=1.87
+ $X2=0 $Y2=0
cc_470 N_A_27_47#_c_352_n N_A_2266_413#_c_1801_n 0.00621924f $X=11.24 $Y=1.99
+ $X2=0 $Y2=0
cc_471 N_A_27_47#_c_363_n N_A_2266_413#_c_1801_n 0.00260872f $X=11.245 $Y=1.87
+ $X2=0 $Y2=0
cc_472 N_A_27_47#_c_346_n N_A_2266_413#_c_1801_n 3.11257e-19 $X=11.235 $Y=1.32
+ $X2=0 $Y2=0
cc_473 N_A_27_47#_c_347_n N_A_2266_413#_c_1801_n 0.00456497f $X=11.21 $Y=1.41
+ $X2=0 $Y2=0
cc_474 N_A_27_47#_M1021_g N_A_2266_413#_c_1805_n 0.013125f $X=11.995 $Y=0.415
+ $X2=0 $Y2=0
cc_475 N_A_27_47#_M1021_g N_A_2266_413#_c_1787_n 0.00856983f $X=11.995 $Y=0.415
+ $X2=0 $Y2=0
cc_476 N_A_27_47#_c_490_p N_VPWR_M1007_d 7.14517e-19 $X=0.78 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_477 N_A_27_47#_c_359_n N_VPWR_M1007_d 0.00186599f $X=0.915 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_478 N_A_27_47#_c_358_n N_VPWR_M1006_d 0.00160392f $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_479 N_A_27_47#_c_360_n N_VPWR_M1028_d 0.00540134f $X=11.075 $Y=1.87 $X2=0
+ $Y2=0
cc_480 N_A_27_47#_c_349_n N_VPWR_c_1918_n 0.00966647f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_481 N_A_27_47#_c_354_n N_VPWR_c_1918_n 0.00694587f $X=0.665 $Y=1.88 $X2=0
+ $Y2=0
cc_482 N_A_27_47#_c_490_p N_VPWR_c_1918_n 0.0133392f $X=0.78 $Y=1.795 $X2=0
+ $Y2=0
cc_483 N_A_27_47#_c_357_n N_VPWR_c_1918_n 0.0246493f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_484 N_A_27_47#_c_359_n N_VPWR_c_1918_n 0.00323377f $X=0.915 $Y=1.87 $X2=0
+ $Y2=0
cc_485 N_A_27_47#_c_358_n N_VPWR_c_1919_n 0.0201046f $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_486 N_A_27_47#_c_358_n N_VPWR_c_1920_n 0.0156853f $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_487 N_A_27_47#_c_358_n N_VPWR_c_1921_n 0.00159236f $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_488 N_A_27_47#_c_350_n N_VPWR_c_1922_n 0.00451183f $X=8.47 $Y=1.99 $X2=0
+ $Y2=0
cc_489 N_A_27_47#_c_360_n N_VPWR_c_1923_n 0.0123459f $X=11.075 $Y=1.87 $X2=0
+ $Y2=0
cc_490 N_A_27_47#_c_360_n N_VPWR_c_1924_n 0.0110731f $X=11.075 $Y=1.87 $X2=0
+ $Y2=0
cc_491 N_A_27_47#_c_354_n N_VPWR_c_1936_n 0.00180073f $X=0.665 $Y=1.88 $X2=0
+ $Y2=0
cc_492 N_A_27_47#_c_357_n N_VPWR_c_1936_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_493 N_A_27_47#_c_349_n N_VPWR_c_1937_n 0.00590576f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_494 N_A_27_47#_c_352_n N_VPWR_c_1939_n 0.00517771f $X=11.24 $Y=1.99 $X2=0
+ $Y2=0
cc_495 N_A_27_47#_c_347_n N_VPWR_c_1939_n 0.00157744f $X=11.21 $Y=1.41 $X2=0
+ $Y2=0
cc_496 N_A_27_47#_c_349_n N_VPWR_c_1917_n 0.00665321f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_497 N_A_27_47#_c_350_n N_VPWR_c_1917_n 0.0063841f $X=8.47 $Y=1.99 $X2=0 $Y2=0
cc_498 N_A_27_47#_c_352_n N_VPWR_c_1917_n 0.00670492f $X=11.24 $Y=1.99 $X2=0
+ $Y2=0
cc_499 N_A_27_47#_c_354_n N_VPWR_c_1917_n 0.00424724f $X=0.665 $Y=1.88 $X2=0
+ $Y2=0
cc_500 N_A_27_47#_c_357_n N_VPWR_c_1917_n 0.00646745f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_501 N_A_27_47#_c_358_n N_VPWR_c_1917_n 0.350505f $X=8.285 $Y=1.87 $X2=0 $Y2=0
cc_502 N_A_27_47#_c_359_n N_VPWR_c_1917_n 0.0145686f $X=0.915 $Y=1.87 $X2=0
+ $Y2=0
cc_503 N_A_27_47#_c_360_n N_VPWR_c_1917_n 0.11717f $X=11.075 $Y=1.87 $X2=0 $Y2=0
cc_504 N_A_27_47#_c_361_n N_VPWR_c_1917_n 0.0169341f $X=8.625 $Y=1.87 $X2=0
+ $Y2=0
cc_505 N_A_27_47#_c_363_n N_VPWR_c_1917_n 0.0186701f $X=11.245 $Y=1.87 $X2=0
+ $Y2=0
cc_506 N_A_27_47#_c_347_n N_VPWR_c_1917_n 0.0010813f $X=11.21 $Y=1.41 $X2=0
+ $Y2=0
cc_507 N_A_27_47#_c_358_n N_A_319_47#_c_2152_n 0.0202026f $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_508 N_A_27_47#_c_358_n N_A_319_47#_c_2145_n 0.00810658f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_509 N_A_27_47#_c_358_n N_A_319_47#_c_2154_n 0.0246407f $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_510 N_A_27_47#_c_358_n N_A_319_47#_c_2146_n 0.00322049f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_511 N_A_27_47#_M1001_g N_A_319_47#_c_2151_n 0.00147169f $X=0.99 $Y=0.445
+ $X2=0 $Y2=0
cc_512 N_A_27_47#_c_358_n A_409_369# 0.00326461f $X=8.285 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_513 N_A_27_47#_c_358_n A_787_369# 0.00545759f $X=8.285 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_514 N_A_27_47#_c_358_n N_A_985_47#_M1030_d 8.03832e-19 $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_515 N_A_27_47#_c_358_n N_A_985_47#_M1014_d 0.00130039f $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_516 N_A_27_47#_c_358_n N_A_985_47#_c_2269_n 0.0118087f $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_517 N_A_27_47#_c_358_n N_A_985_47#_c_2270_n 0.00875376f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_518 N_A_27_47#_M1013_g N_A_985_47#_c_2260_n 0.00568611f $X=8.075 $Y=0.415
+ $X2=0 $Y2=0
cc_519 N_A_27_47#_c_342_n N_A_985_47#_c_2260_n 0.0143664f $X=8.285 $Y=0.845
+ $X2=0 $Y2=0
cc_520 N_A_27_47#_c_343_n N_A_985_47#_c_2260_n 0.00171528f $X=8.065 $Y=0.87
+ $X2=0 $Y2=0
cc_521 N_A_27_47#_c_344_n N_A_985_47#_c_2260_n 0.00573062f $X=8.37 $Y=1.655
+ $X2=0 $Y2=0
cc_522 N_A_27_47#_c_358_n N_A_985_47#_c_2282_n 0.0130137f $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_523 N_A_27_47#_c_361_n N_A_985_47#_c_2282_n 3.07396e-19 $X=8.625 $Y=1.87
+ $X2=0 $Y2=0
cc_524 N_A_27_47#_c_362_n N_A_985_47#_c_2282_n 0.0033501f $X=8.43 $Y=1.87 $X2=0
+ $Y2=0
cc_525 N_A_27_47#_c_358_n N_A_985_47#_c_2271_n 0.0014312f $X=8.285 $Y=1.87 $X2=0
+ $Y2=0
cc_526 N_A_27_47#_c_358_n N_A_985_47#_c_2286_n 0.00255293f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_527 N_A_27_47#_c_358_n N_A_985_47#_c_2264_n 0.00597671f $X=8.285 $Y=1.87
+ $X2=0 $Y2=0
cc_528 N_A_27_47#_c_361_n N_A_985_47#_c_2264_n 2.82202e-19 $X=8.625 $Y=1.87
+ $X2=0 $Y2=0
cc_529 N_A_27_47#_c_362_n N_A_985_47#_c_2264_n 0.00325205f $X=8.43 $Y=1.87 $X2=0
+ $Y2=0
cc_530 N_A_27_47#_M1013_g N_A_985_47#_c_2268_n 0.0071201f $X=8.075 $Y=0.415
+ $X2=0 $Y2=0
cc_531 N_A_27_47#_c_342_n N_A_985_47#_c_2268_n 0.00131254f $X=8.285 $Y=0.845
+ $X2=0 $Y2=0
cc_532 N_A_27_47#_c_343_n N_A_985_47#_c_2268_n 4.36817e-19 $X=8.065 $Y=0.87
+ $X2=0 $Y2=0
cc_533 N_A_27_47#_c_339_n N_VGND_M1037_d 0.00226918f $X=0.665 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_534 N_A_27_47#_c_597_p N_VGND_c_2462_n 0.00725596f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_535 N_A_27_47#_c_339_n N_VGND_c_2462_n 0.00244154f $X=0.665 $Y=0.72 $X2=0
+ $Y2=0
cc_536 N_A_27_47#_M1001_g N_VGND_c_2463_n 0.00585385f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_537 N_A_27_47#_M1013_g N_VGND_c_2465_n 0.00433784f $X=8.075 $Y=0.415 $X2=0
+ $Y2=0
cc_538 N_A_27_47#_c_342_n N_VGND_c_2465_n 0.00293266f $X=8.285 $Y=0.845 $X2=0
+ $Y2=0
cc_539 N_A_27_47#_c_343_n N_VGND_c_2465_n 0.00108996f $X=8.065 $Y=0.87 $X2=0
+ $Y2=0
cc_540 N_A_27_47#_M1021_g N_VGND_c_2466_n 0.00373071f $X=11.995 $Y=0.415 $X2=0
+ $Y2=0
cc_541 N_A_27_47#_M1037_s N_VGND_c_2469_n 0.00437169f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_542 N_A_27_47#_M1001_g N_VGND_c_2469_n 0.0120602f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_543 N_A_27_47#_M1013_g N_VGND_c_2469_n 0.00733227f $X=8.075 $Y=0.415 $X2=0
+ $Y2=0
cc_544 N_A_27_47#_M1021_g N_VGND_c_2469_n 0.00596419f $X=11.995 $Y=0.415 $X2=0
+ $Y2=0
cc_545 N_A_27_47#_c_597_p N_VGND_c_2469_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_546 N_A_27_47#_c_339_n N_VGND_c_2469_n 0.00626967f $X=0.665 $Y=0.72 $X2=0
+ $Y2=0
cc_547 N_A_27_47#_c_342_n N_VGND_c_2469_n 0.00234902f $X=8.285 $Y=0.845 $X2=0
+ $Y2=0
cc_548 N_A_27_47#_c_343_n N_VGND_c_2469_n 0.0011282f $X=8.065 $Y=0.87 $X2=0
+ $Y2=0
cc_549 N_A_27_47#_M1001_g N_VGND_c_2470_n 0.00317372f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_550 N_A_27_47#_c_597_p N_VGND_c_2470_n 0.00895866f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_551 N_A_27_47#_c_339_n N_VGND_c_2470_n 0.0228245f $X=0.665 $Y=0.72 $X2=0
+ $Y2=0
cc_552 N_A_27_47#_c_345_n N_VGND_c_2470_n 6.84019e-19 $X=0.99 $Y=1.235 $X2=0
+ $Y2=0
cc_553 N_D_c_621_n N_A_455_324#_c_669_n 0.0474773f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_554 N_D_c_616_n N_A_455_324#_c_671_n 0.00977109f $X=1.89 $Y=1.475 $X2=0 $Y2=0
cc_555 D N_A_455_324#_c_671_n 0.00118701f $X=1.97 $Y=1.105 $X2=0 $Y2=0
cc_556 N_D_c_616_n N_A_455_324#_c_665_n 4.78431e-19 $X=1.89 $Y=1.475 $X2=0 $Y2=0
cc_557 D N_A_455_324#_c_665_n 0.00974886f $X=1.97 $Y=1.105 $X2=0 $Y2=0
cc_558 N_D_c_616_n N_A_455_324#_c_674_n 0.0043232f $X=1.89 $Y=1.475 $X2=0 $Y2=0
cc_559 D N_A_455_324#_c_674_n 0.001526f $X=1.97 $Y=1.105 $X2=0 $Y2=0
cc_560 N_D_M1043_g N_DE_M1045_g 0.0343711f $X=1.99 $Y=0.445 $X2=0 $Y2=0
cc_561 D N_DE_M1045_g 0.00266183f $X=1.97 $Y=1.105 $X2=0 $Y2=0
cc_562 N_D_c_619_n N_DE_c_766_n 0.0343711f $X=1.88 $Y=1.145 $X2=0 $Y2=0
cc_563 N_D_c_616_n DE 0.00110395f $X=1.89 $Y=1.475 $X2=0 $Y2=0
cc_564 N_D_M1043_g DE 3.92989e-19 $X=1.99 $Y=0.445 $X2=0 $Y2=0
cc_565 D DE 0.049516f $X=1.97 $Y=1.105 $X2=0 $Y2=0
cc_566 N_D_c_616_n N_A_211_363#_c_1346_n 0.00483009f $X=1.89 $Y=1.475 $X2=0
+ $Y2=0
cc_567 D N_A_211_363#_c_1346_n 0.0330428f $X=1.97 $Y=1.105 $X2=0 $Y2=0
cc_568 N_D_c_621_n N_VPWR_c_1919_n 0.00298943f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_569 N_D_c_621_n N_VPWR_c_1937_n 0.00673617f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_570 N_D_c_621_n N_VPWR_c_1917_n 0.00846956f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_571 N_D_c_616_n N_A_319_47#_c_2152_n 0.00345208f $X=1.89 $Y=1.475 $X2=0 $Y2=0
cc_572 N_D_c_621_n N_A_319_47#_c_2152_n 0.00992339f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_573 D N_A_319_47#_c_2152_n 0.00531736f $X=1.97 $Y=1.105 $X2=0 $Y2=0
cc_574 N_D_c_616_n N_A_319_47#_c_2145_n 0.00210858f $X=1.89 $Y=1.475 $X2=0 $Y2=0
cc_575 N_D_c_621_n N_A_319_47#_c_2145_n 0.00257719f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_576 N_D_M1043_g N_A_319_47#_c_2145_n 0.00680859f $X=1.99 $Y=0.445 $X2=0 $Y2=0
cc_577 D N_A_319_47#_c_2145_n 0.0722342f $X=1.97 $Y=1.105 $X2=0 $Y2=0
cc_578 N_D_c_619_n N_A_319_47#_c_2145_n 0.00771276f $X=1.88 $Y=1.145 $X2=0 $Y2=0
cc_579 N_D_M1043_g N_A_319_47#_c_2148_n 7.24971e-19 $X=1.99 $Y=0.445 $X2=0 $Y2=0
cc_580 N_D_M1043_g N_A_319_47#_c_2149_n 0.00388429f $X=1.99 $Y=0.445 $X2=0 $Y2=0
cc_581 D N_A_319_47#_c_2149_n 0.0156758f $X=1.97 $Y=1.105 $X2=0 $Y2=0
cc_582 N_D_c_619_n N_A_319_47#_c_2149_n 0.00198591f $X=1.88 $Y=1.145 $X2=0 $Y2=0
cc_583 D N_A_319_47#_c_2151_n 0.00399016f $X=1.97 $Y=1.105 $X2=0 $Y2=0
cc_584 N_D_c_619_n N_A_319_47#_c_2151_n 0.00238625f $X=1.88 $Y=1.145 $X2=0 $Y2=0
cc_585 N_D_M1043_g N_VGND_c_2446_n 0.00209795f $X=1.99 $Y=0.445 $X2=0 $Y2=0
cc_586 N_D_M1043_g N_VGND_c_2463_n 0.00585385f $X=1.99 $Y=0.445 $X2=0 $Y2=0
cc_587 N_D_M1043_g N_VGND_c_2469_n 0.00614789f $X=1.99 $Y=0.445 $X2=0 $Y2=0
cc_588 N_A_455_324#_c_664_n N_DE_M1045_g 0.00504062f $X=3.12 $Y=0.51 $X2=0 $Y2=0
cc_589 N_A_455_324#_c_665_n N_DE_c_762_n 0.005738f $X=3.132 $Y=1.355 $X2=0 $Y2=0
cc_590 N_A_455_324#_c_674_n N_DE_c_762_n 0.0080968f $X=2.78 $Y=1.52 $X2=0 $Y2=0
cc_591 N_A_455_324#_c_668_n N_DE_c_762_n 0.0178991f $X=3.132 $Y=1.01 $X2=0 $Y2=0
cc_592 N_A_455_324#_c_665_n N_DE_c_763_n 0.0181037f $X=3.132 $Y=1.355 $X2=0
+ $Y2=0
cc_593 N_A_455_324#_c_666_n N_DE_c_763_n 0.00751785f $X=3.8 $Y=1.01 $X2=0 $Y2=0
cc_594 N_A_455_324#_c_674_n N_DE_c_763_n 0.0152811f $X=2.78 $Y=1.52 $X2=0 $Y2=0
cc_595 N_A_455_324#_c_668_n N_DE_c_763_n 0.00317696f $X=3.132 $Y=1.01 $X2=0
+ $Y2=0
cc_596 N_A_455_324#_c_672_n N_DE_c_769_n 0.00953445f $X=3.12 $Y=1.99 $X2=0 $Y2=0
cc_597 N_A_455_324#_M1035_g N_DE_M1034_g 0.014951f $X=3.82 $Y=0.445 $X2=0 $Y2=0
cc_598 N_A_455_324#_c_664_n N_DE_M1034_g 0.00976426f $X=3.12 $Y=0.51 $X2=0 $Y2=0
cc_599 N_A_455_324#_c_666_n N_DE_M1034_g 0.00266577f $X=3.8 $Y=1.01 $X2=0 $Y2=0
cc_600 N_A_455_324#_c_667_n N_DE_M1034_g 0.0213613f $X=3.8 $Y=1.01 $X2=0 $Y2=0
cc_601 N_A_455_324#_c_666_n N_DE_c_770_n 0.00553997f $X=3.8 $Y=1.01 $X2=0 $Y2=0
cc_602 N_A_455_324#_c_667_n N_DE_c_770_n 0.0147305f $X=3.8 $Y=1.01 $X2=0 $Y2=0
cc_603 N_A_455_324#_c_672_n N_DE_c_771_n 5.45483e-19 $X=3.12 $Y=1.99 $X2=0 $Y2=0
cc_604 N_A_455_324#_c_666_n N_DE_c_765_n 0.00402661f $X=3.8 $Y=1.01 $X2=0 $Y2=0
cc_605 N_A_455_324#_c_668_n N_DE_c_765_n 8.39412e-19 $X=3.132 $Y=1.01 $X2=0
+ $Y2=0
cc_606 N_A_455_324#_c_672_n N_DE_c_772_n 0.00187267f $X=3.12 $Y=1.99 $X2=0 $Y2=0
cc_607 N_A_455_324#_c_665_n N_DE_c_772_n 0.00994144f $X=3.132 $Y=1.355 $X2=0
+ $Y2=0
cc_608 N_A_455_324#_c_672_n N_DE_c_773_n 2.30649e-19 $X=3.12 $Y=1.99 $X2=0 $Y2=0
cc_609 N_A_455_324#_c_665_n N_DE_c_773_n 4.99807e-19 $X=3.132 $Y=1.355 $X2=0
+ $Y2=0
cc_610 N_A_455_324#_c_671_n N_DE_c_766_n 0.00825572f $X=2.455 $Y=1.695 $X2=0
+ $Y2=0
cc_611 N_A_455_324#_c_674_n N_DE_c_766_n 0.00254194f $X=2.78 $Y=1.52 $X2=0 $Y2=0
cc_612 N_A_455_324#_c_668_n N_DE_c_766_n 6.98791e-19 $X=3.132 $Y=1.01 $X2=0
+ $Y2=0
cc_613 N_A_455_324#_c_670_n DE 0.00173211f $X=2.615 $Y=1.695 $X2=0 $Y2=0
cc_614 N_A_455_324#_c_671_n DE 0.00333636f $X=2.455 $Y=1.695 $X2=0 $Y2=0
cc_615 N_A_455_324#_c_664_n DE 0.00560441f $X=3.12 $Y=0.51 $X2=0 $Y2=0
cc_616 N_A_455_324#_c_665_n DE 0.014318f $X=3.132 $Y=1.355 $X2=0 $Y2=0
cc_617 N_A_455_324#_c_674_n DE 0.00224128f $X=2.78 $Y=1.52 $X2=0 $Y2=0
cc_618 N_A_455_324#_c_668_n DE 0.023993f $X=3.132 $Y=1.01 $X2=0 $Y2=0
cc_619 N_A_455_324#_M1035_g N_A_851_264#_M1009_g 0.0183299f $X=3.82 $Y=0.445
+ $X2=0 $Y2=0
cc_620 N_A_455_324#_c_667_n N_A_851_264#_M1009_g 0.00870265f $X=3.8 $Y=1.01
+ $X2=0 $Y2=0
cc_621 N_A_455_324#_M1035_g N_A_851_264#_c_866_n 0.00210513f $X=3.82 $Y=0.445
+ $X2=0 $Y2=0
cc_622 N_A_455_324#_c_666_n N_A_851_264#_c_866_n 0.00394871f $X=3.8 $Y=1.01
+ $X2=0 $Y2=0
cc_623 N_A_455_324#_c_667_n N_A_851_264#_c_866_n 0.00250375f $X=3.8 $Y=1.01
+ $X2=0 $Y2=0
cc_624 N_A_455_324#_M1035_g N_A_851_264#_c_867_n 0.00298582f $X=3.82 $Y=0.445
+ $X2=0 $Y2=0
cc_625 N_A_455_324#_c_666_n N_A_851_264#_c_867_n 0.0199538f $X=3.8 $Y=1.01 $X2=0
+ $Y2=0
cc_626 N_A_455_324#_c_667_n N_A_851_264#_c_867_n 0.00281276f $X=3.8 $Y=1.01
+ $X2=0 $Y2=0
cc_627 N_A_455_324#_c_671_n N_A_211_363#_c_1346_n 0.00242983f $X=2.455 $Y=1.695
+ $X2=0 $Y2=0
cc_628 N_A_455_324#_c_672_n N_A_211_363#_c_1346_n 3.18139e-19 $X=3.12 $Y=1.99
+ $X2=0 $Y2=0
cc_629 N_A_455_324#_c_665_n N_A_211_363#_c_1346_n 0.0326294f $X=3.132 $Y=1.355
+ $X2=0 $Y2=0
cc_630 N_A_455_324#_c_666_n N_A_211_363#_c_1346_n 0.0195636f $X=3.8 $Y=1.01
+ $X2=0 $Y2=0
cc_631 N_A_455_324#_c_667_n N_A_211_363#_c_1346_n 0.00256519f $X=3.8 $Y=1.01
+ $X2=0 $Y2=0
cc_632 N_A_455_324#_c_674_n N_A_211_363#_c_1346_n 0.00247375f $X=2.78 $Y=1.52
+ $X2=0 $Y2=0
cc_633 N_A_455_324#_c_669_n N_VPWR_c_1919_n 0.0201841f $X=2.365 $Y=1.77 $X2=0
+ $Y2=0
cc_634 N_A_455_324#_c_670_n N_VPWR_c_1919_n 0.00958044f $X=2.615 $Y=1.695 $X2=0
+ $Y2=0
cc_635 N_A_455_324#_c_672_n N_VPWR_c_1919_n 0.0409813f $X=3.12 $Y=1.99 $X2=0
+ $Y2=0
cc_636 N_A_455_324#_c_665_n N_VPWR_c_1919_n 0.00458578f $X=3.132 $Y=1.355 $X2=0
+ $Y2=0
cc_637 N_A_455_324#_c_672_n N_VPWR_c_1920_n 0.03428f $X=3.12 $Y=1.99 $X2=0 $Y2=0
cc_638 N_A_455_324#_c_666_n N_VPWR_c_1920_n 0.00271398f $X=3.8 $Y=1.01 $X2=0
+ $Y2=0
cc_639 N_A_455_324#_c_672_n N_VPWR_c_1930_n 0.0168164f $X=3.12 $Y=1.99 $X2=0
+ $Y2=0
cc_640 N_A_455_324#_c_669_n N_VPWR_c_1937_n 0.00427505f $X=2.365 $Y=1.77 $X2=0
+ $Y2=0
cc_641 N_A_455_324#_M1006_s N_VPWR_c_1917_n 0.00180737f $X=2.995 $Y=1.845 $X2=0
+ $Y2=0
cc_642 N_A_455_324#_c_669_n N_VPWR_c_1917_n 0.0040398f $X=2.365 $Y=1.77 $X2=0
+ $Y2=0
cc_643 N_A_455_324#_c_672_n N_VPWR_c_1917_n 0.00583478f $X=3.12 $Y=1.99 $X2=0
+ $Y2=0
cc_644 N_A_455_324#_c_669_n N_A_319_47#_c_2152_n 0.00157386f $X=2.365 $Y=1.77
+ $X2=0 $Y2=0
cc_645 N_A_455_324#_M1035_g N_A_319_47#_c_2176_n 2.12706e-19 $X=3.82 $Y=0.445
+ $X2=0 $Y2=0
cc_646 N_A_455_324#_M1034_s N_A_319_47#_c_2149_n 0.00140325f $X=2.995 $Y=0.235
+ $X2=0 $Y2=0
cc_647 N_A_455_324#_M1035_g N_A_319_47#_c_2149_n 0.00442128f $X=3.82 $Y=0.445
+ $X2=0 $Y2=0
cc_648 N_A_455_324#_c_664_n N_A_319_47#_c_2149_n 0.0182289f $X=3.12 $Y=0.51
+ $X2=0 $Y2=0
cc_649 N_A_455_324#_c_666_n N_A_319_47#_c_2149_n 0.0111442f $X=3.8 $Y=1.01 $X2=0
+ $Y2=0
cc_650 N_A_455_324#_c_667_n N_A_319_47#_c_2149_n 0.00213412f $X=3.8 $Y=1.01
+ $X2=0 $Y2=0
cc_651 N_A_455_324#_c_668_n N_A_319_47#_c_2149_n 0.00380715f $X=3.132 $Y=1.01
+ $X2=0 $Y2=0
cc_652 N_A_455_324#_M1035_g N_A_319_47#_c_2150_n 0.00251793f $X=3.82 $Y=0.445
+ $X2=0 $Y2=0
cc_653 N_A_455_324#_c_664_n N_VGND_c_2446_n 0.0165538f $X=3.12 $Y=0.51 $X2=0
+ $Y2=0
cc_654 N_A_455_324#_c_664_n N_VGND_c_2447_n 0.0157007f $X=3.12 $Y=0.51 $X2=0
+ $Y2=0
cc_655 N_A_455_324#_M1035_g N_VGND_c_2448_n 0.0130232f $X=3.82 $Y=0.445 $X2=0
+ $Y2=0
cc_656 N_A_455_324#_c_664_n N_VGND_c_2448_n 0.0241012f $X=3.12 $Y=0.51 $X2=0
+ $Y2=0
cc_657 N_A_455_324#_c_666_n N_VGND_c_2448_n 0.0179132f $X=3.8 $Y=1.01 $X2=0
+ $Y2=0
cc_658 N_A_455_324#_c_667_n N_VGND_c_2448_n 0.00159308f $X=3.8 $Y=1.01 $X2=0
+ $Y2=0
cc_659 N_A_455_324#_M1035_g N_VGND_c_2464_n 0.00505556f $X=3.82 $Y=0.445 $X2=0
+ $Y2=0
cc_660 N_A_455_324#_M1034_s N_VGND_c_2469_n 0.00156059f $X=2.995 $Y=0.235 $X2=0
+ $Y2=0
cc_661 N_A_455_324#_M1035_g N_VGND_c_2469_n 0.0039983f $X=3.82 $Y=0.445 $X2=0
+ $Y2=0
cc_662 N_A_455_324#_c_664_n N_VGND_c_2469_n 0.00215984f $X=3.12 $Y=0.51 $X2=0
+ $Y2=0
cc_663 N_DE_c_771_n N_A_851_264#_c_869_n 0.0270745f $X=3.845 $Y=1.77 $X2=0 $Y2=0
cc_664 N_DE_c_773_n N_A_851_264#_c_869_n 0.0130125f $X=3.845 $Y=1.535 $X2=0
+ $Y2=0
cc_665 N_DE_c_763_n N_A_851_264#_c_876_n 0.00332959f $X=3.355 $Y=1.46 $X2=0
+ $Y2=0
cc_666 N_DE_c_773_n N_A_851_264#_c_876_n 0.00395406f $X=3.845 $Y=1.535 $X2=0
+ $Y2=0
cc_667 N_DE_c_763_n N_A_851_264#_c_867_n 0.00312649f $X=3.355 $Y=1.46 $X2=0
+ $Y2=0
cc_668 N_DE_c_770_n N_A_211_363#_c_1346_n 0.0033956f $X=3.745 $Y=1.535 $X2=0
+ $Y2=0
cc_669 N_DE_c_772_n N_A_211_363#_c_1346_n 0.00384371f $X=3.355 $Y=1.535 $X2=0
+ $Y2=0
cc_670 N_DE_c_773_n N_A_211_363#_c_1346_n 0.00469043f $X=3.845 $Y=1.535 $X2=0
+ $Y2=0
cc_671 N_DE_c_766_n N_A_211_363#_c_1346_n 7.08986e-19 $X=2.655 $Y=0.992 $X2=0
+ $Y2=0
cc_672 DE N_A_211_363#_c_1346_n 0.0162302f $X=2.515 $Y=0.95 $X2=0 $Y2=0
cc_673 N_DE_c_769_n N_VPWR_c_1919_n 0.00294979f $X=3.355 $Y=1.77 $X2=0 $Y2=0
cc_674 DE N_VPWR_c_1919_n 0.00211801f $X=2.515 $Y=0.95 $X2=0 $Y2=0
cc_675 N_DE_c_769_n N_VPWR_c_1920_n 0.00603594f $X=3.355 $Y=1.77 $X2=0 $Y2=0
cc_676 N_DE_c_770_n N_VPWR_c_1920_n 0.00424078f $X=3.745 $Y=1.535 $X2=0 $Y2=0
cc_677 N_DE_c_771_n N_VPWR_c_1920_n 0.00406636f $X=3.845 $Y=1.77 $X2=0 $Y2=0
cc_678 N_DE_c_769_n N_VPWR_c_1930_n 0.00674661f $X=3.355 $Y=1.77 $X2=0 $Y2=0
cc_679 N_DE_c_771_n N_VPWR_c_1938_n 0.00702461f $X=3.845 $Y=1.77 $X2=0 $Y2=0
cc_680 N_DE_c_769_n N_VPWR_c_1917_n 0.00853099f $X=3.355 $Y=1.77 $X2=0 $Y2=0
cc_681 N_DE_c_771_n N_VPWR_c_1917_n 0.00761288f $X=3.845 $Y=1.77 $X2=0 $Y2=0
cc_682 N_DE_c_771_n N_A_319_47#_c_2154_n 0.00340986f $X=3.845 $Y=1.77 $X2=0
+ $Y2=0
cc_683 N_DE_M1045_g N_A_319_47#_c_2149_n 0.00479706f $X=2.35 $Y=0.445 $X2=0
+ $Y2=0
cc_684 N_DE_c_762_n N_A_319_47#_c_2149_n 0.00452289f $X=3.255 $Y=0.925 $X2=0
+ $Y2=0
cc_685 N_DE_M1034_g N_A_319_47#_c_2149_n 0.00130833f $X=3.38 $Y=0.445 $X2=0
+ $Y2=0
cc_686 DE N_A_319_47#_c_2149_n 0.0132392f $X=2.515 $Y=0.95 $X2=0 $Y2=0
cc_687 N_DE_M1045_g N_VGND_c_2446_n 0.0112128f $X=2.35 $Y=0.445 $X2=0 $Y2=0
cc_688 N_DE_c_762_n N_VGND_c_2446_n 5.49262e-19 $X=3.255 $Y=0.925 $X2=0 $Y2=0
cc_689 N_DE_M1034_g N_VGND_c_2446_n 0.00184778f $X=3.38 $Y=0.445 $X2=0 $Y2=0
cc_690 N_DE_c_766_n N_VGND_c_2446_n 0.00120611f $X=2.655 $Y=0.992 $X2=0 $Y2=0
cc_691 DE N_VGND_c_2446_n 0.0170561f $X=2.515 $Y=0.95 $X2=0 $Y2=0
cc_692 N_DE_M1034_g N_VGND_c_2447_n 0.00310428f $X=3.38 $Y=0.445 $X2=0 $Y2=0
cc_693 N_DE_M1034_g N_VGND_c_2448_n 0.0111028f $X=3.38 $Y=0.445 $X2=0 $Y2=0
cc_694 N_DE_M1045_g N_VGND_c_2463_n 0.00427505f $X=2.35 $Y=0.445 $X2=0 $Y2=0
cc_695 N_DE_M1045_g N_VGND_c_2469_n 0.00301124f $X=2.35 $Y=0.445 $X2=0 $Y2=0
cc_696 N_DE_M1034_g N_VGND_c_2469_n 0.00381833f $X=3.38 $Y=0.445 $X2=0 $Y2=0
cc_697 N_A_851_264#_M1009_g N_A_955_21#_c_1083_n 0.0204071f $X=4.43 $Y=0.445
+ $X2=0 $Y2=0
cc_698 N_A_851_264#_c_865_n N_A_955_21#_c_1084_n 0.00846539f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_699 N_A_851_264#_c_865_n N_A_955_21#_c_1085_n 0.00395832f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_700 N_A_851_264#_c_865_n N_A_955_21#_c_1088_n 0.00285622f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_701 N_A_851_264#_c_865_n N_A_955_21#_c_1092_n 0.00443266f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_702 N_A_851_264#_c_865_n N_A_955_21#_c_1093_n 0.0229786f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_703 N_A_851_264#_c_865_n N_SCD_M1038_g 0.00388453f $X=14.385 $Y=0.85 $X2=0
+ $Y2=0
cc_704 N_A_851_264#_c_865_n SCD 0.0113481f $X=14.385 $Y=0.85 $X2=0 $Y2=0
cc_705 N_A_851_264#_c_869_n N_SCE_c_1248_n 0.00823699f $X=4.405 $Y=1.77
+ $X2=-0.19 $Y2=-0.24
cc_706 N_A_851_264#_c_865_n N_SCE_M1015_g 0.00310007f $X=14.385 $Y=0.85 $X2=0
+ $Y2=0
cc_707 N_A_851_264#_c_865_n N_SCE_M1024_g 0.00427016f $X=14.385 $Y=0.85 $X2=0
+ $Y2=0
cc_708 N_A_851_264#_c_869_n N_SCE_c_1251_n 0.0169332f $X=4.405 $Y=1.77 $X2=0
+ $Y2=0
cc_709 N_A_851_264#_c_876_n N_SCE_c_1251_n 2.79151e-19 $X=4.39 $Y=1.485 $X2=0
+ $Y2=0
cc_710 N_A_851_264#_c_865_n N_SCE_c_1251_n 0.00280829f $X=14.385 $Y=0.85 $X2=0
+ $Y2=0
cc_711 N_A_851_264#_c_865_n SCE 0.00498401f $X=14.385 $Y=0.85 $X2=0 $Y2=0
cc_712 N_A_851_264#_c_865_n N_SCE_c_1247_n 3.73597e-19 $X=14.385 $Y=0.85 $X2=0
+ $Y2=0
cc_713 N_A_851_264#_c_865_n N_A_211_363#_c_1333_n 0.00111623f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_714 N_A_851_264#_c_865_n N_A_211_363#_M1042_g 0.00533369f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_715 N_A_851_264#_c_852_n N_A_211_363#_c_1345_n 0.0133138f $X=12.38 $Y=1.89
+ $X2=0 $Y2=0
cc_716 N_A_851_264#_c_872_n N_A_211_363#_c_1345_n 0.014514f $X=12.38 $Y=1.99
+ $X2=0 $Y2=0
cc_717 N_A_851_264#_c_865_n N_A_211_363#_c_1336_n 0.033982f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_718 N_A_851_264#_c_865_n N_A_211_363#_c_1337_n 0.00490197f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_719 N_A_851_264#_c_869_n N_A_211_363#_c_1346_n 0.00127021f $X=4.405 $Y=1.77
+ $X2=0 $Y2=0
cc_720 N_A_851_264#_c_876_n N_A_211_363#_c_1346_n 0.0232082f $X=4.39 $Y=1.485
+ $X2=0 $Y2=0
cc_721 N_A_851_264#_c_865_n N_A_211_363#_c_1346_n 0.150485f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_722 N_A_851_264#_c_866_n N_A_211_363#_c_1346_n 0.0132881f $X=4.335 $Y=0.85
+ $X2=0 $Y2=0
cc_723 N_A_851_264#_c_867_n N_A_211_363#_c_1346_n 3.15466e-19 $X=4.19 $Y=0.85
+ $X2=0 $Y2=0
cc_724 N_A_851_264#_c_865_n N_A_211_363#_c_1348_n 0.14356f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_725 N_A_851_264#_c_865_n N_A_211_363#_c_1349_n 0.0152007f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_726 N_A_851_264#_c_865_n N_A_211_363#_c_1397_n 0.0143644f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_727 N_A_851_264#_c_852_n N_A_211_363#_c_1338_n 0.00179343f $X=12.38 $Y=1.89
+ $X2=0 $Y2=0
cc_728 N_A_851_264#_c_865_n N_A_211_363#_c_1339_n 0.00135618f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_729 N_A_851_264#_c_865_n N_A_211_363#_c_1340_n 0.00127009f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_730 N_A_851_264#_c_865_n N_A_1787_159#_M1010_g 0.00591182f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_731 N_A_851_264#_c_865_n N_A_1787_159#_c_1550_n 0.00757538f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_732 N_A_851_264#_c_865_n N_A_1787_159#_c_1552_n 0.0600767f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_733 N_A_851_264#_c_865_n N_A_1787_159#_c_1554_n 0.012477f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_734 N_A_851_264#_c_865_n N_A_1787_159#_c_1556_n 0.0137823f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_735 N_A_851_264#_c_865_n N_A_1787_159#_c_1557_n 0.00300541f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_736 N_A_851_264#_c_865_n N_A_1611_413#_c_1691_n 0.00826559f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_737 N_A_851_264#_c_865_n N_A_1611_413#_c_1677_n 0.0155494f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_738 N_A_851_264#_c_865_n N_A_1611_413#_c_1678_n 0.00637281f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_739 N_A_851_264#_c_862_n N_A_2266_413#_c_1788_n 0.0249886f $X=14.52 $Y=1.99
+ $X2=0 $Y2=0
cc_740 N_A_851_264#_c_863_n N_A_2266_413#_c_1788_n 0.0118216f $X=14.155 $Y=1.055
+ $X2=0 $Y2=0
cc_741 N_A_851_264#_c_864_n N_A_2266_413#_c_1788_n 0.00378647f $X=14.525
+ $Y=1.055 $X2=0 $Y2=0
cc_742 N_A_851_264#_c_863_n N_A_2266_413#_M1018_g 0.0101663f $X=14.155 $Y=1.055
+ $X2=0 $Y2=0
cc_743 N_A_851_264#_c_864_n N_A_2266_413#_M1018_g 0.00355346f $X=14.525 $Y=1.055
+ $X2=0 $Y2=0
cc_744 N_A_851_264#_c_868_n N_A_2266_413#_M1018_g 0.0141022f $X=14.53 $Y=0.385
+ $X2=0 $Y2=0
cc_745 N_A_851_264#_c_862_n N_A_2266_413#_c_1789_n 0.00940588f $X=14.52 $Y=1.99
+ $X2=0 $Y2=0
cc_746 N_A_851_264#_c_862_n N_A_2266_413#_c_1783_n 0.0164317f $X=14.52 $Y=1.99
+ $X2=0 $Y2=0
cc_747 N_A_851_264#_c_864_n N_A_2266_413#_c_1783_n 0.0107146f $X=14.525 $Y=1.055
+ $X2=0 $Y2=0
cc_748 N_A_851_264#_c_864_n N_A_2266_413#_c_1784_n 2.95806e-19 $X=14.525
+ $Y=1.055 $X2=0 $Y2=0
cc_749 N_A_851_264#_c_862_n N_A_2266_413#_c_1792_n 4.30725e-19 $X=14.52 $Y=1.99
+ $X2=0 $Y2=0
cc_750 N_A_851_264#_c_862_n N_A_2266_413#_c_1786_n 2.53909e-19 $X=14.52 $Y=1.99
+ $X2=0 $Y2=0
cc_751 N_A_851_264#_c_872_n N_A_2266_413#_c_1801_n 0.00754404f $X=12.38 $Y=1.99
+ $X2=0 $Y2=0
cc_752 N_A_851_264#_c_865_n N_A_2266_413#_c_1805_n 0.00756627f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_753 N_A_851_264#_c_852_n N_A_2266_413#_c_1795_n 0.00412925f $X=12.38 $Y=1.89
+ $X2=0 $Y2=0
cc_754 N_A_851_264#_c_872_n N_A_2266_413#_c_1795_n 0.00170274f $X=12.38 $Y=1.99
+ $X2=0 $Y2=0
cc_755 N_A_851_264#_c_854_n N_A_2266_413#_c_1795_n 5.69782e-19 $X=12.815
+ $Y=1.127 $X2=0 $Y2=0
cc_756 N_A_851_264#_c_855_n N_A_2266_413#_c_1795_n 0.00654381f $X=12.915 $Y=1.41
+ $X2=0 $Y2=0
cc_757 N_A_851_264#_c_858_n N_A_2266_413#_c_1795_n 0.00991573f $X=13.385 $Y=1.41
+ $X2=0 $Y2=0
cc_758 N_A_851_264#_c_852_n N_A_2266_413#_c_1796_n 0.00128524f $X=12.38 $Y=1.89
+ $X2=0 $Y2=0
cc_759 N_A_851_264#_c_872_n N_A_2266_413#_c_1796_n 7.1525e-19 $X=12.38 $Y=1.99
+ $X2=0 $Y2=0
cc_760 N_A_851_264#_c_852_n N_A_2266_413#_c_1787_n 0.0200266f $X=12.38 $Y=1.89
+ $X2=0 $Y2=0
cc_761 N_A_851_264#_c_872_n N_A_2266_413#_c_1787_n 0.00753412f $X=12.38 $Y=1.99
+ $X2=0 $Y2=0
cc_762 N_A_851_264#_M1004_g N_A_2266_413#_c_1787_n 0.00648134f $X=12.47 $Y=0.445
+ $X2=0 $Y2=0
cc_763 N_A_851_264#_c_855_n N_A_2266_413#_c_1787_n 0.00118373f $X=12.915 $Y=1.41
+ $X2=0 $Y2=0
cc_764 N_A_851_264#_c_861_n N_A_2266_413#_c_1787_n 0.0104811f $X=12.412 $Y=1.127
+ $X2=0 $Y2=0
cc_765 N_A_851_264#_c_865_n N_A_2266_413#_c_1787_n 0.0253607f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_766 N_A_851_264#_c_860_n N_A_2266_413#_c_1798_n 3.4957e-19 $X=14.02 $Y=1.127
+ $X2=0 $Y2=0
cc_767 N_A_851_264#_c_862_n N_A_2266_413#_c_1798_n 0.00757769f $X=14.52 $Y=1.99
+ $X2=0 $Y2=0
cc_768 N_A_851_264#_c_864_n N_A_2266_413#_c_1798_n 0.00147962f $X=14.525
+ $Y=1.055 $X2=0 $Y2=0
cc_769 N_A_851_264#_c_858_n N_A_2266_413#_c_1799_n 0.00638217f $X=13.385 $Y=1.41
+ $X2=0 $Y2=0
cc_770 N_A_851_264#_c_860_n N_A_2266_413#_c_1799_n 0.0118216f $X=14.02 $Y=1.127
+ $X2=0 $Y2=0
cc_771 N_A_851_264#_c_862_n N_A_2266_413#_c_1799_n 0.0019835f $X=14.52 $Y=1.99
+ $X2=0 $Y2=0
cc_772 N_A_851_264#_c_864_n N_A_2266_413#_c_1799_n 0.00120686f $X=14.525
+ $Y=1.055 $X2=0 $Y2=0
cc_773 N_A_851_264#_c_865_n N_A_2266_413#_c_1799_n 2.03294e-19 $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_774 N_A_851_264#_c_860_n N_A_2266_413#_c_1800_n 8.89189e-19 $X=14.02 $Y=1.127
+ $X2=0 $Y2=0
cc_775 N_A_851_264#_c_862_n N_A_2266_413#_c_1800_n 0.0310392f $X=14.52 $Y=1.99
+ $X2=0 $Y2=0
cc_776 N_A_851_264#_c_864_n N_A_2266_413#_c_1800_n 0.00423209f $X=14.525
+ $Y=1.055 $X2=0 $Y2=0
cc_777 N_A_851_264#_c_852_n N_VPWR_c_1925_n 0.00368287f $X=12.38 $Y=1.89 $X2=0
+ $Y2=0
cc_778 N_A_851_264#_c_872_n N_VPWR_c_1925_n 0.00817671f $X=12.38 $Y=1.99 $X2=0
+ $Y2=0
cc_779 N_A_851_264#_c_854_n N_VPWR_c_1925_n 0.00373031f $X=12.815 $Y=1.127 $X2=0
+ $Y2=0
cc_780 N_A_851_264#_c_855_n N_VPWR_c_1925_n 0.00572061f $X=12.915 $Y=1.41 $X2=0
+ $Y2=0
cc_781 N_A_851_264#_c_865_n N_VPWR_c_1925_n 0.00406719f $X=14.385 $Y=0.85 $X2=0
+ $Y2=0
cc_782 N_A_851_264#_c_855_n N_VPWR_c_1926_n 0.00597712f $X=12.915 $Y=1.41 $X2=0
+ $Y2=0
cc_783 N_A_851_264#_c_858_n N_VPWR_c_1926_n 0.00673617f $X=13.385 $Y=1.41 $X2=0
+ $Y2=0
cc_784 N_A_851_264#_c_858_n N_VPWR_c_1927_n 0.0163679f $X=13.385 $Y=1.41 $X2=0
+ $Y2=0
cc_785 N_A_851_264#_c_862_n N_VPWR_c_1927_n 0.0194681f $X=14.52 $Y=1.99 $X2=0
+ $Y2=0
cc_786 N_A_851_264#_c_865_n N_VPWR_c_1927_n 0.00706095f $X=14.385 $Y=0.85 $X2=0
+ $Y2=0
cc_787 N_A_851_264#_c_862_n N_VPWR_c_1928_n 0.0627047f $X=14.52 $Y=1.99 $X2=0
+ $Y2=0
cc_788 N_A_851_264#_c_869_n N_VPWR_c_1938_n 0.00597712f $X=4.405 $Y=1.77 $X2=0
+ $Y2=0
cc_789 N_A_851_264#_c_872_n N_VPWR_c_1939_n 0.00609153f $X=12.38 $Y=1.99 $X2=0
+ $Y2=0
cc_790 N_A_851_264#_c_862_n N_VPWR_c_1940_n 0.0217628f $X=14.52 $Y=1.99 $X2=0
+ $Y2=0
cc_791 N_A_851_264#_M1005_s N_VPWR_c_1917_n 0.00225715f $X=14.395 $Y=1.845 $X2=0
+ $Y2=0
cc_792 N_A_851_264#_c_869_n N_VPWR_c_1917_n 0.00725925f $X=4.405 $Y=1.77 $X2=0
+ $Y2=0
cc_793 N_A_851_264#_c_872_n N_VPWR_c_1917_n 0.00759045f $X=12.38 $Y=1.99 $X2=0
+ $Y2=0
cc_794 N_A_851_264#_c_855_n N_VPWR_c_1917_n 0.00691969f $X=12.915 $Y=1.41 $X2=0
+ $Y2=0
cc_795 N_A_851_264#_c_858_n N_VPWR_c_1917_n 0.00845433f $X=13.385 $Y=1.41 $X2=0
+ $Y2=0
cc_796 N_A_851_264#_c_862_n N_VPWR_c_1917_n 0.0128576f $X=14.52 $Y=1.99 $X2=0
+ $Y2=0
cc_797 N_A_851_264#_c_869_n N_A_319_47#_c_2154_n 0.0191483f $X=4.405 $Y=1.77
+ $X2=0 $Y2=0
cc_798 N_A_851_264#_c_876_n N_A_319_47#_c_2154_n 0.00639471f $X=4.39 $Y=1.485
+ $X2=0 $Y2=0
cc_799 N_A_851_264#_c_869_n N_A_319_47#_c_2146_n 0.00620991f $X=4.405 $Y=1.77
+ $X2=0 $Y2=0
cc_800 N_A_851_264#_M1009_g N_A_319_47#_c_2146_n 0.00253365f $X=4.43 $Y=0.445
+ $X2=0 $Y2=0
cc_801 N_A_851_264#_c_876_n N_A_319_47#_c_2146_n 0.0240379f $X=4.39 $Y=1.485
+ $X2=0 $Y2=0
cc_802 N_A_851_264#_c_867_n N_A_319_47#_c_2146_n 0.00481225f $X=4.19 $Y=0.85
+ $X2=0 $Y2=0
cc_803 N_A_851_264#_c_869_n N_A_319_47#_c_2147_n 0.00197416f $X=4.405 $Y=1.77
+ $X2=0 $Y2=0
cc_804 N_A_851_264#_M1009_g N_A_319_47#_c_2147_n 0.00656396f $X=4.43 $Y=0.445
+ $X2=0 $Y2=0
cc_805 N_A_851_264#_c_876_n N_A_319_47#_c_2147_n 0.00565f $X=4.39 $Y=1.485 $X2=0
+ $Y2=0
cc_806 N_A_851_264#_c_865_n N_A_319_47#_c_2147_n 0.00430154f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_807 N_A_851_264#_M1009_g N_A_319_47#_c_2176_n 0.00114831f $X=4.43 $Y=0.445
+ $X2=0 $Y2=0
cc_808 N_A_851_264#_c_865_n N_A_319_47#_c_2176_n 0.0293733f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_809 N_A_851_264#_M1009_g N_A_319_47#_c_2149_n 0.00282075f $X=4.43 $Y=0.445
+ $X2=0 $Y2=0
cc_810 N_A_851_264#_c_865_n N_A_319_47#_c_2149_n 0.00739417f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_811 N_A_851_264#_c_866_n N_A_319_47#_c_2149_n 0.0273854f $X=4.335 $Y=0.85
+ $X2=0 $Y2=0
cc_812 N_A_851_264#_c_867_n N_A_319_47#_c_2149_n 0.00264974f $X=4.19 $Y=0.85
+ $X2=0 $Y2=0
cc_813 N_A_851_264#_M1009_g N_A_319_47#_c_2150_n 0.0177941f $X=4.43 $Y=0.445
+ $X2=0 $Y2=0
cc_814 N_A_851_264#_c_865_n N_A_319_47#_c_2150_n 0.0200579f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_815 N_A_851_264#_c_866_n N_A_319_47#_c_2150_n 0.0027459f $X=4.335 $Y=0.85
+ $X2=0 $Y2=0
cc_816 N_A_851_264#_c_867_n N_A_319_47#_c_2150_n 0.0331876f $X=4.19 $Y=0.85
+ $X2=0 $Y2=0
cc_817 N_A_851_264#_c_865_n N_A_985_47#_M1024_d 0.00303818f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_818 N_A_851_264#_c_865_n N_A_985_47#_c_2260_n 0.027397f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_819 N_A_851_264#_c_865_n N_A_985_47#_c_2261_n 0.00745895f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_820 N_A_851_264#_M1009_g N_A_985_47#_c_2262_n 0.00169605f $X=4.43 $Y=0.445
+ $X2=0 $Y2=0
cc_821 N_A_851_264#_c_865_n N_A_985_47#_c_2262_n 0.0100836f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_822 N_A_851_264#_c_865_n N_A_985_47#_c_2265_n 0.0301322f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_823 N_A_851_264#_c_865_n N_A_985_47#_c_2266_n 0.0299403f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_824 N_A_851_264#_c_865_n N_A_985_47#_c_2267_n 0.158651f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_825 N_A_851_264#_c_865_n N_A_985_47#_c_2268_n 0.00623535f $X=14.385 $Y=0.85
+ $X2=0 $Y2=0
cc_826 N_A_851_264#_c_865_n N_Q_N_M1017_s 2.55492e-19 $X=14.385 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_827 N_A_851_264#_c_855_n N_Q_N_c_2398_n 0.0205156f $X=12.915 $Y=1.41 $X2=0
+ $Y2=0
cc_828 N_A_851_264#_c_858_n N_Q_N_c_2398_n 0.0206869f $X=13.385 $Y=1.41 $X2=0
+ $Y2=0
cc_829 N_A_851_264#_M1017_g N_Q_N_c_2396_n 0.00409836f $X=13.005 $Y=0.56 $X2=0
+ $Y2=0
cc_830 N_A_851_264#_c_857_n N_Q_N_c_2396_n 0.00472753f $X=13.285 $Y=1.127 $X2=0
+ $Y2=0
cc_831 N_A_851_264#_c_858_n N_Q_N_c_2396_n 0.00186059f $X=13.385 $Y=1.41 $X2=0
+ $Y2=0
cc_832 N_A_851_264#_M1033_g N_Q_N_c_2396_n 0.0119689f $X=13.475 $Y=0.56 $X2=0
+ $Y2=0
cc_833 N_A_851_264#_c_863_n N_Q_N_c_2396_n 4.62445e-19 $X=14.155 $Y=1.055 $X2=0
+ $Y2=0
cc_834 N_A_851_264#_c_864_n N_Q_N_c_2396_n 0.00812593f $X=14.525 $Y=1.055 $X2=0
+ $Y2=0
cc_835 N_A_851_264#_c_865_n N_Q_N_c_2396_n 0.0315548f $X=14.385 $Y=0.85 $X2=0
+ $Y2=0
cc_836 N_A_851_264#_c_852_n Q_N 0.00105285f $X=12.38 $Y=1.89 $X2=0 $Y2=0
cc_837 N_A_851_264#_c_855_n Q_N 0.0117602f $X=12.915 $Y=1.41 $X2=0 $Y2=0
cc_838 N_A_851_264#_c_857_n Q_N 0.00554273f $X=13.285 $Y=1.127 $X2=0 $Y2=0
cc_839 N_A_851_264#_c_858_n Q_N 0.0150068f $X=13.385 $Y=1.41 $X2=0 $Y2=0
cc_840 N_A_851_264#_c_865_n Q_N 0.00763366f $X=14.385 $Y=0.85 $X2=0 $Y2=0
cc_841 N_A_851_264#_c_862_n N_Q_c_2426_n 0.00630592f $X=14.52 $Y=1.99 $X2=0
+ $Y2=0
cc_842 N_A_851_264#_c_864_n N_Q_c_2426_n 0.00861483f $X=14.525 $Y=1.055 $X2=0
+ $Y2=0
cc_843 N_A_851_264#_c_865_n N_VGND_M1015_d 0.00436703f $X=14.385 $Y=0.85 $X2=0
+ $Y2=0
cc_844 N_A_851_264#_c_865_n N_VGND_M1004_d 6.81311e-19 $X=14.385 $Y=0.85 $X2=0
+ $Y2=0
cc_845 N_A_851_264#_c_865_n N_VGND_M1033_d 0.0014194f $X=14.385 $Y=0.85 $X2=0
+ $Y2=0
cc_846 N_A_851_264#_M1009_g N_VGND_c_2448_n 0.00274629f $X=4.43 $Y=0.445 $X2=0
+ $Y2=0
cc_847 N_A_851_264#_c_865_n N_VGND_c_2449_n 0.0125025f $X=14.385 $Y=0.85 $X2=0
+ $Y2=0
cc_848 N_A_851_264#_c_865_n N_VGND_c_2450_n 0.00212198f $X=14.385 $Y=0.85 $X2=0
+ $Y2=0
cc_849 N_A_851_264#_c_865_n N_VGND_c_2451_n 0.00455022f $X=14.385 $Y=0.85 $X2=0
+ $Y2=0
cc_850 N_A_851_264#_M1004_g N_VGND_c_2452_n 0.0102933f $X=12.47 $Y=0.445 $X2=0
+ $Y2=0
cc_851 N_A_851_264#_c_854_n N_VGND_c_2452_n 0.00667183f $X=12.815 $Y=1.127 $X2=0
+ $Y2=0
cc_852 N_A_851_264#_M1017_g N_VGND_c_2452_n 0.00324684f $X=13.005 $Y=0.56 $X2=0
+ $Y2=0
cc_853 N_A_851_264#_c_865_n N_VGND_c_2452_n 0.0171232f $X=14.385 $Y=0.85 $X2=0
+ $Y2=0
cc_854 N_A_851_264#_M1033_g N_VGND_c_2453_n 0.00676439f $X=13.475 $Y=0.56 $X2=0
+ $Y2=0
cc_855 N_A_851_264#_c_860_n N_VGND_c_2453_n 0.00742348f $X=14.02 $Y=1.127 $X2=0
+ $Y2=0
cc_856 N_A_851_264#_c_864_n N_VGND_c_2453_n 6.20383e-19 $X=14.525 $Y=1.055 $X2=0
+ $Y2=0
cc_857 N_A_851_264#_c_865_n N_VGND_c_2453_n 0.0177642f $X=14.385 $Y=0.85 $X2=0
+ $Y2=0
cc_858 N_A_851_264#_c_1063_p N_VGND_c_2453_n 2.98782e-19 $X=14.53 $Y=0.85 $X2=0
+ $Y2=0
cc_859 N_A_851_264#_c_868_n N_VGND_c_2453_n 0.0242201f $X=14.53 $Y=0.385 $X2=0
+ $Y2=0
cc_860 N_A_851_264#_c_864_n N_VGND_c_2454_n 5.29946e-19 $X=14.525 $Y=1.055 $X2=0
+ $Y2=0
cc_861 N_A_851_264#_c_1063_p N_VGND_c_2454_n 0.00115041f $X=14.53 $Y=0.85 $X2=0
+ $Y2=0
cc_862 N_A_851_264#_c_868_n N_VGND_c_2454_n 0.0385837f $X=14.53 $Y=0.385 $X2=0
+ $Y2=0
cc_863 N_A_851_264#_M1017_g N_VGND_c_2458_n 0.00585385f $X=13.005 $Y=0.56 $X2=0
+ $Y2=0
cc_864 N_A_851_264#_M1033_g N_VGND_c_2458_n 0.00541359f $X=13.475 $Y=0.56 $X2=0
+ $Y2=0
cc_865 N_A_851_264#_M1009_g N_VGND_c_2464_n 0.00495816f $X=4.43 $Y=0.445 $X2=0
+ $Y2=0
cc_866 N_A_851_264#_c_867_n N_VGND_c_2464_n 0.00260398f $X=4.19 $Y=0.85 $X2=0
+ $Y2=0
cc_867 N_A_851_264#_M1004_g N_VGND_c_2466_n 0.00585385f $X=12.47 $Y=0.445 $X2=0
+ $Y2=0
cc_868 N_A_851_264#_c_868_n N_VGND_c_2467_n 0.021656f $X=14.53 $Y=0.385 $X2=0
+ $Y2=0
cc_869 N_A_851_264#_M1018_s N_VGND_c_2469_n 0.00166412f $X=14.405 $Y=0.235 $X2=0
+ $Y2=0
cc_870 N_A_851_264#_M1009_g N_VGND_c_2469_n 0.0055221f $X=4.43 $Y=0.445 $X2=0
+ $Y2=0
cc_871 N_A_851_264#_M1004_g N_VGND_c_2469_n 0.00685062f $X=12.47 $Y=0.445 $X2=0
+ $Y2=0
cc_872 N_A_851_264#_M1017_g N_VGND_c_2469_n 0.00662332f $X=13.005 $Y=0.56 $X2=0
+ $Y2=0
cc_873 N_A_851_264#_M1033_g N_VGND_c_2469_n 0.00756836f $X=13.475 $Y=0.56 $X2=0
+ $Y2=0
cc_874 N_A_851_264#_c_865_n N_VGND_c_2469_n 0.331019f $X=14.385 $Y=0.85 $X2=0
+ $Y2=0
cc_875 N_A_851_264#_c_1063_p N_VGND_c_2469_n 0.014516f $X=14.53 $Y=0.85 $X2=0
+ $Y2=0
cc_876 N_A_851_264#_c_868_n N_VGND_c_2469_n 0.00617083f $X=14.53 $Y=0.385 $X2=0
+ $Y2=0
cc_877 N_A_851_264#_c_865_n A_1373_119# 0.00414878f $X=14.385 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_878 N_A_955_21#_c_1087_n N_SCD_c_1201_n 0.0542844f $X=7.32 $Y=1.77 $X2=-0.19
+ $Y2=-0.24
cc_879 N_A_955_21#_c_1091_n N_SCD_c_1201_n 0.00134654f $X=6.14 $Y=1.835
+ $X2=-0.19 $Y2=-0.24
cc_880 N_A_955_21#_c_1096_n N_SCD_c_1201_n 0.0169246f $X=7.12 $Y=1.92 $X2=-0.19
+ $Y2=-0.24
cc_881 N_A_955_21#_c_1092_n N_SCD_c_1201_n 0.0035277f $X=7.235 $Y=1.52 $X2=-0.19
+ $Y2=-0.24
cc_882 N_A_955_21#_c_1098_n N_SCD_c_1201_n 8.24051e-19 $X=5.955 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_883 N_A_955_21#_c_1090_n N_SCD_M1038_g 0.00109976f $X=6.06 $Y=0.75 $X2=0
+ $Y2=0
cc_884 N_A_955_21#_c_1087_n SCD 0.00166333f $X=7.32 $Y=1.77 $X2=0 $Y2=0
cc_885 N_A_955_21#_c_1091_n SCD 0.034515f $X=6.14 $Y=1.835 $X2=0 $Y2=0
cc_886 N_A_955_21#_c_1096_n SCD 0.0344424f $X=7.12 $Y=1.92 $X2=0 $Y2=0
cc_887 N_A_955_21#_c_1092_n SCD 0.0233244f $X=7.235 $Y=1.52 $X2=0 $Y2=0
cc_888 N_A_955_21#_c_1084_n N_SCE_c_1241_n 0.0087278f $X=5.63 $Y=0.84 $X2=0
+ $Y2=0
cc_889 N_A_955_21#_c_1091_n N_SCE_c_1250_n 0.00320653f $X=6.14 $Y=1.835 $X2=0
+ $Y2=0
cc_890 N_A_955_21#_c_1096_n N_SCE_c_1250_n 0.00647449f $X=7.12 $Y=1.92 $X2=0
+ $Y2=0
cc_891 N_A_955_21#_c_1098_n N_SCE_c_1250_n 0.0117419f $X=5.955 $Y=2 $X2=0 $Y2=0
cc_892 N_A_955_21#_c_1086_n N_SCE_M1015_g 0.00660962f $X=5.705 $Y=0.765 $X2=0
+ $Y2=0
cc_893 N_A_955_21#_c_1088_n N_SCE_M1015_g 0.00589644f $X=5.895 $Y=0.385 $X2=0
+ $Y2=0
cc_894 N_A_955_21#_c_1090_n N_SCE_M1015_g 0.00377036f $X=6.06 $Y=0.75 $X2=0
+ $Y2=0
cc_895 N_A_955_21#_c_1091_n N_SCE_M1015_g 0.00575433f $X=6.14 $Y=1.835 $X2=0
+ $Y2=0
cc_896 N_A_955_21#_c_1093_n N_SCE_M1015_g 0.00174526f $X=6.06 $Y=0.935 $X2=0
+ $Y2=0
cc_897 N_A_955_21#_c_1088_n N_SCE_c_1244_n 2.57001e-19 $X=5.895 $Y=0.385 $X2=0
+ $Y2=0
cc_898 N_A_955_21#_c_1089_n N_SCE_c_1244_n 0.0145232f $X=5.765 $Y=0.34 $X2=0
+ $Y2=0
cc_899 N_A_955_21#_c_1087_n N_SCE_M1024_g 0.00852628f $X=7.32 $Y=1.77 $X2=0
+ $Y2=0
cc_900 N_A_955_21#_c_1096_n N_SCE_M1024_g 5.19778e-19 $X=7.12 $Y=1.92 $X2=0
+ $Y2=0
cc_901 N_A_955_21#_c_1092_n N_SCE_M1024_g 7.94182e-19 $X=7.235 $Y=1.52 $X2=0
+ $Y2=0
cc_902 N_A_955_21#_c_1085_n N_SCE_c_1251_n 0.0087278f $X=4.925 $Y=0.84 $X2=0
+ $Y2=0
cc_903 N_A_955_21#_c_1084_n SCE 0.0021051f $X=5.63 $Y=0.84 $X2=0 $Y2=0
cc_904 N_A_955_21#_c_1088_n SCE 0.00399999f $X=5.895 $Y=0.385 $X2=0 $Y2=0
cc_905 N_A_955_21#_c_1089_n SCE 6.16455e-19 $X=5.765 $Y=0.34 $X2=0 $Y2=0
cc_906 N_A_955_21#_c_1091_n SCE 0.0370038f $X=6.14 $Y=1.835 $X2=0 $Y2=0
cc_907 N_A_955_21#_c_1098_n SCE 0.00528494f $X=5.955 $Y=2 $X2=0 $Y2=0
cc_908 N_A_955_21#_c_1084_n N_SCE_c_1247_n 0.00692221f $X=5.63 $Y=0.84 $X2=0
+ $Y2=0
cc_909 N_A_955_21#_c_1091_n N_SCE_c_1247_n 0.0277865f $X=6.14 $Y=1.835 $X2=0
+ $Y2=0
cc_910 N_A_955_21#_c_1096_n N_SCE_c_1247_n 0.00152823f $X=7.12 $Y=1.92 $X2=0
+ $Y2=0
cc_911 N_A_955_21#_c_1098_n N_SCE_c_1247_n 0.00370055f $X=5.955 $Y=2 $X2=0 $Y2=0
cc_912 N_A_955_21#_c_1093_n N_SCE_c_1247_n 0.0057535f $X=6.06 $Y=0.935 $X2=0
+ $Y2=0
cc_913 N_A_955_21#_c_1087_n N_A_211_363#_c_1342_n 0.0122891f $X=7.32 $Y=1.77
+ $X2=0 $Y2=0
cc_914 N_A_955_21#_c_1087_n N_A_211_363#_c_1343_n 0.0121931f $X=7.32 $Y=1.77
+ $X2=0 $Y2=0
cc_915 N_A_955_21#_c_1085_n N_A_211_363#_c_1346_n 7.61895e-19 $X=4.925 $Y=0.84
+ $X2=0 $Y2=0
cc_916 N_A_955_21#_c_1087_n N_A_211_363#_c_1346_n 0.0029882f $X=7.32 $Y=1.77
+ $X2=0 $Y2=0
cc_917 N_A_955_21#_c_1091_n N_A_211_363#_c_1346_n 0.0129769f $X=6.14 $Y=1.835
+ $X2=0 $Y2=0
cc_918 N_A_955_21#_c_1096_n N_A_211_363#_c_1346_n 0.00367981f $X=7.12 $Y=1.92
+ $X2=0 $Y2=0
cc_919 N_A_955_21#_c_1092_n N_A_211_363#_c_1346_n 0.0148575f $X=7.235 $Y=1.52
+ $X2=0 $Y2=0
cc_920 N_A_955_21#_c_1098_n N_A_211_363#_c_1346_n 0.00120533f $X=5.955 $Y=2
+ $X2=0 $Y2=0
cc_921 N_A_955_21#_c_1093_n N_A_211_363#_c_1346_n 0.00398102f $X=6.06 $Y=0.935
+ $X2=0 $Y2=0
cc_922 N_A_955_21#_c_1087_n N_A_211_363#_c_1340_n 0.00361127f $X=7.32 $Y=1.77
+ $X2=0 $Y2=0
cc_923 N_A_955_21#_c_1096_n N_VPWR_M1022_d 0.00366079f $X=7.12 $Y=1.92 $X2=0
+ $Y2=0
cc_924 N_A_955_21#_c_1096_n N_VPWR_c_1921_n 0.0206935f $X=7.12 $Y=1.92 $X2=0
+ $Y2=0
cc_925 N_A_955_21#_c_1098_n N_VPWR_c_1921_n 0.0185696f $X=5.955 $Y=2 $X2=0 $Y2=0
cc_926 N_A_955_21#_c_1087_n N_VPWR_c_1922_n 0.00563362f $X=7.32 $Y=1.77 $X2=0
+ $Y2=0
cc_927 N_A_955_21#_c_1096_n N_VPWR_c_1922_n 0.00906057f $X=7.12 $Y=1.92 $X2=0
+ $Y2=0
cc_928 N_A_955_21#_c_1096_n N_VPWR_c_1938_n 0.00137879f $X=7.12 $Y=1.92 $X2=0
+ $Y2=0
cc_929 N_A_955_21#_c_1098_n N_VPWR_c_1938_n 0.0230749f $X=5.955 $Y=2 $X2=0 $Y2=0
cc_930 N_A_955_21#_M1022_s N_VPWR_c_1917_n 0.00182584f $X=5.83 $Y=1.845 $X2=0
+ $Y2=0
cc_931 N_A_955_21#_c_1087_n N_VPWR_c_1917_n 0.00739939f $X=7.32 $Y=1.77 $X2=0
+ $Y2=0
cc_932 N_A_955_21#_c_1096_n N_VPWR_c_1917_n 0.00947732f $X=7.12 $Y=1.92 $X2=0
+ $Y2=0
cc_933 N_A_955_21#_c_1098_n N_VPWR_c_1917_n 0.00711001f $X=5.955 $Y=2 $X2=0
+ $Y2=0
cc_934 N_A_955_21#_c_1085_n N_A_319_47#_c_2147_n 0.00354861f $X=4.925 $Y=0.84
+ $X2=0 $Y2=0
cc_935 N_A_955_21#_c_1083_n N_A_319_47#_c_2150_n 0.00294306f $X=4.85 $Y=0.765
+ $X2=0 $Y2=0
cc_936 N_A_955_21#_c_1098_n N_A_985_47#_c_2269_n 0.00597833f $X=5.955 $Y=2 $X2=0
+ $Y2=0
cc_937 N_A_955_21#_c_1098_n N_A_985_47#_c_2270_n 0.0202314f $X=5.955 $Y=2 $X2=0
+ $Y2=0
cc_938 N_A_955_21#_c_1084_n N_A_985_47#_c_2261_n 0.0099502f $X=5.63 $Y=0.84
+ $X2=0 $Y2=0
cc_939 N_A_955_21#_c_1086_n N_A_985_47#_c_2261_n 0.00123232f $X=5.705 $Y=0.765
+ $X2=0 $Y2=0
cc_940 N_A_955_21#_c_1090_n N_A_985_47#_c_2261_n 0.00324948f $X=6.06 $Y=0.75
+ $X2=0 $Y2=0
cc_941 N_A_955_21#_c_1084_n N_A_985_47#_c_2262_n 0.00718124f $X=5.63 $Y=0.84
+ $X2=0 $Y2=0
cc_942 N_A_955_21#_c_1093_n N_A_985_47#_c_2262_n 0.00324948f $X=6.06 $Y=0.935
+ $X2=0 $Y2=0
cc_943 N_A_955_21#_c_1087_n N_A_985_47#_c_2263_n 0.00292257f $X=7.32 $Y=1.77
+ $X2=0 $Y2=0
cc_944 N_A_955_21#_c_1092_n N_A_985_47#_c_2263_n 0.00529702f $X=7.235 $Y=1.52
+ $X2=0 $Y2=0
cc_945 N_A_955_21#_c_1087_n N_A_985_47#_c_2264_n 0.00866347f $X=7.32 $Y=1.77
+ $X2=0 $Y2=0
cc_946 N_A_955_21#_c_1096_n N_A_985_47#_c_2264_n 0.0123117f $X=7.12 $Y=1.92
+ $X2=0 $Y2=0
cc_947 N_A_955_21#_c_1092_n N_A_985_47#_c_2264_n 0.0339761f $X=7.235 $Y=1.52
+ $X2=0 $Y2=0
cc_948 N_A_955_21#_c_1083_n N_A_985_47#_c_2265_n 9.60356e-19 $X=4.85 $Y=0.765
+ $X2=0 $Y2=0
cc_949 N_A_955_21#_c_1086_n N_A_985_47#_c_2265_n 7.02746e-19 $X=5.705 $Y=0.765
+ $X2=0 $Y2=0
cc_950 N_A_955_21#_c_1084_n N_A_985_47#_c_2267_n 0.00350009f $X=5.63 $Y=0.84
+ $X2=0 $Y2=0
cc_951 N_A_955_21#_c_1086_n N_A_985_47#_c_2267_n 0.00252516f $X=5.705 $Y=0.765
+ $X2=0 $Y2=0
cc_952 N_A_955_21#_c_1088_n N_A_985_47#_c_2267_n 0.0306342f $X=5.895 $Y=0.385
+ $X2=0 $Y2=0
cc_953 N_A_955_21#_c_1090_n N_A_985_47#_c_2267_n 0.0105203f $X=6.06 $Y=0.75
+ $X2=0 $Y2=0
cc_954 N_A_955_21#_c_1083_n N_A_985_47#_c_2320_n 0.00282475f $X=4.85 $Y=0.765
+ $X2=0 $Y2=0
cc_955 N_A_955_21#_c_1086_n N_A_985_47#_c_2320_n 0.00172165f $X=5.705 $Y=0.765
+ $X2=0 $Y2=0
cc_956 N_A_955_21#_c_1088_n N_A_985_47#_c_2320_n 0.0202274f $X=5.895 $Y=0.385
+ $X2=0 $Y2=0
cc_957 N_A_955_21#_c_1089_n N_A_985_47#_c_2320_n 5.32913e-19 $X=5.765 $Y=0.34
+ $X2=0 $Y2=0
cc_958 N_A_955_21#_c_1096_n A_1376_369# 0.00449554f $X=7.12 $Y=1.92 $X2=-0.19
+ $Y2=-0.24
cc_959 N_A_955_21#_c_1088_n N_VGND_c_2449_n 0.0157484f $X=5.895 $Y=0.385 $X2=0
+ $Y2=0
cc_960 N_A_955_21#_c_1089_n N_VGND_c_2449_n 4.47621e-19 $X=5.765 $Y=0.34 $X2=0
+ $Y2=0
cc_961 N_A_955_21#_c_1090_n N_VGND_c_2449_n 0.0222116f $X=6.06 $Y=0.75 $X2=0
+ $Y2=0
cc_962 N_A_955_21#_c_1083_n N_VGND_c_2464_n 0.00585385f $X=4.85 $Y=0.765 $X2=0
+ $Y2=0
cc_963 N_A_955_21#_c_1084_n N_VGND_c_2464_n 0.00239942f $X=5.63 $Y=0.84 $X2=0
+ $Y2=0
cc_964 N_A_955_21#_c_1088_n N_VGND_c_2464_n 0.0578663f $X=5.895 $Y=0.385 $X2=0
+ $Y2=0
cc_965 N_A_955_21#_c_1089_n N_VGND_c_2464_n 0.00544529f $X=5.765 $Y=0.34 $X2=0
+ $Y2=0
cc_966 N_A_955_21#_c_1083_n N_VGND_c_2469_n 0.00741933f $X=4.85 $Y=0.765 $X2=0
+ $Y2=0
cc_967 N_A_955_21#_c_1088_n N_VGND_c_2469_n 0.00751944f $X=5.895 $Y=0.385 $X2=0
+ $Y2=0
cc_968 N_A_955_21#_c_1089_n N_VGND_c_2469_n 0.00692302f $X=5.765 $Y=0.34 $X2=0
+ $Y2=0
cc_969 N_SCD_c_1201_n N_SCE_c_1250_n 0.0222607f $X=6.79 $Y=1.77 $X2=0 $Y2=0
cc_970 N_SCD_M1038_g N_SCE_M1015_g 0.0140582f $X=6.79 $Y=0.805 $X2=0 $Y2=0
cc_971 N_SCD_M1038_g N_SCE_c_1243_n 0.0101836f $X=6.79 $Y=0.805 $X2=0 $Y2=0
cc_972 N_SCD_M1038_g N_SCE_M1024_g 0.0431259f $X=6.79 $Y=0.805 $X2=0 $Y2=0
cc_973 SCD N_SCE_M1024_g 3.47742e-19 $X=6.58 $Y=1.105 $X2=0 $Y2=0
cc_974 N_SCD_c_1201_n N_SCE_c_1247_n 0.0184356f $X=6.79 $Y=1.77 $X2=0 $Y2=0
cc_975 N_SCD_M1038_g N_SCE_c_1247_n 0.00286662f $X=6.79 $Y=0.805 $X2=0 $Y2=0
cc_976 SCD N_SCE_c_1247_n 0.00462329f $X=6.58 $Y=1.105 $X2=0 $Y2=0
cc_977 SCD N_A_211_363#_c_1346_n 0.0270775f $X=6.58 $Y=1.105 $X2=0 $Y2=0
cc_978 N_SCD_c_1201_n N_VPWR_c_1921_n 0.0055053f $X=6.79 $Y=1.77 $X2=0 $Y2=0
cc_979 N_SCD_c_1201_n N_VPWR_c_1922_n 0.00523784f $X=6.79 $Y=1.77 $X2=0 $Y2=0
cc_980 N_SCD_c_1201_n N_VPWR_c_1917_n 0.00687597f $X=6.79 $Y=1.77 $X2=0 $Y2=0
cc_981 N_SCD_M1038_g N_A_985_47#_c_2263_n 2.44187e-19 $X=6.79 $Y=0.805 $X2=0
+ $Y2=0
cc_982 SCD N_A_985_47#_c_2263_n 0.00423655f $X=6.58 $Y=1.105 $X2=0 $Y2=0
cc_983 N_SCD_M1038_g N_A_985_47#_c_2264_n 7.62122e-19 $X=6.79 $Y=0.805 $X2=0
+ $Y2=0
cc_984 SCD N_A_985_47#_c_2264_n 0.0058585f $X=6.58 $Y=1.105 $X2=0 $Y2=0
cc_985 N_SCD_M1038_g N_A_985_47#_c_2266_n 2.03985e-19 $X=6.79 $Y=0.805 $X2=0
+ $Y2=0
cc_986 N_SCD_M1038_g N_A_985_47#_c_2267_n 0.00301141f $X=6.79 $Y=0.805 $X2=0
+ $Y2=0
cc_987 N_SCD_c_1201_n N_VGND_c_2449_n 4.32649e-19 $X=6.79 $Y=1.77 $X2=0 $Y2=0
cc_988 N_SCD_M1038_g N_VGND_c_2449_n 0.00223007f $X=6.79 $Y=0.805 $X2=0 $Y2=0
cc_989 SCD N_VGND_c_2449_n 0.0146735f $X=6.58 $Y=1.105 $X2=0 $Y2=0
cc_990 N_SCE_c_1241_n N_A_211_363#_c_1346_n 0.00674772f $X=5.57 $Y=1.5 $X2=0
+ $Y2=0
cc_991 N_SCE_M1024_g N_A_211_363#_c_1346_n 5.39536e-19 $X=7.15 $Y=0.805 $X2=0
+ $Y2=0
cc_992 N_SCE_c_1251_n N_A_211_363#_c_1346_n 0.00334076f $X=4.915 $Y=1.5 $X2=0
+ $Y2=0
cc_993 SCE N_A_211_363#_c_1346_n 0.0167072f $X=5.67 $Y=1.43 $X2=0 $Y2=0
cc_994 N_SCE_c_1247_n N_A_211_363#_c_1346_n 0.00653411f $X=6.195 $Y=1.43 $X2=0
+ $Y2=0
cc_995 N_SCE_c_1250_n N_VPWR_c_1921_n 0.00645414f $X=6.195 $Y=1.77 $X2=0 $Y2=0
cc_996 N_SCE_c_1248_n N_VPWR_c_1938_n 0.00663173f $X=4.915 $Y=1.77 $X2=0 $Y2=0
cc_997 N_SCE_c_1250_n N_VPWR_c_1938_n 0.00512079f $X=6.195 $Y=1.77 $X2=0 $Y2=0
cc_998 N_SCE_c_1248_n N_VPWR_c_1917_n 0.00862708f $X=4.915 $Y=1.77 $X2=0 $Y2=0
cc_999 N_SCE_c_1250_n N_VPWR_c_1917_n 0.00800836f $X=6.195 $Y=1.77 $X2=0 $Y2=0
cc_1000 N_SCE_c_1248_n N_A_319_47#_c_2154_n 0.00350959f $X=4.915 $Y=1.77 $X2=0
+ $Y2=0
cc_1001 N_SCE_c_1248_n N_A_319_47#_c_2146_n 0.00122634f $X=4.915 $Y=1.77 $X2=0
+ $Y2=0
cc_1002 N_SCE_c_1251_n N_A_319_47#_c_2146_n 0.00833804f $X=4.915 $Y=1.5 $X2=0
+ $Y2=0
cc_1003 N_SCE_c_1241_n N_A_985_47#_c_2269_n 0.00386238f $X=5.57 $Y=1.5 $X2=0
+ $Y2=0
cc_1004 N_SCE_M1024_g N_A_985_47#_c_2260_n 0.0111092f $X=7.15 $Y=0.805 $X2=0
+ $Y2=0
cc_1005 N_SCE_c_1251_n N_A_985_47#_c_2261_n 7.45598e-19 $X=4.915 $Y=1.5 $X2=0
+ $Y2=0
cc_1006 N_SCE_c_1248_n N_A_985_47#_c_2262_n 0.00297796f $X=4.915 $Y=1.77 $X2=0
+ $Y2=0
cc_1007 N_SCE_c_1241_n N_A_985_47#_c_2262_n 0.0129434f $X=5.57 $Y=1.5 $X2=0
+ $Y2=0
cc_1008 N_SCE_c_1251_n N_A_985_47#_c_2262_n 0.00448589f $X=4.915 $Y=1.5 $X2=0
+ $Y2=0
cc_1009 SCE N_A_985_47#_c_2262_n 0.0208239f $X=5.67 $Y=1.43 $X2=0 $Y2=0
cc_1010 N_SCE_c_1247_n N_A_985_47#_c_2262_n 0.00286812f $X=6.195 $Y=1.43 $X2=0
+ $Y2=0
cc_1011 N_SCE_M1024_g N_A_985_47#_c_2266_n 0.00369264f $X=7.15 $Y=0.805 $X2=0
+ $Y2=0
cc_1012 N_SCE_M1015_g N_A_985_47#_c_2267_n 0.00415982f $X=6.27 $Y=0.805 $X2=0
+ $Y2=0
cc_1013 N_SCE_c_1243_n N_A_985_47#_c_2267_n 0.00232706f $X=7.075 $Y=0.18 $X2=0
+ $Y2=0
cc_1014 N_SCE_M1024_g N_A_985_47#_c_2267_n 0.00482768f $X=7.15 $Y=0.805 $X2=0
+ $Y2=0
cc_1015 N_SCE_M1024_g N_A_985_47#_c_2268_n 0.00808626f $X=7.15 $Y=0.805 $X2=0
+ $Y2=0
cc_1016 N_SCE_M1015_g N_VGND_c_2449_n 0.00618563f $X=6.27 $Y=0.805 $X2=0 $Y2=0
cc_1017 N_SCE_c_1243_n N_VGND_c_2449_n 0.0207417f $X=7.075 $Y=0.18 $X2=0 $Y2=0
cc_1018 N_SCE_M1024_g N_VGND_c_2449_n 0.00409214f $X=7.15 $Y=0.805 $X2=0 $Y2=0
cc_1019 N_SCE_c_1244_n N_VGND_c_2464_n 0.00922468f $X=6.345 $Y=0.18 $X2=0 $Y2=0
cc_1020 N_SCE_c_1243_n N_VGND_c_2465_n 0.0195638f $X=7.075 $Y=0.18 $X2=0 $Y2=0
cc_1021 N_SCE_c_1243_n N_VGND_c_2469_n 0.0155555f $X=7.075 $Y=0.18 $X2=0 $Y2=0
cc_1022 N_SCE_c_1244_n N_VGND_c_2469_n 0.00517505f $X=6.345 $Y=0.18 $X2=0 $Y2=0
cc_1023 N_A_211_363#_c_1333_n N_A_1787_159#_c_1547_n 0.0139941f $X=8.54 $Y=1.29
+ $X2=0 $Y2=0
cc_1024 N_A_211_363#_c_1348_n N_A_1787_159#_c_1547_n 0.00186506f $X=11.545
+ $Y=1.53 $X2=0 $Y2=0
cc_1025 N_A_211_363#_M1042_g N_A_1787_159#_M1040_g 0.0190058f $X=8.615 $Y=0.415
+ $X2=0 $Y2=0
cc_1026 N_A_211_363#_c_1348_n N_A_1787_159#_c_1560_n 0.00886951f $X=11.545
+ $Y=1.53 $X2=0 $Y2=0
cc_1027 N_A_211_363#_c_1335_n N_A_1787_159#_M1010_g 0.0184231f $X=11.315
+ $Y=0.705 $X2=0 $Y2=0
cc_1028 N_A_211_363#_c_1336_n N_A_1787_159#_M1010_g 0.00191476f $X=11.475
+ $Y=0.87 $X2=0 $Y2=0
cc_1029 N_A_211_363#_c_1337_n N_A_1787_159#_c_1550_n 0.0184231f $X=11.475
+ $Y=0.87 $X2=0 $Y2=0
cc_1030 N_A_211_363#_c_1348_n N_A_1787_159#_c_1550_n 0.00123775f $X=11.545
+ $Y=1.53 $X2=0 $Y2=0
cc_1031 N_A_211_363#_c_1338_n N_A_1787_159#_c_1550_n 2.46861e-19 $X=11.715
+ $Y=1.53 $X2=0 $Y2=0
cc_1032 N_A_211_363#_c_1348_n N_A_1787_159#_c_1551_n 0.00252648f $X=11.545
+ $Y=1.53 $X2=0 $Y2=0
cc_1033 N_A_211_363#_c_1348_n N_A_1787_159#_c_1552_n 0.00787458f $X=11.545
+ $Y=1.53 $X2=0 $Y2=0
cc_1034 N_A_211_363#_c_1348_n N_A_1787_159#_c_1564_n 0.0290415f $X=11.545
+ $Y=1.53 $X2=0 $Y2=0
cc_1035 N_A_211_363#_c_1348_n N_A_1787_159#_c_1554_n 0.0182403f $X=11.545
+ $Y=1.53 $X2=0 $Y2=0
cc_1036 N_A_211_363#_c_1348_n N_A_1787_159#_c_1556_n 9.1448e-19 $X=11.545
+ $Y=1.53 $X2=0 $Y2=0
cc_1037 N_A_211_363#_M1042_g N_A_1787_159#_c_1557_n 0.0139941f $X=8.615 $Y=0.415
+ $X2=0 $Y2=0
cc_1038 N_A_211_363#_c_1348_n N_A_1611_413#_c_1675_n 8.02119e-19 $X=11.545
+ $Y=1.53 $X2=0 $Y2=0
cc_1039 N_A_211_363#_c_1348_n N_A_1611_413#_c_1676_n 0.00281761f $X=11.545
+ $Y=1.53 $X2=0 $Y2=0
cc_1040 N_A_211_363#_c_1343_n N_A_1611_413#_c_1686_n 0.0046816f $X=7.965 $Y=1.99
+ $X2=0 $Y2=0
cc_1041 N_A_211_363#_c_1339_n N_A_1611_413#_c_1686_n 0.00145976f $X=7.965
+ $Y=1.35 $X2=0 $Y2=0
cc_1042 N_A_211_363#_c_1340_n N_A_1611_413#_c_1686_n 0.00117048f $X=8.18 $Y=1.35
+ $X2=0 $Y2=0
cc_1043 N_A_211_363#_c_1333_n N_A_1611_413#_c_1691_n 0.00171584f $X=8.54 $Y=1.29
+ $X2=0 $Y2=0
cc_1044 N_A_211_363#_M1042_g N_A_1611_413#_c_1691_n 0.0159788f $X=8.615 $Y=0.415
+ $X2=0 $Y2=0
cc_1045 N_A_211_363#_M1042_g N_A_1611_413#_c_1677_n 0.00891723f $X=8.615
+ $Y=0.415 $X2=0 $Y2=0
cc_1046 N_A_211_363#_c_1348_n N_A_1611_413#_c_1682_n 0.00508278f $X=11.545
+ $Y=1.53 $X2=0 $Y2=0
cc_1047 N_A_211_363#_c_1333_n N_A_1611_413#_c_1678_n 5.91184e-19 $X=8.54 $Y=1.29
+ $X2=0 $Y2=0
cc_1048 N_A_211_363#_c_1348_n N_A_1611_413#_c_1678_n 0.0393222f $X=11.545
+ $Y=1.53 $X2=0 $Y2=0
cc_1049 N_A_211_363#_c_1345_n N_A_2266_413#_c_1801_n 0.0143369f $X=11.71 $Y=1.99
+ $X2=0 $Y2=0
cc_1050 N_A_211_363#_c_1348_n N_A_2266_413#_c_1801_n 0.00391921f $X=11.545
+ $Y=1.53 $X2=0 $Y2=0
cc_1051 N_A_211_363#_c_1397_n N_A_2266_413#_c_1801_n 0.00120832f $X=11.715
+ $Y=1.53 $X2=0 $Y2=0
cc_1052 N_A_211_363#_c_1338_n N_A_2266_413#_c_1801_n 0.02356f $X=11.715 $Y=1.53
+ $X2=0 $Y2=0
cc_1053 N_A_211_363#_c_1336_n N_A_2266_413#_c_1805_n 0.0330221f $X=11.475
+ $Y=0.87 $X2=0 $Y2=0
cc_1054 N_A_211_363#_c_1337_n N_A_2266_413#_c_1805_n 0.00134485f $X=11.475
+ $Y=0.87 $X2=0 $Y2=0
cc_1055 N_A_211_363#_c_1345_n N_A_2266_413#_c_1796_n 0.00233263f $X=11.71
+ $Y=1.99 $X2=0 $Y2=0
cc_1056 N_A_211_363#_c_1338_n N_A_2266_413#_c_1796_n 0.00722817f $X=11.715
+ $Y=1.53 $X2=0 $Y2=0
cc_1057 N_A_211_363#_c_1345_n N_A_2266_413#_c_1787_n 0.00576207f $X=11.71
+ $Y=1.99 $X2=0 $Y2=0
cc_1058 N_A_211_363#_c_1336_n N_A_2266_413#_c_1787_n 0.0801552f $X=11.475
+ $Y=0.87 $X2=0 $Y2=0
cc_1059 N_A_211_363#_c_1397_n N_A_2266_413#_c_1787_n 0.00162538f $X=11.715
+ $Y=1.53 $X2=0 $Y2=0
cc_1060 N_A_211_363#_c_1341_n N_VPWR_c_1918_n 0.0202126f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_1061 N_A_211_363#_c_1346_n N_VPWR_c_1919_n 0.00168188f $X=7.825 $Y=1.53 $X2=0
+ $Y2=0
cc_1062 N_A_211_363#_c_1346_n N_VPWR_c_1920_n 7.40558e-19 $X=7.825 $Y=1.53 $X2=0
+ $Y2=0
cc_1063 N_A_211_363#_c_1343_n N_VPWR_c_1922_n 0.00646384f $X=7.965 $Y=1.99 $X2=0
+ $Y2=0
cc_1064 N_A_211_363#_c_1348_n N_VPWR_c_1923_n 8.15834e-19 $X=11.545 $Y=1.53
+ $X2=0 $Y2=0
cc_1065 N_A_211_363#_c_1341_n N_VPWR_c_1937_n 0.0120448f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_1066 N_A_211_363#_c_1345_n N_VPWR_c_1939_n 0.00455772f $X=11.71 $Y=1.99 $X2=0
+ $Y2=0
cc_1067 N_A_211_363#_c_1343_n N_VPWR_c_1917_n 0.00776738f $X=7.965 $Y=1.99 $X2=0
+ $Y2=0
cc_1068 N_A_211_363#_c_1345_n N_VPWR_c_1917_n 0.00666932f $X=11.71 $Y=1.99 $X2=0
+ $Y2=0
cc_1069 N_A_211_363#_c_1341_n N_VPWR_c_1917_n 0.00308197f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_1070 N_A_211_363#_c_1346_n N_A_319_47#_c_2152_n 0.00102404f $X=7.825 $Y=1.53
+ $X2=0 $Y2=0
cc_1071 N_A_211_363#_c_1346_n N_A_319_47#_c_2145_n 0.0170715f $X=7.825 $Y=1.53
+ $X2=0 $Y2=0
cc_1072 N_A_211_363#_c_1347_n N_A_319_47#_c_2145_n 0.00283132f $X=1.345 $Y=1.53
+ $X2=0 $Y2=0
cc_1073 N_A_211_363#_c_1341_n N_A_319_47#_c_2145_n 0.145282f $X=1.2 $Y=0.51
+ $X2=0 $Y2=0
cc_1074 N_A_211_363#_c_1346_n N_A_319_47#_c_2154_n 9.16782e-19 $X=7.825 $Y=1.53
+ $X2=0 $Y2=0
cc_1075 N_A_211_363#_c_1346_n N_A_319_47#_c_2146_n 0.0129523f $X=7.825 $Y=1.53
+ $X2=0 $Y2=0
cc_1076 N_A_211_363#_c_1346_n N_A_319_47#_c_2147_n 0.00293129f $X=7.825 $Y=1.53
+ $X2=0 $Y2=0
cc_1077 N_A_211_363#_c_1341_n N_A_319_47#_c_2148_n 0.00796831f $X=1.2 $Y=0.51
+ $X2=0 $Y2=0
cc_1078 N_A_211_363#_c_1341_n N_A_319_47#_c_2151_n 0.0117897f $X=1.2 $Y=0.51
+ $X2=0 $Y2=0
cc_1079 N_A_211_363#_c_1346_n N_A_985_47#_c_2269_n 0.00360434f $X=7.825 $Y=1.53
+ $X2=0 $Y2=0
cc_1080 N_A_211_363#_c_1342_n N_A_985_47#_c_2282_n 0.00153446f $X=7.965 $Y=1.89
+ $X2=0 $Y2=0
cc_1081 N_A_211_363#_c_1346_n N_A_985_47#_c_2282_n 4.75993e-19 $X=7.825 $Y=1.53
+ $X2=0 $Y2=0
cc_1082 N_A_211_363#_c_1343_n N_A_985_47#_c_2346_n 0.00943842f $X=7.965 $Y=1.99
+ $X2=0 $Y2=0
cc_1083 N_A_211_363#_c_1346_n N_A_985_47#_c_2262_n 0.0139678f $X=7.825 $Y=1.53
+ $X2=0 $Y2=0
cc_1084 N_A_211_363#_c_1346_n N_A_985_47#_c_2263_n 0.00592292f $X=7.825 $Y=1.53
+ $X2=0 $Y2=0
cc_1085 N_A_211_363#_c_1339_n N_A_985_47#_c_2263_n 0.0424828f $X=7.965 $Y=1.35
+ $X2=0 $Y2=0
cc_1086 N_A_211_363#_c_1342_n N_A_985_47#_c_2264_n 0.00314461f $X=7.965 $Y=1.89
+ $X2=0 $Y2=0
cc_1087 N_A_211_363#_c_1346_n N_A_985_47#_c_2264_n 0.0128597f $X=7.825 $Y=1.53
+ $X2=0 $Y2=0
cc_1088 N_A_211_363#_c_1349_n N_A_985_47#_c_2264_n 0.00263822f $X=8.165 $Y=1.53
+ $X2=0 $Y2=0
cc_1089 N_A_211_363#_c_1340_n N_A_985_47#_c_2264_n 0.00516969f $X=8.18 $Y=1.35
+ $X2=0 $Y2=0
cc_1090 N_A_211_363#_c_1339_n N_A_985_47#_c_2268_n 2.86271e-19 $X=7.965 $Y=1.35
+ $X2=0 $Y2=0
cc_1091 N_A_211_363#_c_1340_n N_A_985_47#_c_2268_n 0.00207603f $X=8.18 $Y=1.35
+ $X2=0 $Y2=0
cc_1092 N_A_211_363#_M1042_g N_VGND_c_2450_n 0.00129001f $X=8.615 $Y=0.415 $X2=0
+ $Y2=0
cc_1093 N_A_211_363#_c_1341_n N_VGND_c_2463_n 0.00732874f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_1094 N_A_211_363#_M1042_g N_VGND_c_2465_n 0.00357877f $X=8.615 $Y=0.415 $X2=0
+ $Y2=0
cc_1095 N_A_211_363#_c_1335_n N_VGND_c_2466_n 0.00585385f $X=11.315 $Y=0.705
+ $X2=0 $Y2=0
cc_1096 N_A_211_363#_c_1336_n N_VGND_c_2466_n 2.78187e-19 $X=11.475 $Y=0.87
+ $X2=0 $Y2=0
cc_1097 N_A_211_363#_c_1337_n N_VGND_c_2466_n 2.25106e-19 $X=11.475 $Y=0.87
+ $X2=0 $Y2=0
cc_1098 N_A_211_363#_M1001_d N_VGND_c_2469_n 0.00535012f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_1099 N_A_211_363#_M1042_g N_VGND_c_2469_n 0.00580066f $X=8.615 $Y=0.415 $X2=0
+ $Y2=0
cc_1100 N_A_211_363#_c_1335_n N_VGND_c_2469_n 0.00718386f $X=11.315 $Y=0.705
+ $X2=0 $Y2=0
cc_1101 N_A_211_363#_c_1336_n N_VGND_c_2469_n 0.00121732f $X=11.475 $Y=0.87
+ $X2=0 $Y2=0
cc_1102 N_A_211_363#_c_1341_n N_VGND_c_2469_n 0.00616598f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_1103 N_A_1787_159#_c_1552_n N_A_1611_413#_c_1672_n 0.00747237f $X=9.765
+ $Y=0.915 $X2=0 $Y2=0
cc_1104 N_A_1787_159#_c_1554_n N_A_1611_413#_c_1672_n 2.82106e-19 $X=10.645
+ $Y=1.21 $X2=0 $Y2=0
cc_1105 N_A_1787_159#_c_1555_n N_A_1611_413#_c_1672_n 0.00149808f $X=10.645
+ $Y=1.21 $X2=0 $Y2=0
cc_1106 N_A_1787_159#_c_1547_n N_A_1611_413#_c_1679_n 0.00425243f $X=9.035
+ $Y=1.89 $X2=0 $Y2=0
cc_1107 N_A_1787_159#_c_1559_n N_A_1611_413#_c_1679_n 0.00717803f $X=9.035
+ $Y=1.99 $X2=0 $Y2=0
cc_1108 N_A_1787_159#_c_1564_n N_A_1611_413#_c_1679_n 0.0159286f $X=9.98 $Y=1.88
+ $X2=0 $Y2=0
cc_1109 N_A_1787_159#_M1040_g N_A_1611_413#_c_1673_n 0.00927877f $X=9.145
+ $Y=0.445 $X2=0 $Y2=0
cc_1110 N_A_1787_159#_c_1550_n N_A_1611_413#_c_1673_n 0.00146207f $X=10.707
+ $Y=1.045 $X2=0 $Y2=0
cc_1111 N_A_1787_159#_c_1552_n N_A_1611_413#_c_1673_n 0.00531123f $X=9.765
+ $Y=0.915 $X2=0 $Y2=0
cc_1112 N_A_1787_159#_c_1553_n N_A_1611_413#_c_1673_n 0.0135961f $X=10.05
+ $Y=0.39 $X2=0 $Y2=0
cc_1113 N_A_1787_159#_c_1557_n N_A_1611_413#_c_1673_n 0.00413802f $X=9.145
+ $Y=0.93 $X2=0 $Y2=0
cc_1114 N_A_1787_159#_c_1547_n N_A_1611_413#_c_1674_n 0.00484954f $X=9.035
+ $Y=1.89 $X2=0 $Y2=0
cc_1115 N_A_1787_159#_c_1552_n N_A_1611_413#_c_1674_n 0.0148713f $X=9.765
+ $Y=0.915 $X2=0 $Y2=0
cc_1116 N_A_1787_159#_c_1555_n N_A_1611_413#_c_1674_n 0.00146207f $X=10.645
+ $Y=1.21 $X2=0 $Y2=0
cc_1117 N_A_1787_159#_c_1556_n N_A_1611_413#_c_1674_n 2.59308e-19 $X=9.305
+ $Y=0.93 $X2=0 $Y2=0
cc_1118 N_A_1787_159#_c_1557_n N_A_1611_413#_c_1674_n 0.0050046f $X=9.145
+ $Y=0.93 $X2=0 $Y2=0
cc_1119 N_A_1787_159#_c_1547_n N_A_1611_413#_c_1675_n 0.0175058f $X=9.035
+ $Y=1.89 $X2=0 $Y2=0
cc_1120 N_A_1787_159#_c_1552_n N_A_1611_413#_c_1675_n 0.00455719f $X=9.765
+ $Y=0.915 $X2=0 $Y2=0
cc_1121 N_A_1787_159#_c_1557_n N_A_1611_413#_c_1675_n 5.95332e-19 $X=9.145
+ $Y=0.93 $X2=0 $Y2=0
cc_1122 N_A_1787_159#_c_1547_n N_A_1611_413#_c_1676_n 0.002305f $X=9.035 $Y=1.89
+ $X2=0 $Y2=0
cc_1123 N_A_1787_159#_c_1551_n N_A_1611_413#_c_1676_n 0.00149808f $X=10.672
+ $Y=1.375 $X2=0 $Y2=0
cc_1124 N_A_1787_159#_c_1552_n N_A_1611_413#_c_1676_n 0.00386856f $X=9.765
+ $Y=0.915 $X2=0 $Y2=0
cc_1125 N_A_1787_159#_c_1564_n N_A_1611_413#_c_1676_n 0.011301f $X=9.98 $Y=1.88
+ $X2=0 $Y2=0
cc_1126 N_A_1787_159#_c_1559_n N_A_1611_413#_c_1686_n 0.0108944f $X=9.035
+ $Y=1.99 $X2=0 $Y2=0
cc_1127 N_A_1787_159#_M1040_g N_A_1611_413#_c_1691_n 0.00290399f $X=9.145
+ $Y=0.445 $X2=0 $Y2=0
cc_1128 N_A_1787_159#_M1040_g N_A_1611_413#_c_1677_n 0.00424924f $X=9.145
+ $Y=0.445 $X2=0 $Y2=0
cc_1129 N_A_1787_159#_c_1556_n N_A_1611_413#_c_1677_n 0.0223112f $X=9.305
+ $Y=0.93 $X2=0 $Y2=0
cc_1130 N_A_1787_159#_c_1557_n N_A_1611_413#_c_1677_n 0.00632916f $X=9.145
+ $Y=0.93 $X2=0 $Y2=0
cc_1131 N_A_1787_159#_c_1547_n N_A_1611_413#_c_1682_n 0.00946574f $X=9.035
+ $Y=1.89 $X2=0 $Y2=0
cc_1132 N_A_1787_159#_c_1559_n N_A_1611_413#_c_1682_n 0.0100449f $X=9.035
+ $Y=1.99 $X2=0 $Y2=0
cc_1133 N_A_1787_159#_c_1564_n N_A_1611_413#_c_1682_n 0.00704799f $X=9.98
+ $Y=1.88 $X2=0 $Y2=0
cc_1134 N_A_1787_159#_c_1547_n N_A_1611_413#_c_1678_n 0.0157314f $X=9.035
+ $Y=1.89 $X2=0 $Y2=0
cc_1135 N_A_1787_159#_c_1552_n N_A_1611_413#_c_1678_n 0.0419277f $X=9.765
+ $Y=0.915 $X2=0 $Y2=0
cc_1136 N_A_1787_159#_c_1556_n N_A_1611_413#_c_1678_n 0.0141151f $X=9.305
+ $Y=0.93 $X2=0 $Y2=0
cc_1137 N_A_1787_159#_c_1557_n N_A_1611_413#_c_1678_n 0.0019926f $X=9.145
+ $Y=0.93 $X2=0 $Y2=0
cc_1138 N_A_1787_159#_c_1561_n N_A_2266_413#_c_1801_n 6.12204e-19 $X=10.735
+ $Y=1.99 $X2=0 $Y2=0
cc_1139 N_A_1787_159#_c_1559_n N_VPWR_c_1922_n 0.00453517f $X=9.035 $Y=1.99
+ $X2=0 $Y2=0
cc_1140 N_A_1787_159#_c_1547_n N_VPWR_c_1923_n 4.7516e-19 $X=9.035 $Y=1.89 $X2=0
+ $Y2=0
cc_1141 N_A_1787_159#_c_1559_n N_VPWR_c_1923_n 0.00594375f $X=9.035 $Y=1.99
+ $X2=0 $Y2=0
cc_1142 N_A_1787_159#_c_1564_n N_VPWR_c_1923_n 0.0472096f $X=9.98 $Y=1.88 $X2=0
+ $Y2=0
cc_1143 N_A_1787_159#_c_1561_n N_VPWR_c_1924_n 0.00531521f $X=10.735 $Y=1.99
+ $X2=0 $Y2=0
cc_1144 N_A_1787_159#_c_1564_n N_VPWR_c_1924_n 0.0258793f $X=9.98 $Y=1.88 $X2=0
+ $Y2=0
cc_1145 N_A_1787_159#_c_1564_n N_VPWR_c_1932_n 0.0244686f $X=9.98 $Y=1.88 $X2=0
+ $Y2=0
cc_1146 N_A_1787_159#_c_1561_n N_VPWR_c_1939_n 0.00721387f $X=10.735 $Y=1.99
+ $X2=0 $Y2=0
cc_1147 N_A_1787_159#_M1000_d N_VPWR_c_1917_n 0.00179197f $X=9.835 $Y=1.735
+ $X2=0 $Y2=0
cc_1148 N_A_1787_159#_c_1559_n N_VPWR_c_1917_n 0.00684226f $X=9.035 $Y=1.99
+ $X2=0 $Y2=0
cc_1149 N_A_1787_159#_c_1561_n N_VPWR_c_1917_n 0.00888708f $X=10.735 $Y=1.99
+ $X2=0 $Y2=0
cc_1150 N_A_1787_159#_c_1564_n N_VPWR_c_1917_n 0.00675092f $X=9.98 $Y=1.88 $X2=0
+ $Y2=0
cc_1151 N_A_1787_159#_c_1552_n N_VGND_M1040_d 0.00396111f $X=9.765 $Y=0.915
+ $X2=0 $Y2=0
cc_1152 N_A_1787_159#_M1040_g N_VGND_c_2450_n 0.0111851f $X=9.145 $Y=0.445 $X2=0
+ $Y2=0
cc_1153 N_A_1787_159#_c_1553_n N_VGND_c_2450_n 0.0225643f $X=10.05 $Y=0.39 $X2=0
+ $Y2=0
cc_1154 N_A_1787_159#_c_1556_n N_VGND_c_2450_n 0.0224132f $X=9.305 $Y=0.93 $X2=0
+ $Y2=0
cc_1155 N_A_1787_159#_c_1557_n N_VGND_c_2450_n 8.00172e-19 $X=9.145 $Y=0.93
+ $X2=0 $Y2=0
cc_1156 N_A_1787_159#_M1010_g N_VGND_c_2451_n 0.00506681f $X=10.83 $Y=0.445
+ $X2=0 $Y2=0
cc_1157 N_A_1787_159#_c_1550_n N_VGND_c_2451_n 0.00385985f $X=10.707 $Y=1.045
+ $X2=0 $Y2=0
cc_1158 N_A_1787_159#_c_1553_n N_VGND_c_2451_n 0.0239787f $X=10.05 $Y=0.39 $X2=0
+ $Y2=0
cc_1159 N_A_1787_159#_c_1554_n N_VGND_c_2451_n 0.00509394f $X=10.645 $Y=1.21
+ $X2=0 $Y2=0
cc_1160 N_A_1787_159#_c_1553_n N_VGND_c_2456_n 0.0295782f $X=10.05 $Y=0.39 $X2=0
+ $Y2=0
cc_1161 N_A_1787_159#_M1040_g N_VGND_c_2465_n 0.00427505f $X=9.145 $Y=0.445
+ $X2=0 $Y2=0
cc_1162 N_A_1787_159#_M1010_g N_VGND_c_2466_n 0.00585385f $X=10.83 $Y=0.445
+ $X2=0 $Y2=0
cc_1163 N_A_1787_159#_M1047_d N_VGND_c_2469_n 0.00172424f $X=9.915 $Y=0.235
+ $X2=0 $Y2=0
cc_1164 N_A_1787_159#_M1040_g N_VGND_c_2469_n 0.00390784f $X=9.145 $Y=0.445
+ $X2=0 $Y2=0
cc_1165 N_A_1787_159#_M1010_g N_VGND_c_2469_n 0.00782735f $X=10.83 $Y=0.445
+ $X2=0 $Y2=0
cc_1166 N_A_1787_159#_c_1552_n N_VGND_c_2469_n 0.00454361f $X=9.765 $Y=0.915
+ $X2=0 $Y2=0
cc_1167 N_A_1787_159#_c_1553_n N_VGND_c_2469_n 0.00795407f $X=10.05 $Y=0.39
+ $X2=0 $Y2=0
cc_1168 N_A_1787_159#_c_1556_n N_VGND_c_2469_n 0.00354771f $X=9.305 $Y=0.93
+ $X2=0 $Y2=0
cc_1169 N_A_1787_159#_c_1557_n N_VGND_c_2469_n 7.19298e-19 $X=9.145 $Y=0.93
+ $X2=0 $Y2=0
cc_1170 N_A_1611_413#_c_1686_n N_VPWR_M1028_d 0.00203143f $X=8.97 $Y=2.275 $X2=0
+ $Y2=0
cc_1171 N_A_1611_413#_c_1682_n N_VPWR_M1028_d 0.00102868f $X=9.08 $Y=2.175 $X2=0
+ $Y2=0
cc_1172 N_A_1611_413#_c_1686_n N_VPWR_c_1922_n 0.0432828f $X=8.97 $Y=2.275 $X2=0
+ $Y2=0
cc_1173 N_A_1611_413#_c_1679_n N_VPWR_c_1923_n 0.00526378f $X=9.745 $Y=1.66
+ $X2=0 $Y2=0
cc_1174 N_A_1611_413#_c_1675_n N_VPWR_c_1923_n 0.00133139f $X=9.645 $Y=1.41
+ $X2=0 $Y2=0
cc_1175 N_A_1611_413#_c_1686_n N_VPWR_c_1923_n 0.0166341f $X=8.97 $Y=2.275 $X2=0
+ $Y2=0
cc_1176 N_A_1611_413#_c_1682_n N_VPWR_c_1923_n 0.0253391f $X=9.08 $Y=2.175 $X2=0
+ $Y2=0
cc_1177 N_A_1611_413#_c_1678_n N_VPWR_c_1923_n 0.0109124f $X=9.08 $Y=1.41 $X2=0
+ $Y2=0
cc_1178 N_A_1611_413#_c_1679_n N_VPWR_c_1924_n 0.00289293f $X=9.745 $Y=1.66
+ $X2=0 $Y2=0
cc_1179 N_A_1611_413#_c_1679_n N_VPWR_c_1932_n 0.00597712f $X=9.745 $Y=1.66
+ $X2=0 $Y2=0
cc_1180 N_A_1611_413#_M1027_d N_VPWR_c_1917_n 0.00219504f $X=8.055 $Y=2.065
+ $X2=0 $Y2=0
cc_1181 N_A_1611_413#_c_1679_n N_VPWR_c_1917_n 0.00853572f $X=9.745 $Y=1.66
+ $X2=0 $Y2=0
cc_1182 N_A_1611_413#_c_1686_n N_VPWR_c_1917_n 0.0182363f $X=8.97 $Y=2.275 $X2=0
+ $Y2=0
cc_1183 N_A_1611_413#_c_1686_n N_A_985_47#_c_2286_n 0.0138511f $X=8.97 $Y=2.275
+ $X2=0 $Y2=0
cc_1184 N_A_1611_413#_c_1691_n N_A_985_47#_c_2266_n 6.17684e-19 $X=8.695 $Y=0.41
+ $X2=0 $Y2=0
cc_1185 N_A_1611_413#_c_1691_n N_A_985_47#_c_2268_n 0.0213204f $X=8.695 $Y=0.41
+ $X2=0 $Y2=0
cc_1186 N_A_1611_413#_c_1686_n A_1712_413# 0.00620654f $X=8.97 $Y=2.275
+ $X2=-0.19 $Y2=-0.24
cc_1187 N_A_1611_413#_c_1673_n N_VGND_c_2450_n 0.0055661f $X=9.78 $Y=0.95 $X2=0
+ $Y2=0
cc_1188 N_A_1611_413#_c_1691_n N_VGND_c_2450_n 0.0158772f $X=8.695 $Y=0.41 $X2=0
+ $Y2=0
cc_1189 N_A_1611_413#_c_1673_n N_VGND_c_2451_n 0.00214573f $X=9.78 $Y=0.95 $X2=0
+ $Y2=0
cc_1190 N_A_1611_413#_c_1673_n N_VGND_c_2456_n 0.00359186f $X=9.78 $Y=0.95 $X2=0
+ $Y2=0
cc_1191 N_A_1611_413#_c_1691_n N_VGND_c_2465_n 0.0427858f $X=8.695 $Y=0.41 $X2=0
+ $Y2=0
cc_1192 N_A_1611_413#_M1013_d N_VGND_c_2469_n 0.00256974f $X=8.15 $Y=0.235 $X2=0
+ $Y2=0
cc_1193 N_A_1611_413#_c_1673_n N_VGND_c_2469_n 0.00707393f $X=9.78 $Y=0.95 $X2=0
+ $Y2=0
cc_1194 N_A_1611_413#_c_1691_n N_VGND_c_2469_n 0.0124989f $X=8.695 $Y=0.41 $X2=0
+ $Y2=0
cc_1195 N_A_1611_413#_c_1691_n A_1738_47# 0.00469801f $X=8.695 $Y=0.41 $X2=-0.19
+ $Y2=-0.24
cc_1196 N_A_1611_413#_c_1677_n A_1738_47# 0.00105811f $X=8.78 $Y=1.315 $X2=-0.19
+ $Y2=-0.24
cc_1197 N_A_2266_413#_c_1795_n N_VPWR_M1039_d 0.00456215f $X=13.925 $Y=1.87
+ $X2=0 $Y2=0
cc_1198 N_A_2266_413#_c_1795_n N_VPWR_M1020_d 0.00191899f $X=13.925 $Y=1.87
+ $X2=0 $Y2=0
cc_1199 N_A_2266_413#_c_1801_n N_VPWR_c_1924_n 0.00580135f $X=12.125 $Y=2.26
+ $X2=0 $Y2=0
cc_1200 N_A_2266_413#_c_1801_n N_VPWR_c_1925_n 0.0122267f $X=12.125 $Y=2.26
+ $X2=0 $Y2=0
cc_1201 N_A_2266_413#_c_1795_n N_VPWR_c_1925_n 0.0155412f $X=13.925 $Y=1.87
+ $X2=0 $Y2=0
cc_1202 N_A_2266_413#_c_1796_n N_VPWR_c_1925_n 0.00221058f $X=12.395 $Y=1.87
+ $X2=0 $Y2=0
cc_1203 N_A_2266_413#_c_1787_n N_VPWR_c_1925_n 0.0373338f $X=12.25 $Y=1.87 $X2=0
+ $Y2=0
cc_1204 N_A_2266_413#_c_1795_n N_VPWR_c_1927_n 0.0204489f $X=13.925 $Y=1.87
+ $X2=0 $Y2=0
cc_1205 N_A_2266_413#_c_1798_n N_VPWR_c_1927_n 0.0026849f $X=14.07 $Y=1.87 $X2=0
+ $Y2=0
cc_1206 N_A_2266_413#_c_1799_n N_VPWR_c_1927_n 0.00429662f $X=14.07 $Y=1.542
+ $X2=0 $Y2=0
cc_1207 N_A_2266_413#_c_1800_n N_VPWR_c_1927_n 0.0311566f $X=14.07 $Y=1.74 $X2=0
+ $Y2=0
cc_1208 N_A_2266_413#_c_1789_n N_VPWR_c_1928_n 0.0096327f $X=14.765 $Y=1.77
+ $X2=0 $Y2=0
cc_1209 N_A_2266_413#_c_1782_n N_VPWR_c_1928_n 0.00717329f $X=15.2 $Y=1.16 $X2=0
+ $Y2=0
cc_1210 N_A_2266_413#_c_1783_n N_VPWR_c_1928_n 0.00317663f $X=14.865 $Y=1.16
+ $X2=0 $Y2=0
cc_1211 N_A_2266_413#_c_1792_n N_VPWR_c_1928_n 0.00710796f $X=15.3 $Y=1.41 $X2=0
+ $Y2=0
cc_1212 N_A_2266_413#_c_1793_n N_VPWR_c_1929_n 0.00987746f $X=15.77 $Y=1.41
+ $X2=0 $Y2=0
cc_1213 N_A_2266_413#_c_1792_n N_VPWR_c_1934_n 0.00601967f $X=15.3 $Y=1.41 $X2=0
+ $Y2=0
cc_1214 N_A_2266_413#_c_1793_n N_VPWR_c_1934_n 0.00674789f $X=15.77 $Y=1.41
+ $X2=0 $Y2=0
cc_1215 N_A_2266_413#_c_1801_n N_VPWR_c_1939_n 0.0382384f $X=12.125 $Y=2.26
+ $X2=0 $Y2=0
cc_1216 N_A_2266_413#_c_1789_n N_VPWR_c_1940_n 0.00673617f $X=14.765 $Y=1.77
+ $X2=0 $Y2=0
cc_1217 N_A_2266_413#_c_1800_n N_VPWR_c_1940_n 0.00385228f $X=14.07 $Y=1.74
+ $X2=0 $Y2=0
cc_1218 N_A_2266_413#_M1003_d N_VPWR_c_1917_n 0.0023091f $X=11.33 $Y=2.065 $X2=0
+ $Y2=0
cc_1219 N_A_2266_413#_c_1789_n N_VPWR_c_1917_n 0.0133664f $X=14.765 $Y=1.77
+ $X2=0 $Y2=0
cc_1220 N_A_2266_413#_c_1792_n N_VPWR_c_1917_n 0.0101591f $X=15.3 $Y=1.41 $X2=0
+ $Y2=0
cc_1221 N_A_2266_413#_c_1793_n N_VPWR_c_1917_n 0.0129392f $X=15.77 $Y=1.41 $X2=0
+ $Y2=0
cc_1222 N_A_2266_413#_c_1801_n N_VPWR_c_1917_n 0.029528f $X=12.125 $Y=2.26 $X2=0
+ $Y2=0
cc_1223 N_A_2266_413#_c_1795_n N_VPWR_c_1917_n 0.0714889f $X=13.925 $Y=1.87
+ $X2=0 $Y2=0
cc_1224 N_A_2266_413#_c_1796_n N_VPWR_c_1917_n 0.0147314f $X=12.395 $Y=1.87
+ $X2=0 $Y2=0
cc_1225 N_A_2266_413#_c_1798_n N_VPWR_c_1917_n 0.0154783f $X=14.07 $Y=1.87 $X2=0
+ $Y2=0
cc_1226 N_A_2266_413#_c_1799_n N_VPWR_c_1917_n 2.34088e-19 $X=14.07 $Y=1.542
+ $X2=0 $Y2=0
cc_1227 N_A_2266_413#_c_1800_n N_VPWR_c_1917_n 0.00276764f $X=14.07 $Y=1.74
+ $X2=0 $Y2=0
cc_1228 N_A_2266_413#_c_1801_n A_2360_413# 0.0121391f $X=12.125 $Y=2.26
+ $X2=-0.19 $Y2=-0.24
cc_1229 N_A_2266_413#_c_1787_n A_2360_413# 0.00136401f $X=12.25 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_1230 N_A_2266_413#_c_1795_n N_Q_N_c_2398_n 0.0371266f $X=13.925 $Y=1.87 $X2=0
+ $Y2=0
cc_1231 N_A_2266_413#_c_1799_n N_Q_N_c_2398_n 3.06319e-19 $X=14.07 $Y=1.542
+ $X2=0 $Y2=0
cc_1232 N_A_2266_413#_c_1795_n Q_N 0.00353799f $X=13.925 $Y=1.87 $X2=0 $Y2=0
cc_1233 N_A_2266_413#_c_1787_n Q_N 0.0120831f $X=12.25 $Y=1.87 $X2=0 $Y2=0
cc_1234 N_A_2266_413#_M1018_g N_Q_c_2426_n 4.34333e-19 $X=14.74 $Y=0.445 $X2=0
+ $Y2=0
cc_1235 N_A_2266_413#_c_1783_n N_Q_c_2426_n 5.67364e-19 $X=14.865 $Y=1.16 $X2=0
+ $Y2=0
cc_1236 N_A_2266_413#_c_1784_n N_Q_c_2426_n 0.0103604f $X=15.275 $Y=0.995 $X2=0
+ $Y2=0
cc_1237 N_A_2266_413#_c_1792_n N_Q_c_2426_n 0.016307f $X=15.3 $Y=1.41 $X2=0
+ $Y2=0
cc_1238 N_A_2266_413#_c_1793_n N_Q_c_2426_n 0.0152578f $X=15.77 $Y=1.41 $X2=0
+ $Y2=0
cc_1239 N_A_2266_413#_c_1785_n N_Q_c_2426_n 0.003026f $X=15.795 $Y=0.995 $X2=0
+ $Y2=0
cc_1240 N_A_2266_413#_c_1786_n N_Q_c_2426_n 0.0550089f $X=15.77 $Y=1.202 $X2=0
+ $Y2=0
cc_1241 N_A_2266_413#_c_1787_n N_VGND_c_2452_n 0.0166666f $X=12.25 $Y=1.87 $X2=0
+ $Y2=0
cc_1242 N_A_2266_413#_M1018_g N_VGND_c_2454_n 0.00861999f $X=14.74 $Y=0.445
+ $X2=0 $Y2=0
cc_1243 N_A_2266_413#_c_1782_n N_VGND_c_2454_n 0.00620326f $X=15.2 $Y=1.16 $X2=0
+ $Y2=0
cc_1244 N_A_2266_413#_c_1784_n N_VGND_c_2454_n 0.00307023f $X=15.275 $Y=0.995
+ $X2=0 $Y2=0
cc_1245 N_A_2266_413#_c_1785_n N_VGND_c_2455_n 0.00485044f $X=15.795 $Y=0.995
+ $X2=0 $Y2=0
cc_1246 N_A_2266_413#_c_1784_n N_VGND_c_2460_n 0.00541359f $X=15.275 $Y=0.995
+ $X2=0 $Y2=0
cc_1247 N_A_2266_413#_c_1785_n N_VGND_c_2460_n 0.00585385f $X=15.795 $Y=0.995
+ $X2=0 $Y2=0
cc_1248 N_A_2266_413#_c_1805_n N_VGND_c_2466_n 0.0389555f $X=12.125 $Y=0.432
+ $X2=0 $Y2=0
cc_1249 N_A_2266_413#_M1018_g N_VGND_c_2467_n 0.00541359f $X=14.74 $Y=0.445
+ $X2=0 $Y2=0
cc_1250 N_A_2266_413#_M1012_d N_VGND_c_2469_n 0.00365658f $X=11.39 $Y=0.235
+ $X2=0 $Y2=0
cc_1251 N_A_2266_413#_M1018_g N_VGND_c_2469_n 0.0113055f $X=14.74 $Y=0.445 $X2=0
+ $Y2=0
cc_1252 N_A_2266_413#_c_1784_n N_VGND_c_2469_n 0.0100187f $X=15.275 $Y=0.995
+ $X2=0 $Y2=0
cc_1253 N_A_2266_413#_c_1785_n N_VGND_c_2469_n 0.0119211f $X=15.795 $Y=0.995
+ $X2=0 $Y2=0
cc_1254 N_A_2266_413#_c_1805_n N_VGND_c_2469_n 0.0157066f $X=12.125 $Y=0.432
+ $X2=0 $Y2=0
cc_1255 N_A_2266_413#_c_1805_n A_2414_47# 0.00341113f $X=12.125 $Y=0.432
+ $X2=-0.19 $Y2=-0.24
cc_1256 N_A_2266_413#_c_1787_n A_2414_47# 5.79628e-19 $X=12.25 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_1257 N_VPWR_c_1917_n N_A_319_47#_M1023_s 0.00179197f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1258 N_VPWR_c_1917_n N_A_319_47#_M1026_d 0.0022105f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1259 N_VPWR_c_1919_n N_A_319_47#_c_2152_n 0.0176356f $X=2.6 $Y=2 $X2=0 $Y2=0
cc_1260 N_VPWR_c_1937_n N_A_319_47#_c_2152_n 0.0280576f $X=2.385 $Y=2.72 $X2=0
+ $Y2=0
cc_1261 N_VPWR_c_1917_n N_A_319_47#_c_2152_n 0.00773304f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1262 N_VPWR_c_1938_n N_A_319_47#_c_2154_n 0.0238693f $X=6.35 $Y=2.72 $X2=0
+ $Y2=0
cc_1263 N_VPWR_c_1917_n N_A_319_47#_c_2154_n 0.00740377f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1264 N_VPWR_c_1917_n A_409_369# 0.00330845f $X=16.33 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1265 N_VPWR_c_1917_n A_787_369# 0.00546614f $X=16.33 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1266 N_VPWR_c_1917_n N_A_985_47#_M1030_d 0.00236402f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1267 N_VPWR_c_1917_n N_A_985_47#_M1014_d 0.00411682f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1268 N_VPWR_c_1938_n N_A_985_47#_c_2271_n 0.0221045f $X=6.35 $Y=2.72 $X2=0
+ $Y2=0
cc_1269 N_VPWR_c_1917_n N_A_985_47#_c_2271_n 0.0059727f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1270 N_VPWR_c_1922_n N_A_985_47#_c_2286_n 0.0225312f $X=9.36 $Y=2.72 $X2=0
+ $Y2=0
cc_1271 N_VPWR_c_1917_n N_A_985_47#_c_2286_n 0.00594985f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1272 N_VPWR_c_1917_n A_1376_369# 0.00328349f $X=16.33 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1273 N_VPWR_c_1917_n A_1712_413# 0.00261173f $X=16.33 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1274 N_VPWR_c_1917_n A_2165_413# 0.00449658f $X=16.33 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1275 N_VPWR_c_1917_n A_2360_413# 0.00384691f $X=16.33 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1276 N_VPWR_c_1917_n N_Q_N_M1011_s 0.00190235f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_1277 N_VPWR_c_1925_n N_Q_N_c_2398_n 0.0711485f $X=12.68 $Y=1.66 $X2=0 $Y2=0
cc_1278 N_VPWR_c_1926_n N_Q_N_c_2398_n 0.0223557f $X=13.535 $Y=2.72 $X2=0 $Y2=0
cc_1279 N_VPWR_c_1927_n N_Q_N_c_2398_n 0.0610963f $X=13.62 $Y=1.63 $X2=0 $Y2=0
cc_1280 N_VPWR_c_1917_n N_Q_N_c_2398_n 0.00667536f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_1281 N_VPWR_c_1917_n N_Q_M1008_s 0.00234265f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_1282 N_VPWR_c_1928_n N_Q_c_2426_n 0.0730475f $X=15.065 $Y=1.63 $X2=0 $Y2=0
cc_1283 N_VPWR_c_1929_n N_Q_c_2426_n 0.0603669f $X=16.015 $Y=1.63 $X2=0 $Y2=0
cc_1284 N_VPWR_c_1934_n N_Q_c_2426_n 0.0173701f $X=15.92 $Y=2.72 $X2=0 $Y2=0
cc_1285 N_VPWR_c_1917_n N_Q_c_2426_n 0.0136769f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_1286 N_VPWR_c_1925_n N_VGND_c_2452_n 0.0025448f $X=12.68 $Y=1.66 $X2=0 $Y2=0
cc_1287 N_VPWR_c_1927_n N_VGND_c_2453_n 0.0028497f $X=13.62 $Y=1.63 $X2=0 $Y2=0
cc_1288 N_VPWR_c_1928_n N_VGND_c_2454_n 0.00932678f $X=15.065 $Y=1.63 $X2=0
+ $Y2=0
cc_1289 N_VPWR_c_1929_n N_VGND_c_2455_n 0.0104453f $X=16.015 $Y=1.63 $X2=0 $Y2=0
cc_1290 N_A_319_47#_c_2146_n N_A_985_47#_c_2269_n 0.0207307f $X=4.645 $Y=1.82
+ $X2=0 $Y2=0
cc_1291 N_A_319_47#_c_2154_n N_A_985_47#_c_2270_n 0.0207307f $X=4.64 $Y=2 $X2=0
+ $Y2=0
cc_1292 N_A_319_47#_c_2147_n N_A_985_47#_c_2262_n 0.0207307f $X=4.655 $Y=1.15
+ $X2=0 $Y2=0
cc_1293 N_A_319_47#_c_2150_n N_A_985_47#_c_2262_n 0.0063392f $X=4.64 $Y=0.445
+ $X2=0 $Y2=0
cc_1294 N_A_319_47#_c_2176_n N_A_985_47#_c_2265_n 0.0259367f $X=4.62 $Y=0.51
+ $X2=0 $Y2=0
cc_1295 N_A_319_47#_c_2150_n N_A_985_47#_c_2265_n 8.5984e-19 $X=4.64 $Y=0.445
+ $X2=0 $Y2=0
cc_1296 N_A_319_47#_c_2176_n N_A_985_47#_c_2320_n 7.7591e-19 $X=4.62 $Y=0.51
+ $X2=0 $Y2=0
cc_1297 N_A_319_47#_c_2150_n N_A_985_47#_c_2320_n 0.024338f $X=4.64 $Y=0.445
+ $X2=0 $Y2=0
cc_1298 N_A_319_47#_c_2149_n N_VGND_M1045_d 0.00246892f $X=4.425 $Y=0.51 $X2=0
+ $Y2=0
cc_1299 N_A_319_47#_c_2149_n N_VGND_c_2446_n 0.0162997f $X=4.425 $Y=0.51 $X2=0
+ $Y2=0
cc_1300 N_A_319_47#_c_2151_n N_VGND_c_2446_n 0.00382991f $X=1.72 $Y=0.415 $X2=0
+ $Y2=0
cc_1301 N_A_319_47#_c_2149_n N_VGND_c_2447_n 0.00221983f $X=4.425 $Y=0.51 $X2=0
+ $Y2=0
cc_1302 N_A_319_47#_c_2149_n N_VGND_c_2448_n 0.0244754f $X=4.425 $Y=0.51 $X2=0
+ $Y2=0
cc_1303 N_A_319_47#_c_2148_n N_VGND_c_2463_n 6.17783e-19 $X=1.685 $Y=0.51 $X2=0
+ $Y2=0
cc_1304 N_A_319_47#_c_2149_n N_VGND_c_2463_n 0.00254779f $X=4.425 $Y=0.51 $X2=0
+ $Y2=0
cc_1305 N_A_319_47#_c_2151_n N_VGND_c_2463_n 0.0274021f $X=1.72 $Y=0.415 $X2=0
+ $Y2=0
cc_1306 N_A_319_47#_c_2176_n N_VGND_c_2464_n 2.16231e-19 $X=4.62 $Y=0.51 $X2=0
+ $Y2=0
cc_1307 N_A_319_47#_c_2149_n N_VGND_c_2464_n 0.00317176f $X=4.425 $Y=0.51 $X2=0
+ $Y2=0
cc_1308 N_A_319_47#_c_2150_n N_VGND_c_2464_n 0.0186145f $X=4.64 $Y=0.445 $X2=0
+ $Y2=0
cc_1309 N_A_319_47#_M1043_s N_VGND_c_2469_n 0.00141593f $X=1.595 $Y=0.235 $X2=0
+ $Y2=0
cc_1310 N_A_319_47#_M1009_d N_VGND_c_2469_n 0.00123074f $X=4.505 $Y=0.235 $X2=0
+ $Y2=0
cc_1311 N_A_319_47#_c_2148_n N_VGND_c_2469_n 0.329589f $X=1.685 $Y=0.51 $X2=0
+ $Y2=0
cc_1312 N_A_319_47#_c_2150_n N_VGND_c_2469_n 0.00300386f $X=4.64 $Y=0.445 $X2=0
+ $Y2=0
cc_1313 N_A_319_47#_c_2151_n N_VGND_c_2469_n 0.00378066f $X=1.72 $Y=0.415 $X2=0
+ $Y2=0
cc_1314 N_A_319_47#_c_2149_n A_413_47# 0.00649316f $X=4.425 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_1315 N_A_319_47#_c_2149_n A_779_47# 0.00963532f $X=4.425 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_1316 N_A_985_47#_c_2260_n N_VGND_c_2449_n 0.00463496f $X=7.505 $Y=0.98 $X2=0
+ $Y2=0
cc_1317 N_A_985_47#_c_2266_n N_VGND_c_2449_n 9.38714e-19 $X=7.4 $Y=0.51 $X2=0
+ $Y2=0
cc_1318 N_A_985_47#_c_2267_n N_VGND_c_2449_n 0.0191789f $X=7.205 $Y=0.51 $X2=0
+ $Y2=0
cc_1319 N_A_985_47#_c_2268_n N_VGND_c_2449_n 0.00783393f $X=7.755 $Y=0.41 $X2=0
+ $Y2=0
cc_1320 N_A_985_47#_c_2261_n N_VGND_c_2464_n 9.76595e-19 $X=5.125 $Y=0.825 $X2=0
+ $Y2=0
cc_1321 N_A_985_47#_c_2265_n N_VGND_c_2464_n 0.00139545f $X=5.245 $Y=0.51 $X2=0
+ $Y2=0
cc_1322 N_A_985_47#_c_2267_n N_VGND_c_2464_n 0.00170949f $X=7.205 $Y=0.51 $X2=0
+ $Y2=0
cc_1323 N_A_985_47#_c_2320_n N_VGND_c_2464_n 0.0138434f $X=5.11 $Y=0.445 $X2=0
+ $Y2=0
cc_1324 N_A_985_47#_c_2267_n N_VGND_c_2465_n 0.00315872f $X=7.205 $Y=0.51 $X2=0
+ $Y2=0
cc_1325 N_A_985_47#_c_2268_n N_VGND_c_2465_n 0.0410021f $X=7.755 $Y=0.41 $X2=0
+ $Y2=0
cc_1326 N_A_985_47#_M1019_d N_VGND_c_2469_n 0.00166838f $X=4.925 $Y=0.235 $X2=0
+ $Y2=0
cc_1327 N_A_985_47#_M1024_d N_VGND_c_2469_n 0.00412777f $X=7.225 $Y=0.595 $X2=0
+ $Y2=0
cc_1328 N_A_985_47#_c_2265_n N_VGND_c_2469_n 0.259273f $X=5.245 $Y=0.51 $X2=0
+ $Y2=0
cc_1329 N_A_985_47#_c_2320_n N_VGND_c_2469_n 0.00190201f $X=5.11 $Y=0.445 $X2=0
+ $Y2=0
cc_1330 N_A_985_47#_c_2268_n N_VGND_c_2469_n 0.00878695f $X=7.755 $Y=0.41 $X2=0
+ $Y2=0
cc_1331 N_Q_N_c_2396_n N_VGND_c_2452_n 0.00373017f $X=13.265 $Y=0.395 $X2=0
+ $Y2=0
cc_1332 N_Q_N_c_2396_n N_VGND_c_2453_n 0.0388684f $X=13.265 $Y=0.395 $X2=0 $Y2=0
cc_1333 N_Q_N_c_2396_n N_VGND_c_2458_n 0.0197303f $X=13.265 $Y=0.395 $X2=0 $Y2=0
cc_1334 N_Q_N_M1017_s N_VGND_c_2469_n 0.00225609f $X=13.08 $Y=0.235 $X2=0 $Y2=0
cc_1335 N_Q_N_c_2396_n N_VGND_c_2469_n 0.00592003f $X=13.265 $Y=0.395 $X2=0
+ $Y2=0
cc_1336 N_Q_c_2426_n N_VGND_c_2454_n 0.0252834f $X=15.535 $Y=0.395 $X2=0 $Y2=0
cc_1337 N_Q_c_2426_n N_VGND_c_2455_n 9.65365e-19 $X=15.535 $Y=0.395 $X2=0 $Y2=0
cc_1338 N_Q_c_2426_n N_VGND_c_2460_n 0.0232464f $X=15.535 $Y=0.395 $X2=0 $Y2=0
cc_1339 N_Q_M1031_s N_VGND_c_2469_n 0.00364931f $X=15.35 $Y=0.235 $X2=0 $Y2=0
cc_1340 N_Q_c_2426_n N_VGND_c_2469_n 0.0143524f $X=15.535 $Y=0.395 $X2=0 $Y2=0
cc_1341 N_VGND_c_2469_n A_413_47# 0.00154859f $X=16.33 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1342 N_VGND_c_2469_n A_779_47# 0.00333367f $X=16.33 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1343 N_VGND_c_2469_n A_1738_47# 0.00376746f $X=16.33 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1344 N_VGND_c_2469_n A_2181_47# 0.00481883f $X=16.33 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1345 N_VGND_c_2469_n A_2414_47# 0.00235079f $X=16.33 $Y=0 $X2=-0.19 $Y2=-0.24
