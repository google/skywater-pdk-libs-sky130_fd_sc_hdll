* File: sky130_fd_sc_hdll__a31o_4.pxi.spice
* Created: Wed Sep  2 08:20:06 2020
* 
x_PM_SKY130_FD_SC_HDLL__A31O_4%A3 N_A3_c_91_n N_A3_M1002_g N_A3_c_92_n
+ N_A3_M1016_g N_A3_c_93_n N_A3_M1019_g N_A3_c_94_n N_A3_M1007_g N_A3_c_99_n
+ N_A3_c_95_n A3 A3 N_A3_c_96_n PM_SKY130_FD_SC_HDLL__A31O_4%A3
x_PM_SKY130_FD_SC_HDLL__A31O_4%A2 N_A2_c_172_n N_A2_M1000_g N_A2_c_173_n
+ N_A2_M1001_g N_A2_c_174_n N_A2_M1011_g N_A2_c_175_n N_A2_M1014_g N_A2_c_176_n
+ N_A2_c_177_n N_A2_c_178_n A2 A2 N_A2_c_179_n PM_SKY130_FD_SC_HDLL__A31O_4%A2
x_PM_SKY130_FD_SC_HDLL__A31O_4%A1 N_A1_M1005_g N_A1_c_250_n N_A1_M1015_g
+ N_A1_c_251_n N_A1_M1022_g N_A1_M1017_g A1 N_A1_c_249_n
+ PM_SKY130_FD_SC_HDLL__A31O_4%A1
x_PM_SKY130_FD_SC_HDLL__A31O_4%B1 N_B1_c_290_n N_B1_M1012_g N_B1_c_296_n
+ N_B1_M1009_g N_B1_c_291_n N_B1_M1021_g N_B1_c_297_n N_B1_M1018_g N_B1_c_292_n
+ N_B1_c_313_p N_B1_c_293_n B1 B1 N_B1_c_295_n PM_SKY130_FD_SC_HDLL__A31O_4%B1
x_PM_SKY130_FD_SC_HDLL__A31O_4%A_297_47# N_A_297_47#_M1005_s N_A_297_47#_M1012_s
+ N_A_297_47#_M1009_s N_A_297_47#_c_363_n N_A_297_47#_M1003_g
+ N_A_297_47#_c_356_n N_A_297_47#_M1004_g N_A_297_47#_c_364_n
+ N_A_297_47#_M1006_g N_A_297_47#_c_357_n N_A_297_47#_M1008_g
+ N_A_297_47#_c_365_n N_A_297_47#_M1013_g N_A_297_47#_c_358_n
+ N_A_297_47#_M1010_g N_A_297_47#_c_366_n N_A_297_47#_M1020_g
+ N_A_297_47#_c_359_n N_A_297_47#_M1023_g N_A_297_47#_c_383_n
+ N_A_297_47#_c_372_n N_A_297_47#_c_375_n N_A_297_47#_c_360_n
+ N_A_297_47#_c_379_n N_A_297_47#_c_368_n N_A_297_47#_c_361_n
+ N_A_297_47#_c_458_p N_A_297_47#_c_380_n N_A_297_47#_c_415_n
+ N_A_297_47#_c_370_n N_A_297_47#_c_362_n PM_SKY130_FD_SC_HDLL__A31O_4%A_297_47#
x_PM_SKY130_FD_SC_HDLL__A31O_4%A_27_297# N_A_27_297#_M1002_d N_A_27_297#_M1000_d
+ N_A_27_297#_M1022_d N_A_27_297#_M1007_d N_A_27_297#_M1018_d
+ N_A_27_297#_c_512_n N_A_27_297#_c_515_n N_A_27_297#_c_516_n
+ N_A_27_297#_c_519_n N_A_27_297#_c_520_n N_A_27_297#_c_530_n
+ N_A_27_297#_c_521_n N_A_27_297#_c_539_n N_A_27_297#_c_522_n
+ N_A_27_297#_c_524_n N_A_27_297#_c_525_n PM_SKY130_FD_SC_HDLL__A31O_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A31O_4%VPWR N_VPWR_M1002_s N_VPWR_M1015_s N_VPWR_M1011_s
+ N_VPWR_M1003_s N_VPWR_M1006_s N_VPWR_M1020_s N_VPWR_c_574_n N_VPWR_c_575_n
+ N_VPWR_c_576_n N_VPWR_c_577_n N_VPWR_c_578_n N_VPWR_c_579_n N_VPWR_c_580_n
+ N_VPWR_c_581_n N_VPWR_c_582_n N_VPWR_c_583_n N_VPWR_c_584_n VPWR
+ N_VPWR_c_585_n N_VPWR_c_586_n N_VPWR_c_587_n N_VPWR_c_588_n N_VPWR_c_589_n
+ N_VPWR_c_590_n N_VPWR_c_591_n N_VPWR_c_573_n PM_SKY130_FD_SC_HDLL__A31O_4%VPWR
x_PM_SKY130_FD_SC_HDLL__A31O_4%X N_X_M1004_s N_X_M1010_s N_X_M1003_d N_X_M1013_d
+ N_X_c_698_n N_X_c_702_n N_X_c_705_n X X X X N_X_c_693_n X
+ PM_SKY130_FD_SC_HDLL__A31O_4%X
x_PM_SKY130_FD_SC_HDLL__A31O_4%VGND N_VGND_M1016_d N_VGND_M1019_d N_VGND_M1021_d
+ N_VGND_M1008_d N_VGND_M1023_d N_VGND_c_750_n N_VGND_c_751_n N_VGND_c_752_n
+ N_VGND_c_753_n N_VGND_c_754_n N_VGND_c_755_n N_VGND_c_756_n N_VGND_c_757_n
+ VGND N_VGND_c_758_n N_VGND_c_759_n N_VGND_c_760_n N_VGND_c_761_n
+ N_VGND_c_762_n N_VGND_c_763_n PM_SKY130_FD_SC_HDLL__A31O_4%VGND
cc_1 VNB N_A3_c_91_n 0.0361459f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_A3_c_92_n 0.0221349f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_3 VNB N_A3_c_93_n 0.0177217f $X=-0.19 $Y=-0.24 $X2=2.88 $Y2=0.995
cc_4 VNB N_A3_c_94_n 0.0227872f $X=-0.19 $Y=-0.24 $X2=2.905 $Y2=1.41
cc_5 VNB N_A3_c_95_n 0.00396283f $X=-0.19 $Y=-0.24 $X2=2.94 $Y2=1.16
cc_6 VNB N_A3_c_96_n 0.0103665f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_7 VNB N_A2_c_172_n 0.0220745f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_8 VNB N_A2_c_173_n 0.0156441f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_9 VNB N_A2_c_174_n 0.0234647f $X=-0.19 $Y=-0.24 $X2=2.88 $Y2=0.995
cc_10 VNB N_A2_c_175_n 0.0168332f $X=-0.19 $Y=-0.24 $X2=2.905 $Y2=1.41
cc_11 VNB N_A2_c_176_n 0.00671002f $X=-0.19 $Y=-0.24 $X2=2.775 $Y2=1.53
cc_12 VNB N_A2_c_177_n 0.00173313f $X=-0.19 $Y=-0.24 $X2=2.94 $Y2=1.16
cc_13 VNB N_A2_c_178_n 0.00392492f $X=-0.19 $Y=-0.24 $X2=2.965 $Y2=1.53
cc_14 VNB N_A2_c_179_n 0.00796308f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A1_M1005_g 0.0185044f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_16 VNB N_A1_M1017_g 0.0189364f $X=-0.19 $Y=-0.24 $X2=2.775 $Y2=1.53
cc_17 VNB N_A1_c_249_n 0.0403121f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_18 VNB N_B1_c_290_n 0.0172134f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_19 VNB N_B1_c_291_n 0.0198684f $X=-0.19 $Y=-0.24 $X2=2.88 $Y2=0.995
cc_20 VNB N_B1_c_292_n 0.0349501f $X=-0.19 $Y=-0.24 $X2=2.775 $Y2=1.53
cc_21 VNB N_B1_c_293_n 0.0321423f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_22 VNB B1 0.00318716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_B1_c_295_n 0.00281408f $X=-0.19 $Y=-0.24 $X2=0.335 $Y2=1.16
cc_24 VNB N_A_297_47#_c_356_n 0.0201722f $X=-0.19 $Y=-0.24 $X2=2.775 $Y2=1.53
cc_25 VNB N_A_297_47#_c_357_n 0.0164634f $X=-0.19 $Y=-0.24 $X2=2.965 $Y2=1.53
cc_26 VNB N_A_297_47#_c_358_n 0.0169705f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_27 VNB N_A_297_47#_c_359_n 0.0186035f $X=-0.19 $Y=-0.24 $X2=0.335 $Y2=1.19
cc_28 VNB N_A_297_47#_c_360_n 9.7053e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_297_47#_c_361_n 0.00872112f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_297_47#_c_362_n 0.0821127f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_573_n 0.288713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_X_c_693_n 0.0089973f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB X 0.0231184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_750_n 0.0110531f $X=-0.19 $Y=-0.24 $X2=2.94 $Y2=1.16
cc_35 VNB N_VGND_c_751_n 0.00682035f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_752_n 0.00293557f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_37 VNB N_VGND_c_753_n 0.00214417f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_38 VNB N_VGND_c_754_n 0.0138375f $X=-0.19 $Y=-0.24 $X2=2.965 $Y2=1.16
cc_39 VNB N_VGND_c_755_n 0.0128151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_756_n 0.0197881f $X=-0.19 $Y=-0.24 $X2=0.335 $Y2=1.53
cc_41 VNB N_VGND_c_757_n 0.00573782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_758_n 0.0692035f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_759_n 0.0230558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_760_n 0.0143274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_761_n 0.00531951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_762_n 0.016985f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_763_n 0.336125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VPB N_A3_c_91_n 0.0319872f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_49 VPB N_A3_c_94_n 0.0261522f $X=-0.19 $Y=1.305 $X2=2.905 $Y2=1.41
cc_50 VPB N_A3_c_99_n 0.0197497f $X=-0.19 $Y=1.305 $X2=2.775 $Y2=1.53
cc_51 VPB N_A3_c_95_n 0.00306676f $X=-0.19 $Y=1.305 $X2=2.94 $Y2=1.16
cc_52 VPB N_A3_c_96_n 0.00682521f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_53 VPB N_A2_c_172_n 0.0255737f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_54 VPB N_A2_c_174_n 0.0259688f $X=-0.19 $Y=1.305 $X2=2.88 $Y2=0.995
cc_55 VPB N_A1_c_250_n 0.015555f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_56 VPB N_A1_c_251_n 0.0158343f $X=-0.19 $Y=1.305 $X2=2.88 $Y2=0.56
cc_57 VPB N_A1_c_249_n 0.0129133f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_58 VPB N_B1_c_296_n 0.0165222f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_59 VPB N_B1_c_297_n 0.0195993f $X=-0.19 $Y=1.305 $X2=2.905 $Y2=1.41
cc_60 VPB N_B1_c_292_n 0.0217433f $X=-0.19 $Y=1.305 $X2=2.775 $Y2=1.53
cc_61 VPB N_A_297_47#_c_363_n 0.0187827f $X=-0.19 $Y=1.305 $X2=2.905 $Y2=1.41
cc_62 VPB N_A_297_47#_c_364_n 0.0158086f $X=-0.19 $Y=1.305 $X2=2.94 $Y2=1.16
cc_63 VPB N_A_297_47#_c_365_n 0.0160912f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_64 VPB N_A_297_47#_c_366_n 0.0181162f $X=-0.19 $Y=1.305 $X2=2.965 $Y2=1.16
cc_65 VPB N_A_297_47#_c_360_n 0.00124954f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_297_47#_c_368_n 0.0201957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_297_47#_c_361_n 0.00226921f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_297_47#_c_370_n 0.00103601f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_297_47#_c_362_n 0.0534932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_574_n 4.04661e-19 $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_71 VPB N_VPWR_c_575_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_72 VPB N_VPWR_c_576_n 0.00277739f $X=-0.19 $Y=1.305 $X2=0.335 $Y2=1.16
cc_73 VPB N_VPWR_c_577_n 0.00702898f $X=-0.19 $Y=1.305 $X2=0.335 $Y2=1.53
cc_74 VPB N_VPWR_c_578_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_579_n 0.0139576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_580_n 0.0172009f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_581_n 0.0439436f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_582_n 0.00513801f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_583_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_584_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_585_n 0.0159043f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_586_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_587_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_588_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_589_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_590_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_591_n 0.00580385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_573_n 0.0569477f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB X 0.00912754f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_90 VPB X 0.0209855f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 N_A3_c_91_n N_A2_c_172_n 0.0616598f $X=0.495 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_92 N_A3_c_99_n N_A2_c_172_n 0.0152534f $X=2.775 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_93 N_A3_c_96_n N_A2_c_172_n 0.00127905f $X=0.36 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_94 N_A3_c_92_n N_A2_c_173_n 0.0348584f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A3_c_94_n N_A2_c_174_n 0.0534287f $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A3_c_99_n N_A2_c_174_n 0.0152708f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_97 N_A3_c_95_n N_A2_c_174_n 0.00455123f $X=2.94 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A3_c_93_n N_A2_c_175_n 0.0310384f $X=2.88 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A3_c_99_n N_A2_c_176_n 0.0159379f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_100 N_A3_c_93_n N_A2_c_177_n 8.37473e-19 $X=2.88 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A3_c_94_n N_A2_c_178_n 6.942e-19 $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A3_c_99_n N_A2_c_178_n 0.0270622f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_103 N_A3_c_95_n N_A2_c_178_n 0.0145726f $X=2.94 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A3_c_92_n N_A2_c_179_n 0.00735811f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A3_c_99_n N_A2_c_179_n 0.0375279f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_106 N_A3_c_96_n N_A2_c_179_n 0.0123636f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A3_c_99_n N_A1_c_250_n 0.0132009f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_108 N_A3_c_99_n N_A1_c_251_n 0.0135647f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_109 N_A3_c_99_n A1 0.0285404f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_110 N_A3_c_99_n N_A1_c_249_n 0.00767784f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_111 N_A3_c_93_n N_B1_c_290_n 0.0222991f $X=2.88 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_112 N_A3_c_94_n N_B1_c_296_n 0.0269891f $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A3_c_95_n N_B1_c_296_n 0.00169995f $X=2.94 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A3_c_94_n N_B1_c_292_n 0.0252561f $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A3_c_95_n N_B1_c_292_n 0.00269313f $X=2.94 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A3_c_93_n N_A_297_47#_c_372_n 0.0115038f $X=2.88 $Y=0.995 $X2=0 $Y2=0
cc_117 N_A3_c_94_n N_A_297_47#_c_372_n 0.00410811f $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A3_c_95_n N_A_297_47#_c_372_n 0.022384f $X=2.94 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A3_c_93_n N_A_297_47#_c_375_n 9.57275e-19 $X=2.88 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A3_c_93_n N_A_297_47#_c_360_n 5.82448e-19 $X=2.88 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A3_c_94_n N_A_297_47#_c_360_n 8.04969e-19 $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A3_c_95_n N_A_297_47#_c_360_n 0.019459f $X=2.94 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A3_c_94_n N_A_297_47#_c_379_n 9.54699e-19 $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A3_c_99_n N_A_297_47#_c_380_n 0.005232f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_125 N_A3_c_95_n N_A_297_47#_c_370_n 0.00864607f $X=2.94 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A3_c_96_n N_A_27_297#_M1002_d 0.00904073f $X=0.36 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_127 N_A3_c_99_n N_A_27_297#_M1000_d 0.00180713f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_128 N_A3_c_99_n N_A_27_297#_M1022_d 0.00180713f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_129 N_A3_c_95_n N_A_27_297#_M1007_d 0.00253723f $X=2.94 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A3_c_91_n N_A_27_297#_c_512_n 0.0106355f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A3_c_99_n N_A_27_297#_c_512_n 0.0291258f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_132 N_A3_c_96_n N_A_27_297#_c_512_n 0.00898813f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A3_c_99_n N_A_27_297#_c_515_n 0.0373345f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_134 N_A3_c_94_n N_A_27_297#_c_516_n 0.0139214f $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A3_c_99_n N_A_27_297#_c_516_n 0.029417f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_136 N_A3_c_95_n N_A_27_297#_c_516_n 0.0184442f $X=2.94 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A3_c_95_n N_A_27_297#_c_519_n 0.00345721f $X=2.94 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A3_c_94_n N_A_27_297#_c_520_n 0.00544471f $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A3_c_94_n N_A_27_297#_c_521_n 0.00186382f $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A3_c_91_n N_A_27_297#_c_522_n 5.03339e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A3_c_96_n N_A_27_297#_c_522_n 0.0150699f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A3_c_99_n N_A_27_297#_c_524_n 0.013831f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_143 N_A3_c_99_n N_A_27_297#_c_525_n 0.013831f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_144 N_A3_c_99_n N_VPWR_M1002_s 0.00187547f $X=2.775 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_145 N_A3_c_99_n N_VPWR_M1015_s 0.00187547f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_146 N_A3_c_99_n N_VPWR_M1011_s 0.00251484f $X=2.775 $Y=1.53 $X2=0 $Y2=0
cc_147 N_A3_c_91_n N_VPWR_c_574_n 0.0138595f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A3_c_94_n N_VPWR_c_576_n 0.00508294f $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A3_c_94_n N_VPWR_c_581_n 0.00702461f $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A3_c_91_n N_VPWR_c_585_n 0.00427505f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A3_c_91_n N_VPWR_c_573_n 0.00485802f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A3_c_94_n N_VPWR_c_573_n 0.0074134f $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A3_c_91_n N_VGND_c_751_n 0.00305311f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A3_c_92_n N_VGND_c_751_n 0.0146609f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A3_c_96_n N_VGND_c_751_n 0.0149476f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A3_c_93_n N_VGND_c_752_n 0.0121748f $X=2.88 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A3_c_92_n N_VGND_c_758_n 0.00585385f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A3_c_93_n N_VGND_c_758_n 0.00419163f $X=2.88 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A3_c_92_n N_VGND_c_763_n 0.0118856f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A3_c_93_n N_VGND_c_763_n 0.00502958f $X=2.88 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A2_c_172_n N_A1_M1005_g 0.0217285f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A2_c_173_n N_A1_M1005_g 0.0439542f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A2_c_176_n N_A1_M1005_g 0.0127248f $X=2.185 $Y=0.82 $X2=0 $Y2=0
cc_164 N_A2_c_179_n N_A1_M1005_g 0.00675544f $X=1.015 $Y=0.82 $X2=0 $Y2=0
cc_165 N_A2_c_172_n N_A1_c_250_n 0.0224794f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A2_c_174_n N_A1_c_251_n 0.0224794f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A2_c_174_n N_A1_M1017_g 0.0219835f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A2_c_175_n N_A1_M1017_g 0.0357406f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A2_c_176_n N_A1_M1017_g 0.0128837f $X=2.185 $Y=0.82 $X2=0 $Y2=0
cc_170 N_A2_c_177_n N_A1_M1017_g 0.00353848f $X=2.277 $Y=1.075 $X2=0 $Y2=0
cc_171 N_A2_c_176_n A1 0.0288426f $X=2.185 $Y=0.82 $X2=0 $Y2=0
cc_172 N_A2_c_178_n A1 0.00985923f $X=2.35 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A2_c_179_n A1 0.0145535f $X=1.015 $Y=0.82 $X2=0 $Y2=0
cc_174 N_A2_c_172_n N_A1_c_249_n 0.00466095f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A2_c_174_n N_A1_c_249_n 0.00466095f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A2_c_176_n N_A1_c_249_n 0.00433688f $X=2.185 $Y=0.82 $X2=0 $Y2=0
cc_177 N_A2_c_178_n N_A1_c_249_n 0.00163312f $X=2.35 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A2_c_176_n N_A_297_47#_M1005_s 0.00274732f $X=2.185 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_179 N_A2_c_173_n N_A_297_47#_c_383_n 8.22884e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A2_c_174_n N_A_297_47#_c_383_n 0.0012867f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A2_c_175_n N_A_297_47#_c_383_n 0.0113149f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A2_c_176_n N_A_297_47#_c_383_n 0.0474694f $X=2.185 $Y=0.82 $X2=0 $Y2=0
cc_183 N_A2_c_178_n N_A_297_47#_c_383_n 0.00489356f $X=2.35 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A2_c_175_n N_A_297_47#_c_380_n 0.00506771f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A2_c_176_n N_A_297_47#_c_380_n 0.00839452f $X=2.185 $Y=0.82 $X2=0 $Y2=0
cc_186 N_A2_c_172_n N_A_27_297#_c_512_n 0.0110707f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_187 N_A2_c_174_n N_A_27_297#_c_516_n 0.0109757f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A2_c_172_n N_VPWR_c_574_n 0.0092641f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A2_c_172_n N_VPWR_c_575_n 5.73683e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_190 N_A2_c_174_n N_VPWR_c_575_n 5.29587e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_191 N_A2_c_174_n N_VPWR_c_576_n 0.0122152f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_192 N_A2_c_172_n N_VPWR_c_586_n 0.00622633f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A2_c_174_n N_VPWR_c_587_n 0.00427505f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A2_c_172_n N_VPWR_c_573_n 0.00550537f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A2_c_174_n N_VPWR_c_573_n 0.0039718f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A2_c_179_n N_VGND_c_751_n 0.00680222f $X=1.015 $Y=0.82 $X2=0 $Y2=0
cc_197 N_A2_c_175_n N_VGND_c_752_n 0.00165449f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A2_c_173_n N_VGND_c_758_n 0.00439071f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A2_c_175_n N_VGND_c_758_n 0.00385416f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A2_c_176_n N_VGND_c_758_n 0.00233008f $X=2.185 $Y=0.82 $X2=0 $Y2=0
cc_201 N_A2_c_179_n N_VGND_c_758_n 0.00630807f $X=1.015 $Y=0.82 $X2=0 $Y2=0
cc_202 N_A2_c_173_n N_VGND_c_763_n 0.00630006f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A2_c_175_n N_VGND_c_763_n 0.00570859f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A2_c_176_n N_VGND_c_763_n 0.00579003f $X=2.185 $Y=0.82 $X2=0 $Y2=0
cc_205 N_A2_c_179_n N_VGND_c_763_n 0.0124413f $X=1.015 $Y=0.82 $X2=0 $Y2=0
cc_206 N_A2_c_179_n A_119_47# 0.00357645f $X=1.015 $Y=0.82 $X2=-0.19 $Y2=-0.24
cc_207 N_A2_c_176_n A_213_47# 8.08198e-19 $X=2.185 $Y=0.82 $X2=-0.19 $Y2=-0.24
cc_208 N_A2_c_179_n A_213_47# 0.00301714f $X=1.015 $Y=0.82 $X2=-0.19 $Y2=-0.24
cc_209 N_A2_c_176_n A_401_47# 0.00213995f $X=2.185 $Y=0.82 $X2=-0.19 $Y2=-0.24
cc_210 N_A1_M1005_g N_A_297_47#_c_383_n 0.00417689f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_211 N_A1_M1017_g N_A_297_47#_c_383_n 0.0087553f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_212 N_A1_c_250_n N_A_27_297#_c_515_n 0.0106972f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_213 N_A1_c_251_n N_A_27_297#_c_515_n 0.0111137f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A1_c_250_n N_VPWR_c_574_n 5.29587e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A1_c_250_n N_VPWR_c_575_n 0.0122621f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A1_c_251_n N_VPWR_c_575_n 0.00931793f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_217 N_A1_c_251_n N_VPWR_c_576_n 5.73683e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A1_c_250_n N_VPWR_c_586_n 0.00427505f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_219 N_A1_c_251_n N_VPWR_c_587_n 0.00622633f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_220 N_A1_c_250_n N_VPWR_c_573_n 0.0039718f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_221 N_A1_c_251_n N_VPWR_c_573_n 0.00550537f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_222 N_A1_M1005_g N_VGND_c_758_n 0.00428448f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_223 N_A1_M1017_g N_VGND_c_758_n 0.00385416f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_224 N_A1_M1005_g N_VGND_c_763_n 0.00625518f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_225 N_A1_M1017_g N_VGND_c_763_n 0.00578596f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_226 B1 N_A_297_47#_c_356_n 0.00617258f $X=4.23 $Y=0.765 $X2=0 $Y2=0
cc_227 N_B1_c_290_n N_A_297_47#_c_372_n 0.0125447f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_228 N_B1_c_290_n N_A_297_47#_c_375_n 0.00623123f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_229 N_B1_c_291_n N_A_297_47#_c_375_n 0.0101243f $X=3.88 $Y=0.995 $X2=0 $Y2=0
cc_230 N_B1_c_290_n N_A_297_47#_c_360_n 0.00344877f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_231 N_B1_c_296_n N_A_297_47#_c_360_n 0.0010867f $X=3.435 $Y=1.41 $X2=0 $Y2=0
cc_232 N_B1_c_291_n N_A_297_47#_c_360_n 0.00133936f $X=3.88 $Y=0.995 $X2=0 $Y2=0
cc_233 N_B1_c_297_n N_A_297_47#_c_360_n 0.00104655f $X=3.905 $Y=1.41 $X2=0 $Y2=0
cc_234 N_B1_c_292_n N_A_297_47#_c_360_n 0.0293747f $X=4.005 $Y=1.16 $X2=0 $Y2=0
cc_235 N_B1_c_313_p N_A_297_47#_c_360_n 0.0124749f $X=4.215 $Y=1.18 $X2=0 $Y2=0
cc_236 B1 N_A_297_47#_c_360_n 0.00686896f $X=4.23 $Y=0.765 $X2=0 $Y2=0
cc_237 N_B1_c_296_n N_A_297_47#_c_379_n 0.00948509f $X=3.435 $Y=1.41 $X2=0 $Y2=0
cc_238 N_B1_c_297_n N_A_297_47#_c_379_n 0.0117744f $X=3.905 $Y=1.41 $X2=0 $Y2=0
cc_239 N_B1_c_297_n N_A_297_47#_c_368_n 0.0159635f $X=3.905 $Y=1.41 $X2=0 $Y2=0
cc_240 N_B1_c_292_n N_A_297_47#_c_368_n 2.68516e-19 $X=4.005 $Y=1.16 $X2=0 $Y2=0
cc_241 N_B1_c_313_p N_A_297_47#_c_368_n 0.0207343f $X=4.215 $Y=1.18 $X2=0 $Y2=0
cc_242 N_B1_c_293_n N_A_297_47#_c_368_n 0.00651034f $X=4.14 $Y=1.16 $X2=0 $Y2=0
cc_243 N_B1_c_295_n N_A_297_47#_c_368_n 0.0194532f $X=4.335 $Y=1.075 $X2=0 $Y2=0
cc_244 N_B1_c_297_n N_A_297_47#_c_361_n 0.00126653f $X=3.905 $Y=1.41 $X2=0 $Y2=0
cc_245 N_B1_c_292_n N_A_297_47#_c_361_n 0.00259612f $X=4.005 $Y=1.16 $X2=0 $Y2=0
cc_246 N_B1_c_293_n N_A_297_47#_c_361_n 8.66819e-19 $X=4.14 $Y=1.16 $X2=0 $Y2=0
cc_247 B1 N_A_297_47#_c_361_n 0.00558062f $X=4.23 $Y=0.765 $X2=0 $Y2=0
cc_248 N_B1_c_295_n N_A_297_47#_c_361_n 0.0157706f $X=4.335 $Y=1.075 $X2=0 $Y2=0
cc_249 N_B1_c_290_n N_A_297_47#_c_415_n 4.64231e-19 $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_250 N_B1_c_291_n N_A_297_47#_c_415_n 0.00388853f $X=3.88 $Y=0.995 $X2=0 $Y2=0
cc_251 N_B1_c_292_n N_A_297_47#_c_415_n 5.69051e-19 $X=4.005 $Y=1.16 $X2=0 $Y2=0
cc_252 B1 N_A_297_47#_c_415_n 0.00493855f $X=4.23 $Y=0.765 $X2=0 $Y2=0
cc_253 N_B1_c_296_n N_A_297_47#_c_370_n 0.00333566f $X=3.435 $Y=1.41 $X2=0 $Y2=0
cc_254 N_B1_c_297_n N_A_297_47#_c_370_n 0.00119404f $X=3.905 $Y=1.41 $X2=0 $Y2=0
cc_255 N_B1_c_292_n N_A_297_47#_c_370_n 0.00421912f $X=4.005 $Y=1.16 $X2=0 $Y2=0
cc_256 N_B1_c_293_n N_A_297_47#_c_362_n 0.00631965f $X=4.14 $Y=1.16 $X2=0 $Y2=0
cc_257 B1 N_A_297_47#_c_362_n 3.10443e-19 $X=4.23 $Y=0.765 $X2=0 $Y2=0
cc_258 N_B1_c_295_n N_A_297_47#_c_362_n 7.16737e-19 $X=4.335 $Y=1.075 $X2=0
+ $Y2=0
cc_259 N_B1_c_296_n N_A_27_297#_c_530_n 0.0122328f $X=3.435 $Y=1.41 $X2=0 $Y2=0
cc_260 N_B1_c_297_n N_A_27_297#_c_530_n 0.0112564f $X=3.905 $Y=1.41 $X2=0 $Y2=0
cc_261 N_B1_c_297_n N_VPWR_c_577_n 0.00233477f $X=3.905 $Y=1.41 $X2=0 $Y2=0
cc_262 N_B1_c_296_n N_VPWR_c_581_n 0.00429453f $X=3.435 $Y=1.41 $X2=0 $Y2=0
cc_263 N_B1_c_297_n N_VPWR_c_581_n 0.00429453f $X=3.905 $Y=1.41 $X2=0 $Y2=0
cc_264 N_B1_c_296_n N_VPWR_c_573_n 0.00622611f $X=3.435 $Y=1.41 $X2=0 $Y2=0
cc_265 N_B1_c_297_n N_VPWR_c_573_n 0.00734734f $X=3.905 $Y=1.41 $X2=0 $Y2=0
cc_266 B1 X 0.00298276f $X=4.23 $Y=0.765 $X2=0 $Y2=0
cc_267 B1 N_VGND_M1021_d 0.0077898f $X=4.23 $Y=0.765 $X2=0 $Y2=0
cc_268 N_B1_c_290_n N_VGND_c_752_n 0.00304107f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_269 N_B1_c_290_n N_VGND_c_759_n 0.00422176f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_270 N_B1_c_291_n N_VGND_c_759_n 0.00542953f $X=3.88 $Y=0.995 $X2=0 $Y2=0
cc_271 N_B1_c_291_n N_VGND_c_762_n 0.0117864f $X=3.88 $Y=0.995 $X2=0 $Y2=0
cc_272 N_B1_c_313_p N_VGND_c_762_n 0.00267041f $X=4.215 $Y=1.18 $X2=0 $Y2=0
cc_273 N_B1_c_293_n N_VGND_c_762_n 0.00190917f $X=4.14 $Y=1.16 $X2=0 $Y2=0
cc_274 B1 N_VGND_c_762_n 0.0193611f $X=4.23 $Y=0.765 $X2=0 $Y2=0
cc_275 N_B1_c_290_n N_VGND_c_763_n 0.00607052f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_276 N_B1_c_291_n N_VGND_c_763_n 0.0112069f $X=3.88 $Y=0.995 $X2=0 $Y2=0
cc_277 B1 N_VGND_c_763_n 0.00100025f $X=4.23 $Y=0.765 $X2=0 $Y2=0
cc_278 N_A_297_47#_c_368_n N_A_27_297#_M1018_d 0.00404268f $X=4.65 $Y=1.54 $X2=0
+ $Y2=0
cc_279 N_A_297_47#_c_379_n N_A_27_297#_c_519_n 0.0141783f $X=3.67 $Y=1.63 $X2=0
+ $Y2=0
cc_280 N_A_297_47#_c_379_n N_A_27_297#_c_520_n 0.0119085f $X=3.67 $Y=1.63 $X2=0
+ $Y2=0
cc_281 N_A_297_47#_M1009_s N_A_27_297#_c_530_n 0.00356935f $X=3.525 $Y=1.485
+ $X2=0 $Y2=0
cc_282 N_A_297_47#_c_363_n N_A_27_297#_c_530_n 5.00696e-19 $X=4.895 $Y=1.41
+ $X2=0 $Y2=0
cc_283 N_A_297_47#_c_379_n N_A_27_297#_c_530_n 0.0186403f $X=3.67 $Y=1.63 $X2=0
+ $Y2=0
cc_284 N_A_297_47#_c_368_n N_A_27_297#_c_530_n 0.00346334f $X=4.65 $Y=1.54 $X2=0
+ $Y2=0
cc_285 N_A_297_47#_c_363_n N_A_27_297#_c_539_n 0.00626522f $X=4.895 $Y=1.41
+ $X2=0 $Y2=0
cc_286 N_A_297_47#_c_379_n N_A_27_297#_c_539_n 0.0195867f $X=3.67 $Y=1.63 $X2=0
+ $Y2=0
cc_287 N_A_297_47#_c_368_n N_A_27_297#_c_539_n 0.0136517f $X=4.65 $Y=1.54 $X2=0
+ $Y2=0
cc_288 N_A_297_47#_c_368_n N_VPWR_M1003_s 0.00299939f $X=4.65 $Y=1.54 $X2=0
+ $Y2=0
cc_289 N_A_297_47#_c_361_n N_VPWR_M1003_s 0.00221654f $X=4.82 $Y=1.16 $X2=0
+ $Y2=0
cc_290 N_A_297_47#_c_363_n N_VPWR_c_577_n 0.0113301f $X=4.895 $Y=1.41 $X2=0
+ $Y2=0
cc_291 N_A_297_47#_c_364_n N_VPWR_c_577_n 5.27036e-19 $X=5.365 $Y=1.41 $X2=0
+ $Y2=0
cc_292 N_A_297_47#_c_368_n N_VPWR_c_577_n 0.0057537f $X=4.65 $Y=1.54 $X2=0 $Y2=0
cc_293 N_A_297_47#_c_361_n N_VPWR_c_577_n 0.00435779f $X=4.82 $Y=1.16 $X2=0
+ $Y2=0
cc_294 N_A_297_47#_c_363_n N_VPWR_c_578_n 5.73683e-19 $X=4.895 $Y=1.41 $X2=0
+ $Y2=0
cc_295 N_A_297_47#_c_364_n N_VPWR_c_578_n 0.0122621f $X=5.365 $Y=1.41 $X2=0
+ $Y2=0
cc_296 N_A_297_47#_c_365_n N_VPWR_c_578_n 0.00931793f $X=5.835 $Y=1.41 $X2=0
+ $Y2=0
cc_297 N_A_297_47#_c_366_n N_VPWR_c_578_n 5.29587e-19 $X=6.305 $Y=1.41 $X2=0
+ $Y2=0
cc_298 N_A_297_47#_c_365_n N_VPWR_c_580_n 5.73683e-19 $X=5.835 $Y=1.41 $X2=0
+ $Y2=0
cc_299 N_A_297_47#_c_366_n N_VPWR_c_580_n 0.0139334f $X=6.305 $Y=1.41 $X2=0
+ $Y2=0
cc_300 N_A_297_47#_c_363_n N_VPWR_c_583_n 0.00622633f $X=4.895 $Y=1.41 $X2=0
+ $Y2=0
cc_301 N_A_297_47#_c_364_n N_VPWR_c_583_n 0.00427505f $X=5.365 $Y=1.41 $X2=0
+ $Y2=0
cc_302 N_A_297_47#_c_365_n N_VPWR_c_588_n 0.00622633f $X=5.835 $Y=1.41 $X2=0
+ $Y2=0
cc_303 N_A_297_47#_c_366_n N_VPWR_c_588_n 0.00427505f $X=6.305 $Y=1.41 $X2=0
+ $Y2=0
cc_304 N_A_297_47#_M1009_s N_VPWR_c_573_n 0.00232895f $X=3.525 $Y=1.485 $X2=0
+ $Y2=0
cc_305 N_A_297_47#_c_363_n N_VPWR_c_573_n 0.00889328f $X=4.895 $Y=1.41 $X2=0
+ $Y2=0
cc_306 N_A_297_47#_c_364_n N_VPWR_c_573_n 0.00394659f $X=5.365 $Y=1.41 $X2=0
+ $Y2=0
cc_307 N_A_297_47#_c_365_n N_VPWR_c_573_n 0.00548015f $X=5.835 $Y=1.41 $X2=0
+ $Y2=0
cc_308 N_A_297_47#_c_366_n N_VPWR_c_573_n 0.00394659f $X=6.305 $Y=1.41 $X2=0
+ $Y2=0
cc_309 N_A_297_47#_c_364_n N_X_c_698_n 0.0124816f $X=5.365 $Y=1.41 $X2=0 $Y2=0
cc_310 N_A_297_47#_c_365_n N_X_c_698_n 0.0128982f $X=5.835 $Y=1.41 $X2=0 $Y2=0
cc_311 N_A_297_47#_c_458_p N_X_c_698_n 0.0213602f $X=6.06 $Y=1.16 $X2=0 $Y2=0
cc_312 N_A_297_47#_c_362_n N_X_c_698_n 0.00495647f $X=6.305 $Y=1.202 $X2=0 $Y2=0
cc_313 N_A_297_47#_c_363_n N_X_c_702_n 0.0106472f $X=4.895 $Y=1.41 $X2=0 $Y2=0
cc_314 N_A_297_47#_c_458_p N_X_c_702_n 0.00913747f $X=6.06 $Y=1.16 $X2=0 $Y2=0
cc_315 N_A_297_47#_c_362_n N_X_c_702_n 0.00429043f $X=6.305 $Y=1.202 $X2=0 $Y2=0
cc_316 N_A_297_47#_c_458_p N_X_c_705_n 0.00649754f $X=6.06 $Y=1.16 $X2=0 $Y2=0
cc_317 N_A_297_47#_c_362_n N_X_c_705_n 0.0033896f $X=6.305 $Y=1.202 $X2=0 $Y2=0
cc_318 N_A_297_47#_c_356_n X 0.00970467f $X=4.92 $Y=0.995 $X2=0 $Y2=0
cc_319 N_A_297_47#_c_357_n X 0.00932305f $X=5.39 $Y=0.995 $X2=0 $Y2=0
cc_320 N_A_297_47#_c_358_n X 0.0101325f $X=5.86 $Y=0.995 $X2=0 $Y2=0
cc_321 N_A_297_47#_c_359_n X 0.01215f $X=6.33 $Y=0.995 $X2=0 $Y2=0
cc_322 N_A_297_47#_c_458_p X 0.0933211f $X=6.06 $Y=1.16 $X2=0 $Y2=0
cc_323 N_A_297_47#_c_362_n X 0.00941663f $X=6.305 $Y=1.202 $X2=0 $Y2=0
cc_324 N_A_297_47#_c_366_n X 0.0148171f $X=6.305 $Y=1.41 $X2=0 $Y2=0
cc_325 N_A_297_47#_c_458_p X 0.00544776f $X=6.06 $Y=1.16 $X2=0 $Y2=0
cc_326 N_A_297_47#_c_366_n X 0.0129979f $X=6.305 $Y=1.41 $X2=0 $Y2=0
cc_327 N_A_297_47#_c_359_n X 0.0177202f $X=6.33 $Y=0.995 $X2=0 $Y2=0
cc_328 N_A_297_47#_c_458_p X 0.0210694f $X=6.06 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A_297_47#_c_372_n N_VGND_M1019_d 0.00900157f $X=3.455 $Y=0.785 $X2=0
+ $Y2=0
cc_330 N_A_297_47#_c_372_n N_VGND_c_752_n 0.0209753f $X=3.455 $Y=0.785 $X2=0
+ $Y2=0
cc_331 N_A_297_47#_c_356_n N_VGND_c_753_n 0.00240574f $X=4.92 $Y=0.995 $X2=0
+ $Y2=0
cc_332 N_A_297_47#_c_357_n N_VGND_c_753_n 0.013167f $X=5.39 $Y=0.995 $X2=0 $Y2=0
cc_333 N_A_297_47#_c_358_n N_VGND_c_753_n 0.00162962f $X=5.86 $Y=0.995 $X2=0
+ $Y2=0
cc_334 N_A_297_47#_c_358_n N_VGND_c_755_n 0.00132036f $X=5.86 $Y=0.995 $X2=0
+ $Y2=0
cc_335 N_A_297_47#_c_359_n N_VGND_c_755_n 0.0128441f $X=6.33 $Y=0.995 $X2=0
+ $Y2=0
cc_336 N_A_297_47#_c_356_n N_VGND_c_756_n 0.00490967f $X=4.92 $Y=0.995 $X2=0
+ $Y2=0
cc_337 N_A_297_47#_c_357_n N_VGND_c_756_n 0.00199015f $X=5.39 $Y=0.995 $X2=0
+ $Y2=0
cc_338 N_A_297_47#_c_383_n N_VGND_c_758_n 0.0337641f $X=2.6 $Y=0.48 $X2=0 $Y2=0
cc_339 N_A_297_47#_c_372_n N_VGND_c_758_n 0.00233045f $X=3.455 $Y=0.785 $X2=0
+ $Y2=0
cc_340 N_A_297_47#_c_380_n N_VGND_c_758_n 0.00567506f $X=2.685 $Y=0.48 $X2=0
+ $Y2=0
cc_341 N_A_297_47#_c_372_n N_VGND_c_759_n 0.00209524f $X=3.455 $Y=0.785 $X2=0
+ $Y2=0
cc_342 N_A_297_47#_c_375_n N_VGND_c_759_n 0.0177822f $X=3.67 $Y=0.38 $X2=0 $Y2=0
cc_343 N_A_297_47#_c_358_n N_VGND_c_760_n 0.00428022f $X=5.86 $Y=0.995 $X2=0
+ $Y2=0
cc_344 N_A_297_47#_c_359_n N_VGND_c_760_n 0.00199015f $X=6.33 $Y=0.995 $X2=0
+ $Y2=0
cc_345 N_A_297_47#_c_356_n N_VGND_c_762_n 0.0165399f $X=4.92 $Y=0.995 $X2=0
+ $Y2=0
cc_346 N_A_297_47#_c_375_n N_VGND_c_762_n 0.0142237f $X=3.67 $Y=0.38 $X2=0 $Y2=0
cc_347 N_A_297_47#_c_361_n N_VGND_c_762_n 6.07707e-19 $X=4.82 $Y=1.16 $X2=0
+ $Y2=0
cc_348 N_A_297_47#_M1005_s N_VGND_c_763_n 0.00323338f $X=1.485 $Y=0.235 $X2=0
+ $Y2=0
cc_349 N_A_297_47#_M1012_s N_VGND_c_763_n 0.00258107f $X=3.485 $Y=0.235 $X2=0
+ $Y2=0
cc_350 N_A_297_47#_c_356_n N_VGND_c_763_n 0.00938888f $X=4.92 $Y=0.995 $X2=0
+ $Y2=0
cc_351 N_A_297_47#_c_357_n N_VGND_c_763_n 0.00278819f $X=5.39 $Y=0.995 $X2=0
+ $Y2=0
cc_352 N_A_297_47#_c_358_n N_VGND_c_763_n 0.005943f $X=5.86 $Y=0.995 $X2=0 $Y2=0
cc_353 N_A_297_47#_c_359_n N_VGND_c_763_n 0.00278819f $X=6.33 $Y=0.995 $X2=0
+ $Y2=0
cc_354 N_A_297_47#_c_383_n N_VGND_c_763_n 0.0372568f $X=2.6 $Y=0.48 $X2=0 $Y2=0
cc_355 N_A_297_47#_c_372_n N_VGND_c_763_n 0.00941058f $X=3.455 $Y=0.785 $X2=0
+ $Y2=0
cc_356 N_A_297_47#_c_375_n N_VGND_c_763_n 0.013813f $X=3.67 $Y=0.38 $X2=0 $Y2=0
cc_357 N_A_297_47#_c_380_n N_VGND_c_763_n 0.00590183f $X=2.685 $Y=0.48 $X2=0
+ $Y2=0
cc_358 N_A_297_47#_c_383_n A_401_47# 0.00466265f $X=2.6 $Y=0.48 $X2=-0.19
+ $Y2=-0.24
cc_359 N_A_297_47#_c_383_n A_495_47# 0.00313334f $X=2.6 $Y=0.48 $X2=-0.19
+ $Y2=-0.24
cc_360 N_A_297_47#_c_380_n A_495_47# 0.00922746f $X=2.685 $Y=0.48 $X2=-0.19
+ $Y2=-0.24
cc_361 N_A_27_297#_c_512_n N_VPWR_M1002_s 0.00369247f $X=1.115 $Y=1.87 $X2=0.495
+ $Y2=1.41
cc_362 N_A_27_297#_c_515_n N_VPWR_M1015_s 0.0034955f $X=2.055 $Y=1.87 $X2=0.495
+ $Y2=1.985
cc_363 N_A_27_297#_c_516_n N_VPWR_M1011_s 0.00495707f $X=3.115 $Y=1.87 $X2=0.495
+ $Y2=1.985
cc_364 N_A_27_297#_c_512_n N_VPWR_c_574_n 0.0203395f $X=1.115 $Y=1.87 $X2=0.145
+ $Y2=1.105
cc_365 N_A_27_297#_c_522_n N_VPWR_c_574_n 0.0253827f $X=0.26 $Y=1.95 $X2=0.145
+ $Y2=1.105
cc_366 N_A_27_297#_c_524_n N_VPWR_c_574_n 0.0208108f $X=1.2 $Y=1.95 $X2=0.145
+ $Y2=1.105
cc_367 N_A_27_297#_c_515_n N_VPWR_c_575_n 0.0203395f $X=2.055 $Y=1.87 $X2=0.41
+ $Y2=1.16
cc_368 N_A_27_297#_c_524_n N_VPWR_c_575_n 0.0253827f $X=1.2 $Y=1.95 $X2=0.41
+ $Y2=1.16
cc_369 N_A_27_297#_c_525_n N_VPWR_c_575_n 0.0208108f $X=2.14 $Y=1.95 $X2=0.41
+ $Y2=1.16
cc_370 N_A_27_297#_c_516_n N_VPWR_c_576_n 0.0237178f $X=3.115 $Y=1.87 $X2=0.335
+ $Y2=1.16
cc_371 N_A_27_297#_c_525_n N_VPWR_c_576_n 0.0253827f $X=2.14 $Y=1.95 $X2=0.335
+ $Y2=1.16
cc_372 N_A_27_297#_c_530_n N_VPWR_c_577_n 0.010563f $X=4.055 $Y=2.38 $X2=0.335
+ $Y2=1.53
cc_373 N_A_27_297#_c_539_n N_VPWR_c_577_n 0.00949735f $X=4.14 $Y=1.96 $X2=0.335
+ $Y2=1.53
cc_374 N_A_27_297#_c_530_n N_VPWR_c_581_n 0.0534449f $X=4.055 $Y=2.38 $X2=0
+ $Y2=0
cc_375 N_A_27_297#_c_521_n N_VPWR_c_581_n 0.0119545f $X=3.285 $Y=2.38 $X2=0
+ $Y2=0
cc_376 N_A_27_297#_c_522_n N_VPWR_c_585_n 0.0118139f $X=0.26 $Y=1.95 $X2=0 $Y2=0
cc_377 N_A_27_297#_c_524_n N_VPWR_c_586_n 0.0118139f $X=1.2 $Y=1.95 $X2=0 $Y2=0
cc_378 N_A_27_297#_c_525_n N_VPWR_c_587_n 0.0118139f $X=2.14 $Y=1.95 $X2=0 $Y2=0
cc_379 N_A_27_297#_M1002_d N_VPWR_c_573_n 0.00391905f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_380 N_A_27_297#_M1000_d N_VPWR_c_573_n 0.00295369f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_381 N_A_27_297#_M1022_d N_VPWR_c_573_n 0.00295369f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_382 N_A_27_297#_M1007_d N_VPWR_c_573_n 0.00347077f $X=2.995 $Y=1.485 $X2=0
+ $Y2=0
cc_383 N_A_27_297#_M1018_d N_VPWR_c_573_n 0.00356385f $X=3.995 $Y=1.485 $X2=0
+ $Y2=0
cc_384 N_A_27_297#_c_512_n N_VPWR_c_573_n 0.0134894f $X=1.115 $Y=1.87 $X2=0
+ $Y2=0
cc_385 N_A_27_297#_c_515_n N_VPWR_c_573_n 0.0134894f $X=2.055 $Y=1.87 $X2=0
+ $Y2=0
cc_386 N_A_27_297#_c_516_n N_VPWR_c_573_n 0.0178182f $X=3.115 $Y=1.87 $X2=0
+ $Y2=0
cc_387 N_A_27_297#_c_530_n N_VPWR_c_573_n 0.0334226f $X=4.055 $Y=2.38 $X2=0
+ $Y2=0
cc_388 N_A_27_297#_c_521_n N_VPWR_c_573_n 0.006547f $X=3.285 $Y=2.38 $X2=0 $Y2=0
cc_389 N_A_27_297#_c_522_n N_VPWR_c_573_n 0.00646998f $X=0.26 $Y=1.95 $X2=0
+ $Y2=0
cc_390 N_A_27_297#_c_524_n N_VPWR_c_573_n 0.00646998f $X=1.2 $Y=1.95 $X2=0 $Y2=0
cc_391 N_A_27_297#_c_525_n N_VPWR_c_573_n 0.00646998f $X=2.14 $Y=1.95 $X2=0
+ $Y2=0
cc_392 N_VPWR_c_573_n N_X_M1003_d 0.00295281f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_393 N_VPWR_c_573_n N_X_M1013_d 0.00295369f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_394 N_VPWR_M1006_s N_X_c_698_n 0.00437458f $X=5.455 $Y=1.485 $X2=0 $Y2=0
cc_395 N_VPWR_c_578_n N_X_c_698_n 0.0203395f $X=5.6 $Y=2.21 $X2=0 $Y2=0
cc_396 N_VPWR_c_573_n N_X_c_698_n 0.0134894f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_397 N_VPWR_c_577_n N_X_c_702_n 0.0205843f $X=4.66 $Y=2.21 $X2=0 $Y2=0
cc_398 N_VPWR_c_578_n N_X_c_702_n 0.0253827f $X=5.6 $Y=2.21 $X2=0 $Y2=0
cc_399 N_VPWR_c_583_n N_X_c_702_n 0.0118139f $X=5.385 $Y=2.72 $X2=0 $Y2=0
cc_400 N_VPWR_c_573_n N_X_c_702_n 0.0100827f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_401 N_VPWR_c_578_n N_X_c_705_n 0.0208108f $X=5.6 $Y=2.21 $X2=0 $Y2=0
cc_402 N_VPWR_c_580_n N_X_c_705_n 0.0253827f $X=6.54 $Y=2.21 $X2=0 $Y2=0
cc_403 N_VPWR_c_588_n N_X_c_705_n 0.0118139f $X=6.325 $Y=2.72 $X2=0 $Y2=0
cc_404 N_VPWR_c_573_n N_X_c_705_n 0.00646998f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_405 N_VPWR_M1020_s X 0.00810545f $X=6.395 $Y=1.485 $X2=0 $Y2=0
cc_406 N_VPWR_c_579_n X 0.00118135f $X=6.515 $Y=2.635 $X2=0 $Y2=0
cc_407 N_VPWR_c_580_n X 0.0260263f $X=6.54 $Y=2.21 $X2=0 $Y2=0
cc_408 N_VPWR_c_573_n X 0.00881384f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_409 N_VPWR_M1020_s X 0.00488235f $X=6.395 $Y=1.485 $X2=0 $Y2=0
cc_410 X N_VGND_M1008_d 0.00398932f $X=6.585 $Y=0.765 $X2=0 $Y2=0
cc_411 X N_VGND_M1023_d 0.00590716f $X=6.585 $Y=0.765 $X2=0 $Y2=0
cc_412 N_X_c_693_n N_VGND_M1023_d 0.00160749f $X=6.682 $Y=0.825 $X2=0 $Y2=0
cc_413 X N_VGND_M1023_d 9.58474e-19 $X=6.655 $Y=0.85 $X2=0 $Y2=0
cc_414 X N_VGND_c_753_n 0.0214497f $X=6.585 $Y=0.765 $X2=0 $Y2=0
cc_415 N_X_c_693_n N_VGND_c_754_n 0.00146581f $X=6.682 $Y=0.825 $X2=0 $Y2=0
cc_416 X N_VGND_c_755_n 0.0150449f $X=6.585 $Y=0.765 $X2=0 $Y2=0
cc_417 N_X_c_693_n N_VGND_c_755_n 0.0102203f $X=6.682 $Y=0.825 $X2=0 $Y2=0
cc_418 X N_VGND_c_756_n 0.00698859f $X=6.585 $Y=0.765 $X2=0 $Y2=0
cc_419 X N_VGND_c_760_n 0.00810266f $X=6.585 $Y=0.765 $X2=0 $Y2=0
cc_420 N_X_M1004_s N_VGND_c_763_n 0.00384841f $X=4.995 $Y=0.235 $X2=0 $Y2=0
cc_421 N_X_M1010_s N_VGND_c_763_n 0.00384841f $X=5.935 $Y=0.235 $X2=0 $Y2=0
cc_422 X N_VGND_c_763_n 0.0297642f $X=6.585 $Y=0.765 $X2=0 $Y2=0
cc_423 N_X_c_693_n N_VGND_c_763_n 0.00284807f $X=6.682 $Y=0.825 $X2=0 $Y2=0
cc_424 N_VGND_c_763_n A_119_47# 0.00956279f $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24
cc_425 N_VGND_c_763_n A_213_47# 0.00353464f $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24
cc_426 N_VGND_c_763_n A_401_47# 0.00279644f $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24
cc_427 N_VGND_c_763_n A_495_47# 0.00300108f $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24
