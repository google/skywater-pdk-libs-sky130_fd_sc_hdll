* File: sky130_fd_sc_hdll__nand2_16.spice
* Created: Thu Aug 27 19:12:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nand2_16.pex.spice"
.subckt sky130_fd_sc_hdll__nand2_16  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1004 N_A_27_47#_M1004_d N_B_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75014.8 A=0.0975 P=1.6 MULT=1
MM1005 N_A_27_47#_M1005_d N_B_M1005_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75014.3 A=0.0975 P=1.6 MULT=1
MM1014 N_A_27_47#_M1005_d N_B_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.1
+ SB=75013.9 A=0.0975 P=1.6 MULT=1
MM1016 N_A_27_47#_M1016_d N_B_M1016_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.6
+ SB=75013.3 A=0.0975 P=1.6 MULT=1
MM1020 N_A_27_47#_M1016_d N_B_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.1
+ SB=75012.9 A=0.0975 P=1.6 MULT=1
MM1025 N_A_27_47#_M1025_d N_B_M1025_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.6
+ SB=75012.4 A=0.0975 P=1.6 MULT=1
MM1034 N_A_27_47#_M1025_d N_B_M1034_g N_VGND_M1034_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003
+ SB=75012 A=0.0975 P=1.6 MULT=1
MM1035 N_A_27_47#_M1035_d N_B_M1035_g N_VGND_M1034_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.5
+ SB=75011.5 A=0.0975 P=1.6 MULT=1
MM1039 N_A_27_47#_M1035_d N_B_M1039_g N_VGND_M1039_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.9
+ SB=75011 A=0.0975 P=1.6 MULT=1
MM1040 N_A_27_47#_M1040_d N_B_M1040_g N_VGND_M1039_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.5
+ SB=75010.5 A=0.0975 P=1.6 MULT=1
MM1046 N_A_27_47#_M1040_d N_B_M1046_g N_VGND_M1046_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.9
+ SB=75010.1 A=0.0975 P=1.6 MULT=1
MM1053 N_A_27_47#_M1053_d N_B_M1053_g N_VGND_M1046_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75005.4
+ SB=75009.6 A=0.0975 P=1.6 MULT=1
MM1055 N_A_27_47#_M1053_d N_B_M1055_g N_VGND_M1055_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75005.8
+ SB=75009.2 A=0.0975 P=1.6 MULT=1
MM1056 N_A_27_47#_M1056_d N_B_M1056_g N_VGND_M1055_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75006.3
+ SB=75008.6 A=0.0975 P=1.6 MULT=1
MM1057 N_A_27_47#_M1056_d N_B_M1057_g N_VGND_M1057_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75006.8
+ SB=75008.2 A=0.0975 P=1.6 MULT=1
MM1058 N_A_27_47#_M1058_d N_B_M1058_g N_VGND_M1057_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75007.3
+ SB=75007.7 A=0.0975 P=1.6 MULT=1
MM1001 N_Y_M1001_d N_A_M1001_g N_A_27_47#_M1058_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75007.7
+ SB=75007.3 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1001_d N_A_M1006_g N_A_27_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75008.2
+ SB=75006.8 A=0.0975 P=1.6 MULT=1
MM1011 N_Y_M1011_d N_A_M1011_g N_A_27_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75008.6
+ SB=75006.3 A=0.0975 P=1.6 MULT=1
MM1017 N_Y_M1011_d N_A_M1017_g N_A_27_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75009.2
+ SB=75005.8 A=0.0975 P=1.6 MULT=1
MM1018 N_Y_M1018_d N_A_M1018_g N_A_27_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75009.6
+ SB=75005.4 A=0.0975 P=1.6 MULT=1
MM1024 N_Y_M1018_d N_A_M1024_g N_A_27_47#_M1024_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75010.1
+ SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1026 N_Y_M1026_d N_A_M1026_g N_A_27_47#_M1024_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75010.5
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1027 N_Y_M1026_d N_A_M1027_g N_A_27_47#_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75011
+ SB=75004 A=0.0975 P=1.6 MULT=1
MM1030 N_Y_M1030_d N_A_M1030_g N_A_27_47#_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75011.5
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1032 N_Y_M1030_d N_A_M1032_g N_A_27_47#_M1032_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75012
+ SB=75003 A=0.0975 P=1.6 MULT=1
MM1036 N_Y_M1036_d N_A_M1036_g N_A_27_47#_M1032_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75012.4
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1043 N_Y_M1036_d N_A_M1043_g N_A_27_47#_M1043_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75012.9
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1044 N_Y_M1044_d N_A_M1044_g N_A_27_47#_M1043_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75013.3
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1047 N_Y_M1044_d N_A_M1047_g N_A_27_47#_M1047_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75013.9
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1059 N_Y_M1059_d N_A_M1059_g N_A_27_47#_M1047_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75014.3
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1062 N_Y_M1059_d N_A_M1062_g N_A_27_47#_M1062_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.169 PD=1.02 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75014.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_B_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90014.7 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_B_M1002_g N_Y_M1000_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.6
+ SB=90014.3 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1002_d N_B_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.1
+ SB=90013.8 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_B_M1009_g N_Y_M1007_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.6
+ SB=90013.3 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1009_d N_B_M1010_g N_Y_M1010_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.1
+ SB=90012.9 A=0.18 P=2.36 MULT=1
MM1015 N_VPWR_M1015_d N_B_M1015_g N_Y_M1010_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.5
+ SB=90012.4 A=0.18 P=2.36 MULT=1
MM1019 N_VPWR_M1015_d N_B_M1019_g N_Y_M1019_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90011.9 A=0.18 P=2.36 MULT=1
MM1028 N_VPWR_M1028_d N_B_M1028_g N_Y_M1019_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003.5
+ SB=90011.5 A=0.18 P=2.36 MULT=1
MM1033 N_VPWR_M1028_d N_B_M1033_g N_Y_M1033_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003.9
+ SB=90011 A=0.18 P=2.36 MULT=1
MM1037 N_VPWR_M1037_d N_B_M1037_g N_Y_M1033_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90004.4
+ SB=90010.5 A=0.18 P=2.36 MULT=1
MM1042 N_VPWR_M1037_d N_B_M1042_g N_Y_M1042_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90004.9
+ SB=90010 A=0.18 P=2.36 MULT=1
MM1045 N_VPWR_M1045_d N_B_M1045_g N_Y_M1042_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90005.3
+ SB=90009.6 A=0.18 P=2.36 MULT=1
MM1050 N_VPWR_M1045_d N_B_M1050_g N_Y_M1050_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90005.8
+ SB=90009.1 A=0.18 P=2.36 MULT=1
MM1051 N_VPWR_M1051_d N_B_M1051_g N_Y_M1050_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90006.3
+ SB=90008.6 A=0.18 P=2.36 MULT=1
MM1054 N_VPWR_M1051_d N_B_M1054_g N_Y_M1054_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90006.8
+ SB=90008.2 A=0.18 P=2.36 MULT=1
MM1060 N_VPWR_M1060_d N_B_M1060_g N_Y_M1054_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90007.2
+ SB=90007.7 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1060_d N_A_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90007.7
+ SB=90007.2 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90008.2
+ SB=90006.8 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1008_d N_A_M1012_g N_Y_M1012_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90008.6
+ SB=90006.3 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1013_d N_A_M1013_g N_Y_M1012_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90009.1
+ SB=90005.8 A=0.18 P=2.36 MULT=1
MM1021 N_VPWR_M1013_d N_A_M1021_g N_Y_M1021_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90009.6
+ SB=90005.3 A=0.18 P=2.36 MULT=1
MM1022 N_VPWR_M1022_d N_A_M1022_g N_Y_M1021_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90010
+ SB=90004.9 A=0.18 P=2.36 MULT=1
MM1023 N_VPWR_M1022_d N_A_M1023_g N_Y_M1023_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90010.5
+ SB=90004.4 A=0.18 P=2.36 MULT=1
MM1029 N_VPWR_M1029_d N_A_M1029_g N_Y_M1023_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90011
+ SB=90003.9 A=0.18 P=2.36 MULT=1
MM1031 N_VPWR_M1029_d N_A_M1031_g N_Y_M1031_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90011.5
+ SB=90003.5 A=0.18 P=2.36 MULT=1
MM1038 N_VPWR_M1038_d N_A_M1038_g N_Y_M1031_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90011.9
+ SB=90003 A=0.18 P=2.36 MULT=1
MM1041 N_VPWR_M1038_d N_A_M1041_g N_Y_M1041_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90012.4
+ SB=90002.5 A=0.18 P=2.36 MULT=1
MM1048 N_VPWR_M1048_d N_A_M1048_g N_Y_M1041_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90012.9
+ SB=90002.1 A=0.18 P=2.36 MULT=1
MM1049 N_VPWR_M1048_d N_A_M1049_g N_Y_M1049_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90013.3
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1052 N_VPWR_M1052_d N_A_M1052_g N_Y_M1049_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90013.8
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1061 N_VPWR_M1052_d N_A_M1061_g N_Y_M1061_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90014.3
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1063 N_VPWR_M1063_d N_A_M1063_g N_Y_M1061_s VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90014.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX64_noxref VNB VPB NWDIODE A=25.7121 P=35.25
*
.include "sky130_fd_sc_hdll__nand2_16.pxi.spice"
*
.ends
*
*
