* File: sky130_fd_sc_hdll__muxb8to1_2.pxi.spice
* Created: Thu Aug 27 19:12:13 2020
* 
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[0] N_D[0]_M1003_g N_D[0]_M1019_g
+ N_D[0]_M1053_g N_D[0]_M1034_g D[0] N_D[0]_c_429_n N_D[0]_c_430_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[0]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_278_265# N_A_278_265#_M1043_s
+ N_A_278_265#_M1008_s N_A_278_265#_M1006_g N_A_278_265#_c_477_n
+ N_A_278_265#_c_478_n N_A_278_265#_M1013_g N_A_278_265#_c_472_n
+ N_A_278_265#_c_473_n N_A_278_265#_c_480_n N_A_278_265#_c_474_n
+ N_A_278_265#_c_475_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_278_265#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[0] N_S[0]_c_549_n N_S[0]_M1017_g
+ N_S[0]_c_550_n N_S[0]_c_551_n N_S[0]_c_552_n N_S[0]_M1020_g N_S[0]_c_553_n
+ N_S[0]_c_554_n N_S[0]_c_555_n N_S[0]_c_556_n N_S[0]_c_557_n N_S[0]_M1008_g
+ N_S[0]_c_558_n N_S[0]_M1043_g N_S[0]_c_559_n S[0]
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[0]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[1] N_S[1]_c_614_n N_S[1]_M1035_g
+ N_S[1]_c_615_n N_S[1]_M1045_g N_S[1]_c_616_n N_S[1]_c_617_n N_S[1]_c_618_n
+ N_S[1]_c_619_n N_S[1]_c_620_n N_S[1]_M1015_g N_S[1]_c_621_n N_S[1]_c_622_n
+ N_S[1]_M1018_g N_S[1]_c_623_n S[1] PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[1]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_701_47# N_A_701_47#_M1035_d
+ N_A_701_47#_M1045_d N_A_701_47#_M1040_g N_A_701_47#_c_681_n
+ N_A_701_47#_c_676_n N_A_701_47#_M1056_g N_A_701_47#_c_684_n
+ N_A_701_47#_c_677_n N_A_701_47#_c_678_n N_A_701_47#_c_679_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_701_47#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[1] N_D[1]_M1022_g N_D[1]_M1036_g
+ N_D[1]_M1051_g N_D[1]_M1049_g D[1] N_D[1]_c_755_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[1]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[2] N_D[2]_M1000_g N_D[2]_M1057_g
+ N_D[2]_M1063_g N_D[2]_M1060_g D[2] N_D[2]_c_807_n N_D[2]_c_808_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[2]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_1566_265# N_A_1566_265#_M1077_s
+ N_A_1566_265#_M1067_s N_A_1566_265#_M1004_g N_A_1566_265#_c_862_n
+ N_A_1566_265#_c_863_n N_A_1566_265#_M1061_g N_A_1566_265#_c_857_n
+ N_A_1566_265#_c_858_n N_A_1566_265#_c_865_n N_A_1566_265#_c_859_n
+ N_A_1566_265#_c_860_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_1566_265#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[2] N_S[2]_c_935_n N_S[2]_M1058_g
+ N_S[2]_c_936_n N_S[2]_c_937_n N_S[2]_c_938_n N_S[2]_M1076_g N_S[2]_c_939_n
+ N_S[2]_c_940_n N_S[2]_c_941_n N_S[2]_c_942_n N_S[2]_c_943_n N_S[2]_M1067_g
+ N_S[2]_c_944_n N_S[2]_M1077_g N_S[2]_c_945_n S[2]
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[2]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[3] N_S[3]_c_1000_n N_S[3]_M1009_g
+ N_S[3]_c_1001_n N_S[3]_M1023_g N_S[3]_c_1002_n N_S[3]_c_1003_n N_S[3]_c_1004_n
+ N_S[3]_c_1005_n N_S[3]_c_1006_n N_S[3]_M1052_g N_S[3]_c_1007_n N_S[3]_c_1008_n
+ N_S[3]_M1065_g N_S[3]_c_1009_n S[3] PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[3]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_1989_47# N_A_1989_47#_M1009_d
+ N_A_1989_47#_M1023_d N_A_1989_47#_M1005_g N_A_1989_47#_c_1067_n
+ N_A_1989_47#_c_1062_n N_A_1989_47#_M1062_g N_A_1989_47#_c_1070_n
+ N_A_1989_47#_c_1063_n N_A_1989_47#_c_1064_n N_A_1989_47#_c_1065_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_1989_47#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[3] N_D[3]_M1001_g N_D[3]_M1012_g
+ N_D[3]_M1078_g N_D[3]_M1068_g D[3] N_D[3]_c_1141_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[3]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[4] N_D[4]_M1014_g N_D[4]_M1031_g
+ N_D[4]_M1048_g N_D[4]_M1037_g D[4] N_D[4]_c_1193_n N_D[4]_c_1194_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[4]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_2854_265# N_A_2854_265#_M1032_s
+ N_A_2854_265#_M1002_s N_A_2854_265#_M1016_g N_A_2854_265#_c_1248_n
+ N_A_2854_265#_c_1249_n N_A_2854_265#_M1041_g N_A_2854_265#_c_1243_n
+ N_A_2854_265#_c_1244_n N_A_2854_265#_c_1251_n N_A_2854_265#_c_1245_n
+ N_A_2854_265#_c_1246_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_2854_265#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[4] N_S[4]_c_1321_n N_S[4]_M1021_g
+ N_S[4]_c_1322_n N_S[4]_c_1323_n N_S[4]_c_1324_n N_S[4]_M1044_g N_S[4]_c_1325_n
+ N_S[4]_c_1326_n N_S[4]_c_1327_n N_S[4]_c_1328_n N_S[4]_c_1329_n N_S[4]_M1002_g
+ N_S[4]_c_1330_n N_S[4]_M1032_g N_S[4]_c_1331_n S[4]
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[4]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[5] N_S[5]_c_1386_n N_S[5]_M1050_g
+ N_S[5]_c_1387_n N_S[5]_M1028_g N_S[5]_c_1388_n N_S[5]_c_1389_n N_S[5]_c_1390_n
+ N_S[5]_c_1391_n N_S[5]_c_1392_n N_S[5]_M1010_g N_S[5]_c_1393_n N_S[5]_c_1394_n
+ N_S[5]_M1026_g N_S[5]_c_1395_n S[5] PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[5]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_3277_47# N_A_3277_47#_M1050_d
+ N_A_3277_47#_M1028_d N_A_3277_47#_M1024_g N_A_3277_47#_c_1453_n
+ N_A_3277_47#_c_1448_n N_A_3277_47#_M1042_g N_A_3277_47#_c_1456_n
+ N_A_3277_47#_c_1449_n N_A_3277_47#_c_1450_n N_A_3277_47#_c_1451_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_3277_47#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[5] N_D[5]_M1025_g N_D[5]_M1047_g
+ N_D[5]_M1054_g N_D[5]_M1038_g D[5] N_D[5]_c_1527_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[5]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[6] N_D[6]_M1029_g N_D[6]_M1070_g
+ N_D[6]_M1079_g N_D[6]_M1072_g D[6] N_D[6]_c_1579_n N_D[6]_c_1580_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[6]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_4142_265# N_A_4142_265#_M1075_s
+ N_A_4142_265#_M1039_s N_A_4142_265#_M1033_g N_A_4142_265#_c_1634_n
+ N_A_4142_265#_c_1635_n N_A_4142_265#_M1046_g N_A_4142_265#_c_1629_n
+ N_A_4142_265#_c_1630_n N_A_4142_265#_c_1637_n N_A_4142_265#_c_1631_n
+ N_A_4142_265#_c_1632_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_4142_265#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[6] N_S[6]_c_1707_n N_S[6]_M1059_g
+ N_S[6]_c_1708_n N_S[6]_c_1709_n N_S[6]_c_1710_n N_S[6]_M1074_g N_S[6]_c_1711_n
+ N_S[6]_c_1712_n N_S[6]_c_1713_n N_S[6]_c_1714_n N_S[6]_c_1715_n N_S[6]_M1039_g
+ N_S[6]_c_1716_n N_S[6]_M1075_g N_S[6]_c_1717_n S[6]
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[6]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[7] N_S[7]_c_1772_n N_S[7]_M1007_g
+ N_S[7]_c_1773_n N_S[7]_M1066_g N_S[7]_c_1774_n N_S[7]_c_1775_n N_S[7]_c_1776_n
+ N_S[7]_c_1777_n N_S[7]_c_1778_n N_S[7]_M1055_g N_S[7]_c_1779_n N_S[7]_c_1780_n
+ N_S[7]_M1071_g N_S[7]_c_1781_n S[7] PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[7]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_4565_47# N_A_4565_47#_M1007_d
+ N_A_4565_47#_M1066_d N_A_4565_47#_M1064_g N_A_4565_47#_c_1839_n
+ N_A_4565_47#_c_1834_n N_A_4565_47#_M1073_g N_A_4565_47#_c_1842_n
+ N_A_4565_47#_c_1835_n N_A_4565_47#_c_1836_n N_A_4565_47#_c_1837_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_4565_47#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[7] N_D[7]_M1030_g N_D[7]_M1011_g
+ N_D[7]_M1027_g N_D[7]_M1069_g D[7] N_D[7]_c_1912_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[7]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_27_297# N_A_27_297#_M1003_d
+ N_A_27_297#_M1034_d N_A_27_297#_M1013_d N_A_27_297#_c_1953_n
+ N_A_27_297#_c_1959_n N_A_27_297#_c_1963_n N_A_27_297#_c_1967_n
+ N_A_27_297#_c_1975_p N_A_27_297#_c_1954_n N_A_27_297#_c_1955_n
+ N_A_27_297#_c_1956_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%VPWR N_VPWR_M1003_s N_VPWR_M1008_d
+ N_VPWR_M1022_s N_VPWR_M1000_d N_VPWR_M1067_d N_VPWR_M1001_d N_VPWR_M1014_s
+ N_VPWR_M1002_d N_VPWR_M1025_s N_VPWR_M1029_s N_VPWR_M1039_d N_VPWR_M1030_s
+ N_VPWR_c_2001_n N_VPWR_c_2002_n N_VPWR_c_2003_n N_VPWR_c_2004_n
+ N_VPWR_c_2005_n N_VPWR_c_2006_n N_VPWR_c_2007_n N_VPWR_c_2008_n
+ N_VPWR_c_2009_n N_VPWR_c_2010_n N_VPWR_c_2011_n N_VPWR_c_2012_n
+ N_VPWR_c_2041_n N_VPWR_c_2013_n N_VPWR_c_2014_n N_VPWR_c_2077_n
+ N_VPWR_c_2085_n N_VPWR_c_2015_n N_VPWR_c_2016_n N_VPWR_c_2121_n
+ N_VPWR_c_2129_n N_VPWR_c_2017_n N_VPWR_c_2018_n N_VPWR_c_2165_n
+ N_VPWR_c_2173_n N_VPWR_c_2019_n N_VPWR_c_2020_n N_VPWR_c_2209_n VPWR VPWR VPWR
+ VPWR VPWR VPWR VPWR VPWR N_VPWR_c_2022_n N_VPWR_c_2023_n N_VPWR_c_2024_n
+ N_VPWR_c_2025_n N_VPWR_c_2026_n N_VPWR_c_2027_n N_VPWR_c_2028_n
+ N_VPWR_c_2029_n N_VPWR_c_2030_n N_VPWR_c_2031_n N_VPWR_c_2032_n
+ N_VPWR_c_2033_n N_VPWR_c_2034_n N_VPWR_c_2035_n N_VPWR_c_2036_n
+ N_VPWR_c_2037_n N_VPWR_c_2038_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%VPWR
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%Z N_Z_M1017_s N_Z_M1015_s N_Z_M1058_d
+ N_Z_M1052_d N_Z_M1021_d N_Z_M1010_d N_Z_M1059_d N_Z_M1055_d N_Z_M1006_s
+ N_Z_M1040_s N_Z_M1004_d N_Z_M1005_d N_Z_M1016_s N_Z_M1024_s N_Z_M1033_s
+ N_Z_M1064_s N_Z_c_2368_n N_Z_c_2369_n N_Z_c_2370_n N_Z_c_2371_n N_Z_c_2372_n
+ N_Z_c_2373_n N_Z_c_2374_n N_Z_c_2375_n N_Z_c_2384_n N_Z_c_2410_n N_Z_c_2385_n
+ N_Z_c_2441_n N_Z_c_2386_n N_Z_c_2473_n N_Z_c_2387_n N_Z_c_2504_n N_Z_c_2388_n
+ N_Z_c_2536_n N_Z_c_2389_n N_Z_c_2567_n N_Z_c_2390_n N_Z_c_2599_n Z Z Z Z Z Z Z
+ Z N_Z_c_2411_n N_Z_c_2376_n N_Z_c_2442_n N_Z_c_2377_n N_Z_c_2474_n
+ N_Z_c_2378_n N_Z_c_2505_n N_Z_c_2379_n N_Z_c_2537_n N_Z_c_2380_n N_Z_c_2568_n
+ N_Z_c_2381_n N_Z_c_2600_n N_Z_c_2382_n N_Z_c_2630_n N_Z_c_2383_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%Z
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_824_333# N_A_824_333#_M1040_d
+ N_A_824_333#_M1056_d N_A_824_333#_M1049_d N_A_824_333#_c_2850_n
+ N_A_824_333#_c_2858_n N_A_824_333#_c_2860_n N_A_824_333#_c_2861_n
+ N_A_824_333#_c_2864_n N_A_824_333#_c_2862_n N_A_824_333#_c_2851_n
+ N_A_824_333#_c_2852_n N_A_824_333#_c_2853_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_824_333#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_1315_297# N_A_1315_297#_M1000_s
+ N_A_1315_297#_M1060_s N_A_1315_297#_M1061_s N_A_1315_297#_c_2909_n
+ N_A_1315_297#_c_2915_n N_A_1315_297#_c_2919_n N_A_1315_297#_c_2923_n
+ N_A_1315_297#_c_2938_n N_A_1315_297#_c_2910_n N_A_1315_297#_c_2911_n
+ N_A_1315_297#_c_2912_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_1315_297#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_2112_333# N_A_2112_333#_M1005_s
+ N_A_2112_333#_M1062_s N_A_2112_333#_M1068_s N_A_2112_333#_c_2966_n
+ N_A_2112_333#_c_2974_n N_A_2112_333#_c_2976_n N_A_2112_333#_c_2977_n
+ N_A_2112_333#_c_2980_n N_A_2112_333#_c_2978_n N_A_2112_333#_c_2967_n
+ N_A_2112_333#_c_2968_n N_A_2112_333#_c_2969_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_2112_333#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_2603_297# N_A_2603_297#_M1014_d
+ N_A_2603_297#_M1037_d N_A_2603_297#_M1041_d N_A_2603_297#_c_3025_n
+ N_A_2603_297#_c_3031_n N_A_2603_297#_c_3035_n N_A_2603_297#_c_3039_n
+ N_A_2603_297#_c_3054_n N_A_2603_297#_c_3026_n N_A_2603_297#_c_3027_n
+ N_A_2603_297#_c_3028_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_2603_297#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_3400_333# N_A_3400_333#_M1024_d
+ N_A_3400_333#_M1042_d N_A_3400_333#_M1038_d N_A_3400_333#_c_3082_n
+ N_A_3400_333#_c_3090_n N_A_3400_333#_c_3092_n N_A_3400_333#_c_3093_n
+ N_A_3400_333#_c_3096_n N_A_3400_333#_c_3094_n N_A_3400_333#_c_3083_n
+ N_A_3400_333#_c_3084_n N_A_3400_333#_c_3085_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_3400_333#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_3891_297# N_A_3891_297#_M1029_d
+ N_A_3891_297#_M1072_d N_A_3891_297#_M1046_d N_A_3891_297#_c_3141_n
+ N_A_3891_297#_c_3147_n N_A_3891_297#_c_3151_n N_A_3891_297#_c_3155_n
+ N_A_3891_297#_c_3170_n N_A_3891_297#_c_3142_n N_A_3891_297#_c_3143_n
+ N_A_3891_297#_c_3144_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_3891_297#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_4688_333# N_A_4688_333#_M1064_d
+ N_A_4688_333#_M1073_d N_A_4688_333#_M1069_d N_A_4688_333#_c_3198_n
+ N_A_4688_333#_c_3206_n N_A_4688_333#_c_3208_n N_A_4688_333#_c_3209_n
+ N_A_4688_333#_c_3212_n N_A_4688_333#_c_3210_n N_A_4688_333#_c_3199_n
+ N_A_4688_333#_c_3200_n N_A_4688_333#_c_3201_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_4688_333#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_27_47# N_A_27_47#_M1019_d
+ N_A_27_47#_M1053_d N_A_27_47#_M1020_d N_A_27_47#_c_3250_n N_A_27_47#_c_3247_n
+ N_A_27_47#_c_3248_n N_A_27_47#_c_3279_p N_A_27_47#_c_3249_n
+ N_A_27_47#_c_3260_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%VGND N_VGND_M1019_s N_VGND_M1043_d
+ N_VGND_M1036_d N_VGND_M1057_s N_VGND_M1077_d N_VGND_M1012_s N_VGND_M1031_d
+ N_VGND_M1032_d N_VGND_M1047_d N_VGND_M1070_d N_VGND_M1075_d N_VGND_M1011_s
+ N_VGND_c_3289_n N_VGND_c_3290_n N_VGND_c_3291_n N_VGND_c_3292_n
+ N_VGND_c_3293_n N_VGND_c_3294_n N_VGND_c_3295_n N_VGND_c_3296_n
+ N_VGND_c_3297_n N_VGND_c_3298_n N_VGND_c_3299_n N_VGND_c_3300_n
+ N_VGND_c_3301_n N_VGND_c_3302_n N_VGND_c_3303_n N_VGND_c_3304_n
+ N_VGND_c_3305_n N_VGND_c_3306_n N_VGND_c_3307_n N_VGND_c_3308_n
+ N_VGND_c_3309_n N_VGND_c_3310_n N_VGND_c_3311_n N_VGND_c_3312_n
+ N_VGND_c_3313_n VGND VGND VGND VGND VGND VGND VGND VGND N_VGND_c_3315_n
+ N_VGND_c_3316_n N_VGND_c_3317_n N_VGND_c_3318_n N_VGND_c_3319_n
+ N_VGND_c_3320_n N_VGND_c_3321_n N_VGND_c_3322_n N_VGND_c_3323_n
+ N_VGND_c_3324_n N_VGND_c_3325_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%VGND
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_845_69# N_A_845_69#_M1015_d
+ N_A_845_69#_M1018_d N_A_845_69#_M1051_s N_A_845_69#_c_3578_n
+ N_A_845_69#_c_3574_n N_A_845_69#_c_3575_n N_A_845_69#_c_3611_n
+ N_A_845_69#_c_3576_n N_A_845_69#_c_3577_n N_A_845_69#_c_3596_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_845_69#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_1315_47# N_A_1315_47#_M1057_d
+ N_A_1315_47#_M1063_d N_A_1315_47#_M1076_s N_A_1315_47#_c_3625_n
+ N_A_1315_47#_c_3622_n N_A_1315_47#_c_3623_n N_A_1315_47#_c_3660_n
+ N_A_1315_47#_c_3624_n N_A_1315_47#_c_3635_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_1315_47#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_2133_69# N_A_2133_69#_M1052_s
+ N_A_2133_69#_M1065_s N_A_2133_69#_M1078_d N_A_2133_69#_c_3670_n
+ N_A_2133_69#_c_3666_n N_A_2133_69#_c_3667_n N_A_2133_69#_c_3703_n
+ N_A_2133_69#_c_3668_n N_A_2133_69#_c_3669_n N_A_2133_69#_c_3688_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_2133_69#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_2603_47# N_A_2603_47#_M1031_s
+ N_A_2603_47#_M1048_s N_A_2603_47#_M1044_s N_A_2603_47#_c_3717_n
+ N_A_2603_47#_c_3714_n N_A_2603_47#_c_3715_n N_A_2603_47#_c_3752_n
+ N_A_2603_47#_c_3716_n N_A_2603_47#_c_3727_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_2603_47#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_3421_69# N_A_3421_69#_M1010_s
+ N_A_3421_69#_M1026_s N_A_3421_69#_M1054_s N_A_3421_69#_c_3762_n
+ N_A_3421_69#_c_3758_n N_A_3421_69#_c_3759_n N_A_3421_69#_c_3795_n
+ N_A_3421_69#_c_3760_n N_A_3421_69#_c_3761_n N_A_3421_69#_c_3780_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_3421_69#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_3891_47# N_A_3891_47#_M1070_s
+ N_A_3891_47#_M1079_s N_A_3891_47#_M1074_s N_A_3891_47#_c_3809_n
+ N_A_3891_47#_c_3806_n N_A_3891_47#_c_3807_n N_A_3891_47#_c_3844_n
+ N_A_3891_47#_c_3808_n N_A_3891_47#_c_3819_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_3891_47#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_4709_69# N_A_4709_69#_M1055_s
+ N_A_4709_69#_M1071_s N_A_4709_69#_M1027_d N_A_4709_69#_c_3854_n
+ N_A_4709_69#_c_3850_n N_A_4709_69#_c_3851_n N_A_4709_69#_c_3887_n
+ N_A_4709_69#_c_3852_n N_A_4709_69#_c_3853_n N_A_4709_69#_c_3872_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_4709_69#
cc_1 VNB N_D[0]_M1003_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_2 VNB N_D[0]_M1019_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_3 VNB N_D[0]_M1053_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_4 VNB N_D[0]_M1034_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_5 VNB N_D[0]_c_429_n 0.0128835f $X=-0.19 $Y=-0.24 $X2=0.75 $Y2=1.16
cc_6 VNB N_D[0]_c_430_n 0.0571683f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_7 VNB N_A_278_265#_c_472_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_8 VNB N_A_278_265#_c_473_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_278_265#_c_474_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_10 VNB N_A_278_265#_c_475_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_S[0]_c_549_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_12 VNB N_S[0]_c_550_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_S[0]_c_551_n 0.0101495f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.025
cc_14 VNB N_S[0]_c_552_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_15 VNB N_S[0]_c_553_n 0.032124f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_16 VNB N_S[0]_c_554_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_S[0]_c_555_n 0.0222544f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_18 VNB N_S[0]_c_556_n 0.0073997f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_19 VNB N_S[0]_c_557_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_20 VNB N_S[0]_c_558_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_S[0]_c_559_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_22 VNB S[0] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_S[1]_c_614_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_24 VNB N_S[1]_c_615_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_S[1]_c_616_n 0.0296541f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_26 VNB N_S[1]_c_617_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_27 VNB N_S[1]_c_618_n 0.0214653f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_28 VNB N_S[1]_c_619_n 0.0106587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_S[1]_c_620_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_30 VNB N_S[1]_c_621_n 0.0254151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_S[1]_c_622_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_S[1]_c_623_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_33 VNB S[1] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_701_47#_c_676_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_701_47#_c_677_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_701_47#_c_678_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_37 VNB N_A_701_47#_c_679_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_38 VNB N_D[1]_M1022_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_39 VNB N_D[1]_M1036_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_40 VNB N_D[1]_M1051_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_41 VNB N_D[1]_M1049_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_42 VNB D[1] 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_43 VNB N_D[1]_c_755_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_44 VNB N_D[2]_M1000_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_45 VNB N_D[2]_M1057_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_46 VNB N_D[2]_M1063_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_47 VNB N_D[2]_M1060_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_48 VNB N_D[2]_c_807_n 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.75 $Y2=1.16
cc_49 VNB N_D[2]_c_808_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_50 VNB N_A_1566_265#_c_857_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.105
cc_51 VNB N_A_1566_265#_c_858_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_1566_265#_c_859_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_53 VNB N_A_1566_265#_c_860_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_S[2]_c_935_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_55 VNB N_S[2]_c_936_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_S[2]_c_937_n 0.0101495f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.025
cc_57 VNB N_S[2]_c_938_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_58 VNB N_S[2]_c_939_n 0.032124f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_59 VNB N_S[2]_c_940_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_S[2]_c_941_n 0.0222544f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_61 VNB N_S[2]_c_942_n 0.0073997f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_62 VNB N_S[2]_c_943_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_63 VNB N_S[2]_c_944_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_S[2]_c_945_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_65 VNB S[2] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_S[3]_c_1000_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_67 VNB N_S[3]_c_1001_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_S[3]_c_1002_n 0.0296541f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_69 VNB N_S[3]_c_1003_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_70 VNB N_S[3]_c_1004_n 0.0214653f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_71 VNB N_S[3]_c_1005_n 0.0106587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_S[3]_c_1006_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_73 VNB N_S[3]_c_1007_n 0.0254151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_S[3]_c_1008_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_S[3]_c_1009_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_76 VNB S[3] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1989_47#_c_1062_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1989_47#_c_1063_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_1989_47#_c_1064_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_80 VNB N_A_1989_47#_c_1065_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_81 VNB N_D[3]_M1001_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_82 VNB N_D[3]_M1012_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_83 VNB N_D[3]_M1078_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_84 VNB N_D[3]_M1068_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_85 VNB D[3] 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_86 VNB N_D[3]_c_1141_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_87 VNB N_D[4]_M1014_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_88 VNB N_D[4]_M1031_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_89 VNB N_D[4]_M1048_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_90 VNB N_D[4]_M1037_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_91 VNB N_D[4]_c_1193_n 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.75 $Y2=1.16
cc_92 VNB N_D[4]_c_1194_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_93 VNB N_A_2854_265#_c_1243_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.105
cc_94 VNB N_A_2854_265#_c_1244_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_A_2854_265#_c_1245_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_96 VNB N_A_2854_265#_c_1246_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_S[4]_c_1321_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_98 VNB N_S[4]_c_1322_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_S[4]_c_1323_n 0.0101495f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.025
cc_100 VNB N_S[4]_c_1324_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_101 VNB N_S[4]_c_1325_n 0.032124f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_102 VNB N_S[4]_c_1326_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_S[4]_c_1327_n 0.0222544f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_104 VNB N_S[4]_c_1328_n 0.0073997f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_105 VNB N_S[4]_c_1329_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_106 VNB N_S[4]_c_1330_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_S[4]_c_1331_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_108 VNB S[4] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_S[5]_c_1386_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_110 VNB N_S[5]_c_1387_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_S[5]_c_1388_n 0.0296541f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_112 VNB N_S[5]_c_1389_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_113 VNB N_S[5]_c_1390_n 0.0214653f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_114 VNB N_S[5]_c_1391_n 0.0106587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_S[5]_c_1392_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_116 VNB N_S[5]_c_1393_n 0.0254151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_S[5]_c_1394_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_S[5]_c_1395_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_119 VNB S[5] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_A_3277_47#_c_1448_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_A_3277_47#_c_1449_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_A_3277_47#_c_1450_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_123 VNB N_A_3277_47#_c_1451_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_124 VNB N_D[5]_M1025_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_125 VNB N_D[5]_M1047_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_126 VNB N_D[5]_M1054_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_127 VNB N_D[5]_M1038_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_128 VNB D[5] 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_129 VNB N_D[5]_c_1527_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_130 VNB N_D[6]_M1029_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_131 VNB N_D[6]_M1070_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_132 VNB N_D[6]_M1079_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_133 VNB N_D[6]_M1072_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_134 VNB N_D[6]_c_1579_n 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.75 $Y2=1.16
cc_135 VNB N_D[6]_c_1580_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_136 VNB N_A_4142_265#_c_1629_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.105
cc_137 VNB N_A_4142_265#_c_1630_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_138 VNB N_A_4142_265#_c_1631_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94
+ $Y2=1.16
cc_139 VNB N_A_4142_265#_c_1632_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_140 VNB N_S[6]_c_1707_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_141 VNB N_S[6]_c_1708_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_142 VNB N_S[6]_c_1709_n 0.0101495f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.025
cc_143 VNB N_S[6]_c_1710_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_144 VNB N_S[6]_c_1711_n 0.032124f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_145 VNB N_S[6]_c_1712_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_146 VNB N_S[6]_c_1713_n 0.0222544f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_147 VNB N_S[6]_c_1714_n 0.0073997f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_148 VNB N_S[6]_c_1715_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_149 VNB N_S[6]_c_1716_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_150 VNB N_S[6]_c_1717_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_151 VNB S[6] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_152 VNB N_S[7]_c_1772_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_153 VNB N_S[7]_c_1773_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_154 VNB N_S[7]_c_1774_n 0.0296541f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_155 VNB N_S[7]_c_1775_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_156 VNB N_S[7]_c_1776_n 0.0214653f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_157 VNB N_S[7]_c_1777_n 0.0106587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_158 VNB N_S[7]_c_1778_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_159 VNB N_S[7]_c_1779_n 0.0254151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_160 VNB N_S[7]_c_1780_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_161 VNB N_S[7]_c_1781_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_162 VNB S[7] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_163 VNB N_A_4565_47#_c_1834_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_164 VNB N_A_4565_47#_c_1835_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_165 VNB N_A_4565_47#_c_1836_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_166 VNB N_A_4565_47#_c_1837_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_167 VNB N_D[7]_M1030_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_168 VNB N_D[7]_M1011_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_169 VNB N_D[7]_M1027_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_170 VNB N_D[7]_M1069_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_171 VNB D[7] 0.0128835f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_172 VNB N_D[7]_c_1912_n 0.0571683f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_173 VNB VPWR 1.06677f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_174 VNB N_Z_c_2368_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_175 VNB N_Z_c_2369_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_176 VNB N_Z_c_2370_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_177 VNB N_Z_c_2371_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_178 VNB N_Z_c_2372_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_179 VNB N_Z_c_2373_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_180 VNB N_Z_c_2374_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_181 VNB N_Z_c_2375_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_182 VNB N_Z_c_2376_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_183 VNB N_Z_c_2377_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_184 VNB N_Z_c_2378_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_185 VNB N_Z_c_2379_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_186 VNB N_Z_c_2380_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_187 VNB N_Z_c_2381_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_188 VNB N_Z_c_2382_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_189 VNB N_Z_c_2383_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_190 VNB N_A_27_47#_c_3247_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_191 VNB N_A_27_47#_c_3248_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_192 VNB N_A_27_47#_c_3249_n 0.0034739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_193 VNB N_VGND_c_3289_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_194 VNB N_VGND_c_3290_n 0.00516508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_195 VNB N_VGND_c_3291_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_196 VNB N_VGND_c_3292_n 0.0332577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_197 VNB N_VGND_c_3293_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_198 VNB N_VGND_c_3294_n 0.00516508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_199 VNB N_VGND_c_3295_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_200 VNB N_VGND_c_3296_n 0.0332577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_201 VNB N_VGND_c_3297_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_202 VNB N_VGND_c_3298_n 0.00516508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_203 VNB N_VGND_c_3299_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_204 VNB N_VGND_c_3300_n 0.0332577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_205 VNB N_VGND_c_3301_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_206 VNB N_VGND_c_3302_n 0.00516508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_207 VNB N_VGND_c_3303_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_208 VNB N_VGND_c_3304_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_209 VNB N_VGND_c_3305_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_210 VNB N_VGND_c_3306_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_211 VNB N_VGND_c_3307_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_212 VNB N_VGND_c_3308_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_213 VNB N_VGND_c_3309_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_214 VNB N_VGND_c_3310_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_215 VNB N_VGND_c_3311_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_216 VNB N_VGND_c_3312_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_217 VNB N_VGND_c_3313_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_218 VNB VGND 1.17536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_219 VNB N_VGND_c_3315_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_220 VNB N_VGND_c_3316_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_221 VNB N_VGND_c_3317_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_222 VNB N_VGND_c_3318_n 0.0188039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_223 VNB N_VGND_c_3319_n 0.0229085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_224 VNB N_VGND_c_3320_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_225 VNB N_VGND_c_3321_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_226 VNB N_VGND_c_3322_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_227 VNB N_VGND_c_3323_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_228 VNB N_VGND_c_3324_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_229 VNB N_VGND_c_3325_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_230 VNB N_A_845_69#_c_3574_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_231 VNB N_A_845_69#_c_3575_n 0.00109213f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_232 VNB N_A_845_69#_c_3576_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_233 VNB N_A_845_69#_c_3577_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_234 VNB N_A_1315_47#_c_3622_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_235 VNB N_A_1315_47#_c_3623_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_236 VNB N_A_1315_47#_c_3624_n 0.0034739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_237 VNB N_A_2133_69#_c_3666_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_238 VNB N_A_2133_69#_c_3667_n 0.00109213f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_239 VNB N_A_2133_69#_c_3668_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_240 VNB N_A_2133_69#_c_3669_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_241 VNB N_A_2603_47#_c_3714_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_242 VNB N_A_2603_47#_c_3715_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_243 VNB N_A_2603_47#_c_3716_n 0.0034739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_244 VNB N_A_3421_69#_c_3758_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_245 VNB N_A_3421_69#_c_3759_n 0.00109213f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_246 VNB N_A_3421_69#_c_3760_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_247 VNB N_A_3421_69#_c_3761_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_248 VNB N_A_3891_47#_c_3806_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_249 VNB N_A_3891_47#_c_3807_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_250 VNB N_A_3891_47#_c_3808_n 0.0034739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_251 VNB N_A_4709_69#_c_3850_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_252 VNB N_A_4709_69#_c_3851_n 0.00109213f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_253 VNB N_A_4709_69#_c_3852_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_254 VNB N_A_4709_69#_c_3853_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_255 VPB N_D[0]_M1003_g 0.0296461f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_256 VPB N_D[0]_M1034_g 0.0229174f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_257 VPB N_D[0]_c_429_n 0.00632455f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_258 VPB N_A_278_265#_M1006_g 0.0234575f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_259 VPB N_A_278_265#_c_477_n 0.0152663f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_260 VPB N_A_278_265#_c_478_n 0.0114291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_261 VPB N_A_278_265#_M1013_g 0.0267037f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_262 VPB N_A_278_265#_c_480_n 0.0080424f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_263 VPB N_A_278_265#_c_474_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_264 VPB N_A_278_265#_c_475_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_265 VPB N_S[0]_c_557_n 0.0295425f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_266 VPB N_S[1]_c_615_n 0.0295425f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_267 VPB N_A_701_47#_M1040_g 0.0267037f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_268 VPB N_A_701_47#_c_681_n 0.0265655f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_269 VPB N_A_701_47#_c_676_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_270 VPB N_A_701_47#_M1056_g 0.0234575f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_271 VPB N_A_701_47#_c_684_n 0.0080424f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_272 VPB N_A_701_47#_c_679_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_273 VPB N_D[1]_M1022_g 0.0229174f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_274 VPB N_D[1]_M1049_g 0.0296461f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_275 VPB D[1] 0.00525107f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_276 VPB N_D[2]_M1000_g 0.0296461f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_277 VPB N_D[2]_M1060_g 0.0229174f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_278 VPB N_D[2]_c_807_n 0.00525107f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_279 VPB N_A_1566_265#_M1004_g 0.0234575f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_280 VPB N_A_1566_265#_c_862_n 0.0152663f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_281 VPB N_A_1566_265#_c_863_n 0.0112992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_282 VPB N_A_1566_265#_M1061_g 0.0267037f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_283 VPB N_A_1566_265#_c_865_n 0.0080424f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_284 VPB N_A_1566_265#_c_859_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_285 VPB N_A_1566_265#_c_860_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_286 VPB N_S[2]_c_943_n 0.0295425f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_287 VPB N_S[3]_c_1001_n 0.0295425f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_288 VPB N_A_1989_47#_M1005_g 0.0267037f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_289 VPB N_A_1989_47#_c_1067_n 0.0265655f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_290 VPB N_A_1989_47#_c_1062_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_291 VPB N_A_1989_47#_M1062_g 0.0234575f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_292 VPB N_A_1989_47#_c_1070_n 0.0080424f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_293 VPB N_A_1989_47#_c_1065_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_294 VPB N_D[3]_M1001_g 0.0229174f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_295 VPB N_D[3]_M1068_g 0.0296461f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_296 VPB D[3] 0.00525107f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_297 VPB N_D[4]_M1014_g 0.0296461f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_298 VPB N_D[4]_M1037_g 0.0229174f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_299 VPB N_D[4]_c_1193_n 0.00525107f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_300 VPB N_A_2854_265#_M1016_g 0.0234575f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_301 VPB N_A_2854_265#_c_1248_n 0.0152663f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_302 VPB N_A_2854_265#_c_1249_n 0.0112992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_303 VPB N_A_2854_265#_M1041_g 0.0267037f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_304 VPB N_A_2854_265#_c_1251_n 0.0080424f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_305 VPB N_A_2854_265#_c_1245_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_306 VPB N_A_2854_265#_c_1246_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_307 VPB N_S[4]_c_1329_n 0.0295425f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_308 VPB N_S[5]_c_1387_n 0.0295425f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_309 VPB N_A_3277_47#_M1024_g 0.0267037f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_310 VPB N_A_3277_47#_c_1453_n 0.0265655f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_311 VPB N_A_3277_47#_c_1448_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_312 VPB N_A_3277_47#_M1042_g 0.0234575f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_313 VPB N_A_3277_47#_c_1456_n 0.0080424f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_314 VPB N_A_3277_47#_c_1451_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_315 VPB N_D[5]_M1025_g 0.0229174f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_316 VPB N_D[5]_M1038_g 0.0296461f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_317 VPB D[5] 0.00525107f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_318 VPB N_D[6]_M1029_g 0.0296461f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_319 VPB N_D[6]_M1072_g 0.0229174f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_320 VPB N_D[6]_c_1579_n 0.00525107f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_321 VPB N_A_4142_265#_M1033_g 0.0234575f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_322 VPB N_A_4142_265#_c_1634_n 0.0152663f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_323 VPB N_A_4142_265#_c_1635_n 0.0112992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_324 VPB N_A_4142_265#_M1046_g 0.0267037f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_325 VPB N_A_4142_265#_c_1637_n 0.0080424f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_326 VPB N_A_4142_265#_c_1631_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_327 VPB N_A_4142_265#_c_1632_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_328 VPB N_S[6]_c_1715_n 0.0295425f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_329 VPB N_S[7]_c_1773_n 0.0295425f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_330 VPB N_A_4565_47#_M1064_g 0.0267037f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_331 VPB N_A_4565_47#_c_1839_n 0.0266954f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_332 VPB N_A_4565_47#_c_1834_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_333 VPB N_A_4565_47#_M1073_g 0.0234575f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_334 VPB N_A_4565_47#_c_1842_n 0.0080424f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_335 VPB N_A_4565_47#_c_1837_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_336 VPB N_D[7]_M1030_g 0.0229174f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_337 VPB N_D[7]_M1069_g 0.0296461f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_338 VPB D[7] 0.00632455f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_339 VPB N_A_27_297#_c_1953_n 0.0075508f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_340 VPB N_A_27_297#_c_1954_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_341 VPB N_A_27_297#_c_1955_n 0.0101553f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_342 VPB N_A_27_297#_c_1956_n 0.0207852f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_343 VPB N_VPWR_c_2001_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_344 VPB N_VPWR_c_2002_n 0.0147403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_345 VPB N_VPWR_c_2003_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_346 VPB N_VPWR_c_2004_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_347 VPB N_VPWR_c_2005_n 0.0147403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_348 VPB N_VPWR_c_2006_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_349 VPB N_VPWR_c_2007_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_350 VPB N_VPWR_c_2008_n 0.0147403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_351 VPB N_VPWR_c_2009_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_352 VPB N_VPWR_c_2010_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_353 VPB N_VPWR_c_2011_n 0.0147403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_354 VPB N_VPWR_c_2012_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_355 VPB N_VPWR_c_2013_n 0.0531719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_356 VPB N_VPWR_c_2014_n 0.00631862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_357 VPB N_VPWR_c_2015_n 0.0531719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_358 VPB N_VPWR_c_2016_n 0.00631862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_359 VPB N_VPWR_c_2017_n 0.0531719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_360 VPB N_VPWR_c_2018_n 0.00631862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_361 VPB N_VPWR_c_2019_n 0.0531719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_362 VPB N_VPWR_c_2020_n 0.00631862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_363 VPB VPWR 0.0875596f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_364 VPB N_VPWR_c_2022_n 0.0177253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_365 VPB N_VPWR_c_2023_n 0.0531719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_366 VPB N_VPWR_c_2024_n 0.0311005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_367 VPB N_VPWR_c_2025_n 0.0531719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_368 VPB N_VPWR_c_2026_n 0.0311005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_369 VPB N_VPWR_c_2027_n 0.0531719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_370 VPB N_VPWR_c_2028_n 0.0311005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_371 VPB N_VPWR_c_2029_n 0.0531719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_372 VPB N_VPWR_c_2030_n 0.0177253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_373 VPB N_VPWR_c_2031_n 0.00455763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_374 VPB N_VPWR_c_2032_n 0.00455763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_375 VPB N_VPWR_c_2033_n 0.00455763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_376 VPB N_VPWR_c_2034_n 0.00455763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_377 VPB N_VPWR_c_2035_n 0.00455763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_378 VPB N_VPWR_c_2036_n 0.00455763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_379 VPB N_VPWR_c_2037_n 0.00455763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_380 VPB N_VPWR_c_2038_n 0.00455763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_381 VPB N_Z_c_2384_n 0.0098056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_382 VPB N_Z_c_2385_n 0.00920862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_383 VPB N_Z_c_2386_n 0.0098056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_384 VPB N_Z_c_2387_n 0.00920862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_385 VPB N_Z_c_2388_n 0.0098056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_386 VPB N_Z_c_2389_n 0.00920862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_387 VPB N_Z_c_2390_n 0.0098056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_388 VPB N_Z_c_2376_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_389 VPB N_Z_c_2377_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_390 VPB N_Z_c_2378_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_391 VPB N_Z_c_2379_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_392 VPB N_Z_c_2380_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_393 VPB N_Z_c_2381_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_394 VPB N_Z_c_2382_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_395 VPB N_Z_c_2383_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_396 VPB N_A_824_333#_c_2850_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_397 VPB N_A_824_333#_c_2851_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_398 VPB N_A_824_333#_c_2852_n 0.00256593f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_399 VPB N_A_824_333#_c_2853_n 0.00433305f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_400 VPB N_A_1315_297#_c_2909_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=0.56
cc_401 VPB N_A_1315_297#_c_2910_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_402 VPB N_A_1315_297#_c_2911_n 0.00256593f $X=-0.19 $Y=1.305 $X2=0.75
+ $Y2=1.16
cc_403 VPB N_A_1315_297#_c_2912_n 0.00433305f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=1.16
cc_404 VPB N_A_2112_333#_c_2966_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_405 VPB N_A_2112_333#_c_2967_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_406 VPB N_A_2112_333#_c_2968_n 0.00256593f $X=-0.19 $Y=1.305 $X2=0.75
+ $Y2=1.16
cc_407 VPB N_A_2112_333#_c_2969_n 0.00433305f $X=-0.19 $Y=1.305 $X2=0.75
+ $Y2=1.16
cc_408 VPB N_A_2603_297#_c_3025_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=0.56
cc_409 VPB N_A_2603_297#_c_3026_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_410 VPB N_A_2603_297#_c_3027_n 0.00256593f $X=-0.19 $Y=1.305 $X2=0.75
+ $Y2=1.16
cc_411 VPB N_A_2603_297#_c_3028_n 0.00433305f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=1.16
cc_412 VPB N_A_3400_333#_c_3082_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_413 VPB N_A_3400_333#_c_3083_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_414 VPB N_A_3400_333#_c_3084_n 0.00256593f $X=-0.19 $Y=1.305 $X2=0.75
+ $Y2=1.16
cc_415 VPB N_A_3400_333#_c_3085_n 0.00433305f $X=-0.19 $Y=1.305 $X2=0.75
+ $Y2=1.16
cc_416 VPB N_A_3891_297#_c_3141_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=0.56
cc_417 VPB N_A_3891_297#_c_3142_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_418 VPB N_A_3891_297#_c_3143_n 0.00256593f $X=-0.19 $Y=1.305 $X2=0.75
+ $Y2=1.16
cc_419 VPB N_A_3891_297#_c_3144_n 0.00433305f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=1.16
cc_420 VPB N_A_4688_333#_c_3198_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_421 VPB N_A_4688_333#_c_3199_n 0.0075508f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_422 VPB N_A_4688_333#_c_3200_n 0.0101553f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_423 VPB N_A_4688_333#_c_3201_n 0.0207852f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_424 N_D[0]_M1034_g N_A_278_265#_M1006_g 0.0232231f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_425 N_D[0]_M1034_g N_A_278_265#_c_478_n 0.00671996f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_426 N_D[0]_M1053_g N_S[0]_c_551_n 0.0165585f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_427 N_D[0]_c_429_n N_A_27_297#_c_1953_n 0.0235932f $X=0.75 $Y=1.16 $X2=0
+ $Y2=0
cc_428 N_D[0]_c_430_n N_A_27_297#_c_1953_n 9.6385e-19 $X=0.965 $Y=1.16 $X2=0
+ $Y2=0
cc_429 N_D[0]_M1003_g N_A_27_297#_c_1959_n 0.0142998f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_430 N_D[0]_M1034_g N_A_27_297#_c_1959_n 0.0174487f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_431 N_D[0]_c_429_n N_A_27_297#_c_1959_n 0.0339353f $X=0.75 $Y=1.16 $X2=0
+ $Y2=0
cc_432 N_D[0]_c_430_n N_A_27_297#_c_1959_n 7.13708e-19 $X=0.965 $Y=1.16 $X2=0
+ $Y2=0
cc_433 N_D[0]_M1034_g N_A_27_297#_c_1963_n 0.00557487f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_434 N_D[0]_M1003_g N_A_27_297#_c_1955_n 0.00329008f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_435 N_D[0]_M1003_g N_VPWR_c_2001_n 0.0031734f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_436 N_D[0]_M1034_g N_VPWR_c_2001_n 0.00919666f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_437 N_D[0]_M1003_g N_VPWR_c_2041_n 0.00363183f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_438 N_D[0]_M1034_g N_VPWR_c_2041_n 0.00343746f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_439 N_D[0]_M1034_g N_VPWR_c_2013_n 0.00622633f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_440 N_D[0]_M1003_g VPWR 0.0120316f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_441 N_D[0]_M1034_g VPWR 0.0105515f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_442 N_D[0]_M1003_g N_VPWR_c_2022_n 0.00652917f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_443 N_D[0]_M1053_g N_Z_c_2376_n 8.13311e-19 $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_444 N_D[0]_M1034_g N_Z_c_2376_n 0.00112534f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_445 N_D[0]_c_429_n N_Z_c_2376_n 0.00742792f $X=0.75 $Y=1.16 $X2=0 $Y2=0
cc_446 N_D[0]_c_430_n N_Z_c_2376_n 0.00583073f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_447 N_D[0]_M1019_g N_A_27_47#_c_3250_n 0.00633603f $X=0.52 $Y=0.56 $X2=0
+ $Y2=0
cc_448 N_D[0]_M1053_g N_A_27_47#_c_3250_n 5.29024e-19 $X=0.94 $Y=0.56 $X2=0
+ $Y2=0
cc_449 N_D[0]_M1019_g N_A_27_47#_c_3247_n 0.0084485f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_450 N_D[0]_M1053_g N_A_27_47#_c_3247_n 0.0125955f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_451 N_D[0]_c_429_n N_A_27_47#_c_3247_n 0.0274027f $X=0.75 $Y=1.16 $X2=0 $Y2=0
cc_452 N_D[0]_c_430_n N_A_27_47#_c_3247_n 0.00321151f $X=0.965 $Y=1.16 $X2=0
+ $Y2=0
cc_453 N_D[0]_M1019_g N_A_27_47#_c_3248_n 8.68782e-19 $X=0.52 $Y=0.56 $X2=0
+ $Y2=0
cc_454 N_D[0]_c_429_n N_A_27_47#_c_3248_n 0.024456f $X=0.75 $Y=1.16 $X2=0 $Y2=0
cc_455 N_D[0]_c_430_n N_A_27_47#_c_3248_n 0.00464565f $X=0.965 $Y=1.16 $X2=0
+ $Y2=0
cc_456 N_D[0]_M1019_g N_VGND_c_3289_n 0.0030929f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_457 N_D[0]_M1053_g N_VGND_c_3289_n 0.00300333f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_458 N_D[0]_M1053_g N_VGND_c_3304_n 0.00436487f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_459 N_D[0]_M1019_g VGND 0.00697949f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_460 N_D[0]_M1053_g VGND 0.00600262f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_461 N_D[0]_M1019_g N_VGND_c_3319_n 0.00430643f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_462 N_A_278_265#_c_478_n N_S[0]_c_549_n 0.00779314f $X=1.58 $Y=1.4 $X2=-0.19
+ $Y2=-0.24
cc_463 N_A_278_265#_c_477_n N_S[0]_c_552_n 0.00810157f $X=1.87 $Y=1.4 $X2=0
+ $Y2=0
cc_464 N_A_278_265#_c_473_n N_S[0]_c_552_n 7.04048e-19 $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_465 N_A_278_265#_c_472_n N_S[0]_c_554_n 0.0100587f $X=2.43 $Y=0.755 $X2=0
+ $Y2=0
cc_466 N_A_278_265#_c_473_n N_S[0]_c_554_n 0.00267287f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_467 N_A_278_265#_c_472_n N_S[0]_c_555_n 0.0105766f $X=2.43 $Y=0.755 $X2=0
+ $Y2=0
cc_468 N_A_278_265#_c_473_n N_S[0]_c_555_n 0.0090765f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_469 N_A_278_265#_c_474_n N_S[0]_c_555_n 0.00742826f $X=2.715 $Y=1.63 $X2=0
+ $Y2=0
cc_470 N_A_278_265#_c_473_n N_S[0]_c_556_n 0.00445422f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_471 N_A_278_265#_c_474_n N_S[0]_c_556_n 4.25171e-19 $X=2.715 $Y=1.63 $X2=0
+ $Y2=0
cc_472 N_A_278_265#_c_475_n N_S[0]_c_556_n 0.00920672f $X=1.96 $Y=1.34 $X2=0
+ $Y2=0
cc_473 N_A_278_265#_c_473_n N_S[0]_c_557_n 0.00205356f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_474 N_A_278_265#_c_480_n N_S[0]_c_557_n 0.00862444f $X=2.715 $Y=2.31 $X2=0
+ $Y2=0
cc_475 N_A_278_265#_c_474_n N_S[0]_c_557_n 0.00828481f $X=2.715 $Y=1.63 $X2=0
+ $Y2=0
cc_476 N_A_278_265#_c_475_n N_S[0]_c_557_n 0.00692516f $X=1.96 $Y=1.34 $X2=0
+ $Y2=0
cc_477 N_A_278_265#_c_473_n N_S[0]_c_558_n 0.00149517f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_478 N_A_278_265#_c_472_n S[0] 0.0061421f $X=2.43 $Y=0.755 $X2=0 $Y2=0
cc_479 N_A_278_265#_c_473_n S[0] 0.0101733f $X=2.43 $Y=1.205 $X2=0 $Y2=0
cc_480 N_A_278_265#_c_474_n S[0] 0.0127184f $X=2.715 $Y=1.63 $X2=0 $Y2=0
cc_481 N_A_278_265#_c_475_n S[0] 3.07062e-19 $X=1.96 $Y=1.34 $X2=0 $Y2=0
cc_482 N_A_278_265#_M1006_g N_A_27_297#_c_1959_n 0.00176121f $X=1.49 $Y=2.075
+ $X2=0 $Y2=0
cc_483 N_A_278_265#_M1006_g N_A_27_297#_c_1963_n 0.00736707f $X=1.49 $Y=2.075
+ $X2=0 $Y2=0
cc_484 N_A_278_265#_M1006_g N_A_27_297#_c_1967_n 0.0128147f $X=1.49 $Y=2.075
+ $X2=0 $Y2=0
cc_485 N_A_278_265#_M1013_g N_A_27_297#_c_1967_n 0.00971609f $X=1.96 $Y=2.075
+ $X2=0 $Y2=0
cc_486 N_A_278_265#_c_480_n N_A_27_297#_c_1967_n 0.010563f $X=2.715 $Y=2.31
+ $X2=0 $Y2=0
cc_487 N_A_278_265#_M1013_g N_A_27_297#_c_1954_n 0.00745341f $X=1.96 $Y=2.075
+ $X2=0 $Y2=0
cc_488 N_A_278_265#_c_480_n N_A_27_297#_c_1954_n 0.0347621f $X=2.715 $Y=2.31
+ $X2=0 $Y2=0
cc_489 N_A_278_265#_c_474_n N_A_27_297#_c_1954_n 0.0132748f $X=2.715 $Y=1.63
+ $X2=0 $Y2=0
cc_490 N_A_278_265#_c_475_n N_A_27_297#_c_1954_n 0.00133381f $X=1.96 $Y=1.34
+ $X2=0 $Y2=0
cc_491 N_A_278_265#_M1006_g N_VPWR_c_2001_n 0.00107974f $X=1.49 $Y=2.075 $X2=0
+ $Y2=0
cc_492 N_A_278_265#_c_480_n N_VPWR_c_2002_n 0.0321301f $X=2.715 $Y=2.31 $X2=0
+ $Y2=0
cc_493 N_A_278_265#_c_474_n N_VPWR_c_2002_n 0.00732952f $X=2.715 $Y=1.63 $X2=0
+ $Y2=0
cc_494 N_A_278_265#_M1006_g N_VPWR_c_2013_n 0.00429453f $X=1.49 $Y=2.075 $X2=0
+ $Y2=0
cc_495 N_A_278_265#_M1013_g N_VPWR_c_2013_n 0.00429453f $X=1.96 $Y=2.075 $X2=0
+ $Y2=0
cc_496 N_A_278_265#_c_480_n N_VPWR_c_2013_n 0.0210596f $X=2.715 $Y=2.31 $X2=0
+ $Y2=0
cc_497 N_A_278_265#_M1008_s VPWR 0.00179197f $X=2.59 $Y=1.485 $X2=0 $Y2=0
cc_498 N_A_278_265#_M1006_g VPWR 0.00617598f $X=1.49 $Y=2.075 $X2=0 $Y2=0
cc_499 N_A_278_265#_M1013_g VPWR 0.00728421f $X=1.96 $Y=2.075 $X2=0 $Y2=0
cc_500 N_A_278_265#_c_480_n VPWR 0.00594162f $X=2.715 $Y=2.31 $X2=0 $Y2=0
cc_501 N_A_278_265#_c_477_n N_Z_c_2368_n 0.00168443f $X=1.87 $Y=1.4 $X2=0 $Y2=0
cc_502 N_A_278_265#_c_478_n N_Z_c_2368_n 0.00180308f $X=1.58 $Y=1.4 $X2=0 $Y2=0
cc_503 N_A_278_265#_c_473_n N_Z_c_2368_n 0.0033343f $X=2.43 $Y=1.205 $X2=0 $Y2=0
cc_504 N_A_278_265#_M1013_g N_Z_c_2384_n 0.00753886f $X=1.96 $Y=2.075 $X2=0
+ $Y2=0
cc_505 N_A_278_265#_c_480_n N_Z_c_2384_n 0.0308332f $X=2.715 $Y=2.31 $X2=0 $Y2=0
cc_506 N_A_278_265#_c_474_n N_Z_c_2384_n 0.0132841f $X=2.715 $Y=1.63 $X2=0 $Y2=0
cc_507 N_A_278_265#_c_475_n N_Z_c_2384_n 9.57301e-19 $X=1.96 $Y=1.34 $X2=0 $Y2=0
cc_508 N_A_278_265#_M1006_g N_Z_c_2410_n 0.00635853f $X=1.49 $Y=2.075 $X2=0
+ $Y2=0
cc_509 N_A_278_265#_M1006_g N_Z_c_2411_n 0.0105371f $X=1.49 $Y=2.075 $X2=0 $Y2=0
cc_510 N_A_278_265#_c_477_n N_Z_c_2411_n 8.37785e-19 $X=1.87 $Y=1.4 $X2=0 $Y2=0
cc_511 N_A_278_265#_M1013_g N_Z_c_2411_n 0.00635536f $X=1.96 $Y=2.075 $X2=0
+ $Y2=0
cc_512 N_A_278_265#_M1006_g N_Z_c_2376_n 0.00268051f $X=1.49 $Y=2.075 $X2=0
+ $Y2=0
cc_513 N_A_278_265#_c_477_n N_Z_c_2376_n 0.0140509f $X=1.87 $Y=1.4 $X2=0 $Y2=0
cc_514 N_A_278_265#_M1013_g N_Z_c_2376_n 0.00476154f $X=1.96 $Y=2.075 $X2=0
+ $Y2=0
cc_515 N_A_278_265#_c_473_n N_Z_c_2376_n 0.00967956f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_516 N_A_278_265#_c_474_n N_Z_c_2376_n 0.0117695f $X=2.715 $Y=1.63 $X2=0 $Y2=0
cc_517 N_A_278_265#_c_475_n N_Z_c_2376_n 7.26438e-19 $X=1.96 $Y=1.34 $X2=0 $Y2=0
cc_518 N_A_278_265#_c_472_n N_A_27_47#_c_3249_n 0.00358194f $X=2.43 $Y=0.755
+ $X2=0 $Y2=0
cc_519 N_A_278_265#_c_472_n N_A_27_47#_c_3260_n 0.0185512f $X=2.43 $Y=0.755
+ $X2=0 $Y2=0
cc_520 N_A_278_265#_c_473_n N_A_27_47#_c_3260_n 0.00101918f $X=2.43 $Y=1.205
+ $X2=0 $Y2=0
cc_521 N_A_278_265#_c_474_n N_A_27_47#_c_3260_n 0.00285813f $X=2.715 $Y=1.63
+ $X2=0 $Y2=0
cc_522 N_A_278_265#_c_475_n N_A_27_47#_c_3260_n 0.00308807f $X=1.96 $Y=1.34
+ $X2=0 $Y2=0
cc_523 N_A_278_265#_c_472_n N_VGND_c_3304_n 0.0173492f $X=2.43 $Y=0.755 $X2=0
+ $Y2=0
cc_524 N_A_278_265#_M1043_s VGND 0.00250855f $X=2.675 $Y=0.235 $X2=0 $Y2=0
cc_525 N_A_278_265#_c_472_n VGND 0.0186564f $X=2.43 $Y=0.755 $X2=0 $Y2=0
cc_526 N_S[0]_c_558_n N_S[1]_c_614_n 0.0133556f $X=3.01 $Y=0.845 $X2=-0.19
+ $Y2=-0.24
cc_527 N_S[0]_c_557_n N_S[1]_c_615_n 0.0418422f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_528 S[0] N_S[1]_c_615_n 8.74983e-19 $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_529 N_S[0]_c_557_n S[1] 8.74983e-19 $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_530 S[0] S[1] 0.0208489f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_531 N_S[0]_c_557_n N_VPWR_c_2002_n 0.00456891f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_532 S[0] N_VPWR_c_2002_n 0.00569857f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_533 N_S[0]_c_557_n N_VPWR_c_2013_n 0.00673617f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_534 N_S[0]_c_557_n VPWR 0.00852379f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_535 N_S[0]_c_549_n N_Z_c_2368_n 0.00413022f $X=1.46 $Y=0.255 $X2=0 $Y2=0
cc_536 N_S[0]_c_552_n N_Z_c_2368_n 0.00495983f $X=1.88 $Y=0.255 $X2=0 $Y2=0
cc_537 N_S[0]_c_554_n N_Z_c_2368_n 4.25992e-19 $X=2.365 $Y=0.845 $X2=0 $Y2=0
cc_538 N_S[0]_c_557_n N_Z_c_2384_n 0.00513674f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_539 S[0] N_Z_c_2384_n 0.00545567f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_540 N_S[0]_c_549_n N_Z_c_2376_n 0.00199103f $X=1.46 $Y=0.255 $X2=0 $Y2=0
cc_541 N_S[0]_c_552_n N_Z_c_2376_n 0.00133607f $X=1.88 $Y=0.255 $X2=0 $Y2=0
cc_542 N_S[0]_c_549_n N_A_27_47#_c_3247_n 0.00139422f $X=1.46 $Y=0.255 $X2=0
+ $Y2=0
cc_543 N_S[0]_c_549_n N_A_27_47#_c_3249_n 0.0132844f $X=1.46 $Y=0.255 $X2=0
+ $Y2=0
cc_544 N_S[0]_c_550_n N_A_27_47#_c_3249_n 0.00211351f $X=1.805 $Y=0.18 $X2=0
+ $Y2=0
cc_545 N_S[0]_c_552_n N_A_27_47#_c_3249_n 0.0126455f $X=1.88 $Y=0.255 $X2=0
+ $Y2=0
cc_546 N_S[0]_c_553_n N_A_27_47#_c_3249_n 0.00436105f $X=2.29 $Y=0.18 $X2=0
+ $Y2=0
cc_547 N_S[0]_c_554_n N_A_27_47#_c_3249_n 0.00349455f $X=2.365 $Y=0.845 $X2=0
+ $Y2=0
cc_548 N_S[0]_c_554_n N_A_27_47#_c_3260_n 0.00295202f $X=2.365 $Y=0.845 $X2=0
+ $Y2=0
cc_549 N_S[0]_c_558_n N_VGND_c_3290_n 0.00330937f $X=3.01 $Y=0.845 $X2=0 $Y2=0
cc_550 N_S[0]_c_551_n N_VGND_c_3304_n 0.0271255f $X=1.535 $Y=0.18 $X2=0 $Y2=0
cc_551 N_S[0]_c_558_n N_VGND_c_3304_n 0.00585385f $X=3.01 $Y=0.845 $X2=0 $Y2=0
cc_552 N_S[0]_c_550_n VGND 0.00642387f $X=1.805 $Y=0.18 $X2=0 $Y2=0
cc_553 N_S[0]_c_551_n VGND 0.00474746f $X=1.535 $Y=0.18 $X2=0 $Y2=0
cc_554 N_S[0]_c_553_n VGND 0.0193094f $X=2.29 $Y=0.18 $X2=0 $Y2=0
cc_555 N_S[0]_c_558_n VGND 0.0111218f $X=3.01 $Y=0.845 $X2=0 $Y2=0
cc_556 N_S[0]_c_559_n VGND 0.00366655f $X=1.88 $Y=0.18 $X2=0 $Y2=0
cc_557 N_S[1]_c_622_n N_A_701_47#_c_681_n 0.00779314f $X=4.98 $Y=0.255 $X2=0
+ $Y2=0
cc_558 N_S[1]_c_615_n N_A_701_47#_c_676_n 0.00692516f $X=3.49 $Y=1.41 $X2=0
+ $Y2=0
cc_559 N_S[1]_c_616_n N_A_701_47#_c_676_n 0.00920672f $X=4 $Y=0.92 $X2=0 $Y2=0
cc_560 N_S[1]_c_620_n N_A_701_47#_c_676_n 0.00810157f $X=4.56 $Y=0.255 $X2=0
+ $Y2=0
cc_561 S[1] N_A_701_47#_c_676_n 3.07062e-19 $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_562 N_S[1]_c_615_n N_A_701_47#_c_684_n 0.00862444f $X=3.49 $Y=1.41 $X2=0
+ $Y2=0
cc_563 N_S[1]_c_614_n N_A_701_47#_c_677_n 0.00149517f $X=3.43 $Y=0.845 $X2=0
+ $Y2=0
cc_564 N_S[1]_c_615_n N_A_701_47#_c_677_n 0.00205356f $X=3.49 $Y=1.41 $X2=0
+ $Y2=0
cc_565 N_S[1]_c_616_n N_A_701_47#_c_677_n 0.0135307f $X=4 $Y=0.92 $X2=0 $Y2=0
cc_566 N_S[1]_c_617_n N_A_701_47#_c_677_n 0.00267287f $X=4.075 $Y=0.845 $X2=0
+ $Y2=0
cc_567 N_S[1]_c_620_n N_A_701_47#_c_677_n 7.04048e-19 $X=4.56 $Y=0.255 $X2=0
+ $Y2=0
cc_568 S[1] N_A_701_47#_c_677_n 0.0101733f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_569 N_S[1]_c_615_n N_A_701_47#_c_678_n 0.0105766f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_570 N_S[1]_c_617_n N_A_701_47#_c_678_n 0.0100587f $X=4.075 $Y=0.845 $X2=0
+ $Y2=0
cc_571 S[1] N_A_701_47#_c_678_n 0.0061421f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_572 N_S[1]_c_615_n N_A_701_47#_c_679_n 0.00828481f $X=3.49 $Y=1.41 $X2=0
+ $Y2=0
cc_573 N_S[1]_c_616_n N_A_701_47#_c_679_n 0.00785343f $X=4 $Y=0.92 $X2=0 $Y2=0
cc_574 S[1] N_A_701_47#_c_679_n 0.0127184f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_575 N_S[1]_c_621_n N_D[1]_M1036_g 0.0165585f $X=4.905 $Y=0.18 $X2=0 $Y2=0
cc_576 N_S[1]_c_615_n N_VPWR_c_2002_n 0.00456891f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_577 S[1] N_VPWR_c_2002_n 0.00569857f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_578 N_S[1]_c_615_n VPWR 0.00852379f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_579 N_S[1]_c_615_n N_VPWR_c_2023_n 0.00673617f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_580 N_S[1]_c_617_n N_Z_c_2369_n 4.25992e-19 $X=4.075 $Y=0.845 $X2=0 $Y2=0
cc_581 N_S[1]_c_620_n N_Z_c_2369_n 0.00495983f $X=4.56 $Y=0.255 $X2=0 $Y2=0
cc_582 N_S[1]_c_622_n N_Z_c_2369_n 0.00413022f $X=4.98 $Y=0.255 $X2=0 $Y2=0
cc_583 N_S[1]_c_615_n N_Z_c_2384_n 0.00513674f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_584 S[1] N_Z_c_2384_n 0.00545567f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_585 N_S[1]_c_620_n N_Z_c_2377_n 0.00133607f $X=4.56 $Y=0.255 $X2=0 $Y2=0
cc_586 N_S[1]_c_622_n N_Z_c_2377_n 0.00199103f $X=4.98 $Y=0.255 $X2=0 $Y2=0
cc_587 N_S[1]_c_614_n N_VGND_c_3290_n 0.00330937f $X=3.43 $Y=0.845 $X2=0 $Y2=0
cc_588 N_S[1]_c_614_n VGND 0.0111218f $X=3.43 $Y=0.845 $X2=0 $Y2=0
cc_589 N_S[1]_c_618_n VGND 0.0119932f $X=4.485 $Y=0.18 $X2=0 $Y2=0
cc_590 N_S[1]_c_619_n VGND 0.00731624f $X=4.15 $Y=0.18 $X2=0 $Y2=0
cc_591 N_S[1]_c_621_n VGND 0.0111713f $X=4.905 $Y=0.18 $X2=0 $Y2=0
cc_592 N_S[1]_c_623_n VGND 0.00366655f $X=4.56 $Y=0.18 $X2=0 $Y2=0
cc_593 N_S[1]_c_614_n N_VGND_c_3315_n 0.00585385f $X=3.43 $Y=0.845 $X2=0 $Y2=0
cc_594 N_S[1]_c_619_n N_VGND_c_3315_n 0.0271255f $X=4.15 $Y=0.18 $X2=0 $Y2=0
cc_595 N_S[1]_c_617_n N_A_845_69#_c_3578_n 0.00295202f $X=4.075 $Y=0.845 $X2=0
+ $Y2=0
cc_596 N_S[1]_c_620_n N_A_845_69#_c_3574_n 0.0126455f $X=4.56 $Y=0.255 $X2=0
+ $Y2=0
cc_597 N_S[1]_c_621_n N_A_845_69#_c_3574_n 0.00211351f $X=4.905 $Y=0.18 $X2=0
+ $Y2=0
cc_598 N_S[1]_c_622_n N_A_845_69#_c_3574_n 0.0132844f $X=4.98 $Y=0.255 $X2=0
+ $Y2=0
cc_599 N_S[1]_c_617_n N_A_845_69#_c_3575_n 0.00349455f $X=4.075 $Y=0.845 $X2=0
+ $Y2=0
cc_600 N_S[1]_c_618_n N_A_845_69#_c_3575_n 0.00436105f $X=4.485 $Y=0.18 $X2=0
+ $Y2=0
cc_601 N_S[1]_c_622_n N_A_845_69#_c_3577_n 0.00139422f $X=4.98 $Y=0.255 $X2=0
+ $Y2=0
cc_602 N_A_701_47#_c_681_n N_D[1]_M1022_g 0.00671996f $X=4.86 $Y=1.4 $X2=0 $Y2=0
cc_603 N_A_701_47#_M1056_g N_D[1]_M1022_g 0.0241475f $X=4.95 $Y=2.075 $X2=0
+ $Y2=0
cc_604 N_A_701_47#_c_684_n N_VPWR_c_2002_n 0.0321301f $X=3.725 $Y=2.31 $X2=0
+ $Y2=0
cc_605 N_A_701_47#_c_679_n N_VPWR_c_2002_n 0.00732952f $X=4.01 $Y=1.42 $X2=0
+ $Y2=0
cc_606 N_A_701_47#_M1056_g N_VPWR_c_2003_n 0.00107974f $X=4.95 $Y=2.075 $X2=0
+ $Y2=0
cc_607 N_A_701_47#_M1045_d VPWR 0.00179197f $X=3.58 $Y=1.485 $X2=0 $Y2=0
cc_608 N_A_701_47#_M1040_g VPWR 0.00728421f $X=4.48 $Y=2.075 $X2=0 $Y2=0
cc_609 N_A_701_47#_M1056_g VPWR 0.00615305f $X=4.95 $Y=2.075 $X2=0 $Y2=0
cc_610 N_A_701_47#_c_684_n VPWR 0.00594162f $X=3.725 $Y=2.31 $X2=0 $Y2=0
cc_611 N_A_701_47#_M1040_g N_VPWR_c_2023_n 0.00429453f $X=4.48 $Y=2.075 $X2=0
+ $Y2=0
cc_612 N_A_701_47#_M1056_g N_VPWR_c_2023_n 0.00429453f $X=4.95 $Y=2.075 $X2=0
+ $Y2=0
cc_613 N_A_701_47#_c_684_n N_VPWR_c_2023_n 0.0210596f $X=3.725 $Y=2.31 $X2=0
+ $Y2=0
cc_614 N_A_701_47#_c_681_n N_Z_c_2369_n 0.00348752f $X=4.86 $Y=1.4 $X2=0 $Y2=0
cc_615 N_A_701_47#_c_677_n N_Z_c_2369_n 0.0033343f $X=4.01 $Y=1.205 $X2=0 $Y2=0
cc_616 N_A_701_47#_M1040_g N_Z_c_2384_n 0.00753886f $X=4.48 $Y=2.075 $X2=0 $Y2=0
cc_617 N_A_701_47#_c_676_n N_Z_c_2384_n 9.57301e-19 $X=4.57 $Y=1.4 $X2=0 $Y2=0
cc_618 N_A_701_47#_c_684_n N_Z_c_2384_n 0.0308332f $X=3.725 $Y=2.31 $X2=0 $Y2=0
cc_619 N_A_701_47#_c_679_n N_Z_c_2384_n 0.0132841f $X=4.01 $Y=1.42 $X2=0 $Y2=0
cc_620 N_A_701_47#_M1056_g N_Z_c_2385_n 0.00411531f $X=4.95 $Y=2.075 $X2=0 $Y2=0
cc_621 N_A_701_47#_M1056_g N_Z_c_2441_n 0.00513826f $X=4.95 $Y=2.075 $X2=0 $Y2=0
cc_622 N_A_701_47#_M1040_g N_Z_c_2442_n 0.00635536f $X=4.48 $Y=2.075 $X2=0 $Y2=0
cc_623 N_A_701_47#_c_681_n N_Z_c_2442_n 8.37785e-19 $X=4.86 $Y=1.4 $X2=0 $Y2=0
cc_624 N_A_701_47#_M1056_g N_Z_c_2442_n 0.0105371f $X=4.95 $Y=2.075 $X2=0 $Y2=0
cc_625 N_A_701_47#_M1040_g N_Z_c_2377_n 0.00476154f $X=4.48 $Y=2.075 $X2=0 $Y2=0
cc_626 N_A_701_47#_c_681_n N_Z_c_2377_n 0.0140509f $X=4.86 $Y=1.4 $X2=0 $Y2=0
cc_627 N_A_701_47#_c_676_n N_Z_c_2377_n 7.26438e-19 $X=4.57 $Y=1.4 $X2=0 $Y2=0
cc_628 N_A_701_47#_M1056_g N_Z_c_2377_n 0.00268051f $X=4.95 $Y=2.075 $X2=0 $Y2=0
cc_629 N_A_701_47#_c_677_n N_Z_c_2377_n 0.00967956f $X=4.01 $Y=1.205 $X2=0 $Y2=0
cc_630 N_A_701_47#_c_679_n N_Z_c_2377_n 0.0117695f $X=4.01 $Y=1.42 $X2=0 $Y2=0
cc_631 N_A_701_47#_M1040_g N_A_824_333#_c_2850_n 0.00745341f $X=4.48 $Y=2.075
+ $X2=0 $Y2=0
cc_632 N_A_701_47#_c_676_n N_A_824_333#_c_2850_n 0.00133381f $X=4.57 $Y=1.4
+ $X2=0 $Y2=0
cc_633 N_A_701_47#_c_684_n N_A_824_333#_c_2850_n 0.0347621f $X=3.725 $Y=2.31
+ $X2=0 $Y2=0
cc_634 N_A_701_47#_c_679_n N_A_824_333#_c_2850_n 0.0132748f $X=4.01 $Y=1.42
+ $X2=0 $Y2=0
cc_635 N_A_701_47#_M1040_g N_A_824_333#_c_2858_n 0.00971609f $X=4.48 $Y=2.075
+ $X2=0 $Y2=0
cc_636 N_A_701_47#_M1056_g N_A_824_333#_c_2858_n 0.0111338f $X=4.95 $Y=2.075
+ $X2=0 $Y2=0
cc_637 N_A_701_47#_c_684_n N_A_824_333#_c_2860_n 0.010563f $X=3.725 $Y=2.31
+ $X2=0 $Y2=0
cc_638 N_A_701_47#_M1056_g N_A_824_333#_c_2861_n 0.00717732f $X=4.95 $Y=2.075
+ $X2=0 $Y2=0
cc_639 N_A_701_47#_M1056_g N_A_824_333#_c_2862_n 0.00176121f $X=4.95 $Y=2.075
+ $X2=0 $Y2=0
cc_640 N_A_701_47#_M1035_d VGND 0.00250855f $X=3.505 $Y=0.235 $X2=0 $Y2=0
cc_641 N_A_701_47#_c_678_n VGND 0.0186564f $X=3.64 $Y=0.495 $X2=0 $Y2=0
cc_642 N_A_701_47#_c_678_n N_VGND_c_3315_n 0.0173492f $X=3.64 $Y=0.495 $X2=0
+ $Y2=0
cc_643 N_A_701_47#_c_676_n N_A_845_69#_c_3578_n 0.00308807f $X=4.57 $Y=1.4 $X2=0
+ $Y2=0
cc_644 N_A_701_47#_c_677_n N_A_845_69#_c_3578_n 0.00101918f $X=4.01 $Y=1.205
+ $X2=0 $Y2=0
cc_645 N_A_701_47#_c_678_n N_A_845_69#_c_3578_n 0.0185512f $X=3.64 $Y=0.495
+ $X2=0 $Y2=0
cc_646 N_A_701_47#_c_679_n N_A_845_69#_c_3578_n 0.00285813f $X=4.01 $Y=1.42
+ $X2=0 $Y2=0
cc_647 N_A_701_47#_c_678_n N_A_845_69#_c_3575_n 0.00358194f $X=3.64 $Y=0.495
+ $X2=0 $Y2=0
cc_648 D[1] N_D[2]_c_807_n 0.0231965f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_649 N_D[1]_c_755_n N_D[2]_c_807_n 7.85936e-19 $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_650 D[1] N_D[2]_c_808_n 7.85936e-19 $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_651 N_D[1]_c_755_n N_D[2]_c_808_n 0.00603597f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_652 N_D[1]_M1022_g N_VPWR_c_2003_n 0.00919666f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_653 N_D[1]_M1049_g N_VPWR_c_2003_n 0.0031734f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_654 N_D[1]_M1022_g N_VPWR_c_2077_n 0.00295119f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_655 N_D[1]_M1049_g N_VPWR_c_2077_n 0.00314707f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_656 N_D[1]_M1022_g VPWR 0.00588601f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_657 N_D[1]_M1049_g VPWR 0.00822554f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_658 N_D[1]_M1022_g N_VPWR_c_2023_n 0.00622633f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_659 N_D[1]_M1049_g N_VPWR_c_2024_n 0.00652917f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_660 N_D[1]_M1022_g N_Z_c_2385_n 0.00431834f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_661 N_D[1]_M1049_g N_Z_c_2385_n 0.00406261f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_662 D[1] N_Z_c_2385_n 0.00125914f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_663 N_D[1]_M1022_g N_Z_c_2377_n 0.00112534f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_664 N_D[1]_M1036_g N_Z_c_2377_n 8.13311e-19 $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_665 D[1] N_Z_c_2377_n 0.00742792f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_666 N_D[1]_c_755_n N_Z_c_2377_n 0.00583073f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_667 N_D[1]_M1022_g N_A_824_333#_c_2861_n 0.00541465f $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_668 N_D[1]_M1022_g N_A_824_333#_c_2864_n 0.0127833f $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_669 N_D[1]_M1049_g N_A_824_333#_c_2864_n 0.0101085f $X=5.945 $Y=1.985 $X2=0
+ $Y2=0
cc_670 D[1] N_A_824_333#_c_2864_n 0.0323774f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_671 N_D[1]_c_755_n N_A_824_333#_c_2864_n 7.13708e-19 $X=6.03 $Y=1.16 $X2=0
+ $Y2=0
cc_672 D[1] N_A_824_333#_c_2851_n 0.0226682f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_673 N_D[1]_c_755_n N_A_824_333#_c_2851_n 9.6385e-19 $X=6.03 $Y=1.16 $X2=0
+ $Y2=0
cc_674 N_D[1]_M1049_g N_A_824_333#_c_2852_n 0.00325722f $X=5.945 $Y=1.985 $X2=0
+ $Y2=0
cc_675 N_D[1]_M1036_g N_VGND_c_3291_n 0.00300333f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_676 N_D[1]_M1051_g N_VGND_c_3291_n 0.0030929f $X=5.92 $Y=0.56 $X2=0 $Y2=0
cc_677 N_D[1]_M1051_g N_VGND_c_3292_n 0.00430643f $X=5.92 $Y=0.56 $X2=0 $Y2=0
cc_678 N_D[1]_M1036_g VGND 0.00600262f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_679 N_D[1]_M1051_g VGND 0.00733187f $X=5.92 $Y=0.56 $X2=0 $Y2=0
cc_680 N_D[1]_M1036_g N_VGND_c_3315_n 0.00436487f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_681 N_D[1]_M1036_g N_A_845_69#_c_3576_n 0.0114493f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_682 N_D[1]_M1051_g N_A_845_69#_c_3576_n 0.00931728f $X=5.92 $Y=0.56 $X2=0
+ $Y2=0
cc_683 D[1] N_A_845_69#_c_3576_n 0.0518587f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_684 N_D[1]_c_755_n N_A_845_69#_c_3576_n 0.00665175f $X=6.03 $Y=1.16 $X2=0
+ $Y2=0
cc_685 N_D[1]_M1036_g N_A_845_69#_c_3577_n 0.00114614f $X=5.5 $Y=0.56 $X2=0
+ $Y2=0
cc_686 N_D[1]_c_755_n N_A_845_69#_c_3577_n 0.00120541f $X=6.03 $Y=1.16 $X2=0
+ $Y2=0
cc_687 N_D[1]_M1036_g N_A_845_69#_c_3596_n 5.29024e-19 $X=5.5 $Y=0.56 $X2=0
+ $Y2=0
cc_688 N_D[1]_M1051_g N_A_845_69#_c_3596_n 0.00633603f $X=5.92 $Y=0.56 $X2=0
+ $Y2=0
cc_689 N_D[2]_M1060_g N_A_1566_265#_M1004_g 0.0241475f $X=7.405 $Y=1.985 $X2=0
+ $Y2=0
cc_690 N_D[2]_M1060_g N_A_1566_265#_c_863_n 0.00671996f $X=7.405 $Y=1.985 $X2=0
+ $Y2=0
cc_691 N_D[2]_M1063_g N_S[2]_c_937_n 0.0165585f $X=7.38 $Y=0.56 $X2=0 $Y2=0
cc_692 N_D[2]_M1000_g N_VPWR_c_2004_n 0.0031734f $X=6.935 $Y=1.985 $X2=0 $Y2=0
cc_693 N_D[2]_M1060_g N_VPWR_c_2004_n 0.00919666f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_694 N_D[2]_M1000_g N_VPWR_c_2085_n 0.00314707f $X=6.935 $Y=1.985 $X2=0 $Y2=0
cc_695 N_D[2]_M1060_g N_VPWR_c_2085_n 0.00295119f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_696 N_D[2]_M1060_g N_VPWR_c_2015_n 0.00622633f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_697 N_D[2]_M1000_g VPWR 0.00822554f $X=6.935 $Y=1.985 $X2=0 $Y2=0
cc_698 N_D[2]_M1060_g VPWR 0.00588601f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_699 N_D[2]_M1000_g N_VPWR_c_2024_n 0.00652917f $X=6.935 $Y=1.985 $X2=0 $Y2=0
cc_700 N_D[2]_M1000_g N_Z_c_2385_n 0.00406261f $X=6.935 $Y=1.985 $X2=0 $Y2=0
cc_701 N_D[2]_M1060_g N_Z_c_2385_n 0.00431834f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_702 N_D[2]_c_807_n N_Z_c_2385_n 0.00125914f $X=7.19 $Y=1.16 $X2=0 $Y2=0
cc_703 N_D[2]_M1063_g N_Z_c_2378_n 8.13311e-19 $X=7.38 $Y=0.56 $X2=0 $Y2=0
cc_704 N_D[2]_M1060_g N_Z_c_2378_n 0.00112534f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_705 N_D[2]_c_807_n N_Z_c_2378_n 0.00742792f $X=7.19 $Y=1.16 $X2=0 $Y2=0
cc_706 N_D[2]_c_808_n N_Z_c_2378_n 0.00583073f $X=7.405 $Y=1.16 $X2=0 $Y2=0
cc_707 N_D[2]_c_807_n N_A_1315_297#_c_2909_n 0.0226682f $X=7.19 $Y=1.16 $X2=0
+ $Y2=0
cc_708 N_D[2]_c_808_n N_A_1315_297#_c_2909_n 9.6385e-19 $X=7.405 $Y=1.16 $X2=0
+ $Y2=0
cc_709 N_D[2]_M1000_g N_A_1315_297#_c_2915_n 0.0101085f $X=6.935 $Y=1.985 $X2=0
+ $Y2=0
cc_710 N_D[2]_M1060_g N_A_1315_297#_c_2915_n 0.0127833f $X=7.405 $Y=1.985 $X2=0
+ $Y2=0
cc_711 N_D[2]_c_807_n N_A_1315_297#_c_2915_n 0.0323774f $X=7.19 $Y=1.16 $X2=0
+ $Y2=0
cc_712 N_D[2]_c_808_n N_A_1315_297#_c_2915_n 7.13708e-19 $X=7.405 $Y=1.16 $X2=0
+ $Y2=0
cc_713 N_D[2]_M1060_g N_A_1315_297#_c_2919_n 0.00541465f $X=7.405 $Y=1.985 $X2=0
+ $Y2=0
cc_714 N_D[2]_M1000_g N_A_1315_297#_c_2911_n 0.00325722f $X=6.935 $Y=1.985 $X2=0
+ $Y2=0
cc_715 N_D[2]_M1057_g N_VGND_c_3292_n 0.00430643f $X=6.96 $Y=0.56 $X2=0 $Y2=0
cc_716 N_D[2]_M1057_g N_VGND_c_3293_n 0.0030929f $X=6.96 $Y=0.56 $X2=0 $Y2=0
cc_717 N_D[2]_M1063_g N_VGND_c_3293_n 0.00300333f $X=7.38 $Y=0.56 $X2=0 $Y2=0
cc_718 N_D[2]_M1063_g N_VGND_c_3306_n 0.00436487f $X=7.38 $Y=0.56 $X2=0 $Y2=0
cc_719 N_D[2]_M1057_g VGND 0.00733187f $X=6.96 $Y=0.56 $X2=0 $Y2=0
cc_720 N_D[2]_M1063_g VGND 0.00600262f $X=7.38 $Y=0.56 $X2=0 $Y2=0
cc_721 N_D[2]_M1057_g N_A_1315_47#_c_3625_n 0.00633603f $X=6.96 $Y=0.56 $X2=0
+ $Y2=0
cc_722 N_D[2]_M1063_g N_A_1315_47#_c_3625_n 5.29024e-19 $X=7.38 $Y=0.56 $X2=0
+ $Y2=0
cc_723 N_D[2]_M1057_g N_A_1315_47#_c_3622_n 0.0084485f $X=6.96 $Y=0.56 $X2=0
+ $Y2=0
cc_724 N_D[2]_M1063_g N_A_1315_47#_c_3622_n 0.0125955f $X=7.38 $Y=0.56 $X2=0
+ $Y2=0
cc_725 N_D[2]_c_807_n N_A_1315_47#_c_3622_n 0.0274027f $X=7.19 $Y=1.16 $X2=0
+ $Y2=0
cc_726 N_D[2]_c_808_n N_A_1315_47#_c_3622_n 0.00321151f $X=7.405 $Y=1.16 $X2=0
+ $Y2=0
cc_727 N_D[2]_M1057_g N_A_1315_47#_c_3623_n 8.68782e-19 $X=6.96 $Y=0.56 $X2=0
+ $Y2=0
cc_728 N_D[2]_c_807_n N_A_1315_47#_c_3623_n 0.024456f $X=7.19 $Y=1.16 $X2=0
+ $Y2=0
cc_729 N_D[2]_c_808_n N_A_1315_47#_c_3623_n 0.00464565f $X=7.405 $Y=1.16 $X2=0
+ $Y2=0
cc_730 N_A_1566_265#_c_863_n N_S[2]_c_935_n 0.00779314f $X=8.02 $Y=1.4 $X2=-0.19
+ $Y2=-0.24
cc_731 N_A_1566_265#_c_862_n N_S[2]_c_938_n 0.00810157f $X=8.31 $Y=1.4 $X2=0
+ $Y2=0
cc_732 N_A_1566_265#_c_858_n N_S[2]_c_938_n 7.04048e-19 $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_733 N_A_1566_265#_c_857_n N_S[2]_c_940_n 0.0100587f $X=8.87 $Y=0.755 $X2=0
+ $Y2=0
cc_734 N_A_1566_265#_c_858_n N_S[2]_c_940_n 0.00267287f $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_735 N_A_1566_265#_c_857_n N_S[2]_c_941_n 0.0105766f $X=8.87 $Y=0.755 $X2=0
+ $Y2=0
cc_736 N_A_1566_265#_c_858_n N_S[2]_c_941_n 0.0090765f $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_737 N_A_1566_265#_c_859_n N_S[2]_c_941_n 0.00742826f $X=9.155 $Y=1.63 $X2=0
+ $Y2=0
cc_738 N_A_1566_265#_c_858_n N_S[2]_c_942_n 0.00445422f $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_739 N_A_1566_265#_c_859_n N_S[2]_c_942_n 4.25171e-19 $X=9.155 $Y=1.63 $X2=0
+ $Y2=0
cc_740 N_A_1566_265#_c_860_n N_S[2]_c_942_n 0.00920672f $X=8.4 $Y=1.34 $X2=0
+ $Y2=0
cc_741 N_A_1566_265#_c_858_n N_S[2]_c_943_n 0.00205356f $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_742 N_A_1566_265#_c_865_n N_S[2]_c_943_n 0.00862444f $X=9.155 $Y=2.31 $X2=0
+ $Y2=0
cc_743 N_A_1566_265#_c_859_n N_S[2]_c_943_n 0.00828481f $X=9.155 $Y=1.63 $X2=0
+ $Y2=0
cc_744 N_A_1566_265#_c_860_n N_S[2]_c_943_n 0.00692516f $X=8.4 $Y=1.34 $X2=0
+ $Y2=0
cc_745 N_A_1566_265#_c_858_n N_S[2]_c_944_n 0.00149517f $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_746 N_A_1566_265#_c_857_n S[2] 0.0061421f $X=8.87 $Y=0.755 $X2=0 $Y2=0
cc_747 N_A_1566_265#_c_858_n S[2] 0.0101733f $X=8.87 $Y=1.205 $X2=0 $Y2=0
cc_748 N_A_1566_265#_c_859_n S[2] 0.0127184f $X=9.155 $Y=1.63 $X2=0 $Y2=0
cc_749 N_A_1566_265#_c_860_n S[2] 3.07062e-19 $X=8.4 $Y=1.34 $X2=0 $Y2=0
cc_750 N_A_1566_265#_M1004_g N_VPWR_c_2004_n 0.00107974f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_751 N_A_1566_265#_c_865_n N_VPWR_c_2005_n 0.0321301f $X=9.155 $Y=2.31 $X2=0
+ $Y2=0
cc_752 N_A_1566_265#_c_859_n N_VPWR_c_2005_n 0.00732952f $X=9.155 $Y=1.63 $X2=0
+ $Y2=0
cc_753 N_A_1566_265#_M1004_g N_VPWR_c_2015_n 0.00429453f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_754 N_A_1566_265#_M1061_g N_VPWR_c_2015_n 0.00429453f $X=8.4 $Y=2.075 $X2=0
+ $Y2=0
cc_755 N_A_1566_265#_c_865_n N_VPWR_c_2015_n 0.0210596f $X=9.155 $Y=2.31 $X2=0
+ $Y2=0
cc_756 N_A_1566_265#_M1067_s VPWR 0.00179197f $X=9.03 $Y=1.485 $X2=0 $Y2=0
cc_757 N_A_1566_265#_M1004_g VPWR 0.00615305f $X=7.93 $Y=2.075 $X2=0 $Y2=0
cc_758 N_A_1566_265#_M1061_g VPWR 0.00728421f $X=8.4 $Y=2.075 $X2=0 $Y2=0
cc_759 N_A_1566_265#_c_865_n VPWR 0.00594162f $X=9.155 $Y=2.31 $X2=0 $Y2=0
cc_760 N_A_1566_265#_c_862_n N_Z_c_2370_n 0.00168443f $X=8.31 $Y=1.4 $X2=0 $Y2=0
cc_761 N_A_1566_265#_c_863_n N_Z_c_2370_n 0.00180308f $X=8.02 $Y=1.4 $X2=0 $Y2=0
cc_762 N_A_1566_265#_c_858_n N_Z_c_2370_n 0.0033343f $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_763 N_A_1566_265#_M1004_g N_Z_c_2385_n 0.00411531f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_764 N_A_1566_265#_M1061_g N_Z_c_2386_n 0.00753886f $X=8.4 $Y=2.075 $X2=0
+ $Y2=0
cc_765 N_A_1566_265#_c_865_n N_Z_c_2386_n 0.0308332f $X=9.155 $Y=2.31 $X2=0
+ $Y2=0
cc_766 N_A_1566_265#_c_859_n N_Z_c_2386_n 0.0132841f $X=9.155 $Y=1.63 $X2=0
+ $Y2=0
cc_767 N_A_1566_265#_c_860_n N_Z_c_2386_n 9.57301e-19 $X=8.4 $Y=1.34 $X2=0 $Y2=0
cc_768 N_A_1566_265#_M1004_g N_Z_c_2473_n 0.00513826f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_769 N_A_1566_265#_M1004_g N_Z_c_2474_n 0.0105371f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_770 N_A_1566_265#_c_862_n N_Z_c_2474_n 8.37785e-19 $X=8.31 $Y=1.4 $X2=0 $Y2=0
cc_771 N_A_1566_265#_M1061_g N_Z_c_2474_n 0.00635536f $X=8.4 $Y=2.075 $X2=0
+ $Y2=0
cc_772 N_A_1566_265#_M1004_g N_Z_c_2378_n 0.00268051f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_773 N_A_1566_265#_c_862_n N_Z_c_2378_n 0.0140509f $X=8.31 $Y=1.4 $X2=0 $Y2=0
cc_774 N_A_1566_265#_M1061_g N_Z_c_2378_n 0.00476154f $X=8.4 $Y=2.075 $X2=0
+ $Y2=0
cc_775 N_A_1566_265#_c_858_n N_Z_c_2378_n 0.00967956f $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_776 N_A_1566_265#_c_859_n N_Z_c_2378_n 0.0117695f $X=9.155 $Y=1.63 $X2=0
+ $Y2=0
cc_777 N_A_1566_265#_c_860_n N_Z_c_2378_n 7.26438e-19 $X=8.4 $Y=1.34 $X2=0 $Y2=0
cc_778 N_A_1566_265#_M1004_g N_A_1315_297#_c_2915_n 0.00176121f $X=7.93 $Y=2.075
+ $X2=0 $Y2=0
cc_779 N_A_1566_265#_M1004_g N_A_1315_297#_c_2919_n 0.00717732f $X=7.93 $Y=2.075
+ $X2=0 $Y2=0
cc_780 N_A_1566_265#_M1004_g N_A_1315_297#_c_2923_n 0.0111338f $X=7.93 $Y=2.075
+ $X2=0 $Y2=0
cc_781 N_A_1566_265#_M1061_g N_A_1315_297#_c_2923_n 0.00971609f $X=8.4 $Y=2.075
+ $X2=0 $Y2=0
cc_782 N_A_1566_265#_c_865_n N_A_1315_297#_c_2923_n 0.010563f $X=9.155 $Y=2.31
+ $X2=0 $Y2=0
cc_783 N_A_1566_265#_M1061_g N_A_1315_297#_c_2910_n 0.00745341f $X=8.4 $Y=2.075
+ $X2=0 $Y2=0
cc_784 N_A_1566_265#_c_865_n N_A_1315_297#_c_2910_n 0.0347621f $X=9.155 $Y=2.31
+ $X2=0 $Y2=0
cc_785 N_A_1566_265#_c_859_n N_A_1315_297#_c_2910_n 0.0132748f $X=9.155 $Y=1.63
+ $X2=0 $Y2=0
cc_786 N_A_1566_265#_c_860_n N_A_1315_297#_c_2910_n 0.00133381f $X=8.4 $Y=1.34
+ $X2=0 $Y2=0
cc_787 N_A_1566_265#_c_857_n N_VGND_c_3306_n 0.0173492f $X=8.87 $Y=0.755 $X2=0
+ $Y2=0
cc_788 N_A_1566_265#_M1077_s VGND 0.00250855f $X=9.115 $Y=0.235 $X2=0 $Y2=0
cc_789 N_A_1566_265#_c_857_n VGND 0.0186564f $X=8.87 $Y=0.755 $X2=0 $Y2=0
cc_790 N_A_1566_265#_c_857_n N_A_1315_47#_c_3624_n 0.00358194f $X=8.87 $Y=0.755
+ $X2=0 $Y2=0
cc_791 N_A_1566_265#_c_857_n N_A_1315_47#_c_3635_n 0.0185512f $X=8.87 $Y=0.755
+ $X2=0 $Y2=0
cc_792 N_A_1566_265#_c_858_n N_A_1315_47#_c_3635_n 0.00101918f $X=8.87 $Y=1.205
+ $X2=0 $Y2=0
cc_793 N_A_1566_265#_c_859_n N_A_1315_47#_c_3635_n 0.00285813f $X=9.155 $Y=1.63
+ $X2=0 $Y2=0
cc_794 N_A_1566_265#_c_860_n N_A_1315_47#_c_3635_n 0.00308807f $X=8.4 $Y=1.34
+ $X2=0 $Y2=0
cc_795 N_S[2]_c_944_n N_S[3]_c_1000_n 0.0133556f $X=9.45 $Y=0.845 $X2=-0.19
+ $Y2=-0.24
cc_796 N_S[2]_c_943_n N_S[3]_c_1001_n 0.0418422f $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_797 S[2] N_S[3]_c_1001_n 8.74983e-19 $X=9.345 $Y=1.105 $X2=0 $Y2=0
cc_798 N_S[2]_c_943_n S[3] 8.74983e-19 $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_799 S[2] S[3] 0.0208489f $X=9.345 $Y=1.105 $X2=0 $Y2=0
cc_800 N_S[2]_c_943_n N_VPWR_c_2005_n 0.00456891f $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_801 S[2] N_VPWR_c_2005_n 0.00569857f $X=9.345 $Y=1.105 $X2=0 $Y2=0
cc_802 N_S[2]_c_943_n N_VPWR_c_2015_n 0.00673617f $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_803 N_S[2]_c_943_n VPWR 0.00852379f $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_804 N_S[2]_c_935_n N_Z_c_2370_n 0.00413022f $X=7.9 $Y=0.255 $X2=0 $Y2=0
cc_805 N_S[2]_c_938_n N_Z_c_2370_n 0.00495983f $X=8.32 $Y=0.255 $X2=0 $Y2=0
cc_806 N_S[2]_c_940_n N_Z_c_2370_n 4.25992e-19 $X=8.805 $Y=0.845 $X2=0 $Y2=0
cc_807 N_S[2]_c_943_n N_Z_c_2386_n 0.00513674f $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_808 S[2] N_Z_c_2386_n 0.00545567f $X=9.345 $Y=1.105 $X2=0 $Y2=0
cc_809 N_S[2]_c_935_n N_Z_c_2378_n 0.00199103f $X=7.9 $Y=0.255 $X2=0 $Y2=0
cc_810 N_S[2]_c_938_n N_Z_c_2378_n 0.00133607f $X=8.32 $Y=0.255 $X2=0 $Y2=0
cc_811 N_S[2]_c_944_n N_VGND_c_3294_n 0.00330937f $X=9.45 $Y=0.845 $X2=0 $Y2=0
cc_812 N_S[2]_c_937_n N_VGND_c_3306_n 0.0271255f $X=7.975 $Y=0.18 $X2=0 $Y2=0
cc_813 N_S[2]_c_944_n N_VGND_c_3306_n 0.00585385f $X=9.45 $Y=0.845 $X2=0 $Y2=0
cc_814 N_S[2]_c_936_n VGND 0.00642387f $X=8.245 $Y=0.18 $X2=0 $Y2=0
cc_815 N_S[2]_c_937_n VGND 0.00474746f $X=7.975 $Y=0.18 $X2=0 $Y2=0
cc_816 N_S[2]_c_939_n VGND 0.0193094f $X=8.73 $Y=0.18 $X2=0 $Y2=0
cc_817 N_S[2]_c_944_n VGND 0.0111218f $X=9.45 $Y=0.845 $X2=0 $Y2=0
cc_818 N_S[2]_c_945_n VGND 0.00366655f $X=8.32 $Y=0.18 $X2=0 $Y2=0
cc_819 N_S[2]_c_935_n N_A_1315_47#_c_3622_n 0.00139422f $X=7.9 $Y=0.255 $X2=0
+ $Y2=0
cc_820 N_S[2]_c_935_n N_A_1315_47#_c_3624_n 0.0132844f $X=7.9 $Y=0.255 $X2=0
+ $Y2=0
cc_821 N_S[2]_c_936_n N_A_1315_47#_c_3624_n 0.00211351f $X=8.245 $Y=0.18 $X2=0
+ $Y2=0
cc_822 N_S[2]_c_938_n N_A_1315_47#_c_3624_n 0.0126455f $X=8.32 $Y=0.255 $X2=0
+ $Y2=0
cc_823 N_S[2]_c_939_n N_A_1315_47#_c_3624_n 0.00436105f $X=8.73 $Y=0.18 $X2=0
+ $Y2=0
cc_824 N_S[2]_c_940_n N_A_1315_47#_c_3624_n 0.00349455f $X=8.805 $Y=0.845 $X2=0
+ $Y2=0
cc_825 N_S[2]_c_940_n N_A_1315_47#_c_3635_n 0.00295202f $X=8.805 $Y=0.845 $X2=0
+ $Y2=0
cc_826 N_S[3]_c_1008_n N_A_1989_47#_c_1067_n 0.00779314f $X=11.42 $Y=0.255 $X2=0
+ $Y2=0
cc_827 N_S[3]_c_1001_n N_A_1989_47#_c_1062_n 0.00692516f $X=9.93 $Y=1.41 $X2=0
+ $Y2=0
cc_828 N_S[3]_c_1002_n N_A_1989_47#_c_1062_n 0.00920672f $X=10.44 $Y=0.92 $X2=0
+ $Y2=0
cc_829 N_S[3]_c_1006_n N_A_1989_47#_c_1062_n 0.00810157f $X=11 $Y=0.255 $X2=0
+ $Y2=0
cc_830 S[3] N_A_1989_47#_c_1062_n 3.07062e-19 $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_831 N_S[3]_c_1001_n N_A_1989_47#_c_1070_n 0.00862444f $X=9.93 $Y=1.41 $X2=0
+ $Y2=0
cc_832 N_S[3]_c_1000_n N_A_1989_47#_c_1063_n 0.00149517f $X=9.87 $Y=0.845 $X2=0
+ $Y2=0
cc_833 N_S[3]_c_1001_n N_A_1989_47#_c_1063_n 0.00205356f $X=9.93 $Y=1.41 $X2=0
+ $Y2=0
cc_834 N_S[3]_c_1002_n N_A_1989_47#_c_1063_n 0.0135307f $X=10.44 $Y=0.92 $X2=0
+ $Y2=0
cc_835 N_S[3]_c_1003_n N_A_1989_47#_c_1063_n 0.00267287f $X=10.515 $Y=0.845
+ $X2=0 $Y2=0
cc_836 N_S[3]_c_1006_n N_A_1989_47#_c_1063_n 7.04048e-19 $X=11 $Y=0.255 $X2=0
+ $Y2=0
cc_837 S[3] N_A_1989_47#_c_1063_n 0.0101733f $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_838 N_S[3]_c_1001_n N_A_1989_47#_c_1064_n 0.0105766f $X=9.93 $Y=1.41 $X2=0
+ $Y2=0
cc_839 N_S[3]_c_1003_n N_A_1989_47#_c_1064_n 0.0100587f $X=10.515 $Y=0.845 $X2=0
+ $Y2=0
cc_840 S[3] N_A_1989_47#_c_1064_n 0.0061421f $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_841 N_S[3]_c_1001_n N_A_1989_47#_c_1065_n 0.00828481f $X=9.93 $Y=1.41 $X2=0
+ $Y2=0
cc_842 N_S[3]_c_1002_n N_A_1989_47#_c_1065_n 0.00785343f $X=10.44 $Y=0.92 $X2=0
+ $Y2=0
cc_843 S[3] N_A_1989_47#_c_1065_n 0.0127184f $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_844 N_S[3]_c_1007_n N_D[3]_M1012_g 0.0165585f $X=11.345 $Y=0.18 $X2=0 $Y2=0
cc_845 N_S[3]_c_1001_n N_VPWR_c_2005_n 0.00456891f $X=9.93 $Y=1.41 $X2=0 $Y2=0
cc_846 S[3] N_VPWR_c_2005_n 0.00569857f $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_847 N_S[3]_c_1001_n VPWR 0.00852379f $X=9.93 $Y=1.41 $X2=0 $Y2=0
cc_848 N_S[3]_c_1001_n N_VPWR_c_2025_n 0.00673617f $X=9.93 $Y=1.41 $X2=0 $Y2=0
cc_849 N_S[3]_c_1003_n N_Z_c_2371_n 4.25992e-19 $X=10.515 $Y=0.845 $X2=0 $Y2=0
cc_850 N_S[3]_c_1006_n N_Z_c_2371_n 0.00495983f $X=11 $Y=0.255 $X2=0 $Y2=0
cc_851 N_S[3]_c_1008_n N_Z_c_2371_n 0.00413022f $X=11.42 $Y=0.255 $X2=0 $Y2=0
cc_852 N_S[3]_c_1001_n N_Z_c_2386_n 0.00513674f $X=9.93 $Y=1.41 $X2=0 $Y2=0
cc_853 S[3] N_Z_c_2386_n 0.00545567f $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_854 N_S[3]_c_1006_n N_Z_c_2379_n 0.00133607f $X=11 $Y=0.255 $X2=0 $Y2=0
cc_855 N_S[3]_c_1008_n N_Z_c_2379_n 0.00199103f $X=11.42 $Y=0.255 $X2=0 $Y2=0
cc_856 N_S[3]_c_1000_n N_VGND_c_3294_n 0.00330937f $X=9.87 $Y=0.845 $X2=0 $Y2=0
cc_857 N_S[3]_c_1000_n VGND 0.0111218f $X=9.87 $Y=0.845 $X2=0 $Y2=0
cc_858 N_S[3]_c_1004_n VGND 0.0119932f $X=10.925 $Y=0.18 $X2=0 $Y2=0
cc_859 N_S[3]_c_1005_n VGND 0.00731624f $X=10.59 $Y=0.18 $X2=0 $Y2=0
cc_860 N_S[3]_c_1007_n VGND 0.0111713f $X=11.345 $Y=0.18 $X2=0 $Y2=0
cc_861 N_S[3]_c_1009_n VGND 0.00366655f $X=11 $Y=0.18 $X2=0 $Y2=0
cc_862 N_S[3]_c_1000_n N_VGND_c_3316_n 0.00585385f $X=9.87 $Y=0.845 $X2=0 $Y2=0
cc_863 N_S[3]_c_1005_n N_VGND_c_3316_n 0.0271255f $X=10.59 $Y=0.18 $X2=0 $Y2=0
cc_864 N_S[3]_c_1003_n N_A_2133_69#_c_3670_n 0.00295202f $X=10.515 $Y=0.845
+ $X2=0 $Y2=0
cc_865 N_S[3]_c_1006_n N_A_2133_69#_c_3666_n 0.0126455f $X=11 $Y=0.255 $X2=0
+ $Y2=0
cc_866 N_S[3]_c_1007_n N_A_2133_69#_c_3666_n 0.00211351f $X=11.345 $Y=0.18 $X2=0
+ $Y2=0
cc_867 N_S[3]_c_1008_n N_A_2133_69#_c_3666_n 0.0132844f $X=11.42 $Y=0.255 $X2=0
+ $Y2=0
cc_868 N_S[3]_c_1003_n N_A_2133_69#_c_3667_n 0.00349455f $X=10.515 $Y=0.845
+ $X2=0 $Y2=0
cc_869 N_S[3]_c_1004_n N_A_2133_69#_c_3667_n 0.00436105f $X=10.925 $Y=0.18 $X2=0
+ $Y2=0
cc_870 N_S[3]_c_1008_n N_A_2133_69#_c_3669_n 0.00139422f $X=11.42 $Y=0.255 $X2=0
+ $Y2=0
cc_871 N_A_1989_47#_c_1067_n N_D[3]_M1001_g 0.00671996f $X=11.3 $Y=1.4 $X2=0
+ $Y2=0
cc_872 N_A_1989_47#_M1062_g N_D[3]_M1001_g 0.0241475f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_873 N_A_1989_47#_c_1070_n N_VPWR_c_2005_n 0.0321301f $X=10.165 $Y=2.31 $X2=0
+ $Y2=0
cc_874 N_A_1989_47#_c_1065_n N_VPWR_c_2005_n 0.00732952f $X=10.45 $Y=1.42 $X2=0
+ $Y2=0
cc_875 N_A_1989_47#_M1062_g N_VPWR_c_2006_n 0.00107974f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_876 N_A_1989_47#_M1023_d VPWR 0.00179197f $X=10.02 $Y=1.485 $X2=0 $Y2=0
cc_877 N_A_1989_47#_M1005_g VPWR 0.00728421f $X=10.92 $Y=2.075 $X2=0 $Y2=0
cc_878 N_A_1989_47#_M1062_g VPWR 0.00615305f $X=11.39 $Y=2.075 $X2=0 $Y2=0
cc_879 N_A_1989_47#_c_1070_n VPWR 0.00594162f $X=10.165 $Y=2.31 $X2=0 $Y2=0
cc_880 N_A_1989_47#_M1005_g N_VPWR_c_2025_n 0.00429453f $X=10.92 $Y=2.075 $X2=0
+ $Y2=0
cc_881 N_A_1989_47#_M1062_g N_VPWR_c_2025_n 0.00429453f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_882 N_A_1989_47#_c_1070_n N_VPWR_c_2025_n 0.0210596f $X=10.165 $Y=2.31 $X2=0
+ $Y2=0
cc_883 N_A_1989_47#_c_1067_n N_Z_c_2371_n 0.00348752f $X=11.3 $Y=1.4 $X2=0 $Y2=0
cc_884 N_A_1989_47#_c_1063_n N_Z_c_2371_n 0.0033343f $X=10.45 $Y=1.205 $X2=0
+ $Y2=0
cc_885 N_A_1989_47#_M1005_g N_Z_c_2386_n 0.00753886f $X=10.92 $Y=2.075 $X2=0
+ $Y2=0
cc_886 N_A_1989_47#_c_1062_n N_Z_c_2386_n 9.57301e-19 $X=11.01 $Y=1.4 $X2=0
+ $Y2=0
cc_887 N_A_1989_47#_c_1070_n N_Z_c_2386_n 0.0308332f $X=10.165 $Y=2.31 $X2=0
+ $Y2=0
cc_888 N_A_1989_47#_c_1065_n N_Z_c_2386_n 0.0132841f $X=10.45 $Y=1.42 $X2=0
+ $Y2=0
cc_889 N_A_1989_47#_M1062_g N_Z_c_2387_n 0.00411531f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_890 N_A_1989_47#_M1062_g N_Z_c_2504_n 0.00513826f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_891 N_A_1989_47#_M1005_g N_Z_c_2505_n 0.00635536f $X=10.92 $Y=2.075 $X2=0
+ $Y2=0
cc_892 N_A_1989_47#_c_1067_n N_Z_c_2505_n 8.37785e-19 $X=11.3 $Y=1.4 $X2=0 $Y2=0
cc_893 N_A_1989_47#_M1062_g N_Z_c_2505_n 0.0105371f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_894 N_A_1989_47#_M1005_g N_Z_c_2379_n 0.00476154f $X=10.92 $Y=2.075 $X2=0
+ $Y2=0
cc_895 N_A_1989_47#_c_1067_n N_Z_c_2379_n 0.0140509f $X=11.3 $Y=1.4 $X2=0 $Y2=0
cc_896 N_A_1989_47#_c_1062_n N_Z_c_2379_n 7.26438e-19 $X=11.01 $Y=1.4 $X2=0
+ $Y2=0
cc_897 N_A_1989_47#_M1062_g N_Z_c_2379_n 0.00268051f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_898 N_A_1989_47#_c_1063_n N_Z_c_2379_n 0.00967956f $X=10.45 $Y=1.205 $X2=0
+ $Y2=0
cc_899 N_A_1989_47#_c_1065_n N_Z_c_2379_n 0.0117695f $X=10.45 $Y=1.42 $X2=0
+ $Y2=0
cc_900 N_A_1989_47#_M1005_g N_A_2112_333#_c_2966_n 0.00745341f $X=10.92 $Y=2.075
+ $X2=0 $Y2=0
cc_901 N_A_1989_47#_c_1062_n N_A_2112_333#_c_2966_n 0.00133381f $X=11.01 $Y=1.4
+ $X2=0 $Y2=0
cc_902 N_A_1989_47#_c_1070_n N_A_2112_333#_c_2966_n 0.0347621f $X=10.165 $Y=2.31
+ $X2=0 $Y2=0
cc_903 N_A_1989_47#_c_1065_n N_A_2112_333#_c_2966_n 0.0132748f $X=10.45 $Y=1.42
+ $X2=0 $Y2=0
cc_904 N_A_1989_47#_M1005_g N_A_2112_333#_c_2974_n 0.00971609f $X=10.92 $Y=2.075
+ $X2=0 $Y2=0
cc_905 N_A_1989_47#_M1062_g N_A_2112_333#_c_2974_n 0.0111338f $X=11.39 $Y=2.075
+ $X2=0 $Y2=0
cc_906 N_A_1989_47#_c_1070_n N_A_2112_333#_c_2976_n 0.010563f $X=10.165 $Y=2.31
+ $X2=0 $Y2=0
cc_907 N_A_1989_47#_M1062_g N_A_2112_333#_c_2977_n 0.00717732f $X=11.39 $Y=2.075
+ $X2=0 $Y2=0
cc_908 N_A_1989_47#_M1062_g N_A_2112_333#_c_2978_n 0.00176121f $X=11.39 $Y=2.075
+ $X2=0 $Y2=0
cc_909 N_A_1989_47#_M1009_d VGND 0.00250855f $X=9.945 $Y=0.235 $X2=0 $Y2=0
cc_910 N_A_1989_47#_c_1064_n VGND 0.0186564f $X=10.08 $Y=0.495 $X2=0 $Y2=0
cc_911 N_A_1989_47#_c_1064_n N_VGND_c_3316_n 0.0173492f $X=10.08 $Y=0.495 $X2=0
+ $Y2=0
cc_912 N_A_1989_47#_c_1062_n N_A_2133_69#_c_3670_n 0.00308807f $X=11.01 $Y=1.4
+ $X2=0 $Y2=0
cc_913 N_A_1989_47#_c_1063_n N_A_2133_69#_c_3670_n 0.00101918f $X=10.45 $Y=1.205
+ $X2=0 $Y2=0
cc_914 N_A_1989_47#_c_1064_n N_A_2133_69#_c_3670_n 0.0185512f $X=10.08 $Y=0.495
+ $X2=0 $Y2=0
cc_915 N_A_1989_47#_c_1065_n N_A_2133_69#_c_3670_n 0.00285813f $X=10.45 $Y=1.42
+ $X2=0 $Y2=0
cc_916 N_A_1989_47#_c_1064_n N_A_2133_69#_c_3667_n 0.00358194f $X=10.08 $Y=0.495
+ $X2=0 $Y2=0
cc_917 D[3] N_D[4]_c_1193_n 0.0231965f $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_918 N_D[3]_c_1141_n N_D[4]_c_1193_n 7.85936e-19 $X=12.47 $Y=1.16 $X2=0 $Y2=0
cc_919 D[3] N_D[4]_c_1194_n 7.85936e-19 $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_920 N_D[3]_c_1141_n N_D[4]_c_1194_n 0.00603597f $X=12.47 $Y=1.16 $X2=0 $Y2=0
cc_921 N_D[3]_M1001_g N_VPWR_c_2006_n 0.00919666f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_922 N_D[3]_M1068_g N_VPWR_c_2006_n 0.0031734f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_923 N_D[3]_M1001_g N_VPWR_c_2121_n 0.00295119f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_924 N_D[3]_M1068_g N_VPWR_c_2121_n 0.00314707f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_925 N_D[3]_M1001_g VPWR 0.00588601f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_926 N_D[3]_M1068_g VPWR 0.00822554f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_927 N_D[3]_M1001_g N_VPWR_c_2025_n 0.00622633f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_928 N_D[3]_M1068_g N_VPWR_c_2026_n 0.00652917f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_929 N_D[3]_M1001_g N_Z_c_2387_n 0.00431834f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_930 N_D[3]_M1068_g N_Z_c_2387_n 0.00406261f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_931 D[3] N_Z_c_2387_n 0.00125914f $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_932 N_D[3]_M1001_g N_Z_c_2379_n 0.00112534f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_933 N_D[3]_M1012_g N_Z_c_2379_n 8.13311e-19 $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_934 D[3] N_Z_c_2379_n 0.00742792f $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_935 N_D[3]_c_1141_n N_Z_c_2379_n 0.00583073f $X=12.47 $Y=1.16 $X2=0 $Y2=0
cc_936 N_D[3]_M1001_g N_A_2112_333#_c_2977_n 0.00541465f $X=11.915 $Y=1.985
+ $X2=0 $Y2=0
cc_937 N_D[3]_M1001_g N_A_2112_333#_c_2980_n 0.0127833f $X=11.915 $Y=1.985 $X2=0
+ $Y2=0
cc_938 N_D[3]_M1068_g N_A_2112_333#_c_2980_n 0.0101085f $X=12.385 $Y=1.985 $X2=0
+ $Y2=0
cc_939 D[3] N_A_2112_333#_c_2980_n 0.0323774f $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_940 N_D[3]_c_1141_n N_A_2112_333#_c_2980_n 7.13708e-19 $X=12.47 $Y=1.16 $X2=0
+ $Y2=0
cc_941 D[3] N_A_2112_333#_c_2967_n 0.0226682f $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_942 N_D[3]_c_1141_n N_A_2112_333#_c_2967_n 9.6385e-19 $X=12.47 $Y=1.16 $X2=0
+ $Y2=0
cc_943 N_D[3]_M1068_g N_A_2112_333#_c_2968_n 0.00325722f $X=12.385 $Y=1.985
+ $X2=0 $Y2=0
cc_944 N_D[3]_M1012_g N_VGND_c_3295_n 0.00300333f $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_945 N_D[3]_M1078_g N_VGND_c_3295_n 0.0030929f $X=12.36 $Y=0.56 $X2=0 $Y2=0
cc_946 N_D[3]_M1078_g N_VGND_c_3296_n 0.00430643f $X=12.36 $Y=0.56 $X2=0 $Y2=0
cc_947 N_D[3]_M1012_g VGND 0.00600262f $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_948 N_D[3]_M1078_g VGND 0.00733187f $X=12.36 $Y=0.56 $X2=0 $Y2=0
cc_949 N_D[3]_M1012_g N_VGND_c_3316_n 0.00436487f $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_950 N_D[3]_M1012_g N_A_2133_69#_c_3668_n 0.0114493f $X=11.94 $Y=0.56 $X2=0
+ $Y2=0
cc_951 N_D[3]_M1078_g N_A_2133_69#_c_3668_n 0.00931728f $X=12.36 $Y=0.56 $X2=0
+ $Y2=0
cc_952 D[3] N_A_2133_69#_c_3668_n 0.0518587f $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_953 N_D[3]_c_1141_n N_A_2133_69#_c_3668_n 0.00665175f $X=12.47 $Y=1.16 $X2=0
+ $Y2=0
cc_954 N_D[3]_M1012_g N_A_2133_69#_c_3669_n 0.00114614f $X=11.94 $Y=0.56 $X2=0
+ $Y2=0
cc_955 N_D[3]_c_1141_n N_A_2133_69#_c_3669_n 0.00120541f $X=12.47 $Y=1.16 $X2=0
+ $Y2=0
cc_956 N_D[3]_M1012_g N_A_2133_69#_c_3688_n 5.29024e-19 $X=11.94 $Y=0.56 $X2=0
+ $Y2=0
cc_957 N_D[3]_M1078_g N_A_2133_69#_c_3688_n 0.00633603f $X=12.36 $Y=0.56 $X2=0
+ $Y2=0
cc_958 N_D[4]_M1037_g N_A_2854_265#_M1016_g 0.0241475f $X=13.845 $Y=1.985 $X2=0
+ $Y2=0
cc_959 N_D[4]_M1037_g N_A_2854_265#_c_1249_n 0.00671996f $X=13.845 $Y=1.985
+ $X2=0 $Y2=0
cc_960 N_D[4]_M1048_g N_S[4]_c_1323_n 0.0165585f $X=13.82 $Y=0.56 $X2=0 $Y2=0
cc_961 N_D[4]_M1014_g N_VPWR_c_2007_n 0.0031734f $X=13.375 $Y=1.985 $X2=0 $Y2=0
cc_962 N_D[4]_M1037_g N_VPWR_c_2007_n 0.00919666f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_963 N_D[4]_M1014_g N_VPWR_c_2129_n 0.00314707f $X=13.375 $Y=1.985 $X2=0 $Y2=0
cc_964 N_D[4]_M1037_g N_VPWR_c_2129_n 0.00295119f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_965 N_D[4]_M1037_g N_VPWR_c_2017_n 0.00622633f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_966 N_D[4]_M1014_g VPWR 0.00822554f $X=13.375 $Y=1.985 $X2=0 $Y2=0
cc_967 N_D[4]_M1037_g VPWR 0.00588601f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_968 N_D[4]_M1014_g N_VPWR_c_2026_n 0.00652917f $X=13.375 $Y=1.985 $X2=0 $Y2=0
cc_969 N_D[4]_M1014_g N_Z_c_2387_n 0.00406261f $X=13.375 $Y=1.985 $X2=0 $Y2=0
cc_970 N_D[4]_M1037_g N_Z_c_2387_n 0.00431834f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_971 N_D[4]_c_1193_n N_Z_c_2387_n 0.00125914f $X=13.63 $Y=1.16 $X2=0 $Y2=0
cc_972 N_D[4]_M1048_g N_Z_c_2380_n 8.13311e-19 $X=13.82 $Y=0.56 $X2=0 $Y2=0
cc_973 N_D[4]_M1037_g N_Z_c_2380_n 0.00112534f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_974 N_D[4]_c_1193_n N_Z_c_2380_n 0.00742792f $X=13.63 $Y=1.16 $X2=0 $Y2=0
cc_975 N_D[4]_c_1194_n N_Z_c_2380_n 0.00583073f $X=13.845 $Y=1.16 $X2=0 $Y2=0
cc_976 N_D[4]_c_1193_n N_A_2603_297#_c_3025_n 0.0226682f $X=13.63 $Y=1.16 $X2=0
+ $Y2=0
cc_977 N_D[4]_c_1194_n N_A_2603_297#_c_3025_n 9.6385e-19 $X=13.845 $Y=1.16 $X2=0
+ $Y2=0
cc_978 N_D[4]_M1014_g N_A_2603_297#_c_3031_n 0.0101085f $X=13.375 $Y=1.985 $X2=0
+ $Y2=0
cc_979 N_D[4]_M1037_g N_A_2603_297#_c_3031_n 0.0127833f $X=13.845 $Y=1.985 $X2=0
+ $Y2=0
cc_980 N_D[4]_c_1193_n N_A_2603_297#_c_3031_n 0.0323774f $X=13.63 $Y=1.16 $X2=0
+ $Y2=0
cc_981 N_D[4]_c_1194_n N_A_2603_297#_c_3031_n 7.13708e-19 $X=13.845 $Y=1.16
+ $X2=0 $Y2=0
cc_982 N_D[4]_M1037_g N_A_2603_297#_c_3035_n 0.00541465f $X=13.845 $Y=1.985
+ $X2=0 $Y2=0
cc_983 N_D[4]_M1014_g N_A_2603_297#_c_3027_n 0.00325722f $X=13.375 $Y=1.985
+ $X2=0 $Y2=0
cc_984 N_D[4]_M1031_g N_VGND_c_3296_n 0.00430643f $X=13.4 $Y=0.56 $X2=0 $Y2=0
cc_985 N_D[4]_M1031_g N_VGND_c_3297_n 0.0030929f $X=13.4 $Y=0.56 $X2=0 $Y2=0
cc_986 N_D[4]_M1048_g N_VGND_c_3297_n 0.00300333f $X=13.82 $Y=0.56 $X2=0 $Y2=0
cc_987 N_D[4]_M1048_g N_VGND_c_3308_n 0.00436487f $X=13.82 $Y=0.56 $X2=0 $Y2=0
cc_988 N_D[4]_M1031_g VGND 0.00733187f $X=13.4 $Y=0.56 $X2=0 $Y2=0
cc_989 N_D[4]_M1048_g VGND 0.00600262f $X=13.82 $Y=0.56 $X2=0 $Y2=0
cc_990 N_D[4]_M1031_g N_A_2603_47#_c_3717_n 0.00633603f $X=13.4 $Y=0.56 $X2=0
+ $Y2=0
cc_991 N_D[4]_M1048_g N_A_2603_47#_c_3717_n 5.29024e-19 $X=13.82 $Y=0.56 $X2=0
+ $Y2=0
cc_992 N_D[4]_M1031_g N_A_2603_47#_c_3714_n 0.0084485f $X=13.4 $Y=0.56 $X2=0
+ $Y2=0
cc_993 N_D[4]_M1048_g N_A_2603_47#_c_3714_n 0.0125955f $X=13.82 $Y=0.56 $X2=0
+ $Y2=0
cc_994 N_D[4]_c_1193_n N_A_2603_47#_c_3714_n 0.0274027f $X=13.63 $Y=1.16 $X2=0
+ $Y2=0
cc_995 N_D[4]_c_1194_n N_A_2603_47#_c_3714_n 0.00321151f $X=13.845 $Y=1.16 $X2=0
+ $Y2=0
cc_996 N_D[4]_M1031_g N_A_2603_47#_c_3715_n 8.68782e-19 $X=13.4 $Y=0.56 $X2=0
+ $Y2=0
cc_997 N_D[4]_c_1193_n N_A_2603_47#_c_3715_n 0.024456f $X=13.63 $Y=1.16 $X2=0
+ $Y2=0
cc_998 N_D[4]_c_1194_n N_A_2603_47#_c_3715_n 0.00464565f $X=13.845 $Y=1.16 $X2=0
+ $Y2=0
cc_999 N_A_2854_265#_c_1249_n N_S[4]_c_1321_n 0.00779314f $X=14.46 $Y=1.4
+ $X2=-0.19 $Y2=-0.24
cc_1000 N_A_2854_265#_c_1248_n N_S[4]_c_1324_n 0.00810157f $X=14.75 $Y=1.4 $X2=0
+ $Y2=0
cc_1001 N_A_2854_265#_c_1244_n N_S[4]_c_1324_n 7.04048e-19 $X=15.31 $Y=1.205
+ $X2=0 $Y2=0
cc_1002 N_A_2854_265#_c_1243_n N_S[4]_c_1326_n 0.0100587f $X=15.31 $Y=0.755
+ $X2=0 $Y2=0
cc_1003 N_A_2854_265#_c_1244_n N_S[4]_c_1326_n 0.00267287f $X=15.31 $Y=1.205
+ $X2=0 $Y2=0
cc_1004 N_A_2854_265#_c_1243_n N_S[4]_c_1327_n 0.0105766f $X=15.31 $Y=0.755
+ $X2=0 $Y2=0
cc_1005 N_A_2854_265#_c_1244_n N_S[4]_c_1327_n 0.0090765f $X=15.31 $Y=1.205
+ $X2=0 $Y2=0
cc_1006 N_A_2854_265#_c_1245_n N_S[4]_c_1327_n 0.00742826f $X=15.595 $Y=1.63
+ $X2=0 $Y2=0
cc_1007 N_A_2854_265#_c_1244_n N_S[4]_c_1328_n 0.00445422f $X=15.31 $Y=1.205
+ $X2=0 $Y2=0
cc_1008 N_A_2854_265#_c_1245_n N_S[4]_c_1328_n 4.25171e-19 $X=15.595 $Y=1.63
+ $X2=0 $Y2=0
cc_1009 N_A_2854_265#_c_1246_n N_S[4]_c_1328_n 0.00920672f $X=14.84 $Y=1.34
+ $X2=0 $Y2=0
cc_1010 N_A_2854_265#_c_1244_n N_S[4]_c_1329_n 0.00205356f $X=15.31 $Y=1.205
+ $X2=0 $Y2=0
cc_1011 N_A_2854_265#_c_1251_n N_S[4]_c_1329_n 0.00862444f $X=15.595 $Y=2.31
+ $X2=0 $Y2=0
cc_1012 N_A_2854_265#_c_1245_n N_S[4]_c_1329_n 0.00828481f $X=15.595 $Y=1.63
+ $X2=0 $Y2=0
cc_1013 N_A_2854_265#_c_1246_n N_S[4]_c_1329_n 0.00692516f $X=14.84 $Y=1.34
+ $X2=0 $Y2=0
cc_1014 N_A_2854_265#_c_1244_n N_S[4]_c_1330_n 0.00149517f $X=15.31 $Y=1.205
+ $X2=0 $Y2=0
cc_1015 N_A_2854_265#_c_1243_n S[4] 0.0061421f $X=15.31 $Y=0.755 $X2=0 $Y2=0
cc_1016 N_A_2854_265#_c_1244_n S[4] 0.0101733f $X=15.31 $Y=1.205 $X2=0 $Y2=0
cc_1017 N_A_2854_265#_c_1245_n S[4] 0.0127184f $X=15.595 $Y=1.63 $X2=0 $Y2=0
cc_1018 N_A_2854_265#_c_1246_n S[4] 3.07062e-19 $X=14.84 $Y=1.34 $X2=0 $Y2=0
cc_1019 N_A_2854_265#_M1016_g N_VPWR_c_2007_n 0.00107974f $X=14.37 $Y=2.075
+ $X2=0 $Y2=0
cc_1020 N_A_2854_265#_c_1251_n N_VPWR_c_2008_n 0.0321301f $X=15.595 $Y=2.31
+ $X2=0 $Y2=0
cc_1021 N_A_2854_265#_c_1245_n N_VPWR_c_2008_n 0.00732952f $X=15.595 $Y=1.63
+ $X2=0 $Y2=0
cc_1022 N_A_2854_265#_M1016_g N_VPWR_c_2017_n 0.00429453f $X=14.37 $Y=2.075
+ $X2=0 $Y2=0
cc_1023 N_A_2854_265#_M1041_g N_VPWR_c_2017_n 0.00429453f $X=14.84 $Y=2.075
+ $X2=0 $Y2=0
cc_1024 N_A_2854_265#_c_1251_n N_VPWR_c_2017_n 0.0210596f $X=15.595 $Y=2.31
+ $X2=0 $Y2=0
cc_1025 N_A_2854_265#_M1002_s VPWR 0.00179197f $X=15.47 $Y=1.485 $X2=0 $Y2=0
cc_1026 N_A_2854_265#_M1016_g VPWR 0.00615305f $X=14.37 $Y=2.075 $X2=0 $Y2=0
cc_1027 N_A_2854_265#_M1041_g VPWR 0.00728421f $X=14.84 $Y=2.075 $X2=0 $Y2=0
cc_1028 N_A_2854_265#_c_1251_n VPWR 0.00594162f $X=15.595 $Y=2.31 $X2=0 $Y2=0
cc_1029 N_A_2854_265#_c_1248_n N_Z_c_2372_n 0.00168443f $X=14.75 $Y=1.4 $X2=0
+ $Y2=0
cc_1030 N_A_2854_265#_c_1249_n N_Z_c_2372_n 0.00180308f $X=14.46 $Y=1.4 $X2=0
+ $Y2=0
cc_1031 N_A_2854_265#_c_1244_n N_Z_c_2372_n 0.0033343f $X=15.31 $Y=1.205 $X2=0
+ $Y2=0
cc_1032 N_A_2854_265#_M1016_g N_Z_c_2387_n 0.00411531f $X=14.37 $Y=2.075 $X2=0
+ $Y2=0
cc_1033 N_A_2854_265#_M1041_g N_Z_c_2388_n 0.00753886f $X=14.84 $Y=2.075 $X2=0
+ $Y2=0
cc_1034 N_A_2854_265#_c_1251_n N_Z_c_2388_n 0.0308332f $X=15.595 $Y=2.31 $X2=0
+ $Y2=0
cc_1035 N_A_2854_265#_c_1245_n N_Z_c_2388_n 0.0132841f $X=15.595 $Y=1.63 $X2=0
+ $Y2=0
cc_1036 N_A_2854_265#_c_1246_n N_Z_c_2388_n 9.57301e-19 $X=14.84 $Y=1.34 $X2=0
+ $Y2=0
cc_1037 N_A_2854_265#_M1016_g N_Z_c_2536_n 0.00513826f $X=14.37 $Y=2.075 $X2=0
+ $Y2=0
cc_1038 N_A_2854_265#_M1016_g N_Z_c_2537_n 0.0105371f $X=14.37 $Y=2.075 $X2=0
+ $Y2=0
cc_1039 N_A_2854_265#_c_1248_n N_Z_c_2537_n 8.37785e-19 $X=14.75 $Y=1.4 $X2=0
+ $Y2=0
cc_1040 N_A_2854_265#_M1041_g N_Z_c_2537_n 0.00635536f $X=14.84 $Y=2.075 $X2=0
+ $Y2=0
cc_1041 N_A_2854_265#_M1016_g N_Z_c_2380_n 0.00268051f $X=14.37 $Y=2.075 $X2=0
+ $Y2=0
cc_1042 N_A_2854_265#_c_1248_n N_Z_c_2380_n 0.0140509f $X=14.75 $Y=1.4 $X2=0
+ $Y2=0
cc_1043 N_A_2854_265#_M1041_g N_Z_c_2380_n 0.00476154f $X=14.84 $Y=2.075 $X2=0
+ $Y2=0
cc_1044 N_A_2854_265#_c_1244_n N_Z_c_2380_n 0.00967956f $X=15.31 $Y=1.205 $X2=0
+ $Y2=0
cc_1045 N_A_2854_265#_c_1245_n N_Z_c_2380_n 0.0117695f $X=15.595 $Y=1.63 $X2=0
+ $Y2=0
cc_1046 N_A_2854_265#_c_1246_n N_Z_c_2380_n 7.26438e-19 $X=14.84 $Y=1.34 $X2=0
+ $Y2=0
cc_1047 N_A_2854_265#_M1016_g N_A_2603_297#_c_3031_n 0.00176121f $X=14.37
+ $Y=2.075 $X2=0 $Y2=0
cc_1048 N_A_2854_265#_M1016_g N_A_2603_297#_c_3035_n 0.00717732f $X=14.37
+ $Y=2.075 $X2=0 $Y2=0
cc_1049 N_A_2854_265#_M1016_g N_A_2603_297#_c_3039_n 0.0111338f $X=14.37
+ $Y=2.075 $X2=0 $Y2=0
cc_1050 N_A_2854_265#_M1041_g N_A_2603_297#_c_3039_n 0.00971609f $X=14.84
+ $Y=2.075 $X2=0 $Y2=0
cc_1051 N_A_2854_265#_c_1251_n N_A_2603_297#_c_3039_n 0.010563f $X=15.595
+ $Y=2.31 $X2=0 $Y2=0
cc_1052 N_A_2854_265#_M1041_g N_A_2603_297#_c_3026_n 0.00745341f $X=14.84
+ $Y=2.075 $X2=0 $Y2=0
cc_1053 N_A_2854_265#_c_1251_n N_A_2603_297#_c_3026_n 0.0347621f $X=15.595
+ $Y=2.31 $X2=0 $Y2=0
cc_1054 N_A_2854_265#_c_1245_n N_A_2603_297#_c_3026_n 0.0132748f $X=15.595
+ $Y=1.63 $X2=0 $Y2=0
cc_1055 N_A_2854_265#_c_1246_n N_A_2603_297#_c_3026_n 0.00133381f $X=14.84
+ $Y=1.34 $X2=0 $Y2=0
cc_1056 N_A_2854_265#_c_1243_n N_VGND_c_3308_n 0.0173492f $X=15.31 $Y=0.755
+ $X2=0 $Y2=0
cc_1057 N_A_2854_265#_M1032_s VGND 0.00250855f $X=15.555 $Y=0.235 $X2=0 $Y2=0
cc_1058 N_A_2854_265#_c_1243_n VGND 0.0186564f $X=15.31 $Y=0.755 $X2=0 $Y2=0
cc_1059 N_A_2854_265#_c_1243_n N_A_2603_47#_c_3716_n 0.00358194f $X=15.31
+ $Y=0.755 $X2=0 $Y2=0
cc_1060 N_A_2854_265#_c_1243_n N_A_2603_47#_c_3727_n 0.0185512f $X=15.31
+ $Y=0.755 $X2=0 $Y2=0
cc_1061 N_A_2854_265#_c_1244_n N_A_2603_47#_c_3727_n 0.00101918f $X=15.31
+ $Y=1.205 $X2=0 $Y2=0
cc_1062 N_A_2854_265#_c_1245_n N_A_2603_47#_c_3727_n 0.00285813f $X=15.595
+ $Y=1.63 $X2=0 $Y2=0
cc_1063 N_A_2854_265#_c_1246_n N_A_2603_47#_c_3727_n 0.00308807f $X=14.84
+ $Y=1.34 $X2=0 $Y2=0
cc_1064 N_S[4]_c_1330_n N_S[5]_c_1386_n 0.0133556f $X=15.89 $Y=0.845 $X2=-0.19
+ $Y2=-0.24
cc_1065 N_S[4]_c_1329_n N_S[5]_c_1387_n 0.0418422f $X=15.83 $Y=1.41 $X2=0 $Y2=0
cc_1066 S[4] N_S[5]_c_1387_n 8.74983e-19 $X=15.785 $Y=1.105 $X2=0 $Y2=0
cc_1067 N_S[4]_c_1329_n S[5] 8.74983e-19 $X=15.83 $Y=1.41 $X2=0 $Y2=0
cc_1068 S[4] S[5] 0.0208489f $X=15.785 $Y=1.105 $X2=0 $Y2=0
cc_1069 N_S[4]_c_1329_n N_VPWR_c_2008_n 0.00456891f $X=15.83 $Y=1.41 $X2=0 $Y2=0
cc_1070 S[4] N_VPWR_c_2008_n 0.00569857f $X=15.785 $Y=1.105 $X2=0 $Y2=0
cc_1071 N_S[4]_c_1329_n N_VPWR_c_2017_n 0.00673617f $X=15.83 $Y=1.41 $X2=0 $Y2=0
cc_1072 N_S[4]_c_1329_n VPWR 0.00852379f $X=15.83 $Y=1.41 $X2=0 $Y2=0
cc_1073 N_S[4]_c_1321_n N_Z_c_2372_n 0.00413022f $X=14.34 $Y=0.255 $X2=0 $Y2=0
cc_1074 N_S[4]_c_1324_n N_Z_c_2372_n 0.00495983f $X=14.76 $Y=0.255 $X2=0 $Y2=0
cc_1075 N_S[4]_c_1326_n N_Z_c_2372_n 4.25992e-19 $X=15.245 $Y=0.845 $X2=0 $Y2=0
cc_1076 N_S[4]_c_1329_n N_Z_c_2388_n 0.00513674f $X=15.83 $Y=1.41 $X2=0 $Y2=0
cc_1077 S[4] N_Z_c_2388_n 0.00545567f $X=15.785 $Y=1.105 $X2=0 $Y2=0
cc_1078 N_S[4]_c_1321_n N_Z_c_2380_n 0.00199103f $X=14.34 $Y=0.255 $X2=0 $Y2=0
cc_1079 N_S[4]_c_1324_n N_Z_c_2380_n 0.00133607f $X=14.76 $Y=0.255 $X2=0 $Y2=0
cc_1080 N_S[4]_c_1330_n N_VGND_c_3298_n 0.00330937f $X=15.89 $Y=0.845 $X2=0
+ $Y2=0
cc_1081 N_S[4]_c_1323_n N_VGND_c_3308_n 0.0271255f $X=14.415 $Y=0.18 $X2=0 $Y2=0
cc_1082 N_S[4]_c_1330_n N_VGND_c_3308_n 0.00585385f $X=15.89 $Y=0.845 $X2=0
+ $Y2=0
cc_1083 N_S[4]_c_1322_n VGND 0.00642387f $X=14.685 $Y=0.18 $X2=0 $Y2=0
cc_1084 N_S[4]_c_1323_n VGND 0.00474746f $X=14.415 $Y=0.18 $X2=0 $Y2=0
cc_1085 N_S[4]_c_1325_n VGND 0.0193094f $X=15.17 $Y=0.18 $X2=0 $Y2=0
cc_1086 N_S[4]_c_1330_n VGND 0.0111218f $X=15.89 $Y=0.845 $X2=0 $Y2=0
cc_1087 N_S[4]_c_1331_n VGND 0.00366655f $X=14.76 $Y=0.18 $X2=0 $Y2=0
cc_1088 N_S[4]_c_1321_n N_A_2603_47#_c_3714_n 0.00139422f $X=14.34 $Y=0.255
+ $X2=0 $Y2=0
cc_1089 N_S[4]_c_1321_n N_A_2603_47#_c_3716_n 0.0132844f $X=14.34 $Y=0.255 $X2=0
+ $Y2=0
cc_1090 N_S[4]_c_1322_n N_A_2603_47#_c_3716_n 0.00211351f $X=14.685 $Y=0.18
+ $X2=0 $Y2=0
cc_1091 N_S[4]_c_1324_n N_A_2603_47#_c_3716_n 0.0126455f $X=14.76 $Y=0.255 $X2=0
+ $Y2=0
cc_1092 N_S[4]_c_1325_n N_A_2603_47#_c_3716_n 0.00436105f $X=15.17 $Y=0.18 $X2=0
+ $Y2=0
cc_1093 N_S[4]_c_1326_n N_A_2603_47#_c_3716_n 0.00349455f $X=15.245 $Y=0.845
+ $X2=0 $Y2=0
cc_1094 N_S[4]_c_1326_n N_A_2603_47#_c_3727_n 0.00295202f $X=15.245 $Y=0.845
+ $X2=0 $Y2=0
cc_1095 N_S[5]_c_1394_n N_A_3277_47#_c_1453_n 0.00779314f $X=17.86 $Y=0.255
+ $X2=0 $Y2=0
cc_1096 N_S[5]_c_1387_n N_A_3277_47#_c_1448_n 0.00692516f $X=16.37 $Y=1.41 $X2=0
+ $Y2=0
cc_1097 N_S[5]_c_1388_n N_A_3277_47#_c_1448_n 0.00920672f $X=16.88 $Y=0.92 $X2=0
+ $Y2=0
cc_1098 N_S[5]_c_1392_n N_A_3277_47#_c_1448_n 0.00810157f $X=17.44 $Y=0.255
+ $X2=0 $Y2=0
cc_1099 S[5] N_A_3277_47#_c_1448_n 3.07062e-19 $X=16.245 $Y=1.105 $X2=0 $Y2=0
cc_1100 N_S[5]_c_1387_n N_A_3277_47#_c_1456_n 0.00862444f $X=16.37 $Y=1.41 $X2=0
+ $Y2=0
cc_1101 N_S[5]_c_1386_n N_A_3277_47#_c_1449_n 0.00149517f $X=16.31 $Y=0.845
+ $X2=0 $Y2=0
cc_1102 N_S[5]_c_1387_n N_A_3277_47#_c_1449_n 0.00205356f $X=16.37 $Y=1.41 $X2=0
+ $Y2=0
cc_1103 N_S[5]_c_1388_n N_A_3277_47#_c_1449_n 0.0135307f $X=16.88 $Y=0.92 $X2=0
+ $Y2=0
cc_1104 N_S[5]_c_1389_n N_A_3277_47#_c_1449_n 0.00267287f $X=16.955 $Y=0.845
+ $X2=0 $Y2=0
cc_1105 N_S[5]_c_1392_n N_A_3277_47#_c_1449_n 7.04048e-19 $X=17.44 $Y=0.255
+ $X2=0 $Y2=0
cc_1106 S[5] N_A_3277_47#_c_1449_n 0.0101733f $X=16.245 $Y=1.105 $X2=0 $Y2=0
cc_1107 N_S[5]_c_1387_n N_A_3277_47#_c_1450_n 0.0105766f $X=16.37 $Y=1.41 $X2=0
+ $Y2=0
cc_1108 N_S[5]_c_1389_n N_A_3277_47#_c_1450_n 0.0100587f $X=16.955 $Y=0.845
+ $X2=0 $Y2=0
cc_1109 S[5] N_A_3277_47#_c_1450_n 0.0061421f $X=16.245 $Y=1.105 $X2=0 $Y2=0
cc_1110 N_S[5]_c_1387_n N_A_3277_47#_c_1451_n 0.00828481f $X=16.37 $Y=1.41 $X2=0
+ $Y2=0
cc_1111 N_S[5]_c_1388_n N_A_3277_47#_c_1451_n 0.00785343f $X=16.88 $Y=0.92 $X2=0
+ $Y2=0
cc_1112 S[5] N_A_3277_47#_c_1451_n 0.0127184f $X=16.245 $Y=1.105 $X2=0 $Y2=0
cc_1113 N_S[5]_c_1393_n N_D[5]_M1047_g 0.0165585f $X=17.785 $Y=0.18 $X2=0 $Y2=0
cc_1114 N_S[5]_c_1387_n N_VPWR_c_2008_n 0.00456891f $X=16.37 $Y=1.41 $X2=0 $Y2=0
cc_1115 S[5] N_VPWR_c_2008_n 0.00569857f $X=16.245 $Y=1.105 $X2=0 $Y2=0
cc_1116 N_S[5]_c_1387_n VPWR 0.00852379f $X=16.37 $Y=1.41 $X2=0 $Y2=0
cc_1117 N_S[5]_c_1387_n N_VPWR_c_2027_n 0.00673617f $X=16.37 $Y=1.41 $X2=0 $Y2=0
cc_1118 N_S[5]_c_1389_n N_Z_c_2373_n 4.25992e-19 $X=16.955 $Y=0.845 $X2=0 $Y2=0
cc_1119 N_S[5]_c_1392_n N_Z_c_2373_n 0.00495983f $X=17.44 $Y=0.255 $X2=0 $Y2=0
cc_1120 N_S[5]_c_1394_n N_Z_c_2373_n 0.00413022f $X=17.86 $Y=0.255 $X2=0 $Y2=0
cc_1121 N_S[5]_c_1387_n N_Z_c_2388_n 0.00513674f $X=16.37 $Y=1.41 $X2=0 $Y2=0
cc_1122 S[5] N_Z_c_2388_n 0.00545567f $X=16.245 $Y=1.105 $X2=0 $Y2=0
cc_1123 N_S[5]_c_1392_n N_Z_c_2381_n 0.00133607f $X=17.44 $Y=0.255 $X2=0 $Y2=0
cc_1124 N_S[5]_c_1394_n N_Z_c_2381_n 0.00199103f $X=17.86 $Y=0.255 $X2=0 $Y2=0
cc_1125 N_S[5]_c_1386_n N_VGND_c_3298_n 0.00330937f $X=16.31 $Y=0.845 $X2=0
+ $Y2=0
cc_1126 N_S[5]_c_1386_n VGND 0.0111218f $X=16.31 $Y=0.845 $X2=0 $Y2=0
cc_1127 N_S[5]_c_1390_n VGND 0.0119932f $X=17.365 $Y=0.18 $X2=0 $Y2=0
cc_1128 N_S[5]_c_1391_n VGND 0.00731624f $X=17.03 $Y=0.18 $X2=0 $Y2=0
cc_1129 N_S[5]_c_1393_n VGND 0.0111713f $X=17.785 $Y=0.18 $X2=0 $Y2=0
cc_1130 N_S[5]_c_1395_n VGND 0.00366655f $X=17.44 $Y=0.18 $X2=0 $Y2=0
cc_1131 N_S[5]_c_1386_n N_VGND_c_3317_n 0.00585385f $X=16.31 $Y=0.845 $X2=0
+ $Y2=0
cc_1132 N_S[5]_c_1391_n N_VGND_c_3317_n 0.0271255f $X=17.03 $Y=0.18 $X2=0 $Y2=0
cc_1133 N_S[5]_c_1389_n N_A_3421_69#_c_3762_n 0.00295202f $X=16.955 $Y=0.845
+ $X2=0 $Y2=0
cc_1134 N_S[5]_c_1392_n N_A_3421_69#_c_3758_n 0.0126455f $X=17.44 $Y=0.255 $X2=0
+ $Y2=0
cc_1135 N_S[5]_c_1393_n N_A_3421_69#_c_3758_n 0.00211351f $X=17.785 $Y=0.18
+ $X2=0 $Y2=0
cc_1136 N_S[5]_c_1394_n N_A_3421_69#_c_3758_n 0.0132844f $X=17.86 $Y=0.255 $X2=0
+ $Y2=0
cc_1137 N_S[5]_c_1389_n N_A_3421_69#_c_3759_n 0.00349455f $X=16.955 $Y=0.845
+ $X2=0 $Y2=0
cc_1138 N_S[5]_c_1390_n N_A_3421_69#_c_3759_n 0.00436105f $X=17.365 $Y=0.18
+ $X2=0 $Y2=0
cc_1139 N_S[5]_c_1394_n N_A_3421_69#_c_3761_n 0.00139422f $X=17.86 $Y=0.255
+ $X2=0 $Y2=0
cc_1140 N_A_3277_47#_c_1453_n N_D[5]_M1025_g 0.00671996f $X=17.74 $Y=1.4 $X2=0
+ $Y2=0
cc_1141 N_A_3277_47#_M1042_g N_D[5]_M1025_g 0.0241475f $X=17.83 $Y=2.075 $X2=0
+ $Y2=0
cc_1142 N_A_3277_47#_c_1456_n N_VPWR_c_2008_n 0.0321301f $X=16.605 $Y=2.31 $X2=0
+ $Y2=0
cc_1143 N_A_3277_47#_c_1451_n N_VPWR_c_2008_n 0.00732952f $X=16.89 $Y=1.42 $X2=0
+ $Y2=0
cc_1144 N_A_3277_47#_M1042_g N_VPWR_c_2009_n 0.00107974f $X=17.83 $Y=2.075 $X2=0
+ $Y2=0
cc_1145 N_A_3277_47#_M1028_d VPWR 0.00179197f $X=16.46 $Y=1.485 $X2=0 $Y2=0
cc_1146 N_A_3277_47#_M1024_g VPWR 0.00728421f $X=17.36 $Y=2.075 $X2=0 $Y2=0
cc_1147 N_A_3277_47#_M1042_g VPWR 0.00615305f $X=17.83 $Y=2.075 $X2=0 $Y2=0
cc_1148 N_A_3277_47#_c_1456_n VPWR 0.00594162f $X=16.605 $Y=2.31 $X2=0 $Y2=0
cc_1149 N_A_3277_47#_M1024_g N_VPWR_c_2027_n 0.00429453f $X=17.36 $Y=2.075 $X2=0
+ $Y2=0
cc_1150 N_A_3277_47#_M1042_g N_VPWR_c_2027_n 0.00429453f $X=17.83 $Y=2.075 $X2=0
+ $Y2=0
cc_1151 N_A_3277_47#_c_1456_n N_VPWR_c_2027_n 0.0210596f $X=16.605 $Y=2.31 $X2=0
+ $Y2=0
cc_1152 N_A_3277_47#_c_1453_n N_Z_c_2373_n 0.00348752f $X=17.74 $Y=1.4 $X2=0
+ $Y2=0
cc_1153 N_A_3277_47#_c_1449_n N_Z_c_2373_n 0.0033343f $X=16.89 $Y=1.205 $X2=0
+ $Y2=0
cc_1154 N_A_3277_47#_M1024_g N_Z_c_2388_n 0.00753886f $X=17.36 $Y=2.075 $X2=0
+ $Y2=0
cc_1155 N_A_3277_47#_c_1448_n N_Z_c_2388_n 9.57301e-19 $X=17.45 $Y=1.4 $X2=0
+ $Y2=0
cc_1156 N_A_3277_47#_c_1456_n N_Z_c_2388_n 0.0308332f $X=16.605 $Y=2.31 $X2=0
+ $Y2=0
cc_1157 N_A_3277_47#_c_1451_n N_Z_c_2388_n 0.0132841f $X=16.89 $Y=1.42 $X2=0
+ $Y2=0
cc_1158 N_A_3277_47#_M1042_g N_Z_c_2389_n 0.00411531f $X=17.83 $Y=2.075 $X2=0
+ $Y2=0
cc_1159 N_A_3277_47#_M1042_g N_Z_c_2567_n 0.00513826f $X=17.83 $Y=2.075 $X2=0
+ $Y2=0
cc_1160 N_A_3277_47#_M1024_g N_Z_c_2568_n 0.00635536f $X=17.36 $Y=2.075 $X2=0
+ $Y2=0
cc_1161 N_A_3277_47#_c_1453_n N_Z_c_2568_n 8.37785e-19 $X=17.74 $Y=1.4 $X2=0
+ $Y2=0
cc_1162 N_A_3277_47#_M1042_g N_Z_c_2568_n 0.0105371f $X=17.83 $Y=2.075 $X2=0
+ $Y2=0
cc_1163 N_A_3277_47#_M1024_g N_Z_c_2381_n 0.00476154f $X=17.36 $Y=2.075 $X2=0
+ $Y2=0
cc_1164 N_A_3277_47#_c_1453_n N_Z_c_2381_n 0.0140509f $X=17.74 $Y=1.4 $X2=0
+ $Y2=0
cc_1165 N_A_3277_47#_c_1448_n N_Z_c_2381_n 7.26438e-19 $X=17.45 $Y=1.4 $X2=0
+ $Y2=0
cc_1166 N_A_3277_47#_M1042_g N_Z_c_2381_n 0.00268051f $X=17.83 $Y=2.075 $X2=0
+ $Y2=0
cc_1167 N_A_3277_47#_c_1449_n N_Z_c_2381_n 0.00967956f $X=16.89 $Y=1.205 $X2=0
+ $Y2=0
cc_1168 N_A_3277_47#_c_1451_n N_Z_c_2381_n 0.0117695f $X=16.89 $Y=1.42 $X2=0
+ $Y2=0
cc_1169 N_A_3277_47#_M1024_g N_A_3400_333#_c_3082_n 0.00745341f $X=17.36
+ $Y=2.075 $X2=0 $Y2=0
cc_1170 N_A_3277_47#_c_1448_n N_A_3400_333#_c_3082_n 0.00133381f $X=17.45 $Y=1.4
+ $X2=0 $Y2=0
cc_1171 N_A_3277_47#_c_1456_n N_A_3400_333#_c_3082_n 0.0347621f $X=16.605
+ $Y=2.31 $X2=0 $Y2=0
cc_1172 N_A_3277_47#_c_1451_n N_A_3400_333#_c_3082_n 0.0132748f $X=16.89 $Y=1.42
+ $X2=0 $Y2=0
cc_1173 N_A_3277_47#_M1024_g N_A_3400_333#_c_3090_n 0.00971609f $X=17.36
+ $Y=2.075 $X2=0 $Y2=0
cc_1174 N_A_3277_47#_M1042_g N_A_3400_333#_c_3090_n 0.0111338f $X=17.83 $Y=2.075
+ $X2=0 $Y2=0
cc_1175 N_A_3277_47#_c_1456_n N_A_3400_333#_c_3092_n 0.010563f $X=16.605 $Y=2.31
+ $X2=0 $Y2=0
cc_1176 N_A_3277_47#_M1042_g N_A_3400_333#_c_3093_n 0.00717732f $X=17.83
+ $Y=2.075 $X2=0 $Y2=0
cc_1177 N_A_3277_47#_M1042_g N_A_3400_333#_c_3094_n 0.00176121f $X=17.83
+ $Y=2.075 $X2=0 $Y2=0
cc_1178 N_A_3277_47#_M1050_d VGND 0.00250855f $X=16.385 $Y=0.235 $X2=0 $Y2=0
cc_1179 N_A_3277_47#_c_1450_n VGND 0.0186564f $X=16.52 $Y=0.495 $X2=0 $Y2=0
cc_1180 N_A_3277_47#_c_1450_n N_VGND_c_3317_n 0.0173492f $X=16.52 $Y=0.495 $X2=0
+ $Y2=0
cc_1181 N_A_3277_47#_c_1448_n N_A_3421_69#_c_3762_n 0.00308807f $X=17.45 $Y=1.4
+ $X2=0 $Y2=0
cc_1182 N_A_3277_47#_c_1449_n N_A_3421_69#_c_3762_n 0.00101918f $X=16.89
+ $Y=1.205 $X2=0 $Y2=0
cc_1183 N_A_3277_47#_c_1450_n N_A_3421_69#_c_3762_n 0.0185512f $X=16.52 $Y=0.495
+ $X2=0 $Y2=0
cc_1184 N_A_3277_47#_c_1451_n N_A_3421_69#_c_3762_n 0.00285813f $X=16.89 $Y=1.42
+ $X2=0 $Y2=0
cc_1185 N_A_3277_47#_c_1450_n N_A_3421_69#_c_3759_n 0.00358194f $X=16.52
+ $Y=0.495 $X2=0 $Y2=0
cc_1186 D[5] N_D[6]_c_1579_n 0.0231965f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_1187 N_D[5]_c_1527_n N_D[6]_c_1579_n 7.85936e-19 $X=18.91 $Y=1.16 $X2=0 $Y2=0
cc_1188 D[5] N_D[6]_c_1580_n 7.85936e-19 $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_1189 N_D[5]_c_1527_n N_D[6]_c_1580_n 0.00603597f $X=18.91 $Y=1.16 $X2=0 $Y2=0
cc_1190 N_D[5]_M1025_g N_VPWR_c_2009_n 0.00919666f $X=18.355 $Y=1.985 $X2=0
+ $Y2=0
cc_1191 N_D[5]_M1038_g N_VPWR_c_2009_n 0.0031734f $X=18.825 $Y=1.985 $X2=0 $Y2=0
cc_1192 N_D[5]_M1025_g N_VPWR_c_2165_n 0.00295119f $X=18.355 $Y=1.985 $X2=0
+ $Y2=0
cc_1193 N_D[5]_M1038_g N_VPWR_c_2165_n 0.00314707f $X=18.825 $Y=1.985 $X2=0
+ $Y2=0
cc_1194 N_D[5]_M1025_g VPWR 0.00588601f $X=18.355 $Y=1.985 $X2=0 $Y2=0
cc_1195 N_D[5]_M1038_g VPWR 0.00822554f $X=18.825 $Y=1.985 $X2=0 $Y2=0
cc_1196 N_D[5]_M1025_g N_VPWR_c_2027_n 0.00622633f $X=18.355 $Y=1.985 $X2=0
+ $Y2=0
cc_1197 N_D[5]_M1038_g N_VPWR_c_2028_n 0.00652917f $X=18.825 $Y=1.985 $X2=0
+ $Y2=0
cc_1198 N_D[5]_M1025_g N_Z_c_2389_n 0.00431834f $X=18.355 $Y=1.985 $X2=0 $Y2=0
cc_1199 N_D[5]_M1038_g N_Z_c_2389_n 0.00406261f $X=18.825 $Y=1.985 $X2=0 $Y2=0
cc_1200 D[5] N_Z_c_2389_n 0.00125914f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_1201 N_D[5]_M1025_g N_Z_c_2381_n 0.00112534f $X=18.355 $Y=1.985 $X2=0 $Y2=0
cc_1202 N_D[5]_M1047_g N_Z_c_2381_n 8.13311e-19 $X=18.38 $Y=0.56 $X2=0 $Y2=0
cc_1203 D[5] N_Z_c_2381_n 0.00742792f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_1204 N_D[5]_c_1527_n N_Z_c_2381_n 0.00583073f $X=18.91 $Y=1.16 $X2=0 $Y2=0
cc_1205 N_D[5]_M1025_g N_A_3400_333#_c_3093_n 0.00541465f $X=18.355 $Y=1.985
+ $X2=0 $Y2=0
cc_1206 N_D[5]_M1025_g N_A_3400_333#_c_3096_n 0.0127833f $X=18.355 $Y=1.985
+ $X2=0 $Y2=0
cc_1207 N_D[5]_M1038_g N_A_3400_333#_c_3096_n 0.0101085f $X=18.825 $Y=1.985
+ $X2=0 $Y2=0
cc_1208 D[5] N_A_3400_333#_c_3096_n 0.0323774f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_1209 N_D[5]_c_1527_n N_A_3400_333#_c_3096_n 7.13708e-19 $X=18.91 $Y=1.16
+ $X2=0 $Y2=0
cc_1210 D[5] N_A_3400_333#_c_3083_n 0.0226682f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_1211 N_D[5]_c_1527_n N_A_3400_333#_c_3083_n 9.6385e-19 $X=18.91 $Y=1.16 $X2=0
+ $Y2=0
cc_1212 N_D[5]_M1038_g N_A_3400_333#_c_3084_n 0.00325722f $X=18.825 $Y=1.985
+ $X2=0 $Y2=0
cc_1213 N_D[5]_M1047_g N_VGND_c_3299_n 0.00300333f $X=18.38 $Y=0.56 $X2=0 $Y2=0
cc_1214 N_D[5]_M1054_g N_VGND_c_3299_n 0.0030929f $X=18.8 $Y=0.56 $X2=0 $Y2=0
cc_1215 N_D[5]_M1054_g N_VGND_c_3300_n 0.00430643f $X=18.8 $Y=0.56 $X2=0 $Y2=0
cc_1216 N_D[5]_M1047_g VGND 0.00600262f $X=18.38 $Y=0.56 $X2=0 $Y2=0
cc_1217 N_D[5]_M1054_g VGND 0.00733187f $X=18.8 $Y=0.56 $X2=0 $Y2=0
cc_1218 N_D[5]_M1047_g N_VGND_c_3317_n 0.00436487f $X=18.38 $Y=0.56 $X2=0 $Y2=0
cc_1219 N_D[5]_M1047_g N_A_3421_69#_c_3760_n 0.0114493f $X=18.38 $Y=0.56 $X2=0
+ $Y2=0
cc_1220 N_D[5]_M1054_g N_A_3421_69#_c_3760_n 0.00931728f $X=18.8 $Y=0.56 $X2=0
+ $Y2=0
cc_1221 D[5] N_A_3421_69#_c_3760_n 0.0518587f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_1222 N_D[5]_c_1527_n N_A_3421_69#_c_3760_n 0.00665175f $X=18.91 $Y=1.16 $X2=0
+ $Y2=0
cc_1223 N_D[5]_M1047_g N_A_3421_69#_c_3761_n 0.00114614f $X=18.38 $Y=0.56 $X2=0
+ $Y2=0
cc_1224 N_D[5]_c_1527_n N_A_3421_69#_c_3761_n 0.00120541f $X=18.91 $Y=1.16 $X2=0
+ $Y2=0
cc_1225 N_D[5]_M1047_g N_A_3421_69#_c_3780_n 5.29024e-19 $X=18.38 $Y=0.56 $X2=0
+ $Y2=0
cc_1226 N_D[5]_M1054_g N_A_3421_69#_c_3780_n 0.00633603f $X=18.8 $Y=0.56 $X2=0
+ $Y2=0
cc_1227 N_D[6]_M1072_g N_A_4142_265#_M1033_g 0.0241475f $X=20.285 $Y=1.985 $X2=0
+ $Y2=0
cc_1228 N_D[6]_M1072_g N_A_4142_265#_c_1635_n 0.00671996f $X=20.285 $Y=1.985
+ $X2=0 $Y2=0
cc_1229 N_D[6]_M1079_g N_S[6]_c_1709_n 0.0165585f $X=20.26 $Y=0.56 $X2=0 $Y2=0
cc_1230 N_D[6]_M1029_g N_VPWR_c_2010_n 0.0031734f $X=19.815 $Y=1.985 $X2=0 $Y2=0
cc_1231 N_D[6]_M1072_g N_VPWR_c_2010_n 0.00919666f $X=20.285 $Y=1.985 $X2=0
+ $Y2=0
cc_1232 N_D[6]_M1029_g N_VPWR_c_2173_n 0.00314707f $X=19.815 $Y=1.985 $X2=0
+ $Y2=0
cc_1233 N_D[6]_M1072_g N_VPWR_c_2173_n 0.00295119f $X=20.285 $Y=1.985 $X2=0
+ $Y2=0
cc_1234 N_D[6]_M1072_g N_VPWR_c_2019_n 0.00622633f $X=20.285 $Y=1.985 $X2=0
+ $Y2=0
cc_1235 N_D[6]_M1029_g VPWR 0.00822554f $X=19.815 $Y=1.985 $X2=0 $Y2=0
cc_1236 N_D[6]_M1072_g VPWR 0.00588601f $X=20.285 $Y=1.985 $X2=0 $Y2=0
cc_1237 N_D[6]_M1029_g N_VPWR_c_2028_n 0.00652917f $X=19.815 $Y=1.985 $X2=0
+ $Y2=0
cc_1238 N_D[6]_M1029_g N_Z_c_2389_n 0.00406261f $X=19.815 $Y=1.985 $X2=0 $Y2=0
cc_1239 N_D[6]_M1072_g N_Z_c_2389_n 0.00431834f $X=20.285 $Y=1.985 $X2=0 $Y2=0
cc_1240 N_D[6]_c_1579_n N_Z_c_2389_n 0.00125914f $X=20.07 $Y=1.16 $X2=0 $Y2=0
cc_1241 N_D[6]_M1079_g N_Z_c_2382_n 8.13311e-19 $X=20.26 $Y=0.56 $X2=0 $Y2=0
cc_1242 N_D[6]_M1072_g N_Z_c_2382_n 0.00112534f $X=20.285 $Y=1.985 $X2=0 $Y2=0
cc_1243 N_D[6]_c_1579_n N_Z_c_2382_n 0.00742792f $X=20.07 $Y=1.16 $X2=0 $Y2=0
cc_1244 N_D[6]_c_1580_n N_Z_c_2382_n 0.00583073f $X=20.285 $Y=1.16 $X2=0 $Y2=0
cc_1245 N_D[6]_c_1579_n N_A_3891_297#_c_3141_n 0.0226682f $X=20.07 $Y=1.16 $X2=0
+ $Y2=0
cc_1246 N_D[6]_c_1580_n N_A_3891_297#_c_3141_n 9.6385e-19 $X=20.285 $Y=1.16
+ $X2=0 $Y2=0
cc_1247 N_D[6]_M1029_g N_A_3891_297#_c_3147_n 0.0101085f $X=19.815 $Y=1.985
+ $X2=0 $Y2=0
cc_1248 N_D[6]_M1072_g N_A_3891_297#_c_3147_n 0.0127833f $X=20.285 $Y=1.985
+ $X2=0 $Y2=0
cc_1249 N_D[6]_c_1579_n N_A_3891_297#_c_3147_n 0.0323774f $X=20.07 $Y=1.16 $X2=0
+ $Y2=0
cc_1250 N_D[6]_c_1580_n N_A_3891_297#_c_3147_n 7.13708e-19 $X=20.285 $Y=1.16
+ $X2=0 $Y2=0
cc_1251 N_D[6]_M1072_g N_A_3891_297#_c_3151_n 0.00541465f $X=20.285 $Y=1.985
+ $X2=0 $Y2=0
cc_1252 N_D[6]_M1029_g N_A_3891_297#_c_3143_n 0.00325722f $X=19.815 $Y=1.985
+ $X2=0 $Y2=0
cc_1253 N_D[6]_M1070_g N_VGND_c_3300_n 0.00430643f $X=19.84 $Y=0.56 $X2=0 $Y2=0
cc_1254 N_D[6]_M1070_g N_VGND_c_3301_n 0.0030929f $X=19.84 $Y=0.56 $X2=0 $Y2=0
cc_1255 N_D[6]_M1079_g N_VGND_c_3301_n 0.00300333f $X=20.26 $Y=0.56 $X2=0 $Y2=0
cc_1256 N_D[6]_M1079_g N_VGND_c_3310_n 0.00436487f $X=20.26 $Y=0.56 $X2=0 $Y2=0
cc_1257 N_D[6]_M1070_g VGND 0.00733187f $X=19.84 $Y=0.56 $X2=0 $Y2=0
cc_1258 N_D[6]_M1079_g VGND 0.00600262f $X=20.26 $Y=0.56 $X2=0 $Y2=0
cc_1259 N_D[6]_M1070_g N_A_3891_47#_c_3809_n 0.00633603f $X=19.84 $Y=0.56 $X2=0
+ $Y2=0
cc_1260 N_D[6]_M1079_g N_A_3891_47#_c_3809_n 5.29024e-19 $X=20.26 $Y=0.56 $X2=0
+ $Y2=0
cc_1261 N_D[6]_M1070_g N_A_3891_47#_c_3806_n 0.0084485f $X=19.84 $Y=0.56 $X2=0
+ $Y2=0
cc_1262 N_D[6]_M1079_g N_A_3891_47#_c_3806_n 0.0125955f $X=20.26 $Y=0.56 $X2=0
+ $Y2=0
cc_1263 N_D[6]_c_1579_n N_A_3891_47#_c_3806_n 0.0274027f $X=20.07 $Y=1.16 $X2=0
+ $Y2=0
cc_1264 N_D[6]_c_1580_n N_A_3891_47#_c_3806_n 0.00321151f $X=20.285 $Y=1.16
+ $X2=0 $Y2=0
cc_1265 N_D[6]_M1070_g N_A_3891_47#_c_3807_n 8.68782e-19 $X=19.84 $Y=0.56 $X2=0
+ $Y2=0
cc_1266 N_D[6]_c_1579_n N_A_3891_47#_c_3807_n 0.024456f $X=20.07 $Y=1.16 $X2=0
+ $Y2=0
cc_1267 N_D[6]_c_1580_n N_A_3891_47#_c_3807_n 0.00464565f $X=20.285 $Y=1.16
+ $X2=0 $Y2=0
cc_1268 N_A_4142_265#_c_1635_n N_S[6]_c_1707_n 0.00779314f $X=20.9 $Y=1.4
+ $X2=-0.19 $Y2=-0.24
cc_1269 N_A_4142_265#_c_1634_n N_S[6]_c_1710_n 0.00810157f $X=21.19 $Y=1.4 $X2=0
+ $Y2=0
cc_1270 N_A_4142_265#_c_1630_n N_S[6]_c_1710_n 7.04048e-19 $X=21.75 $Y=1.205
+ $X2=0 $Y2=0
cc_1271 N_A_4142_265#_c_1629_n N_S[6]_c_1712_n 0.0100587f $X=21.75 $Y=0.755
+ $X2=0 $Y2=0
cc_1272 N_A_4142_265#_c_1630_n N_S[6]_c_1712_n 0.00267287f $X=21.75 $Y=1.205
+ $X2=0 $Y2=0
cc_1273 N_A_4142_265#_c_1629_n N_S[6]_c_1713_n 0.0105766f $X=21.75 $Y=0.755
+ $X2=0 $Y2=0
cc_1274 N_A_4142_265#_c_1630_n N_S[6]_c_1713_n 0.0090765f $X=21.75 $Y=1.205
+ $X2=0 $Y2=0
cc_1275 N_A_4142_265#_c_1631_n N_S[6]_c_1713_n 0.00742826f $X=22.035 $Y=1.63
+ $X2=0 $Y2=0
cc_1276 N_A_4142_265#_c_1630_n N_S[6]_c_1714_n 0.00445422f $X=21.75 $Y=1.205
+ $X2=0 $Y2=0
cc_1277 N_A_4142_265#_c_1631_n N_S[6]_c_1714_n 4.25171e-19 $X=22.035 $Y=1.63
+ $X2=0 $Y2=0
cc_1278 N_A_4142_265#_c_1632_n N_S[6]_c_1714_n 0.00920672f $X=21.28 $Y=1.34
+ $X2=0 $Y2=0
cc_1279 N_A_4142_265#_c_1630_n N_S[6]_c_1715_n 0.00205356f $X=21.75 $Y=1.205
+ $X2=0 $Y2=0
cc_1280 N_A_4142_265#_c_1637_n N_S[6]_c_1715_n 0.00862444f $X=22.035 $Y=2.31
+ $X2=0 $Y2=0
cc_1281 N_A_4142_265#_c_1631_n N_S[6]_c_1715_n 0.00828481f $X=22.035 $Y=1.63
+ $X2=0 $Y2=0
cc_1282 N_A_4142_265#_c_1632_n N_S[6]_c_1715_n 0.00692516f $X=21.28 $Y=1.34
+ $X2=0 $Y2=0
cc_1283 N_A_4142_265#_c_1630_n N_S[6]_c_1716_n 0.00149517f $X=21.75 $Y=1.205
+ $X2=0 $Y2=0
cc_1284 N_A_4142_265#_c_1629_n S[6] 0.0061421f $X=21.75 $Y=0.755 $X2=0 $Y2=0
cc_1285 N_A_4142_265#_c_1630_n S[6] 0.0101733f $X=21.75 $Y=1.205 $X2=0 $Y2=0
cc_1286 N_A_4142_265#_c_1631_n S[6] 0.0127184f $X=22.035 $Y=1.63 $X2=0 $Y2=0
cc_1287 N_A_4142_265#_c_1632_n S[6] 3.07062e-19 $X=21.28 $Y=1.34 $X2=0 $Y2=0
cc_1288 N_A_4142_265#_M1033_g N_VPWR_c_2010_n 0.00107974f $X=20.81 $Y=2.075
+ $X2=0 $Y2=0
cc_1289 N_A_4142_265#_c_1637_n N_VPWR_c_2011_n 0.0321301f $X=22.035 $Y=2.31
+ $X2=0 $Y2=0
cc_1290 N_A_4142_265#_c_1631_n N_VPWR_c_2011_n 0.00732952f $X=22.035 $Y=1.63
+ $X2=0 $Y2=0
cc_1291 N_A_4142_265#_M1033_g N_VPWR_c_2019_n 0.00429453f $X=20.81 $Y=2.075
+ $X2=0 $Y2=0
cc_1292 N_A_4142_265#_M1046_g N_VPWR_c_2019_n 0.00429453f $X=21.28 $Y=2.075
+ $X2=0 $Y2=0
cc_1293 N_A_4142_265#_c_1637_n N_VPWR_c_2019_n 0.0210596f $X=22.035 $Y=2.31
+ $X2=0 $Y2=0
cc_1294 N_A_4142_265#_M1039_s VPWR 0.00179197f $X=21.91 $Y=1.485 $X2=0 $Y2=0
cc_1295 N_A_4142_265#_M1033_g VPWR 0.00615305f $X=20.81 $Y=2.075 $X2=0 $Y2=0
cc_1296 N_A_4142_265#_M1046_g VPWR 0.00728421f $X=21.28 $Y=2.075 $X2=0 $Y2=0
cc_1297 N_A_4142_265#_c_1637_n VPWR 0.00594162f $X=22.035 $Y=2.31 $X2=0 $Y2=0
cc_1298 N_A_4142_265#_c_1634_n N_Z_c_2374_n 0.00168443f $X=21.19 $Y=1.4 $X2=0
+ $Y2=0
cc_1299 N_A_4142_265#_c_1635_n N_Z_c_2374_n 0.00180308f $X=20.9 $Y=1.4 $X2=0
+ $Y2=0
cc_1300 N_A_4142_265#_c_1630_n N_Z_c_2374_n 0.0033343f $X=21.75 $Y=1.205 $X2=0
+ $Y2=0
cc_1301 N_A_4142_265#_M1033_g N_Z_c_2389_n 0.00411531f $X=20.81 $Y=2.075 $X2=0
+ $Y2=0
cc_1302 N_A_4142_265#_M1046_g N_Z_c_2390_n 0.00753886f $X=21.28 $Y=2.075 $X2=0
+ $Y2=0
cc_1303 N_A_4142_265#_c_1637_n N_Z_c_2390_n 0.0308332f $X=22.035 $Y=2.31 $X2=0
+ $Y2=0
cc_1304 N_A_4142_265#_c_1631_n N_Z_c_2390_n 0.0132841f $X=22.035 $Y=1.63 $X2=0
+ $Y2=0
cc_1305 N_A_4142_265#_c_1632_n N_Z_c_2390_n 9.57301e-19 $X=21.28 $Y=1.34 $X2=0
+ $Y2=0
cc_1306 N_A_4142_265#_M1033_g N_Z_c_2599_n 0.00513826f $X=20.81 $Y=2.075 $X2=0
+ $Y2=0
cc_1307 N_A_4142_265#_M1033_g N_Z_c_2600_n 0.0105371f $X=20.81 $Y=2.075 $X2=0
+ $Y2=0
cc_1308 N_A_4142_265#_c_1634_n N_Z_c_2600_n 8.37785e-19 $X=21.19 $Y=1.4 $X2=0
+ $Y2=0
cc_1309 N_A_4142_265#_M1046_g N_Z_c_2600_n 0.00635536f $X=21.28 $Y=2.075 $X2=0
+ $Y2=0
cc_1310 N_A_4142_265#_M1033_g N_Z_c_2382_n 0.00268051f $X=20.81 $Y=2.075 $X2=0
+ $Y2=0
cc_1311 N_A_4142_265#_c_1634_n N_Z_c_2382_n 0.0140509f $X=21.19 $Y=1.4 $X2=0
+ $Y2=0
cc_1312 N_A_4142_265#_M1046_g N_Z_c_2382_n 0.00476154f $X=21.28 $Y=2.075 $X2=0
+ $Y2=0
cc_1313 N_A_4142_265#_c_1630_n N_Z_c_2382_n 0.00967956f $X=21.75 $Y=1.205 $X2=0
+ $Y2=0
cc_1314 N_A_4142_265#_c_1631_n N_Z_c_2382_n 0.0117695f $X=22.035 $Y=1.63 $X2=0
+ $Y2=0
cc_1315 N_A_4142_265#_c_1632_n N_Z_c_2382_n 7.26438e-19 $X=21.28 $Y=1.34 $X2=0
+ $Y2=0
cc_1316 N_A_4142_265#_M1033_g N_A_3891_297#_c_3147_n 0.00176121f $X=20.81
+ $Y=2.075 $X2=0 $Y2=0
cc_1317 N_A_4142_265#_M1033_g N_A_3891_297#_c_3151_n 0.00717732f $X=20.81
+ $Y=2.075 $X2=0 $Y2=0
cc_1318 N_A_4142_265#_M1033_g N_A_3891_297#_c_3155_n 0.0111338f $X=20.81
+ $Y=2.075 $X2=0 $Y2=0
cc_1319 N_A_4142_265#_M1046_g N_A_3891_297#_c_3155_n 0.00971609f $X=21.28
+ $Y=2.075 $X2=0 $Y2=0
cc_1320 N_A_4142_265#_c_1637_n N_A_3891_297#_c_3155_n 0.010563f $X=22.035
+ $Y=2.31 $X2=0 $Y2=0
cc_1321 N_A_4142_265#_M1046_g N_A_3891_297#_c_3142_n 0.00745341f $X=21.28
+ $Y=2.075 $X2=0 $Y2=0
cc_1322 N_A_4142_265#_c_1637_n N_A_3891_297#_c_3142_n 0.0347621f $X=22.035
+ $Y=2.31 $X2=0 $Y2=0
cc_1323 N_A_4142_265#_c_1631_n N_A_3891_297#_c_3142_n 0.0132748f $X=22.035
+ $Y=1.63 $X2=0 $Y2=0
cc_1324 N_A_4142_265#_c_1632_n N_A_3891_297#_c_3142_n 0.00133381f $X=21.28
+ $Y=1.34 $X2=0 $Y2=0
cc_1325 N_A_4142_265#_c_1629_n N_VGND_c_3310_n 0.0173492f $X=21.75 $Y=0.755
+ $X2=0 $Y2=0
cc_1326 N_A_4142_265#_M1075_s VGND 0.00250855f $X=21.995 $Y=0.235 $X2=0 $Y2=0
cc_1327 N_A_4142_265#_c_1629_n VGND 0.0186564f $X=21.75 $Y=0.755 $X2=0 $Y2=0
cc_1328 N_A_4142_265#_c_1629_n N_A_3891_47#_c_3808_n 0.00358194f $X=21.75
+ $Y=0.755 $X2=0 $Y2=0
cc_1329 N_A_4142_265#_c_1629_n N_A_3891_47#_c_3819_n 0.0185512f $X=21.75
+ $Y=0.755 $X2=0 $Y2=0
cc_1330 N_A_4142_265#_c_1630_n N_A_3891_47#_c_3819_n 0.00101918f $X=21.75
+ $Y=1.205 $X2=0 $Y2=0
cc_1331 N_A_4142_265#_c_1631_n N_A_3891_47#_c_3819_n 0.00285813f $X=22.035
+ $Y=1.63 $X2=0 $Y2=0
cc_1332 N_A_4142_265#_c_1632_n N_A_3891_47#_c_3819_n 0.00308807f $X=21.28
+ $Y=1.34 $X2=0 $Y2=0
cc_1333 N_S[6]_c_1716_n N_S[7]_c_1772_n 0.0133556f $X=22.33 $Y=0.845 $X2=-0.19
+ $Y2=-0.24
cc_1334 N_S[6]_c_1715_n N_S[7]_c_1773_n 0.0418422f $X=22.27 $Y=1.41 $X2=0 $Y2=0
cc_1335 S[6] N_S[7]_c_1773_n 8.74983e-19 $X=22.225 $Y=1.105 $X2=0 $Y2=0
cc_1336 N_S[6]_c_1715_n S[7] 8.74983e-19 $X=22.27 $Y=1.41 $X2=0 $Y2=0
cc_1337 S[6] S[7] 0.0208489f $X=22.225 $Y=1.105 $X2=0 $Y2=0
cc_1338 N_S[6]_c_1715_n N_VPWR_c_2011_n 0.00456891f $X=22.27 $Y=1.41 $X2=0 $Y2=0
cc_1339 S[6] N_VPWR_c_2011_n 0.00569857f $X=22.225 $Y=1.105 $X2=0 $Y2=0
cc_1340 N_S[6]_c_1715_n N_VPWR_c_2019_n 0.00673617f $X=22.27 $Y=1.41 $X2=0 $Y2=0
cc_1341 N_S[6]_c_1715_n VPWR 0.00852379f $X=22.27 $Y=1.41 $X2=0 $Y2=0
cc_1342 N_S[6]_c_1707_n N_Z_c_2374_n 0.00413022f $X=20.78 $Y=0.255 $X2=0 $Y2=0
cc_1343 N_S[6]_c_1710_n N_Z_c_2374_n 0.00495983f $X=21.2 $Y=0.255 $X2=0 $Y2=0
cc_1344 N_S[6]_c_1712_n N_Z_c_2374_n 4.25992e-19 $X=21.685 $Y=0.845 $X2=0 $Y2=0
cc_1345 N_S[6]_c_1715_n N_Z_c_2390_n 0.00513674f $X=22.27 $Y=1.41 $X2=0 $Y2=0
cc_1346 S[6] N_Z_c_2390_n 0.00545567f $X=22.225 $Y=1.105 $X2=0 $Y2=0
cc_1347 N_S[6]_c_1707_n N_Z_c_2382_n 0.00199103f $X=20.78 $Y=0.255 $X2=0 $Y2=0
cc_1348 N_S[6]_c_1710_n N_Z_c_2382_n 0.00133607f $X=21.2 $Y=0.255 $X2=0 $Y2=0
cc_1349 N_S[6]_c_1716_n N_VGND_c_3302_n 0.00330937f $X=22.33 $Y=0.845 $X2=0
+ $Y2=0
cc_1350 N_S[6]_c_1709_n N_VGND_c_3310_n 0.0271255f $X=20.855 $Y=0.18 $X2=0 $Y2=0
cc_1351 N_S[6]_c_1716_n N_VGND_c_3310_n 0.00585385f $X=22.33 $Y=0.845 $X2=0
+ $Y2=0
cc_1352 N_S[6]_c_1708_n VGND 0.00642387f $X=21.125 $Y=0.18 $X2=0 $Y2=0
cc_1353 N_S[6]_c_1709_n VGND 0.00474746f $X=20.855 $Y=0.18 $X2=0 $Y2=0
cc_1354 N_S[6]_c_1711_n VGND 0.0193094f $X=21.61 $Y=0.18 $X2=0 $Y2=0
cc_1355 N_S[6]_c_1716_n VGND 0.0111218f $X=22.33 $Y=0.845 $X2=0 $Y2=0
cc_1356 N_S[6]_c_1717_n VGND 0.00366655f $X=21.2 $Y=0.18 $X2=0 $Y2=0
cc_1357 N_S[6]_c_1707_n N_A_3891_47#_c_3806_n 0.00139422f $X=20.78 $Y=0.255
+ $X2=0 $Y2=0
cc_1358 N_S[6]_c_1707_n N_A_3891_47#_c_3808_n 0.0132844f $X=20.78 $Y=0.255 $X2=0
+ $Y2=0
cc_1359 N_S[6]_c_1708_n N_A_3891_47#_c_3808_n 0.00211351f $X=21.125 $Y=0.18
+ $X2=0 $Y2=0
cc_1360 N_S[6]_c_1710_n N_A_3891_47#_c_3808_n 0.0126455f $X=21.2 $Y=0.255 $X2=0
+ $Y2=0
cc_1361 N_S[6]_c_1711_n N_A_3891_47#_c_3808_n 0.00436105f $X=21.61 $Y=0.18 $X2=0
+ $Y2=0
cc_1362 N_S[6]_c_1712_n N_A_3891_47#_c_3808_n 0.00349455f $X=21.685 $Y=0.845
+ $X2=0 $Y2=0
cc_1363 N_S[6]_c_1712_n N_A_3891_47#_c_3819_n 0.00295202f $X=21.685 $Y=0.845
+ $X2=0 $Y2=0
cc_1364 N_S[7]_c_1780_n N_A_4565_47#_c_1839_n 0.00779314f $X=24.3 $Y=0.255 $X2=0
+ $Y2=0
cc_1365 N_S[7]_c_1773_n N_A_4565_47#_c_1834_n 0.00692516f $X=22.81 $Y=1.41 $X2=0
+ $Y2=0
cc_1366 N_S[7]_c_1774_n N_A_4565_47#_c_1834_n 0.00920672f $X=23.32 $Y=0.92 $X2=0
+ $Y2=0
cc_1367 N_S[7]_c_1778_n N_A_4565_47#_c_1834_n 0.00810157f $X=23.88 $Y=0.255
+ $X2=0 $Y2=0
cc_1368 S[7] N_A_4565_47#_c_1834_n 3.07062e-19 $X=22.685 $Y=1.105 $X2=0 $Y2=0
cc_1369 N_S[7]_c_1773_n N_A_4565_47#_c_1842_n 0.00862444f $X=22.81 $Y=1.41 $X2=0
+ $Y2=0
cc_1370 N_S[7]_c_1772_n N_A_4565_47#_c_1835_n 0.00149517f $X=22.75 $Y=0.845
+ $X2=0 $Y2=0
cc_1371 N_S[7]_c_1773_n N_A_4565_47#_c_1835_n 0.00205356f $X=22.81 $Y=1.41 $X2=0
+ $Y2=0
cc_1372 N_S[7]_c_1774_n N_A_4565_47#_c_1835_n 0.0135307f $X=23.32 $Y=0.92 $X2=0
+ $Y2=0
cc_1373 N_S[7]_c_1775_n N_A_4565_47#_c_1835_n 0.00267287f $X=23.395 $Y=0.845
+ $X2=0 $Y2=0
cc_1374 N_S[7]_c_1778_n N_A_4565_47#_c_1835_n 7.04048e-19 $X=23.88 $Y=0.255
+ $X2=0 $Y2=0
cc_1375 S[7] N_A_4565_47#_c_1835_n 0.0101733f $X=22.685 $Y=1.105 $X2=0 $Y2=0
cc_1376 N_S[7]_c_1773_n N_A_4565_47#_c_1836_n 0.0105766f $X=22.81 $Y=1.41 $X2=0
+ $Y2=0
cc_1377 N_S[7]_c_1775_n N_A_4565_47#_c_1836_n 0.0100587f $X=23.395 $Y=0.845
+ $X2=0 $Y2=0
cc_1378 S[7] N_A_4565_47#_c_1836_n 0.0061421f $X=22.685 $Y=1.105 $X2=0 $Y2=0
cc_1379 N_S[7]_c_1773_n N_A_4565_47#_c_1837_n 0.00828481f $X=22.81 $Y=1.41 $X2=0
+ $Y2=0
cc_1380 N_S[7]_c_1774_n N_A_4565_47#_c_1837_n 0.00785343f $X=23.32 $Y=0.92 $X2=0
+ $Y2=0
cc_1381 S[7] N_A_4565_47#_c_1837_n 0.0127184f $X=22.685 $Y=1.105 $X2=0 $Y2=0
cc_1382 N_S[7]_c_1779_n N_D[7]_M1011_g 0.0165585f $X=24.225 $Y=0.18 $X2=0 $Y2=0
cc_1383 N_S[7]_c_1773_n N_VPWR_c_2011_n 0.00456891f $X=22.81 $Y=1.41 $X2=0 $Y2=0
cc_1384 S[7] N_VPWR_c_2011_n 0.00569857f $X=22.685 $Y=1.105 $X2=0 $Y2=0
cc_1385 N_S[7]_c_1773_n VPWR 0.00852379f $X=22.81 $Y=1.41 $X2=0 $Y2=0
cc_1386 N_S[7]_c_1773_n N_VPWR_c_2029_n 0.00673617f $X=22.81 $Y=1.41 $X2=0 $Y2=0
cc_1387 N_S[7]_c_1775_n N_Z_c_2375_n 4.25992e-19 $X=23.395 $Y=0.845 $X2=0 $Y2=0
cc_1388 N_S[7]_c_1778_n N_Z_c_2375_n 0.00495983f $X=23.88 $Y=0.255 $X2=0 $Y2=0
cc_1389 N_S[7]_c_1780_n N_Z_c_2375_n 0.00413022f $X=24.3 $Y=0.255 $X2=0 $Y2=0
cc_1390 N_S[7]_c_1773_n N_Z_c_2390_n 0.00513674f $X=22.81 $Y=1.41 $X2=0 $Y2=0
cc_1391 S[7] N_Z_c_2390_n 0.00545567f $X=22.685 $Y=1.105 $X2=0 $Y2=0
cc_1392 N_S[7]_c_1778_n N_Z_c_2383_n 0.00133607f $X=23.88 $Y=0.255 $X2=0 $Y2=0
cc_1393 N_S[7]_c_1780_n N_Z_c_2383_n 0.00199103f $X=24.3 $Y=0.255 $X2=0 $Y2=0
cc_1394 N_S[7]_c_1772_n N_VGND_c_3302_n 0.00330937f $X=22.75 $Y=0.845 $X2=0
+ $Y2=0
cc_1395 N_S[7]_c_1772_n N_VGND_c_3312_n 0.00585385f $X=22.75 $Y=0.845 $X2=0
+ $Y2=0
cc_1396 N_S[7]_c_1777_n N_VGND_c_3312_n 0.0271255f $X=23.47 $Y=0.18 $X2=0 $Y2=0
cc_1397 N_S[7]_c_1772_n VGND 0.0111218f $X=22.75 $Y=0.845 $X2=0 $Y2=0
cc_1398 N_S[7]_c_1776_n VGND 0.0119932f $X=23.805 $Y=0.18 $X2=0 $Y2=0
cc_1399 N_S[7]_c_1777_n VGND 0.00731624f $X=23.47 $Y=0.18 $X2=0 $Y2=0
cc_1400 N_S[7]_c_1779_n VGND 0.0111713f $X=24.225 $Y=0.18 $X2=0 $Y2=0
cc_1401 N_S[7]_c_1781_n VGND 0.00366655f $X=23.88 $Y=0.18 $X2=0 $Y2=0
cc_1402 N_S[7]_c_1775_n N_A_4709_69#_c_3854_n 0.00295202f $X=23.395 $Y=0.845
+ $X2=0 $Y2=0
cc_1403 N_S[7]_c_1778_n N_A_4709_69#_c_3850_n 0.0126455f $X=23.88 $Y=0.255 $X2=0
+ $Y2=0
cc_1404 N_S[7]_c_1779_n N_A_4709_69#_c_3850_n 0.00211351f $X=24.225 $Y=0.18
+ $X2=0 $Y2=0
cc_1405 N_S[7]_c_1780_n N_A_4709_69#_c_3850_n 0.0132844f $X=24.3 $Y=0.255 $X2=0
+ $Y2=0
cc_1406 N_S[7]_c_1775_n N_A_4709_69#_c_3851_n 0.00349455f $X=23.395 $Y=0.845
+ $X2=0 $Y2=0
cc_1407 N_S[7]_c_1776_n N_A_4709_69#_c_3851_n 0.00436105f $X=23.805 $Y=0.18
+ $X2=0 $Y2=0
cc_1408 N_S[7]_c_1780_n N_A_4709_69#_c_3853_n 0.00139422f $X=24.3 $Y=0.255 $X2=0
+ $Y2=0
cc_1409 N_A_4565_47#_c_1839_n N_D[7]_M1030_g 0.00671996f $X=24.18 $Y=1.4 $X2=0
+ $Y2=0
cc_1410 N_A_4565_47#_M1073_g N_D[7]_M1030_g 0.0232231f $X=24.27 $Y=2.075 $X2=0
+ $Y2=0
cc_1411 N_A_4565_47#_c_1842_n N_VPWR_c_2011_n 0.0321301f $X=23.045 $Y=2.31 $X2=0
+ $Y2=0
cc_1412 N_A_4565_47#_c_1837_n N_VPWR_c_2011_n 0.00732952f $X=23.33 $Y=1.42 $X2=0
+ $Y2=0
cc_1413 N_A_4565_47#_M1073_g N_VPWR_c_2012_n 0.00107974f $X=24.27 $Y=2.075 $X2=0
+ $Y2=0
cc_1414 N_A_4565_47#_M1066_d VPWR 0.00179197f $X=22.9 $Y=1.485 $X2=0 $Y2=0
cc_1415 N_A_4565_47#_M1064_g VPWR 0.00728421f $X=23.8 $Y=2.075 $X2=0 $Y2=0
cc_1416 N_A_4565_47#_M1073_g VPWR 0.00617598f $X=24.27 $Y=2.075 $X2=0 $Y2=0
cc_1417 N_A_4565_47#_c_1842_n VPWR 0.00594162f $X=23.045 $Y=2.31 $X2=0 $Y2=0
cc_1418 N_A_4565_47#_M1064_g N_VPWR_c_2029_n 0.00429453f $X=23.8 $Y=2.075 $X2=0
+ $Y2=0
cc_1419 N_A_4565_47#_M1073_g N_VPWR_c_2029_n 0.00429453f $X=24.27 $Y=2.075 $X2=0
+ $Y2=0
cc_1420 N_A_4565_47#_c_1842_n N_VPWR_c_2029_n 0.0210596f $X=23.045 $Y=2.31 $X2=0
+ $Y2=0
cc_1421 N_A_4565_47#_c_1839_n N_Z_c_2375_n 0.00348752f $X=24.18 $Y=1.4 $X2=0
+ $Y2=0
cc_1422 N_A_4565_47#_c_1835_n N_Z_c_2375_n 0.0033343f $X=23.33 $Y=1.205 $X2=0
+ $Y2=0
cc_1423 N_A_4565_47#_M1064_g N_Z_c_2390_n 0.00753886f $X=23.8 $Y=2.075 $X2=0
+ $Y2=0
cc_1424 N_A_4565_47#_c_1834_n N_Z_c_2390_n 9.57301e-19 $X=23.89 $Y=1.4 $X2=0
+ $Y2=0
cc_1425 N_A_4565_47#_c_1842_n N_Z_c_2390_n 0.0308332f $X=23.045 $Y=2.31 $X2=0
+ $Y2=0
cc_1426 N_A_4565_47#_c_1837_n N_Z_c_2390_n 0.0132841f $X=23.33 $Y=1.42 $X2=0
+ $Y2=0
cc_1427 N_A_4565_47#_M1073_g Z 0.00635853f $X=24.27 $Y=2.075 $X2=0 $Y2=0
cc_1428 N_A_4565_47#_M1064_g N_Z_c_2630_n 0.00635536f $X=23.8 $Y=2.075 $X2=0
+ $Y2=0
cc_1429 N_A_4565_47#_c_1839_n N_Z_c_2630_n 8.37785e-19 $X=24.18 $Y=1.4 $X2=0
+ $Y2=0
cc_1430 N_A_4565_47#_M1073_g N_Z_c_2630_n 0.0105371f $X=24.27 $Y=2.075 $X2=0
+ $Y2=0
cc_1431 N_A_4565_47#_M1064_g N_Z_c_2383_n 0.00476154f $X=23.8 $Y=2.075 $X2=0
+ $Y2=0
cc_1432 N_A_4565_47#_c_1839_n N_Z_c_2383_n 0.0140509f $X=24.18 $Y=1.4 $X2=0
+ $Y2=0
cc_1433 N_A_4565_47#_c_1834_n N_Z_c_2383_n 7.26438e-19 $X=23.89 $Y=1.4 $X2=0
+ $Y2=0
cc_1434 N_A_4565_47#_M1073_g N_Z_c_2383_n 0.00268051f $X=24.27 $Y=2.075 $X2=0
+ $Y2=0
cc_1435 N_A_4565_47#_c_1835_n N_Z_c_2383_n 0.00967956f $X=23.33 $Y=1.205 $X2=0
+ $Y2=0
cc_1436 N_A_4565_47#_c_1837_n N_Z_c_2383_n 0.0117695f $X=23.33 $Y=1.42 $X2=0
+ $Y2=0
cc_1437 N_A_4565_47#_M1064_g N_A_4688_333#_c_3198_n 0.00745341f $X=23.8 $Y=2.075
+ $X2=0 $Y2=0
cc_1438 N_A_4565_47#_c_1834_n N_A_4688_333#_c_3198_n 0.00133381f $X=23.89 $Y=1.4
+ $X2=0 $Y2=0
cc_1439 N_A_4565_47#_c_1842_n N_A_4688_333#_c_3198_n 0.0347621f $X=23.045
+ $Y=2.31 $X2=0 $Y2=0
cc_1440 N_A_4565_47#_c_1837_n N_A_4688_333#_c_3198_n 0.0132748f $X=23.33 $Y=1.42
+ $X2=0 $Y2=0
cc_1441 N_A_4565_47#_M1064_g N_A_4688_333#_c_3206_n 0.00971609f $X=23.8 $Y=2.075
+ $X2=0 $Y2=0
cc_1442 N_A_4565_47#_M1073_g N_A_4688_333#_c_3206_n 0.0128147f $X=24.27 $Y=2.075
+ $X2=0 $Y2=0
cc_1443 N_A_4565_47#_c_1842_n N_A_4688_333#_c_3208_n 0.010563f $X=23.045 $Y=2.31
+ $X2=0 $Y2=0
cc_1444 N_A_4565_47#_M1073_g N_A_4688_333#_c_3209_n 0.00736707f $X=24.27
+ $Y=2.075 $X2=0 $Y2=0
cc_1445 N_A_4565_47#_M1073_g N_A_4688_333#_c_3210_n 0.00176121f $X=24.27
+ $Y=2.075 $X2=0 $Y2=0
cc_1446 N_A_4565_47#_c_1836_n N_VGND_c_3312_n 0.0173492f $X=22.96 $Y=0.495 $X2=0
+ $Y2=0
cc_1447 N_A_4565_47#_M1007_d VGND 0.00250855f $X=22.825 $Y=0.235 $X2=0 $Y2=0
cc_1448 N_A_4565_47#_c_1836_n VGND 0.0186564f $X=22.96 $Y=0.495 $X2=0 $Y2=0
cc_1449 N_A_4565_47#_c_1834_n N_A_4709_69#_c_3854_n 0.00308807f $X=23.89 $Y=1.4
+ $X2=0 $Y2=0
cc_1450 N_A_4565_47#_c_1835_n N_A_4709_69#_c_3854_n 0.00101918f $X=23.33
+ $Y=1.205 $X2=0 $Y2=0
cc_1451 N_A_4565_47#_c_1836_n N_A_4709_69#_c_3854_n 0.0185512f $X=22.96 $Y=0.495
+ $X2=0 $Y2=0
cc_1452 N_A_4565_47#_c_1837_n N_A_4709_69#_c_3854_n 0.00285813f $X=23.33 $Y=1.42
+ $X2=0 $Y2=0
cc_1453 N_A_4565_47#_c_1836_n N_A_4709_69#_c_3851_n 0.00358194f $X=22.96
+ $Y=0.495 $X2=0 $Y2=0
cc_1454 N_D[7]_M1030_g N_VPWR_c_2012_n 0.00919666f $X=24.795 $Y=1.985 $X2=0
+ $Y2=0
cc_1455 N_D[7]_M1069_g N_VPWR_c_2012_n 0.0031734f $X=25.265 $Y=1.985 $X2=0 $Y2=0
cc_1456 N_D[7]_M1030_g N_VPWR_c_2209_n 0.00343746f $X=24.795 $Y=1.985 $X2=0
+ $Y2=0
cc_1457 N_D[7]_M1069_g N_VPWR_c_2209_n 0.00363183f $X=25.265 $Y=1.985 $X2=0
+ $Y2=0
cc_1458 N_D[7]_M1030_g VPWR 0.0105515f $X=24.795 $Y=1.985 $X2=0 $Y2=0
cc_1459 N_D[7]_M1069_g VPWR 0.0120316f $X=25.265 $Y=1.985 $X2=0 $Y2=0
cc_1460 N_D[7]_M1030_g N_VPWR_c_2029_n 0.00622633f $X=24.795 $Y=1.985 $X2=0
+ $Y2=0
cc_1461 N_D[7]_M1069_g N_VPWR_c_2030_n 0.00652917f $X=25.265 $Y=1.985 $X2=0
+ $Y2=0
cc_1462 N_D[7]_M1030_g N_Z_c_2383_n 0.00112534f $X=24.795 $Y=1.985 $X2=0 $Y2=0
cc_1463 N_D[7]_M1011_g N_Z_c_2383_n 8.13311e-19 $X=24.82 $Y=0.56 $X2=0 $Y2=0
cc_1464 D[7] N_Z_c_2383_n 0.00742792f $X=25.445 $Y=1.105 $X2=0 $Y2=0
cc_1465 N_D[7]_c_1912_n N_Z_c_2383_n 0.00583073f $X=25.35 $Y=1.16 $X2=0 $Y2=0
cc_1466 N_D[7]_M1030_g N_A_4688_333#_c_3209_n 0.00557487f $X=24.795 $Y=1.985
+ $X2=0 $Y2=0
cc_1467 N_D[7]_M1030_g N_A_4688_333#_c_3212_n 0.0174487f $X=24.795 $Y=1.985
+ $X2=0 $Y2=0
cc_1468 N_D[7]_M1069_g N_A_4688_333#_c_3212_n 0.0142998f $X=25.265 $Y=1.985
+ $X2=0 $Y2=0
cc_1469 D[7] N_A_4688_333#_c_3212_n 0.0339353f $X=25.445 $Y=1.105 $X2=0 $Y2=0
cc_1470 N_D[7]_c_1912_n N_A_4688_333#_c_3212_n 7.13708e-19 $X=25.35 $Y=1.16
+ $X2=0 $Y2=0
cc_1471 D[7] N_A_4688_333#_c_3199_n 0.0235932f $X=25.445 $Y=1.105 $X2=0 $Y2=0
cc_1472 N_D[7]_c_1912_n N_A_4688_333#_c_3199_n 9.6385e-19 $X=25.35 $Y=1.16 $X2=0
+ $Y2=0
cc_1473 N_D[7]_M1069_g N_A_4688_333#_c_3200_n 0.00329008f $X=25.265 $Y=1.985
+ $X2=0 $Y2=0
cc_1474 N_D[7]_M1011_g N_VGND_c_3303_n 0.00300333f $X=24.82 $Y=0.56 $X2=0 $Y2=0
cc_1475 N_D[7]_M1027_g N_VGND_c_3303_n 0.0030929f $X=25.24 $Y=0.56 $X2=0 $Y2=0
cc_1476 N_D[7]_M1011_g N_VGND_c_3312_n 0.00436487f $X=24.82 $Y=0.56 $X2=0 $Y2=0
cc_1477 N_D[7]_M1011_g VGND 0.00600262f $X=24.82 $Y=0.56 $X2=0 $Y2=0
cc_1478 N_D[7]_M1027_g VGND 0.00697949f $X=25.24 $Y=0.56 $X2=0 $Y2=0
cc_1479 N_D[7]_M1027_g N_VGND_c_3318_n 0.00430643f $X=25.24 $Y=0.56 $X2=0 $Y2=0
cc_1480 N_D[7]_M1011_g N_A_4709_69#_c_3852_n 0.0114493f $X=24.82 $Y=0.56 $X2=0
+ $Y2=0
cc_1481 N_D[7]_M1027_g N_A_4709_69#_c_3852_n 0.00931728f $X=25.24 $Y=0.56 $X2=0
+ $Y2=0
cc_1482 D[7] N_A_4709_69#_c_3852_n 0.0518587f $X=25.445 $Y=1.105 $X2=0 $Y2=0
cc_1483 N_D[7]_c_1912_n N_A_4709_69#_c_3852_n 0.00665175f $X=25.35 $Y=1.16 $X2=0
+ $Y2=0
cc_1484 N_D[7]_M1011_g N_A_4709_69#_c_3853_n 0.00114614f $X=24.82 $Y=0.56 $X2=0
+ $Y2=0
cc_1485 N_D[7]_c_1912_n N_A_4709_69#_c_3853_n 0.00120541f $X=25.35 $Y=1.16 $X2=0
+ $Y2=0
cc_1486 N_D[7]_M1011_g N_A_4709_69#_c_3872_n 5.29024e-19 $X=24.82 $Y=0.56 $X2=0
+ $Y2=0
cc_1487 N_D[7]_M1027_g N_A_4709_69#_c_3872_n 0.00633603f $X=25.24 $Y=0.56 $X2=0
+ $Y2=0
cc_1488 N_A_27_297#_c_1959_n N_VPWR_M1003_s 0.00350459f $X=1.115 $Y=1.58
+ $X2=-0.19 $Y2=1.305
cc_1489 N_A_27_297#_c_1975_p N_VPWR_c_2001_n 0.0114322f $X=1.285 $Y=2.38 $X2=0
+ $Y2=0
cc_1490 N_A_27_297#_c_1959_n N_VPWR_c_2041_n 0.0170301f $X=1.115 $Y=1.58 $X2=0
+ $Y2=0
cc_1491 N_A_27_297#_c_1963_n N_VPWR_c_2041_n 0.0272234f $X=1.2 $Y=1.78 $X2=0
+ $Y2=0
cc_1492 N_A_27_297#_c_1967_n N_VPWR_c_2013_n 0.0569572f $X=2.11 $Y=2.38 $X2=0
+ $Y2=0
cc_1493 N_A_27_297#_c_1975_p N_VPWR_c_2013_n 0.0119545f $X=1.285 $Y=2.38 $X2=0
+ $Y2=0
cc_1494 N_A_27_297#_M1003_d VPWR 0.00217517f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_1495 N_A_27_297#_M1034_d VPWR 0.00481062f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_1496 N_A_27_297#_M1013_d VPWR 0.00210318f $X=2.05 $Y=1.665 $X2=0 $Y2=0
cc_1497 N_A_27_297#_c_1967_n VPWR 0.0196248f $X=2.11 $Y=2.38 $X2=0 $Y2=0
cc_1498 N_A_27_297#_c_1975_p VPWR 0.006547f $X=1.285 $Y=2.38 $X2=0 $Y2=0
cc_1499 N_A_27_297#_c_1955_n VPWR 0.0124483f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_1500 N_A_27_297#_c_1955_n N_VPWR_c_2022_n 0.020978f $X=0.26 $Y=2.34 $X2=0
+ $Y2=0
cc_1501 N_A_27_297#_c_1967_n N_Z_M1006_s 0.00341588f $X=2.11 $Y=2.38 $X2=0 $Y2=0
cc_1502 N_A_27_297#_M1013_d N_Z_c_2384_n 0.00237684f $X=2.05 $Y=1.665 $X2=0
+ $Y2=0
cc_1503 N_A_27_297#_c_1967_n N_Z_c_2384_n 0.00494997f $X=2.11 $Y=2.38 $X2=0
+ $Y2=0
cc_1504 N_A_27_297#_c_1954_n N_Z_c_2384_n 0.0132602f $X=2.195 $Y=1.81 $X2=0
+ $Y2=0
cc_1505 N_A_27_297#_c_1963_n N_Z_c_2410_n 0.0062686f $X=1.2 $Y=1.78 $X2=0 $Y2=0
cc_1506 N_A_27_297#_c_1967_n N_Z_c_2410_n 8.66896e-19 $X=2.11 $Y=2.38 $X2=0
+ $Y2=0
cc_1507 N_A_27_297#_c_1954_n N_Z_c_2410_n 4.86317e-19 $X=2.195 $Y=1.81 $X2=0
+ $Y2=0
cc_1508 N_A_27_297#_c_1963_n N_Z_c_2411_n 0.0235305f $X=1.2 $Y=1.78 $X2=0 $Y2=0
cc_1509 N_A_27_297#_c_1967_n N_Z_c_2411_n 0.0211175f $X=2.11 $Y=2.38 $X2=0 $Y2=0
cc_1510 N_A_27_297#_c_1954_n N_Z_c_2411_n 0.0212802f $X=2.195 $Y=1.81 $X2=0
+ $Y2=0
cc_1511 N_A_27_297#_c_1959_n N_Z_c_2376_n 0.00930189f $X=1.115 $Y=1.58 $X2=0
+ $Y2=0
cc_1512 N_A_27_297#_c_1954_n N_Z_c_2376_n 0.00468052f $X=2.195 $Y=1.81 $X2=0
+ $Y2=0
cc_1513 N_A_27_297#_c_1959_n N_A_27_47#_c_3247_n 0.0110288f $X=1.115 $Y=1.58
+ $X2=0 $Y2=0
cc_1514 VPWR N_Z_M1006_s 0.00187512f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1515 VPWR N_Z_M1040_s 0.00187512f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1516 VPWR N_Z_M1004_d 0.00187512f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1517 VPWR N_Z_M1005_d 0.00187512f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1518 VPWR N_Z_M1016_s 0.00187512f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1519 VPWR N_Z_M1024_s 0.00187512f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1520 VPWR N_Z_M1033_s 0.00187512f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1521 VPWR N_Z_M1064_s 0.00187512f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1522 N_VPWR_M1008_d N_Z_c_2384_n 5.82057e-19 $X=3.04 $Y=1.485 $X2=0 $Y2=0
cc_1523 N_VPWR_c_2002_n N_Z_c_2384_n 0.0287846f $X=3.22 $Y=1.63 $X2=0 $Y2=0
cc_1524 VPWR N_Z_c_2384_n 0.138617f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1525 VPWR N_Z_c_2410_n 0.0144354f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1526 N_VPWR_M1022_s N_Z_c_2385_n 0.00219731f $X=5.565 $Y=1.485 $X2=0 $Y2=0
cc_1527 N_VPWR_M1000_d N_Z_c_2385_n 0.00219731f $X=7.025 $Y=1.485 $X2=0 $Y2=0
cc_1528 N_VPWR_c_2077_n N_Z_c_2385_n 0.0159439f $X=5.71 $Y=1.94 $X2=0 $Y2=0
cc_1529 N_VPWR_c_2085_n N_Z_c_2385_n 0.0159439f $X=7.17 $Y=1.94 $X2=0 $Y2=0
cc_1530 VPWR N_Z_c_2385_n 0.136626f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1531 VPWR N_Z_c_2441_n 0.0144354f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1532 N_VPWR_M1067_d N_Z_c_2386_n 5.82057e-19 $X=9.48 $Y=1.485 $X2=0 $Y2=0
cc_1533 N_VPWR_c_2005_n N_Z_c_2386_n 0.0287846f $X=9.66 $Y=1.63 $X2=0 $Y2=0
cc_1534 VPWR N_Z_c_2386_n 0.138617f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1535 VPWR N_Z_c_2473_n 0.0144354f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1536 N_VPWR_M1001_d N_Z_c_2387_n 0.00219731f $X=12.005 $Y=1.485 $X2=0 $Y2=0
cc_1537 N_VPWR_M1014_s N_Z_c_2387_n 0.00219731f $X=13.465 $Y=1.485 $X2=0 $Y2=0
cc_1538 N_VPWR_c_2121_n N_Z_c_2387_n 0.0159439f $X=12.15 $Y=1.94 $X2=0 $Y2=0
cc_1539 N_VPWR_c_2129_n N_Z_c_2387_n 0.0159439f $X=13.61 $Y=1.94 $X2=0 $Y2=0
cc_1540 VPWR N_Z_c_2387_n 0.136626f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1541 VPWR N_Z_c_2504_n 0.0144354f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1542 N_VPWR_M1002_d N_Z_c_2388_n 5.82057e-19 $X=15.92 $Y=1.485 $X2=0 $Y2=0
cc_1543 N_VPWR_c_2008_n N_Z_c_2388_n 0.0287846f $X=16.1 $Y=1.63 $X2=0 $Y2=0
cc_1544 VPWR N_Z_c_2388_n 0.138617f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1545 VPWR N_Z_c_2536_n 0.0144354f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1546 N_VPWR_M1025_s N_Z_c_2389_n 0.00219731f $X=18.445 $Y=1.485 $X2=0 $Y2=0
cc_1547 N_VPWR_M1029_s N_Z_c_2389_n 0.00219731f $X=19.905 $Y=1.485 $X2=0 $Y2=0
cc_1548 N_VPWR_c_2165_n N_Z_c_2389_n 0.0159439f $X=18.59 $Y=1.94 $X2=0 $Y2=0
cc_1549 N_VPWR_c_2173_n N_Z_c_2389_n 0.0159439f $X=20.05 $Y=1.94 $X2=0 $Y2=0
cc_1550 VPWR N_Z_c_2389_n 0.136626f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1551 VPWR N_Z_c_2567_n 0.0144354f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1552 N_VPWR_M1039_d N_Z_c_2390_n 5.82057e-19 $X=22.36 $Y=1.485 $X2=0 $Y2=0
cc_1553 N_VPWR_c_2011_n N_Z_c_2390_n 0.0287846f $X=22.54 $Y=1.63 $X2=0 $Y2=0
cc_1554 VPWR N_Z_c_2390_n 0.138617f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1555 VPWR N_Z_c_2599_n 0.0144354f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1556 VPWR Z 0.0144354f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1557 VPWR N_A_824_333#_M1040_d 0.00210318f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=-0.24
cc_1558 VPWR N_A_824_333#_M1056_d 0.00273129f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1559 VPWR N_A_824_333#_M1049_d 0.00179197f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1560 N_VPWR_c_2003_n N_A_824_333#_c_2858_n 0.0114322f $X=5.71 $Y=2.34 $X2=0
+ $Y2=0
cc_1561 VPWR N_A_824_333#_c_2858_n 0.0161639f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1562 N_VPWR_c_2023_n N_A_824_333#_c_2858_n 0.0570268f $X=5.545 $Y=2.72 $X2=0
+ $Y2=0
cc_1563 VPWR N_A_824_333#_c_2860_n 0.0031082f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1564 N_VPWR_c_2023_n N_A_824_333#_c_2860_n 0.0118848f $X=5.545 $Y=2.72 $X2=0
+ $Y2=0
cc_1565 N_VPWR_c_2077_n N_A_824_333#_c_2861_n 0.0265477f $X=5.71 $Y=1.94 $X2=0
+ $Y2=0
cc_1566 N_VPWR_M1022_s N_A_824_333#_c_2864_n 0.00331615f $X=5.565 $Y=1.485 $X2=0
+ $Y2=0
cc_1567 N_VPWR_c_2077_n N_A_824_333#_c_2864_n 0.0158304f $X=5.71 $Y=1.94 $X2=0
+ $Y2=0
cc_1568 VPWR N_A_824_333#_c_2852_n 0.00591741f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1569 N_VPWR_c_2024_n N_A_824_333#_c_2852_n 0.020978f $X=7.035 $Y=2.72 $X2=0
+ $Y2=0
cc_1570 N_VPWR_c_2077_n N_A_824_333#_c_2853_n 0.0115021f $X=5.71 $Y=1.94 $X2=0
+ $Y2=0
cc_1571 VPWR N_A_1315_297#_M1000_s 0.00179197f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=-0.24
cc_1572 VPWR N_A_1315_297#_M1060_s 0.00273129f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1573 VPWR N_A_1315_297#_M1061_s 0.00210318f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1574 N_VPWR_M1000_d N_A_1315_297#_c_2915_n 0.00331615f $X=7.025 $Y=1.485
+ $X2=0 $Y2=0
cc_1575 N_VPWR_c_2085_n N_A_1315_297#_c_2915_n 0.0158304f $X=7.17 $Y=1.94 $X2=0
+ $Y2=0
cc_1576 N_VPWR_c_2085_n N_A_1315_297#_c_2919_n 0.0265477f $X=7.17 $Y=1.94 $X2=0
+ $Y2=0
cc_1577 N_VPWR_c_2015_n N_A_1315_297#_c_2923_n 0.0569572f $X=9.495 $Y=2.72 $X2=0
+ $Y2=0
cc_1578 VPWR N_A_1315_297#_c_2923_n 0.0161535f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1579 N_VPWR_c_2004_n N_A_1315_297#_c_2938_n 0.0114322f $X=7.17 $Y=2.34 $X2=0
+ $Y2=0
cc_1580 N_VPWR_c_2015_n N_A_1315_297#_c_2938_n 0.0119545f $X=9.495 $Y=2.72 $X2=0
+ $Y2=0
cc_1581 VPWR N_A_1315_297#_c_2938_n 0.00311866f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1582 VPWR N_A_1315_297#_c_2911_n 0.00591741f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1583 N_VPWR_c_2024_n N_A_1315_297#_c_2911_n 0.020978f $X=7.035 $Y=2.72 $X2=0
+ $Y2=0
cc_1584 N_VPWR_c_2085_n N_A_1315_297#_c_2912_n 0.0115021f $X=7.17 $Y=1.94 $X2=0
+ $Y2=0
cc_1585 VPWR N_A_2112_333#_M1005_s 0.00210318f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=-0.24
cc_1586 VPWR N_A_2112_333#_M1062_s 0.00273129f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1587 VPWR N_A_2112_333#_M1068_s 0.00179197f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1588 N_VPWR_c_2006_n N_A_2112_333#_c_2974_n 0.0114322f $X=12.15 $Y=2.34 $X2=0
+ $Y2=0
cc_1589 VPWR N_A_2112_333#_c_2974_n 0.0161639f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1590 N_VPWR_c_2025_n N_A_2112_333#_c_2974_n 0.0570268f $X=11.985 $Y=2.72
+ $X2=0 $Y2=0
cc_1591 VPWR N_A_2112_333#_c_2976_n 0.0031082f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1592 N_VPWR_c_2025_n N_A_2112_333#_c_2976_n 0.0118848f $X=11.985 $Y=2.72
+ $X2=0 $Y2=0
cc_1593 N_VPWR_c_2121_n N_A_2112_333#_c_2977_n 0.0265477f $X=12.15 $Y=1.94 $X2=0
+ $Y2=0
cc_1594 N_VPWR_M1001_d N_A_2112_333#_c_2980_n 0.00331615f $X=12.005 $Y=1.485
+ $X2=0 $Y2=0
cc_1595 N_VPWR_c_2121_n N_A_2112_333#_c_2980_n 0.0158304f $X=12.15 $Y=1.94 $X2=0
+ $Y2=0
cc_1596 VPWR N_A_2112_333#_c_2968_n 0.00591741f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1597 N_VPWR_c_2026_n N_A_2112_333#_c_2968_n 0.020978f $X=13.475 $Y=2.72 $X2=0
+ $Y2=0
cc_1598 N_VPWR_c_2121_n N_A_2112_333#_c_2969_n 0.0115021f $X=12.15 $Y=1.94 $X2=0
+ $Y2=0
cc_1599 VPWR N_A_2603_297#_M1014_d 0.00179197f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=-0.24
cc_1600 VPWR N_A_2603_297#_M1037_d 0.00273129f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1601 VPWR N_A_2603_297#_M1041_d 0.00210318f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1602 N_VPWR_M1014_s N_A_2603_297#_c_3031_n 0.00331615f $X=13.465 $Y=1.485
+ $X2=0 $Y2=0
cc_1603 N_VPWR_c_2129_n N_A_2603_297#_c_3031_n 0.0158304f $X=13.61 $Y=1.94 $X2=0
+ $Y2=0
cc_1604 N_VPWR_c_2129_n N_A_2603_297#_c_3035_n 0.0265477f $X=13.61 $Y=1.94 $X2=0
+ $Y2=0
cc_1605 N_VPWR_c_2017_n N_A_2603_297#_c_3039_n 0.0569572f $X=15.935 $Y=2.72
+ $X2=0 $Y2=0
cc_1606 VPWR N_A_2603_297#_c_3039_n 0.0161535f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1607 N_VPWR_c_2007_n N_A_2603_297#_c_3054_n 0.0114322f $X=13.61 $Y=2.34 $X2=0
+ $Y2=0
cc_1608 N_VPWR_c_2017_n N_A_2603_297#_c_3054_n 0.0119545f $X=15.935 $Y=2.72
+ $X2=0 $Y2=0
cc_1609 VPWR N_A_2603_297#_c_3054_n 0.00311866f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1610 VPWR N_A_2603_297#_c_3027_n 0.00591741f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1611 N_VPWR_c_2026_n N_A_2603_297#_c_3027_n 0.020978f $X=13.475 $Y=2.72 $X2=0
+ $Y2=0
cc_1612 N_VPWR_c_2129_n N_A_2603_297#_c_3028_n 0.0115021f $X=13.61 $Y=1.94 $X2=0
+ $Y2=0
cc_1613 VPWR N_A_3400_333#_M1024_d 0.00210318f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=-0.24
cc_1614 VPWR N_A_3400_333#_M1042_d 0.00273129f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1615 VPWR N_A_3400_333#_M1038_d 0.00179197f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1616 N_VPWR_c_2009_n N_A_3400_333#_c_3090_n 0.0114322f $X=18.59 $Y=2.34 $X2=0
+ $Y2=0
cc_1617 VPWR N_A_3400_333#_c_3090_n 0.0161639f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1618 N_VPWR_c_2027_n N_A_3400_333#_c_3090_n 0.0570268f $X=18.425 $Y=2.72
+ $X2=0 $Y2=0
cc_1619 VPWR N_A_3400_333#_c_3092_n 0.0031082f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1620 N_VPWR_c_2027_n N_A_3400_333#_c_3092_n 0.0118848f $X=18.425 $Y=2.72
+ $X2=0 $Y2=0
cc_1621 N_VPWR_c_2165_n N_A_3400_333#_c_3093_n 0.0265477f $X=18.59 $Y=1.94 $X2=0
+ $Y2=0
cc_1622 N_VPWR_M1025_s N_A_3400_333#_c_3096_n 0.00331615f $X=18.445 $Y=1.485
+ $X2=0 $Y2=0
cc_1623 N_VPWR_c_2165_n N_A_3400_333#_c_3096_n 0.0158304f $X=18.59 $Y=1.94 $X2=0
+ $Y2=0
cc_1624 VPWR N_A_3400_333#_c_3084_n 0.00591741f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1625 N_VPWR_c_2028_n N_A_3400_333#_c_3084_n 0.020978f $X=19.915 $Y=2.72 $X2=0
+ $Y2=0
cc_1626 N_VPWR_c_2165_n N_A_3400_333#_c_3085_n 0.0115021f $X=18.59 $Y=1.94 $X2=0
+ $Y2=0
cc_1627 VPWR N_A_3891_297#_M1029_d 0.00179197f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=-0.24
cc_1628 VPWR N_A_3891_297#_M1072_d 0.00273129f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1629 VPWR N_A_3891_297#_M1046_d 0.00210318f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1630 N_VPWR_M1029_s N_A_3891_297#_c_3147_n 0.00331615f $X=19.905 $Y=1.485
+ $X2=0 $Y2=0
cc_1631 N_VPWR_c_2173_n N_A_3891_297#_c_3147_n 0.0158304f $X=20.05 $Y=1.94 $X2=0
+ $Y2=0
cc_1632 N_VPWR_c_2173_n N_A_3891_297#_c_3151_n 0.0265477f $X=20.05 $Y=1.94 $X2=0
+ $Y2=0
cc_1633 N_VPWR_c_2019_n N_A_3891_297#_c_3155_n 0.0569572f $X=22.375 $Y=2.72
+ $X2=0 $Y2=0
cc_1634 VPWR N_A_3891_297#_c_3155_n 0.0161535f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1635 N_VPWR_c_2010_n N_A_3891_297#_c_3170_n 0.0114322f $X=20.05 $Y=2.34 $X2=0
+ $Y2=0
cc_1636 N_VPWR_c_2019_n N_A_3891_297#_c_3170_n 0.0119545f $X=22.375 $Y=2.72
+ $X2=0 $Y2=0
cc_1637 VPWR N_A_3891_297#_c_3170_n 0.00311866f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1638 VPWR N_A_3891_297#_c_3143_n 0.00591741f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1639 N_VPWR_c_2028_n N_A_3891_297#_c_3143_n 0.020978f $X=19.915 $Y=2.72 $X2=0
+ $Y2=0
cc_1640 N_VPWR_c_2173_n N_A_3891_297#_c_3144_n 0.0115021f $X=20.05 $Y=1.94 $X2=0
+ $Y2=0
cc_1641 VPWR N_A_4688_333#_M1064_d 0.00210318f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=-0.24
cc_1642 VPWR N_A_4688_333#_M1073_d 0.00481062f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1643 VPWR N_A_4688_333#_M1069_d 0.00217517f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1644 N_VPWR_c_2012_n N_A_4688_333#_c_3206_n 0.0114322f $X=25.03 $Y=2.34 $X2=0
+ $Y2=0
cc_1645 VPWR N_A_4688_333#_c_3206_n 0.0230635f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1646 N_VPWR_c_2029_n N_A_4688_333#_c_3206_n 0.0570268f $X=24.865 $Y=2.72
+ $X2=0 $Y2=0
cc_1647 VPWR N_A_4688_333#_c_3208_n 0.0031082f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1648 N_VPWR_c_2029_n N_A_4688_333#_c_3208_n 0.0118848f $X=24.865 $Y=2.72
+ $X2=0 $Y2=0
cc_1649 N_VPWR_c_2209_n N_A_4688_333#_c_3209_n 0.0272234f $X=25.03 $Y=1.94 $X2=0
+ $Y2=0
cc_1650 N_VPWR_M1030_s N_A_4688_333#_c_3212_n 0.00350459f $X=24.885 $Y=1.485
+ $X2=0 $Y2=0
cc_1651 N_VPWR_c_2209_n N_A_4688_333#_c_3212_n 0.0170301f $X=25.03 $Y=1.94 $X2=0
+ $Y2=0
cc_1652 VPWR N_A_4688_333#_c_3200_n 0.0124483f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1653 N_VPWR_c_2030_n N_A_4688_333#_c_3200_n 0.020978f $X=25.53 $Y=2.72 $X2=0
+ $Y2=0
cc_1654 N_Z_c_2384_n N_A_824_333#_M1040_d 0.00237684f $X=4.685 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_1655 N_Z_c_2385_n N_A_824_333#_M1056_d 0.00645967f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_1656 N_Z_c_2384_n N_A_824_333#_c_2850_n 0.0132602f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_1657 N_Z_c_2441_n N_A_824_333#_c_2850_n 4.86317e-19 $X=4.975 $Y=1.87 $X2=0
+ $Y2=0
cc_1658 N_Z_c_2442_n N_A_824_333#_c_2850_n 0.0212802f $X=4.83 $Y=1.87 $X2=0
+ $Y2=0
cc_1659 N_Z_c_2377_n N_A_824_333#_c_2850_n 0.00468052f $X=4.76 $Y=1.755 $X2=0
+ $Y2=0
cc_1660 N_Z_M1040_s N_A_824_333#_c_2858_n 0.00341588f $X=4.57 $Y=1.665 $X2=0
+ $Y2=0
cc_1661 N_Z_c_2384_n N_A_824_333#_c_2858_n 0.00494997f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_1662 N_Z_c_2385_n N_A_824_333#_c_2858_n 0.00415493f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_1663 N_Z_c_2441_n N_A_824_333#_c_2858_n 8.66896e-19 $X=4.975 $Y=1.87 $X2=0
+ $Y2=0
cc_1664 N_Z_c_2442_n N_A_824_333#_c_2858_n 0.0211175f $X=4.83 $Y=1.87 $X2=0
+ $Y2=0
cc_1665 N_Z_c_2385_n N_A_824_333#_c_2861_n 0.0190087f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_1666 N_Z_c_2441_n N_A_824_333#_c_2861_n 0.00221246f $X=4.975 $Y=1.87 $X2=0
+ $Y2=0
cc_1667 N_Z_c_2442_n N_A_824_333#_c_2861_n 0.024193f $X=4.83 $Y=1.87 $X2=0 $Y2=0
cc_1668 N_Z_c_2385_n N_A_824_333#_c_2864_n 0.0237468f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_1669 N_Z_c_2377_n N_A_824_333#_c_2862_n 0.00930189f $X=4.76 $Y=1.755 $X2=0
+ $Y2=0
cc_1670 N_Z_c_2385_n N_A_824_333#_c_2852_n 3.2447e-19 $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_1671 N_Z_c_2385_n N_A_824_333#_c_2853_n 0.0219733f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_1672 N_Z_c_2385_n N_A_1315_297#_M1060_s 0.00645967f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_1673 N_Z_c_2386_n N_A_1315_297#_M1061_s 0.00237684f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_1674 N_Z_c_2385_n N_A_1315_297#_c_2915_n 0.0237468f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_1675 N_Z_c_2378_n N_A_1315_297#_c_2915_n 0.00930189f $X=8.12 $Y=1.755 $X2=0
+ $Y2=0
cc_1676 N_Z_c_2385_n N_A_1315_297#_c_2919_n 0.0190087f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_1677 N_Z_c_2473_n N_A_1315_297#_c_2919_n 0.00221246f $X=8.195 $Y=1.87 $X2=0
+ $Y2=0
cc_1678 N_Z_c_2474_n N_A_1315_297#_c_2919_n 0.024193f $X=8.05 $Y=1.87 $X2=0
+ $Y2=0
cc_1679 N_Z_M1004_d N_A_1315_297#_c_2923_n 0.00341588f $X=8.02 $Y=1.665 $X2=0
+ $Y2=0
cc_1680 N_Z_c_2385_n N_A_1315_297#_c_2923_n 0.00415493f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_1681 N_Z_c_2386_n N_A_1315_297#_c_2923_n 0.00494997f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_1682 N_Z_c_2473_n N_A_1315_297#_c_2923_n 8.66896e-19 $X=8.195 $Y=1.87 $X2=0
+ $Y2=0
cc_1683 N_Z_c_2474_n N_A_1315_297#_c_2923_n 0.0211175f $X=8.05 $Y=1.87 $X2=0
+ $Y2=0
cc_1684 N_Z_c_2386_n N_A_1315_297#_c_2910_n 0.0132602f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_1685 N_Z_c_2473_n N_A_1315_297#_c_2910_n 4.86317e-19 $X=8.195 $Y=1.87 $X2=0
+ $Y2=0
cc_1686 N_Z_c_2474_n N_A_1315_297#_c_2910_n 0.0212802f $X=8.05 $Y=1.87 $X2=0
+ $Y2=0
cc_1687 N_Z_c_2378_n N_A_1315_297#_c_2910_n 0.00468052f $X=8.12 $Y=1.755 $X2=0
+ $Y2=0
cc_1688 N_Z_c_2385_n N_A_1315_297#_c_2911_n 3.2447e-19 $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_1689 N_Z_c_2385_n N_A_1315_297#_c_2912_n 0.0219733f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_1690 N_Z_c_2386_n N_A_2112_333#_M1005_s 0.00237684f $X=11.125 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_1691 N_Z_c_2387_n N_A_2112_333#_M1062_s 0.00645967f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_1692 N_Z_c_2386_n N_A_2112_333#_c_2966_n 0.0132602f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_1693 N_Z_c_2504_n N_A_2112_333#_c_2966_n 4.86317e-19 $X=11.415 $Y=1.87 $X2=0
+ $Y2=0
cc_1694 N_Z_c_2505_n N_A_2112_333#_c_2966_n 0.0212802f $X=11.27 $Y=1.87 $X2=0
+ $Y2=0
cc_1695 N_Z_c_2379_n N_A_2112_333#_c_2966_n 0.00468052f $X=11.2 $Y=1.755 $X2=0
+ $Y2=0
cc_1696 N_Z_M1005_d N_A_2112_333#_c_2974_n 0.00341588f $X=11.01 $Y=1.665 $X2=0
+ $Y2=0
cc_1697 N_Z_c_2386_n N_A_2112_333#_c_2974_n 0.00494997f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_1698 N_Z_c_2387_n N_A_2112_333#_c_2974_n 0.00415493f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_1699 N_Z_c_2504_n N_A_2112_333#_c_2974_n 8.66896e-19 $X=11.415 $Y=1.87 $X2=0
+ $Y2=0
cc_1700 N_Z_c_2505_n N_A_2112_333#_c_2974_n 0.0211175f $X=11.27 $Y=1.87 $X2=0
+ $Y2=0
cc_1701 N_Z_c_2387_n N_A_2112_333#_c_2977_n 0.0190087f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_1702 N_Z_c_2504_n N_A_2112_333#_c_2977_n 0.00221246f $X=11.415 $Y=1.87 $X2=0
+ $Y2=0
cc_1703 N_Z_c_2505_n N_A_2112_333#_c_2977_n 0.024193f $X=11.27 $Y=1.87 $X2=0
+ $Y2=0
cc_1704 N_Z_c_2387_n N_A_2112_333#_c_2980_n 0.0237468f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_1705 N_Z_c_2379_n N_A_2112_333#_c_2978_n 0.00930189f $X=11.2 $Y=1.755 $X2=0
+ $Y2=0
cc_1706 N_Z_c_2387_n N_A_2112_333#_c_2968_n 3.2447e-19 $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_1707 N_Z_c_2387_n N_A_2112_333#_c_2969_n 0.0219733f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_1708 N_Z_c_2387_n N_A_2603_297#_M1037_d 0.00645967f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_1709 N_Z_c_2388_n N_A_2603_297#_M1041_d 0.00237684f $X=17.565 $Y=1.87 $X2=0
+ $Y2=0
cc_1710 N_Z_c_2387_n N_A_2603_297#_c_3031_n 0.0237468f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_1711 N_Z_c_2380_n N_A_2603_297#_c_3031_n 0.00930189f $X=14.56 $Y=1.755 $X2=0
+ $Y2=0
cc_1712 N_Z_c_2387_n N_A_2603_297#_c_3035_n 0.0190087f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_1713 N_Z_c_2536_n N_A_2603_297#_c_3035_n 0.00221246f $X=14.635 $Y=1.87 $X2=0
+ $Y2=0
cc_1714 N_Z_c_2537_n N_A_2603_297#_c_3035_n 0.024193f $X=14.49 $Y=1.87 $X2=0
+ $Y2=0
cc_1715 N_Z_M1016_s N_A_2603_297#_c_3039_n 0.00341588f $X=14.46 $Y=1.665 $X2=0
+ $Y2=0
cc_1716 N_Z_c_2387_n N_A_2603_297#_c_3039_n 0.00415493f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_1717 N_Z_c_2388_n N_A_2603_297#_c_3039_n 0.00494997f $X=17.565 $Y=1.87 $X2=0
+ $Y2=0
cc_1718 N_Z_c_2536_n N_A_2603_297#_c_3039_n 8.66896e-19 $X=14.635 $Y=1.87 $X2=0
+ $Y2=0
cc_1719 N_Z_c_2537_n N_A_2603_297#_c_3039_n 0.0211175f $X=14.49 $Y=1.87 $X2=0
+ $Y2=0
cc_1720 N_Z_c_2388_n N_A_2603_297#_c_3026_n 0.0132602f $X=17.565 $Y=1.87 $X2=0
+ $Y2=0
cc_1721 N_Z_c_2536_n N_A_2603_297#_c_3026_n 4.86317e-19 $X=14.635 $Y=1.87 $X2=0
+ $Y2=0
cc_1722 N_Z_c_2537_n N_A_2603_297#_c_3026_n 0.0212802f $X=14.49 $Y=1.87 $X2=0
+ $Y2=0
cc_1723 N_Z_c_2380_n N_A_2603_297#_c_3026_n 0.00468052f $X=14.56 $Y=1.755 $X2=0
+ $Y2=0
cc_1724 N_Z_c_2387_n N_A_2603_297#_c_3027_n 3.2447e-19 $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_1725 N_Z_c_2387_n N_A_2603_297#_c_3028_n 0.0219733f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_1726 N_Z_c_2388_n N_A_3400_333#_M1024_d 0.00237684f $X=17.565 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_1727 N_Z_c_2389_n N_A_3400_333#_M1042_d 0.00645967f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_1728 N_Z_c_2388_n N_A_3400_333#_c_3082_n 0.0132602f $X=17.565 $Y=1.87 $X2=0
+ $Y2=0
cc_1729 N_Z_c_2567_n N_A_3400_333#_c_3082_n 4.86317e-19 $X=17.855 $Y=1.87 $X2=0
+ $Y2=0
cc_1730 N_Z_c_2568_n N_A_3400_333#_c_3082_n 0.0212802f $X=17.71 $Y=1.87 $X2=0
+ $Y2=0
cc_1731 N_Z_c_2381_n N_A_3400_333#_c_3082_n 0.00468052f $X=17.64 $Y=1.755 $X2=0
+ $Y2=0
cc_1732 N_Z_M1024_s N_A_3400_333#_c_3090_n 0.00341588f $X=17.45 $Y=1.665 $X2=0
+ $Y2=0
cc_1733 N_Z_c_2388_n N_A_3400_333#_c_3090_n 0.00494997f $X=17.565 $Y=1.87 $X2=0
+ $Y2=0
cc_1734 N_Z_c_2389_n N_A_3400_333#_c_3090_n 0.00415493f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_1735 N_Z_c_2567_n N_A_3400_333#_c_3090_n 8.66896e-19 $X=17.855 $Y=1.87 $X2=0
+ $Y2=0
cc_1736 N_Z_c_2568_n N_A_3400_333#_c_3090_n 0.0211175f $X=17.71 $Y=1.87 $X2=0
+ $Y2=0
cc_1737 N_Z_c_2389_n N_A_3400_333#_c_3093_n 0.0190087f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_1738 N_Z_c_2567_n N_A_3400_333#_c_3093_n 0.00221246f $X=17.855 $Y=1.87 $X2=0
+ $Y2=0
cc_1739 N_Z_c_2568_n N_A_3400_333#_c_3093_n 0.024193f $X=17.71 $Y=1.87 $X2=0
+ $Y2=0
cc_1740 N_Z_c_2389_n N_A_3400_333#_c_3096_n 0.0237468f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_1741 N_Z_c_2381_n N_A_3400_333#_c_3094_n 0.00930189f $X=17.64 $Y=1.755 $X2=0
+ $Y2=0
cc_1742 N_Z_c_2389_n N_A_3400_333#_c_3084_n 3.2447e-19 $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_1743 N_Z_c_2389_n N_A_3400_333#_c_3085_n 0.0219733f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_1744 N_Z_c_2389_n N_A_3891_297#_M1072_d 0.00645967f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_1745 N_Z_c_2390_n N_A_3891_297#_M1046_d 0.00237684f $X=24.005 $Y=1.87 $X2=0
+ $Y2=0
cc_1746 N_Z_c_2389_n N_A_3891_297#_c_3147_n 0.0237468f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_1747 N_Z_c_2382_n N_A_3891_297#_c_3147_n 0.00930189f $X=21 $Y=1.755 $X2=0
+ $Y2=0
cc_1748 N_Z_c_2389_n N_A_3891_297#_c_3151_n 0.0190087f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_1749 N_Z_c_2599_n N_A_3891_297#_c_3151_n 0.00221246f $X=21.075 $Y=1.87 $X2=0
+ $Y2=0
cc_1750 N_Z_c_2600_n N_A_3891_297#_c_3151_n 0.024193f $X=20.93 $Y=1.87 $X2=0
+ $Y2=0
cc_1751 N_Z_M1033_s N_A_3891_297#_c_3155_n 0.00341588f $X=20.9 $Y=1.665 $X2=0
+ $Y2=0
cc_1752 N_Z_c_2389_n N_A_3891_297#_c_3155_n 0.00415493f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_1753 N_Z_c_2390_n N_A_3891_297#_c_3155_n 0.00494997f $X=24.005 $Y=1.87 $X2=0
+ $Y2=0
cc_1754 N_Z_c_2599_n N_A_3891_297#_c_3155_n 8.66896e-19 $X=21.075 $Y=1.87 $X2=0
+ $Y2=0
cc_1755 N_Z_c_2600_n N_A_3891_297#_c_3155_n 0.0211175f $X=20.93 $Y=1.87 $X2=0
+ $Y2=0
cc_1756 N_Z_c_2390_n N_A_3891_297#_c_3142_n 0.0132602f $X=24.005 $Y=1.87 $X2=0
+ $Y2=0
cc_1757 N_Z_c_2599_n N_A_3891_297#_c_3142_n 4.86317e-19 $X=21.075 $Y=1.87 $X2=0
+ $Y2=0
cc_1758 N_Z_c_2600_n N_A_3891_297#_c_3142_n 0.0212802f $X=20.93 $Y=1.87 $X2=0
+ $Y2=0
cc_1759 N_Z_c_2382_n N_A_3891_297#_c_3142_n 0.00468052f $X=21 $Y=1.755 $X2=0
+ $Y2=0
cc_1760 N_Z_c_2389_n N_A_3891_297#_c_3143_n 3.2447e-19 $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_1761 N_Z_c_2389_n N_A_3891_297#_c_3144_n 0.0219733f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_1762 N_Z_c_2390_n N_A_4688_333#_M1064_d 0.00237684f $X=24.005 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_1763 N_Z_c_2390_n N_A_4688_333#_c_3198_n 0.0132602f $X=24.005 $Y=1.87 $X2=0
+ $Y2=0
cc_1764 Z N_A_4688_333#_c_3198_n 4.86317e-19 $X=24.065 $Y=1.785 $X2=0 $Y2=0
cc_1765 N_Z_c_2630_n N_A_4688_333#_c_3198_n 0.0212802f $X=24.15 $Y=1.87 $X2=0
+ $Y2=0
cc_1766 N_Z_c_2383_n N_A_4688_333#_c_3198_n 0.00468052f $X=24.08 $Y=1.755 $X2=0
+ $Y2=0
cc_1767 N_Z_M1064_s N_A_4688_333#_c_3206_n 0.00341588f $X=23.89 $Y=1.665 $X2=0
+ $Y2=0
cc_1768 N_Z_c_2390_n N_A_4688_333#_c_3206_n 0.00494997f $X=24.005 $Y=1.87 $X2=0
+ $Y2=0
cc_1769 Z N_A_4688_333#_c_3206_n 8.66896e-19 $X=24.065 $Y=1.785 $X2=0 $Y2=0
cc_1770 N_Z_c_2630_n N_A_4688_333#_c_3206_n 0.0211175f $X=24.15 $Y=1.87 $X2=0
+ $Y2=0
cc_1771 Z N_A_4688_333#_c_3209_n 0.0062686f $X=24.065 $Y=1.785 $X2=0 $Y2=0
cc_1772 N_Z_c_2630_n N_A_4688_333#_c_3209_n 0.0235305f $X=24.15 $Y=1.87 $X2=0
+ $Y2=0
cc_1773 N_Z_c_2383_n N_A_4688_333#_c_3210_n 0.00930189f $X=24.08 $Y=1.755 $X2=0
+ $Y2=0
cc_1774 N_Z_c_2368_n N_A_27_47#_c_3247_n 0.00729487f $X=1.67 $Y=0.68 $X2=0 $Y2=0
cc_1775 N_Z_c_2376_n N_A_27_47#_c_3247_n 0.00238404f $X=1.68 $Y=1.755 $X2=0
+ $Y2=0
cc_1776 N_Z_M1017_s N_A_27_47#_c_3249_n 0.00165831f $X=1.535 $Y=0.345 $X2=0
+ $Y2=0
cc_1777 N_Z_c_2368_n N_A_27_47#_c_3249_n 0.0156951f $X=1.67 $Y=0.68 $X2=0 $Y2=0
cc_1778 N_Z_M1015_s N_A_845_69#_c_3574_n 0.00165831f $X=4.635 $Y=0.345 $X2=0
+ $Y2=0
cc_1779 N_Z_c_2369_n N_A_845_69#_c_3574_n 0.0156951f $X=4.77 $Y=0.68 $X2=0 $Y2=0
cc_1780 N_Z_c_2369_n N_A_845_69#_c_3577_n 0.00729487f $X=4.77 $Y=0.68 $X2=0
+ $Y2=0
cc_1781 N_Z_c_2377_n N_A_845_69#_c_3577_n 0.00238404f $X=4.76 $Y=1.755 $X2=0
+ $Y2=0
cc_1782 N_Z_c_2370_n N_A_1315_47#_c_3622_n 0.00729487f $X=8.11 $Y=0.68 $X2=0
+ $Y2=0
cc_1783 N_Z_c_2378_n N_A_1315_47#_c_3622_n 0.00238404f $X=8.12 $Y=1.755 $X2=0
+ $Y2=0
cc_1784 N_Z_M1058_d N_A_1315_47#_c_3624_n 0.00165831f $X=7.975 $Y=0.345 $X2=0
+ $Y2=0
cc_1785 N_Z_c_2370_n N_A_1315_47#_c_3624_n 0.0156951f $X=8.11 $Y=0.68 $X2=0
+ $Y2=0
cc_1786 N_Z_M1052_d N_A_2133_69#_c_3666_n 0.00165831f $X=11.075 $Y=0.345 $X2=0
+ $Y2=0
cc_1787 N_Z_c_2371_n N_A_2133_69#_c_3666_n 0.0156951f $X=11.21 $Y=0.68 $X2=0
+ $Y2=0
cc_1788 N_Z_c_2371_n N_A_2133_69#_c_3669_n 0.00729487f $X=11.21 $Y=0.68 $X2=0
+ $Y2=0
cc_1789 N_Z_c_2379_n N_A_2133_69#_c_3669_n 0.00238404f $X=11.2 $Y=1.755 $X2=0
+ $Y2=0
cc_1790 N_Z_c_2372_n N_A_2603_47#_c_3714_n 0.00729487f $X=14.55 $Y=0.68 $X2=0
+ $Y2=0
cc_1791 N_Z_c_2380_n N_A_2603_47#_c_3714_n 0.00238404f $X=14.56 $Y=1.755 $X2=0
+ $Y2=0
cc_1792 N_Z_M1021_d N_A_2603_47#_c_3716_n 0.00165831f $X=14.415 $Y=0.345 $X2=0
+ $Y2=0
cc_1793 N_Z_c_2372_n N_A_2603_47#_c_3716_n 0.0156951f $X=14.55 $Y=0.68 $X2=0
+ $Y2=0
cc_1794 N_Z_M1010_d N_A_3421_69#_c_3758_n 0.00165831f $X=17.515 $Y=0.345 $X2=0
+ $Y2=0
cc_1795 N_Z_c_2373_n N_A_3421_69#_c_3758_n 0.0156951f $X=17.65 $Y=0.68 $X2=0
+ $Y2=0
cc_1796 N_Z_c_2373_n N_A_3421_69#_c_3761_n 0.00729487f $X=17.65 $Y=0.68 $X2=0
+ $Y2=0
cc_1797 N_Z_c_2381_n N_A_3421_69#_c_3761_n 0.00238404f $X=17.64 $Y=1.755 $X2=0
+ $Y2=0
cc_1798 N_Z_c_2374_n N_A_3891_47#_c_3806_n 0.00729487f $X=20.99 $Y=0.68 $X2=0
+ $Y2=0
cc_1799 N_Z_c_2382_n N_A_3891_47#_c_3806_n 0.00238404f $X=21 $Y=1.755 $X2=0
+ $Y2=0
cc_1800 N_Z_M1059_d N_A_3891_47#_c_3808_n 0.00165831f $X=20.855 $Y=0.345 $X2=0
+ $Y2=0
cc_1801 N_Z_c_2374_n N_A_3891_47#_c_3808_n 0.0156951f $X=20.99 $Y=0.68 $X2=0
+ $Y2=0
cc_1802 N_Z_M1055_d N_A_4709_69#_c_3850_n 0.00165831f $X=23.955 $Y=0.345 $X2=0
+ $Y2=0
cc_1803 N_Z_c_2375_n N_A_4709_69#_c_3850_n 0.0156951f $X=24.09 $Y=0.68 $X2=0
+ $Y2=0
cc_1804 N_Z_c_2375_n N_A_4709_69#_c_3853_n 0.00729487f $X=24.09 $Y=0.68 $X2=0
+ $Y2=0
cc_1805 N_Z_c_2383_n N_A_4709_69#_c_3853_n 0.00238404f $X=24.08 $Y=1.755 $X2=0
+ $Y2=0
cc_1806 N_A_824_333#_c_2851_n N_A_1315_297#_c_2909_n 0.0147157f $X=6.195
+ $Y=1.665 $X2=0 $Y2=0
cc_1807 N_A_824_333#_c_2852_n N_A_1315_297#_c_2911_n 0.0296136f $X=6.18 $Y=2.34
+ $X2=0 $Y2=0
cc_1808 N_A_824_333#_c_2853_n N_A_1315_297#_c_2912_n 0.0296136f $X=6.18 $Y=2.21
+ $X2=0 $Y2=0
cc_1809 N_A_824_333#_c_2864_n N_A_845_69#_c_3576_n 0.00251701f $X=6.045 $Y=1.58
+ $X2=0 $Y2=0
cc_1810 N_A_824_333#_c_2864_n N_A_845_69#_c_3577_n 0.00200781f $X=6.045 $Y=1.58
+ $X2=0 $Y2=0
cc_1811 N_A_824_333#_c_2862_n N_A_845_69#_c_3577_n 0.00650395f $X=5.325 $Y=1.58
+ $X2=0 $Y2=0
cc_1812 N_A_1315_297#_c_2915_n N_A_1315_47#_c_3622_n 0.0110288f $X=7.555 $Y=1.58
+ $X2=0 $Y2=0
cc_1813 N_A_2112_333#_c_2967_n N_A_2603_297#_c_3025_n 0.0147157f $X=12.635
+ $Y=1.665 $X2=0 $Y2=0
cc_1814 N_A_2112_333#_c_2968_n N_A_2603_297#_c_3027_n 0.0296136f $X=12.62
+ $Y=2.34 $X2=0 $Y2=0
cc_1815 N_A_2112_333#_c_2969_n N_A_2603_297#_c_3028_n 0.0296136f $X=12.62
+ $Y=2.21 $X2=0 $Y2=0
cc_1816 N_A_2112_333#_c_2980_n N_A_2133_69#_c_3668_n 0.00251701f $X=12.485
+ $Y=1.58 $X2=0 $Y2=0
cc_1817 N_A_2112_333#_c_2980_n N_A_2133_69#_c_3669_n 0.00200781f $X=12.485
+ $Y=1.58 $X2=0 $Y2=0
cc_1818 N_A_2112_333#_c_2978_n N_A_2133_69#_c_3669_n 0.00650395f $X=11.765
+ $Y=1.58 $X2=0 $Y2=0
cc_1819 N_A_2603_297#_c_3031_n N_A_2603_47#_c_3714_n 0.0110288f $X=13.995
+ $Y=1.58 $X2=0 $Y2=0
cc_1820 N_A_3400_333#_c_3083_n N_A_3891_297#_c_3141_n 0.0147157f $X=19.075
+ $Y=1.665 $X2=0 $Y2=0
cc_1821 N_A_3400_333#_c_3084_n N_A_3891_297#_c_3143_n 0.0296136f $X=19.06
+ $Y=2.34 $X2=0 $Y2=0
cc_1822 N_A_3400_333#_c_3085_n N_A_3891_297#_c_3144_n 0.0296136f $X=19.06
+ $Y=2.21 $X2=0 $Y2=0
cc_1823 N_A_3400_333#_c_3096_n N_A_3421_69#_c_3760_n 0.00251701f $X=18.925
+ $Y=1.58 $X2=0 $Y2=0
cc_1824 N_A_3400_333#_c_3096_n N_A_3421_69#_c_3761_n 0.00200781f $X=18.925
+ $Y=1.58 $X2=0 $Y2=0
cc_1825 N_A_3400_333#_c_3094_n N_A_3421_69#_c_3761_n 0.00650395f $X=18.205
+ $Y=1.58 $X2=0 $Y2=0
cc_1826 N_A_3891_297#_c_3147_n N_A_3891_47#_c_3806_n 0.0110288f $X=20.435
+ $Y=1.58 $X2=0 $Y2=0
cc_1827 N_A_4688_333#_c_3212_n N_A_4709_69#_c_3852_n 0.00251701f $X=25.365
+ $Y=1.58 $X2=0 $Y2=0
cc_1828 N_A_4688_333#_c_3212_n N_A_4709_69#_c_3853_n 0.00200781f $X=25.365
+ $Y=1.58 $X2=0 $Y2=0
cc_1829 N_A_4688_333#_c_3210_n N_A_4709_69#_c_3853_n 0.00650395f $X=24.645
+ $Y=1.58 $X2=0 $Y2=0
cc_1830 N_A_27_47#_c_3247_n N_VGND_M1019_s 0.00306532f $X=1.03 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_1831 N_A_27_47#_c_3247_n N_VGND_c_3289_n 0.012179f $X=1.03 $Y=0.8 $X2=0 $Y2=0
cc_1832 N_A_27_47#_c_3247_n N_VGND_c_3304_n 0.00219745f $X=1.03 $Y=0.8 $X2=0
+ $Y2=0
cc_1833 N_A_27_47#_c_3279_p N_VGND_c_3304_n 0.0199987f $X=1.182 $Y=0.425 $X2=0
+ $Y2=0
cc_1834 N_A_27_47#_c_3249_n N_VGND_c_3304_n 0.0535945f $X=2.005 $Y=0.34 $X2=0
+ $Y2=0
cc_1835 N_A_27_47#_M1019_d VGND 0.00288496f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_1836 N_A_27_47#_M1053_d VGND 0.0024283f $X=1.015 $Y=0.235 $X2=0 $Y2=0
cc_1837 N_A_27_47#_c_3250_n VGND 0.0124017f $X=0.31 $Y=0.38 $X2=0 $Y2=0
cc_1838 N_A_27_47#_c_3247_n VGND 0.00838939f $X=1.03 $Y=0.8 $X2=0 $Y2=0
cc_1839 N_A_27_47#_c_3279_p VGND 0.0117415f $X=1.182 $Y=0.425 $X2=0 $Y2=0
cc_1840 N_A_27_47#_c_3249_n VGND 0.0279432f $X=2.005 $Y=0.34 $X2=0 $Y2=0
cc_1841 N_A_27_47#_c_3250_n N_VGND_c_3319_n 0.020879f $X=0.31 $Y=0.38 $X2=0
+ $Y2=0
cc_1842 N_A_27_47#_c_3247_n N_VGND_c_3319_n 0.0020257f $X=1.03 $Y=0.8 $X2=0
+ $Y2=0
cc_1843 VGND N_A_845_69#_M1018_d 0.0024283f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1844 VGND N_A_845_69#_M1051_s 0.00288496f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1845 VGND N_A_845_69#_c_3574_n 0.0222193f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1846 N_VGND_c_3315_n N_A_845_69#_c_3574_n 0.0422314f $X=5.58 $Y=0 $X2=0 $Y2=0
cc_1847 VGND N_A_845_69#_c_3575_n 0.00572388f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1848 N_VGND_c_3315_n N_A_845_69#_c_3575_n 0.0113631f $X=5.58 $Y=0 $X2=0 $Y2=0
cc_1849 VGND N_A_845_69#_c_3611_n 0.0117415f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1850 N_VGND_c_3315_n N_A_845_69#_c_3611_n 0.0199987f $X=5.58 $Y=0 $X2=0 $Y2=0
cc_1851 N_VGND_M1036_d N_A_845_69#_c_3576_n 0.00306532f $X=5.575 $Y=0.235 $X2=0
+ $Y2=0
cc_1852 N_VGND_c_3291_n N_A_845_69#_c_3576_n 0.012179f $X=5.71 $Y=0.38 $X2=0
+ $Y2=0
cc_1853 N_VGND_c_3292_n N_A_845_69#_c_3576_n 0.0020257f $X=7.085 $Y=0 $X2=0
+ $Y2=0
cc_1854 VGND N_A_845_69#_c_3576_n 0.00838939f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1855 N_VGND_c_3315_n N_A_845_69#_c_3576_n 0.00219745f $X=5.58 $Y=0 $X2=0
+ $Y2=0
cc_1856 N_VGND_c_3292_n N_A_845_69#_c_3596_n 0.020879f $X=7.085 $Y=0 $X2=0 $Y2=0
cc_1857 VGND N_A_845_69#_c_3596_n 0.0124017f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1858 VGND N_A_1315_47#_M1057_d 0.00288496f $X=25.445 $Y=-0.085 $X2=-0.19
+ $Y2=-0.24
cc_1859 VGND N_A_1315_47#_M1063_d 0.0024283f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1860 N_VGND_c_3292_n N_A_1315_47#_c_3625_n 0.020879f $X=7.085 $Y=0 $X2=0
+ $Y2=0
cc_1861 VGND N_A_1315_47#_c_3625_n 0.0124017f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1862 N_VGND_M1057_s N_A_1315_47#_c_3622_n 0.00306532f $X=7.035 $Y=0.235 $X2=0
+ $Y2=0
cc_1863 N_VGND_c_3292_n N_A_1315_47#_c_3622_n 0.0020257f $X=7.085 $Y=0 $X2=0
+ $Y2=0
cc_1864 N_VGND_c_3293_n N_A_1315_47#_c_3622_n 0.012179f $X=7.17 $Y=0.38 $X2=0
+ $Y2=0
cc_1865 N_VGND_c_3306_n N_A_1315_47#_c_3622_n 0.00219745f $X=9.535 $Y=0 $X2=0
+ $Y2=0
cc_1866 VGND N_A_1315_47#_c_3622_n 0.00838939f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1867 N_VGND_c_3306_n N_A_1315_47#_c_3660_n 0.0199987f $X=9.535 $Y=0 $X2=0
+ $Y2=0
cc_1868 VGND N_A_1315_47#_c_3660_n 0.0117415f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1869 N_VGND_c_3306_n N_A_1315_47#_c_3624_n 0.0535945f $X=9.535 $Y=0 $X2=0
+ $Y2=0
cc_1870 VGND N_A_1315_47#_c_3624_n 0.0279432f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1871 VGND N_A_2133_69#_M1065_s 0.0024283f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1872 VGND N_A_2133_69#_M1078_d 0.00288496f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1873 VGND N_A_2133_69#_c_3666_n 0.0222193f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1874 N_VGND_c_3316_n N_A_2133_69#_c_3666_n 0.0422314f $X=12.02 $Y=0 $X2=0
+ $Y2=0
cc_1875 VGND N_A_2133_69#_c_3667_n 0.00572388f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1876 N_VGND_c_3316_n N_A_2133_69#_c_3667_n 0.0113631f $X=12.02 $Y=0 $X2=0
+ $Y2=0
cc_1877 VGND N_A_2133_69#_c_3703_n 0.0117415f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1878 N_VGND_c_3316_n N_A_2133_69#_c_3703_n 0.0199987f $X=12.02 $Y=0 $X2=0
+ $Y2=0
cc_1879 N_VGND_M1012_s N_A_2133_69#_c_3668_n 0.00306532f $X=12.015 $Y=0.235
+ $X2=0 $Y2=0
cc_1880 N_VGND_c_3295_n N_A_2133_69#_c_3668_n 0.012179f $X=12.15 $Y=0.38 $X2=0
+ $Y2=0
cc_1881 N_VGND_c_3296_n N_A_2133_69#_c_3668_n 0.0020257f $X=13.525 $Y=0 $X2=0
+ $Y2=0
cc_1882 VGND N_A_2133_69#_c_3668_n 0.00838939f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1883 N_VGND_c_3316_n N_A_2133_69#_c_3668_n 0.00219745f $X=12.02 $Y=0 $X2=0
+ $Y2=0
cc_1884 N_VGND_c_3296_n N_A_2133_69#_c_3688_n 0.020879f $X=13.525 $Y=0 $X2=0
+ $Y2=0
cc_1885 VGND N_A_2133_69#_c_3688_n 0.0124017f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1886 VGND N_A_2603_47#_M1031_s 0.00288496f $X=25.445 $Y=-0.085 $X2=-0.19
+ $Y2=-0.24
cc_1887 VGND N_A_2603_47#_M1048_s 0.0024283f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1888 N_VGND_c_3296_n N_A_2603_47#_c_3717_n 0.020879f $X=13.525 $Y=0 $X2=0
+ $Y2=0
cc_1889 VGND N_A_2603_47#_c_3717_n 0.0124017f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1890 N_VGND_M1031_d N_A_2603_47#_c_3714_n 0.00306532f $X=13.475 $Y=0.235
+ $X2=0 $Y2=0
cc_1891 N_VGND_c_3296_n N_A_2603_47#_c_3714_n 0.0020257f $X=13.525 $Y=0 $X2=0
+ $Y2=0
cc_1892 N_VGND_c_3297_n N_A_2603_47#_c_3714_n 0.012179f $X=13.61 $Y=0.38 $X2=0
+ $Y2=0
cc_1893 N_VGND_c_3308_n N_A_2603_47#_c_3714_n 0.00219745f $X=15.975 $Y=0 $X2=0
+ $Y2=0
cc_1894 VGND N_A_2603_47#_c_3714_n 0.00838939f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1895 N_VGND_c_3308_n N_A_2603_47#_c_3752_n 0.0199987f $X=15.975 $Y=0 $X2=0
+ $Y2=0
cc_1896 VGND N_A_2603_47#_c_3752_n 0.0117415f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1897 N_VGND_c_3308_n N_A_2603_47#_c_3716_n 0.0535945f $X=15.975 $Y=0 $X2=0
+ $Y2=0
cc_1898 VGND N_A_2603_47#_c_3716_n 0.0279432f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1899 VGND N_A_3421_69#_M1026_s 0.0024283f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1900 VGND N_A_3421_69#_M1054_s 0.00288496f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1901 VGND N_A_3421_69#_c_3758_n 0.0222193f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1902 N_VGND_c_3317_n N_A_3421_69#_c_3758_n 0.0422314f $X=18.46 $Y=0 $X2=0
+ $Y2=0
cc_1903 VGND N_A_3421_69#_c_3759_n 0.00572388f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1904 N_VGND_c_3317_n N_A_3421_69#_c_3759_n 0.0113631f $X=18.46 $Y=0 $X2=0
+ $Y2=0
cc_1905 VGND N_A_3421_69#_c_3795_n 0.0117415f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1906 N_VGND_c_3317_n N_A_3421_69#_c_3795_n 0.0199987f $X=18.46 $Y=0 $X2=0
+ $Y2=0
cc_1907 N_VGND_M1047_d N_A_3421_69#_c_3760_n 0.00306532f $X=18.455 $Y=0.235
+ $X2=0 $Y2=0
cc_1908 N_VGND_c_3299_n N_A_3421_69#_c_3760_n 0.012179f $X=18.59 $Y=0.38 $X2=0
+ $Y2=0
cc_1909 N_VGND_c_3300_n N_A_3421_69#_c_3760_n 0.0020257f $X=19.965 $Y=0 $X2=0
+ $Y2=0
cc_1910 VGND N_A_3421_69#_c_3760_n 0.00838939f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1911 N_VGND_c_3317_n N_A_3421_69#_c_3760_n 0.00219745f $X=18.46 $Y=0 $X2=0
+ $Y2=0
cc_1912 N_VGND_c_3300_n N_A_3421_69#_c_3780_n 0.020879f $X=19.965 $Y=0 $X2=0
+ $Y2=0
cc_1913 VGND N_A_3421_69#_c_3780_n 0.0124017f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1914 VGND N_A_3891_47#_M1070_s 0.00288496f $X=25.445 $Y=-0.085 $X2=-0.19
+ $Y2=-0.24
cc_1915 VGND N_A_3891_47#_M1079_s 0.0024283f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1916 N_VGND_c_3300_n N_A_3891_47#_c_3809_n 0.020879f $X=19.965 $Y=0 $X2=0
+ $Y2=0
cc_1917 VGND N_A_3891_47#_c_3809_n 0.0124017f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1918 N_VGND_M1070_d N_A_3891_47#_c_3806_n 0.00306532f $X=19.915 $Y=0.235
+ $X2=0 $Y2=0
cc_1919 N_VGND_c_3300_n N_A_3891_47#_c_3806_n 0.0020257f $X=19.965 $Y=0 $X2=0
+ $Y2=0
cc_1920 N_VGND_c_3301_n N_A_3891_47#_c_3806_n 0.012179f $X=20.05 $Y=0.38 $X2=0
+ $Y2=0
cc_1921 N_VGND_c_3310_n N_A_3891_47#_c_3806_n 0.00219745f $X=22.415 $Y=0 $X2=0
+ $Y2=0
cc_1922 VGND N_A_3891_47#_c_3806_n 0.00838939f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1923 N_VGND_c_3310_n N_A_3891_47#_c_3844_n 0.0199987f $X=22.415 $Y=0 $X2=0
+ $Y2=0
cc_1924 VGND N_A_3891_47#_c_3844_n 0.0117415f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1925 N_VGND_c_3310_n N_A_3891_47#_c_3808_n 0.0535945f $X=22.415 $Y=0 $X2=0
+ $Y2=0
cc_1926 VGND N_A_3891_47#_c_3808_n 0.0279432f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1927 VGND N_A_4709_69#_M1071_s 0.0024283f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1928 VGND N_A_4709_69#_M1027_d 0.00288496f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1929 N_VGND_c_3312_n N_A_4709_69#_c_3850_n 0.0422314f $X=24.9 $Y=0 $X2=0
+ $Y2=0
cc_1930 VGND N_A_4709_69#_c_3850_n 0.0222193f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1931 N_VGND_c_3312_n N_A_4709_69#_c_3851_n 0.0113631f $X=24.9 $Y=0 $X2=0
+ $Y2=0
cc_1932 VGND N_A_4709_69#_c_3851_n 0.00572388f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1933 N_VGND_c_3312_n N_A_4709_69#_c_3887_n 0.0199987f $X=24.9 $Y=0 $X2=0
+ $Y2=0
cc_1934 VGND N_A_4709_69#_c_3887_n 0.0117415f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1935 N_VGND_M1011_s N_A_4709_69#_c_3852_n 0.00306532f $X=24.895 $Y=0.235
+ $X2=0 $Y2=0
cc_1936 N_VGND_c_3303_n N_A_4709_69#_c_3852_n 0.012179f $X=25.03 $Y=0.38 $X2=0
+ $Y2=0
cc_1937 N_VGND_c_3312_n N_A_4709_69#_c_3852_n 0.00219745f $X=24.9 $Y=0 $X2=0
+ $Y2=0
cc_1938 VGND N_A_4709_69#_c_3852_n 0.00838939f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1939 N_VGND_c_3318_n N_A_4709_69#_c_3852_n 0.0020257f $X=25.53 $Y=0 $X2=0
+ $Y2=0
cc_1940 VGND N_A_4709_69#_c_3872_n 0.0124017f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1941 N_VGND_c_3318_n N_A_4709_69#_c_3872_n 0.020879f $X=25.53 $Y=0 $X2=0
+ $Y2=0
cc_1942 N_A_845_69#_c_3596_n N_A_1315_47#_c_3625_n 0.0248576f $X=6.13 $Y=0.38
+ $X2=0 $Y2=0
cc_1943 N_A_845_69#_c_3576_n N_A_1315_47#_c_3623_n 0.0103099f $X=5.965 $Y=0.8
+ $X2=0 $Y2=0
cc_1944 N_A_2133_69#_c_3688_n N_A_2603_47#_c_3717_n 0.0248576f $X=12.57 $Y=0.38
+ $X2=0 $Y2=0
cc_1945 N_A_2133_69#_c_3668_n N_A_2603_47#_c_3715_n 0.0103099f $X=12.405 $Y=0.8
+ $X2=0 $Y2=0
cc_1946 N_A_3421_69#_c_3780_n N_A_3891_47#_c_3809_n 0.0248576f $X=19.01 $Y=0.38
+ $X2=0 $Y2=0
cc_1947 N_A_3421_69#_c_3760_n N_A_3891_47#_c_3807_n 0.0103099f $X=18.845 $Y=0.8
+ $X2=0 $Y2=0
