* File: sky130_fd_sc_hdll__muxb8to1_1.spice
* Created: Wed Sep  2 08:36:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__muxb8to1_1.pex.spice"
.subckt sky130_fd_sc_hdll__muxb8to1_1  VNB VPB D[0] S[0] S[1] D[1] D[2] S[2]
+ S[3] D[3] D[4] S[4] S[5] D[5] D[6] S[6] S[7] D[7] VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* D[7]	D[7]
* S[7]	S[7]
* S[6]	S[6]
* D[6]	D[6]
* D[5]	D[5]
* S[5]	S[5]
* S[4]	S[4]
* D[4]	D[4]
* D[3]	D[3]
* S[3]	S[3]
* S[2]	S[2]
* D[2]	D[2]
* D[1]	D[1]
* S[1]	S[1]
* S[0]	S[0]
* D[0]	D[0]
* VPB	VPB
* VNB	VNB
MM1040 A_109_47# N_D[0]_M1040_g N_VGND_M1040_s VNB NSHORT L=0.15 W=0.65
+ AD=0.111944 AS=0.169 PD=1.08333 PS=1.82 NRD=21.636 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1044 N_Z_M1044_d N_S[0]_M1044_g A_109_47# VNB NSHORT L=0.15 W=0.52 AD=0.1352
+ AS=0.0895556 PD=1.56 PS=0.866667 NRD=0 NRS=27.048 M=1 R=3.46667 SA=75000.7
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1029 N_VGND_M1029_d N_S[0]_M1029_g N_A_184_265#_M1029_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1118 AS=0.1482 PD=0.95 PS=1.61 NRD=17.304 NRS=4.608 M=1 R=3.46667
+ SA=75000.2 SB=75000.8 A=0.078 P=1.34 MULT=1
MM1028 N_A_533_47#_M1028_d N_S[1]_M1028_g N_VGND_M1029_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1482 AS=0.1118 PD=1.61 PS=0.95 NRD=4.608 NRS=17.304 M=1 R=3.46667
+ SA=75000.8 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1014 A_746_47# N_S[1]_M1014_g N_Z_M1014_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0895556 AS=0.1352 PD=0.866667 PS=1.56 NRD=27.048 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1032 N_VGND_M1032_d N_D[1]_M1032_g A_746_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.111944 PD=0.98 PS=1.08333 NRD=4.608 NRS=21.636 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1001 A_937_47# N_D[2]_M1001_g N_VGND_M1032_d VNB NSHORT L=0.15 W=0.65
+ AD=0.111944 AS=0.10725 PD=1.08333 PS=0.98 NRD=21.636 NRS=4.608 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1010 N_Z_M1010_d N_S[2]_M1010_g A_937_47# VNB NSHORT L=0.15 W=0.52 AD=0.1352
+ AS=0.0895556 PD=1.56 PS=0.866667 NRD=0 NRS=27.048 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1042 N_VGND_M1042_d N_S[2]_M1042_g N_A_1012_265#_M1042_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1118 AS=0.1482 PD=0.95 PS=1.61 NRD=17.304 NRS=4.608 M=1 R=3.46667
+ SA=75000.2 SB=75000.8 A=0.078 P=1.34 MULT=1
MM1027 N_A_1361_47#_M1027_d N_S[3]_M1027_g N_VGND_M1042_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1482 AS=0.1118 PD=1.61 PS=0.95 NRD=4.608 NRS=17.304 M=1 R=3.46667
+ SA=75000.8 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1008 A_1574_47# N_S[3]_M1008_g N_Z_M1008_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0895556 AS=0.1352 PD=0.866667 PS=1.56 NRD=27.048 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1039 N_VGND_M1039_d N_D[3]_M1039_g A_1574_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.111944 PD=0.98 PS=1.08333 NRD=4.608 NRS=21.636 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1000 A_1765_47# N_D[4]_M1000_g N_VGND_M1039_d VNB NSHORT L=0.15 W=0.65
+ AD=0.111944 AS=0.10725 PD=1.08333 PS=0.98 NRD=21.636 NRS=4.608 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1018 N_Z_M1018_d N_S[4]_M1018_g A_1765_47# VNB NSHORT L=0.15 W=0.52 AD=0.1352
+ AS=0.0895556 PD=1.56 PS=0.866667 NRD=0 NRS=27.048 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1046 N_VGND_M1046_d N_S[4]_M1046_g N_A_1840_265#_M1046_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1118 AS=0.1482 PD=0.95 PS=1.61 NRD=17.304 NRS=4.608 M=1 R=3.46667
+ SA=75000.2 SB=75000.8 A=0.078 P=1.34 MULT=1
MM1037 N_A_2189_47#_M1037_d N_S[5]_M1037_g N_VGND_M1046_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1482 AS=0.1118 PD=1.61 PS=0.95 NRD=4.608 NRS=17.304 M=1 R=3.46667
+ SA=75000.8 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1012 A_2402_47# N_S[5]_M1012_g N_Z_M1012_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0895556 AS=0.1352 PD=0.866667 PS=1.56 NRD=27.048 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1041 N_VGND_M1041_d N_D[5]_M1041_g A_2402_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.111944 PD=0.98 PS=1.08333 NRD=4.608 NRS=21.636 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1002 A_2593_47# N_D[6]_M1002_g N_VGND_M1041_d VNB NSHORT L=0.15 W=0.65
+ AD=0.111944 AS=0.10725 PD=1.08333 PS=0.98 NRD=21.636 NRS=4.608 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1033 N_Z_M1033_d N_S[6]_M1033_g A_2593_47# VNB NSHORT L=0.15 W=0.52 AD=0.1352
+ AS=0.0895556 PD=1.56 PS=0.866667 NRD=0 NRS=27.048 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1004 N_VGND_M1004_d N_S[6]_M1004_g N_A_2668_265#_M1004_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1118 AS=0.1482 PD=0.95 PS=1.61 NRD=17.304 NRS=4.608 M=1 R=3.46667
+ SA=75000.2 SB=75000.8 A=0.078 P=1.34 MULT=1
MM1047 N_A_3017_47#_M1047_d N_S[7]_M1047_g N_VGND_M1004_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1482 AS=0.1118 PD=1.61 PS=0.95 NRD=4.608 NRS=17.304 M=1 R=3.46667
+ SA=75000.8 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1031 A_3230_47# N_S[7]_M1031_g N_Z_M1031_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0895556 AS=0.1352 PD=0.866667 PS=1.56 NRD=27.048 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.7 A=0.078 P=1.34 MULT=1
MM1043 N_VGND_M1043_d N_D[7]_M1043_g A_3230_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.111944 PD=1.82 PS=1.08333 NRD=0 NRS=21.636 M=1 R=4.33333
+ SA=75000.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1015 A_117_297# N_D[0]_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.27 PD=1.47802 PS=2.54 NRD=24.8417 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1019 N_Z_M1019_d N_A_184_265#_M1019_g A_117_297# VPB PHIGHVT L=0.18 W=0.82
+ AD=0.2214 AS=0.148546 PD=2.18 PS=1.21198 NRD=1.182 NRS=30.2986 M=1 R=4.55556
+ SA=90000.7 SB=90000.2 A=0.1476 P=2 MULT=1
MM1023 N_VPWR_M1023_d N_S[0]_M1023_g N_A_184_265#_M1023_s VPB PHIGHVT L=0.18 W=1
+ AD=0.2 AS=0.27 PD=1.4 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1020 N_A_533_47#_M1020_d N_S[1]_M1020_g N_VPWR_M1023_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.2 PD=2.54 PS=1.4 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90000.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1009 A_734_333# N_A_533_47#_M1009_g N_Z_M1009_s VPB PHIGHVT L=0.18 W=0.82
+ AD=0.148546 AS=0.2214 PD=1.21198 PS=2.18 NRD=30.2986 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.8 A=0.1476 P=2 MULT=1
MM1035 N_VPWR_M1035_d N_D[1]_M1035_g A_734_333# VPB PHIGHVT L=0.18 W=1 AD=0.175
+ AS=0.181154 PD=1.35 PS=1.47802 NRD=6.8753 NRS=24.8417 M=1 R=5.55556 SA=90000.6
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1021 A_945_297# N_D[2]_M1021_g N_VPWR_M1035_d VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.175 PD=1.47802 PS=1.35 NRD=24.8417 NRS=6.8753 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1022 N_Z_M1022_d N_A_1012_265#_M1022_g A_945_297# VPB PHIGHVT L=0.18 W=0.82
+ AD=0.2214 AS=0.148546 PD=2.18 PS=1.21198 NRD=1.182 NRS=30.2986 M=1 R=4.55556
+ SA=90001.8 SB=90000.2 A=0.1476 P=2 MULT=1
MM1025 N_VPWR_M1025_d N_S[2]_M1025_g N_A_1012_265#_M1025_s VPB PHIGHVT L=0.18
+ W=1 AD=0.2 AS=0.27 PD=1.4 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1005 N_A_1361_47#_M1005_d N_S[3]_M1005_g N_VPWR_M1025_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.2 PD=2.54 PS=1.4 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90000.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1013 A_1562_333# N_A_1361_47#_M1013_g N_Z_M1013_s VPB PHIGHVT L=0.18 W=0.82
+ AD=0.148546 AS=0.2214 PD=1.21198 PS=2.18 NRD=30.2986 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.8 A=0.1476 P=2 MULT=1
MM1016 N_VPWR_M1016_d N_D[3]_M1016_g A_1562_333# VPB PHIGHVT L=0.18 W=1 AD=0.175
+ AS=0.181154 PD=1.35 PS=1.47802 NRD=6.8753 NRS=24.8417 M=1 R=5.55556 SA=90000.6
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1003 A_1773_297# N_D[4]_M1003_g N_VPWR_M1016_d VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.175 PD=1.47802 PS=1.35 NRD=24.8417 NRS=6.8753 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1007 N_Z_M1007_d N_A_1840_265#_M1007_g A_1773_297# VPB PHIGHVT L=0.18 W=0.82
+ AD=0.2214 AS=0.148546 PD=2.18 PS=1.21198 NRD=1.182 NRS=30.2986 M=1 R=4.55556
+ SA=90001.8 SB=90000.2 A=0.1476 P=2 MULT=1
MM1038 N_VPWR_M1038_d N_S[4]_M1038_g N_A_1840_265#_M1038_s VPB PHIGHVT L=0.18
+ W=1 AD=0.2 AS=0.27 PD=1.4 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1024 N_A_2189_47#_M1024_d N_S[5]_M1024_g N_VPWR_M1038_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.2 PD=2.54 PS=1.4 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90000.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1030 A_2390_333# N_A_2189_47#_M1030_g N_Z_M1030_s VPB PHIGHVT L=0.18 W=0.82
+ AD=0.148546 AS=0.2214 PD=1.21198 PS=2.18 NRD=30.2986 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.8 A=0.1476 P=2 MULT=1
MM1036 N_VPWR_M1036_d N_D[5]_M1036_g A_2390_333# VPB PHIGHVT L=0.18 W=1 AD=0.175
+ AS=0.181154 PD=1.35 PS=1.47802 NRD=6.8753 NRS=24.8417 M=1 R=5.55556 SA=90000.6
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1017 A_2601_297# N_D[6]_M1017_g N_VPWR_M1036_d VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.175 PD=1.47802 PS=1.35 NRD=24.8417 NRS=6.8753 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1026 N_Z_M1026_d N_A_2668_265#_M1026_g A_2601_297# VPB PHIGHVT L=0.18 W=0.82
+ AD=0.2214 AS=0.148546 PD=2.18 PS=1.21198 NRD=1.182 NRS=30.2986 M=1 R=4.55556
+ SA=90001.8 SB=90000.2 A=0.1476 P=2 MULT=1
MM1034 N_VPWR_M1034_d N_S[6]_M1034_g N_A_2668_265#_M1034_s VPB PHIGHVT L=0.18
+ W=1 AD=0.2 AS=0.27 PD=1.4 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1011 N_A_3017_47#_M1011_d N_S[7]_M1011_g N_VPWR_M1034_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.2 PD=2.54 PS=1.4 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90000.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1045 A_3218_333# N_A_3017_47#_M1045_g N_Z_M1045_s VPB PHIGHVT L=0.18 W=0.82
+ AD=0.148546 AS=0.2214 PD=1.21198 PS=2.18 NRD=30.2986 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.7 A=0.1476 P=2 MULT=1
MM1006 N_VPWR_M1006_d N_D[7]_M1006_g A_3218_333# VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.181154 PD=2.54 PS=1.47802 NRD=0.9653 NRS=24.8417 M=1 R=5.55556 SA=90000.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX48_noxref VNB VPB NWDIODE A=27.927 P=38.01
*
.include "sky130_fd_sc_hdll__muxb8to1_1.pxi.spice"
*
.ends
*
*
