* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__bufbuf_16 A VGND VNB VPB VPWR X
X0 VPWR a_225_47# a_589_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VPWR a_589_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_225_47# a_117_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_589_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 VGND a_589_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 X a_589_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 VGND a_225_47# a_589_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_589_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VPWR a_117_297# a_225_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 a_589_47# a_225_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 X a_589_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_225_47# a_117_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 X a_589_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 a_589_47# a_225_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 X a_589_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_589_47# a_225_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 X a_589_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 X a_589_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_589_47# a_225_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 X a_589_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 X a_589_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_589_47# a_225_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR a_589_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 VPWR a_589_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 X a_589_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 VPWR a_589_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X27 X a_589_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 VGND a_117_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 X a_589_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X30 VPWR a_225_47# a_589_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X31 VGND A a_117_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 X a_589_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 VGND a_589_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 X a_589_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 X a_589_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X36 VGND a_589_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 VPWR a_225_47# a_589_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X38 VGND a_589_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 a_225_47# a_117_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X40 X a_589_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X41 VGND a_589_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X42 VPWR a_589_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X43 VGND a_225_47# a_589_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X44 VGND a_589_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X45 VPWR a_589_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X46 VPWR a_589_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X47 VGND a_589_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X48 a_589_47# a_225_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X49 a_225_47# a_117_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X50 VGND a_225_47# a_589_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X51 VGND a_589_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
