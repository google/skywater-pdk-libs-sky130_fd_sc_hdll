* NGSPICE file created from sky130_fd_sc_hdll__isobufsrc_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__isobufsrc_1 A SLEEP VGND VNB VPB VPWR X
M1000 VGND a_74_47# X VNB nshort w=650000u l=150000u
+  ad=4.23e+11p pd=3.99e+06u as=2.08e+11p ps=1.94e+06u
M1001 a_283_297# SLEEP VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.3e+11p pd=2.46e+06u as=3.288e+11p ps=2.82e+06u
M1002 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_74_47# a_283_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1004 VGND A a_74_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1005 VPWR A a_74_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
.ends

