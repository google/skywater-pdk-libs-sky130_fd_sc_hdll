# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__xor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xor2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 1.075000 0.925000 1.275000 ;
        RECT 0.755000 1.275000 0.925000 1.445000 ;
        RECT 0.755000 1.445000 2.080000 1.615000 ;
        RECT 1.860000 1.075000 3.530000 1.275000 ;
        RECT 1.860000 1.275000 2.080000 1.445000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.105000 1.075000 1.395000 1.120000 ;
        RECT 1.105000 1.120000 4.055000 1.260000 ;
        RECT 1.105000 1.260000 1.395000 1.305000 ;
        RECT 3.765000 1.075000 4.055000 1.120000 ;
        RECT 3.765000 1.260000 4.055000 1.305000 ;
    END
  END B
  PIN VGND
    ANTENNADIFFAREA  1.069250 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  0.925000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  0.806750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.975000 0.645000 4.305000 0.725000 ;
        RECT 3.975000 0.725000 6.350000 0.905000 ;
        RECT 5.385000 0.645000 5.765000 0.725000 ;
        RECT 5.475000 1.415000 6.350000 1.625000 ;
        RECT 5.475000 1.625000 5.725000 2.125000 ;
        RECT 5.985000 0.905000 6.350000 1.415000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.120000  0.725000 1.850000 0.905000 ;
      RECT 0.120000  0.905000 0.290000 1.785000 ;
      RECT 0.120000  1.785000 2.420000 1.955000 ;
      RECT 0.120000  2.135000 0.400000 2.465000 ;
      RECT 0.145000  2.125000 0.315000 2.135000 ;
      RECT 0.190000  0.085000 0.360000 0.555000 ;
      RECT 0.530000  0.255000 0.910000 0.725000 ;
      RECT 0.620000  2.135000 0.870000 2.635000 ;
      RECT 1.090000  2.135000 1.340000 2.295000 ;
      RECT 1.090000  2.295000 2.280000 2.465000 ;
      RECT 1.130000  0.085000 1.300000 0.555000 ;
      RECT 1.145000  1.075000 1.690000 1.275000 ;
      RECT 1.165000  2.125000 1.335000 2.135000 ;
      RECT 1.470000  0.255000 1.850000 0.725000 ;
      RECT 1.560000  1.955000 1.810000 2.125000 ;
      RECT 2.030000  2.135000 2.280000 2.295000 ;
      RECT 2.070000  0.085000 2.240000 0.555000 ;
      RECT 2.250000  1.445000 5.185000 1.615000 ;
      RECT 2.250000  1.615000 2.420000 1.785000 ;
      RECT 2.485000  2.125000 2.800000 2.465000 ;
      RECT 2.510000  0.255000 2.840000 0.725000 ;
      RECT 2.510000  0.725000 3.700000 0.905000 ;
      RECT 2.590000  1.785000 5.255000 1.955000 ;
      RECT 2.590000  1.955000 2.800000 2.125000 ;
      RECT 3.020000  2.135000 3.270000 2.635000 ;
      RECT 3.060000  0.085000 3.230000 0.555000 ;
      RECT 3.400000  0.255000 4.780000 0.475000 ;
      RECT 3.400000  0.475000 3.700000 0.725000 ;
      RECT 3.490000  1.955000 3.740000 2.465000 ;
      RECT 3.720000  1.075000 4.490000 1.275000 ;
      RECT 3.960000  2.135000 4.265000 2.635000 ;
      RECT 4.485000  1.955000 5.255000 2.295000 ;
      RECT 4.485000  2.295000 6.195000 2.465000 ;
      RECT 5.015000  1.075000 5.725000 1.245000 ;
      RECT 5.015000  1.245000 5.185000 1.445000 ;
      RECT 5.045000  0.085000 5.215000 0.555000 ;
      RECT 5.945000  1.795000 6.195000 2.295000 ;
      RECT 5.985000  0.085000 6.155000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.165000  1.105000 1.335000 1.275000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  1.105000 3.995000 1.275000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 0.085000 2.095000 0.375000 2.140000 ;
      RECT 0.085000 2.140000 1.395000 2.280000 ;
      RECT 0.085000 2.280000 0.375000 2.325000 ;
      RECT 1.105000 2.095000 1.395000 2.140000 ;
      RECT 1.105000 2.280000 1.395000 2.325000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor2_2
