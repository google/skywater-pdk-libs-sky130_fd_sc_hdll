* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__and2_6 A B VGND VNB VPB VPWR X
X0 VPWR a_117_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 X a_117_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND a_117_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 X a_117_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR a_117_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 VPWR B a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 X a_117_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 VGND a_117_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X a_117_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_117_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_117_297# A a_293_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND a_117_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 VGND B a_131_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR a_117_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 a_293_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_117_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_131_47# A a_117_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 X a_117_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 X a_117_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
