* File: sky130_fd_sc_hdll__o22ai_1.pex.spice
* Created: Wed Sep  2 08:45:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O22AI_1%B1 1 3 4 6 7 12
r32 12 13 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r33 10 12 33.7665 $w=3.64e-07 $l=2.55e-07 $layer=POLY_cond $X=0.24 $Y=1.202
+ $X2=0.495 $Y2=1.202
r34 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r35 7 11 14.8857 $w=2.38e-07 $l=3.1e-07 $layer=LI1_cond $X=0.205 $Y=0.85
+ $X2=0.205 $Y2=1.16
r36 4 13 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r37 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r38 1 12 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r39 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_1%B2 1 3 4 6 7 11
c36 4 0 3.60226e-19 $X=1.09 $Y=1.41
r37 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.16 $X2=1.14 $Y2=1.16
r38 7 11 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=1.53 $X2=1.2
+ $Y2=1.16
r39 4 10 47.4309 $w=3.07e-07 $l=2.81514e-07 $layer=POLY_cond $X=1.09 $Y=1.41
+ $X2=1.157 $Y2=1.16
r40 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.09 $Y=1.41 $X2=1.09
+ $Y2=1.985
r41 1 10 38.5336 $w=3.07e-07 $l=2.05925e-07 $layer=POLY_cond $X=1.065 $Y=0.995
+ $X2=1.157 $Y2=1.16
r42 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.065 $Y=0.995
+ $X2=1.065 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_1%A2 1 3 4 6 7 8 18 20
c45 18 0 1.62645e-19 $X=2.045 $Y=1.615
c46 8 0 1.97582e-19 $X=1.865 $Y=1.445
r47 18 20 12.444 $w=2.5e-07 $l=2.55e-07 $layer=LI1_cond $X=2.045 $Y=1.615
+ $X2=2.045 $Y2=1.87
r48 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.745
+ $Y=1.16 $X2=1.745 $Y2=1.16
r49 8 18 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.865 $Y=1.53
+ $X2=2.045 $Y2=1.53
r50 7 10 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.865 $Y=1.16
+ $X2=1.745 $Y2=1.16
r51 7 8 10.0212 $w=2.28e-07 $l=2e-07 $layer=LI1_cond $X=1.865 $Y=1.245 $X2=1.865
+ $Y2=1.445
r52 4 11 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=1.83 $Y=1.41
+ $X2=1.77 $Y2=1.16
r53 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.83 $Y=1.41 $X2=1.83
+ $Y2=1.985
r54 1 11 38.578 $w=2.95e-07 $l=1.72337e-07 $layer=POLY_cond $X=1.755 $Y=0.995
+ $X2=1.77 $Y2=1.16
r55 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.755 $Y=0.995
+ $X2=1.755 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_1%A1 1 3 4 6 7 14
r25 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.435
+ $Y=1.16 $X2=2.435 $Y2=1.16
r26 7 14 4.43636 $w=1.98e-07 $l=8e-08 $layer=LI1_cond $X=2.515 $Y=1.175
+ $X2=2.435 $Y2=1.175
r27 4 10 45.1054 $w=3.82e-07 $l=3.02076e-07 $layer=POLY_cond $X=2.24 $Y=1.41
+ $X2=2.355 $Y2=1.16
r28 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.24 $Y=1.41 $X2=2.24
+ $Y2=1.985
r29 1 10 39.2524 $w=3.82e-07 $l=2.24332e-07 $layer=POLY_cond $X=2.215 $Y=0.995
+ $X2=2.355 $Y2=1.16
r30 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.215 $Y=0.995
+ $X2=2.215 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_1%VPWR 1 2 7 9 11 13 17 19 32
r34 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r35 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r36 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r37 23 26 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r38 22 25 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r39 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r40 20 28 3.66972 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r41 20 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r42 19 31 4.67607 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.34 $Y=2.72 $X2=2.55
+ $Y2=2.72
r43 19 25 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.34 $Y=2.72 $X2=2.07
+ $Y2=2.72
r44 17 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r45 17 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r46 13 16 24.4894 $w=3.18e-07 $l=6.8e-07 $layer=LI1_cond $X=2.5 $Y=1.64 $X2=2.5
+ $Y2=2.32
r47 11 31 3.00604 $w=3.2e-07 $l=1.07121e-07 $layer=LI1_cond $X=2.5 $Y=2.635
+ $X2=2.55 $Y2=2.72
r48 11 16 11.3444 $w=3.18e-07 $l=3.15e-07 $layer=LI1_cond $X=2.5 $Y=2.635
+ $X2=2.5 $Y2=2.32
r49 7 28 3.24547 $w=2.1e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.172 $Y2=2.72
r50 7 9 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.24 $Y2=2.34
r51 2 16 400 $w=1.7e-07 $l=9.04599e-07 $layer=licon1_PDIFF $count=1 $X=2.33
+ $Y=1.485 $X2=2.475 $Y2=2.32
r52 2 13 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=2.33
+ $Y=1.485 $X2=2.475 $Y2=1.64
r53 1 9 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_1%Y 1 2 8 9 10 12 15 17
r36 17 20 0.434938 $w=5.48e-07 $l=2e-08 $layer=LI1_cond $X=1.405 $Y=1.94
+ $X2=1.405 $Y2=1.96
r37 15 20 5.43672 $w=5.48e-07 $l=2.5e-07 $layer=LI1_cond $X=1.405 $Y=2.21
+ $X2=1.405 $Y2=1.96
r38 12 14 3.55422 $w=3.98e-07 $l=9.5e-08 $layer=LI1_cond $X=0.695 $Y=0.73
+ $X2=0.695 $Y2=0.825
r39 9 17 6.43462 $w=2.1e-07 $l=2.75e-07 $layer=LI1_cond $X=1.13 $Y=1.94
+ $X2=1.405 $Y2=1.94
r40 9 10 17.9567 $w=2.08e-07 $l=3.4e-07 $layer=LI1_cond $X=1.13 $Y=1.94 $X2=0.79
+ $Y2=1.94
r41 8 10 7.07071 $w=2.1e-07 $l=1.93505e-07 $layer=LI1_cond $X=0.642 $Y=1.835
+ $X2=0.79 $Y2=1.94
r42 8 14 39.4565 $w=2.93e-07 $l=1.01e-06 $layer=LI1_cond $X=0.642 $Y=1.835
+ $X2=0.642 $Y2=0.825
r43 2 20 300 $w=1.7e-07 $l=5.74565e-07 $layer=licon1_PDIFF $count=2 $X=1.18
+ $Y=1.485 $X2=1.4 $Y2=1.96
r44 1 12 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_1%A_27_47# 1 2 3 10 14 15 16 20
r47 18 20 9.0127 $w=3.88e-07 $l=3.05e-07 $layer=LI1_cond $X=2.465 $Y=0.695
+ $X2=2.465 $Y2=0.39
r48 17 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.62 $Y=0.78
+ $X2=1.455 $Y2=0.78
r49 16 18 8.28377 $w=1.7e-07 $l=2.33666e-07 $layer=LI1_cond $X=2.27 $Y=0.78
+ $X2=2.465 $Y2=0.695
r50 16 17 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.27 $Y=0.78
+ $X2=1.62 $Y2=0.78
r51 15 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.455 $Y=0.695
+ $X2=1.455 $Y2=0.78
r52 14 23 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.455 $Y=0.475
+ $X2=1.455 $Y2=0.385
r53 14 15 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.455 $Y=0.475
+ $X2=1.455 $Y2=0.695
r54 10 23 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.29 $Y=0.385
+ $X2=1.455 $Y2=0.385
r55 10 12 63.4646 $w=1.78e-07 $l=1.03e-06 $layer=LI1_cond $X=1.29 $Y=0.385
+ $X2=0.26 $Y2=0.385
r56 3 20 91 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_NDIFF $count=2 $X=2.29
+ $Y=0.235 $X2=2.485 $Y2=0.39
r57 2 25 182 $w=1.7e-07 $l=6.33206e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.235 $X2=1.455 $Y2=0.73
r58 2 23 182 $w=1.7e-07 $l=3.84773e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.235 $X2=1.455 $Y2=0.39
r59 1 12 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_1%VGND 1 6 9 10 11 21 22
r33 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r34 19 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r35 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r36 14 18 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r37 11 19 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r38 11 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r39 9 18 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.61
+ $Y2=0
r40 9 10 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.975
+ $Y2=0
r41 8 21 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.06 $Y=0 $X2=2.53
+ $Y2=0
r42 8 10 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.06 $Y=0 $X2=1.975
+ $Y2=0
r43 4 10 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=0.085
+ $X2=1.975 $Y2=0
r44 4 6 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.975 $Y=0.085
+ $X2=1.975 $Y2=0.36
r45 1 6 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.83
+ $Y=0.235 $X2=1.975 $Y2=0.36
.ends

