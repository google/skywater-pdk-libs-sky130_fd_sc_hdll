# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__and2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and2_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 0.995000 1.535000 1.295000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.615000 1.325000 ;
        RECT 0.435000 1.325000 0.615000 1.465000 ;
        RECT 0.435000 1.465000 1.885000 1.635000 ;
        RECT 1.705000 0.995000 1.965000 1.325000 ;
        RECT 1.705000 1.325000 1.885000 1.465000 ;
    END
  END B
  PIN VGND
    ANTENNADIFFAREA  1.456000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  2.010000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  1.862000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.475000 0.255000 2.745000 0.715000 ;
        RECT 2.475000 0.715000 5.915000 0.885000 ;
        RECT 2.475000 1.445000 5.915000 1.615000 ;
        RECT 2.475000 1.615000 2.745000 2.465000 ;
        RECT 3.415000 0.255000 3.685000 0.715000 ;
        RECT 3.415000 1.615000 3.685000 2.465000 ;
        RECT 4.355000 0.255000 4.625000 0.715000 ;
        RECT 4.355000 1.615000 4.625000 2.465000 ;
        RECT 5.295000 0.255000 5.565000 0.715000 ;
        RECT 5.295000 1.615000 5.565000 2.465000 ;
        RECT 5.495000 0.885000 5.915000 1.445000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.825000 ;
      RECT 0.095000  1.805000 0.395000 2.635000 ;
      RECT 0.565000  1.805000 2.305000 1.975000 ;
      RECT 0.565000  1.975000 0.865000 2.465000 ;
      RECT 1.015000  0.255000 1.345000 0.655000 ;
      RECT 1.015000  0.655000 2.305000 0.825000 ;
      RECT 1.035000  2.145000 1.365000 2.635000 ;
      RECT 1.535000  1.975000 1.805000 2.465000 ;
      RECT 1.940000  0.085000 2.270000 0.485000 ;
      RECT 1.975000  2.160000 2.305000 2.635000 ;
      RECT 2.135000  0.825000 2.305000 1.055000 ;
      RECT 2.135000  1.055000 5.325000 1.265000 ;
      RECT 2.135000  1.265000 2.305000 1.805000 ;
      RECT 2.915000  0.085000 3.245000 0.545000 ;
      RECT 2.915000  1.785000 3.245000 2.635000 ;
      RECT 3.855000  0.085000 4.185000 0.545000 ;
      RECT 3.855000  1.785000 4.185000 2.635000 ;
      RECT 4.795000  0.085000 5.125000 0.545000 ;
      RECT 4.795000  1.785000 5.125000 2.635000 ;
      RECT 5.735000  0.085000 6.065000 0.545000 ;
      RECT 5.735000  1.785000 6.065000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2_8
