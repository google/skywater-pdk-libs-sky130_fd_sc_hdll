* File: sky130_fd_sc_hdll__o2bb2a_2.pxi.spice
* Created: Thu Aug 27 19:21:49 2020
* 
x_PM_SKY130_FD_SC_HDLL__O2BB2A_2%A_84_21# N_A_84_21#_M1004_s N_A_84_21#_M1005_d
+ N_A_84_21#_c_82_n N_A_84_21#_M1003_g N_A_84_21#_c_90_n N_A_84_21#_M1007_g
+ N_A_84_21#_c_83_n N_A_84_21#_M1011_g N_A_84_21#_c_91_n N_A_84_21#_M1013_g
+ N_A_84_21#_c_84_n N_A_84_21#_c_93_n N_A_84_21#_c_106_p N_A_84_21#_c_148_p
+ N_A_84_21#_c_85_n N_A_84_21#_c_95_n N_A_84_21#_c_86_n N_A_84_21#_c_87_n
+ N_A_84_21#_c_88_n N_A_84_21#_c_96_n N_A_84_21#_c_89_n
+ PM_SKY130_FD_SC_HDLL__O2BB2A_2%A_84_21#
x_PM_SKY130_FD_SC_HDLL__O2BB2A_2%A1_N N_A1_N_M1012_g N_A1_N_c_203_n
+ N_A1_N_c_204_n N_A1_N_M1001_g A1_N N_A1_N_c_202_n A1_N
+ PM_SKY130_FD_SC_HDLL__O2BB2A_2%A1_N
x_PM_SKY130_FD_SC_HDLL__O2BB2A_2%A2_N N_A2_N_M1000_g N_A2_N_c_242_n
+ N_A2_N_c_247_n N_A2_N_M1008_g A2_N N_A2_N_c_243_n N_A2_N_c_244_n A2_N
+ PM_SKY130_FD_SC_HDLL__O2BB2A_2%A2_N
x_PM_SKY130_FD_SC_HDLL__O2BB2A_2%A_321_369# N_A_321_369#_M1000_d
+ N_A_321_369#_M1001_d N_A_321_369#_c_288_n N_A_321_369#_M1005_g
+ N_A_321_369#_M1004_g N_A_321_369#_c_290_n N_A_321_369#_c_291_n
+ N_A_321_369#_c_292_n N_A_321_369#_c_286_n N_A_321_369#_c_293_n
+ N_A_321_369#_c_287_n PM_SKY130_FD_SC_HDLL__O2BB2A_2%A_321_369#
x_PM_SKY130_FD_SC_HDLL__O2BB2A_2%B2 N_B2_c_357_n N_B2_c_358_n N_B2_M1009_g
+ N_B2_M1010_g N_B2_c_355_n B2 B2 N_B2_c_356_n B2 N_B2_c_361_n B2
+ PM_SKY130_FD_SC_HDLL__O2BB2A_2%B2
x_PM_SKY130_FD_SC_HDLL__O2BB2A_2%B1 N_B1_M1002_g N_B1_c_408_n N_B1_c_409_n
+ N_B1_M1006_g B1 B1 N_B1_c_407_n B1 PM_SKY130_FD_SC_HDLL__O2BB2A_2%B1
x_PM_SKY130_FD_SC_HDLL__O2BB2A_2%VPWR N_VPWR_M1007_d N_VPWR_M1013_d
+ N_VPWR_M1008_d N_VPWR_M1006_d N_VPWR_c_436_n N_VPWR_c_437_n N_VPWR_c_438_n
+ N_VPWR_c_439_n N_VPWR_c_440_n VPWR N_VPWR_c_441_n N_VPWR_c_442_n
+ N_VPWR_c_443_n N_VPWR_c_444_n N_VPWR_c_445_n N_VPWR_c_435_n VPWR
+ PM_SKY130_FD_SC_HDLL__O2BB2A_2%VPWR
x_PM_SKY130_FD_SC_HDLL__O2BB2A_2%X N_X_M1003_d N_X_M1007_s N_X_c_499_n
+ N_X_c_502_n N_X_c_497_n X N_X_c_514_n PM_SKY130_FD_SC_HDLL__O2BB2A_2%X
x_PM_SKY130_FD_SC_HDLL__O2BB2A_2%VGND N_VGND_M1003_s N_VGND_M1011_s
+ N_VGND_M1010_d N_VGND_c_530_n N_VGND_c_531_n N_VGND_c_532_n N_VGND_c_533_n
+ N_VGND_c_534_n N_VGND_c_535_n N_VGND_c_536_n VGND N_VGND_c_537_n
+ N_VGND_c_538_n N_VGND_c_539_n VGND PM_SKY130_FD_SC_HDLL__O2BB2A_2%VGND
x_PM_SKY130_FD_SC_HDLL__O2BB2A_2%A_627_47# N_A_627_47#_M1004_d
+ N_A_627_47#_M1002_d N_A_627_47#_c_590_n N_A_627_47#_c_591_n
+ N_A_627_47#_c_592_n N_A_627_47#_c_593_n
+ PM_SKY130_FD_SC_HDLL__O2BB2A_2%A_627_47#
cc_1 VNB N_A_84_21#_c_82_n 0.0213429f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.995
cc_2 VNB N_A_84_21#_c_83_n 0.017609f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=0.995
cc_3 VNB N_A_84_21#_c_84_n 0.00380342f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.16
cc_4 VNB N_A_84_21#_c_85_n 5.1593e-19 $X=-0.19 $Y=-0.24 $X2=2.915 $Y2=1.495
cc_5 VNB N_A_84_21#_c_86_n 0.00199768f $X=-0.19 $Y=-0.24 $X2=2.82 $Y2=0.485
cc_6 VNB N_A_84_21#_c_87_n 0.00745463f $X=-0.19 $Y=-0.24 $X2=2.905 $Y2=1.075
cc_7 VNB N_A_84_21#_c_88_n 0.00179548f $X=-0.19 $Y=-0.24 $X2=2.905 $Y2=1.245
cc_8 VNB N_A_84_21#_c_89_n 0.0560668f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.202
cc_9 VNB N_A1_N_M1012_g 0.0309113f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB A1_N 0.009648f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.41
cc_11 VNB N_A1_N_c_202_n 0.023201f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=0.995
cc_12 VNB N_A2_N_c_242_n 0.012989f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A2_N_c_243_n 0.0365109f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.985
cc_14 VNB N_A2_N_c_244_n 0.0209173f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=0.56
cc_15 VNB A2_N 0.00714943f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.985
cc_16 VNB N_A_321_369#_M1004_g 0.05428f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.985
cc_17 VNB N_A_321_369#_c_286_n 0.00382046f $X=-0.19 $Y=-0.24 $X2=1.035 $Y2=1.16
cc_18 VNB N_A_321_369#_c_287_n 0.014905f $X=-0.19 $Y=-0.24 $X2=2.895 $Y2=1.075
cc_19 VNB N_B2_M1010_g 0.0288584f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.56
cc_20 VNB N_B2_c_355_n 0.00551982f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.985
cc_21 VNB N_B2_c_356_n 0.0229754f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.985
cc_22 VNB N_B1_M1002_g 0.0362863f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB B1 0.0115713f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.41
cc_24 VNB N_B1_c_407_n 0.0371145f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.985
cc_25 VNB N_VPWR_c_435_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_X_c_497_n 0.00106626f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=0.56
cc_27 VNB N_VGND_c_530_n 0.0106114f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.41
cc_28 VNB N_VGND_c_531_n 0.0341371f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.985
cc_29 VNB N_VGND_c_532_n 0.0205922f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=0.56
cc_30 VNB N_VGND_c_533_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.985
cc_31 VNB N_VGND_c_534_n 0.00470034f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.16
cc_32 VNB N_VGND_c_535_n 0.0636011f $X=-0.19 $Y=-0.24 $X2=1.285 $Y2=1.885
cc_33 VNB N_VGND_c_536_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=2.83 $Y2=1.97
cc_34 VNB N_VGND_c_537_n 0.0223141f $X=-0.19 $Y=-0.24 $X2=2.82 $Y2=0.485
cc_35 VNB N_VGND_c_538_n 0.24966f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_539_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=3.27 $Y2=2
cc_37 VNB N_A_627_47#_c_590_n 0.00120906f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.56
cc_38 VNB N_A_627_47#_c_591_n 0.0204136f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.985
cc_39 VNB N_A_627_47#_c_592_n 0.003732f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.985
cc_40 VNB N_A_627_47#_c_593_n 0.0164847f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=0.56
cc_41 VPB N_A_84_21#_c_90_n 0.018801f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.41
cc_42 VPB N_A_84_21#_c_91_n 0.0158373f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.41
cc_43 VPB N_A_84_21#_c_84_n 0.00146886f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.16
cc_44 VPB N_A_84_21#_c_93_n 0.0019007f $X=-0.19 $Y=1.305 $X2=1.285 $Y2=1.885
cc_45 VPB N_A_84_21#_c_85_n 4.37229e-19 $X=-0.19 $Y=1.305 $X2=2.915 $Y2=1.495
cc_46 VPB N_A_84_21#_c_95_n 0.0066444f $X=-0.19 $Y=1.305 $X2=1.285 $Y2=1.53
cc_47 VPB N_A_84_21#_c_96_n 0.00719069f $X=-0.19 $Y=1.305 $X2=3.132 $Y2=1.97
cc_48 VPB N_A_84_21#_c_89_n 0.0283171f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.202
cc_49 VPB N_A1_N_c_203_n 0.0215623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A1_N_c_204_n 0.0248325f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=0.995
cc_51 VPB N_A1_N_c_202_n 0.00431928f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=0.995
cc_52 VPB N_A2_N_c_242_n 0.0205577f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A2_N_c_247_n 0.0283773f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_321_369#_c_288_n 0.0194971f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=0.995
cc_55 VPB N_A_321_369#_M1004_g 0.00307141f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.985
cc_56 VPB N_A_321_369#_c_290_n 0.0502722f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=0.56
cc_57 VPB N_A_321_369#_c_291_n 0.0194444f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=0.56
cc_58 VPB N_A_321_369#_c_292_n 0.00965838f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.41
cc_59 VPB N_A_321_369#_c_293_n 0.00803699f $X=-0.19 $Y=1.305 $X2=1.37 $Y2=1.97
cc_60 VPB N_A_321_369#_c_287_n 8.61122e-19 $X=-0.19 $Y=1.305 $X2=2.895 $Y2=1.075
cc_61 VPB N_B2_c_357_n 0.0200365f $X=-0.19 $Y=1.305 $X2=3.125 $Y2=1.845
cc_62 VPB N_B2_c_358_n 0.0230986f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_B2_c_355_n 0.00157619f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.985
cc_64 VPB N_B2_c_356_n 0.00498286f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.985
cc_65 VPB N_B2_c_361_n 0.00938631f $X=-0.19 $Y=1.305 $X2=2.83 $Y2=1.97
cc_66 VPB N_B1_c_408_n 0.0246416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_B1_c_409_n 0.0307014f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=0.995
cc_68 VPB B1 0.0173304f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.41
cc_69 VPB N_B1_c_407_n 0.00828342f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.985
cc_70 VPB N_VPWR_c_436_n 0.0105855f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=0.995
cc_71 VPB N_VPWR_c_437_n 0.0490932f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=0.56
cc_72 VPB N_VPWR_c_438_n 0.0027905f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.16
cc_73 VPB N_VPWR_c_439_n 0.0120619f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_440_n 0.0350731f $X=-0.19 $Y=1.305 $X2=1.285 $Y2=1.885
cc_75 VPB N_VPWR_c_441_n 0.0164234f $X=-0.19 $Y=1.305 $X2=2.895 $Y2=1.075
cc_76 VPB N_VPWR_c_442_n 0.0267798f $X=-0.19 $Y=1.305 $X2=1.285 $Y2=1.53
cc_77 VPB N_VPWR_c_443_n 0.0369579f $X=-0.19 $Y=1.305 $X2=2.857 $Y2=0.69
cc_78 VPB N_VPWR_c_444_n 0.005797f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_445_n 0.0138739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_435_n 0.0449522f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_X_c_497_n 9.46957e-19 $X=-0.19 $Y=1.305 $X2=0.965 $Y2=0.56
cc_82 N_A_84_21#_c_83_n N_A1_N_M1012_g 0.016001f $X=0.965 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A_84_21#_c_91_n N_A1_N_c_203_n 0.0109099f $X=0.99 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_84_21#_c_84_n N_A1_N_c_203_n 0.00238776f $X=1.01 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_84_21#_c_93_n N_A1_N_c_203_n 0.00221821f $X=1.285 $Y=1.885 $X2=0 $Y2=0
cc_86 N_A_84_21#_c_95_n N_A1_N_c_203_n 0.00255969f $X=1.285 $Y=1.53 $X2=0 $Y2=0
cc_87 N_A_84_21#_c_89_n N_A1_N_c_203_n 0.00292843f $X=0.99 $Y=1.202 $X2=0 $Y2=0
cc_88 N_A_84_21#_c_91_n N_A1_N_c_204_n 0.0210246f $X=0.99 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A_84_21#_c_93_n N_A1_N_c_204_n 0.00205417f $X=1.285 $Y=1.885 $X2=0 $Y2=0
cc_90 N_A_84_21#_c_106_p N_A1_N_c_204_n 0.0156443f $X=2.83 $Y=1.97 $X2=0 $Y2=0
cc_91 N_A_84_21#_c_84_n A1_N 0.0158819f $X=1.01 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_84_21#_c_106_p A1_N 0.00357405f $X=2.83 $Y=1.97 $X2=0 $Y2=0
cc_93 N_A_84_21#_c_95_n A1_N 0.00419335f $X=1.285 $Y=1.53 $X2=0 $Y2=0
cc_94 N_A_84_21#_c_89_n A1_N 0.00146165f $X=0.99 $Y=1.202 $X2=0 $Y2=0
cc_95 N_A_84_21#_c_84_n N_A1_N_c_202_n 0.00102326f $X=1.01 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_84_21#_c_89_n N_A1_N_c_202_n 0.0214157f $X=0.99 $Y=1.202 $X2=0 $Y2=0
cc_97 N_A_84_21#_c_106_p N_A2_N_c_247_n 0.0163557f $X=2.83 $Y=1.97 $X2=0 $Y2=0
cc_98 N_A_84_21#_c_96_n N_A2_N_c_247_n 0.00397768f $X=3.132 $Y=1.97 $X2=0 $Y2=0
cc_99 N_A_84_21#_c_83_n A2_N 7.29046e-19 $X=0.965 $Y=0.995 $X2=0 $Y2=0
cc_100 N_A_84_21#_c_106_p N_A_321_369#_M1001_d 0.00963598f $X=2.83 $Y=1.97 $X2=0
+ $Y2=0
cc_101 N_A_84_21#_c_96_n N_A_321_369#_c_288_n 0.0273046f $X=3.132 $Y=1.97 $X2=0
+ $Y2=0
cc_102 N_A_84_21#_c_85_n N_A_321_369#_M1004_g 0.0032526f $X=2.915 $Y=1.495 $X2=0
+ $Y2=0
cc_103 N_A_84_21#_c_86_n N_A_321_369#_M1004_g 0.00983659f $X=2.82 $Y=0.485 $X2=0
+ $Y2=0
cc_104 N_A_84_21#_c_88_n N_A_321_369#_M1004_g 0.00546478f $X=2.905 $Y=1.245
+ $X2=0 $Y2=0
cc_105 N_A_84_21#_c_106_p N_A_321_369#_c_290_n 0.00743538f $X=2.83 $Y=1.97 $X2=0
+ $Y2=0
cc_106 N_A_84_21#_c_85_n N_A_321_369#_c_290_n 0.00572493f $X=2.915 $Y=1.495
+ $X2=0 $Y2=0
cc_107 N_A_84_21#_c_86_n N_A_321_369#_c_290_n 0.00182253f $X=2.82 $Y=0.485 $X2=0
+ $Y2=0
cc_108 N_A_84_21#_c_88_n N_A_321_369#_c_290_n 6.14215e-19 $X=2.905 $Y=1.245
+ $X2=0 $Y2=0
cc_109 N_A_84_21#_c_96_n N_A_321_369#_c_290_n 0.00669585f $X=3.132 $Y=1.97 $X2=0
+ $Y2=0
cc_110 N_A_84_21#_c_85_n N_A_321_369#_c_291_n 0.00449656f $X=2.915 $Y=1.495
+ $X2=0 $Y2=0
cc_111 N_A_84_21#_c_96_n N_A_321_369#_c_291_n 0.0170389f $X=3.132 $Y=1.97 $X2=0
+ $Y2=0
cc_112 N_A_84_21#_c_93_n N_A_321_369#_c_292_n 0.0078685f $X=1.285 $Y=1.885 $X2=0
+ $Y2=0
cc_113 N_A_84_21#_c_106_p N_A_321_369#_c_292_n 0.0563007f $X=2.83 $Y=1.97 $X2=0
+ $Y2=0
cc_114 N_A_84_21#_c_95_n N_A_321_369#_c_292_n 0.0101775f $X=1.285 $Y=1.53 $X2=0
+ $Y2=0
cc_115 N_A_84_21#_c_86_n N_A_321_369#_c_286_n 0.0141488f $X=2.82 $Y=0.485 $X2=0
+ $Y2=0
cc_116 N_A_84_21#_c_106_p N_A_321_369#_c_293_n 0.0214628f $X=2.83 $Y=1.97 $X2=0
+ $Y2=0
cc_117 N_A_84_21#_c_85_n N_A_321_369#_c_293_n 0.00979025f $X=2.915 $Y=1.495
+ $X2=0 $Y2=0
cc_118 N_A_84_21#_c_96_n N_A_321_369#_c_293_n 0.0173771f $X=3.132 $Y=1.97 $X2=0
+ $Y2=0
cc_119 N_A_84_21#_c_85_n N_A_321_369#_c_287_n 0.00602699f $X=2.915 $Y=1.495
+ $X2=0 $Y2=0
cc_120 N_A_84_21#_c_86_n N_A_321_369#_c_287_n 0.00951384f $X=2.82 $Y=0.485 $X2=0
+ $Y2=0
cc_121 N_A_84_21#_c_87_n N_A_321_369#_c_287_n 0.032417f $X=2.905 $Y=1.075 $X2=0
+ $Y2=0
cc_122 N_A_84_21#_c_85_n N_B2_c_357_n 5.39947e-19 $X=2.915 $Y=1.495 $X2=0 $Y2=0
cc_123 N_A_84_21#_c_96_n N_B2_c_357_n 0.00427294f $X=3.132 $Y=1.97 $X2=0 $Y2=0
cc_124 N_A_84_21#_c_96_n N_B2_c_358_n 0.00339757f $X=3.132 $Y=1.97 $X2=0 $Y2=0
cc_125 N_A_84_21#_c_88_n N_B2_c_355_n 0.0163886f $X=2.905 $Y=1.245 $X2=0 $Y2=0
cc_126 N_A_84_21#_c_96_n N_B2_c_355_n 0.0183257f $X=3.132 $Y=1.97 $X2=0 $Y2=0
cc_127 N_A_84_21#_c_88_n N_B2_c_356_n 2.03161e-19 $X=2.905 $Y=1.245 $X2=0 $Y2=0
cc_128 N_A_84_21#_c_96_n N_B2_c_356_n 0.00139774f $X=3.132 $Y=1.97 $X2=0 $Y2=0
cc_129 N_A_84_21#_c_85_n N_B2_c_361_n 0.00427743f $X=2.915 $Y=1.495 $X2=0 $Y2=0
cc_130 N_A_84_21#_c_96_n N_B2_c_361_n 0.0441356f $X=3.132 $Y=1.97 $X2=0 $Y2=0
cc_131 N_A_84_21#_c_93_n N_VPWR_M1013_d 0.00424463f $X=1.285 $Y=1.885 $X2=0
+ $Y2=0
cc_132 N_A_84_21#_c_148_p N_VPWR_M1013_d 0.00422188f $X=1.37 $Y=1.97 $X2=0 $Y2=0
cc_133 N_A_84_21#_c_95_n N_VPWR_M1013_d 0.0021597f $X=1.285 $Y=1.53 $X2=0 $Y2=0
cc_134 N_A_84_21#_c_106_p N_VPWR_M1008_d 0.0160599f $X=2.83 $Y=1.97 $X2=0 $Y2=0
cc_135 N_A_84_21#_c_96_n N_VPWR_M1008_d 0.00188802f $X=3.132 $Y=1.97 $X2=0 $Y2=0
cc_136 N_A_84_21#_c_90_n N_VPWR_c_437_n 0.00791237f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A_84_21#_c_90_n N_VPWR_c_438_n 5.09998e-19 $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_84_21#_c_91_n N_VPWR_c_438_n 0.0108783f $X=0.99 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_84_21#_c_148_p N_VPWR_c_438_n 0.0131715f $X=1.37 $Y=1.97 $X2=0 $Y2=0
cc_140 N_A_84_21#_c_95_n N_VPWR_c_438_n 0.00369081f $X=1.285 $Y=1.53 $X2=0 $Y2=0
cc_141 N_A_84_21#_c_90_n N_VPWR_c_441_n 0.00590121f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_84_21#_c_91_n N_VPWR_c_441_n 0.00427505f $X=0.99 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_84_21#_c_106_p N_VPWR_c_442_n 0.0139796f $X=2.83 $Y=1.97 $X2=0 $Y2=0
cc_144 N_A_84_21#_c_106_p N_VPWR_c_443_n 0.00105858f $X=2.83 $Y=1.97 $X2=0 $Y2=0
cc_145 N_A_84_21#_c_96_n N_VPWR_c_443_n 0.0221356f $X=3.132 $Y=1.97 $X2=0 $Y2=0
cc_146 N_A_84_21#_c_106_p N_VPWR_c_445_n 0.0295056f $X=2.83 $Y=1.97 $X2=0 $Y2=0
cc_147 N_A_84_21#_c_96_n N_VPWR_c_445_n 0.0106951f $X=3.132 $Y=1.97 $X2=0 $Y2=0
cc_148 N_A_84_21#_M1005_d N_VPWR_c_435_n 0.0024999f $X=3.125 $Y=1.845 $X2=0
+ $Y2=0
cc_149 N_A_84_21#_c_90_n N_VPWR_c_435_n 0.0107561f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_84_21#_c_91_n N_VPWR_c_435_n 0.00732977f $X=0.99 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_84_21#_c_106_p N_VPWR_c_435_n 0.0287395f $X=2.83 $Y=1.97 $X2=0 $Y2=0
cc_152 N_A_84_21#_c_148_p N_VPWR_c_435_n 7.95799e-19 $X=1.37 $Y=1.97 $X2=0 $Y2=0
cc_153 N_A_84_21#_c_96_n N_VPWR_c_435_n 0.0201321f $X=3.132 $Y=1.97 $X2=0 $Y2=0
cc_154 N_A_84_21#_c_82_n N_X_c_499_n 0.00674407f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_84_21#_c_83_n N_X_c_499_n 0.00886912f $X=0.965 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A_84_21#_c_89_n N_X_c_499_n 0.00194336f $X=0.99 $Y=1.202 $X2=0 $Y2=0
cc_157 N_A_84_21#_c_90_n N_X_c_502_n 0.00225529f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_84_21#_c_93_n N_X_c_502_n 0.00391171f $X=1.285 $Y=1.885 $X2=0 $Y2=0
cc_159 N_A_84_21#_c_148_p N_X_c_502_n 0.008241f $X=1.37 $Y=1.97 $X2=0 $Y2=0
cc_160 N_A_84_21#_c_89_n N_X_c_502_n 0.00281092f $X=0.99 $Y=1.202 $X2=0 $Y2=0
cc_161 N_A_84_21#_c_82_n N_X_c_497_n 0.00549578f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_84_21#_c_90_n N_X_c_497_n 0.00835766f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A_84_21#_c_83_n N_X_c_497_n 0.00366888f $X=0.965 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_84_21#_c_91_n N_X_c_497_n 0.00289211f $X=0.99 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A_84_21#_c_84_n N_X_c_497_n 0.0321643f $X=1.01 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_84_21#_c_93_n N_X_c_497_n 0.0065201f $X=1.285 $Y=1.885 $X2=0 $Y2=0
cc_167 N_A_84_21#_c_95_n N_X_c_497_n 0.0130579f $X=1.285 $Y=1.53 $X2=0 $Y2=0
cc_168 N_A_84_21#_c_89_n N_X_c_497_n 0.0351273f $X=0.99 $Y=1.202 $X2=0 $Y2=0
cc_169 N_A_84_21#_c_90_n N_X_c_514_n 0.00829631f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_84_21#_c_82_n N_VGND_c_531_n 0.00501374f $X=0.495 $Y=0.995 $X2=0
+ $Y2=0
cc_171 N_A_84_21#_c_82_n N_VGND_c_532_n 0.00533769f $X=0.495 $Y=0.995 $X2=0
+ $Y2=0
cc_172 N_A_84_21#_c_83_n N_VGND_c_532_n 0.00541359f $X=0.965 $Y=0.995 $X2=0
+ $Y2=0
cc_173 N_A_84_21#_c_83_n N_VGND_c_533_n 0.00511555f $X=0.965 $Y=0.995 $X2=0
+ $Y2=0
cc_174 N_A_84_21#_c_84_n N_VGND_c_533_n 5.1142e-19 $X=1.01 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_84_21#_c_89_n N_VGND_c_533_n 0.00215169f $X=0.99 $Y=1.202 $X2=0 $Y2=0
cc_176 N_A_84_21#_c_86_n N_VGND_c_535_n 0.0106665f $X=2.82 $Y=0.485 $X2=0 $Y2=0
cc_177 N_A_84_21#_M1004_s N_VGND_c_538_n 0.00402485f $X=2.695 $Y=0.235 $X2=0
+ $Y2=0
cc_178 N_A_84_21#_c_82_n N_VGND_c_538_n 0.0104335f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_84_21#_c_83_n N_VGND_c_538_n 0.0100908f $X=0.965 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_84_21#_c_86_n N_VGND_c_538_n 0.00899799f $X=2.82 $Y=0.485 $X2=0 $Y2=0
cc_181 N_A_84_21#_c_86_n N_A_627_47#_c_590_n 0.0147414f $X=2.82 $Y=0.485 $X2=0
+ $Y2=0
cc_182 N_A_84_21#_c_87_n N_A_627_47#_c_592_n 0.0124676f $X=2.905 $Y=1.075 $X2=0
+ $Y2=0
cc_183 N_A_84_21#_c_96_n N_A_627_47#_c_592_n 5.82402e-19 $X=3.132 $Y=1.97 $X2=0
+ $Y2=0
cc_184 N_A1_N_c_203_n N_A2_N_c_242_n 0.00691657f $X=1.515 $Y=1.67 $X2=0 $Y2=0
cc_185 A1_N N_A2_N_c_242_n 0.00195818f $X=1.525 $Y=1.095 $X2=0 $Y2=0
cc_186 N_A1_N_c_202_n N_A2_N_c_242_n 0.00944382f $X=1.55 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A1_N_c_204_n N_A2_N_c_247_n 0.0327653f $X=1.515 $Y=1.77 $X2=0 $Y2=0
cc_188 N_A1_N_c_202_n N_A2_N_c_243_n 0.00700696f $X=1.55 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A1_N_M1012_g N_A2_N_c_244_n 0.027093f $X=1.49 $Y=0.445 $X2=0 $Y2=0
cc_190 N_A1_N_M1012_g A2_N 0.0169278f $X=1.49 $Y=0.445 $X2=0 $Y2=0
cc_191 A1_N A2_N 0.0272498f $X=1.525 $Y=1.095 $X2=0 $Y2=0
cc_192 N_A1_N_c_202_n A2_N 0.00506381f $X=1.55 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A1_N_c_203_n N_A_321_369#_c_292_n 0.00648471f $X=1.515 $Y=1.67 $X2=0
+ $Y2=0
cc_194 N_A1_N_c_204_n N_A_321_369#_c_292_n 0.00231468f $X=1.515 $Y=1.77 $X2=0
+ $Y2=0
cc_195 A1_N N_A_321_369#_c_292_n 0.0178762f $X=1.525 $Y=1.095 $X2=0 $Y2=0
cc_196 N_A1_N_c_202_n N_A_321_369#_c_292_n 0.00278096f $X=1.55 $Y=1.16 $X2=0
+ $Y2=0
cc_197 A1_N N_A_321_369#_c_287_n 0.00620734f $X=1.525 $Y=1.095 $X2=0 $Y2=0
cc_198 N_A1_N_c_204_n N_VPWR_c_438_n 0.00449935f $X=1.515 $Y=1.77 $X2=0 $Y2=0
cc_199 N_A1_N_c_204_n N_VPWR_c_442_n 0.00515358f $X=1.515 $Y=1.77 $X2=0 $Y2=0
cc_200 N_A1_N_c_204_n N_VPWR_c_435_n 0.00725759f $X=1.515 $Y=1.77 $X2=0 $Y2=0
cc_201 N_A1_N_M1012_g N_X_c_499_n 3.70255e-19 $X=1.49 $Y=0.445 $X2=0 $Y2=0
cc_202 N_A1_N_M1012_g N_VGND_c_533_n 0.00720949f $X=1.49 $Y=0.445 $X2=0 $Y2=0
cc_203 N_A1_N_M1012_g N_VGND_c_535_n 0.00524503f $X=1.49 $Y=0.445 $X2=0 $Y2=0
cc_204 N_A1_N_M1012_g N_VGND_c_538_n 0.00973453f $X=1.49 $Y=0.445 $X2=0 $Y2=0
cc_205 N_A2_N_c_243_n N_A_321_369#_M1004_g 0.00280896f $X=2.09 $Y=0.935 $X2=0
+ $Y2=0
cc_206 N_A2_N_c_242_n N_A_321_369#_c_290_n 0.0201825f $X=2.125 $Y=1.67 $X2=0
+ $Y2=0
cc_207 N_A2_N_c_247_n N_A_321_369#_c_291_n 8.73107e-19 $X=2.125 $Y=1.77 $X2=0
+ $Y2=0
cc_208 N_A2_N_c_242_n N_A_321_369#_c_292_n 0.011421f $X=2.125 $Y=1.67 $X2=0
+ $Y2=0
cc_209 N_A2_N_c_247_n N_A_321_369#_c_292_n 0.00465586f $X=2.125 $Y=1.77 $X2=0
+ $Y2=0
cc_210 N_A2_N_c_243_n N_A_321_369#_c_292_n 0.00305969f $X=2.09 $Y=0.935 $X2=0
+ $Y2=0
cc_211 A2_N N_A_321_369#_c_292_n 0.0135342f $X=1.64 $Y=0.51 $X2=0 $Y2=0
cc_212 N_A2_N_c_243_n N_A_321_369#_c_286_n 0.00251225f $X=2.09 $Y=0.935 $X2=0
+ $Y2=0
cc_213 N_A2_N_c_244_n N_A_321_369#_c_286_n 0.00299986f $X=2.11 $Y=0.77 $X2=0
+ $Y2=0
cc_214 A2_N N_A_321_369#_c_286_n 0.0242556f $X=1.64 $Y=0.51 $X2=0 $Y2=0
cc_215 N_A2_N_c_242_n N_A_321_369#_c_293_n 2.08609e-19 $X=2.125 $Y=1.67 $X2=0
+ $Y2=0
cc_216 N_A2_N_c_242_n N_A_321_369#_c_287_n 0.0101503f $X=2.125 $Y=1.67 $X2=0
+ $Y2=0
cc_217 N_A2_N_c_243_n N_A_321_369#_c_287_n 0.00392576f $X=2.09 $Y=0.935 $X2=0
+ $Y2=0
cc_218 N_A2_N_c_244_n N_A_321_369#_c_287_n 0.0021185f $X=2.11 $Y=0.77 $X2=0
+ $Y2=0
cc_219 A2_N N_A_321_369#_c_287_n 0.0342232f $X=1.64 $Y=0.51 $X2=0 $Y2=0
cc_220 N_A2_N_c_247_n N_VPWR_c_442_n 0.00515358f $X=2.125 $Y=1.77 $X2=0 $Y2=0
cc_221 N_A2_N_c_247_n N_VPWR_c_445_n 0.0138479f $X=2.125 $Y=1.77 $X2=0 $Y2=0
cc_222 N_A2_N_c_247_n N_VPWR_c_435_n 0.00859375f $X=2.125 $Y=1.77 $X2=0 $Y2=0
cc_223 A2_N N_X_c_499_n 0.00213193f $X=1.64 $Y=0.51 $X2=0 $Y2=0
cc_224 A2_N N_VGND_c_533_n 0.0231205f $X=1.64 $Y=0.51 $X2=0 $Y2=0
cc_225 N_A2_N_c_244_n N_VGND_c_535_n 0.00424763f $X=2.11 $Y=0.77 $X2=0 $Y2=0
cc_226 A2_N N_VGND_c_535_n 0.0151937f $X=1.64 $Y=0.51 $X2=0 $Y2=0
cc_227 N_A2_N_c_244_n N_VGND_c_538_n 0.00758555f $X=2.11 $Y=0.77 $X2=0 $Y2=0
cc_228 A2_N N_VGND_c_538_n 0.01704f $X=1.64 $Y=0.51 $X2=0 $Y2=0
cc_229 A2_N A_313_47# 0.00741641f $X=1.64 $Y=0.51 $X2=-0.19 $Y2=-0.24
cc_230 N_A_321_369#_M1004_g N_B2_c_357_n 0.00976325f $X=3.06 $Y=0.445 $X2=0
+ $Y2=0
cc_231 N_A_321_369#_c_288_n N_B2_c_358_n 0.0088055f $X=3.035 $Y=1.77 $X2=0 $Y2=0
cc_232 N_A_321_369#_c_291_n N_B2_c_358_n 0.00976325f $X=3.035 $Y=1.562 $X2=0
+ $Y2=0
cc_233 N_A_321_369#_M1004_g N_B2_M1010_g 0.0180943f $X=3.06 $Y=0.445 $X2=0 $Y2=0
cc_234 N_A_321_369#_M1004_g N_B2_c_355_n 0.00191788f $X=3.06 $Y=0.445 $X2=0
+ $Y2=0
cc_235 N_A_321_369#_M1004_g N_B2_c_356_n 0.0177879f $X=3.06 $Y=0.445 $X2=0 $Y2=0
cc_236 N_A_321_369#_c_288_n N_VPWR_c_443_n 0.00477138f $X=3.035 $Y=1.77 $X2=0
+ $Y2=0
cc_237 N_A_321_369#_c_288_n N_VPWR_c_445_n 0.0100189f $X=3.035 $Y=1.77 $X2=0
+ $Y2=0
cc_238 N_A_321_369#_M1001_d N_VPWR_c_435_n 0.00522079f $X=1.605 $Y=1.845 $X2=0
+ $Y2=0
cc_239 N_A_321_369#_c_288_n N_VPWR_c_435_n 0.00788748f $X=3.035 $Y=1.77 $X2=0
+ $Y2=0
cc_240 N_A_321_369#_M1004_g N_VGND_c_535_n 0.00585385f $X=3.06 $Y=0.445 $X2=0
+ $Y2=0
cc_241 N_A_321_369#_c_286_n N_VGND_c_535_n 0.0169048f $X=2.395 $Y=0.48 $X2=0
+ $Y2=0
cc_242 N_A_321_369#_M1000_d N_VGND_c_538_n 0.00264183f $X=2.095 $Y=0.235 $X2=0
+ $Y2=0
cc_243 N_A_321_369#_M1004_g N_VGND_c_538_n 0.0123858f $X=3.06 $Y=0.445 $X2=0
+ $Y2=0
cc_244 N_A_321_369#_c_286_n N_VGND_c_538_n 0.0173842f $X=2.395 $Y=0.48 $X2=0
+ $Y2=0
cc_245 N_A_321_369#_M1004_g N_A_627_47#_c_590_n 0.00184177f $X=3.06 $Y=0.445
+ $X2=0 $Y2=0
cc_246 N_A_321_369#_M1004_g N_A_627_47#_c_592_n 0.00174076f $X=3.06 $Y=0.445
+ $X2=0 $Y2=0
cc_247 N_B2_M1010_g N_B1_M1002_g 0.0209374f $X=3.55 $Y=0.445 $X2=0 $Y2=0
cc_248 N_B2_c_357_n N_B1_c_408_n 0.00655745f $X=3.525 $Y=1.67 $X2=0 $Y2=0
cc_249 N_B2_c_361_n N_B1_c_408_n 0.00503188f $X=3.825 $Y=1.915 $X2=0 $Y2=0
cc_250 N_B2_c_358_n N_B1_c_409_n 0.0334012f $X=3.525 $Y=1.77 $X2=0 $Y2=0
cc_251 B2 N_B1_c_409_n 0.0143455f $X=3.805 $Y=2.125 $X2=0 $Y2=0
cc_252 N_B2_c_361_n N_B1_c_409_n 0.00188914f $X=3.825 $Y=1.915 $X2=0 $Y2=0
cc_253 N_B2_c_355_n B1 0.0209246f $X=3.655 $Y=1.2 $X2=0 $Y2=0
cc_254 N_B2_c_356_n B1 2.2964e-19 $X=3.5 $Y=1.16 $X2=0 $Y2=0
cc_255 N_B2_c_361_n B1 0.0240847f $X=3.825 $Y=1.915 $X2=0 $Y2=0
cc_256 N_B2_c_355_n N_B1_c_407_n 0.00192779f $X=3.655 $Y=1.2 $X2=0 $Y2=0
cc_257 N_B2_c_356_n N_B1_c_407_n 0.0165938f $X=3.5 $Y=1.16 $X2=0 $Y2=0
cc_258 N_B2_c_361_n N_VPWR_c_440_n 0.00294081f $X=3.825 $Y=1.915 $X2=0 $Y2=0
cc_259 N_B2_c_358_n N_VPWR_c_443_n 0.00702461f $X=3.525 $Y=1.77 $X2=0 $Y2=0
cc_260 B2 N_VPWR_c_443_n 0.0167213f $X=3.805 $Y=2.125 $X2=0 $Y2=0
cc_261 N_B2_c_358_n N_VPWR_c_435_n 0.0129134f $X=3.525 $Y=1.77 $X2=0 $Y2=0
cc_262 B2 N_VPWR_c_435_n 0.0125469f $X=3.805 $Y=2.125 $X2=0 $Y2=0
cc_263 B2 A_723_369# 0.00889271f $X=3.805 $Y=2.125 $X2=-0.19 $Y2=-0.24
cc_264 N_B2_c_361_n A_723_369# 0.00117124f $X=3.825 $Y=1.915 $X2=-0.19 $Y2=-0.24
cc_265 N_B2_M1010_g N_VGND_c_534_n 0.00276849f $X=3.55 $Y=0.445 $X2=0 $Y2=0
cc_266 N_B2_M1010_g N_VGND_c_535_n 0.00437852f $X=3.55 $Y=0.445 $X2=0 $Y2=0
cc_267 N_B2_M1010_g N_VGND_c_538_n 0.0062849f $X=3.55 $Y=0.445 $X2=0 $Y2=0
cc_268 N_B2_M1010_g N_A_627_47#_c_590_n 9.54201e-19 $X=3.55 $Y=0.445 $X2=0 $Y2=0
cc_269 N_B2_M1010_g N_A_627_47#_c_591_n 0.0127176f $X=3.55 $Y=0.445 $X2=0 $Y2=0
cc_270 N_B2_c_355_n N_A_627_47#_c_591_n 0.0299003f $X=3.655 $Y=1.2 $X2=0 $Y2=0
cc_271 N_B2_c_356_n N_A_627_47#_c_591_n 0.00263703f $X=3.5 $Y=1.16 $X2=0 $Y2=0
cc_272 N_B2_c_355_n N_A_627_47#_c_592_n 0.0181468f $X=3.655 $Y=1.2 $X2=0 $Y2=0
cc_273 N_B2_c_356_n N_A_627_47#_c_592_n 0.00182889f $X=3.5 $Y=1.16 $X2=0 $Y2=0
cc_274 N_B2_M1010_g N_A_627_47#_c_593_n 5.72217e-19 $X=3.55 $Y=0.445 $X2=0 $Y2=0
cc_275 N_B1_c_409_n N_VPWR_c_440_n 0.00562173f $X=4.05 $Y=1.77 $X2=0 $Y2=0
cc_276 B1 N_VPWR_c_440_n 0.0275562f $X=4.165 $Y=1.105 $X2=0 $Y2=0
cc_277 N_B1_c_407_n N_VPWR_c_440_n 8.3577e-19 $X=4.215 $Y=1.16 $X2=0 $Y2=0
cc_278 N_B1_c_409_n N_VPWR_c_443_n 0.00652714f $X=4.05 $Y=1.77 $X2=0 $Y2=0
cc_279 N_B1_c_409_n N_VPWR_c_435_n 0.0123603f $X=4.05 $Y=1.77 $X2=0 $Y2=0
cc_280 N_B1_M1002_g N_VGND_c_534_n 0.0046109f $X=4.025 $Y=0.445 $X2=0 $Y2=0
cc_281 N_B1_M1002_g N_VGND_c_537_n 0.00401347f $X=4.025 $Y=0.445 $X2=0 $Y2=0
cc_282 N_B1_M1002_g N_VGND_c_538_n 0.00681804f $X=4.025 $Y=0.445 $X2=0 $Y2=0
cc_283 N_B1_M1002_g N_A_627_47#_c_591_n 0.0137702f $X=4.025 $Y=0.445 $X2=0 $Y2=0
cc_284 B1 N_A_627_47#_c_591_n 0.0347024f $X=4.165 $Y=1.105 $X2=0 $Y2=0
cc_285 N_B1_c_407_n N_A_627_47#_c_591_n 0.00722528f $X=4.215 $Y=1.16 $X2=0 $Y2=0
cc_286 N_B1_M1002_g N_A_627_47#_c_593_n 0.00998891f $X=4.025 $Y=0.445 $X2=0
+ $Y2=0
cc_287 N_VPWR_c_435_n N_X_M1007_s 0.00439555f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_288 N_VPWR_c_437_n N_X_c_497_n 0.0791229f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_289 N_VPWR_c_438_n N_X_c_514_n 0.0179342f $X=1.225 $Y=2.32 $X2=0 $Y2=0
cc_290 N_VPWR_c_441_n N_X_c_514_n 0.0191238f $X=1.01 $Y=2.72 $X2=0 $Y2=0
cc_291 N_VPWR_c_435_n N_X_c_514_n 0.0112569f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_292 N_VPWR_c_435_n A_723_369# 0.00422001f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_293 N_VPWR_c_437_n N_VGND_c_531_n 0.0111763f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_294 N_X_c_499_n N_VGND_c_531_n 0.0258205f $X=0.755 $Y=0.37 $X2=0 $Y2=0
cc_295 N_X_c_499_n N_VGND_c_532_n 0.0226664f $X=0.755 $Y=0.37 $X2=0 $Y2=0
cc_296 N_X_c_499_n N_VGND_c_533_n 0.030869f $X=0.755 $Y=0.37 $X2=0 $Y2=0
cc_297 N_X_M1003_d N_VGND_c_538_n 0.0025535f $X=0.57 $Y=0.235 $X2=0 $Y2=0
cc_298 N_X_c_499_n N_VGND_c_538_n 0.0142885f $X=0.755 $Y=0.37 $X2=0 $Y2=0
cc_299 N_VGND_c_538_n A_313_47# 0.00354201f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
cc_300 N_VGND_c_538_n N_A_627_47#_M1004_d 0.00542902f $X=4.37 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_301 N_VGND_c_538_n N_A_627_47#_M1002_d 0.00218422f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_302 N_VGND_c_535_n N_A_627_47#_c_590_n 0.0107942f $X=3.675 $Y=0 $X2=0 $Y2=0
cc_303 N_VGND_c_538_n N_A_627_47#_c_590_n 0.00844976f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_304 N_VGND_c_534_n N_A_627_47#_c_591_n 0.0131415f $X=3.76 $Y=0.39 $X2=0 $Y2=0
cc_305 N_VGND_c_535_n N_A_627_47#_c_591_n 0.00337805f $X=3.675 $Y=0 $X2=0 $Y2=0
cc_306 N_VGND_c_537_n N_A_627_47#_c_591_n 0.00246723f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_307 N_VGND_c_538_n N_A_627_47#_c_591_n 0.0103778f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_308 N_VGND_c_534_n N_A_627_47#_c_593_n 0.0175799f $X=3.76 $Y=0.39 $X2=0 $Y2=0
cc_309 N_VGND_c_537_n N_A_627_47#_c_593_n 0.0175487f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_310 N_VGND_c_538_n N_A_627_47#_c_593_n 0.0139114f $X=4.37 $Y=0 $X2=0 $Y2=0
