* NGSPICE file created from sky130_fd_sc_hdll__nor3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__nor3_1 A B C VGND VNB VPB VPWR Y
M1000 a_211_297# B a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u
M1001 Y B VGND VNB nshort w=650000u l=150000u
+  ad=3.77e+11p pd=3.76e+06u as=6.305e+11p ps=4.54e+06u
M1002 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_117_297# C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1004 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A a_211_297# VPB phighvt w=1e+06u l=180000u
+  ad=6.1e+11p pd=3.22e+06u as=0p ps=0u
.ends

