* File: sky130_fd_sc_hdll__conb_1.pxi.spice
* Created: Thu Aug 27 19:03:43 2020
* 
x_PM_SKY130_FD_SC_HDLL__CONB_1%HI HI N_HI_R1_pos N_HI_c_21_n N_HI_c_22_n
+ PM_SKY130_FD_SC_HDLL__CONB_1%HI
x_PM_SKY130_FD_SC_HDLL__CONB_1%VPWR N_VPWR_c_39_n N_VPWR_c_37_n N_VPWR_c_41_n
+ N_VPWR_c_42_n VPWR N_VPWR_R1_neg N_VPWR_c_43_n N_VPWR_c_38_n
+ PM_SKY130_FD_SC_HDLL__CONB_1%VPWR
x_PM_SKY130_FD_SC_HDLL__CONB_1%VGND N_VGND_c_55_n N_VGND_c_56_n N_VGND_c_57_n
+ VGND N_VGND_R0_pos N_VGND_c_58_n N_VGND_c_59_n
+ PM_SKY130_FD_SC_HDLL__CONB_1%VGND
x_PM_SKY130_FD_SC_HDLL__CONB_1%LO LO N_LO_R0_neg N_LO_c_71_n
+ PM_SKY130_FD_SC_HDLL__CONB_1%LO
cc_1 VNB N_HI_c_21_n 0.112124f $X=-0.19 $Y=-0.24 $X2=0.44 $Y2=0.34
cc_2 VNB N_HI_c_22_n 0.0491283f $X=-0.19 $Y=-0.24 $X2=0.44 $Y2=0.34
cc_3 VNB N_VPWR_c_37_n 0.00887735f $X=-0.19 $Y=-0.24 $X2=0.345 $Y2=0.34
cc_4 VNB N_VPWR_c_38_n 0.0609879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_VGND_c_55_n 0.0141225f $X=-0.19 $Y=-0.24 $X2=0.335 $Y2=1.125
cc_6 VNB N_VGND_c_56_n 0.00557157f $X=-0.19 $Y=-0.24 $X2=0.345 $Y2=1.16
cc_7 VNB N_VGND_c_57_n 0.127423f $X=-0.19 $Y=-0.24 $X2=0.345 $Y2=0.34
cc_8 VNB N_VGND_c_58_n 0.0207924f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_VGND_c_59_n 0.110844f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB LO 0.0188723f $X=-0.19 $Y=-0.24 $X2=0.335 $Y2=1.125
cc_11 VNB N_LO_c_71_n 0.00887735f $X=-0.19 $Y=-0.24 $X2=0.44 $Y2=0.34
cc_12 VPB N_HI_c_22_n 0.0207802f $X=-0.19 $Y=1.305 $X2=0.44 $Y2=0.34
cc_13 VPB N_VPWR_c_39_n 0.00596761f $X=-0.19 $Y=1.305 $X2=0.345 $Y2=1.16
cc_14 VPB N_VPWR_c_37_n 0.152023f $X=-0.19 $Y=1.305 $X2=0.345 $Y2=0.34
cc_15 VPB N_VPWR_c_41_n 0.00984754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_16 VPB N_VPWR_c_42_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0.345 $Y2=0.34
cc_17 VPB N_VPWR_c_43_n 0.0207924f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_18 VPB N_VPWR_c_38_n 0.0498604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_19 VPB LO 0.0539991f $X=-0.19 $Y=1.305 $X2=0.335 $Y2=1.125
cc_20 VPB N_LO_c_71_n 0.135079f $X=-0.19 $Y=1.305 $X2=0.44 $Y2=0.34
cc_21 N_HI_c_22_n N_VPWR_c_39_n 0.0279374f $X=0.44 $Y=0.34 $X2=0 $Y2=0
cc_22 N_HI_c_22_n N_VPWR_c_37_n 0.0460163f $X=0.44 $Y=0.34 $X2=0 $Y2=0
cc_23 N_HI_c_21_n N_VGND_c_56_n 0.00412998f $X=0.44 $Y=0.34 $X2=0 $Y2=0
cc_24 N_HI_c_22_n N_VGND_c_56_n 0.0423296f $X=0.44 $Y=0.34 $X2=0 $Y2=0
cc_25 N_HI_c_21_n N_VGND_c_57_n 0.0689999f $X=0.44 $Y=0.34 $X2=0 $Y2=0
cc_26 N_HI_c_22_n N_VGND_c_57_n 0.00677716f $X=0.44 $Y=0.34 $X2=0 $Y2=0
cc_27 N_HI_c_21_n N_VGND_c_58_n 0.0114454f $X=0.44 $Y=0.34 $X2=0 $Y2=0
cc_28 N_HI_c_22_n N_VGND_c_58_n 0.0354508f $X=0.44 $Y=0.34 $X2=0 $Y2=0
cc_29 N_HI_c_21_n N_VGND_c_59_n 0.013733f $X=0.44 $Y=0.34 $X2=0 $Y2=0
cc_30 N_HI_c_22_n N_VGND_c_59_n 0.017754f $X=0.44 $Y=0.34 $X2=0 $Y2=0
cc_31 N_HI_c_21_n LO 8.32646e-19 $X=0.44 $Y=0.34 $X2=-0.19 $Y2=-0.24
cc_32 N_HI_c_22_n LO 0.0735573f $X=0.44 $Y=0.34 $X2=-0.19 $Y2=-0.24
cc_33 N_HI_c_22_n N_LO_c_71_n 0.00181903f $X=0.44 $Y=0.34 $X2=0 $Y2=0
cc_34 N_VPWR_c_39_n LO 0.0478402f $X=0.44 $Y=1.995 $X2=-0.19 $Y2=-0.24
cc_35 N_VPWR_c_37_n LO 0.00798463f $X=0.44 $Y=1.995 $X2=-0.19 $Y2=-0.24
cc_36 N_VPWR_c_43_n LO 0.0354508f $X=1.15 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_37 N_VPWR_c_38_n LO 0.017754f $X=1.15 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_38 N_VPWR_c_39_n N_LO_c_71_n 0.00431607f $X=0.44 $Y=1.995 $X2=0 $Y2=0
cc_39 N_VPWR_c_37_n N_LO_c_71_n 0.0921235f $X=0.44 $Y=1.995 $X2=0 $Y2=0
cc_40 N_VPWR_c_43_n N_LO_c_71_n 0.0114454f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_41 N_VPWR_c_38_n N_LO_c_71_n 0.013733f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_42 N_VGND_c_56_n LO 0.0287839f $X=0.94 $Y=0.32 $X2=-0.19 $Y2=-0.24
cc_43 N_VGND_c_57_n LO 0.0278978f $X=0.94 $Y=0.32 $X2=-0.19 $Y2=-0.24
