* File: sky130_fd_sc_hdll__and4_2.pxi.spice
* Created: Thu Aug 27 18:58:46 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND4_2%A N_A_c_70_n N_A_c_71_n N_A_M1002_g N_A_M1007_g A
+ A A A N_A_c_69_n PM_SKY130_FD_SC_HDLL__AND4_2%A
x_PM_SKY130_FD_SC_HDLL__AND4_2%B N_B_M1006_g N_B_c_105_n N_B_c_106_n N_B_M1008_g
+ B B N_B_c_104_n PM_SKY130_FD_SC_HDLL__AND4_2%B
x_PM_SKY130_FD_SC_HDLL__AND4_2%C N_C_M1009_g N_C_c_143_n N_C_c_144_n N_C_M1003_g
+ C C C N_C_c_142_n PM_SKY130_FD_SC_HDLL__AND4_2%C
x_PM_SKY130_FD_SC_HDLL__AND4_2%D N_D_M1001_g N_D_c_181_n N_D_c_182_n N_D_M1010_g
+ D D N_D_c_180_n PM_SKY130_FD_SC_HDLL__AND4_2%D
x_PM_SKY130_FD_SC_HDLL__AND4_2%A_27_47# N_A_27_47#_M1007_s N_A_27_47#_M1002_d
+ N_A_27_47#_M1003_d N_A_27_47#_c_220_n N_A_27_47#_M1000_g N_A_27_47#_c_225_n
+ N_A_27_47#_M1004_g N_A_27_47#_c_226_n N_A_27_47#_M1011_g N_A_27_47#_c_221_n
+ N_A_27_47#_M1005_g N_A_27_47#_c_222_n N_A_27_47#_c_228_n N_A_27_47#_c_229_n
+ N_A_27_47#_c_230_n N_A_27_47#_c_231_n N_A_27_47#_c_232_n N_A_27_47#_c_223_n
+ N_A_27_47#_c_245_n N_A_27_47#_c_234_n N_A_27_47#_c_224_n
+ PM_SKY130_FD_SC_HDLL__AND4_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__AND4_2%VPWR N_VPWR_M1002_s N_VPWR_M1008_d N_VPWR_M1010_d
+ N_VPWR_M1011_s N_VPWR_c_323_n N_VPWR_c_324_n N_VPWR_c_325_n N_VPWR_c_326_n
+ N_VPWR_c_327_n N_VPWR_c_328_n N_VPWR_c_329_n N_VPWR_c_330_n VPWR
+ N_VPWR_c_331_n N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_322_n
+ PM_SKY130_FD_SC_HDLL__AND4_2%VPWR
x_PM_SKY130_FD_SC_HDLL__AND4_2%X N_X_M1000_s N_X_M1004_d X X X X X X X
+ N_X_c_378_n X PM_SKY130_FD_SC_HDLL__AND4_2%X
x_PM_SKY130_FD_SC_HDLL__AND4_2%VGND N_VGND_M1001_d N_VGND_M1005_d N_VGND_c_408_n
+ N_VGND_c_409_n N_VGND_c_410_n N_VGND_c_411_n N_VGND_c_412_n VGND
+ N_VGND_c_413_n N_VGND_c_414_n PM_SKY130_FD_SC_HDLL__AND4_2%VGND
cc_1 VNB N_A_M1007_g 0.0329646f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB A 0.0123633f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_3 VNB N_A_c_69_n 0.046476f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_4 VNB N_B_M1006_g 0.0260522f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.99
cc_5 VNB B 0.00831098f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_6 VNB N_B_c_104_n 0.0196241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_C_M1009_g 0.0289552f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.99
cc_8 VNB C 0.00439626f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_9 VNB N_C_c_142_n 0.0206952f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_D_M1001_g 0.0319324f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.99
cc_11 VNB D 0.00496168f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_12 VNB N_D_c_180_n 0.0222558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_220_n 0.0194906f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_14 VNB N_A_27_47#_c_221_n 0.0233081f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_15 VNB N_A_27_47#_c_222_n 0.00405332f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_16 VNB N_A_27_47#_c_223_n 3.65887e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_224_n 0.0593945f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_322_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB X 0.00213477f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_408_n 0.00469317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_409_n 0.0118978f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_22 VNB N_VGND_c_410_n 0.0293542f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.785
cc_23 VNB N_VGND_c_411_n 0.0642926f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_412_n 0.00324283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_413_n 0.0211781f $X=-0.19 $Y=-0.24 $X2=0.227 $Y2=1.16
cc_26 VNB N_VGND_c_414_n 0.201178f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VPB N_A_c_70_n 0.0328413f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_28 VPB N_A_c_71_n 0.0252831f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_29 VPB A 0.035367f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_30 VPB N_A_c_69_n 0.0123377f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_31 VPB N_B_c_105_n 0.0315211f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_32 VPB N_B_c_106_n 0.022247f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_33 VPB B 0.00192179f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_34 VPB N_B_c_104_n 0.00304612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_C_c_143_n 0.0317747f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_36 VPB N_C_c_144_n 0.0229263f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_37 VPB C 0.00151812f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_38 VPB N_C_c_142_n 0.00311522f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_D_c_181_n 0.0352253f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_40 VPB N_D_c_182_n 0.025213f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_41 VPB D 0.00127851f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_42 VPB N_D_c_180_n 0.0032159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_47#_c_225_n 0.017701f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.785
cc_44 VPB N_A_27_47#_c_226_n 0.0212262f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_47#_c_222_n 0.00199676f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_46 VPB N_A_27_47#_c_228_n 0.00790718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_27_47#_c_229_n 0.0122537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_27_47#_c_230_n 0.0074586f $X=-0.19 $Y=1.305 $X2=0.227 $Y2=1.53
cc_49 VPB N_A_27_47#_c_231_n 0.00858669f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_47#_c_232_n 0.00400408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_c_223_n 0.00196678f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_47#_c_234_n 0.00580186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_c_224_n 0.0282259f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_323_n 0.0103622f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.785
cc_55 VPB N_VPWR_c_324_n 0.0128547f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_325_n 0.00623254f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_57 VPB N_VPWR_c_326_n 0.00519418f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_58 VPB N_VPWR_c_327_n 0.0119952f $X=-0.19 $Y=1.305 $X2=0.227 $Y2=0.85
cc_59 VPB N_VPWR_c_328_n 0.03142f $X=-0.19 $Y=1.305 $X2=0.227 $Y2=1.16
cc_60 VPB N_VPWR_c_329_n 0.0230609f $X=-0.19 $Y=1.305 $X2=0.227 $Y2=1.87
cc_61 VPB N_VPWR_c_330_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_331_n 0.0156737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_332_n 0.0218683f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_333_n 0.00513801f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_322_n 0.0438995f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB X 9.52925e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 N_A_M1007_g N_B_M1006_g 0.0213875f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_68 N_A_c_70_n N_B_c_105_n 0.0213875f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_69 N_A_c_71_n N_B_c_106_n 0.031614f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_70 N_A_M1007_g B 0.00209584f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_71 N_A_c_69_n N_B_c_104_n 0.0213875f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_c_70_n N_A_27_47#_c_222_n 0.00402997f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_73 N_A_M1007_g N_A_27_47#_c_222_n 0.0141693f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_74 A N_A_27_47#_c_222_n 0.0523938f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_75 N_A_c_69_n N_A_27_47#_c_222_n 0.00912063f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_c_70_n N_A_27_47#_c_228_n 0.00300536f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_77 N_A_c_71_n N_A_27_47#_c_228_n 0.00516374f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_78 A N_A_27_47#_c_228_n 0.0203383f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_79 N_A_c_70_n N_A_27_47#_c_230_n 0.00915498f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_80 A N_A_27_47#_c_230_n 0.0136075f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_81 N_A_M1007_g N_A_27_47#_c_245_n 0.0104905f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_82 A N_A_27_47#_c_245_n 0.0129122f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_83 N_A_c_69_n N_A_27_47#_c_245_n 0.00356085f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_84 A N_VPWR_M1002_s 0.0023304f $X=0.15 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_85 N_A_c_71_n N_VPWR_c_324_n 0.00857735f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_86 A N_VPWR_c_324_n 0.0163288f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_87 N_A_c_71_n N_VPWR_c_325_n 5.87379e-19 $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_88 N_A_c_71_n N_VPWR_c_331_n 0.00643335f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_89 N_A_c_71_n N_VPWR_c_322_n 0.0106848f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_90 A N_VPWR_c_322_n 0.00103325f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_91 N_A_M1007_g N_VGND_c_411_n 0.00357877f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_92 A N_VGND_c_411_n 7.89669e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_93 N_A_M1007_g N_VGND_c_414_n 0.00625228f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_94 A N_VGND_c_414_n 0.00167133f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_95 N_B_M1006_g N_C_M1009_g 0.0302261f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_96 B N_C_M1009_g 0.00627179f $X=1.06 $Y=0.425 $X2=0 $Y2=0
cc_97 N_B_c_105_n N_C_c_143_n 0.0146709f $X=0.965 $Y=1.89 $X2=0 $Y2=0
cc_98 N_B_c_106_n N_C_c_144_n 0.0256038f $X=0.965 $Y=1.99 $X2=0 $Y2=0
cc_99 N_B_M1006_g C 5.20291e-19 $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_100 B C 0.0715341f $X=1.06 $Y=0.425 $X2=0 $Y2=0
cc_101 N_B_c_104_n C 3.16267e-19 $X=1 $Y=1.16 $X2=0 $Y2=0
cc_102 N_B_c_104_n N_C_c_142_n 0.0190095f $X=1 $Y=1.16 $X2=0 $Y2=0
cc_103 N_B_M1006_g N_A_27_47#_c_222_n 0.00229932f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_104 N_B_c_105_n N_A_27_47#_c_222_n 0.00342502f $X=0.965 $Y=1.89 $X2=0 $Y2=0
cc_105 B N_A_27_47#_c_222_n 0.0529471f $X=1.06 $Y=0.425 $X2=0 $Y2=0
cc_106 N_B_c_105_n N_A_27_47#_c_228_n 0.00663212f $X=0.965 $Y=1.89 $X2=0 $Y2=0
cc_107 N_B_c_106_n N_A_27_47#_c_228_n 0.00216043f $X=0.965 $Y=1.99 $X2=0 $Y2=0
cc_108 N_B_c_105_n N_A_27_47#_c_229_n 0.0178401f $X=0.965 $Y=1.89 $X2=0 $Y2=0
cc_109 B N_A_27_47#_c_229_n 0.0299509f $X=1.06 $Y=0.425 $X2=0 $Y2=0
cc_110 N_B_c_104_n N_A_27_47#_c_229_n 4.93463e-19 $X=1 $Y=1.16 $X2=0 $Y2=0
cc_111 N_B_M1006_g N_A_27_47#_c_245_n 0.00466494f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_112 N_B_c_106_n N_VPWR_c_324_n 5.03052e-19 $X=0.965 $Y=1.99 $X2=0 $Y2=0
cc_113 N_B_c_106_n N_VPWR_c_325_n 0.0139697f $X=0.965 $Y=1.99 $X2=0 $Y2=0
cc_114 N_B_c_106_n N_VPWR_c_331_n 0.00643335f $X=0.965 $Y=1.99 $X2=0 $Y2=0
cc_115 N_B_c_106_n N_VPWR_c_322_n 0.0106848f $X=0.965 $Y=1.99 $X2=0 $Y2=0
cc_116 B A_203_47# 0.00456934f $X=1.06 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_117 N_B_M1006_g N_VGND_c_411_n 0.0038979f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_118 B N_VGND_c_411_n 0.0114757f $X=1.06 $Y=0.425 $X2=0 $Y2=0
cc_119 N_B_M1006_g N_VGND_c_414_n 0.00564572f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_120 B N_VGND_c_414_n 0.012494f $X=1.06 $Y=0.425 $X2=0 $Y2=0
cc_121 N_C_M1009_g N_D_M1001_g 0.0319714f $X=1.43 $Y=0.445 $X2=0 $Y2=0
cc_122 C N_D_M1001_g 0.0101175f $X=1.515 $Y=0.425 $X2=0 $Y2=0
cc_123 N_C_c_143_n N_D_c_181_n 0.0142193f $X=1.455 $Y=1.89 $X2=0 $Y2=0
cc_124 N_C_c_144_n N_D_c_182_n 0.0240091f $X=1.455 $Y=1.99 $X2=0 $Y2=0
cc_125 N_C_M1009_g D 2.24815e-19 $X=1.43 $Y=0.445 $X2=0 $Y2=0
cc_126 C D 0.0433432f $X=1.515 $Y=0.425 $X2=0 $Y2=0
cc_127 N_C_c_142_n D 3.27643e-19 $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_128 N_C_c_142_n N_D_c_180_n 0.0202006f $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_129 N_C_c_143_n N_A_27_47#_c_229_n 0.0200091f $X=1.455 $Y=1.89 $X2=0 $Y2=0
cc_130 C N_A_27_47#_c_229_n 0.0125111f $X=1.515 $Y=0.425 $X2=0 $Y2=0
cc_131 N_C_c_143_n N_A_27_47#_c_231_n 0.00746798f $X=1.455 $Y=1.89 $X2=0 $Y2=0
cc_132 N_C_c_144_n N_A_27_47#_c_231_n 8.49449e-19 $X=1.455 $Y=1.99 $X2=0 $Y2=0
cc_133 C N_A_27_47#_c_234_n 0.0123056f $X=1.515 $Y=0.425 $X2=0 $Y2=0
cc_134 N_C_c_142_n N_A_27_47#_c_234_n 4.35311e-19 $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_135 N_C_c_144_n N_VPWR_c_325_n 0.00648748f $X=1.455 $Y=1.99 $X2=0 $Y2=0
cc_136 N_C_c_144_n N_VPWR_c_329_n 0.00721387f $X=1.455 $Y=1.99 $X2=0 $Y2=0
cc_137 N_C_c_144_n N_VPWR_c_322_n 0.0127316f $X=1.455 $Y=1.99 $X2=0 $Y2=0
cc_138 C A_301_47# 0.00531584f $X=1.515 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_139 C N_VGND_c_408_n 0.00407967f $X=1.515 $Y=0.425 $X2=0 $Y2=0
cc_140 N_C_M1009_g N_VGND_c_411_n 0.00455696f $X=1.43 $Y=0.445 $X2=0 $Y2=0
cc_141 C N_VGND_c_411_n 0.00914931f $X=1.515 $Y=0.425 $X2=0 $Y2=0
cc_142 N_C_M1009_g N_VGND_c_414_n 0.00761943f $X=1.43 $Y=0.445 $X2=0 $Y2=0
cc_143 C N_VGND_c_414_n 0.00998001f $X=1.515 $Y=0.425 $X2=0 $Y2=0
cc_144 N_D_M1001_g N_A_27_47#_c_220_n 0.0139869f $X=1.91 $Y=0.445 $X2=0 $Y2=0
cc_145 D N_A_27_47#_c_220_n 0.00434768f $X=1.975 $Y=0.765 $X2=0 $Y2=0
cc_146 N_D_c_181_n N_A_27_47#_c_225_n 0.0109135f $X=1.935 $Y=1.89 $X2=0 $Y2=0
cc_147 N_D_c_182_n N_A_27_47#_c_225_n 0.0072832f $X=1.935 $Y=1.99 $X2=0 $Y2=0
cc_148 N_D_c_181_n N_A_27_47#_c_231_n 0.00633492f $X=1.935 $Y=1.89 $X2=0 $Y2=0
cc_149 N_D_c_182_n N_A_27_47#_c_231_n 0.00101311f $X=1.935 $Y=1.99 $X2=0 $Y2=0
cc_150 N_D_c_181_n N_A_27_47#_c_232_n 0.0210857f $X=1.935 $Y=1.89 $X2=0 $Y2=0
cc_151 D N_A_27_47#_c_232_n 0.0207642f $X=1.975 $Y=0.765 $X2=0 $Y2=0
cc_152 N_D_c_180_n N_A_27_47#_c_232_n 4.93463e-19 $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_153 N_D_c_181_n N_A_27_47#_c_223_n 0.00259923f $X=1.935 $Y=1.89 $X2=0 $Y2=0
cc_154 D N_A_27_47#_c_223_n 0.0146578f $X=1.975 $Y=0.765 $X2=0 $Y2=0
cc_155 N_D_c_180_n N_A_27_47#_c_223_n 3.69664e-19 $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_156 N_D_c_181_n N_A_27_47#_c_224_n 0.00179597f $X=1.935 $Y=1.89 $X2=0 $Y2=0
cc_157 D N_A_27_47#_c_224_n 0.00269093f $X=1.975 $Y=0.765 $X2=0 $Y2=0
cc_158 N_D_c_180_n N_A_27_47#_c_224_n 0.0118831f $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_159 N_D_c_181_n N_VPWR_c_326_n 0.00170115f $X=1.935 $Y=1.89 $X2=0 $Y2=0
cc_160 N_D_c_182_n N_VPWR_c_326_n 0.00816734f $X=1.935 $Y=1.99 $X2=0 $Y2=0
cc_161 N_D_c_182_n N_VPWR_c_329_n 0.00743866f $X=1.935 $Y=1.99 $X2=0 $Y2=0
cc_162 N_D_c_182_n N_VPWR_c_322_n 0.0137061f $X=1.935 $Y=1.99 $X2=0 $Y2=0
cc_163 N_D_M1001_g N_X_c_378_n 9.20006e-19 $X=1.91 $Y=0.445 $X2=0 $Y2=0
cc_164 D N_X_c_378_n 0.00231203f $X=1.975 $Y=0.765 $X2=0 $Y2=0
cc_165 D N_VGND_M1001_d 0.00396695f $X=1.975 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_166 N_D_M1001_g N_VGND_c_408_n 0.00661286f $X=1.91 $Y=0.445 $X2=0 $Y2=0
cc_167 N_D_M1001_g N_VGND_c_411_n 0.00489262f $X=1.91 $Y=0.445 $X2=0 $Y2=0
cc_168 D N_VGND_c_411_n 0.00407684f $X=1.975 $Y=0.765 $X2=0 $Y2=0
cc_169 N_D_M1001_g N_VGND_c_414_n 0.00844242f $X=1.91 $Y=0.445 $X2=0 $Y2=0
cc_170 D N_VGND_c_414_n 0.00689956f $X=1.975 $Y=0.765 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_232_n N_VPWR_M1010_d 0.0191981f $X=2.495 $Y=1.58 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_228_n N_VPWR_c_324_n 0.0127138f $X=0.73 $Y=2.3 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_228_n N_VPWR_c_325_n 0.0334757f $X=0.73 $Y=2.3 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_229_n N_VPWR_c_325_n 0.0208202f $X=1.57 $Y=1.58 $X2=0 $Y2=0
cc_175 N_A_27_47#_c_231_n N_VPWR_c_325_n 0.0220026f $X=1.695 $Y=2.3 $X2=0 $Y2=0
cc_176 N_A_27_47#_c_225_n N_VPWR_c_326_n 0.00528945f $X=2.605 $Y=1.41 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_231_n N_VPWR_c_326_n 0.0199759f $X=1.695 $Y=2.3 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_232_n N_VPWR_c_326_n 0.0201769f $X=2.495 $Y=1.58 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_226_n N_VPWR_c_328_n 0.00486741f $X=3.135 $Y=1.41 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_231_n N_VPWR_c_329_n 0.0152795f $X=1.695 $Y=2.3 $X2=0 $Y2=0
cc_181 N_A_27_47#_c_228_n N_VPWR_c_331_n 0.0118139f $X=0.73 $Y=2.3 $X2=0 $Y2=0
cc_182 N_A_27_47#_c_225_n N_VPWR_c_332_n 0.00597712f $X=2.605 $Y=1.41 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_226_n N_VPWR_c_332_n 0.00658436f $X=3.135 $Y=1.41 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_M1002_d N_VPWR_c_322_n 0.0060606f $X=0.585 $Y=2.065 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_M1003_d N_VPWR_c_322_n 0.0037108f $X=1.545 $Y=2.065 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_225_n N_VPWR_c_322_n 0.0106636f $X=2.605 $Y=1.41 $X2=0 $Y2=0
cc_187 N_A_27_47#_c_226_n N_VPWR_c_322_n 0.0125201f $X=3.135 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_228_n N_VPWR_c_322_n 0.00646998f $X=0.73 $Y=2.3 $X2=0 $Y2=0
cc_189 N_A_27_47#_c_231_n N_VPWR_c_322_n 0.00955092f $X=1.695 $Y=2.3 $X2=0 $Y2=0
cc_190 N_A_27_47#_c_220_n X 0.00311861f $X=2.58 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_27_47#_c_225_n X 0.00464862f $X=2.605 $Y=1.41 $X2=0 $Y2=0
cc_192 N_A_27_47#_c_226_n X 0.0228658f $X=3.135 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_221_n X 0.00708519f $X=3.16 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_27_47#_c_232_n X 0.0136906f $X=2.495 $Y=1.58 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_223_n X 0.0353969f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A_27_47#_c_224_n X 0.0393087f $X=3.135 $Y=1.202 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_220_n N_X_c_378_n 0.00896527f $X=2.58 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_223_n N_X_c_378_n 0.00250298f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A_27_47#_c_224_n N_X_c_378_n 0.00375314f $X=3.135 $Y=1.202 $X2=0 $Y2=0
cc_200 N_A_27_47#_c_225_n X 0.0122029f $X=2.605 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_226_n X 0.0167053f $X=3.135 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A_27_47#_c_232_n X 0.00323636f $X=2.495 $Y=1.58 $X2=0 $Y2=0
cc_203 N_A_27_47#_c_224_n X 0.00331798f $X=3.135 $Y=1.202 $X2=0 $Y2=0
cc_204 N_A_27_47#_c_222_n A_119_47# 6.59066e-19 $X=0.585 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_205 N_A_27_47#_c_245_n A_119_47# 0.00389845f $X=0.585 $Y=0.42 $X2=-0.19
+ $Y2=-0.24
cc_206 N_A_27_47#_c_220_n N_VGND_c_408_n 0.0030265f $X=2.58 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A_27_47#_c_221_n N_VGND_c_410_n 0.00491123f $X=3.16 $Y=0.995 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_c_245_n N_VGND_c_411_n 0.0289623f $X=0.585 $Y=0.42 $X2=0 $Y2=0
cc_209 N_A_27_47#_c_220_n N_VGND_c_413_n 0.00542953f $X=2.58 $Y=0.995 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_221_n N_VGND_c_413_n 0.00585385f $X=3.16 $Y=0.995 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_M1007_s N_VGND_c_414_n 0.00271953f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_220_n N_VGND_c_414_n 0.0103952f $X=2.58 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A_27_47#_c_221_n N_VGND_c_414_n 0.0118925f $X=3.16 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A_27_47#_c_245_n N_VGND_c_414_n 0.0179555f $X=0.585 $Y=0.42 $X2=0 $Y2=0
cc_215 N_VPWR_c_322_n N_X_M1004_d 0.00280243f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_216 N_VPWR_c_326_n X 0.0416608f $X=2.33 $Y=2 $X2=0 $Y2=0
cc_217 N_VPWR_c_332_n X 0.0272312f $X=3.245 $Y=2.72 $X2=0 $Y2=0
cc_218 N_VPWR_c_322_n X 0.0167167f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_219 N_X_c_378_n N_VGND_c_413_n 0.0219969f $X=2.84 $Y=0.38 $X2=0 $Y2=0
cc_220 N_X_M1000_s N_VGND_c_414_n 0.00387469f $X=2.655 $Y=0.235 $X2=0 $Y2=0
cc_221 N_X_c_378_n N_VGND_c_414_n 0.0166401f $X=2.84 $Y=0.38 $X2=0 $Y2=0
cc_222 A_119_47# N_VGND_c_414_n 0.0086256f $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_223 A_203_47# N_VGND_c_414_n 0.00713426f $X=1.015 $Y=0.235 $X2=0 $Y2=0
cc_224 A_301_47# N_VGND_c_414_n 0.00737302f $X=1.505 $Y=0.235 $X2=0 $Y2=0
