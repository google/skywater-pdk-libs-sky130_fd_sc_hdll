* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
X0 a_27_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X1 VGND D a_841_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_641_47# C a_841_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y a_211_413# a_361_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 a_641_47# a_27_47# a_361_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 VGND A_N a_211_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 a_841_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Y a_211_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 a_361_47# a_211_413# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR A_N a_211_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X13 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 a_27_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_361_47# a_27_47# a_641_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_841_47# C a_641_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VPWR a_211_413# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
