* File: sky130_fd_sc_hdll__o21ai_2.spice
* Created: Thu Aug 27 19:19:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o21ai_2.pex.spice"
.subckt sky130_fd_sc_hdll__o21ai_2  VNB VPB A1 A2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1000 N_A_29_47#_M1000_d N_A1_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.20475 AS=0.10725 PD=1.93 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1009 N_A_29_47#_M1009_d N_A2_M1009_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75000.7
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1010 N_A_29_47#_M1009_d N_A2_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.143 PD=0.98 PS=1.09 NRD=9.228 NRS=9.228 M=1 R=4.33333
+ SA=75001.2 SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1008 N_A_29_47#_M1008_d N_A1_M1008_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.143 PD=0.93 PS=1.09 NRD=0 NRS=20.304 M=1 R=4.33333 SA=75001.8
+ SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_B1_M1004_g N_A_29_47#_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.091 PD=0.98 PS=0.93 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75002.2
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1004_d N_B1_M1006_g N_A_29_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.273 PD=0.98 PS=2.14 NRD=0 NRS=28.608 M=1 R=4.33333 SA=75002.7
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1002 N_A_120_297#_M1002_d N_A1_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90002.8 A=0.18 P=2.36 MULT=1
MM1003 N_A_120_297#_M1002_d N_A2_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90002.3 A=0.18 P=2.36 MULT=1
MM1007 N_A_120_297#_M1007_d N_A2_M1007_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.185 AS=0.15 PD=1.37 PS=1.3 NRD=11.8003 NRS=1.9503 M=1 R=5.55556
+ SA=90001.1 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1005 N_A_120_297#_M1007_d N_A1_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.185 AS=0.17 PD=1.37 PS=1.34 NRD=5.8903 NRS=4.9053 M=1 R=5.55556
+ SA=90001.7 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.17 PD=1.3 PS=1.34 NRD=1.9503 NRS=6.8753 M=1 R=5.55556 SA=90002.2
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1011 N_Y_M1001_d N_B1_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.38 PD=1.3 PS=2.76 NRD=1.9503 NRS=22.6353 M=1 R=5.55556 SA=90002.7
+ SB=90000.3 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
pX13_noxref noxref_11 A2 A2 PROBETYPE=1
c_56 VPB 0 8.49032e-20 $X=0.14 $Y=2.635
*
.include "sky130_fd_sc_hdll__o21ai_2.pxi.spice"
*
.ends
*
*
