* File: sky130_fd_sc_hdll__a2bb2o_4.pex.spice
* Created: Thu Aug 27 18:54:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_4%B1 1 3 4 6 7 9 10 12 13 16 20 23 27
c82 16 0 1.00809e-19 $X=1.75 $Y=1.445
c83 13 0 7.96704e-20 $X=1.665 $Y=1.53
c84 7 0 1.85574e-19 $X=1.905 $Y=1.41
c85 4 0 8.54817e-20 $X=0.52 $Y=0.995
r86 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r87 23 33 7.53086 $w=5.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.355 $Y=1.19
+ $X2=0.355 $Y2=1.53
r88 23 27 0.664488 $w=5.38e-07 $l=3e-08 $layer=LI1_cond $X=0.355 $Y=1.19
+ $X2=0.355 $Y2=1.16
r89 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.16 $X2=1.88 $Y2=1.16
r90 17 20 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.75 $Y=1.16
+ $X2=1.88 $Y2=1.16
r91 15 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.75 $Y=1.245
+ $X2=1.75 $Y2=1.16
r92 15 16 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.75 $Y=1.245 $X2=1.75
+ $Y2=1.445
r93 14 33 7.6426 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=0.625 $Y=1.53
+ $X2=0.355 $Y2=1.53
r94 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.665 $Y=1.53
+ $X2=1.75 $Y2=1.445
r95 13 14 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=1.665 $Y=1.53
+ $X2=0.625 $Y2=1.53
r96 10 21 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.905 $Y2=1.16
r97 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r98 7 21 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.16
r99 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r100 4 26 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.435 $Y2=1.16
r101 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=0.56
r102 1 26 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.435 $Y2=1.16
r103 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_4%B2 1 3 4 6 7 9 10 12 13 20 25
c46 25 0 1.85574e-19 $X=1.155 $Y=1.19
c47 10 0 8.861e-20 $X=1.46 $Y=0.995
c48 1 0 1.56165e-19 $X=0.94 $Y=0.995
r49 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.46 $Y2=1.202
r50 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=1.2 $Y=1.202
+ $X2=1.435 $Y2=1.202
r51 18 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2
+ $Y=1.16 $X2=1.2 $Y2=1.16
r52 16 18 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=1.2 $Y2=1.202
r53 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.202
+ $X2=0.965 $Y2=1.202
r54 13 25 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=1.145 $Y=1.175
+ $X2=1.155 $Y2=1.175
r55 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=1.202
r56 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=0.56
r57 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r58 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r59 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r60 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r61 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=1.202
r62 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995 $X2=0.94
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_4%A_455_21# 1 2 3 10 12 13 15 16 18 19 21
+ 22 28 30 31 32 33 37 39 43 45 47 48 56
c137 56 0 1.84956e-19 $X=2.87 $Y=1.202
c138 16 0 4.99794e-20 $X=2.845 $Y=1.41
c139 13 0 2.38703e-19 $X=2.375 $Y=1.41
r140 55 56 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=2.87 $Y2=1.202
r141 54 55 62.0658 $w=3.65e-07 $l=4.7e-07 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.845 $Y2=1.202
r142 53 54 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.202
+ $X2=2.375 $Y2=1.202
r143 48 51 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=1.875
+ $X2=4.54 $Y2=1.96
r144 41 43 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.985 $Y=0.725
+ $X2=4.985 $Y2=0.39
r145 40 47 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.235 $Y=0.815
+ $X2=4.045 $Y2=0.815
r146 39 41 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=4.795 $Y=0.815
+ $X2=4.985 $Y2=0.725
r147 39 40 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.795 $Y=0.815
+ $X2=4.235 $Y2=0.815
r148 35 47 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=4.045 $Y=0.725
+ $X2=4.045 $Y2=0.815
r149 35 37 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.045 $Y=0.725
+ $X2=4.045 $Y2=0.39
r150 34 46 2.30104 $w=1.8e-07 $l=1.7e-07 $layer=LI1_cond $X=3.605 $Y=1.875
+ $X2=3.435 $Y2=1.875
r151 33 48 2.6621 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.415 $Y=1.875
+ $X2=4.54 $Y2=1.875
r152 33 34 49.9091 $w=1.78e-07 $l=8.1e-07 $layer=LI1_cond $X=4.415 $Y=1.875
+ $X2=3.605 $Y2=1.875
r153 31 47 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.855 $Y=0.815
+ $X2=4.045 $Y2=0.815
r154 31 32 25.2626 $w=1.78e-07 $l=4.1e-07 $layer=LI1_cond $X=3.855 $Y=0.815
+ $X2=3.445 $Y2=0.815
r155 30 46 20.2107 $w=2.35e-07 $l=4.20357e-07 $layer=LI1_cond $X=3.35 $Y=1.495
+ $X2=3.435 $Y2=1.875
r156 29 45 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.35 $Y=1.245
+ $X2=3.35 $Y2=1.16
r157 29 30 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=3.35 $Y=1.245
+ $X2=3.35 $Y2=1.495
r158 28 45 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.35 $Y=1.075
+ $X2=3.35 $Y2=1.16
r159 27 32 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=3.35 $Y=0.905
+ $X2=3.445 $Y2=0.815
r160 27 28 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=3.35 $Y=0.905
+ $X2=3.35 $Y2=1.075
r161 25 56 27.7315 $w=3.65e-07 $l=2.1e-07 $layer=POLY_cond $X=3.08 $Y=1.202
+ $X2=2.87 $Y2=1.202
r162 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.08
+ $Y=1.16 $X2=3.08 $Y2=1.16
r163 22 45 1.74598 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.255 $Y=1.16
+ $X2=3.35 $Y2=1.16
r164 22 24 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.255 $Y=1.16
+ $X2=3.08 $Y2=1.16
r165 19 56 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.87 $Y=0.995
+ $X2=2.87 $Y2=1.202
r166 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.87 $Y=0.995
+ $X2=2.87 $Y2=0.56
r167 16 55 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r168 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r169 13 54 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r170 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r171 10 53 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.202
r172 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=0.56
r173 3 51 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.485 $X2=4.54 $Y2=1.96
r174 2 43 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.875
+ $Y=0.235 $X2=5.01 $Y2=0.39
r175 1 37 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.935
+ $Y=0.235 $X2=4.07 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_4%A1_N 1 3 4 6 7 9 10 12 13 16 19
c86 19 0 1.6626e-19 $X=5.29 $Y=1.19
c87 16 0 1.84956e-19 $X=3.78 $Y=1.16
c88 10 0 7.88531e-20 $X=5.27 $Y=0.995
c89 7 0 2.90838e-19 $X=5.245 $Y=1.41
r90 19 28 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=5.275 $Y=1.16
+ $X2=5.275 $Y2=1.53
r91 19 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.25
+ $Y=1.16 $X2=5.25 $Y2=1.16
r92 16 18 14.8487 $w=3.04e-07 $l=3.7e-07 $layer=LI1_cond $X=3.81 $Y=1.16
+ $X2=3.81 $Y2=1.53
r93 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.78
+ $Y=1.16 $X2=3.78 $Y2=1.16
r94 14 18 4.13891 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.005 $Y=1.53
+ $X2=3.81 $Y2=1.53
r95 13 28 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.085 $Y=1.53
+ $X2=5.275 $Y2=1.53
r96 13 14 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=5.085 $Y=1.53
+ $X2=4.005 $Y2=1.53
r97 10 23 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=5.27 $Y=0.995
+ $X2=5.245 $Y2=1.16
r98 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.27 $Y=0.995
+ $X2=5.27 $Y2=0.56
r99 7 23 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.16
r100 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.985
r101 4 17 38.7084 $w=3.43e-07 $l=1.90526e-07 $layer=POLY_cond $X=3.86 $Y=0.995
+ $X2=3.805 $Y2=1.16
r102 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.86 $Y=0.995
+ $X2=3.86 $Y2=0.56
r103 1 17 45.964 $w=3.43e-07 $l=2.64575e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.805 $Y2=1.16
r104 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_4%A2_N 1 3 4 6 7 9 10 12 13 19 20
r49 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.775 $Y=1.202
+ $X2=4.8 $Y2=1.202
r50 18 20 8.24474 $w=3.8e-07 $l=6.5e-08 $layer=POLY_cond $X=4.71 $Y=1.202
+ $X2=4.775 $Y2=1.202
r51 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.71
+ $Y=1.16 $X2=4.71 $Y2=1.16
r52 16 18 51.3711 $w=3.8e-07 $l=4.05e-07 $layer=POLY_cond $X=4.305 $Y=1.202
+ $X2=4.71 $Y2=1.202
r53 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.28 $Y=1.202
+ $X2=4.305 $Y2=1.202
r54 13 19 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=4.37 $Y=1.175
+ $X2=4.71 $Y2=1.175
r55 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.8 $Y=0.995
+ $X2=4.8 $Y2=1.202
r56 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.8 $Y=0.995 $X2=4.8
+ $Y2=0.56
r57 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.202
r58 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
r59 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.202
r60 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.985
r61 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.28 $Y=0.995
+ $X2=4.28 $Y2=1.202
r62 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.28 $Y=0.995 $X2=4.28
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_4%A_203_47# 1 2 3 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 31 33 34 38 41 47 51 55 56 57 63 74 78 81
c169 63 0 1.52229e-19 $X=5.815 $Y=1.53
c170 51 0 1.74092e-19 $X=1.2 $Y=0.73
c171 41 0 1.08203e-19 $X=2.59 $Y=1.415
c172 34 0 1.29925e-20 $X=2.395 $Y=0.82
c173 28 0 1.66154e-19 $X=7.125 $Y=1.41
r174 78 80 11.7175 $w=3.54e-07 $l=3.4e-07 $layer=LI1_cond $X=2.677 $Y=1.62
+ $X2=2.677 $Y2=1.96
r175 74 75 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.125 $Y=1.202
+ $X2=7.15 $Y2=1.202
r176 71 72 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.63 $Y=1.202
+ $X2=6.655 $Y2=1.202
r177 70 71 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=6.185 $Y=1.202
+ $X2=6.63 $Y2=1.202
r178 69 70 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.16 $Y=1.202
+ $X2=6.185 $Y2=1.202
r179 66 67 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.69 $Y=1.202
+ $X2=5.715 $Y2=1.202
r180 64 81 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=5.822 $Y=1.53
+ $X2=5.822 $Y2=1.16
r181 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.815 $Y=1.53
+ $X2=5.815 $Y2=1.53
r182 60 78 3.10169 $w=3.54e-07 $l=9e-08 $layer=LI1_cond $X=2.677 $Y=1.53
+ $X2=2.677 $Y2=1.62
r183 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.785 $Y=1.53
+ $X2=2.785 $Y2=1.53
r184 57 59 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=2.98 $Y=1.53
+ $X2=2.785 $Y2=1.53
r185 56 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.67 $Y=1.53
+ $X2=5.815 $Y2=1.53
r186 56 57 3.3292 $w=1.4e-07 $l=2.69e-06 $layer=MET1_cond $X=5.67 $Y=1.53
+ $X2=2.98 $Y2=1.53
r187 51 53 2.69402 $w=3.83e-07 $l=9e-08 $layer=LI1_cond $X=1.177 $Y=0.73
+ $X2=1.177 $Y2=0.82
r188 48 74 34.336 $w=3.72e-07 $l=2.65e-07 $layer=POLY_cond $X=6.86 $Y=1.202
+ $X2=7.125 $Y2=1.202
r189 48 72 26.5618 $w=3.72e-07 $l=2.05e-07 $layer=POLY_cond $X=6.86 $Y=1.202
+ $X2=6.655 $Y2=1.202
r190 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.86
+ $Y=1.16 $X2=6.86 $Y2=1.16
r191 45 69 10.3656 $w=3.72e-07 $l=8e-08 $layer=POLY_cond $X=6.08 $Y=1.202
+ $X2=6.16 $Y2=1.202
r192 45 67 47.293 $w=3.72e-07 $l=3.65e-07 $layer=POLY_cond $X=6.08 $Y=1.202
+ $X2=5.715 $Y2=1.202
r193 44 47 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=6.08 $Y=1.16
+ $X2=6.86 $Y2=1.16
r194 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.08
+ $Y=1.16 $X2=6.08 $Y2=1.16
r195 42 81 5.38787 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=6.01 $Y=1.16
+ $X2=5.822 $Y2=1.16
r196 42 44 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=6.01 $Y=1.16 $X2=6.08
+ $Y2=1.16
r197 41 60 5.96567 $w=3.54e-07 $l=1.52414e-07 $layer=LI1_cond $X=2.59 $Y=1.415
+ $X2=2.677 $Y2=1.53
r198 40 55 3.19717 $w=2.95e-07 $l=8.74643e-08 $layer=LI1_cond $X=2.59 $Y=0.905
+ $X2=2.585 $Y2=0.82
r199 40 41 26.9351 $w=2.08e-07 $l=5.1e-07 $layer=LI1_cond $X=2.59 $Y=0.905
+ $X2=2.59 $Y2=1.415
r200 36 55 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=0.735
+ $X2=2.585 $Y2=0.82
r201 36 38 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=2.585 $Y=0.735
+ $X2=2.585 $Y2=0.39
r202 35 53 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.37 $Y=0.82
+ $X2=1.177 $Y2=0.82
r203 34 55 3.3845 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=0.82
+ $X2=2.585 $Y2=0.82
r204 34 35 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=2.395 $Y=0.82
+ $X2=1.37 $Y2=0.82
r205 31 75 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.15 $Y=0.995
+ $X2=7.15 $Y2=1.202
r206 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.15 $Y=0.995
+ $X2=7.15 $Y2=0.56
r207 28 74 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.202
r208 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.985
r209 25 72 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.202
r210 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.985
r211 22 71 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=1.202
r212 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=0.56
r213 19 70 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.202
r214 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.985
r215 16 69 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=1.202
r216 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=0.56
r217 13 67 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.202
r218 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.985
r219 10 66 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=1.202
r220 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=0.56
r221 3 80 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.96
r222 3 78 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.62
r223 2 38 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.39
r224 1 51 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_4%A_27_297# 1 2 3 4 15 17 18 21 23 31 33 34
+ 35 36 38
r53 38 40 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.08 $Y=2.3 $X2=3.08
+ $Y2=2.38
r54 33 40 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.955 $Y=2.38
+ $X2=3.08 $Y2=2.38
r55 33 34 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.955 $Y=2.38
+ $X2=2.265 $Y2=2.38
r56 29 36 3.98977 $w=2.3e-07 $l=9.44722e-08 $layer=LI1_cond $X=2.16 $Y=1.785
+ $X2=2.14 $Y2=1.87
r57 29 31 8.71429 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=2.16 $Y=1.785
+ $X2=2.16 $Y2=1.62
r58 26 34 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.14 $Y=2.295
+ $X2=2.265 $Y2=2.38
r59 26 28 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.14 $Y=2.295
+ $X2=2.14 $Y2=1.96
r60 25 36 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=1.955
+ $X2=2.14 $Y2=1.87
r61 25 28 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=2.14 $Y=1.955
+ $X2=2.14 $Y2=1.96
r62 24 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.325 $Y=1.87
+ $X2=1.2 $Y2=1.87
r63 23 36 2.45049 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.015 $Y=1.87
+ $X2=2.14 $Y2=1.87
r64 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.015 $Y=1.87
+ $X2=1.325 $Y2=1.87
r65 19 35 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=1.955
+ $X2=1.2 $Y2=1.87
r66 19 21 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.2 $Y=1.955 $X2=1.2
+ $Y2=1.96
r67 17 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.075 $Y=1.87
+ $X2=1.2 $Y2=1.87
r68 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.075 $Y=1.87
+ $X2=0.385 $Y2=1.87
r69 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.26 $Y=1.955
+ $X2=0.385 $Y2=1.87
r70 13 15 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.26 $Y=1.955
+ $X2=0.26 $Y2=1.96
r71 4 38 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2.3
r72 3 31 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.62
r73 3 28 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.96
r74 2 21 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.96
r75 1 15 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_4%VPWR 1 2 3 4 5 6 21 23 27 31 35 39 43 46
+ 47 49 50 52 53 55 56 57 59 84 85 88 91
r118 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r119 89 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r120 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r121 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r122 82 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r123 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r124 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r125 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r126 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r127 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r128 73 76 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r129 72 75 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r130 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r131 70 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r132 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r133 67 70 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r134 67 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r135 66 69 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r136 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r137 64 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.795 $Y=2.72
+ $X2=1.67 $Y2=2.72
r138 64 66 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.795 $Y=2.72
+ $X2=2.07 $Y2=2.72
r139 59 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.605 $Y=2.72
+ $X2=0.73 $Y2=2.72
r140 59 61 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.605 $Y=2.72
+ $X2=0.23 $Y2=2.72
r141 57 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r142 57 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r143 55 81 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.235 $Y=2.72
+ $X2=7.13 $Y2=2.72
r144 55 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.235 $Y=2.72
+ $X2=7.36 $Y2=2.72
r145 54 84 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.485 $Y=2.72
+ $X2=7.59 $Y2=2.72
r146 54 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.485 $Y=2.72
+ $X2=7.36 $Y2=2.72
r147 52 78 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.295 $Y=2.72
+ $X2=6.21 $Y2=2.72
r148 52 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.295 $Y=2.72
+ $X2=6.42 $Y2=2.72
r149 51 81 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=6.545 $Y=2.72
+ $X2=7.13 $Y2=2.72
r150 51 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.545 $Y=2.72
+ $X2=6.42 $Y2=2.72
r151 49 75 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.355 $Y=2.72
+ $X2=5.29 $Y2=2.72
r152 49 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.355 $Y=2.72
+ $X2=5.48 $Y2=2.72
r153 48 78 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=5.605 $Y=2.72
+ $X2=6.21 $Y2=2.72
r154 48 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.605 $Y=2.72
+ $X2=5.48 $Y2=2.72
r155 46 69 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.475 $Y=2.72
+ $X2=3.45 $Y2=2.72
r156 46 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.475 $Y=2.72
+ $X2=3.6 $Y2=2.72
r157 45 72 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.725 $Y=2.72
+ $X2=3.91 $Y2=2.72
r158 45 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.725 $Y=2.72
+ $X2=3.6 $Y2=2.72
r159 41 56 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=2.635
+ $X2=7.36 $Y2=2.72
r160 41 43 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=7.36 $Y=2.635
+ $X2=7.36 $Y2=1.99
r161 37 53 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=2.72
r162 37 39 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=2.33
r163 33 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2.72
r164 33 35 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=1.96
r165 29 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=2.635
+ $X2=3.6 $Y2=2.72
r166 29 31 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.6 $Y=2.635
+ $X2=3.6 $Y2=2.34
r167 25 91 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.72
r168 25 27 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.3
r169 24 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=0.73 $Y2=2.72
r170 23 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.545 $Y=2.72
+ $X2=1.67 $Y2=2.72
r171 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.545 $Y=2.72
+ $X2=0.855 $Y2=2.72
r172 19 88 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.72
r173 19 21 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.3
r174 6 43 300 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_PDIFF $count=2 $X=7.215
+ $Y=1.485 $X2=7.36 $Y2=1.99
r175 5 39 600 $w=1.7e-07 $l=9.14631e-07 $layer=licon1_PDIFF $count=1 $X=6.275
+ $Y=1.485 $X2=6.42 $Y2=2.33
r176 4 35 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=1.96
r177 3 31 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=3.475
+ $Y=1.485 $X2=3.6 $Y2=2.34
r178 2 27 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.3
r179 1 21 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_4%A_785_297# 1 2 7 11 14
c19 11 0 1.38609e-19 $X=5.01 $Y=1.96
c20 2 0 1.6626e-19 $X=4.865 $Y=1.485
r21 14 16 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.07 $Y=2.3 $X2=4.07
+ $Y2=2.38
r22 9 11 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.01 $Y=2.295
+ $X2=5.01 $Y2=1.96
r23 8 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.195 $Y=2.38
+ $X2=4.07 $Y2=2.38
r24 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.885 $Y=2.38
+ $X2=5.01 $Y2=2.295
r25 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.885 $Y=2.38 $X2=4.195
+ $Y2=2.38
r26 2 11 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=1.96
r27 1 14 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_4%X 1 2 3 4 15 19 21 22 23 24 27 31 33 35
+ 37 38 44 45 48
c80 44 0 1.66154e-19 $X=7.59 $Y=1.19
c81 24 0 7.88531e-20 $X=6.115 $Y=0.815
r82 45 48 2.86169 $w=3.65e-07 $l=1.2e-07 $layer=LI1_cond $X=7.492 $Y=1.535
+ $X2=7.492 $Y2=1.415
r83 44 48 7.1041 $w=3.63e-07 $l=2.25e-07 $layer=LI1_cond $X=7.492 $Y=1.19
+ $X2=7.492 $Y2=1.415
r84 43 44 8.99853 $w=3.63e-07 $l=2.85e-07 $layer=LI1_cond $X=7.492 $Y=0.905
+ $X2=7.492 $Y2=1.19
r85 41 42 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=6.89 $Y=1.62
+ $X2=6.89 $Y2=1.87
r86 38 41 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=1.535
+ $X2=6.89 $Y2=1.62
r87 36 37 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=7.055 $Y=0.815
+ $X2=6.865 $Y2=0.815
r88 35 43 7.89155 $w=1.8e-07 $l=2.22495e-07 $layer=LI1_cond $X=7.31 $Y=0.815
+ $X2=7.492 $Y2=0.905
r89 35 36 15.7121 $w=1.78e-07 $l=2.55e-07 $layer=LI1_cond $X=7.31 $Y=0.815
+ $X2=7.055 $Y2=0.815
r90 34 38 0.964185 $w=2.4e-07 $l=1.25e-07 $layer=LI1_cond $X=7.015 $Y=1.535
+ $X2=6.89 $Y2=1.535
r91 33 45 4.34023 $w=2.4e-07 $l=1.82e-07 $layer=LI1_cond $X=7.31 $Y=1.535
+ $X2=7.492 $Y2=1.535
r92 33 34 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=7.31 $Y=1.535
+ $X2=7.015 $Y2=1.535
r93 29 42 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=1.955
+ $X2=6.89 $Y2=1.87
r94 29 31 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=6.89 $Y=1.955
+ $X2=6.89 $Y2=1.96
r95 25 37 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=6.865 $Y=0.725
+ $X2=6.865 $Y2=0.815
r96 25 27 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.865 $Y=0.725
+ $X2=6.865 $Y2=0.39
r97 23 37 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.675 $Y=0.815
+ $X2=6.865 $Y2=0.815
r98 23 24 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=6.675 $Y=0.815
+ $X2=6.115 $Y2=0.815
r99 21 42 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.765 $Y=1.87
+ $X2=6.89 $Y2=1.87
r100 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.765 $Y=1.87
+ $X2=6.075 $Y2=1.87
r101 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.95 $Y=1.955
+ $X2=6.075 $Y2=1.87
r102 17 19 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=5.95 $Y=1.955
+ $X2=5.95 $Y2=1.96
r103 13 24 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=5.925 $Y=0.725
+ $X2=6.115 $Y2=0.815
r104 13 15 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.925 $Y=0.725
+ $X2=5.925 $Y2=0.39
r105 4 41 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=1.62
r106 4 31 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=1.96
r107 3 19 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=1.96
r108 2 27 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=6.705
+ $Y=0.235 $X2=6.89 $Y2=0.39
r109 1 15 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=5.765
+ $Y=0.235 $X2=5.95 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_4%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44
+ 47 48 50 51 53 54 56 57 58 60 84 85 91 96 99
r125 98 99 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=0.235
+ $X2=3.685 $Y2=0.235
r126 94 98 2.80331 $w=6.38e-07 $l=1.5e-07 $layer=LI1_cond $X=3.45 $Y=0.235
+ $X2=3.6 $Y2=0.235
r127 94 96 15.8366 $w=6.38e-07 $l=4.55e-07 $layer=LI1_cond $X=3.45 $Y=0.235
+ $X2=2.995 $Y2=0.235
r128 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r129 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r130 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r131 82 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=7.59
+ $Y2=0
r132 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r133 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r134 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r135 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r136 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r137 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r138 73 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.45
+ $Y2=0
r139 72 99 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=4.37 $Y=0
+ $X2=3.685 $Y2=0
r140 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r141 69 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r142 69 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r143 68 96 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.99 $Y=0 $X2=2.995
+ $Y2=0
r144 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r145 66 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=0 $X2=2.14
+ $Y2=0
r146 66 68 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.225 $Y=0
+ $X2=2.99 $Y2=0
r147 64 92 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=2.07 $Y2=0
r148 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r149 61 88 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r150 61 63 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r151 60 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0 $X2=2.14
+ $Y2=0
r152 60 63 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=2.055 $Y=0
+ $X2=0.69 $Y2=0
r153 58 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r154 58 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r155 56 81 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.275 $Y=0
+ $X2=7.13 $Y2=0
r156 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.275 $Y=0 $X2=7.36
+ $Y2=0
r157 55 84 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.445 $Y=0
+ $X2=7.59 $Y2=0
r158 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.445 $Y=0 $X2=7.36
+ $Y2=0
r159 53 78 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.335 $Y=0
+ $X2=6.21 $Y2=0
r160 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.335 $Y=0 $X2=6.42
+ $Y2=0
r161 52 81 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=6.505 $Y=0
+ $X2=7.13 $Y2=0
r162 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.505 $Y=0 $X2=6.42
+ $Y2=0
r163 50 75 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=5.395 $Y=0
+ $X2=5.29 $Y2=0
r164 50 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=0 $X2=5.48
+ $Y2=0
r165 49 78 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=5.565 $Y=0
+ $X2=6.21 $Y2=0
r166 49 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=0 $X2=5.48
+ $Y2=0
r167 47 72 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=0 $X2=4.37
+ $Y2=0
r168 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=0 $X2=4.54
+ $Y2=0
r169 46 75 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.625 $Y=0 $X2=5.29
+ $Y2=0
r170 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=0 $X2=4.54
+ $Y2=0
r171 42 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0
r172 42 44 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0.39
r173 38 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0
r174 38 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0.39
r175 34 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0
r176 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.39
r177 30 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0
r178 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0.39
r179 26 91 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0
r180 26 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0.39
r181 22 88 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r182 22 24 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.39
r183 7 44 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.225
+ $Y=0.235 $X2=7.36 $Y2=0.39
r184 6 40 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=6.235
+ $Y=0.235 $X2=6.42 $Y2=0.39
r185 5 36 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.345
+ $Y=0.235 $X2=5.48 $Y2=0.39
r186 4 32 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.355
+ $Y=0.235 $X2=4.54 $Y2=0.39
r187 3 98 91 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_NDIFF $count=2 $X=2.945
+ $Y=0.235 $X2=3.6 $Y2=0.39
r188 2 28 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.39
r189 1 24 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_4%A_119_47# 1 2 7 9 13
c21 9 0 1.43173e-19 $X=0.73 $Y=0.73
r22 11 16 4.05488 $w=2.2e-07 $l=1.5e-07 $layer=LI1_cond $X=0.815 $Y=0.365
+ $X2=0.665 $Y2=0.365
r23 11 13 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=0.815 $Y=0.365
+ $X2=1.67 $Y2=0.365
r24 7 16 2.97358 $w=3e-07 $l=1.1e-07 $layer=LI1_cond $X=0.665 $Y=0.475 $X2=0.665
+ $Y2=0.365
r25 7 9 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=0.665 $Y=0.475
+ $X2=0.665 $Y2=0.73
r26 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.39
r27 1 16 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.39
r28 1 9 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.73
.ends

