* File: sky130_fd_sc_hdll__a31oi_4.pex.spice
* Created: Thu Aug 27 18:55:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A31OI_4%A3 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 27 28 45 54 58
r74 45 46 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=1.93 $Y2=1.202
r75 44 54 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.495 $Y=1.16
+ $X2=1.155 $Y2=1.16
r76 43 45 54.1425 $w=3.65e-07 $l=4.1e-07 $layer=POLY_cond $X=1.495 $Y=1.202
+ $X2=1.905 $Y2=1.202
r77 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.495
+ $Y=1.16 $X2=1.495 $Y2=1.16
r78 41 43 4.62192 $w=3.65e-07 $l=3.5e-08 $layer=POLY_cond $X=1.46 $Y=1.202
+ $X2=1.495 $Y2=1.202
r79 40 41 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.46 $Y2=1.202
r80 39 40 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=0.99 $Y=1.202
+ $X2=1.435 $Y2=1.202
r81 38 39 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r82 37 38 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.965 $Y2=1.202
r83 36 37 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r84 34 36 27.7315 $w=3.65e-07 $l=2.1e-07 $layer=POLY_cond $X=0.285 $Y=1.202
+ $X2=0.495 $Y2=1.202
r85 28 58 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=1.595 $Y=1.16
+ $X2=1.615 $Y2=1.16
r86 28 44 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.595 $Y=1.16
+ $X2=1.495 $Y2=1.16
r87 27 54 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.15 $Y=1.16
+ $X2=1.155 $Y2=1.16
r88 26 27 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=0.695 $Y=1.16
+ $X2=1.15 $Y2=1.16
r89 25 26 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=1.16
+ $X2=0.695 $Y2=1.16
r90 25 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.285
+ $Y=1.16 $X2=0.285 $Y2=1.16
r91 22 46 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r92 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r93 19 45 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r94 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r95 16 41 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=1.202
r96 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=0.56
r97 13 40 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r98 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r99 10 39 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r100 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r101 7 38 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r102 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r103 4 37 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r104 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=0.56
r105 1 36 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r106 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_4%A2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 27 28 45 48 54 57 61
r74 45 46 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.785 $Y=1.202
+ $X2=3.81 $Y2=1.202
r75 44 57 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=3.67 $Y=1.16
+ $X2=3.455 $Y2=1.16
r76 43 45 14.9005 $w=3.72e-07 $l=1.15e-07 $layer=POLY_cond $X=3.67 $Y=1.202
+ $X2=3.785 $Y2=1.202
r77 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.67
+ $Y=1.16 $X2=3.67 $Y2=1.16
r78 41 43 45.9973 $w=3.72e-07 $l=3.55e-07 $layer=POLY_cond $X=3.315 $Y=1.202
+ $X2=3.67 $Y2=1.202
r79 40 41 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.202
+ $X2=3.315 $Y2=1.202
r80 39 40 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=3.29 $Y2=1.202
r81 38 39 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.845 $Y2=1.202
r82 36 38 53.1237 $w=3.72e-07 $l=4.1e-07 $layer=POLY_cond $X=2.41 $Y=1.202
+ $X2=2.82 $Y2=1.202
r83 36 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.41
+ $Y=1.16 $X2=2.41 $Y2=1.16
r84 34 36 4.53495 $w=3.72e-07 $l=3.5e-08 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.41 $Y2=1.202
r85 33 34 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.202
+ $X2=2.375 $Y2=1.202
r86 28 61 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=3.865 $Y=1.16
+ $X2=3.875 $Y2=1.16
r87 28 44 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.865 $Y=1.16
+ $X2=3.67 $Y2=1.16
r88 27 57 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=3.445 $Y=1.16
+ $X2=3.455 $Y2=1.16
r89 27 54 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.445 $Y=1.16
+ $X2=2.995 $Y2=1.16
r90 26 54 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=2.975 $Y=1.16
+ $X2=2.995 $Y2=1.16
r91 25 26 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=2.52 $Y=1.16
+ $X2=2.975 $Y2=1.16
r92 25 48 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.52 $Y=1.16
+ $X2=2.33 $Y2=1.16
r93 22 46 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=1.202
r94 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=0.56
r95 19 45 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.202
r96 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r97 16 41 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.202
r98 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r99 13 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=1.202
r100 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=0.56
r101 10 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r102 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r103 7 38 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=1.202
r104 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=0.56
r105 4 34 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r106 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r107 1 33 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.202
r108 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_4%A1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 23 24 26 27 28 29 30 51 54 57 60
c76 30 0 1.6924e-19 $X=5.67 $Y=1.105
r77 46 47 13.3536 $w=3.79e-07 $l=1.05e-07 $layer=POLY_cond $X=5.685 $Y=1.202
+ $X2=5.79 $Y2=1.202
r78 45 60 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=5.57 $Y=1.16
+ $X2=5.75 $Y2=1.16
r79 45 57 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.57 $Y=1.16
+ $X2=5.315 $Y2=1.16
r80 44 46 14.6253 $w=3.79e-07 $l=1.15e-07 $layer=POLY_cond $X=5.57 $Y=1.202
+ $X2=5.685 $Y2=1.202
r81 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.57
+ $Y=1.16 $X2=5.57 $Y2=1.16
r82 42 44 31.7942 $w=3.79e-07 $l=2.5e-07 $layer=POLY_cond $X=5.32 $Y=1.202
+ $X2=5.57 $Y2=1.202
r83 41 42 13.3536 $w=3.79e-07 $l=1.05e-07 $layer=POLY_cond $X=5.215 $Y=1.202
+ $X2=5.32 $Y2=1.202
r84 40 41 46.4195 $w=3.79e-07 $l=3.65e-07 $layer=POLY_cond $X=4.85 $Y=1.202
+ $X2=5.215 $Y2=1.202
r85 39 40 13.3536 $w=3.79e-07 $l=1.05e-07 $layer=POLY_cond $X=4.745 $Y=1.202
+ $X2=4.85 $Y2=1.202
r86 37 39 55.3219 $w=3.79e-07 $l=4.35e-07 $layer=POLY_cond $X=4.31 $Y=1.202
+ $X2=4.745 $Y2=1.202
r87 35 37 4.45119 $w=3.79e-07 $l=3.5e-08 $layer=POLY_cond $X=4.275 $Y=1.202
+ $X2=4.31 $Y2=1.202
r88 30 60 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=5.755 $Y=1.16
+ $X2=5.75 $Y2=1.16
r89 29 57 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.3 $Y=1.16
+ $X2=5.315 $Y2=1.16
r90 29 54 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=5.3 $Y=1.16
+ $X2=4.855 $Y2=1.16
r91 28 54 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=4.845 $Y=1.16
+ $X2=4.855 $Y2=1.16
r92 28 51 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.845 $Y=1.16
+ $X2=4.395 $Y2=1.16
r93 27 51 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.31 $Y=1.16
+ $X2=4.395 $Y2=1.16
r94 27 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.31
+ $Y=1.16 $X2=4.31 $Y2=1.16
r95 24 26 144.6 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=6.26 $Y=1.01 $X2=6.26
+ $Y2=0.56
r96 23 47 11.055 $w=3.79e-07 $l=9.08295e-08 $layer=POLY_cond $X=5.865 $Y=1.167
+ $X2=5.79 $Y2=1.202
r97 22 24 31.5954 $w=3.15e-07 $l=1.90851e-07 $layer=POLY_cond $X=6.185 $Y=1.167
+ $X2=6.26 $Y2=1.01
r98 22 23 58.6202 $w=3.15e-07 $l=3.2e-07 $layer=POLY_cond $X=6.185 $Y=1.167
+ $X2=5.865 $Y2=1.167
r99 19 47 24.5487 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.79 $Y=0.995
+ $X2=5.79 $Y2=1.202
r100 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.79 $Y=0.995
+ $X2=5.79 $Y2=0.56
r101 16 46 20.1817 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.685 $Y=1.41
+ $X2=5.685 $Y2=1.202
r102 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.685 $Y=1.41
+ $X2=5.685 $Y2=1.985
r103 13 42 24.5487 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.32 $Y=0.995
+ $X2=5.32 $Y2=1.202
r104 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.32 $Y=0.995
+ $X2=5.32 $Y2=0.56
r105 10 41 20.1817 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.215 $Y=1.41
+ $X2=5.215 $Y2=1.202
r106 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.215 $Y=1.41
+ $X2=5.215 $Y2=1.985
r107 7 40 24.5487 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.85 $Y=0.995
+ $X2=4.85 $Y2=1.202
r108 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.85 $Y=0.995
+ $X2=4.85 $Y2=0.56
r109 4 39 20.1817 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.745 $Y=1.41
+ $X2=4.745 $Y2=1.202
r110 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.745 $Y=1.41
+ $X2=4.745 $Y2=1.985
r111 1 35 20.1817 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.275 $Y=1.41
+ $X2=4.275 $Y2=1.202
r112 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.275 $Y=1.41
+ $X2=4.275 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_4%B1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 29 49 54 57 61
c77 49 0 1.6924e-19 $X=8.115 $Y=1.202
r78 54 57 8.09943 $w=6.33e-07 $l=4.3e-07 $layer=LI1_cond $X=6.68 $Y=1.312
+ $X2=7.11 $Y2=1.312
r79 49 50 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=8.115 $Y=1.202
+ $X2=8.14 $Y2=1.202
r80 48 49 57.9703 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=7.67 $Y=1.202
+ $X2=8.115 $Y2=1.202
r81 47 48 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=7.645 $Y=1.202
+ $X2=7.67 $Y2=1.202
r82 45 47 16.2838 $w=3.7e-07 $l=1.25e-07 $layer=POLY_cond $X=7.52 $Y=1.202
+ $X2=7.645 $Y2=1.202
r83 43 45 41.6865 $w=3.7e-07 $l=3.2e-07 $layer=POLY_cond $X=7.2 $Y=1.202
+ $X2=7.52 $Y2=1.202
r84 42 43 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=7.175 $Y=1.202
+ $X2=7.2 $Y2=1.202
r85 41 42 57.9703 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=6.73 $Y=1.202
+ $X2=7.175 $Y2=1.202
r86 40 41 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=6.705 $Y=1.202
+ $X2=6.73 $Y2=1.202
r87 38 40 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=6.68 $Y=1.202
+ $X2=6.705 $Y2=1.202
r88 38 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.68
+ $Y=1.16 $X2=6.68 $Y2=1.16
r89 29 61 1.13015 $w=6.33e-07 $l=6e-08 $layer=LI1_cond $X=7.52 $Y=1.312 $X2=7.46
+ $Y2=1.312
r90 29 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.52
+ $Y=1.16 $X2=7.52 $Y2=1.16
r91 27 61 6.02748 $w=6.33e-07 $l=3.2e-07 $layer=LI1_cond $X=7.14 $Y=1.312
+ $X2=7.46 $Y2=1.312
r92 27 57 0.565076 $w=6.33e-07 $l=3e-08 $layer=LI1_cond $X=7.14 $Y=1.312
+ $X2=7.11 $Y2=1.312
r93 25 54 0.0941794 $w=6.33e-07 $l=5e-09 $layer=LI1_cond $X=6.675 $Y=1.312
+ $X2=6.68 $Y2=1.312
r94 22 50 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.14 $Y=0.995
+ $X2=8.14 $Y2=1.202
r95 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.14 $Y=0.995
+ $X2=8.14 $Y2=0.56
r96 19 49 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.115 $Y=1.41
+ $X2=8.115 $Y2=1.202
r97 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.115 $Y=1.41
+ $X2=8.115 $Y2=1.985
r98 16 48 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.67 $Y=0.995
+ $X2=7.67 $Y2=1.202
r99 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.67 $Y=0.995
+ $X2=7.67 $Y2=0.56
r100 13 47 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.645 $Y=1.41
+ $X2=7.645 $Y2=1.202
r101 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.645 $Y=1.41
+ $X2=7.645 $Y2=1.985
r102 10 43 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.2 $Y=0.995
+ $X2=7.2 $Y2=1.202
r103 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.2 $Y=0.995
+ $X2=7.2 $Y2=0.56
r104 7 42 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.175 $Y=1.41
+ $X2=7.175 $Y2=1.202
r105 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.175 $Y=1.41
+ $X2=7.175 $Y2=1.985
r106 4 41 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.73 $Y=0.995
+ $X2=6.73 $Y2=1.202
r107 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.73 $Y=0.995
+ $X2=6.73 $Y2=0.56
r108 1 40 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.705 $Y=1.41
+ $X2=6.705 $Y2=1.202
r109 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.705 $Y=1.41
+ $X2=6.705 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_4%A_27_297# 1 2 3 4 5 6 7 8 9 30 32 33 36 38
+ 42 44 48 50 54 56 60 62 67 68 69 72 74 76 77 78 79 80
r115 72 82 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.39 $Y=2.255
+ $X2=8.39 $Y2=2.34
r116 72 74 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=8.39 $Y=2.255
+ $X2=8.39 $Y2=1.66
r117 69 71 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=6.005 $Y=2.34
+ $X2=7.41 $Y2=2.34
r118 68 82 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.265 $Y=2.34
+ $X2=8.39 $Y2=2.34
r119 68 71 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=8.265 $Y=2.34
+ $X2=7.41 $Y2=2.34
r120 65 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.92 $Y=2.255
+ $X2=6.005 $Y2=2.34
r121 65 67 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=5.92 $Y=2.255
+ $X2=5.92 $Y2=1.8
r122 64 67 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.92 $Y=1.665
+ $X2=5.92 $Y2=1.8
r123 63 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=1.58
+ $X2=4.98 $Y2=1.58
r124 62 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.835 $Y=1.58
+ $X2=5.92 $Y2=1.665
r125 62 63 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.835 $Y=1.58
+ $X2=5.065 $Y2=1.58
r126 58 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=1.665
+ $X2=4.98 $Y2=1.58
r127 58 60 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.98 $Y=1.665
+ $X2=4.98 $Y2=1.96
r128 57 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=1.58
+ $X2=4.02 $Y2=1.58
r129 56 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=1.58
+ $X2=4.98 $Y2=1.58
r130 56 57 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.895 $Y=1.58
+ $X2=4.105 $Y2=1.58
r131 52 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=1.665
+ $X2=4.02 $Y2=1.58
r132 52 54 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.02 $Y=1.665
+ $X2=4.02 $Y2=1.96
r133 51 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=1.58
+ $X2=3.08 $Y2=1.58
r134 50 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=1.58
+ $X2=4.02 $Y2=1.58
r135 50 51 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.935 $Y=1.58
+ $X2=3.165 $Y2=1.58
r136 46 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=1.665
+ $X2=3.08 $Y2=1.58
r137 46 48 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.08 $Y=1.665
+ $X2=3.08 $Y2=1.96
r138 45 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=1.58
+ $X2=2.14 $Y2=1.58
r139 44 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=1.58
+ $X2=3.08 $Y2=1.58
r140 44 45 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.995 $Y=1.58
+ $X2=2.225 $Y2=1.58
r141 40 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=1.665
+ $X2=2.14 $Y2=1.58
r142 40 42 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.14 $Y=1.665
+ $X2=2.14 $Y2=1.96
r143 39 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=1.58
+ $X2=1.2 $Y2=1.58
r144 38 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=1.58
+ $X2=2.14 $Y2=1.58
r145 38 39 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=1.58
+ $X2=1.285 $Y2=1.58
r146 34 76 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=1.665 $X2=1.2
+ $Y2=1.58
r147 34 36 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=1.665
+ $X2=1.2 $Y2=1.96
r148 32 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=1.58
+ $X2=1.2 $Y2=1.58
r149 32 33 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=1.58
+ $X2=0.345 $Y2=1.58
r150 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.345 $Y2=1.58
r151 28 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=1.96
r152 9 82 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=8.205
+ $Y=1.485 $X2=8.35 $Y2=2.34
r153 9 74 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=8.205
+ $Y=1.485 $X2=8.35 $Y2=1.66
r154 8 71 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.265
+ $Y=1.485 $X2=7.41 $Y2=2.34
r155 7 67 300 $w=1.7e-07 $l=3.80657e-07 $layer=licon1_PDIFF $count=2 $X=5.775
+ $Y=1.485 $X2=5.92 $Y2=1.8
r156 6 60 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.835
+ $Y=1.485 $X2=4.98 $Y2=1.96
r157 5 54 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=1.96
r158 4 48 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=1.96
r159 3 42 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.96
r160 2 36 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.96
r161 1 30 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_4%VPWR 1 2 3 4 5 6 21 25 29 33 35 39 41 43
+ 45 50 55 60 70 71 74 77 80 83 86 89
r127 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r128 89 92 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=5.425 $Y=2.34
+ $X2=5.425 $Y2=2.72
r129 87 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r130 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r131 84 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r132 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r133 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r134 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r135 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r136 70 71 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r137 68 71 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=8.51 $Y2=2.72
r138 68 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r139 67 70 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=5.75 $Y=2.72
+ $X2=8.51 $Y2=2.72
r140 67 68 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r141 65 92 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.615 $Y=2.72
+ $X2=5.425 $Y2=2.72
r142 65 67 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.615 $Y=2.72
+ $X2=5.75 $Y2=2.72
r143 64 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r144 64 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r145 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r146 61 80 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=2.72
+ $X2=2.585 $Y2=2.72
r147 61 63 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.775 $Y=2.72
+ $X2=2.99 $Y2=2.72
r148 60 83 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.335 $Y=2.72
+ $X2=3.525 $Y2=2.72
r149 60 63 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.335 $Y=2.72
+ $X2=2.99 $Y2=2.72
r150 59 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r151 59 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r152 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r153 56 77 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=2.72
+ $X2=1.645 $Y2=2.72
r154 56 58 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.835 $Y=2.72
+ $X2=2.07 $Y2=2.72
r155 55 80 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=2.72
+ $X2=2.585 $Y2=2.72
r156 55 58 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.395 $Y=2.72
+ $X2=2.07 $Y2=2.72
r157 54 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r158 54 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r159 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r160 51 74 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r161 51 53 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r162 50 77 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.645 $Y2=2.72
r163 50 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r164 45 74 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r165 45 47 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r166 43 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r167 43 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r168 42 86 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.675 $Y=2.72
+ $X2=4.485 $Y2=2.72
r169 41 92 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.235 $Y=2.72
+ $X2=5.425 $Y2=2.72
r170 41 42 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.235 $Y=2.72
+ $X2=4.675 $Y2=2.72
r171 37 86 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.485 $Y=2.635
+ $X2=4.485 $Y2=2.72
r172 37 39 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=4.485 $Y=2.635
+ $X2=4.485 $Y2=2
r173 36 83 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.715 $Y=2.72
+ $X2=3.525 $Y2=2.72
r174 35 86 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.295 $Y=2.72
+ $X2=4.485 $Y2=2.72
r175 35 36 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.295 $Y=2.72
+ $X2=3.715 $Y2=2.72
r176 31 83 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=2.635
+ $X2=3.525 $Y2=2.72
r177 31 33 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=3.525 $Y=2.635
+ $X2=3.525 $Y2=2
r178 27 80 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=2.635
+ $X2=2.585 $Y2=2.72
r179 27 29 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.585 $Y=2.635
+ $X2=2.585 $Y2=2
r180 23 77 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=2.635
+ $X2=1.645 $Y2=2.72
r181 23 25 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=1.645 $Y=2.635
+ $X2=1.645 $Y2=2
r182 19 74 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r183 19 21 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2
r184 6 89 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.305
+ $Y=1.485 $X2=5.45 $Y2=2.34
r185 5 39 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.365
+ $Y=1.485 $X2=4.51 $Y2=2
r186 4 33 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2
r187 3 29 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2
r188 2 25 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2
r189 1 21 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_4%Y 1 2 3 4 5 6 7 22 30 36 38 40 44 46 47 48
+ 49 50 58 60 68
r76 58 68 2.16083 $w=2.38e-07 $l=4.5e-08 $layer=LI1_cond $X=7.965 $Y=1.915
+ $X2=7.965 $Y2=1.87
r77 57 60 2.16083 $w=2.38e-07 $l=4.5e-08 $layer=LI1_cond $X=7.965 $Y=0.805
+ $X2=7.965 $Y2=0.85
r78 50 58 2.93484 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=7.965 $Y=2 $X2=7.965
+ $Y2=1.915
r79 50 68 0.960369 $w=2.38e-07 $l=2e-08 $layer=LI1_cond $X=7.965 $Y=1.85
+ $X2=7.965 $Y2=1.87
r80 49 50 15.3659 $w=2.38e-07 $l=3.2e-07 $layer=LI1_cond $X=7.965 $Y=1.53
+ $X2=7.965 $Y2=1.85
r81 48 49 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=7.965 $Y=1.19
+ $X2=7.965 $Y2=1.53
r82 47 57 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=7.965 $Y=0.72
+ $X2=7.965 $Y2=0.805
r83 47 48 15.3659 $w=2.38e-07 $l=3.2e-07 $layer=LI1_cond $X=7.965 $Y=0.87
+ $X2=7.965 $Y2=1.19
r84 47 60 0.960369 $w=2.38e-07 $l=2e-08 $layer=LI1_cond $X=7.965 $Y=0.87
+ $X2=7.965 $Y2=0.85
r85 42 44 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=8.35 $Y=0.635
+ $X2=8.35 $Y2=0.42
r86 41 47 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=8.085 $Y=0.72
+ $X2=7.965 $Y2=0.72
r87 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.265 $Y=0.72
+ $X2=8.35 $Y2=0.635
r88 40 41 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.265 $Y=0.72
+ $X2=8.085 $Y2=0.72
r89 39 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.495 $Y=0.72
+ $X2=7.41 $Y2=0.72
r90 38 47 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.845 $Y=0.72
+ $X2=7.965 $Y2=0.72
r91 38 39 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.845 $Y=0.72
+ $X2=7.495 $Y2=0.72
r92 34 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.41 $Y=0.635
+ $X2=7.41 $Y2=0.72
r93 34 36 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=7.41 $Y=0.635
+ $X2=7.41 $Y2=0.42
r94 30 50 4.1433 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.845 $Y=2 $X2=7.965
+ $Y2=2
r95 30 32 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=7.845 $Y=2 $X2=6.94
+ $Y2=2
r96 27 29 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=5.53 $Y=0.72
+ $X2=6.47 $Y2=0.72
r97 24 27 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=4.59 $Y=0.72
+ $X2=5.53 $Y2=0.72
r98 22 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.325 $Y=0.72
+ $X2=7.41 $Y2=0.72
r99 22 29 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=7.325 $Y=0.72
+ $X2=6.47 $Y2=0.72
r100 7 50 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=7.735
+ $Y=1.485 $X2=7.88 $Y2=2
r101 6 32 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=6.795
+ $Y=1.485 $X2=6.94 $Y2=2
r102 5 44 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=8.215
+ $Y=0.235 $X2=8.35 $Y2=0.42
r103 4 36 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=7.275
+ $Y=0.235 $X2=7.41 $Y2=0.42
r104 3 29 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=6.335
+ $Y=0.235 $X2=6.47 $Y2=0.72
r105 2 27 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=5.395
+ $Y=0.235 $X2=5.53 $Y2=0.72
r106 1 24 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=4.465
+ $Y=0.235 $X2=4.59 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_4%A_27_47# 1 2 3 4 5 18 20 21 24 26 30 36 38
+ 39
r54 34 36 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.08 $Y=0.72
+ $X2=4.02 $Y2=0.72
r55 32 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=0.72
+ $X2=2.14 $Y2=0.72
r56 32 34 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=2.225 $Y=0.72
+ $X2=3.08 $Y2=0.72
r57 28 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.635
+ $X2=2.14 $Y2=0.72
r58 28 30 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.14 $Y=0.635
+ $X2=2.14 $Y2=0.42
r59 27 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=0.72 $X2=1.2
+ $Y2=0.72
r60 26 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0.72
+ $X2=2.14 $Y2=0.72
r61 26 27 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=0.72
+ $X2=1.285 $Y2=0.72
r62 22 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.635 $X2=1.2
+ $Y2=0.72
r63 22 24 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.2 $Y=0.635
+ $X2=1.2 $Y2=0.42
r64 20 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0.72 $X2=1.2
+ $Y2=0.72
r65 20 21 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=0.72
+ $X2=0.345 $Y2=0.72
r66 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r67 16 18 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.42
r68 5 36 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.235 $X2=4.02 $Y2=0.72
r69 4 34 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.72
r70 3 30 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.42
r71 2 24 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.42
r72 1 18 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_4%VGND 1 2 3 4 13 14 20 21 27 29 34 50 51 55
+ 62
r111 62 65 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=1.645 $Y=0
+ $X2=1.645 $Y2=0.38
r112 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r113 55 58 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.38
r114 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r115 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r116 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.51
+ $Y2=0
r117 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r118 45 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.59
+ $Y2=0
r119 44 45 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r120 42 45 1.30889 $w=4.8e-07 $l=4.6e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=6.67
+ $Y2=0
r121 42 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r122 41 44 300.107 $w=1.68e-07 $l=4.6e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=6.67
+ $Y2=0
r123 41 42 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r124 39 62 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=1.645
+ $Y2=0
r125 39 41 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.835 $Y=0
+ $X2=2.07 $Y2=0
r126 38 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r127 38 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r128 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r129 35 55 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r130 35 37 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r131 34 62 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.645
+ $Y2=0
r132 34 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r133 29 55 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r134 29 31 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r135 27 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r136 27 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r137 23 50 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=8.045 $Y=0
+ $X2=8.51 $Y2=0
r138 21 47 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=7.665 $Y=0 $X2=7.59
+ $Y2=0
r139 20 25 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=7.855 $Y=0
+ $X2=7.855 $Y2=0.38
r140 20 23 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.855 $Y=0 $X2=8.045
+ $Y2=0
r141 20 21 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.855 $Y=0 $X2=7.665
+ $Y2=0
r142 16 47 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=7.105 $Y=0
+ $X2=7.59 $Y2=0
r143 14 44 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=6.725 $Y=0 $X2=6.67
+ $Y2=0
r144 13 18 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=6.915 $Y=0
+ $X2=6.915 $Y2=0.38
r145 13 16 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.915 $Y=0 $X2=7.105
+ $Y2=0
r146 13 14 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.915 $Y=0 $X2=6.725
+ $Y2=0
r147 4 25 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.745
+ $Y=0.235 $X2=7.88 $Y2=0.38
r148 3 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.805
+ $Y=0.235 $X2=6.94 $Y2=0.38
r149 2 65 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.38
r150 1 58 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_4%A_485_47# 1 2 3 4 21
r26 19 21 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=5.06 $Y=0.38 $X2=6
+ $Y2=0.38
r27 17 19 98.5134 $w=1.68e-07 $l=1.51e-06 $layer=LI1_cond $X=3.55 $Y=0.38
+ $X2=5.06 $Y2=0.38
r28 14 17 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=2.61 $Y=0.38
+ $X2=3.55 $Y2=0.38
r29 4 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.865
+ $Y=0.235 $X2=6 $Y2=0.38
r30 3 19 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.925
+ $Y=0.235 $X2=5.06 $Y2=0.38
r31 2 17 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.38
r32 1 14 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.38
.ends

