* File: sky130_fd_sc_hdll__o221ai_1.pxi.spice
* Created: Wed Sep  2 08:44:52 2020
* 
x_PM_SKY130_FD_SC_HDLL__O221AI_1%C1 N_C1_c_49_n N_C1_M1001_g N_C1_c_50_n
+ N_C1_M1004_g C1 N_C1_c_51_n PM_SKY130_FD_SC_HDLL__O221AI_1%C1
x_PM_SKY130_FD_SC_HDLL__O221AI_1%B1 N_B1_c_74_n N_B1_M1009_g N_B1_c_75_n
+ N_B1_M1007_g B1 N_B1_c_76_n B1 PM_SKY130_FD_SC_HDLL__O221AI_1%B1
x_PM_SKY130_FD_SC_HDLL__O221AI_1%B2 N_B2_c_99_n N_B2_M1000_g N_B2_c_100_n
+ N_B2_M1005_g B2 B2 PM_SKY130_FD_SC_HDLL__O221AI_1%B2
x_PM_SKY130_FD_SC_HDLL__O221AI_1%A2 N_A2_c_133_n N_A2_M1008_g N_A2_c_134_n
+ N_A2_M1002_g N_A2_c_135_n N_A2_c_136_n N_A2_c_139_n A2
+ PM_SKY130_FD_SC_HDLL__O221AI_1%A2
x_PM_SKY130_FD_SC_HDLL__O221AI_1%A1 N_A1_c_179_n N_A1_M1006_g N_A1_c_180_n
+ N_A1_M1003_g A1 A1 PM_SKY130_FD_SC_HDLL__O221AI_1%A1
x_PM_SKY130_FD_SC_HDLL__O221AI_1%Y N_Y_M1004_s N_Y_M1001_s N_Y_M1000_d
+ N_Y_c_203_n N_Y_c_206_n N_Y_c_207_n N_Y_c_212_n N_Y_c_204_n N_Y_c_217_n
+ N_Y_c_205_n N_Y_c_224_n N_Y_c_238_p N_Y_c_228_n Y Y Y
+ PM_SKY130_FD_SC_HDLL__O221AI_1%Y
x_PM_SKY130_FD_SC_HDLL__O221AI_1%VPWR N_VPWR_M1001_d N_VPWR_M1003_d
+ N_VPWR_c_267_n N_VPWR_c_268_n VPWR N_VPWR_c_269_n N_VPWR_c_270_n
+ N_VPWR_c_271_n N_VPWR_c_266_n PM_SKY130_FD_SC_HDLL__O221AI_1%VPWR
x_PM_SKY130_FD_SC_HDLL__O221AI_1%A_123_47# N_A_123_47#_M1004_d
+ N_A_123_47#_M1007_d N_A_123_47#_c_317_n
+ PM_SKY130_FD_SC_HDLL__O221AI_1%A_123_47#
x_PM_SKY130_FD_SC_HDLL__O221AI_1%A_261_47# N_A_261_47#_M1007_s
+ N_A_261_47#_M1005_d N_A_261_47#_M1006_d N_A_261_47#_c_332_n
+ N_A_261_47#_c_333_n N_A_261_47#_c_334_n N_A_261_47#_c_342_n
+ PM_SKY130_FD_SC_HDLL__O221AI_1%A_261_47#
x_PM_SKY130_FD_SC_HDLL__O221AI_1%VGND N_VGND_M1008_d N_VGND_c_377_n
+ N_VGND_c_378_n N_VGND_c_379_n VGND N_VGND_c_380_n N_VGND_c_381_n
+ PM_SKY130_FD_SC_HDLL__O221AI_1%VGND
cc_1 VNB N_C1_c_49_n 0.0336232f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_2 VNB N_C1_c_50_n 0.0251465f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_3 VNB N_C1_c_51_n 0.013208f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.16
cc_4 VNB N_B1_c_74_n 0.0330519f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_5 VNB N_B1_c_75_n 0.022682f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_6 VNB N_B1_c_76_n 0.00888426f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.16
cc_7 VNB N_B2_c_99_n 0.0215105f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_8 VNB N_B2_c_100_n 0.0181387f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_9 VNB B2 0.00627491f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_10 VNB N_A2_c_133_n 0.0176822f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_11 VNB N_A2_c_134_n 0.0223238f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_12 VNB N_A2_c_135_n 4.82646e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A2_c_136_n 0.0037596f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.16
cc_14 VNB N_A1_c_179_n 0.0222254f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_15 VNB N_A1_c_180_n 0.0388902f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_16 VNB A1 0.00968497f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_17 VNB N_Y_c_203_n 0.011033f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.16
cc_18 VNB N_Y_c_204_n 0.00810425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_Y_c_205_n 0.0110591f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_266_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_123_47#_c_317_n 0.0148006f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.16
cc_22 VNB N_A_261_47#_c_332_n 0.00322242f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.16
cc_23 VNB N_A_261_47#_c_333_n 0.00767792f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_261_47#_c_334_n 0.0168702f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_377_n 0.0046757f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.56
cc_26 VNB N_VGND_c_378_n 0.0722191f $X=-0.19 $Y=-0.24 $X2=0.43 $Y2=1.16
cc_27 VNB N_VGND_c_379_n 0.00324214f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.16
cc_28 VNB N_VGND_c_380_n 0.0191497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_381_n 0.204502f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VPB N_C1_c_49_n 0.0374f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_31 VPB N_C1_c_51_n 0.00220476f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.16
cc_32 VPB N_B1_c_74_n 0.0345199f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_33 VPB N_B1_c_76_n 0.00360343f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.16
cc_34 VPB N_B2_c_99_n 0.02754f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_35 VPB B2 0.00202999f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_36 VPB N_A2_c_134_n 0.0281047f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_37 VPB N_A2_c_135_n 0.00316612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A2_c_139_n 0.00343707f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A1_c_180_n 0.0380946f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_40 VPB N_Y_c_206_n 0.00939401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_Y_c_207_n 0.0294554f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.16
cc_42 VPB N_Y_c_205_n 0.00768942f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_267_n 0.0105255f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_44 VPB N_VPWR_c_268_n 0.0463965f $X=-0.19 $Y=1.305 $X2=0.43 $Y2=1.16
cc_45 VPB N_VPWR_c_269_n 0.0460005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_270_n 0.0175557f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_271_n 0.0205264f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_266_n 0.0439532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 N_C1_c_50_n N_Y_c_203_n 0.0087171f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_50 N_C1_c_49_n N_Y_c_206_n 0.00279548f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_51 N_C1_c_51_n N_Y_c_206_n 0.0238687f $X=0.38 $Y=1.16 $X2=0 $Y2=0
cc_52 N_C1_c_49_n N_Y_c_212_n 0.00273348f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_53 N_C1_c_50_n N_Y_c_212_n 0.016431f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_54 N_C1_c_51_n N_Y_c_212_n 0.00677361f $X=0.38 $Y=1.16 $X2=0 $Y2=0
cc_55 N_C1_c_49_n N_Y_c_204_n 0.00230026f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_56 N_C1_c_51_n N_Y_c_204_n 0.0215583f $X=0.38 $Y=1.16 $X2=0 $Y2=0
cc_57 N_C1_c_49_n N_Y_c_217_n 0.0210161f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_58 N_C1_c_51_n N_Y_c_217_n 0.00511762f $X=0.38 $Y=1.16 $X2=0 $Y2=0
cc_59 N_C1_c_49_n N_Y_c_205_n 0.00327408f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_60 N_C1_c_50_n N_Y_c_205_n 0.0187652f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_61 N_C1_c_51_n N_Y_c_205_n 0.0213426f $X=0.38 $Y=1.16 $X2=0 $Y2=0
cc_62 N_C1_c_49_n N_VPWR_c_270_n 0.00681171f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_63 N_C1_c_49_n N_VPWR_c_271_n 0.0135745f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_64 N_C1_c_49_n N_VPWR_c_266_n 0.0122036f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_65 N_C1_c_50_n N_A_123_47#_c_317_n 0.00726496f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_66 N_C1_c_50_n N_A_261_47#_c_332_n 8.55515e-19 $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_67 N_C1_c_50_n N_VGND_c_378_n 0.00387603f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_68 N_C1_c_50_n N_VGND_c_381_n 0.00783163f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_69 N_B1_c_74_n N_B2_c_99_n 0.0801501f $X=1.665 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_70 N_B1_c_76_n N_B2_c_99_n 2.3951e-19 $X=1.51 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_71 N_B1_c_75_n N_B2_c_100_n 0.0223719f $X=1.69 $Y=0.995 $X2=0 $Y2=0
cc_72 N_B1_c_74_n B2 0.00300535f $X=1.665 $Y=1.41 $X2=0 $Y2=0
cc_73 N_B1_c_76_n B2 0.0232491f $X=1.51 $Y=1.16 $X2=0 $Y2=0
cc_74 N_B1_c_74_n N_Y_c_205_n 0.0010765f $X=1.665 $Y=1.41 $X2=0 $Y2=0
cc_75 N_B1_c_76_n N_Y_c_205_n 0.0273405f $X=1.51 $Y=1.16 $X2=0 $Y2=0
cc_76 N_B1_c_74_n N_Y_c_224_n 0.027895f $X=1.665 $Y=1.41 $X2=0 $Y2=0
cc_77 N_B1_c_76_n N_Y_c_224_n 0.0427987f $X=1.51 $Y=1.16 $X2=0 $Y2=0
cc_78 N_B1_c_74_n Y 0.00976295f $X=1.665 $Y=1.41 $X2=0 $Y2=0
cc_79 N_B1_c_74_n N_VPWR_c_269_n 0.00681171f $X=1.665 $Y=1.41 $X2=0 $Y2=0
cc_80 N_B1_c_74_n N_VPWR_c_271_n 0.0138231f $X=1.665 $Y=1.41 $X2=0 $Y2=0
cc_81 N_B1_c_74_n N_VPWR_c_266_n 0.0113016f $X=1.665 $Y=1.41 $X2=0 $Y2=0
cc_82 N_B1_c_75_n N_A_123_47#_c_317_n 0.0100597f $X=1.69 $Y=0.995 $X2=0 $Y2=0
cc_83 N_B1_c_76_n N_A_123_47#_c_317_n 0.00859171f $X=1.51 $Y=1.16 $X2=0 $Y2=0
cc_84 N_B1_c_74_n N_A_261_47#_c_332_n 0.00542966f $X=1.665 $Y=1.41 $X2=0 $Y2=0
cc_85 N_B1_c_75_n N_A_261_47#_c_332_n 0.0111261f $X=1.69 $Y=0.995 $X2=0 $Y2=0
cc_86 N_B1_c_76_n N_A_261_47#_c_332_n 0.0248151f $X=1.51 $Y=1.16 $X2=0 $Y2=0
cc_87 N_B1_c_75_n N_VGND_c_378_n 0.00368123f $X=1.69 $Y=0.995 $X2=0 $Y2=0
cc_88 N_B1_c_75_n N_VGND_c_381_n 0.00676883f $X=1.69 $Y=0.995 $X2=0 $Y2=0
cc_89 N_B2_c_100_n N_A2_c_133_n 0.0186073f $X=2.16 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_90 N_B2_c_99_n N_A2_c_134_n 0.0371613f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_91 B2 N_A2_c_134_n 0.00105444f $X=1.995 $Y=1.105 $X2=0 $Y2=0
cc_92 N_B2_c_99_n N_A2_c_135_n 0.00222533f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_93 B2 N_A2_c_135_n 0.00371474f $X=1.995 $Y=1.105 $X2=0 $Y2=0
cc_94 N_B2_c_99_n N_A2_c_136_n 5.84928e-19 $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_95 B2 N_A2_c_136_n 0.013542f $X=1.995 $Y=1.105 $X2=0 $Y2=0
cc_96 N_B2_c_99_n N_A2_c_139_n 7.64615e-19 $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_97 B2 N_Y_c_224_n 0.00668775f $X=1.995 $Y=1.105 $X2=0 $Y2=0
cc_98 N_B2_c_99_n N_Y_c_228_n 0.0112095f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_99 B2 N_Y_c_228_n 0.0298737f $X=1.995 $Y=1.105 $X2=0 $Y2=0
cc_100 N_B2_c_99_n Y 0.0108172f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_101 N_B2_c_99_n Y 0.00805122f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_102 N_B2_c_99_n N_VPWR_c_269_n 0.00429201f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_103 N_B2_c_99_n N_VPWR_c_271_n 0.00160636f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_104 N_B2_c_99_n N_VPWR_c_266_n 0.00640674f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_105 N_B2_c_99_n N_A_261_47#_c_332_n 0.00195591f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_106 N_B2_c_100_n N_A_261_47#_c_332_n 0.0103101f $X=2.16 $Y=0.995 $X2=0 $Y2=0
cc_107 B2 N_A_261_47#_c_332_n 0.0310568f $X=1.995 $Y=1.105 $X2=0 $Y2=0
cc_108 N_B2_c_99_n N_A_261_47#_c_342_n 9.04308e-19 $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_109 N_B2_c_100_n N_A_261_47#_c_342_n 9.70164e-19 $X=2.16 $Y=0.995 $X2=0 $Y2=0
cc_110 B2 N_A_261_47#_c_342_n 0.00294124f $X=1.995 $Y=1.105 $X2=0 $Y2=0
cc_111 N_B2_c_100_n N_VGND_c_378_n 0.00426565f $X=2.16 $Y=0.995 $X2=0 $Y2=0
cc_112 N_B2_c_100_n N_VGND_c_381_n 0.0063492f $X=2.16 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A2_c_133_n N_A1_c_179_n 0.0276478f $X=2.72 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_114 N_A2_c_134_n N_A1_c_180_n 0.093099f $X=2.755 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A2_c_135_n N_A1_c_180_n 0.00376404f $X=2.765 $Y=1.445 $X2=0 $Y2=0
cc_116 N_A2_c_136_n N_A1_c_180_n 6.59103e-19 $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A2_c_139_n N_A1_c_180_n 0.00541975f $X=2.99 $Y=1.615 $X2=0 $Y2=0
cc_118 A2 N_A1_c_180_n 0.017655f $X=2.91 $Y=1.785 $X2=0 $Y2=0
cc_119 N_A2_c_134_n A1 2.29876e-19 $X=2.755 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A2_c_136_n A1 0.0163554f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A2_c_139_n A1 0.00415563f $X=2.99 $Y=1.615 $X2=0 $Y2=0
cc_122 N_A2_c_134_n N_Y_c_228_n 0.00153889f $X=2.755 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A2_c_134_n Y 0.0051522f $X=2.755 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A2_c_134_n Y 0.00427606f $X=2.755 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A2_c_139_n N_VPWR_c_268_n 0.0115575f $X=2.99 $Y=1.615 $X2=0 $Y2=0
cc_126 A2 N_VPWR_c_268_n 0.0544438f $X=2.91 $Y=1.785 $X2=0 $Y2=0
cc_127 N_A2_c_134_n N_VPWR_c_269_n 0.00702461f $X=2.755 $Y=1.41 $X2=0 $Y2=0
cc_128 A2 N_VPWR_c_269_n 0.0109773f $X=2.91 $Y=1.785 $X2=0 $Y2=0
cc_129 N_A2_c_134_n N_VPWR_c_266_n 0.0130392f $X=2.755 $Y=1.41 $X2=0 $Y2=0
cc_130 A2 N_VPWR_c_266_n 0.00977549f $X=2.91 $Y=1.785 $X2=0 $Y2=0
cc_131 N_A2_c_139_n A_569_297# 3.43001e-19 $X=2.99 $Y=1.615 $X2=-0.19 $Y2=-0.24
cc_132 A2 A_569_297# 0.00163082f $X=2.91 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_133 N_A2_c_133_n N_A_261_47#_c_333_n 0.01269f $X=2.72 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A2_c_134_n N_A_261_47#_c_333_n 0.00336607f $X=2.755 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A2_c_136_n N_A_261_47#_c_333_n 0.0171794f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A2_c_139_n N_A_261_47#_c_333_n 0.00441919f $X=2.99 $Y=1.615 $X2=0 $Y2=0
cc_137 N_A2_c_133_n N_A_261_47#_c_334_n 5.29341e-19 $X=2.72 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A2_c_133_n N_A_261_47#_c_342_n 0.00502039f $X=2.72 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A2_c_134_n N_A_261_47#_c_342_n 6.24057e-19 $X=2.755 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A2_c_136_n N_A_261_47#_c_342_n 0.00370499f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A2_c_133_n N_VGND_c_377_n 0.00268723f $X=2.72 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A2_c_133_n N_VGND_c_378_n 0.00433717f $X=2.72 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A2_c_133_n N_VGND_c_381_n 0.00623009f $X=2.72 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A1_c_180_n N_VPWR_c_268_n 0.0154615f $X=3.165 $Y=1.41 $X2=0 $Y2=0
cc_145 A1 N_VPWR_c_268_n 0.0202856f $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_146 N_A1_c_180_n N_VPWR_c_269_n 0.00632076f $X=3.165 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A1_c_180_n N_VPWR_c_266_n 0.0115827f $X=3.165 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A1_c_179_n N_A_261_47#_c_333_n 0.00944054f $X=3.14 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A1_c_180_n N_A_261_47#_c_333_n 0.0080738f $X=3.165 $Y=1.41 $X2=0 $Y2=0
cc_150 A1 N_A_261_47#_c_333_n 0.0310137f $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_151 N_A1_c_179_n N_A_261_47#_c_334_n 0.00606965f $X=3.14 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A1_c_179_n N_VGND_c_377_n 0.00268723f $X=3.14 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A1_c_179_n N_VGND_c_380_n 0.00421028f $X=3.14 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A1_c_179_n N_VGND_c_381_n 0.00670066f $X=3.14 $Y=0.995 $X2=0 $Y2=0
cc_155 N_Y_c_217_n N_VPWR_M1001_d 3.69166e-19 $X=0.675 $Y=1.6 $X2=-0.19
+ $Y2=-0.24
cc_156 N_Y_c_205_n N_VPWR_M1001_d 4.7208e-19 $X=0.76 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_157 N_Y_c_224_n N_VPWR_M1001_d 0.025121f $X=1.9 $Y=1.6 $X2=-0.19 $Y2=-0.24
cc_158 N_Y_c_238_p N_VPWR_M1001_d 0.00256112f $X=0.76 $Y=1.6 $X2=-0.19 $Y2=-0.24
cc_159 Y N_VPWR_c_269_n 0.0378492f $X=2.09 $Y=2.21 $X2=0 $Y2=0
cc_160 N_Y_c_207_n N_VPWR_c_270_n 0.0196165f $X=0.28 $Y=1.96 $X2=0 $Y2=0
cc_161 N_Y_c_207_n N_VPWR_c_271_n 0.0373319f $X=0.28 $Y=1.96 $X2=0 $Y2=0
cc_162 N_Y_c_217_n N_VPWR_c_271_n 0.00137348f $X=0.675 $Y=1.6 $X2=0 $Y2=0
cc_163 N_Y_c_224_n N_VPWR_c_271_n 0.055606f $X=1.9 $Y=1.6 $X2=0 $Y2=0
cc_164 N_Y_c_238_p N_VPWR_c_271_n 0.0151701f $X=0.76 $Y=1.6 $X2=0 $Y2=0
cc_165 Y N_VPWR_c_271_n 0.0310773f $X=2 $Y=1.785 $X2=0 $Y2=0
cc_166 N_Y_M1001_s N_VPWR_c_266_n 0.00442207f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_167 N_Y_M1000_d N_VPWR_c_266_n 0.00937374f $X=2.195 $Y=1.485 $X2=0 $Y2=0
cc_168 N_Y_c_207_n N_VPWR_c_266_n 0.0107063f $X=0.28 $Y=1.96 $X2=0 $Y2=0
cc_169 Y N_VPWR_c_266_n 0.0222953f $X=2.09 $Y=2.21 $X2=0 $Y2=0
cc_170 N_Y_c_224_n A_351_297# 0.0043065f $X=1.9 $Y=1.6 $X2=-0.19 $Y2=-0.24
cc_171 N_Y_c_228_n A_351_297# 6.43421e-19 $X=2.182 $Y=1.705 $X2=-0.19 $Y2=-0.24
cc_172 Y A_351_297# 0.00562394f $X=2 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_173 Y A_351_297# 0.00374402f $X=2.09 $Y=2.21 $X2=-0.19 $Y2=-0.24
cc_174 N_Y_c_212_n N_A_123_47#_M1004_d 0.00531769f $X=0.675 $Y=0.735 $X2=-0.19
+ $Y2=-0.24
cc_175 N_Y_c_205_n N_A_123_47#_M1004_d 0.00306019f $X=0.76 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_176 N_Y_c_203_n N_A_123_47#_c_317_n 0.00882843f $X=0.215 $Y=0.645 $X2=0 $Y2=0
cc_177 N_Y_c_212_n N_A_123_47#_c_317_n 0.0196316f $X=0.675 $Y=0.735 $X2=0 $Y2=0
cc_178 N_Y_c_212_n N_A_261_47#_c_332_n 0.00876865f $X=0.675 $Y=0.735 $X2=0 $Y2=0
cc_179 N_Y_c_224_n N_A_261_47#_c_332_n 0.00343876f $X=1.9 $Y=1.6 $X2=0 $Y2=0
cc_180 N_Y_c_228_n N_A_261_47#_c_342_n 0.00442842f $X=2.182 $Y=1.705 $X2=0 $Y2=0
cc_181 N_Y_c_203_n N_VGND_c_378_n 0.0103423f $X=0.215 $Y=0.645 $X2=0 $Y2=0
cc_182 N_Y_c_212_n N_VGND_c_378_n 0.00242085f $X=0.675 $Y=0.735 $X2=0 $Y2=0
cc_183 N_Y_M1004_s N_VGND_c_381_n 0.00321876f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_184 N_Y_c_203_n N_VGND_c_381_n 0.00923165f $X=0.215 $Y=0.645 $X2=0 $Y2=0
cc_185 N_Y_c_212_n N_VGND_c_381_n 0.00480101f $X=0.675 $Y=0.735 $X2=0 $Y2=0
cc_186 N_VPWR_c_266_n A_351_297# 0.00715626f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_187 N_VPWR_c_266_n A_569_297# 0.00226512f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_188 N_A_123_47#_c_317_n N_A_261_47#_M1007_s 0.00633995f $X=1.9 $Y=0.39
+ $X2=-0.19 $Y2=-0.24
cc_189 N_A_123_47#_M1007_d N_A_261_47#_c_332_n 0.00426562f $X=1.765 $Y=0.235
+ $X2=0 $Y2=0
cc_190 N_A_123_47#_c_317_n N_A_261_47#_c_332_n 0.0454185f $X=1.9 $Y=0.39 $X2=0
+ $Y2=0
cc_191 N_A_123_47#_c_317_n N_VGND_c_378_n 0.0702277f $X=1.9 $Y=0.39 $X2=0 $Y2=0
cc_192 N_A_123_47#_M1004_d N_VGND_c_381_n 0.0021262f $X=0.615 $Y=0.235 $X2=0
+ $Y2=0
cc_193 N_A_123_47#_M1007_d N_VGND_c_381_n 0.00266367f $X=1.765 $Y=0.235 $X2=0
+ $Y2=0
cc_194 N_A_123_47#_c_317_n N_VGND_c_381_n 0.0546618f $X=1.9 $Y=0.39 $X2=0 $Y2=0
cc_195 N_A_261_47#_c_333_n N_VGND_M1008_d 0.00429463f $X=3.185 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_196 N_A_261_47#_c_333_n N_VGND_c_377_n 0.012114f $X=3.185 $Y=0.78 $X2=0 $Y2=0
cc_197 N_A_261_47#_c_332_n N_VGND_c_378_n 0.00306767f $X=2.285 $Y=0.735 $X2=0
+ $Y2=0
cc_198 N_A_261_47#_c_333_n N_VGND_c_378_n 0.00345506f $X=3.185 $Y=0.78 $X2=0
+ $Y2=0
cc_199 N_A_261_47#_c_342_n N_VGND_c_378_n 0.0161384f $X=2.37 $Y=0.66 $X2=0 $Y2=0
cc_200 N_A_261_47#_c_333_n N_VGND_c_380_n 0.00211912f $X=3.185 $Y=0.78 $X2=0
+ $Y2=0
cc_201 N_A_261_47#_c_334_n N_VGND_c_380_n 0.021576f $X=3.4 $Y=0.39 $X2=0 $Y2=0
cc_202 N_A_261_47#_M1007_s N_VGND_c_381_n 0.00255063f $X=1.305 $Y=0.235 $X2=0
+ $Y2=0
cc_203 N_A_261_47#_M1005_d N_VGND_c_381_n 0.00387059f $X=2.235 $Y=0.235 $X2=0
+ $Y2=0
cc_204 N_A_261_47#_M1006_d N_VGND_c_381_n 0.00251629f $X=3.215 $Y=0.235 $X2=0
+ $Y2=0
cc_205 N_A_261_47#_c_332_n N_VGND_c_381_n 0.00691149f $X=2.285 $Y=0.735 $X2=0
+ $Y2=0
cc_206 N_A_261_47#_c_333_n N_VGND_c_381_n 0.011534f $X=3.185 $Y=0.78 $X2=0 $Y2=0
cc_207 N_A_261_47#_c_334_n N_VGND_c_381_n 0.0144931f $X=3.4 $Y=0.39 $X2=0 $Y2=0
cc_208 N_A_261_47#_c_342_n N_VGND_c_381_n 0.0103304f $X=2.37 $Y=0.66 $X2=0 $Y2=0
