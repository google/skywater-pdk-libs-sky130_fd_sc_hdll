* File: sky130_fd_sc_hdll__xnor2_1.pex.spice
* Created: Wed Sep  2 08:53:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__XNOR2_1%B 1 3 4 6 7 9 10 12 13 16 17 19 22 27
c83 7 0 8.52358e-20 $X=2.395 $Y=1.41
c84 1 0 1.74411e-19 $X=0.535 $Y=1.41
r85 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r86 22 27 7.27582 $w=5.53e-07 $l=2.85e-07 $layer=LI1_cond $X=0.617 $Y=1.445
+ $X2=0.617 $Y2=1.16
r87 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.43
+ $Y=1.16 $X2=2.43 $Y2=1.16
r88 17 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.165 $Y=1.16
+ $X2=2.43 $Y2=1.16
r89 15 17 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.055 $Y=1.245
+ $X2=2.165 $Y2=1.16
r90 15 16 10.4768 $w=2.18e-07 $l=2e-07 $layer=LI1_cond $X=2.055 $Y=1.245
+ $X2=2.055 $Y2=1.445
r91 14 22 5.72073 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.81 $Y=1.53
+ $X2=0.617 $Y2=1.53
r92 13 16 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.945 $Y=1.53
+ $X2=2.055 $Y2=1.445
r93 13 14 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=1.945 $Y=1.53
+ $X2=0.81 $Y2=1.53
r94 10 20 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.54 $Y=0.995
+ $X2=2.455 $Y2=1.16
r95 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.54 $Y=0.995
+ $X2=2.54 $Y2=0.56
r96 7 20 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.455 $Y2=1.16
r97 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.985
r98 4 26 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.62 $Y=0.995
+ $X2=0.535 $Y2=1.16
r99 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.62 $Y=0.995 $X2=0.62
+ $Y2=0.56
r100 1 26 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=0.535 $Y=1.41
+ $X2=0.535 $Y2=1.16
r101 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.535 $Y=1.41
+ $X2=0.535 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_1%A 1 3 4 6 7 9 10 12 13 19 20 23
c49 20 0 2.59647e-19 $X=1.535 $Y=1.16
c50 10 0 1.73498e-19 $X=1.985 $Y=1.41
r51 19 21 60.5866 $w=3.58e-07 $l=4.5e-07 $layer=POLY_cond $X=1.535 $Y=1.202
+ $X2=1.985 $Y2=1.202
r52 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.535
+ $Y=1.16 $X2=1.535 $Y2=1.16
r53 17 19 4.71229 $w=3.58e-07 $l=3.5e-08 $layer=POLY_cond $X=1.5 $Y=1.202
+ $X2=1.535 $Y2=1.202
r54 16 17 66.6452 $w=3.58e-07 $l=4.95e-07 $layer=POLY_cond $X=1.005 $Y=1.202
+ $X2=1.5 $Y2=1.202
r55 15 16 3.36592 $w=3.58e-07 $l=2.5e-08 $layer=POLY_cond $X=0.98 $Y=1.202
+ $X2=1.005 $Y2=1.202
r56 13 20 19.6864 $w=1.98e-07 $l=3.55e-07 $layer=LI1_cond $X=1.18 $Y=1.175
+ $X2=1.535 $Y2=1.175
r57 13 23 1.66364 $w=1.98e-07 $l=3e-08 $layer=LI1_cond $X=1.18 $Y=1.175 $X2=1.15
+ $Y2=1.175
r58 10 21 18.8375 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.985 $Y=1.41
+ $X2=1.985 $Y2=1.202
r59 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.985 $Y=1.41
+ $X2=1.985 $Y2=1.985
r60 7 17 23.1716 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.5 $Y=0.995 $X2=1.5
+ $Y2=1.202
r61 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.5 $Y=0.995 $X2=1.5
+ $Y2=0.56
r62 4 16 18.8375 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.005 $Y=1.41
+ $X2=1.005 $Y2=1.202
r63 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.005 $Y=1.41
+ $X2=1.005 $Y2=1.985
r64 1 15 23.1716 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.98 $Y=0.995
+ $X2=0.98 $Y2=1.202
r65 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.98 $Y=0.995 $X2=0.98
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_1%A_47_47# 1 2 7 9 10 12 14 15 16 19 21 24
+ 25 26 29 33 36
c96 26 0 1.73498e-19 $X=2.555 $Y=1.5
r97 33 35 16.2536 $w=4.63e-07 $l=4.35e-07 $layer=LI1_cond $X=0.317 $Y=0.39
+ $X2=0.317 $Y2=0.825
r98 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.96
+ $Y=1.16 $X2=2.96 $Y2=1.16
r99 27 29 13.3579 $w=2.18e-07 $l=2.55e-07 $layer=LI1_cond $X=2.985 $Y=1.415
+ $X2=2.985 $Y2=1.16
r100 25 27 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.875 $Y=1.5
+ $X2=2.985 $Y2=1.415
r101 25 26 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.875 $Y=1.5
+ $X2=2.555 $Y2=1.5
r102 23 26 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.445 $Y=1.585
+ $X2=2.555 $Y2=1.5
r103 23 24 10.4768 $w=2.18e-07 $l=2e-07 $layer=LI1_cond $X=2.445 $Y=1.585
+ $X2=2.445 $Y2=1.785
r104 22 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.935 $Y=1.87
+ $X2=0.745 $Y2=1.87
r105 21 24 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.335 $Y=1.87
+ $X2=2.445 $Y2=1.785
r106 21 22 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=2.335 $Y=1.87
+ $X2=0.935 $Y2=1.87
r107 17 36 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=1.955
+ $X2=0.745 $Y2=1.87
r108 17 19 0.151637 $w=3.78e-07 $l=5e-09 $layer=LI1_cond $X=0.745 $Y=1.955
+ $X2=0.745 $Y2=1.96
r109 15 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.555 $Y=1.87
+ $X2=0.745 $Y2=1.87
r110 15 16 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.555 $Y=1.87
+ $X2=0.255 $Y2=1.87
r111 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=1.785
+ $X2=0.255 $Y2=1.87
r112 14 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.17 $Y=1.785
+ $X2=0.17 $Y2=0.825
r113 10 30 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=2.985 $Y2=1.16
r114 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=3.01 $Y2=0.56
r115 7 30 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.925 $Y=1.41
+ $X2=2.985 $Y2=1.16
r116 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.925 $Y=1.41
+ $X2=2.925 $Y2=1.985
r117 2 19 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.625
+ $Y=1.485 $X2=0.77 $Y2=1.96
r118 1 33 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.235
+ $Y=0.235 $X2=0.36 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_1%VPWR 1 2 3 10 12 14 16 18 25 39 42 45
r52 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r53 41 42 9.26921 $w=6.78e-07 $l=8.5e-08 $layer=LI1_cond $X=1.75 $Y=2.465
+ $X2=1.835 $Y2=2.465
r54 37 41 2.46251 $w=6.78e-07 $l=1.4e-07 $layer=LI1_cond $X=1.61 $Y=2.465
+ $X2=1.75 $Y2=2.465
r55 37 39 15.7773 $w=6.78e-07 $l=4.55e-07 $layer=LI1_cond $X=1.61 $Y=2.465
+ $X2=1.155 $Y2=2.465
r56 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r57 32 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r58 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r59 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r60 29 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r61 28 31 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r62 28 42 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=1.835 $Y2=2.72
r63 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r64 25 44 4.24846 $w=1.7e-07 $l=2.82e-07 $layer=LI1_cond $X=3.115 $Y=2.72
+ $X2=3.397 $Y2=2.72
r65 25 31 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.115 $Y=2.72
+ $X2=2.99 $Y2=2.72
r66 24 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r67 23 39 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=1.155 $Y2=2.72
r68 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r69 21 34 4.51997 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.192 $Y2=2.72
r70 21 23 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=1.15 $Y2=2.72
r71 18 24 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r72 18 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r73 14 44 3.26921 $w=3e-07 $l=1.69245e-07 $layer=LI1_cond $X=3.265 $Y=2.635
+ $X2=3.397 $Y2=2.72
r74 14 16 13.2531 $w=2.98e-07 $l=3.45e-07 $layer=LI1_cond $X=3.265 $Y=2.635
+ $X2=3.265 $Y2=2.29
r75 10 34 2.9977 $w=3e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.235 $Y=2.635
+ $X2=0.192 $Y2=2.72
r76 10 12 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.235 $Y=2.635
+ $X2=0.235 $Y2=2.34
r77 3 16 600 $w=1.7e-07 $l=8.92721e-07 $layer=licon1_PDIFF $count=1 $X=3.015
+ $Y=1.485 $X2=3.2 $Y2=2.29
r78 2 41 300 $w=1.7e-07 $l=1.08411e-06 $layer=licon1_PDIFF $count=2 $X=1.095
+ $Y=1.485 $X2=1.75 $Y2=2.29
r79 1 12 600 $w=1.7e-07 $l=9.33863e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.3 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_1%Y 1 2 8 10 14 16 20 22 25 27
r37 22 25 3.75819 $w=2e-07 $l=1.2e-07 $layer=LI1_cond $X=3.475 $Y=1.855
+ $X2=3.355 $Y2=1.855
r38 22 25 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=3.34 $Y=1.855
+ $X2=3.355 $Y2=1.855
r39 22 27 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=3.34 $Y=1.855 $X2=3.3
+ $Y2=1.855
r40 18 20 5.35743 $w=4.78e-07 $l=2.15e-07 $layer=LI1_cond $X=3.26 $Y=0.585
+ $X2=3.475 $Y2=0.585
r41 16 27 22.4591 $w=1.98e-07 $l=4.05e-07 $layer=LI1_cond $X=2.895 $Y=1.855
+ $X2=3.3 $Y2=1.855
r42 12 14 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.69 $Y=2.21
+ $X2=2.81 $Y2=2.21
r43 10 22 3.13183 $w=2.4e-07 $l=1e-07 $layer=LI1_cond $X=3.475 $Y=1.755
+ $X2=3.475 $Y2=1.855
r44 9 20 4.80115 $w=2.4e-07 $l=2.4e-07 $layer=LI1_cond $X=3.475 $Y=0.825
+ $X2=3.475 $Y2=0.585
r45 9 10 44.6572 $w=2.38e-07 $l=9.3e-07 $layer=LI1_cond $X=3.475 $Y=0.825
+ $X2=3.475 $Y2=1.755
r46 8 14 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=2.125
+ $X2=2.81 $Y2=2.21
r47 7 16 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.81 $Y=1.955
+ $X2=2.895 $Y2=1.855
r48 7 8 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.81 $Y=1.955 $X2=2.81
+ $Y2=2.125
r49 2 12 600 $w=1.7e-07 $l=8.21127e-07 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.485 $X2=2.69 $Y2=2.21
r50 1 18 182 $w=1.7e-07 $l=3.97995e-07 $layer=licon1_NDIFF $count=1 $X=3.085
+ $Y=0.235 $X2=3.26 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_1%VGND 1 2 9 12 13 14 15 21 37 38
r46 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r47 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r48 34 37 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r49 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r50 32 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r51 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r52 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r53 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r54 24 28 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r55 21 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r56 21 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r57 17 34 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.495 $Y=0 $X2=2.53
+ $Y2=0
r58 15 31 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.095 $Y=0 $X2=2.07
+ $Y2=0
r59 14 19 11.2363 $w=3.98e-07 $l=3.9e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.295
+ $Y2=0.39
r60 14 17 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.495
+ $Y2=0
r61 14 15 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.095
+ $Y2=0
r62 12 28 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.15
+ $Y2=0
r63 12 13 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.24
+ $Y2=0
r64 11 31 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=1.325 $Y=0 $X2=2.07
+ $Y2=0
r65 11 13 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.325 $Y=0 $X2=1.24
+ $Y2=0
r66 7 13 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.24 $Y=0.085 $X2=1.24
+ $Y2=0
r67 7 9 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.24 $Y=0.085
+ $X2=1.24 $Y2=0.39
r68 2 19 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.155
+ $Y=0.235 $X2=2.28 $Y2=0.39
r69 1 9 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.055
+ $Y=0.235 $X2=1.24 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_1%A_315_47# 1 2 9 11 12 13
r32 13 15 5.30435 $w=2.3e-07 $l=1e-07 $layer=LI1_cond $X=2.78 $Y=0.655 $X2=2.78
+ $Y2=0.555
r33 11 13 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.665 $Y=0.74
+ $X2=2.78 $Y2=0.655
r34 11 12 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=2.665 $Y=0.74
+ $X2=1.875 $Y2=0.74
r35 7 12 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=1.685 $Y=0.655
+ $X2=1.875 $Y2=0.74
r36 7 9 8.03677 $w=3.78e-07 $l=2.65e-07 $layer=LI1_cond $X=1.685 $Y=0.655
+ $X2=1.685 $Y2=0.39
r37 2 15 182 $w=1.7e-07 $l=3.81576e-07 $layer=licon1_NDIFF $count=1 $X=2.615
+ $Y=0.235 $X2=2.75 $Y2=0.555
r38 1 9 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.575
+ $Y=0.235 $X2=1.71 $Y2=0.39
.ends

