* File: sky130_fd_sc_hdll__a2bb2o_2.spice
* Created: Thu Aug 27 18:54:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a2bb2o_2.pex.spice"
.subckt sky130_fd_sc_hdll__a2bb2o_2  VNB VPB A1_N A2_N B2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_82_21#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.104 PD=1.83 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A_82_21#_M1011_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.178416 AS=0.104 PD=1.43972 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1006 N_A_343_47#_M1006_d N_A1_N_M1006_g N_VGND_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.115284 PD=0.74 PS=0.93028 NRD=0 NRS=59.988 M=1 R=2.8
+ SA=75001.3 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A2_N_M1005_g N_A_343_47#_M1006_d VNB NSHORT L=0.15
+ W=0.42 AD=0.15225 AS=0.0672 PD=1.145 PS=0.74 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75001.8 SB=75002 A=0.063 P=1.14 MULT=1
MM1013 N_A_82_21#_M1013_d N_A_343_47#_M1013_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.15225 PD=0.69 PS=1.145 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75002.7 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 A_696_47# N_B2_M1001_g N_A_82_21#_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0567 PD=0.74 PS=0.69 NRD=30 NRS=0 M=1 R=2.8 SA=75003.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_B1_M1012_g A_696_47# VNB NSHORT L=0.15 W=0.42 AD=0.1302
+ AS=0.0672 PD=1.46 PS=0.74 NRD=12.852 NRS=30 M=1 R=2.8 SA=75003.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_82_21#_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.275 PD=1.29 PS=2.55 NRD=0.9653 NRS=1.9503 M=1 R=5.55556
+ SA=90000.2 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1010 N_X_M1000_d N_A_82_21#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.236829 PD=1.29 PS=1.77439 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1008 A_341_297# N_A1_N_M1008_g N_VPWR_M1010_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0736 AS=0.151571 PD=0.87 PS=1.13561 NRD=18.4589 NRS=55.9677 M=1 R=3.55556
+ SA=90001.3 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1002 N_A_343_47#_M1002_d N_A2_N_M1002_g A_341_297# VPB PHIGHVT L=0.18 W=0.64
+ AD=0.176 AS=0.0736 PD=1.83 PS=0.87 NRD=1.5366 NRS=18.4589 M=1 R=3.55556
+ SA=90001.7 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1007 N_A_622_369#_M1007_d N_A_343_47#_M1007_g N_A_82_21#_M1007_s VPB PHIGHVT
+ L=0.18 W=0.64 AD=0.104 AS=0.1728 PD=0.965 PS=1.82 NRD=12.2928 NRS=1.5366 M=1
+ R=3.55556 SA=90000.2 SB=90001.2 A=0.1152 P=1.64 MULT=1
MM1009 N_VPWR_M1009_d N_B2_M1009_g N_A_622_369#_M1007_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.0928 AS=0.104 PD=0.93 PS=0.965 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.7 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1004 N_A_622_369#_M1004_d N_B1_M1004_g N_VPWR_M1009_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90001.2 SB=90000.2 A=0.1152 P=1.64 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
c_73 VPB 0 1.32963e-19 $X=0.125 $Y=2.635
*
.include "sky130_fd_sc_hdll__a2bb2o_2.pxi.spice"
*
.ends
*
*
