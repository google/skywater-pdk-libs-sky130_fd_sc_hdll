* File: sky130_fd_sc_hdll__ebufn_2.spice
* Created: Thu Aug 27 19:07:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__ebufn_2.pex.spice"
.subckt sky130_fd_sc_hdll__ebufn_2  VNB VPB A TE_B VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* TE_B	TE_B
* A	A
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_M1010_g N_A_27_47#_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.08925 AS=0.1092 PD=0.845 PS=1.36 NRD=12.852 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1002 N_A_224_47#_M1002_d N_TE_B_M1002_g N_VGND_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1302 AS=0.08925 PD=1.46 PS=0.845 NRD=12.852 NRS=28.56 M=1 R=2.8
+ SA=75000.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_224_47#_M1001_g N_A_412_47#_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.234 PD=0.92 PS=2.02 NRD=0 NRS=17.532 M=1 R=4.33333
+ SA=75000.3 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1001_d N_A_224_47#_M1004_g N_A_412_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.141375 PD=0.92 PS=1.085 NRD=0 NRS=18.456 M=1 R=4.33333
+ SA=75000.7 SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1005 N_A_412_47#_M1004_s N_A_27_47#_M1005_g N_Z_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.141375 AS=0.12025 PD=1.085 PS=1.02 NRD=10.152 NRS=8.304 M=1
+ R=4.33333 SA=75001.3 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1011 N_A_412_47#_M1011_d N_A_27_47#_M1011_g N_Z_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.8 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_27_47#_M1000_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.1264 AS=0.1728 PD=1.035 PS=1.82 NRD=18.4589 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.8 A=0.1152 P=1.64 MULT=1
MM1006 N_A_224_47#_M1006_d N_TE_B_M1006_g N_VPWR_M1000_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.1264 PD=1.82 PS=1.035 NRD=1.5366 NRS=16.9223 M=1
+ R=3.55556 SA=90000.8 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1007 N_A_340_309#_M1007_d N_TE_B_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.2538 AS=0.1363 PD=2.42 PS=1.23 NRD=1.0441 NRS=1.0441 M=1 R=5.22222
+ SA=90000.2 SB=90002.1 A=0.1692 P=2.24 MULT=1
MM1008 N_A_340_309#_M1008_d N_TE_B_M1008_g N_VPWR_M1007_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.392426 AS=0.1363 PD=1.75887 PS=1.23 NRD=13.6127 NRS=1.0441 M=1
+ R=5.22222 SA=90000.6 SB=90001.7 A=0.1692 P=2.24 MULT=1
MM1003 N_A_340_309#_M1008_d N_A_27_47#_M1003_g N_Z_M1003_s VPB PHIGHVT L=0.18
+ W=1 AD=0.417474 AS=0.145 PD=1.87113 PS=1.29 NRD=15.7403 NRS=0.9653 M=1
+ R=5.55556 SA=90001.6 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1009 N_A_340_309#_M1009_d N_A_27_47#_M1009_g N_Z_M1003_s VPB PHIGHVT L=0.18
+ W=1 AD=0.29 AS=0.145 PD=2.58 PS=1.29 NRD=4.9053 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.9929 P=13.17
pX13_noxref noxref_12 TE_B TE_B PROBETYPE=1
pX14_noxref noxref_13 Z Z PROBETYPE=1
pX15_noxref noxref_14 Z Z PROBETYPE=1
pX16_noxref noxref_15 Z Z PROBETYPE=1
*
.include "sky130_fd_sc_hdll__ebufn_2.pxi.spice"
*
.ends
*
*
