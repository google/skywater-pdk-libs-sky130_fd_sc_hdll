* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
X0 Y A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_485_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR a_1311_21# a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 a_109_47# a_1311_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_493_297# a_1311_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 a_485_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Y A0 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y A0 a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 a_493_297# A1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 a_117_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_485_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Y A1 a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_117_297# A0 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 Y A0 a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 Y A1 a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VPWR a_1311_21# a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 a_109_47# A0 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_493_297# a_1311_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 a_117_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 a_109_47# A0 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 Y A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 VPWR S a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 VGND S a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_109_47# a_1311_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VGND a_1311_21# a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_117_297# A0 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X26 Y A0 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VGND S a_1311_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VPWR S a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 VPWR S a_1311_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X30 VGND S a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 VGND a_1311_21# a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 a_493_297# A1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 a_485_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
