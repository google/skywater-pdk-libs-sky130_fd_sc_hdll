* NGSPICE file created from sky130_fd_sc_hdll__clkinv_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__clkinv_1 A VGND VNB VPB VPWR Y
M1000 VGND A Y VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.323e+11p ps=1.47e+06u
M1001 Y A VPWR VPB phighvt w=840000u l=180000u
+  ad=2.436e+11p pd=2.26e+06u as=4.704e+11p ps=4.48e+06u
M1002 VPWR A Y VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

