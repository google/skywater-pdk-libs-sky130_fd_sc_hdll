* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 VGND A1_N a_313_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND B1 a_627_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 a_723_369# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X6 VPWR a_321_369# a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X7 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VPWR A1_N a_321_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X9 a_84_21# B2 a_723_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X10 a_84_21# a_321_369# a_627_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_313_47# A2_N a_321_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_627_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_321_369# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
.ends
