* File: sky130_fd_sc_hdll__sdfstp_1.spice
* Created: Thu Aug 27 19:27:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__sdfstp_1.pex.spice"
.subckt sky130_fd_sc_hdll__sdfstp_1  VNB VPB SCD SCE D CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* SCE	SCE
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1022 A_119_47# N_SCD_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.42 AD=0.0546
+ AS=0.1302 PD=0.68 PS=1.46 NRD=21.42 NRS=12.852 M=1 R=2.8 SA=75000.2 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1030 N_A_201_47#_M1030_d N_SCE_M1030_g A_119_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0546 PD=0.74 PS=0.68 NRD=0 NRS=21.42 M=1 R=2.8 SA=75000.6
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1029 A_295_47# N_D_M1029_g N_A_201_47#_M1030_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0672 PD=0.69 PS=0.74 NRD=22.848 NRS=12.852 M=1 R=2.8 SA=75001.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_349_21#_M1001_g A_295_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1428 AS=0.0567 PD=1.52 PS=0.69 NRD=21.42 NRS=22.848 M=1 R=2.8 SA=75001.5
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_SCE_M1005_g N_A_349_21#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1302 PD=1.36 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_CLK_M1017_g N_A_693_369#_M1017_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1015 N_A_877_369#_M1015_d N_A_693_369#_M1015_g N_VGND_M1017_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1092 AS=0.0672 PD=1.36 PS=0.74 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1026 N_A_1075_413#_M1026_d N_A_693_369#_M1026_g N_A_201_47#_M1026_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1023 A_1177_47# N_A_877_369#_M1023_g N_A_1075_413#_M1026_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0546 AS=0.0672 PD=0.68 PS=0.74 NRD=21.42 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_1229_21#_M1016_g A_1177_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0546 PD=1.36 PS=0.68 NRD=0 NRS=21.42 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1020 A_1467_47# N_A_1075_413#_M1020_g N_A_1229_21#_M1020_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1512 PD=0.63 PS=1.56 NRD=14.28 NRS=27.132 M=1 R=2.8
+ SA=75000.3 SB=75004.2 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_SET_B_M1024_g A_1467_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0898245 AS=0.0441 PD=0.808302 PS=0.63 NRD=15.708 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75003.9 A=0.063 P=1.14 MULT=1
MM1018 A_1645_47# N_A_1075_413#_M1018_g N_VGND_M1024_d VNB NSHORT L=0.15 W=0.64
+ AD=0.2528 AS=0.136875 PD=1.43 PS=1.2317 NRD=63.744 NRS=8.436 M=1 R=4.26667
+ SA=75000.9 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1007 N_A_1725_329#_M1007_d N_A_877_369#_M1007_g A_1645_47# VNB NSHORT L=0.15
+ W=0.64 AD=0.149857 AS=0.2528 PD=1.3283 PS=1.43 NRD=0 NRS=63.744 M=1 R=4.26667
+ SA=75001.8 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1003 A_1955_47# N_A_693_369#_M1003_g N_A_1725_329#_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0983434 PD=0.63 PS=0.871698 NRD=14.28 NRS=52.848 M=1
+ R=2.8 SA=75002.7 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1027 A_2027_47# N_A_1921_295#_M1027_g A_1955_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.0441 PD=0.8 PS=0.63 NRD=38.568 NRS=14.28 M=1 R=2.8 SA=75003.1
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1031_d N_SET_B_M1031_g A_2027_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0924 AS=0.0798 PD=0.86 PS=0.8 NRD=32.856 NRS=38.568 M=1 R=2.8 SA=75003.6
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1034 N_A_1921_295#_M1034_d N_A_1725_329#_M1034_g N_VGND_M1031_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1596 AS=0.0924 PD=1.6 PS=0.86 NRD=32.856 NRS=12.852 M=1
+ R=2.8 SA=75004.2 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1032 N_VGND_M1032_d N_A_1725_329#_M1032_g N_A_2381_47#_M1032_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0971495 AS=0.1092 PD=0.843925 PS=1.36 NRD=19.992 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1002 N_Q_M1002_d N_A_2381_47#_M1002_g N_VGND_M1032_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.15035 PD=1.82 PS=1.30607 NRD=0 NRS=13.836 M=1 R=4.33333
+ SA=75000.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_VPWR_M1008_d N_SCD_M1008_g N_A_27_369#_M1008_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90001.5 A=0.1152 P=1.64 MULT=1
MM1033 A_211_369# N_SCE_M1033_g N_VPWR_M1008_d VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0736 AS=0.0928 PD=0.87 PS=0.93 NRD=18.4589 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90001.1 A=0.1152 P=1.64 MULT=1
MM1036 N_A_201_47#_M1036_d N_D_M1036_g A_211_369# VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.0736 PD=0.93 PS=0.87 NRD=1.5366 NRS=18.4589 M=1 R=3.55556
+ SA=90001.1 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1021 N_A_27_369#_M1021_d N_A_349_21#_M1021_g N_A_201_47#_M1036_d VPB PHIGHVT
+ L=0.18 W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1
+ R=3.55556 SA=90001.5 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1012 N_VPWR_M1012_d N_SCE_M1012_g N_A_349_21#_M1012_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.1728 PD=1.82 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1039 N_VPWR_M1039_d N_CLK_M1039_g N_A_693_369#_M1039_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1025 N_A_877_369#_M1025_d N_A_693_369#_M1025_g N_VPWR_M1039_d VPB PHIGHVT
+ L=0.18 W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1
+ R=3.55556 SA=90000.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1006 N_A_1075_413#_M1006_d N_A_877_369#_M1006_g N_A_201_47#_M1006_s VPB
+ PHIGHVT L=0.18 W=0.42 AD=0.0609 AS=0.1134 PD=0.71 PS=1.38 NRD=2.3443
+ NRS=2.3443 M=1 R=2.33333 SA=90000.2 SB=90005.2 A=0.0756 P=1.2 MULT=1
MM1037 A_1169_413# N_A_693_369#_M1037_g N_A_1075_413#_M1006_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0798 AS=0.0609 PD=0.8 PS=0.71 NRD=63.3158 NRS=2.3443 M=1 R=2.33333
+ SA=90000.6 SB=90004.7 A=0.0756 P=1.2 MULT=1
MM1038 N_VPWR_M1038_d N_A_1229_21#_M1038_g A_1169_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.1071 AS=0.0798 PD=0.93 PS=0.8 NRD=30.4759 NRS=63.3158 M=1 R=2.33333
+ SA=90001.2 SB=90004.1 A=0.0756 P=1.2 MULT=1
MM1009 N_A_1229_21#_M1009_d N_A_1075_413#_M1009_g N_VPWR_M1038_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.0861 AS=0.1071 PD=0.83 PS=0.93 NRD=14.0658 NRS=77.3816 M=1
+ R=2.33333 SA=90001.9 SB=90003.4 A=0.0756 P=1.2 MULT=1
MM1000 N_VPWR_M1000_d N_SET_B_M1000_g N_A_1229_21#_M1009_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0854 AS=0.0861 PD=0.793333 PS=0.83 NRD=23.443 NRS=46.886 M=1
+ R=2.33333 SA=90002.5 SB=90002.8 A=0.0756 P=1.2 MULT=1
MM1028 A_1643_329# N_A_1075_413#_M1028_g N_VPWR_M1000_d VPB PHIGHVT L=0.18
+ W=0.84 AD=0.0966 AS=0.1708 PD=1.07 PS=1.58667 NRD=14.0658 NRS=4.6886 M=1
+ R=4.66667 SA=90001.6 SB=90001.4 A=0.1512 P=2.04 MULT=1
MM1013 N_A_1725_329#_M1013_d N_A_693_369#_M1013_g A_1643_329# VPB PHIGHVT L=0.18
+ W=0.84 AD=0.1848 AS=0.0966 PD=1.65333 PS=1.07 NRD=26.9693 NRS=14.0658 M=1
+ R=4.66667 SA=90002 SB=90001 A=0.1512 P=2.04 MULT=1
MM1010 A_1841_413# N_A_877_369#_M1010_g N_A_1725_329#_M1013_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0861 AS=0.0924 PD=0.83 PS=0.826667 NRD=70.3487 NRS=2.3443 M=1
+ R=2.33333 SA=90004 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1019 N_VPWR_M1019_d N_A_1921_295#_M1019_g A_1841_413# VPB PHIGHVT L=0.18
+ W=0.42 AD=0.07875 AS=0.0861 PD=0.795 PS=0.83 NRD=42.1974 NRS=70.3487 M=1
+ R=2.33333 SA=90004.6 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1011 N_A_1725_329#_M1011_d N_SET_B_M1011_g N_VPWR_M1019_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.07875 PD=1.38 PS=0.795 NRD=2.3443 NRS=2.3443 M=1
+ R=2.33333 SA=90005.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1014 N_A_1921_295#_M1014_d N_A_1725_329#_M1014_g N_VPWR_M1014_s VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.1134 AS=0.1134 PD=1.38 PS=1.38 NRD=2.3443 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1004 N_VPWR_M1004_d N_A_1725_329#_M1004_g N_A_2381_47#_M1004_s VPB PHIGHVT
+ L=0.18 W=0.64 AD=0.122693 AS=0.1728 PD=1.04976 PS=1.82 NRD=9.2196 NRS=1.5366
+ M=1 R=3.55556 SA=90000.2 SB=90000.7 A=0.1152 P=1.64 MULT=1
MM1035 N_Q_M1035_d N_A_2381_47#_M1035_g N_VPWR_M1004_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.191707 PD=2.54 PS=1.64024 NRD=0.9653 NRS=6.8753 M=1 R=5.55556
+ SA=90000.5 SB=90000.2 A=0.18 P=2.36 MULT=1
DX40_noxref VNB VPB NWDIODE A=22.0206 P=30.65
c_124 VNB 0 1.07953e-19 $X=0.145 $Y=-0.085
c_262 VPB 0 1.96862e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__sdfstp_1.pxi.spice"
*
.ends
*
*
