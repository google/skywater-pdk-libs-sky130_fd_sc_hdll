* File: sky130_fd_sc_hdll__sedfxbp_2.pex.spice
* Created: Thu Aug 27 19:28:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%CLK 1 2 3 5 6 8 13
c37 1 0 2.71124e-20 $X=0.31 $Y=1.325
r38 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r39 6 16 86.4067 $w=2.69e-07 $l=5.05816e-07 $layer=POLY_cond $X=0.52 $Y=0.73
+ $X2=0.355 $Y2=1.16
r40 6 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.445
r41 3 9 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=0.495 $Y=1.665
+ $X2=0.31 $Y2=1.665
r42 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.74
+ $X2=0.495 $Y2=2.135
r43 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.31 $Y=1.59 $X2=0.31
+ $Y2=1.665
r44 1 16 38.9235 $w=2.69e-07 $l=1.86145e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.355 $Y2=1.16
r45 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.31 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_27_47# 1 2 8 9 11 14 18 20 22 24 25 27
+ 28 32 36 40 41 42 45 47 49 52 55 57 58 59 60 61 68 70 76 84 88
c281 68 0 2.41332e-19 $X=8.43 $Y=1.87
c282 60 0 1.92092e-19 $X=11.075 $Y=1.87
c283 58 0 1.69416e-19 $X=8.285 $Y=1.87
c284 52 0 1.6051e-19 $X=8.065 $Y=0.87
c285 49 0 1.43548e-19 $X=8.285 $Y=0.845
c286 45 0 1.77499e-19 $X=0.78 $Y=1.795
c287 42 0 1.03679e-19 $X=0.665 $Y=1.88
r288 87 89 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=11.235 $Y=1.41
+ $X2=11.235 $Y2=1.575
r289 87 88 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.21
+ $Y=1.41 $X2=11.21 $Y2=1.41
r290 84 87 16.2293 $w=3.2e-07 $l=9e-08 $layer=POLY_cond $X=11.235 $Y=1.32
+ $X2=11.235 $Y2=1.41
r291 75 76 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.235
+ $X2=0.99 $Y2=1.235
r292 71 88 22.0885 $w=2.38e-07 $l=4.6e-07 $layer=LI1_cond $X=11.245 $Y=1.87
+ $X2=11.245 $Y2=1.41
r293 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.245 $Y=1.87
+ $X2=11.245 $Y2=1.87
r294 68 95 1.97562 $w=3.48e-07 $l=6e-08 $layer=LI1_cond $X=8.43 $Y=1.83 $X2=8.37
+ $Y2=1.83
r295 68 82 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.54
+ $Y=1.74 $X2=8.54 $Y2=1.74
r296 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.43 $Y=1.87
+ $X2=8.43 $Y2=1.87
r297 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.77 $Y=1.87
+ $X2=0.77 $Y2=1.87
r298 61 67 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=8.625 $Y=1.87
+ $X2=8.43 $Y2=1.87
r299 60 70 0.131507 $w=2.3e-07 $l=1.7e-07 $layer=MET1_cond $X=11.075 $Y=1.87
+ $X2=11.245 $Y2=1.87
r300 60 61 3.03217 $w=1.4e-07 $l=2.45e-06 $layer=MET1_cond $X=11.075 $Y=1.87
+ $X2=8.625 $Y2=1.87
r301 59 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.915 $Y=1.87
+ $X2=0.77 $Y2=1.87
r302 58 67 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.285 $Y=1.87
+ $X2=8.43 $Y2=1.87
r303 58 59 9.12127 $w=1.4e-07 $l=7.37e-06 $layer=MET1_cond $X=8.285 $Y=1.87
+ $X2=0.915 $Y2=1.87
r304 55 95 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=8.37 $Y=1.655
+ $X2=8.37 $Y2=1.83
r305 54 55 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=8.37 $Y=0.955
+ $X2=8.37 $Y2=1.655
r306 52 79 40.861 $w=3.8e-07 $l=1.35e-07 $layer=POLY_cond $X=8.09 $Y=0.87
+ $X2=8.09 $Y2=0.735
r307 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.065
+ $Y=0.87 $X2=8.065 $Y2=0.87
r308 49 54 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=8.285 $Y=0.845
+ $X2=8.37 $Y2=0.955
r309 49 51 11.5244 $w=2.18e-07 $l=2.2e-07 $layer=LI1_cond $X=8.285 $Y=0.845
+ $X2=8.065 $Y2=0.845
r310 48 75 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=0.81 $Y=1.235
+ $X2=0.965 $Y2=1.235
r311 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.81
+ $Y=1.235 $X2=0.81 $Y2=1.235
r312 45 64 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=1.795
+ $X2=0.78 $Y2=1.88
r313 45 47 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.78 $Y=1.795
+ $X2=0.78 $Y2=1.235
r314 44 47 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=0.805
+ $X2=0.78 $Y2=1.235
r315 43 57 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r316 42 64 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.665 $Y=1.88
+ $X2=0.78 $Y2=1.88
r317 42 43 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.665 $Y=1.88
+ $X2=0.345 $Y2=1.88
r318 40 44 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.665 $Y=0.72
+ $X2=0.78 $Y2=0.805
r319 40 41 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.665 $Y=0.72
+ $X2=0.345 $Y2=0.72
r320 34 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r321 34 36 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r322 30 32 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=11.995 $Y=1.245
+ $X2=11.995 $Y2=0.415
r323 29 84 20.4921 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=11.395 $Y=1.32
+ $X2=11.235 $Y2=1.32
r324 28 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.92 $Y=1.32
+ $X2=11.995 $Y2=1.245
r325 28 29 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=11.92 $Y=1.32
+ $X2=11.395 $Y2=1.32
r326 25 27 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=11.24 $Y=1.99
+ $X2=11.24 $Y2=2.275
r327 24 25 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=11.24 $Y=1.89 $X2=11.24
+ $Y2=1.99
r328 24 89 104.447 $w=2e-07 $l=3.15e-07 $layer=POLY_cond $X=11.24 $Y=1.89
+ $X2=11.24 $Y2=1.575
r329 20 82 46.6797 $w=3.23e-07 $l=2.8592e-07 $layer=POLY_cond $X=8.47 $Y=1.99
+ $X2=8.547 $Y2=1.74
r330 20 22 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=8.47 $Y=1.99
+ $X2=8.47 $Y2=2.275
r331 18 79 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.075 $Y=0.415
+ $X2=8.075 $Y2=0.735
r332 12 76 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=1.235
r333 12 14 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=0.445
r334 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.965 $Y=1.74
+ $X2=0.965 $Y2=2.135
r335 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.64 $X2=0.965
+ $Y2=1.74
r336 7 75 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=0.965 $Y=1.37
+ $X2=0.965 $Y2=1.235
r337 7 8 89.5258 $w=2e-07 $l=2.7e-07 $layer=POLY_cond $X=0.965 $Y=1.37 $X2=0.965
+ $Y2=1.64
r338 2 57 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r339 1 36 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%D 2 3 5 8 10 13
r47 13 15 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=1.145
+ $X2=1.89 $Y2=0.98
r48 13 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.88
+ $Y=1.145 $X2=1.88 $Y2=1.145
r49 10 14 2.2356 $w=9.53e-07 $l=1.75e-07 $layer=LI1_cond $X=2.055 $Y=1.242
+ $X2=1.88 $Y2=1.242
r50 8 15 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=1.99 $Y=0.445
+ $X2=1.99 $Y2=0.98
r51 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.955 $Y=1.77
+ $X2=1.955 $Y2=2.165
r52 2 3 49.3715 $w=2.88e-07 $l=3.25883e-07 $layer=POLY_cond $X=1.89 $Y=1.475
+ $X2=1.955 $Y2=1.77
r53 1 13 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=1.89 $Y=1.155 $X2=1.89
+ $Y2=1.145
r54 1 2 52.7581 $w=3.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.89 $Y=1.155 $X2=1.89
+ $Y2=1.475
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_455_324# 1 2 7 9 10 11 14 18 22 25 28
+ 29 33 38
c98 22 0 1.13207e-19 $X=3.12 $Y=0.51
r99 33 41 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.78 $Y=1.52
+ $X2=2.78 $Y2=1.695
r100 32 35 10.7351 $w=3.63e-07 $l=3.4e-07 $layer=LI1_cond $X=2.78 $Y=1.537
+ $X2=3.12 $Y2=1.537
r101 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.78
+ $Y=1.52 $X2=2.78 $Y2=1.52
r102 29 44 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=1.01
+ $X2=3.825 $Y2=0.845
r103 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.8
+ $Y=1.01 $X2=3.8 $Y2=1.01
r104 26 38 0.565906 $w=3.3e-07 $l=1.53e-07 $layer=LI1_cond $X=3.285 $Y=1.01
+ $X2=3.132 $Y2=1.01
r105 26 28 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=3.285 $Y=1.01
+ $X2=3.8 $Y2=1.01
r106 25 35 0.378885 $w=3.63e-07 $l=1.2e-08 $layer=LI1_cond $X=3.132 $Y=1.537
+ $X2=3.12 $Y2=1.537
r107 24 38 6.17543 $w=2.65e-07 $l=1.65e-07 $layer=LI1_cond $X=3.132 $Y=1.175
+ $X2=3.132 $Y2=1.01
r108 24 25 6.8013 $w=3.03e-07 $l=1.8e-07 $layer=LI1_cond $X=3.132 $Y=1.175
+ $X2=3.132 $Y2=1.355
r109 20 38 6.17543 $w=2.65e-07 $l=1.83916e-07 $layer=LI1_cond $X=3.092 $Y=0.845
+ $X2=3.132 $Y2=1.01
r110 20 22 17.1586 $w=2.23e-07 $l=3.35e-07 $layer=LI1_cond $X=3.092 $Y=0.845
+ $X2=3.092 $Y2=0.51
r111 16 35 1.32393 $w=3.3e-07 $l=1.83e-07 $layer=LI1_cond $X=3.12 $Y=1.72
+ $X2=3.12 $Y2=1.537
r112 16 18 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=3.12 $Y=1.72
+ $X2=3.12 $Y2=1.99
r113 14 44 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.82 $Y=0.445
+ $X2=3.82 $Y2=0.845
r114 10 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.615 $Y=1.695
+ $X2=2.78 $Y2=1.695
r115 10 11 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.615 $Y=1.695
+ $X2=2.455 $Y2=1.695
r116 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.365 $Y=1.77
+ $X2=2.455 $Y2=1.695
r117 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.365 $Y=1.77
+ $X2=2.365 $Y2=2.165
r118 2 18 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.995
+ $Y=1.845 $X2=3.12 $Y2=1.99
r119 1 22 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=2.995
+ $Y=0.235 $X2=3.12 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%DE 3 5 8 9 11 14 16 18 20 21 22 23 25 32
+ 35
c90 32 0 1.13207e-19 $X=2.655 $Y=0.992
r91 30 32 54.5718 $w=3.65e-07 $l=2.15e-07 $layer=POLY_cond $X=2.44 $Y=0.992
+ $X2=2.655 $Y2=0.992
r92 30 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.44
+ $Y=1.01 $X2=2.44 $Y2=1.01
r93 25 35 3.33333 $w=3.66e-07 $l=1e-07 $layer=LI1_cond $X=2.545 $Y=0.85
+ $X2=2.545 $Y2=0.95
r94 18 23 78.7283 $w=2e-07 $l=2.35e-07 $layer=POLY_cond $X=3.845 $Y=1.77
+ $X2=3.845 $Y2=1.535
r95 18 20 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.845 $Y=1.77
+ $X2=3.845 $Y2=2.165
r96 17 22 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=3.455 $Y=1.535
+ $X2=3.355 $Y2=1.535
r97 16 23 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=3.745 $Y=1.535
+ $X2=3.845 $Y2=1.535
r98 16 17 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.745 $Y=1.535
+ $X2=3.455 $Y2=1.535
r99 12 21 17.9196 $w=1.75e-07 $l=8.66025e-08 $layer=POLY_cond $X=3.38 $Y=0.85
+ $X2=3.355 $Y2=0.925
r100 12 14 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=3.38 $Y=0.85
+ $X2=3.38 $Y2=0.445
r101 9 22 78.7283 $w=2e-07 $l=2.35e-07 $layer=POLY_cond $X=3.355 $Y=1.77
+ $X2=3.355 $Y2=1.535
r102 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.355 $Y=1.77
+ $X2=3.355 $Y2=2.165
r103 8 22 24.8683 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=3.355 $Y=1.46
+ $X2=3.355 $Y2=1.535
r104 7 21 17.9196 $w=1.75e-07 $l=7.5e-08 $layer=POLY_cond $X=3.355 $Y=1
+ $X2=3.355 $Y2=0.925
r105 7 8 152.525 $w=2e-07 $l=4.6e-07 $layer=POLY_cond $X=3.355 $Y=1 $X2=3.355
+ $Y2=1.46
r106 5 21 7.5188 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=3.255 $Y=0.925
+ $X2=3.355 $Y2=0.925
r107 5 32 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.255 $Y=0.925
+ $X2=2.655 $Y2=0.925
r108 1 30 14.2284 $w=3.65e-07 $l=9e-08 $layer=POLY_cond $X=2.35 $Y=0.992
+ $X2=2.44 $Y2=0.992
r109 1 3 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.35 $Y=0.81 $X2=2.35
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_851_264# 1 2 7 9 12 15 16 18 21 23 25
+ 27 30 32 34 36 39 41 43 48 54 59 61 64 65 68 71 82
c232 64 0 6.12178e-20 $X=14.385 $Y=0.85
c233 59 0 8.50484e-20 $X=14.155 $Y=1.055
c234 16 0 1.42198e-20 $X=12.38 $Y=1.99
c235 12 0 5.64525e-20 $X=4.43 $Y=0.445
r236 72 82 15.7614 $w=3.38e-07 $l=4.65e-07 $layer=LI1_cond $X=14.525 $Y=0.85
+ $X2=14.525 $Y2=0.385
r237 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.53 $Y=0.85
+ $X2=14.53 $Y2=0.85
r238 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.19 $Y=0.85
+ $X2=4.19 $Y2=0.85
r239 65 67 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.335 $Y=0.85
+ $X2=4.19 $Y2=0.85
r240 64 71 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.385 $Y=0.85
+ $X2=14.53 $Y2=0.85
r241 64 65 12.4381 $w=1.4e-07 $l=1.005e-05 $layer=MET1_cond $X=14.385 $Y=0.85
+ $X2=4.335 $Y2=0.85
r242 62 72 1.35582 $w=3.38e-07 $l=4e-08 $layer=LI1_cond $X=14.525 $Y=0.89
+ $X2=14.525 $Y2=0.85
r243 61 62 0.533618 $w=3.4e-07 $l=1.65e-07 $layer=LI1_cond $X=14.525 $Y=1.055
+ $X2=14.525 $Y2=0.89
r244 59 77 15.9965 $w=2.7e-07 $l=7.2e-08 $layer=POLY_cond $X=14.155 $Y=1.055
+ $X2=14.155 $Y2=1.127
r245 58 61 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=14.155 $Y=1.055
+ $X2=14.525 $Y2=1.055
r246 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.155
+ $Y=1.055 $X2=14.155 $Y2=1.055
r247 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.39
+ $Y=1.485 $X2=4.39 $Y2=1.485
r248 51 68 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=4.19 $Y=1.32
+ $X2=4.19 $Y2=0.85
r249 50 54 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=4.19 $Y=1.485 $X2=4.39
+ $Y2=1.485
r250 50 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.19 $Y=1.485
+ $X2=4.19 $Y2=1.32
r251 46 61 0.533618 $w=3.4e-07 $l=1.65e-07 $layer=LI1_cond $X=14.525 $Y=1.22
+ $X2=14.525 $Y2=1.055
r252 46 48 26.0994 $w=3.38e-07 $l=7.7e-07 $layer=LI1_cond $X=14.525 $Y=1.22
+ $X2=14.525 $Y2=1.99
r253 42 45 8.26431 $w=1.85e-07 $l=1.33e-07 $layer=POLY_cond $X=13.55 $Y=1.127
+ $X2=13.417 $Y2=1.127
r254 41 77 11.7477 $w=1.85e-07 $l=1.35e-07 $layer=POLY_cond $X=14.02 $Y=1.127
+ $X2=14.155 $Y2=1.127
r255 41 42 173.629 $w=1.85e-07 $l=4.7e-07 $layer=POLY_cond $X=14.02 $Y=1.127
+ $X2=13.55 $Y2=1.127
r256 37 45 25.1228 $w=2.32e-07 $l=1.17473e-07 $layer=POLY_cond $X=13.475
+ $Y=1.035 $X2=13.417 $Y2=1.127
r257 37 39 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=13.475 $Y=1.035
+ $X2=13.475 $Y2=0.56
r258 34 45 61.3446 $w=2.32e-07 $l=2.98572e-07 $layer=POLY_cond $X=13.385 $Y=1.41
+ $X2=13.417 $Y2=1.127
r259 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=13.385 $Y=1.41
+ $X2=13.385 $Y2=1.985
r260 33 44 8.26431 $w=1.85e-07 $l=1.33e-07 $layer=POLY_cond $X=13.08 $Y=1.127
+ $X2=12.947 $Y2=1.127
r261 32 45 8.26431 $w=1.85e-07 $l=1.32e-07 $layer=POLY_cond $X=13.285 $Y=1.127
+ $X2=13.417 $Y2=1.127
r262 32 33 75.7318 $w=1.85e-07 $l=2.05e-07 $layer=POLY_cond $X=13.285 $Y=1.127
+ $X2=13.08 $Y2=1.127
r263 28 44 25.1228 $w=2.32e-07 $l=1.17473e-07 $layer=POLY_cond $X=13.005
+ $Y=1.035 $X2=12.947 $Y2=1.127
r264 28 30 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=13.005 $Y=1.035
+ $X2=13.005 $Y2=0.56
r265 25 44 61.3446 $w=2.32e-07 $l=2.98572e-07 $layer=POLY_cond $X=12.915 $Y=1.41
+ $X2=12.947 $Y2=1.127
r266 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.915 $Y=1.41
+ $X2=12.915 $Y2=1.985
r267 24 43 4.51672 $w=1.85e-07 $l=1.33e-07 $layer=POLY_cond $X=12.545 $Y=1.127
+ $X2=12.412 $Y2=1.127
r268 23 44 8.26431 $w=1.85e-07 $l=1.32e-07 $layer=POLY_cond $X=12.815 $Y=1.127
+ $X2=12.947 $Y2=1.127
r269 23 24 99.7443 $w=1.85e-07 $l=2.7e-07 $layer=POLY_cond $X=12.815 $Y=1.127
+ $X2=12.545 $Y2=1.127
r270 19 43 21.3708 $w=1.75e-07 $l=1.17473e-07 $layer=POLY_cond $X=12.47 $Y=1.035
+ $X2=12.412 $Y2=1.127
r271 19 21 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=12.47 $Y=1.035
+ $X2=12.47 $Y2=0.445
r272 16 18 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=12.38 $Y=1.99
+ $X2=12.38 $Y2=2.275
r273 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=12.38 $Y=1.89 $X2=12.38
+ $Y2=1.99
r274 14 43 21.3708 $w=1.75e-07 $l=1.07819e-07 $layer=POLY_cond $X=12.38 $Y=1.22
+ $X2=12.412 $Y2=1.127
r275 14 15 222.157 $w=2e-07 $l=6.7e-07 $layer=POLY_cond $X=12.38 $Y=1.22
+ $X2=12.38 $Y2=1.89
r276 10 55 38.6342 $w=2.88e-07 $l=1.72337e-07 $layer=POLY_cond $X=4.43 $Y=1.32
+ $X2=4.415 $Y2=1.485
r277 10 12 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=4.43 $Y=1.32
+ $X2=4.43 $Y2=0.445
r278 7 55 54.4391 $w=2.88e-07 $l=2.89957e-07 $layer=POLY_cond $X=4.405 $Y=1.77
+ $X2=4.415 $Y2=1.485
r279 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=4.405 $Y=1.77
+ $X2=4.405 $Y2=2.165
r280 2 48 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=14.395
+ $Y=1.845 $X2=14.52 $Y2=1.99
r281 1 82 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=14.405
+ $Y=0.235 $X2=14.53 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_955_21# 1 2 7 9 10 11 13 14 16 17 20
+ 26 28 29 33 37 38
c118 28 0 1.97212e-19 $X=6.14 $Y=1.835
c119 20 0 1.41479e-20 $X=5.765 $Y=0.34
c120 14 0 4.70699e-20 $X=7.32 $Y=1.77
r121 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.235
+ $Y=1.52 $X2=7.235 $Y2=1.52
r122 31 33 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=7.245 $Y=1.835
+ $X2=7.245 $Y2=1.52
r123 30 37 2.83584 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=6.225 $Y=1.92
+ $X2=6.007 $Y2=1.92
r124 29 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.12 $Y=1.92
+ $X2=7.245 $Y2=1.835
r125 29 30 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=7.12 $Y=1.92
+ $X2=6.225 $Y2=1.92
r126 28 37 3.64284 $w=2.55e-07 $l=1.70276e-07 $layer=LI1_cond $X=6.14 $Y=1.835
+ $X2=6.007 $Y2=1.92
r127 28 38 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=6.14 $Y=1.835
+ $X2=6.14 $Y2=0.935
r128 24 38 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.06 $Y=0.77
+ $X2=6.06 $Y2=0.935
r129 24 26 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=6.06 $Y=0.77 $X2=6.06
+ $Y2=0.75
r130 23 26 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=6.06 $Y=0.515
+ $X2=6.06 $Y2=0.75
r131 20 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.765 $Y=0.34
+ $X2=5.765 $Y2=0.505
r132 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.765
+ $Y=0.34 $X2=5.765 $Y2=0.34
r133 17 23 6.94204 $w=2.6e-07 $l=2.20624e-07 $layer=LI1_cond $X=5.895 $Y=0.385
+ $X2=6.06 $Y2=0.515
r134 17 19 6.1 $w=2.6e-07 $l=1.3e-07 $layer=LI1_cond $X=5.895 $Y=0.385 $X2=5.765
+ $Y2=0.385
r135 14 34 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=7.32 $Y=1.77
+ $X2=7.26 $Y2=1.52
r136 14 16 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=7.32 $Y=1.77
+ $X2=7.32 $Y2=2.165
r137 13 41 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=5.705 $Y=0.765
+ $X2=5.705 $Y2=0.505
r138 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.63 $Y=0.84
+ $X2=5.705 $Y2=0.765
r139 10 11 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=5.63 $Y=0.84
+ $X2=4.925 $Y2=0.84
r140 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.85 $Y=0.765
+ $X2=4.925 $Y2=0.84
r141 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.85 $Y=0.765
+ $X2=4.85 $Y2=0.445
r142 2 37 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=5.83
+ $Y=1.845 $X2=5.955 $Y2=2
r143 1 26 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=5.935
+ $Y=0.595 $X2=6.06 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%SCD 1 3 6 8
c40 6 0 3.43252e-19 $X=6.79 $Y=0.805
r41 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.705
+ $Y=1.52 $X2=6.705 $Y2=1.52
r42 8 12 7.81596 $w=5.03e-07 $l=3.3e-07 $layer=LI1_cond $X=6.697 $Y=1.19
+ $X2=6.697 $Y2=1.52
r43 4 11 38.578 $w=2.95e-07 $l=1.92678e-07 $layer=POLY_cond $X=6.79 $Y=1.355
+ $X2=6.73 $Y2=1.52
r44 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.79 $Y=1.355 $X2=6.79
+ $Y2=0.805
r45 1 11 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=6.79 $Y=1.77
+ $X2=6.73 $Y2=1.52
r46 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=6.79 $Y=1.77 $X2=6.79
+ $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%SCE 1 3 4 6 8 12 13 14 17 19 21 26 31
c92 19 0 1.69416e-19 $X=4.915 $Y=1.5
r93 26 27 9.85014 $w=3.67e-07 $l=7.5e-08 $layer=POLY_cond $X=6.195 $Y=1.43
+ $X2=6.27 $Y2=1.43
r94 24 26 57.7875 $w=3.67e-07 $l=4.4e-07 $layer=POLY_cond $X=5.755 $Y=1.43
+ $X2=6.195 $Y2=1.43
r95 21 31 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=5.745 $Y=1.44
+ $X2=5.745 $Y2=1.53
r96 21 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.755
+ $Y=1.44 $X2=5.755 $Y2=1.44
r97 15 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.15 $Y=0.255
+ $X2=7.15 $Y2=0.805
r98 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.075 $Y=0.18
+ $X2=7.15 $Y2=0.255
r99 13 14 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=7.075 $Y=0.18
+ $X2=6.345 $Y2=0.18
r100 10 27 23.77 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=6.27 $Y=1.09 $X2=6.27
+ $Y2=1.43
r101 10 12 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.27 $Y=1.09
+ $X2=6.27 $Y2=0.805
r102 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.27 $Y=0.255
+ $X2=6.345 $Y2=0.18
r103 9 12 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.27 $Y=0.255
+ $X2=6.27 $Y2=0.805
r104 6 26 19.4219 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=6.195 $Y=1.77
+ $X2=6.195 $Y2=1.43
r105 6 8 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=6.195 $Y=1.77
+ $X2=6.195 $Y2=2.165
r106 5 19 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=5.015 $Y=1.5 $X2=4.915
+ $Y2=1.5
r107 4 24 41.637 $w=3.67e-07 $l=2.17198e-07 $layer=POLY_cond $X=5.57 $Y=1.5
+ $X2=5.755 $Y2=1.43
r108 4 5 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=5.57 $Y=1.5
+ $X2=5.015 $Y2=1.5
r109 1 19 90.3335 $w=2e-07 $l=2.7e-07 $layer=POLY_cond $X=4.915 $Y=1.77
+ $X2=4.915 $Y2=1.5
r110 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=4.915 $Y=1.77
+ $X2=4.915 $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_211_363# 1 2 8 9 11 12 16 18 20 21 23
+ 26 27 30 31 32 33 42 43 47 49 58
c214 43 0 1.42198e-20 $X=11.715 $Y=1.53
c215 33 0 1.29874e-19 $X=8.165 $Y=1.53
c216 32 0 3.06364e-20 $X=11.545 $Y=1.53
c217 30 0 1.87807e-19 $X=7.825 $Y=1.53
c218 27 0 1.51095e-20 $X=11.475 $Y=0.87
c219 12 0 1.43548e-19 $X=8.54 $Y=1.29
c220 9 0 1.36878e-19 $X=7.965 $Y=1.99
r221 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.77
+ $Y=1.74 $X2=11.77 $Y2=1.74
r222 46 49 59.5246 $w=2.7e-07 $l=2.15e-07 $layer=POLY_cond $X=7.965 $Y=1.35
+ $X2=8.18 $Y2=1.35
r223 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.965
+ $Y=1.35 $X2=7.965 $Y2=1.35
r224 43 56 6.54089 $w=3.68e-07 $l=2.1e-07 $layer=LI1_cond $X=11.72 $Y=1.53
+ $X2=11.72 $Y2=1.74
r225 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.715 $Y=1.53
+ $X2=11.715 $Y2=1.53
r226 40 47 8.82722 $w=2.33e-07 $l=1.8e-07 $layer=LI1_cond $X=7.997 $Y=1.53
+ $X2=7.997 $Y2=1.35
r227 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.995 $Y=1.53
+ $X2=7.995 $Y2=1.53
r228 36 62 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.2 $Y=1.53 $X2=1.2
+ $Y2=1.96
r229 36 58 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.2 $Y=1.53
+ $X2=1.2 $Y2=0.51
r230 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=1.53 $X2=1.2
+ $Y2=1.53
r231 33 39 0.131507 $w=2.3e-07 $l=1.7e-07 $layer=MET1_cond $X=8.165 $Y=1.53
+ $X2=7.995 $Y2=1.53
r232 32 42 0.131507 $w=2.3e-07 $l=1.7e-07 $layer=MET1_cond $X=11.545 $Y=1.53
+ $X2=11.715 $Y2=1.53
r233 32 33 4.18316 $w=1.4e-07 $l=3.38e-06 $layer=MET1_cond $X=11.545 $Y=1.53
+ $X2=8.165 $Y2=1.53
r234 31 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=1.53
+ $X2=1.2 $Y2=1.53
r235 30 39 0.131507 $w=2.3e-07 $l=1.7e-07 $layer=MET1_cond $X=7.825 $Y=1.53
+ $X2=7.995 $Y2=1.53
r236 30 31 8.01979 $w=1.4e-07 $l=6.48e-06 $layer=MET1_cond $X=7.825 $Y=1.53
+ $X2=1.345 $Y2=1.53
r237 29 43 15.4178 $w=3.68e-07 $l=4.95e-07 $layer=LI1_cond $X=11.72 $Y=1.035
+ $X2=11.72 $Y2=1.53
r238 27 50 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=11.475 $Y=0.87
+ $X2=11.315 $Y2=0.87
r239 26 29 4.79917 $w=5.13e-07 $l=1.65e-07 $layer=LI1_cond $X=11.647 $Y=0.87
+ $X2=11.647 $Y2=1.035
r240 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.475
+ $Y=0.87 $X2=11.475 $Y2=0.87
r241 21 55 46.5577 $w=3.26e-07 $l=2.89396e-07 $layer=POLY_cond $X=11.71 $Y=1.99
+ $X2=11.795 $Y2=1.74
r242 21 23 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=11.71 $Y=1.99
+ $X2=11.71 $Y2=2.275
r243 18 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.315 $Y=0.705
+ $X2=11.315 $Y2=0.87
r244 18 20 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=11.315 $Y=0.705
+ $X2=11.315 $Y2=0.415
r245 14 16 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=8.615 $Y=1.215
+ $X2=8.615 $Y2=0.415
r246 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.54 $Y=1.29
+ $X2=8.615 $Y2=1.215
r247 12 49 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=8.54 $Y=1.29
+ $X2=8.18 $Y2=1.29
r248 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.965 $Y=1.99
+ $X2=7.965 $Y2=2.275
r249 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.965 $Y=1.89 $X2=7.965
+ $Y2=1.99
r250 7 46 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=7.965 $Y=1.485
+ $X2=7.965 $Y2=1.35
r251 7 8 134.289 $w=2e-07 $l=4.05e-07 $layer=POLY_cond $X=7.965 $Y=1.485
+ $X2=7.965 $Y2=1.89
r252 2 62 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.815 $X2=1.2 $Y2=1.96
r253 1 58 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_1787_159# 1 2 8 9 11 14 17 18 20 23 27
+ 29 30 34 38 42 43 49 57
c125 42 0 6.25468e-20 $X=10.645 $Y=1.21
c126 9 0 1.04454e-19 $X=9.035 $Y=1.99
r127 51 52 4.69761 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=9.992 $Y=1.21
+ $X2=9.992 $Y2=1.375
r128 47 57 1.11087 $w=2.7e-07 $l=5e-09 $layer=POLY_cond $X=9.14 $Y=0.93
+ $X2=9.145 $Y2=0.93
r129 47 54 23.3282 $w=2.7e-07 $l=1.05e-07 $layer=POLY_cond $X=9.14 $Y=0.93
+ $X2=9.035 $Y2=0.93
r130 46 49 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.14 $Y=0.93
+ $X2=9.305 $Y2=0.93
r131 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.14
+ $Y=0.93 $X2=9.14 $Y2=0.93
r132 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.645
+ $Y=1.21 $X2=10.645 $Y2=1.21
r133 40 51 2.61955 $w=3.3e-07 $l=2.28e-07 $layer=LI1_cond $X=10.22 $Y=1.21
+ $X2=9.992 $Y2=1.21
r134 40 42 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=10.22 $Y=1.21
+ $X2=10.645 $Y2=1.21
r135 38 52 15.3154 $w=3.78e-07 $l=5.05e-07 $layer=LI1_cond $X=9.955 $Y=1.88
+ $X2=9.955 $Y2=1.375
r136 32 34 9.85779 $w=4.53e-07 $l=3.75e-07 $layer=LI1_cond $X=9.992 $Y=0.765
+ $X2=9.992 $Y2=0.39
r137 30 51 7.75479 $w=4.53e-07 $l=2.95e-07 $layer=LI1_cond $X=9.992 $Y=0.915
+ $X2=9.992 $Y2=1.21
r138 30 32 3.94312 $w=4.53e-07 $l=1.5e-07 $layer=LI1_cond $X=9.992 $Y=0.915
+ $X2=9.992 $Y2=0.765
r139 30 49 17.6708 $w=2.98e-07 $l=4.6e-07 $layer=LI1_cond $X=9.765 $Y=0.915
+ $X2=9.305 $Y2=0.915
r140 28 43 0.532654 $w=3.25e-07 $l=3e-09 $layer=POLY_cond $X=10.672 $Y=1.213
+ $X2=10.672 $Y2=1.21
r141 28 29 37.2436 $w=3.25e-07 $l=1.62e-07 $layer=POLY_cond $X=10.672 $Y=1.213
+ $X2=10.672 $Y2=1.375
r142 27 43 29.296 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=10.672 $Y=1.045
+ $X2=10.672 $Y2=1.21
r143 26 27 43.5133 $w=3.25e-07 $l=1.5e-07 $layer=POLY_cond $X=10.707 $Y=0.895
+ $X2=10.707 $Y2=1.045
r144 23 26 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=10.83 $Y=0.445
+ $X2=10.83 $Y2=0.895
r145 18 20 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=10.735 $Y=1.99
+ $X2=10.735 $Y2=2.275
r146 17 18 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=10.735 $Y=1.89
+ $X2=10.735 $Y2=1.99
r147 17 29 170.762 $w=2e-07 $l=5.15e-07 $layer=POLY_cond $X=10.735 $Y=1.89
+ $X2=10.735 $Y2=1.375
r148 12 57 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.145 $Y=0.795
+ $X2=9.145 $Y2=0.93
r149 12 14 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.145 $Y=0.795
+ $X2=9.145 $Y2=0.445
r150 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=9.035 $Y=1.99
+ $X2=9.035 $Y2=2.275
r151 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=9.035 $Y=1.89 $X2=9.035
+ $Y2=1.99
r152 7 54 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=9.035 $Y=1.065
+ $X2=9.035 $Y2=0.93
r153 7 8 273.551 $w=2e-07 $l=8.25e-07 $layer=POLY_cond $X=9.035 $Y=1.065
+ $X2=9.035 $Y2=1.89
r154 2 38 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=9.835
+ $Y=1.735 $X2=9.98 $Y2=1.88
r155 1 34 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=9.915
+ $Y=0.235 $X2=10.05 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_1611_413# 1 2 8 9 11 14 15 16 17 18 19
+ 23 28 30 32
c109 28 0 1.48265e-19 $X=8.78 $Y=1.315
c110 18 0 1.92092e-19 $X=9.745 $Y=1.467
c111 16 0 6.25468e-20 $X=9.78 $Y=1.1
r112 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.51
+ $Y=1.41 $X2=9.51 $Y2=1.41
r113 32 34 21.4122 $w=2.45e-07 $l=4.3e-07 $layer=LI1_cond $X=9.08 $Y=1.41
+ $X2=9.51 $Y2=1.41
r114 29 32 1.3646 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=9.08 $Y=1.575
+ $X2=9.08 $Y2=1.41
r115 29 30 31.4303 $w=2.18e-07 $l=6e-07 $layer=LI1_cond $X=9.08 $Y=1.575
+ $X2=9.08 $Y2=2.175
r116 28 32 14.9388 $w=2.45e-07 $l=3e-07 $layer=LI1_cond $X=8.78 $Y=1.41 $X2=9.08
+ $Y2=1.41
r117 27 28 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=8.78 $Y=0.565
+ $X2=8.78 $Y2=1.315
r118 23 27 7.59919 $w=3.1e-07 $l=1.92873e-07 $layer=LI1_cond $X=8.695 $Y=0.41
+ $X2=8.78 $Y2=0.565
r119 23 25 13.3832 $w=3.08e-07 $l=3.6e-07 $layer=LI1_cond $X=8.695 $Y=0.41
+ $X2=8.335 $Y2=0.41
r120 19 30 6.83662 $w=2e-07 $l=1.51987e-07 $layer=LI1_cond $X=8.97 $Y=2.275
+ $X2=9.08 $Y2=2.175
r121 19 21 41.8682 $w=1.98e-07 $l=7.55e-07 $layer=LI1_cond $X=8.97 $Y=2.275
+ $X2=8.215 $Y2=2.275
r122 17 35 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=9.645 $Y=1.41
+ $X2=9.51 $Y2=1.41
r123 17 18 0.448535 $w=2.7e-07 $l=1.253e-07 $layer=POLY_cond $X=9.645 $Y=1.41
+ $X2=9.745 $Y2=1.467
r124 15 16 54.0301 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=9.78 $Y=0.95 $X2=9.78
+ $Y2=1.1
r125 14 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=9.84 $Y=0.555
+ $X2=9.84 $Y2=0.95
r126 9 18 27.0491 $w=1.9e-07 $l=1.93e-07 $layer=POLY_cond $X=9.745 $Y=1.66
+ $X2=9.745 $Y2=1.467
r127 9 11 120.5 $w=1.8e-07 $l=4.5e-07 $layer=POLY_cond $X=9.745 $Y=1.66
+ $X2=9.745 $Y2=2.11
r128 8 18 27.0491 $w=1.9e-07 $l=1.92e-07 $layer=POLY_cond $X=9.745 $Y=1.275
+ $X2=9.745 $Y2=1.467
r129 8 16 58.026 $w=2e-07 $l=1.75e-07 $layer=POLY_cond $X=9.745 $Y=1.275
+ $X2=9.745 $Y2=1.1
r130 2 21 600 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_PDIFF $count=1 $X=8.055
+ $Y=2.065 $X2=8.215 $Y2=2.275
r131 1 25 182 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_NDIFF $count=1 $X=8.15
+ $Y=0.235 $X2=8.335 $Y2=0.41
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_2266_413# 1 2 7 11 13 15 16 17 18 20
+ 21 23 24 26 27 29 35 37 41 47 48 51 54 57 61
r136 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.07
+ $Y=1.74 $X2=14.07 $Y2=1.74
r137 57 60 43.9904 $w=2.7e-07 $l=1.98e-07 $layer=POLY_cond $X=14.07 $Y=1.542
+ $X2=14.07 $Y2=1.74
r138 54 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.07 $Y=1.87
+ $X2=14.07 $Y2=1.87
r139 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.25 $Y=1.87
+ $X2=12.25 $Y2=1.87
r140 48 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.395 $Y=1.87
+ $X2=12.25 $Y2=1.87
r141 47 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.925 $Y=1.87
+ $X2=14.07 $Y2=1.87
r142 47 48 1.89356 $w=1.4e-07 $l=1.53e-06 $layer=MET1_cond $X=13.925 $Y=1.87
+ $X2=12.395 $Y2=1.87
r143 46 51 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=12.25 $Y=2.165
+ $X2=12.25 $Y2=1.87
r144 45 51 61.5405 $w=2.48e-07 $l=1.335e-06 $layer=LI1_cond $X=12.25 $Y=0.535
+ $X2=12.25 $Y2=1.87
r145 41 45 6.90357 $w=2.05e-07 $l=1.68819e-07 $layer=LI1_cond $X=12.125 $Y=0.432
+ $X2=12.25 $Y2=0.535
r146 41 43 28.9446 $w=2.03e-07 $l=5.35e-07 $layer=LI1_cond $X=12.125 $Y=0.432
+ $X2=11.59 $Y2=0.432
r147 37 46 6.98266 $w=1.9e-07 $l=1.65831e-07 $layer=LI1_cond $X=12.125 $Y=2.26
+ $X2=12.25 $Y2=2.165
r148 37 39 37.9426 $w=1.88e-07 $l=6.5e-07 $layer=LI1_cond $X=12.125 $Y=2.26
+ $X2=11.475 $Y2=2.26
r149 35 36 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=15.77 $Y=1.202
+ $X2=15.795 $Y2=1.202
r150 34 35 59.6158 $w=3.8e-07 $l=4.7e-07 $layer=POLY_cond $X=15.3 $Y=1.202
+ $X2=15.77 $Y2=1.202
r151 33 34 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=15.275 $Y=1.202
+ $X2=15.3 $Y2=1.202
r152 27 36 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=15.795 $Y=0.995
+ $X2=15.795 $Y2=1.202
r153 27 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=15.795 $Y=0.995
+ $X2=15.795 $Y2=0.56
r154 24 35 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=15.77 $Y=1.41
+ $X2=15.77 $Y2=1.202
r155 24 26 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.77 $Y=1.41
+ $X2=15.77 $Y2=1.985
r156 21 34 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=15.3 $Y=1.41
+ $X2=15.3 $Y2=1.202
r157 21 23 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.3 $Y=1.41
+ $X2=15.3 $Y2=1.985
r158 18 33 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=15.275 $Y=0.995
+ $X2=15.275 $Y2=1.202
r159 18 20 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=15.275 $Y=0.995
+ $X2=15.275 $Y2=0.56
r160 17 32 126.662 $w=2e-07 $l=3.82e-07 $layer=POLY_cond $X=14.765 $Y=1.16
+ $X2=14.765 $Y2=1.542
r161 17 31 59.0037 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=14.765 $Y=1.16
+ $X2=14.765 $Y2=0.995
r162 16 33 10.4773 $w=3.8e-07 $l=9.3675e-08 $layer=POLY_cond $X=15.2 $Y=1.16
+ $X2=15.275 $Y2=1.202
r163 16 17 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=15.2 $Y=1.16
+ $X2=14.865 $Y2=1.16
r164 13 32 76.4073 $w=2e-07 $l=2.28e-07 $layer=POLY_cond $X=14.765 $Y=1.77
+ $X2=14.765 $Y2=1.542
r165 13 15 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=14.765 $Y=1.77
+ $X2=14.765 $Y2=2.165
r166 11 31 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=14.74 $Y=0.445
+ $X2=14.74 $Y2=0.995
r167 8 57 7.22716 $w=2.25e-07 $l=1.35e-07 $layer=POLY_cond $X=14.205 $Y=1.542
+ $X2=14.07 $Y2=1.542
r168 7 32 0.0601136 $w=2.25e-07 $l=1e-07 $layer=POLY_cond $X=14.665 $Y=1.542
+ $X2=14.765 $Y2=1.542
r169 7 8 131.195 $w=2.25e-07 $l=4.6e-07 $layer=POLY_cond $X=14.665 $Y=1.542
+ $X2=14.205 $Y2=1.542
r170 2 39 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=11.33
+ $Y=2.065 $X2=11.475 $Y2=2.26
r171 1 43 182 $w=1.7e-07 $l=2.82843e-07 $layer=licon1_NDIFF $count=1 $X=11.39
+ $Y=0.235 $X2=11.59 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 45 47
+ 51 55 59 63 67 73 79 84 85 87 88 90 91 92 94 99 111 122 126 136 137 140 143
+ 146 149 152 155 158
c228 137 0 1.77499e-19 $X=16.33 $Y=2.72
c229 1 0 1.03679e-19 $X=0.585 $Y=1.815
r230 158 159 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.95 $Y=2.72
+ $X2=14.95 $Y2=2.72
r231 155 156 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.57 $Y=2.72
+ $X2=13.57 $Y2=2.72
r232 153 156 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=13.57 $Y2=2.72
r233 152 153 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r234 149 150 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r235 147 150 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=9.43 $Y2=2.72
r236 146 147 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r237 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r238 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r239 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.33 $Y=2.72
+ $X2=16.33 $Y2=2.72
r240 134 137 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.87 $Y=2.72
+ $X2=16.33 $Y2=2.72
r241 134 159 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=15.87 $Y=2.72
+ $X2=14.95 $Y2=2.72
r242 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.87 $Y=2.72
+ $X2=15.87 $Y2=2.72
r243 131 158 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=15.15 $Y=2.72
+ $X2=15.032 $Y2=2.72
r244 131 133 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=15.15 $Y=2.72
+ $X2=15.87 $Y2=2.72
r245 130 159 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=14.03 $Y=2.72
+ $X2=14.95 $Y2=2.72
r246 130 156 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.03 $Y=2.72
+ $X2=13.57 $Y2=2.72
r247 129 130 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.03 $Y=2.72
+ $X2=14.03 $Y2=2.72
r248 127 155 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.785 $Y=2.72
+ $X2=13.66 $Y2=2.72
r249 127 129 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=13.785 $Y=2.72
+ $X2=14.03 $Y2=2.72
r250 126 158 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=14.915 $Y=2.72
+ $X2=15.032 $Y2=2.72
r251 126 129 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=14.915 $Y=2.72
+ $X2=14.03 $Y2=2.72
r252 125 153 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=12.65 $Y2=2.72
r253 124 125 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r254 122 152 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.595 $Y=2.72
+ $X2=12.68 $Y2=2.72
r255 122 124 116.455 $w=1.68e-07 $l=1.785e-06 $layer=LI1_cond $X=12.595 $Y=2.72
+ $X2=10.81 $Y2=2.72
r256 121 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=10.81 $Y2=2.72
r257 121 150 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=9.43 $Y2=2.72
r258 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r259 118 149 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=9.595 $Y=2.72
+ $X2=9.477 $Y2=2.72
r260 118 120 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=9.595 $Y=2.72
+ $X2=10.35 $Y2=2.72
r261 117 147 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r262 116 117 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r263 114 117 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=6.21 $Y2=2.72
r264 113 116 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=6.21 $Y2=2.72
r265 113 114 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r266 111 146 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=6.35 $Y=2.72
+ $X2=6.522 $Y2=2.72
r267 111 116 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.35 $Y=2.72
+ $X2=6.21 $Y2=2.72
r268 110 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r269 110 144 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r270 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r271 107 143 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.765 $Y=2.72
+ $X2=2.575 $Y2=2.72
r272 107 109 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=2.765 $Y=2.72
+ $X2=3.45 $Y2=2.72
r273 106 144 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r274 105 106 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r275 103 106 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r276 103 141 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r277 102 105 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r278 102 103 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r279 100 140 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r280 100 102 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r281 99 143 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.385 $Y=2.72
+ $X2=2.575 $Y2=2.72
r282 99 105 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.385 $Y=2.72
+ $X2=2.07 $Y2=2.72
r283 94 140 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r284 94 96 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r285 92 141 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r286 92 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r287 90 133 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=15.92 $Y=2.72
+ $X2=15.87 $Y2=2.72
r288 90 91 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=15.92 $Y=2.72
+ $X2=16.05 $Y2=2.72
r289 89 136 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=16.18 $Y=2.72
+ $X2=16.33 $Y2=2.72
r290 89 91 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=16.18 $Y=2.72
+ $X2=16.05 $Y2=2.72
r291 87 120 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=10.355 $Y=2.72
+ $X2=10.35 $Y2=2.72
r292 87 88 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=10.355 $Y=2.72
+ $X2=10.5 $Y2=2.72
r293 86 124 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.645 $Y=2.72
+ $X2=10.81 $Y2=2.72
r294 86 88 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=10.645 $Y=2.72
+ $X2=10.5 $Y2=2.72
r295 84 109 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.515 $Y=2.72
+ $X2=3.45 $Y2=2.72
r296 84 85 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=3.515 $Y=2.72
+ $X2=3.612 $Y2=2.72
r297 83 113 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.71 $Y=2.72
+ $X2=3.91 $Y2=2.72
r298 83 85 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=3.71 $Y=2.72
+ $X2=3.612 $Y2=2.72
r299 79 82 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=16.05 $Y=1.63
+ $X2=16.05 $Y2=2.31
r300 77 91 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=16.05 $Y=2.635
+ $X2=16.05 $Y2=2.72
r301 77 82 14.4055 $w=2.58e-07 $l=3.25e-07 $layer=LI1_cond $X=16.05 $Y=2.635
+ $X2=16.05 $Y2=2.31
r302 73 76 16.6736 $w=2.33e-07 $l=3.4e-07 $layer=LI1_cond $X=15.032 $Y=1.63
+ $X2=15.032 $Y2=1.97
r303 71 158 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=15.032 $Y=2.635
+ $X2=15.032 $Y2=2.72
r304 71 76 32.6117 $w=2.33e-07 $l=6.65e-07 $layer=LI1_cond $X=15.032 $Y=2.635
+ $X2=15.032 $Y2=1.97
r305 67 70 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=13.66 $Y=1.63
+ $X2=13.66 $Y2=2.31
r306 65 155 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.66 $Y=2.635
+ $X2=13.66 $Y2=2.72
r307 65 70 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=13.66 $Y=2.635
+ $X2=13.66 $Y2=2.31
r308 64 152 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.765 $Y=2.72
+ $X2=12.68 $Y2=2.72
r309 63 155 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.535 $Y=2.72
+ $X2=13.66 $Y2=2.72
r310 63 64 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=13.535 $Y=2.72
+ $X2=12.765 $Y2=2.72
r311 59 62 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=12.68 $Y=1.66
+ $X2=12.68 $Y2=2.34
r312 57 152 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.68 $Y=2.635
+ $X2=12.68 $Y2=2.72
r313 57 62 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.68 $Y=2.635
+ $X2=12.68 $Y2=2.34
r314 53 88 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=10.5 $Y=2.635
+ $X2=10.5 $Y2=2.72
r315 53 55 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=10.5 $Y=2.635
+ $X2=10.5 $Y2=2.275
r316 49 149 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=9.477 $Y=2.635
+ $X2=9.477 $Y2=2.72
r317 49 51 31.1405 $w=2.33e-07 $l=6.35e-07 $layer=LI1_cond $X=9.477 $Y=2.635
+ $X2=9.477 $Y2=2
r318 48 146 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=6.695 $Y=2.72
+ $X2=6.522 $Y2=2.72
r319 47 149 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=9.36 $Y=2.72
+ $X2=9.477 $Y2=2.72
r320 47 48 173.866 $w=1.68e-07 $l=2.665e-06 $layer=LI1_cond $X=9.36 $Y=2.72
+ $X2=6.695 $Y2=2.72
r321 43 146 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=6.522 $Y=2.635
+ $X2=6.522 $Y2=2.72
r322 43 45 9.85422 $w=3.43e-07 $l=2.95e-07 $layer=LI1_cond $X=6.522 $Y=2.635
+ $X2=6.522 $Y2=2.34
r323 39 85 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.612 $Y=2.635
+ $X2=3.612 $Y2=2.72
r324 39 41 36.6853 $w=1.93e-07 $l=6.45e-07 $layer=LI1_cond $X=3.612 $Y=2.635
+ $X2=3.612 $Y2=1.99
r325 35 143 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.575 $Y=2.635
+ $X2=2.575 $Y2=2.72
r326 35 37 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.575 $Y=2.635
+ $X2=2.575 $Y2=2
r327 31 140 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r328 31 33 12.5859 $w=3.78e-07 $l=4.15e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.22
r329 10 82 400 $w=1.7e-07 $l=8.99166e-07 $layer=licon1_PDIFF $count=1 $X=15.86
+ $Y=1.485 $X2=16.015 $Y2=2.31
r330 10 79 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=15.86
+ $Y=1.485 $X2=16.015 $Y2=1.63
r331 9 76 300 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=2 $X=14.855
+ $Y=1.845 $X2=15.065 $Y2=1.97
r332 9 73 600 $w=1.7e-07 $l=3.02283e-07 $layer=licon1_PDIFF $count=1 $X=14.855
+ $Y=1.845 $X2=15.065 $Y2=1.63
r333 8 70 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=13.475
+ $Y=1.485 $X2=13.62 $Y2=2.31
r334 8 67 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=13.475
+ $Y=1.485 $X2=13.62 $Y2=1.63
r335 7 62 400 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_PDIFF $count=1 $X=12.47
+ $Y=2.065 $X2=12.68 $Y2=2.34
r336 7 59 400 $w=1.7e-07 $l=4.99074e-07 $layer=licon1_PDIFF $count=1 $X=12.47
+ $Y=2.065 $X2=12.68 $Y2=1.66
r337 6 55 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=10.375
+ $Y=2.065 $X2=10.5 $Y2=2.275
r338 5 51 300 $w=1.7e-07 $l=3.86135e-07 $layer=licon1_PDIFF $count=2 $X=9.125
+ $Y=2.065 $X2=9.48 $Y2=2
r339 4 45 600 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_PDIFF $count=1 $X=6.285
+ $Y=1.845 $X2=6.49 $Y2=2.34
r340 3 41 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=3.445
+ $Y=1.845 $X2=3.6 $Y2=1.99
r341 2 37 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=2.455
+ $Y=1.845 $X2=2.6 $Y2=2
r342 1 33 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.815 $X2=0.73 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_319_47# 1 2 3 4 20 21 24 25 29 36 38
+ 40 43 48
r111 38 40 0.13119 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=4.62 $Y=0.51
+ $X2=4.425 $Y2=0.51
r112 38 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.62 $Y=0.51
+ $X2=4.62 $Y2=0.51
r113 36 40 2.34588 $w=1.85e-07 $l=2.74e-06 $layer=MET1_cond $X=1.685 $Y=0.487
+ $X2=4.425 $Y2=0.487
r114 34 48 7.97845 $w=2.58e-07 $l=1.8e-07 $layer=LI1_cond $X=1.54 $Y=0.385
+ $X2=1.72 $Y2=0.385
r115 33 36 0.0991101 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.54 $Y=0.51
+ $X2=1.685 $Y2=0.51
r116 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.54 $Y=0.51
+ $X2=1.54 $Y2=0.51
r117 28 43 19.2674 $w=3.18e-07 $l=5.35e-07 $layer=LI1_cond $X=4.605 $Y=0.98
+ $X2=4.605 $Y2=0.445
r118 28 29 8.64032 $w=3.18e-07 $l=1.7e-07 $layer=LI1_cond $X=4.655 $Y=0.98
+ $X2=4.655 $Y2=1.15
r119 25 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.78 $Y=1.82
+ $X2=4.78 $Y2=1.15
r120 24 25 9.22819 $w=4.38e-07 $l=1.8e-07 $layer=LI1_cond $X=4.645 $Y=2
+ $X2=4.645 $Y2=1.82
r121 20 21 7.04283 $w=4.28e-07 $l=1e-07 $layer=LI1_cond $X=1.67 $Y=1.99 $X2=1.67
+ $Y2=1.89
r122 13 34 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.54 $Y=0.515
+ $X2=1.54 $Y2=0.385
r123 13 21 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=1.54 $Y=0.515
+ $X2=1.54 $Y2=1.89
r124 4 24 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=4.495
+ $Y=1.845 $X2=4.64 $Y2=2
r125 3 20 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.595
+ $Y=1.845 $X2=1.72 $Y2=1.99
r126 2 43 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=4.505
+ $Y=0.235 $X2=4.64 $Y2=0.445
r127 1 48 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.72 $Y2=0.415
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%A_985_47# 1 2 3 4 15 18 20 23 26 29 31
+ 34 35 37 40 47 49 51 54 60
c128 49 0 1.67078e-19 $X=7.4 $Y=0.51
c129 29 0 5.64525e-20 $X=5.125 $Y=0.825
r130 49 51 0.13119 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=7.4 $Y=0.51
+ $X2=7.205 $Y2=0.51
r131 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.4 $Y=0.51 $X2=7.4
+ $Y2=0.51
r132 47 51 1.67808 $w=1.85e-07 $l=1.96e-06 $layer=MET1_cond $X=5.245 $Y=0.487
+ $X2=7.205 $Y2=0.487
r133 44 47 0.0991101 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.1 $Y=0.51
+ $X2=5.245 $Y2=0.51
r134 44 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.1 $Y=0.51 $X2=5.1
+ $Y2=0.51
r135 37 38 7.33994 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=7.625 $Y=2.34
+ $X2=7.625 $Y2=2.15
r136 35 40 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.625 $Y=1.185
+ $X2=7.625 $Y2=1.865
r137 31 32 4.83766 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=5.2 $Y=2.34 $X2=5.2
+ $Y2=2.21
r138 29 34 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.17 $Y=0.825
+ $X2=5.17 $Y2=1.785
r139 28 54 11.0909 $w=1.98e-07 $l=2e-07 $layer=LI1_cond $X=5.095 $Y=0.645
+ $X2=5.095 $Y2=0.445
r140 28 29 10.2632 $w=1.98e-07 $l=1.8e-07 $layer=LI1_cond $X=5.125 $Y=0.645
+ $X2=5.125 $Y2=0.825
r141 26 38 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=7.665 $Y=2
+ $X2=7.665 $Y2=2.15
r142 23 40 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=7.665 $Y=1.99
+ $X2=7.665 $Y2=1.865
r143 23 26 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=7.665 $Y=1.99
+ $X2=7.665 $Y2=2
r144 20 35 9.81506 $w=4.08e-07 $l=2.05e-07 $layer=LI1_cond $X=7.505 $Y=0.98
+ $X2=7.505 $Y2=1.185
r145 19 60 9.29389 $w=3.08e-07 $l=2.5e-07 $layer=LI1_cond $X=7.505 $Y=0.41
+ $X2=7.755 $Y2=0.41
r146 19 50 3.90344 $w=3.08e-07 $l=1.05e-07 $layer=LI1_cond $X=7.505 $Y=0.41
+ $X2=7.4 $Y2=0.41
r147 19 20 11.665 $w=4.08e-07 $l=4.15e-07 $layer=LI1_cond $X=7.505 $Y=0.565
+ $X2=7.505 $Y2=0.98
r148 18 32 8.64332 $w=2.78e-07 $l=2.1e-07 $layer=LI1_cond $X=5.225 $Y=2
+ $X2=5.225 $Y2=2.21
r149 15 34 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=5.225 $Y=1.925
+ $X2=5.225 $Y2=1.785
r150 15 18 3.0869 $w=2.78e-07 $l=7.5e-08 $layer=LI1_cond $X=5.225 $Y=1.925
+ $X2=5.225 $Y2=2
r151 4 37 600 $w=1.7e-07 $l=5.92832e-07 $layer=licon1_PDIFF $count=1 $X=7.41
+ $Y=1.845 $X2=7.625 $Y2=2.34
r152 4 26 600 $w=1.7e-07 $l=2.82046e-07 $layer=licon1_PDIFF $count=1 $X=7.41
+ $Y=1.845 $X2=7.625 $Y2=2
r153 3 31 600 $w=1.7e-07 $l=5.84423e-07 $layer=licon1_PDIFF $count=1 $X=5.005
+ $Y=1.845 $X2=5.2 $Y2=2.34
r154 3 18 600 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_PDIFF $count=1 $X=5.005
+ $Y=1.845 $X2=5.2 $Y2=2
r155 2 60 91 $w=1.7e-07 $l=6.15589e-07 $layer=licon1_NDIFF $count=2 $X=7.225
+ $Y=0.595 $X2=7.755 $Y2=0.41
r156 1 54 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=4.925
+ $Y=0.235 $X2=5.11 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%Q_N 1 2 9 15 17
r30 17 22 3.33383 $w=4.93e-07 $l=1.1e-07 $layer=LI1_cond $X=13.182 $Y=1.19
+ $X2=13.182 $Y2=1.3
r31 17 21 4.35249 $w=4.93e-07 $l=1.25e-07 $layer=LI1_cond $X=13.182 $Y=1.19
+ $X2=13.182 $Y2=1.065
r32 15 21 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=13.265 $Y=0.395
+ $X2=13.265 $Y2=1.065
r33 9 11 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=13.125 $Y=1.63
+ $X2=13.125 $Y2=2.31
r34 9 22 10.0081 $w=3.78e-07 $l=3.3e-07 $layer=LI1_cond $X=13.125 $Y=1.63
+ $X2=13.125 $Y2=1.3
r35 2 11 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=13.005
+ $Y=1.485 $X2=13.15 $Y2=2.31
r36 2 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=13.005
+ $Y=1.485 $X2=13.15 $Y2=1.63
r37 1 15 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=13.08
+ $Y=0.235 $X2=13.265 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%Q 1 2 7 10
r20 15 17 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=15.51 $Y=1.63
+ $X2=15.51 $Y2=2.31
r21 7 15 13.3441 $w=3.78e-07 $l=4.4e-07 $layer=LI1_cond $X=15.51 $Y=1.19
+ $X2=15.51 $Y2=1.63
r22 7 10 24.1103 $w=3.78e-07 $l=7.95e-07 $layer=LI1_cond $X=15.51 $Y=1.19
+ $X2=15.51 $Y2=0.395
r23 2 17 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=15.39
+ $Y=1.485 $X2=15.535 $Y2=2.31
r24 2 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=15.39
+ $Y=1.485 $X2=15.535 $Y2=1.63
r25 1 10 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=15.35
+ $Y=0.235 $X2=15.535 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HDLL__SEDFXBP_2%VGND 1 2 3 4 5 6 7 8 9 10 33 35 39 43 47
+ 51 55 61 65 71 74 75 77 78 80 81 82 84 89 97 105 114 122 131 132 136 142 145
+ 148 151 154 157
c234 132 0 1.88263e-19 $X=16.33 $Y=0
c235 105 0 1.67078e-19 $X=9.18 $Y=0
c236 61 0 8.50484e-20 $X=13.735 $Y=0.395
c237 43 0 1.87807e-19 $X=6.53 $Y=0.74
r238 157 158 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.95 $Y=0
+ $X2=14.95 $Y2=0
r239 154 155 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r240 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r241 148 149 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r242 145 146 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r243 143 146 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.45 $Y2=0
r244 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r245 136 139 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.38
r246 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r247 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.33 $Y=0
+ $X2=16.33 $Y2=0
r248 129 132 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.87 $Y=0
+ $X2=16.33 $Y2=0
r249 129 158 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=15.87 $Y=0
+ $X2=14.95 $Y2=0
r250 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.87 $Y=0
+ $X2=15.87 $Y2=0
r251 126 157 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=15.15 $Y=0
+ $X2=15.032 $Y2=0
r252 126 128 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=15.15 $Y=0
+ $X2=15.87 $Y2=0
r253 125 158 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=14.03 $Y=0
+ $X2=14.95 $Y2=0
r254 124 125 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.03 $Y=0
+ $X2=14.03 $Y2=0
r255 122 157 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=14.915 $Y=0
+ $X2=15.032 $Y2=0
r256 122 124 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=14.915 $Y=0
+ $X2=14.03 $Y2=0
r257 121 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=14.03 $Y2=0
r258 121 155 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=12.65 $Y2=0
r259 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r260 118 154 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.88 $Y=0
+ $X2=12.755 $Y2=0
r261 118 120 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=12.88 $Y=0
+ $X2=13.57 $Y2=0
r262 117 155 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=12.65 $Y2=0
r263 116 117 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r264 114 154 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.63 $Y=0
+ $X2=12.755 $Y2=0
r265 114 116 118.738 $w=1.68e-07 $l=1.82e-06 $layer=LI1_cond $X=12.63 $Y=0
+ $X2=10.81 $Y2=0
r266 113 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=10.81 $Y2=0
r267 113 152 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=9.43 $Y2=0
r268 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r269 110 151 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=9.575 $Y=0
+ $X2=9.377 $Y2=0
r270 110 112 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=9.575 $Y=0
+ $X2=10.35 $Y2=0
r271 109 152 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.43 $Y2=0
r272 109 149 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=6.67 $Y2=0
r273 108 109 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r274 106 148 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.695 $Y=0
+ $X2=6.57 $Y2=0
r275 106 108 148.422 $w=1.68e-07 $l=2.275e-06 $layer=LI1_cond $X=6.695 $Y=0
+ $X2=8.97 $Y2=0
r276 105 151 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=9.18 $Y=0
+ $X2=9.377 $Y2=0
r277 105 108 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.18 $Y=0
+ $X2=8.97 $Y2=0
r278 104 149 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=6.67 $Y2=0
r279 103 104 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r280 101 104 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=6.21 $Y2=0
r281 101 146 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=3.45 $Y2=0
r282 100 103 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=3.91 $Y=0
+ $X2=6.21 $Y2=0
r283 100 101 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r284 98 145 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.765 $Y=0
+ $X2=3.575 $Y2=0
r285 98 100 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.765 $Y=0
+ $X2=3.91 $Y2=0
r286 97 148 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.445 $Y=0
+ $X2=6.57 $Y2=0
r287 97 103 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.445 $Y=0
+ $X2=6.21 $Y2=0
r288 96 143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=2.53 $Y2=0
r289 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r290 93 96 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r291 93 137 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r292 92 95 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r293 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r294 90 136 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=0.705 $Y2=0
r295 90 92 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r296 89 142 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.385 $Y=0
+ $X2=2.575 $Y2=0
r297 89 95 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.385 $Y=0
+ $X2=2.07 $Y2=0
r298 84 136 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.705 $Y2=0
r299 84 86 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r300 82 137 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r301 82 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r302 80 128 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=15.92 $Y=0 $X2=15.87
+ $Y2=0
r303 80 81 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=15.92 $Y=0 $X2=16.05
+ $Y2=0
r304 79 131 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=16.18 $Y=0
+ $X2=16.33 $Y2=0
r305 79 81 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=16.18 $Y=0 $X2=16.05
+ $Y2=0
r306 77 120 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=13.65 $Y=0 $X2=13.57
+ $Y2=0
r307 77 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.65 $Y=0
+ $X2=13.775 $Y2=0
r308 76 124 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=13.9 $Y=0
+ $X2=14.03 $Y2=0
r309 76 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.9 $Y=0
+ $X2=13.775 $Y2=0
r310 74 112 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=10.45 $Y=0 $X2=10.35
+ $Y2=0
r311 74 75 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=10.45 $Y=0
+ $X2=10.587 $Y2=0
r312 73 116 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=10.725 $Y=0
+ $X2=10.81 $Y2=0
r313 73 75 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=10.725 $Y=0
+ $X2=10.587 $Y2=0
r314 69 81 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=16.05 $Y=0.085
+ $X2=16.05 $Y2=0
r315 69 71 13.7407 $w=2.58e-07 $l=3.1e-07 $layer=LI1_cond $X=16.05 $Y=0.085
+ $X2=16.05 $Y2=0.395
r316 65 67 16.6736 $w=2.33e-07 $l=3.4e-07 $layer=LI1_cond $X=15.032 $Y=0.395
+ $X2=15.032 $Y2=0.735
r317 63 157 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=15.032 $Y=0.085
+ $X2=15.032 $Y2=0
r318 63 65 15.2024 $w=2.33e-07 $l=3.1e-07 $layer=LI1_cond $X=15.032 $Y=0.085
+ $X2=15.032 $Y2=0.395
r319 59 78 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.775 $Y=0.085
+ $X2=13.775 $Y2=0
r320 59 61 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=13.775 $Y=0.085
+ $X2=13.775 $Y2=0.395
r321 55 57 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=12.755 $Y=0.395
+ $X2=12.755 $Y2=0.735
r322 53 154 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.755 $Y=0.085
+ $X2=12.755 $Y2=0
r323 53 55 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=12.755 $Y=0.085
+ $X2=12.755 $Y2=0.395
r324 49 75 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=10.587 $Y=0.085
+ $X2=10.587 $Y2=0
r325 49 51 15.2961 $w=2.73e-07 $l=3.65e-07 $layer=LI1_cond $X=10.587 $Y=0.085
+ $X2=10.587 $Y2=0.45
r326 45 151 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=9.377 $Y=0.085
+ $X2=9.377 $Y2=0
r327 45 47 9.77388 $w=3.93e-07 $l=3.35e-07 $layer=LI1_cond $X=9.377 $Y=0.085
+ $X2=9.377 $Y2=0.42
r328 41 148 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.57 $Y=0.085
+ $X2=6.57 $Y2=0
r329 41 43 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=6.57 $Y=0.085
+ $X2=6.57 $Y2=0.74
r330 37 145 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.575 $Y=0.085
+ $X2=3.575 $Y2=0
r331 37 39 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.575 $Y=0.085
+ $X2=3.575 $Y2=0.445
r332 36 142 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.765 $Y=0
+ $X2=2.575 $Y2=0
r333 35 145 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.385 $Y=0
+ $X2=3.575 $Y2=0
r334 35 36 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.385 $Y=0
+ $X2=2.765 $Y2=0
r335 31 142 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.575 $Y=0.085
+ $X2=2.575 $Y2=0
r336 31 33 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=2.575 $Y=0.085
+ $X2=2.575 $Y2=0.38
r337 10 71 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=15.87
+ $Y=0.235 $X2=16.015 $Y2=0.395
r338 9 67 182 $w=1.7e-07 $l=6.12372e-07 $layer=licon1_NDIFF $count=1 $X=14.815
+ $Y=0.235 $X2=15.065 $Y2=0.735
r339 9 65 182 $w=1.7e-07 $l=3.20156e-07 $layer=licon1_NDIFF $count=1 $X=14.815
+ $Y=0.235 $X2=15.065 $Y2=0.395
r340 8 61 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=13.55
+ $Y=0.235 $X2=13.735 $Y2=0.395
r341 7 57 182 $w=1.7e-07 $l=6.12372e-07 $layer=licon1_NDIFF $count=1 $X=12.545
+ $Y=0.235 $X2=12.795 $Y2=0.735
r342 7 55 182 $w=1.7e-07 $l=3.20156e-07 $layer=licon1_NDIFF $count=1 $X=12.545
+ $Y=0.235 $X2=12.795 $Y2=0.395
r343 6 51 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=10.445
+ $Y=0.235 $X2=10.57 $Y2=0.45
r344 5 47 182 $w=1.7e-07 $l=2.66927e-07 $layer=licon1_NDIFF $count=1 $X=9.22
+ $Y=0.235 $X2=9.41 $Y2=0.42
r345 4 43 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=6.345
+ $Y=0.595 $X2=6.53 $Y2=0.74
r346 3 39 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.455
+ $Y=0.235 $X2=3.6 $Y2=0.445
r347 2 33 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.6 $Y2=0.38
r348 1 139 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

