* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 Y a_120_297# a_396_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND B1 a_396_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR A1_N a_120_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 a_396_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND A1_N a_122_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_122_47# A2_N a_120_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR a_120_297# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 a_492_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 a_120_297# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 Y B2 a_492_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
