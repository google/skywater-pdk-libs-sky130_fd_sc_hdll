* NGSPICE file created from sky130_fd_sc_hdll__clkbuf_12.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__clkbuf_12 A VGND VNB VPB VPWR X
M1000 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=2.57e+12p pd=2.314e+07u as=1.74e+12p ps=1.548e+07u
M1001 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=6.804e+11p pd=8.28e+06u as=1.3482e+12p ps=1.398e+07u
M1002 VPWR A a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1003 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A a_117_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.268e+11p ps=2.76e+06u
M1010 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_117_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_117_297# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_117_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND A a_117_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_117_297# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

