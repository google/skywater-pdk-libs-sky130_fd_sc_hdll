* File: sky130_fd_sc_hdll__ebufn_8.spice
* Created: Thu Aug 27 19:07:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__ebufn_8.pex.spice"
.subckt sky130_fd_sc_hdll__ebufn_8  VNB VPB A TE_B VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* TE_B	TE_B
* A	A
* VPB	VPB
* VNB	VNB
MM1013 N_A_124_297#_M1013_d N_A_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.22425 PD=0.97 PS=1.99 NRD=0 NRS=11.076 M=1 R=4.33333 SA=75000.3
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1026 N_A_124_297#_M1013_d N_A_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.115375 PD=0.97 PS=1.005 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1007 N_A_321_47#_M1007_d N_TE_B_M1007_g N_VGND_M1026_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.115375 PD=1.92 PS=1.005 NRD=8.304 NRS=14.76 M=1
+ R=4.33333 SA=75001.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1009 N_A_485_47#_M1009_d N_A_321_47#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.12025 PD=1.92 PS=1.02 NRD=8.304 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75007.9 A=0.0975 P=1.6 MULT=1
MM1010 N_A_485_47#_M1010_d N_A_321_47#_M1010_g N_VGND_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.12025 PD=1.02 PS=1.02 NRD=8.304 NRS=8.304 M=1 R=4.33333
+ SA=75000.8 SB=75007.4 A=0.0975 P=1.6 MULT=1
MM1018 N_A_485_47#_M1010_d N_A_321_47#_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.12025 PD=1.02 PS=1.02 NRD=8.304 NRS=8.304 M=1 R=4.33333
+ SA=75001.3 SB=75006.9 A=0.0975 P=1.6 MULT=1
MM1019 N_A_485_47#_M1019_d N_A_321_47#_M1019_g N_VGND_M1018_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.12025 PD=1.02 PS=1.02 NRD=8.304 NRS=8.304 M=1 R=4.33333
+ SA=75001.8 SB=75006.4 A=0.0975 P=1.6 MULT=1
MM1022 N_A_485_47#_M1019_d N_A_321_47#_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.12025 PD=1.02 PS=1.02 NRD=8.304 NRS=8.304 M=1 R=4.33333
+ SA=75002.3 SB=75005.8 A=0.0975 P=1.6 MULT=1
MM1032 N_A_485_47#_M1032_d N_A_321_47#_M1032_g N_VGND_M1022_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.12025 PD=1.02 PS=1.02 NRD=8.304 NRS=8.304 M=1 R=4.33333
+ SA=75002.8 SB=75005.3 A=0.0975 P=1.6 MULT=1
MM1034 N_A_485_47#_M1032_d N_A_321_47#_M1034_g N_VGND_M1034_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.12025 PD=1.02 PS=1.02 NRD=8.304 NRS=8.304 M=1 R=4.33333
+ SA=75003.4 SB=75004.8 A=0.0975 P=1.6 MULT=1
MM1036 N_A_485_47#_M1036_d N_A_321_47#_M1036_g N_VGND_M1034_s VNB NSHORT L=0.15
+ W=0.65 AD=0.1885 AS=0.12025 PD=1.23 PS=1.02 NRD=33.228 NRS=8.304 M=1 R=4.33333
+ SA=75003.9 SB=75004.3 A=0.0975 P=1.6 MULT=1
MM1004 N_A_485_47#_M1036_d N_A_124_297#_M1004_g N_Z_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.1885 AS=0.104 PD=1.23 PS=0.97 NRD=22.152 NRS=8.304 M=1 R=4.33333
+ SA=75004.6 SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1011 N_A_485_47#_M1011_d N_A_124_297#_M1011_g N_Z_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75005.1 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1023 N_A_485_47#_M1011_d N_A_124_297#_M1023_g N_Z_M1023_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75005.5 SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1024 N_A_485_47#_M1024_d N_A_124_297#_M1024_g N_Z_M1023_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75006 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1025 N_A_485_47#_M1024_d N_A_124_297#_M1025_g N_Z_M1025_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75006.5 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1027 N_A_485_47#_M1027_d N_A_124_297#_M1027_g N_Z_M1025_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75007 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1029 N_A_485_47#_M1027_d N_A_124_297#_M1029_g N_Z_M1029_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75007.4 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1037 N_A_485_47#_M1037_d N_A_124_297#_M1037_g N_Z_M1029_s VNB NSHORT L=0.15
+ W=0.65 AD=0.182 AS=0.12025 PD=1.86 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75007.9 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g N_A_124_297#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.305 AS=0.145 PD=2.61 PS=1.29 NRD=3.9203 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1033 N_VPWR_M1033_d N_A_M1033_g N_A_124_297#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1875 AS=0.145 PD=1.375 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1014 N_A_321_47#_M1014_d N_TE_B_M1014_g N_VPWR_M1033_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.1875 PD=2.54 PS=1.375 NRD=0.9653 NRS=17.73 M=1 R=5.55556
+ SA=90001.2 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_TE_B_M1000_g N_A_437_309#_M1000_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1598 AS=0.2538 PD=1.28 PS=2.42 NRD=1.0441 NRS=1.0441 M=1 R=5.22222
+ SA=90000.2 SB=90008.1 A=0.1692 P=2.24 MULT=1
MM1001 N_VPWR_M1000_d N_TE_B_M1001_g N_A_437_309#_M1001_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1598 AS=0.1598 PD=1.28 PS=1.28 NRD=11.5245 NRS=1.0441 M=1
+ R=5.22222 SA=90000.7 SB=90007.6 A=0.1692 P=2.24 MULT=1
MM1002 N_VPWR_M1002_d N_TE_B_M1002_g N_A_437_309#_M1001_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1598 AS=0.1598 PD=1.28 PS=1.28 NRD=1.0441 NRS=11.5245 M=1
+ R=5.22222 SA=90001.2 SB=90007.1 A=0.1692 P=2.24 MULT=1
MM1003 N_VPWR_M1002_d N_TE_B_M1003_g N_A_437_309#_M1003_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1598 AS=0.1598 PD=1.28 PS=1.28 NRD=11.5245 NRS=1.0441 M=1
+ R=5.22222 SA=90001.7 SB=90006.6 A=0.1692 P=2.24 MULT=1
MM1006 N_VPWR_M1006_d N_TE_B_M1006_g N_A_437_309#_M1003_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1598 AS=0.1598 PD=1.28 PS=1.28 NRD=1.0441 NRS=11.5245 M=1
+ R=5.22222 SA=90002.3 SB=90006.1 A=0.1692 P=2.24 MULT=1
MM1012 N_VPWR_M1006_d N_TE_B_M1012_g N_A_437_309#_M1012_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1598 AS=0.1598 PD=1.28 PS=1.28 NRD=11.5245 NRS=1.0441 M=1
+ R=5.22222 SA=90002.8 SB=90005.5 A=0.1692 P=2.24 MULT=1
MM1016 N_VPWR_M1016_d N_TE_B_M1016_g N_A_437_309#_M1012_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1598 AS=0.1598 PD=1.28 PS=1.28 NRD=1.0441 NRS=11.5245 M=1
+ R=5.22222 SA=90003.3 SB=90005 A=0.1692 P=2.24 MULT=1
MM1021 N_VPWR_M1016_d N_TE_B_M1021_g N_A_437_309#_M1021_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1598 AS=0.404539 PD=1.28 PS=1.78309 NRD=11.5245 NRS=18.8529 M=1
+ R=5.22222 SA=90003.8 SB=90004.5 A=0.1692 P=2.24 MULT=1
MM1008 N_A_437_309#_M1021_s N_A_124_297#_M1008_g N_Z_M1008_s VPB PHIGHVT L=0.18
+ W=1 AD=0.430361 AS=0.145 PD=1.89691 PS=1.29 NRD=15.7403 NRS=0.9653 M=1
+ R=5.55556 SA=90004.6 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1015 N_A_437_309#_M1015_d N_A_124_297#_M1015_g N_Z_M1008_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.1 SB=90003 A=0.18 P=2.36 MULT=1
MM1017 N_A_437_309#_M1015_d N_A_124_297#_M1017_g N_Z_M1017_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.5 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1020 N_A_437_309#_M1020_d N_A_124_297#_M1020_g N_Z_M1017_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90006 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1028 N_A_437_309#_M1020_d N_A_124_297#_M1028_g N_Z_M1028_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90006.5 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1030 N_A_437_309#_M1030_d N_A_124_297#_M1030_g N_Z_M1028_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90006.9 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1031 N_A_437_309#_M1030_d N_A_124_297#_M1031_g N_Z_M1031_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90007.4 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1035 N_A_437_309#_M1035_d N_A_124_297#_M1035_g N_Z_M1031_s VPB PHIGHVT L=0.18
+ W=1 AD=0.29 AS=0.145 PD=2.58 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90007.9 SB=90000.2 A=0.18 P=2.36 MULT=1
DX38_noxref VNB VPB NWDIODE A=18.3291 P=26.05
pX39_noxref noxref_12 TE_B TE_B PROBETYPE=1
pX40_noxref noxref_13 TE_B TE_B PROBETYPE=1
*
.include "sky130_fd_sc_hdll__ebufn_8.pxi.spice"
*
.ends
*
*
