* File: sky130_fd_sc_hdll__nand4_2.spice
* Created: Wed Sep  2 08:38:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nand4_2.pex.spice"
.subckt sky130_fd_sc_hdll__nand4_2  VNB VPB D C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1002 N_A_27_47#_M1002_d N_D_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1012 N_A_27_47#_M1012_d N_D_M1012_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1005 N_A_297_47#_M1005_d N_C_M1005_g N_A_27_47#_M1012_d VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1013 N_A_297_47#_M1005_d N_C_M1013_g N_A_27_47#_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.182 PD=1.02 PS=1.86 NRD=8.304 NRS=2.76 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_511_47#_M1004_d N_B_M1004_g N_A_297_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.247 AS=0.104 PD=2.06 PS=0.97 NRD=11.988 NRS=0 M=1 R=4.33333
+ SA=75000.3 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1010 N_A_511_47#_M1010_d N_B_M1010_g N_A_297_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.8 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1007 N_A_511_47#_M1010_d N_A_M1007_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.2
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1008 N_A_511_47#_M1008_d N_A_M1008_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2665 AS=0.104 PD=2.12 PS=0.97 NRD=23.076 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_D_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90004.2 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_D_M1009_g N_Y_M1000_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.6
+ SB=90003.8 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1009_d N_C_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.1
+ SB=90003.3 A=0.18 P=2.36 MULT=1
MM1015 N_VPWR_M1015_d N_C_M1015_g N_Y_M1011_s VPB PHIGHVT L=0.18 W=1 AD=0.225
+ AS=0.145 PD=1.45 PS=1.29 NRD=16.7253 NRS=0.9653 M=1 R=5.55556 SA=90001.6
+ SB=90002.8 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1015_d N_B_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1 AD=0.225
+ AS=0.145 PD=1.45 PS=1.29 NRD=16.7253 NRS=0.9653 M=1 R=5.55556 SA=90002.2
+ SB=90002.2 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_B_M1006_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1 AD=0.37
+ AS=0.145 PD=1.74 PS=1.29 NRD=44.3053 NRS=0.9653 M=1 R=5.55556 SA=90002.7
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g N_VPWR_M1006_d VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.37 PD=1.29 PS=1.74 NRD=0.9653 NRS=46.2753 M=1 R=5.55556 SA=90003.6
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1014 N_Y_M1003_d N_A_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.43 PD=1.29 PS=2.86 NRD=0.9653 NRS=16.7253 M=1 R=5.55556 SA=90004.1
+ SB=90000.3 A=0.18 P=2.36 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.7312 P=14.09
*
.include "sky130_fd_sc_hdll__nand4_2.pxi.spice"
*
.ends
*
*
