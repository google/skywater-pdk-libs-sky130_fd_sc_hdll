* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
X0 a_331_413# a_27_410# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_27_410# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND D_N a_216_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR a_331_413# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 a_331_413# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND a_331_413# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND a_216_93# a_331_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_527_297# B a_609_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X8 a_27_410# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X9 VGND B a_331_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR D_N a_216_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X11 a_609_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X12 a_331_413# a_216_93# a_421_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X13 a_421_413# a_27_410# a_527_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
.ends
