* File: sky130_fd_sc_hdll__xor2_1.pxi.spice
* Created: Thu Aug 27 19:29:45 2020
* 
x_PM_SKY130_FD_SC_HDLL__XOR2_1%B N_B_c_55_n N_B_M1006_g N_B_c_56_n N_B_M1002_g
+ N_B_c_57_n N_B_M1005_g N_B_c_58_n N_B_M1008_g N_B_c_59_n N_B_c_60_n N_B_c_65_n
+ B N_B_c_61_n PM_SKY130_FD_SC_HDLL__XOR2_1%B
x_PM_SKY130_FD_SC_HDLL__XOR2_1%A N_A_c_131_n N_A_M1003_g N_A_c_134_n N_A_M1000_g
+ N_A_c_135_n N_A_M1009_g N_A_c_132_n N_A_M1007_g A N_A_c_133_n
+ PM_SKY130_FD_SC_HDLL__XOR2_1%A
x_PM_SKY130_FD_SC_HDLL__XOR2_1%A_35_297# N_A_35_297#_M1002_d N_A_35_297#_M1006_s
+ N_A_35_297#_c_179_n N_A_35_297#_M1001_g N_A_35_297#_c_174_n
+ N_A_35_297#_M1004_g N_A_35_297#_c_180_n N_A_35_297#_c_181_n
+ N_A_35_297#_c_188_n N_A_35_297#_c_175_n N_A_35_297#_c_238_p
+ N_A_35_297#_c_190_n N_A_35_297#_c_176_n N_A_35_297#_c_177_n
+ N_A_35_297#_c_202_n N_A_35_297#_c_178_n PM_SKY130_FD_SC_HDLL__XOR2_1%A_35_297#
x_PM_SKY130_FD_SC_HDLL__XOR2_1%VPWR N_VPWR_M1000_d N_VPWR_M1005_d N_VPWR_c_257_n
+ N_VPWR_c_258_n N_VPWR_c_259_n N_VPWR_c_260_n N_VPWR_c_261_n N_VPWR_c_262_n
+ VPWR N_VPWR_c_263_n N_VPWR_c_256_n PM_SKY130_FD_SC_HDLL__XOR2_1%VPWR
x_PM_SKY130_FD_SC_HDLL__XOR2_1%A_315_297# N_A_315_297#_M1009_d
+ N_A_315_297#_M1001_s N_A_315_297#_c_300_n N_A_315_297#_c_306_n
+ N_A_315_297#_c_301_n PM_SKY130_FD_SC_HDLL__XOR2_1%A_315_297#
x_PM_SKY130_FD_SC_HDLL__XOR2_1%X N_X_M1008_d N_X_M1001_d N_X_c_328_n N_X_c_324_n
+ X X PM_SKY130_FD_SC_HDLL__XOR2_1%X
x_PM_SKY130_FD_SC_HDLL__XOR2_1%VGND N_VGND_M1002_s N_VGND_M1003_d N_VGND_M1004_d
+ N_VGND_c_349_n N_VGND_c_350_n N_VGND_c_351_n N_VGND_c_352_n N_VGND_c_353_n
+ VGND N_VGND_c_354_n N_VGND_c_355_n N_VGND_c_356_n N_VGND_c_357_n
+ PM_SKY130_FD_SC_HDLL__XOR2_1%VGND
cc_1 VNB N_B_c_55_n 0.0243341f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.41
cc_2 VNB N_B_c_56_n 0.0197111f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=0.995
cc_3 VNB N_B_c_57_n 0.0223939f $X=-0.19 $Y=-0.24 $X2=1.965 $Y2=1.41
cc_4 VNB N_B_c_58_n 0.0206055f $X=-0.19 $Y=-0.24 $X2=1.99 $Y2=0.995
cc_5 VNB N_B_c_59_n 6.88268e-19 $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.445
cc_6 VNB N_B_c_60_n 0.00589395f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.16
cc_7 VNB N_B_c_61_n 0.00709878f $X=-0.19 $Y=-0.24 $X2=0.57 $Y2=1.16
cc_8 VNB N_A_c_131_n 0.0170298f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.41
cc_9 VNB N_A_c_132_n 0.0177205f $X=-0.19 $Y=-0.24 $X2=1.99 $Y2=0.995
cc_10 VNB N_A_c_133_n 0.0371053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_35_297#_c_174_n 0.0231874f $X=-0.19 $Y=-0.24 $X2=1.99 $Y2=0.995
cc_12 VNB N_A_35_297#_c_175_n 0.00850627f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_35_297#_c_176_n 0.00531955f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.16
cc_14 VNB N_A_35_297#_c_177_n 0.0222346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_35_297#_c_178_n 0.0435543f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.445
cc_16 VNB N_VPWR_c_256_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_X_c_324_n 0.0135385f $X=-0.19 $Y=-0.24 $X2=1.99 $Y2=0.56
cc_18 VNB N_VGND_c_349_n 0.0126079f $X=-0.19 $Y=-0.24 $X2=1.99 $Y2=0.995
cc_19 VNB N_VGND_c_350_n 0.0145224f $X=-0.19 $Y=-0.24 $X2=1.99 $Y2=0.56
cc_20 VNB N_VGND_c_351_n 0.00299877f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_352_n 0.0120854f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.16
cc_22 VNB N_VGND_c_353_n 0.0362482f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_354_n 0.0139516f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_355_n 0.0464433f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.16
cc_25 VNB N_VGND_c_356_n 0.00603303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_357_n 0.201385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VPB N_B_c_55_n 0.0286696f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=1.41
cc_28 VPB N_B_c_57_n 0.0318203f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=1.41
cc_29 VPB N_B_c_59_n 0.00130718f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=1.445
cc_30 VPB N_B_c_65_n 0.00629631f $X=-0.19 $Y=1.305 $X2=1.72 $Y2=1.53
cc_31 VPB B 3.66229e-19 $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.445
cc_32 VPB N_B_c_61_n 0.00272548f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=1.16
cc_33 VPB N_A_c_134_n 0.0160347f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=0.995
cc_34 VPB N_A_c_135_n 0.0160346f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=1.41
cc_35 VPB N_A_c_133_n 0.0193513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_35_297#_c_179_n 0.0244382f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=1.41
cc_37 VPB N_A_35_297#_c_180_n 0.00782983f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=1.16
cc_38 VPB N_A_35_297#_c_181_n 0.0207996f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=1.16
cc_39 VPB N_A_35_297#_c_176_n 0.00348787f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=1.16
cc_40 VPB N_A_35_297#_c_177_n 0.0196401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_35_297#_c_178_n 0.0207778f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.445
cc_42 VPB N_VPWR_c_257_n 0.00469739f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=1.985
cc_43 VPB N_VPWR_c_258_n 0.00474148f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=1.245
cc_44 VPB N_VPWR_c_259_n 0.035534f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_260_n 0.00324069f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=1.16
cc_46 VPB N_VPWR_c_261_n 0.0209591f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=1.16
cc_47 VPB N_VPWR_c_262_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_263_n 0.0397991f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_256_n 0.0492091f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_315_297#_c_300_n 0.00731822f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=1.985
cc_51 VPB N_A_315_297#_c_301_n 0.0117534f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_X_c_324_n 0.00214401f $X=-0.19 $Y=1.305 $X2=1.99 $Y2=0.56
cc_53 VPB X 0.0367116f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=1.245
cc_54 VPB X 0.0183038f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=1.16
cc_55 N_B_c_56_n N_A_c_131_n 0.0233733f $X=0.56 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_56 N_B_c_55_n N_A_c_134_n 0.0500536f $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_57 N_B_c_65_n N_A_c_134_n 0.0178438f $X=1.72 $Y=1.53 $X2=0 $Y2=0
cc_58 N_B_c_61_n N_A_c_134_n 8.42217e-19 $X=0.57 $Y=1.16 $X2=0 $Y2=0
cc_59 N_B_c_57_n N_A_c_135_n 0.0212654f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_60 N_B_c_59_n N_A_c_135_n 7.37913e-19 $X=1.805 $Y=1.445 $X2=0 $Y2=0
cc_61 N_B_c_65_n N_A_c_135_n 0.0163362f $X=1.72 $Y=1.53 $X2=0 $Y2=0
cc_62 N_B_c_58_n N_A_c_132_n 0.0353115f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_63 N_B_c_55_n A 2.01976e-19 $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_64 N_B_c_59_n A 0.00187374f $X=1.805 $Y=1.445 $X2=0 $Y2=0
cc_65 N_B_c_60_n A 0.0117085f $X=1.93 $Y=1.16 $X2=0 $Y2=0
cc_66 N_B_c_65_n A 0.0384921f $X=1.72 $Y=1.53 $X2=0 $Y2=0
cc_67 N_B_c_61_n A 0.0157167f $X=0.57 $Y=1.16 $X2=0 $Y2=0
cc_68 N_B_c_55_n N_A_c_133_n 0.0251372f $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_69 N_B_c_57_n N_A_c_133_n 0.026093f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_70 N_B_c_59_n N_A_c_133_n 0.00317065f $X=1.805 $Y=1.445 $X2=0 $Y2=0
cc_71 N_B_c_60_n N_A_c_133_n 0.00127117f $X=1.93 $Y=1.16 $X2=0 $Y2=0
cc_72 N_B_c_65_n N_A_c_133_n 0.00810508f $X=1.72 $Y=1.53 $X2=0 $Y2=0
cc_73 N_B_c_61_n N_A_c_133_n 0.00675021f $X=0.57 $Y=1.16 $X2=0 $Y2=0
cc_74 N_B_c_55_n N_A_35_297#_c_180_n 0.00431969f $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_75 B N_A_35_297#_c_180_n 0.00159714f $X=0.655 $Y=1.445 $X2=0 $Y2=0
cc_76 N_B_c_55_n N_A_35_297#_c_181_n 0.0094805f $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_77 N_B_c_56_n N_A_35_297#_c_188_n 0.0130275f $X=0.56 $Y=0.995 $X2=0 $Y2=0
cc_78 N_B_c_61_n N_A_35_297#_c_188_n 0.0159787f $X=0.57 $Y=1.16 $X2=0 $Y2=0
cc_79 N_B_c_57_n N_A_35_297#_c_190_n 0.00279205f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_80 N_B_c_58_n N_A_35_297#_c_190_n 0.0131484f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_81 N_B_c_60_n N_A_35_297#_c_190_n 0.0198815f $X=1.93 $Y=1.16 $X2=0 $Y2=0
cc_82 N_B_c_65_n N_A_35_297#_c_190_n 0.0070073f $X=1.72 $Y=1.53 $X2=0 $Y2=0
cc_83 N_B_c_57_n N_A_35_297#_c_176_n 0.00122617f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_84 N_B_c_58_n N_A_35_297#_c_176_n 0.0058744f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_85 N_B_c_59_n N_A_35_297#_c_176_n 0.00218954f $X=1.805 $Y=1.445 $X2=0 $Y2=0
cc_86 N_B_c_60_n N_A_35_297#_c_176_n 0.00829779f $X=1.93 $Y=1.16 $X2=0 $Y2=0
cc_87 N_B_c_55_n N_A_35_297#_c_177_n 0.010044f $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_88 N_B_c_56_n N_A_35_297#_c_177_n 0.00542458f $X=0.56 $Y=0.995 $X2=0 $Y2=0
cc_89 B N_A_35_297#_c_177_n 0.008073f $X=0.655 $Y=1.445 $X2=0 $Y2=0
cc_90 N_B_c_61_n N_A_35_297#_c_177_n 0.0357971f $X=0.57 $Y=1.16 $X2=0 $Y2=0
cc_91 N_B_c_65_n N_A_35_297#_c_202_n 0.00250422f $X=1.72 $Y=1.53 $X2=0 $Y2=0
cc_92 N_B_c_61_n N_A_35_297#_c_202_n 0.00754392f $X=0.57 $Y=1.16 $X2=0 $Y2=0
cc_93 N_B_c_57_n N_A_35_297#_c_178_n 0.0074115f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_94 N_B_c_60_n N_A_35_297#_c_178_n 7.46431e-19 $X=1.93 $Y=1.16 $X2=0 $Y2=0
cc_95 N_B_c_65_n A_125_297# 0.00351031f $X=1.72 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_96 B A_125_297# 0.00410451f $X=0.655 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_97 N_B_c_65_n N_VPWR_M1000_d 0.00178587f $X=1.72 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_98 N_B_c_65_n N_VPWR_c_257_n 0.0136682f $X=1.72 $Y=1.53 $X2=0 $Y2=0
cc_99 N_B_c_57_n N_VPWR_c_258_n 0.00592966f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_100 N_B_c_55_n N_VPWR_c_259_n 0.00673617f $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_101 N_B_c_57_n N_VPWR_c_261_n 0.00688798f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_102 N_B_c_55_n N_VPWR_c_256_n 0.0130168f $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_103 N_B_c_57_n N_VPWR_c_256_n 0.00830105f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_104 N_B_c_65_n N_A_315_297#_M1009_d 0.00197851f $X=1.72 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_105 N_B_c_57_n N_A_315_297#_c_300_n 0.014638f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_106 N_B_c_60_n N_A_315_297#_c_300_n 0.00666299f $X=1.93 $Y=1.16 $X2=0 $Y2=0
cc_107 N_B_c_65_n N_A_315_297#_c_300_n 2.89797e-19 $X=1.72 $Y=1.53 $X2=0 $Y2=0
cc_108 N_B_c_57_n N_A_315_297#_c_306_n 0.00795433f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_109 N_B_c_65_n N_A_315_297#_c_306_n 0.0216384f $X=1.72 $Y=1.53 $X2=0 $Y2=0
cc_110 N_B_c_57_n N_A_315_297#_c_301_n 0.00338109f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_111 N_B_c_58_n N_X_c_328_n 0.00694695f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_112 N_B_c_56_n N_VGND_c_350_n 0.00332197f $X=0.56 $Y=0.995 $X2=0 $Y2=0
cc_113 N_B_c_56_n N_VGND_c_351_n 7.28296e-19 $X=0.56 $Y=0.995 $X2=0 $Y2=0
cc_114 N_B_c_56_n N_VGND_c_354_n 0.00428022f $X=0.56 $Y=0.995 $X2=0 $Y2=0
cc_115 N_B_c_58_n N_VGND_c_355_n 0.00370116f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_116 N_B_c_56_n N_VGND_c_357_n 0.00676791f $X=0.56 $Y=0.995 $X2=0 $Y2=0
cc_117 N_B_c_58_n N_VGND_c_357_n 0.00675389f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A_c_134_n N_A_35_297#_c_180_n 0.00313866f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_c_131_n N_A_35_297#_c_190_n 0.0125083f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A_c_132_n N_A_35_297#_c_190_n 0.0140611f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_121 A N_A_35_297#_c_190_n 0.02527f $X=1.175 $Y=1.105 $X2=0 $Y2=0
cc_122 N_A_c_133_n N_A_35_297#_c_190_n 0.00443538f $X=1.485 $Y=1.202 $X2=0 $Y2=0
cc_123 N_A_c_134_n N_VPWR_c_257_n 0.0163121f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A_c_135_n N_VPWR_c_257_n 0.00488595f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A_c_134_n N_VPWR_c_259_n 0.00702461f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A_c_135_n N_VPWR_c_261_n 0.00597712f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A_c_134_n N_VPWR_c_256_n 0.0126382f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A_c_135_n N_VPWR_c_256_n 0.0100435f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_c_135_n N_A_315_297#_c_306_n 0.0110607f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_c_131_n N_VGND_c_351_n 0.00776987f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_c_132_n N_VGND_c_351_n 0.00325012f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_c_131_n N_VGND_c_354_n 0.00341689f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_c_132_n N_VGND_c_355_n 0.00428022f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_c_131_n N_VGND_c_357_n 0.0040799f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_c_132_n N_VGND_c_357_n 0.00610074f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_35_297#_c_179_n N_VPWR_c_258_n 0.00228722f $X=2.955 $Y=1.41 $X2=0
+ $Y2=0
cc_137 N_A_35_297#_c_181_n N_VPWR_c_259_n 0.0246443f $X=0.3 $Y=2 $X2=0 $Y2=0
cc_138 N_A_35_297#_c_179_n N_VPWR_c_263_n 0.00702461f $X=2.955 $Y=1.41 $X2=0
+ $Y2=0
cc_139 N_A_35_297#_M1006_s N_VPWR_c_256_n 0.00217517f $X=0.175 $Y=1.485 $X2=0
+ $Y2=0
cc_140 N_A_35_297#_c_179_n N_VPWR_c_256_n 0.0150744f $X=2.955 $Y=1.41 $X2=0
+ $Y2=0
cc_141 N_A_35_297#_c_181_n N_VPWR_c_256_n 0.0143981f $X=0.3 $Y=2 $X2=0 $Y2=0
cc_142 N_A_35_297#_c_176_n N_A_315_297#_c_301_n 0.00936215f $X=2.66 $Y=1.16
+ $X2=0 $Y2=0
cc_143 N_A_35_297#_c_178_n N_A_315_297#_c_301_n 0.00426664f $X=2.955 $Y=1.202
+ $X2=0 $Y2=0
cc_144 N_A_35_297#_c_190_n N_X_M1008_d 0.0264339f $X=2.515 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_145 N_A_35_297#_c_176_n N_X_M1008_d 0.00139844f $X=2.66 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_146 N_A_35_297#_c_174_n N_X_c_328_n 0.0109707f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_35_297#_c_190_n N_X_c_328_n 0.0545166f $X=2.515 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A_35_297#_c_178_n N_X_c_328_n 0.00439655f $X=2.955 $Y=1.202 $X2=0 $Y2=0
cc_149 N_A_35_297#_c_174_n N_X_c_324_n 0.0219177f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A_35_297#_c_190_n N_X_c_324_n 0.0134183f $X=2.515 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A_35_297#_c_176_n N_X_c_324_n 0.035203f $X=2.66 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_35_297#_c_178_n N_X_c_324_n 0.0166498f $X=2.955 $Y=1.202 $X2=0 $Y2=0
cc_153 N_A_35_297#_c_179_n X 0.0245578f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_35_297#_c_179_n X 0.0153559f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_35_297#_c_178_n X 0.00408656f $X=2.955 $Y=1.202 $X2=0 $Y2=0
cc_156 N_A_35_297#_c_188_n N_VGND_M1002_s 0.00872414f $X=0.685 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_157 N_A_35_297#_c_175_n N_VGND_M1002_s 0.00162757f $X=0.255 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_158 N_A_35_297#_c_177_n N_VGND_M1002_s 9.73118e-19 $X=0.275 $Y=1.785
+ $X2=-0.19 $Y2=-0.24
cc_159 N_A_35_297#_c_190_n N_VGND_M1003_d 0.00547059f $X=2.515 $Y=0.74 $X2=0
+ $Y2=0
cc_160 N_A_35_297#_c_175_n N_VGND_c_349_n 9.77208e-19 $X=0.255 $Y=0.74 $X2=0
+ $Y2=0
cc_161 N_A_35_297#_c_188_n N_VGND_c_350_n 0.0125954f $X=0.685 $Y=0.74 $X2=0
+ $Y2=0
cc_162 N_A_35_297#_c_175_n N_VGND_c_350_n 0.00971556f $X=0.255 $Y=0.74 $X2=0
+ $Y2=0
cc_163 N_A_35_297#_c_238_p N_VGND_c_351_n 0.00999963f $X=0.77 $Y=0.5 $X2=0 $Y2=0
cc_164 N_A_35_297#_c_190_n N_VGND_c_351_n 0.0206198f $X=2.515 $Y=0.74 $X2=0
+ $Y2=0
cc_165 N_A_35_297#_c_174_n N_VGND_c_353_n 0.0103911f $X=2.98 $Y=0.995 $X2=0
+ $Y2=0
cc_166 N_A_35_297#_c_188_n N_VGND_c_354_n 0.0029785f $X=0.685 $Y=0.74 $X2=0
+ $Y2=0
cc_167 N_A_35_297#_c_238_p N_VGND_c_354_n 0.00747591f $X=0.77 $Y=0.5 $X2=0 $Y2=0
cc_168 N_A_35_297#_c_190_n N_VGND_c_354_n 0.00241682f $X=2.515 $Y=0.74 $X2=0
+ $Y2=0
cc_169 N_A_35_297#_c_174_n N_VGND_c_355_n 0.0036993f $X=2.98 $Y=0.995 $X2=0
+ $Y2=0
cc_170 N_A_35_297#_c_190_n N_VGND_c_355_n 0.00687326f $X=2.515 $Y=0.74 $X2=0
+ $Y2=0
cc_171 N_A_35_297#_M1002_d N_VGND_c_357_n 0.00271058f $X=0.635 $Y=0.235 $X2=0
+ $Y2=0
cc_172 N_A_35_297#_c_174_n N_VGND_c_357_n 0.00782537f $X=2.98 $Y=0.995 $X2=0
+ $Y2=0
cc_173 N_A_35_297#_c_188_n N_VGND_c_357_n 0.00624268f $X=0.685 $Y=0.74 $X2=0
+ $Y2=0
cc_174 N_A_35_297#_c_175_n N_VGND_c_357_n 0.0021233f $X=0.255 $Y=0.74 $X2=0
+ $Y2=0
cc_175 N_A_35_297#_c_238_p N_VGND_c_357_n 0.00613703f $X=0.77 $Y=0.5 $X2=0 $Y2=0
cc_176 N_A_35_297#_c_190_n N_VGND_c_357_n 0.0193926f $X=2.515 $Y=0.74 $X2=0
+ $Y2=0
cc_177 N_A_35_297#_c_190_n A_317_47# 0.00698512f $X=2.515 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_178 A_125_297# N_VPWR_c_256_n 0.0128237f $X=0.625 $Y=1.485 $X2=0 $Y2=0
cc_179 N_VPWR_c_256_n N_A_315_297#_M1009_d 0.00239291f $X=3.45 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_180 N_VPWR_c_256_n N_A_315_297#_M1001_s 0.00252233f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_181 N_VPWR_M1005_d N_A_315_297#_c_300_n 0.0106576f $X=2.055 $Y=1.485 $X2=0
+ $Y2=0
cc_182 N_VPWR_c_258_n N_A_315_297#_c_300_n 0.0132786f $X=2.2 $Y=2.29 $X2=0 $Y2=0
cc_183 N_VPWR_c_256_n N_A_315_297#_c_300_n 0.0140433f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_184 N_VPWR_c_257_n N_A_315_297#_c_306_n 0.0513974f $X=1.25 $Y=1.95 $X2=0
+ $Y2=0
cc_185 N_VPWR_c_258_n N_A_315_297#_c_306_n 0.0201136f $X=2.2 $Y=2.29 $X2=0 $Y2=0
cc_186 N_VPWR_c_261_n N_A_315_297#_c_306_n 0.0223771f $X=2.115 $Y=2.72 $X2=0
+ $Y2=0
cc_187 N_VPWR_c_256_n N_A_315_297#_c_306_n 0.0140558f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_188 N_VPWR_c_258_n N_A_315_297#_c_301_n 0.0269205f $X=2.2 $Y=2.29 $X2=0 $Y2=0
cc_189 N_VPWR_c_263_n N_A_315_297#_c_301_n 0.0265761f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_190 N_VPWR_c_256_n N_A_315_297#_c_301_n 0.0153277f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_191 N_VPWR_c_256_n N_X_M1001_d 0.00994238f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_192 N_VPWR_c_263_n X 0.0224293f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_193 N_VPWR_c_256_n X 0.0122467f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_194 N_X_c_324_n N_VGND_c_353_n 0.0184437f $X=3 $Y=1.365 $X2=0 $Y2=0
cc_195 X N_VGND_c_353_n 0.0124789f $X=3.405 $Y=1.53 $X2=0 $Y2=0
cc_196 N_X_c_328_n N_VGND_c_355_n 0.0518793f $X=2.915 $Y=0.4 $X2=0 $Y2=0
cc_197 N_X_M1008_d N_VGND_c_357_n 0.00696094f $X=2.065 $Y=0.235 $X2=0 $Y2=0
cc_198 N_X_c_328_n N_VGND_c_357_n 0.0419897f $X=2.915 $Y=0.4 $X2=0 $Y2=0
cc_199 N_VGND_c_357_n A_317_47# 0.00381757f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
