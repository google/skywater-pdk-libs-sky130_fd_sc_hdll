* NGSPICE file created from sky130_fd_sc_hdll__or3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__or3_1 A B C VGND VNB VPB VPWR X
M1000 X a_29_53# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=4.95e+11p pd=2.99e+06u as=3.107e+11p ps=2.72e+06u
M1001 VGND C a_29_53# VNB nshort w=420000u l=150000u
+  ad=3.4965e+11p pd=3.46e+06u as=2.856e+11p ps=3.04e+06u
M1002 a_119_297# C a_29_53# VPB phighvt w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=1.134e+11p ps=1.38e+06u
M1003 VPWR A a_203_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.428e+11p ps=1.52e+06u
M1004 X a_29_53# VGND VNB nshort w=650000u l=150000u
+  ad=3.1525e+11p pd=2.27e+06u as=0p ps=0u
M1005 VGND A a_29_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_203_297# B a_119_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_29_53# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

