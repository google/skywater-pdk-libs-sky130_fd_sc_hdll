* File: sky130_fd_sc_hdll__clkinv_12.pex.spice
* Created: Thu Aug 27 19:02:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKINV_12%A 1 3 4 6 7 9 10 12 15 19 21 23 24 26 29
+ 33 35 37 38 40 43 47 49 51 52 54 57 61 63 65 66 68 71 75 77 79 80 82 85 89 91
+ 93 94 96 97 99 100 102 103 138 139
r263 139 140 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=8.015 $Y=1.202
+ $X2=8.485 $Y2=1.202
r264 137 139 33.4905 $w=3.67e-07 $l=2.55e-07 $layer=POLY_cond $X=7.76 $Y=1.202
+ $X2=8.015 $Y2=1.202
r265 137 138 13.2073 $w=1.7e-07 $l=1.87e-06 $layer=licon1_POLY $count=11 $X=7.76
+ $Y=1.16 $X2=7.76 $Y2=1.16
r266 135 137 28.2371 $w=3.67e-07 $l=2.15e-07 $layer=POLY_cond $X=7.545 $Y=1.202
+ $X2=7.76 $Y2=1.202
r267 134 135 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=7.075 $Y=1.202
+ $X2=7.545 $Y2=1.202
r268 133 134 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=7.05 $Y=1.202
+ $X2=7.075 $Y2=1.202
r269 132 133 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=6.63 $Y=1.202
+ $X2=7.05 $Y2=1.202
r270 131 132 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=6.605 $Y=1.202
+ $X2=6.63 $Y2=1.202
r271 130 131 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=6.135 $Y=1.202
+ $X2=6.605 $Y2=1.202
r272 129 130 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=6.11 $Y=1.202
+ $X2=6.135 $Y2=1.202
r273 128 129 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=5.69 $Y=1.202
+ $X2=6.11 $Y2=1.202
r274 127 128 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=5.665 $Y=1.202
+ $X2=5.69 $Y2=1.202
r275 126 127 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=5.195 $Y=1.202
+ $X2=5.665 $Y2=1.202
r276 125 126 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=5.17 $Y=1.202
+ $X2=5.195 $Y2=1.202
r277 124 125 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=4.75 $Y=1.202
+ $X2=5.17 $Y2=1.202
r278 123 124 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=4.725 $Y=1.202
+ $X2=4.75 $Y2=1.202
r279 122 123 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=4.255 $Y=1.202
+ $X2=4.725 $Y2=1.202
r280 121 122 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=4.23 $Y=1.202
+ $X2=4.255 $Y2=1.202
r281 120 121 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=3.81 $Y=1.202
+ $X2=4.23 $Y2=1.202
r282 119 120 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=3.785 $Y=1.202
+ $X2=3.81 $Y2=1.202
r283 118 119 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=3.315 $Y=1.202
+ $X2=3.785 $Y2=1.202
r284 117 118 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.202
+ $X2=3.315 $Y2=1.202
r285 116 117 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=2.87 $Y=1.202
+ $X2=3.29 $Y2=1.202
r286 115 116 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=2.87 $Y2=1.202
r287 114 115 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.845 $Y2=1.202
r288 113 114 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.202
+ $X2=2.375 $Y2=1.202
r289 112 113 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=1.93 $Y=1.202
+ $X2=2.35 $Y2=1.202
r290 111 112 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=1.93 $Y2=1.202
r291 110 111 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.905 $Y2=1.202
r292 109 110 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=1.435 $Y2=1.202
r293 107 109 45.3106 $w=3.67e-07 $l=3.45e-07 $layer=POLY_cond $X=0.62 $Y=1.202
+ $X2=0.965 $Y2=1.202
r294 107 108 13.2073 $w=1.7e-07 $l=1.87e-06 $layer=licon1_POLY $count=11 $X=0.62
+ $Y=1.16 $X2=0.62 $Y2=1.16
r295 105 107 16.4169 $w=3.67e-07 $l=1.25e-07 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.62 $Y2=1.202
r296 103 138 153.207 $w=2.53e-07 $l=3.39e-06 $layer=LI1_cond $X=4.37 $Y=1.162
+ $X2=7.76 $Y2=1.162
r297 103 108 169.477 $w=2.53e-07 $l=3.75e-06 $layer=LI1_cond $X=4.37 $Y=1.162
+ $X2=0.62 $Y2=1.162
r298 100 140 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.485 $Y=1.41
+ $X2=8.485 $Y2=1.202
r299 100 102 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.485 $Y=1.41
+ $X2=8.485 $Y2=1.985
r300 97 139 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.015 $Y=1.41
+ $X2=8.015 $Y2=1.202
r301 97 99 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.015 $Y=1.41
+ $X2=8.015 $Y2=1.985
r302 94 135 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.202
r303 94 96 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.985
r304 91 134 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.202
r305 91 93 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.985
r306 87 133 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.05 $Y=0.995
+ $X2=7.05 $Y2=1.202
r307 87 89 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.05 $Y=0.995
+ $X2=7.05 $Y2=0.445
r308 83 132 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=1.202
r309 83 85 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=0.445
r310 80 131 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.202
r311 80 82 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.985
r312 77 130 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.202
r313 77 79 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.985
r314 73 129 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.11 $Y=0.995
+ $X2=6.11 $Y2=1.202
r315 73 75 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.11 $Y=0.995
+ $X2=6.11 $Y2=0.445
r316 69 128 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=1.202
r317 69 71 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=0.445
r318 66 127 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.202
r319 66 68 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.985
r320 63 126 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.202
r321 63 65 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.985
r322 59 125 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.17 $Y=0.995
+ $X2=5.17 $Y2=1.202
r323 59 61 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.17 $Y=0.995
+ $X2=5.17 $Y2=0.445
r324 55 124 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.75 $Y=0.995
+ $X2=4.75 $Y2=1.202
r325 55 57 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.75 $Y=0.995
+ $X2=4.75 $Y2=0.445
r326 52 123 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.202
r327 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.985
r328 49 122 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.202
r329 49 51 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.985
r330 45 121 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.23 $Y=0.995
+ $X2=4.23 $Y2=1.202
r331 45 47 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.23 $Y=0.995
+ $X2=4.23 $Y2=0.445
r332 41 120 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=1.202
r333 41 43 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=0.445
r334 38 119 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.202
r335 38 40 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r336 35 118 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.202
r337 35 37 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r338 31 117 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=1.202
r339 31 33 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=0.445
r340 27 116 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.87 $Y=0.995
+ $X2=2.87 $Y2=1.202
r341 27 29 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.87 $Y=0.995
+ $X2=2.87 $Y2=0.445
r342 24 115 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r343 24 26 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r344 21 114 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r345 21 23 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r346 17 113 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.202
r347 17 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=0.445
r348 13 112 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r349 13 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.445
r350 10 111 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r351 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r352 7 110 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r353 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r354 4 109 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r355 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r356 1 105 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r357 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_12%VPWR 1 2 3 4 5 6 7 8 9 10 31 33 37 41 43
+ 47 49 53 55 59 61 65 69 73 77 80 81 83 84 86 87 88 90 95 111 112 118 121 124
+ 127 130 133
r153 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r154 131 134 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r155 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r156 128 131 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r157 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r158 125 128 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r159 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r160 122 125 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r161 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r162 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r163 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r164 109 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.97 $Y2=2.72
r165 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r166 106 109 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r167 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r168 103 106 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r169 103 134 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=5.75 $Y2=2.72
r170 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r171 100 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.065 $Y=2.72
+ $X2=5.9 $Y2=2.72
r172 100 102 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=6.065 $Y=2.72
+ $X2=6.67 $Y2=2.72
r173 99 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r174 99 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r175 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r176 96 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.2 $Y2=2.72
r177 96 98 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.61 $Y2=2.72
r178 95 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=2.72
+ $X2=2.14 $Y2=2.72
r179 95 98 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.975 $Y=2.72
+ $X2=1.61 $Y2=2.72
r180 94 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r181 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r182 91 115 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r183 91 93 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r184 90 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=1.2 $Y2=2.72
r185 90 93 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=0.69 $Y2=2.72
r186 88 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r187 88 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r188 86 108 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=8.555 $Y=2.72
+ $X2=8.51 $Y2=2.72
r189 86 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.555 $Y=2.72
+ $X2=8.72 $Y2=2.72
r190 85 111 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=2.72
+ $X2=8.97 $Y2=2.72
r191 85 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.885 $Y=2.72
+ $X2=8.72 $Y2=2.72
r192 83 105 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=7.615 $Y=2.72
+ $X2=7.59 $Y2=2.72
r193 83 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.615 $Y=2.72
+ $X2=7.78 $Y2=2.72
r194 82 108 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=7.945 $Y=2.72
+ $X2=8.51 $Y2=2.72
r195 82 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.945 $Y=2.72
+ $X2=7.78 $Y2=2.72
r196 80 102 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.675 $Y=2.72
+ $X2=6.67 $Y2=2.72
r197 80 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=2.72
+ $X2=6.84 $Y2=2.72
r198 79 105 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=7.005 $Y=2.72
+ $X2=7.59 $Y2=2.72
r199 79 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.005 $Y=2.72
+ $X2=6.84 $Y2=2.72
r200 75 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.72 $Y=2.635
+ $X2=8.72 $Y2=2.72
r201 75 77 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=8.72 $Y=2.635
+ $X2=8.72 $Y2=1.925
r202 71 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.78 $Y=2.635
+ $X2=7.78 $Y2=2.72
r203 71 73 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=7.78 $Y=2.635
+ $X2=7.78 $Y2=1.925
r204 67 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=2.635
+ $X2=6.84 $Y2=2.72
r205 67 69 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=6.84 $Y=2.635
+ $X2=6.84 $Y2=1.925
r206 63 133 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=2.635
+ $X2=5.9 $Y2=2.72
r207 63 65 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=5.9 $Y=2.635 $X2=5.9
+ $Y2=1.925
r208 62 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=2.72
+ $X2=4.96 $Y2=2.72
r209 61 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.735 $Y=2.72
+ $X2=5.9 $Y2=2.72
r210 61 62 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.735 $Y=2.72
+ $X2=5.125 $Y2=2.72
r211 57 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=2.72
r212 57 59 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=1.925
r213 56 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=2.72
+ $X2=4.02 $Y2=2.72
r214 55 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=2.72
+ $X2=4.96 $Y2=2.72
r215 55 56 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.795 $Y=2.72
+ $X2=4.185 $Y2=2.72
r216 51 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=2.72
r217 51 53 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=1.925
r218 50 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=2.72
+ $X2=3.08 $Y2=2.72
r219 49 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=2.72
+ $X2=4.02 $Y2=2.72
r220 49 50 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.855 $Y=2.72
+ $X2=3.245 $Y2=2.72
r221 45 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2.72
r222 45 47 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=1.925
r223 44 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=2.72
+ $X2=2.14 $Y2=2.72
r224 43 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=3.08 $Y2=2.72
r225 43 44 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=2.305 $Y2=2.72
r226 39 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.72
r227 39 41 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=1.925
r228 35 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.72
r229 35 37 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=1.925
r230 31 115 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r231 31 33 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=1.925
r232 10 77 300 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_PDIFF $count=2 $X=8.575
+ $Y=1.485 $X2=8.72 $Y2=1.925
r233 9 73 300 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_PDIFF $count=2 $X=7.635
+ $Y=1.485 $X2=7.78 $Y2=1.925
r234 8 69 300 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_PDIFF $count=2 $X=6.695
+ $Y=1.485 $X2=6.84 $Y2=1.925
r235 7 65 300 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_PDIFF $count=2 $X=5.755
+ $Y=1.485 $X2=5.9 $Y2=1.925
r236 6 59 300 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=1.925
r237 5 53 300 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=1.925
r238 4 47 300 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=1.925
r239 3 41 300 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.925
r240 2 37 300 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.925
r241 1 33 300 $w=1.7e-07 $l=4.98598e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.925
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_12%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 47
+ 48 49 50 51 54 56 60 62 66 68 72 74 78 80 84 86 90 92 96 98 102 104 108 110
+ 114 116 120 122 126 128 132 134 138 141 143 144 146 147 149 150 152 153 155
+ 156 158 159 161 165 166
r263 163 166 5.81876 $w=5.53e-07 $l=2.7e-07 $layer=LI1_cond $X=8.377 $Y=1.46
+ $X2=8.377 $Y2=1.19
r264 163 165 2.35019 $w=4.12e-07 $l=8.5e-08 $layer=LI1_cond $X=8.377 $Y=1.46
+ $X2=8.377 $Y2=1.545
r265 162 166 7.00406 $w=5.53e-07 $l=3.25e-07 $layer=LI1_cond $X=8.377 $Y=0.865
+ $X2=8.377 $Y2=1.19
r266 136 165 2.35019 $w=4.12e-07 $l=1.64085e-07 $layer=LI1_cond $X=8.25 $Y=1.63
+ $X2=8.377 $Y2=1.545
r267 136 138 28.5977 $w=2.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.25 $Y=1.63
+ $X2=8.25 $Y2=2.3
r268 135 161 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.445 $Y=1.545
+ $X2=7.31 $Y2=1.545
r269 134 165 4.66114 $w=1.7e-07 $l=2.77e-07 $layer=LI1_cond $X=8.1 $Y=1.545
+ $X2=8.377 $Y2=1.545
r270 134 135 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=8.1 $Y=1.545
+ $X2=7.445 $Y2=1.545
r271 130 161 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.31 $Y=1.63
+ $X2=7.31 $Y2=1.545
r272 130 132 28.5977 $w=2.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.31 $Y=1.63
+ $X2=7.31 $Y2=2.3
r273 129 159 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.975 $Y=0.78
+ $X2=6.84 $Y2=0.78
r274 128 162 9.6854 $w=1.7e-07 $l=3.16661e-07 $layer=LI1_cond $X=8.1 $Y=0.78
+ $X2=8.377 $Y2=0.865
r275 128 129 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=8.1 $Y=0.78
+ $X2=6.975 $Y2=0.78
r276 124 159 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=0.695
+ $X2=6.84 $Y2=0.78
r277 124 126 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.84 $Y=0.695
+ $X2=6.84 $Y2=0.445
r278 123 158 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.505 $Y=1.545
+ $X2=6.37 $Y2=1.545
r279 122 161 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.175 $Y=1.545
+ $X2=7.31 $Y2=1.545
r280 122 123 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.175 $Y=1.545
+ $X2=6.505 $Y2=1.545
r281 118 158 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.37 $Y=1.63
+ $X2=6.37 $Y2=1.545
r282 118 120 28.5977 $w=2.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.37 $Y=1.63
+ $X2=6.37 $Y2=2.3
r283 117 156 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.035 $Y=0.78
+ $X2=5.9 $Y2=0.78
r284 116 159 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.705 $Y=0.78
+ $X2=6.84 $Y2=0.78
r285 116 117 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.705 $Y=0.78
+ $X2=6.035 $Y2=0.78
r286 112 156 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=0.695
+ $X2=5.9 $Y2=0.78
r287 112 114 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.9 $Y=0.695
+ $X2=5.9 $Y2=0.445
r288 111 155 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.565 $Y=1.545
+ $X2=5.43 $Y2=1.545
r289 110 158 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.235 $Y=1.545
+ $X2=6.37 $Y2=1.545
r290 110 111 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.235 $Y=1.545
+ $X2=5.565 $Y2=1.545
r291 106 155 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.43 $Y=1.63
+ $X2=5.43 $Y2=1.545
r292 106 108 28.5977 $w=2.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.43 $Y=1.63
+ $X2=5.43 $Y2=2.3
r293 105 153 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.095 $Y=0.78
+ $X2=4.96 $Y2=0.78
r294 104 156 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.765 $Y=0.78
+ $X2=5.9 $Y2=0.78
r295 104 105 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.765 $Y=0.78
+ $X2=5.095 $Y2=0.78
r296 100 153 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=0.695
+ $X2=4.96 $Y2=0.78
r297 100 102 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.96 $Y=0.695
+ $X2=4.96 $Y2=0.445
r298 99 152 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.625 $Y=1.545
+ $X2=4.49 $Y2=1.545
r299 98 155 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.295 $Y=1.545
+ $X2=5.43 $Y2=1.545
r300 98 99 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.295 $Y=1.545
+ $X2=4.625 $Y2=1.545
r301 94 152 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=1.63
+ $X2=4.49 $Y2=1.545
r302 94 96 28.5977 $w=2.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.49 $Y=1.63
+ $X2=4.49 $Y2=2.3
r303 93 150 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.155 $Y=0.78
+ $X2=4.02 $Y2=0.78
r304 92 153 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.825 $Y=0.78
+ $X2=4.96 $Y2=0.78
r305 92 93 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.825 $Y=0.78
+ $X2=4.155 $Y2=0.78
r306 88 150 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.695
+ $X2=4.02 $Y2=0.78
r307 88 90 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.02 $Y=0.695
+ $X2=4.02 $Y2=0.445
r308 87 149 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.685 $Y=1.545
+ $X2=3.55 $Y2=1.545
r309 86 152 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.355 $Y=1.545
+ $X2=4.49 $Y2=1.545
r310 86 87 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.355 $Y=1.545
+ $X2=3.685 $Y2=1.545
r311 82 149 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=1.63
+ $X2=3.55 $Y2=1.545
r312 82 84 28.5977 $w=2.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.55 $Y=1.63
+ $X2=3.55 $Y2=2.3
r313 81 147 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.215 $Y=0.78
+ $X2=3.08 $Y2=0.78
r314 80 150 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.885 $Y=0.78
+ $X2=4.02 $Y2=0.78
r315 80 81 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.885 $Y=0.78
+ $X2=3.215 $Y2=0.78
r316 76 147 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.695
+ $X2=3.08 $Y2=0.78
r317 76 78 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.08 $Y=0.695
+ $X2=3.08 $Y2=0.445
r318 75 146 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.745 $Y=1.545
+ $X2=2.61 $Y2=1.545
r319 74 149 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.415 $Y=1.545
+ $X2=3.55 $Y2=1.545
r320 74 75 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.415 $Y=1.545
+ $X2=2.745 $Y2=1.545
r321 70 146 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=1.63
+ $X2=2.61 $Y2=1.545
r322 70 72 28.5977 $w=2.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.61 $Y=1.63
+ $X2=2.61 $Y2=2.3
r323 69 144 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.275 $Y=0.78
+ $X2=2.14 $Y2=0.78
r324 68 147 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.945 $Y=0.78
+ $X2=3.08 $Y2=0.78
r325 68 69 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.945 $Y=0.78
+ $X2=2.275 $Y2=0.78
r326 64 144 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.695
+ $X2=2.14 $Y2=0.78
r327 64 66 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.14 $Y=0.695
+ $X2=2.14 $Y2=0.445
r328 63 143 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.805 $Y=1.545
+ $X2=1.67 $Y2=1.545
r329 62 146 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.475 $Y=1.545
+ $X2=2.61 $Y2=1.545
r330 62 63 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.475 $Y=1.545
+ $X2=1.805 $Y2=1.545
r331 58 143 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=1.63
+ $X2=1.67 $Y2=1.545
r332 58 60 28.5977 $w=2.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.67 $Y=1.63
+ $X2=1.67 $Y2=2.3
r333 57 141 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.865 $Y=1.545
+ $X2=0.73 $Y2=1.545
r334 56 143 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.535 $Y=1.545
+ $X2=1.67 $Y2=1.545
r335 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.535 $Y=1.545
+ $X2=0.865 $Y2=1.545
r336 52 141 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.63
+ $X2=0.73 $Y2=1.545
r337 52 54 28.5977 $w=2.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.73 $Y=1.63
+ $X2=0.73 $Y2=2.3
r338 50 141 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.595 $Y=1.545
+ $X2=0.73 $Y2=1.545
r339 50 51 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.595 $Y=1.545
+ $X2=0.285 $Y2=1.545
r340 48 144 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.005 $Y=0.78
+ $X2=2.14 $Y2=0.78
r341 48 49 112.214 $w=1.68e-07 $l=1.72e-06 $layer=LI1_cond $X=2.005 $Y=0.78
+ $X2=0.285 $Y2=0.78
r342 47 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.2 $Y=1.46
+ $X2=0.285 $Y2=1.545
r343 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.2 $Y=0.865
+ $X2=0.285 $Y2=0.78
r344 46 47 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=0.2 $Y=0.865
+ $X2=0.2 $Y2=1.46
r345 15 165 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.105
+ $Y=1.485 $X2=8.25 $Y2=1.62
r346 15 138 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=8.105
+ $Y=1.485 $X2=8.25 $Y2=2.3
r347 14 161 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.165
+ $Y=1.485 $X2=7.31 $Y2=1.62
r348 14 132 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=7.165
+ $Y=1.485 $X2=7.31 $Y2=2.3
r349 13 158 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.225
+ $Y=1.485 $X2=6.37 $Y2=1.62
r350 13 120 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=6.225
+ $Y=1.485 $X2=6.37 $Y2=2.3
r351 12 155 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=1.62
r352 12 108 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=2.3
r353 11 152 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=1.62
r354 11 96 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=2.3
r355 10 149 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.62
r356 10 84 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2.3
r357 9 146 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.62
r358 9 72 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.3
r359 8 143 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.62
r360 8 60 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.3
r361 7 141 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.62
r362 7 54 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.3
r363 6 126 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=6.705
+ $Y=0.235 $X2=6.84 $Y2=0.445
r364 5 114 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=5.765
+ $Y=0.235 $X2=5.9 $Y2=0.445
r365 4 102 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=4.825
+ $Y=0.235 $X2=4.96 $Y2=0.445
r366 3 90 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.235 $X2=4.02 $Y2=0.445
r367 2 78 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=2.945
+ $Y=0.235 $X2=3.08 $Y2=0.445
r368 1 66 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_12%VGND 1 2 3 4 5 6 7 24 26 30 32 36 38 42
+ 44 48 50 60 75 76 81 84 86 89 92 95 98 103 106
r105 105 106 10.2213 $w=6.08e-07 $l=1.65e-07 $layer=LI1_cond $X=7.65 $Y=0.22
+ $X2=7.815 $Y2=0.22
r106 101 105 1.17647 $w=6.08e-07 $l=6e-08 $layer=LI1_cond $X=7.59 $Y=0.22
+ $X2=7.65 $Y2=0.22
r107 101 103 15.7115 $w=6.08e-07 $l=4.45e-07 $layer=LI1_cond $X=7.59 $Y=0.22
+ $X2=7.145 $Y2=0.22
r108 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r109 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r110 96 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r111 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r112 93 96 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r113 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r114 90 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r115 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r116 87 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r117 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r118 83 84 10.2213 $w=6.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.67 $Y=0.22
+ $X2=1.835 $Y2=0.22
r119 79 83 1.17647 $w=6.08e-07 $l=6e-08 $layer=LI1_cond $X=1.61 $Y=0.22 $X2=1.67
+ $Y2=0.22
r120 79 81 15.7115 $w=6.08e-07 $l=4.45e-07 $layer=LI1_cond $X=1.61 $Y=0.22
+ $X2=1.165 $Y2=0.22
r121 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r122 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r123 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=8.97
+ $Y2=0
r124 73 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=7.59 $Y2=0
r125 72 75 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.05 $Y=0 $X2=8.97
+ $Y2=0
r126 72 106 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=8.05 $Y=0
+ $X2=7.815 $Y2=0
r127 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r128 69 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=7.59 $Y2=0
r129 69 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=6.21
+ $Y2=0
r130 68 103 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=7.13 $Y=0
+ $X2=7.145 $Y2=0
r131 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r132 66 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.535 $Y=0 $X2=6.37
+ $Y2=0
r133 66 68 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=6.535 $Y=0
+ $X2=7.13 $Y2=0
r134 64 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r135 64 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r136 63 84 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.07 $Y=0
+ $X2=1.835 $Y2=0
r137 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r138 60 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.61
+ $Y2=0
r139 60 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.445 $Y=0
+ $X2=2.07 $Y2=0
r140 59 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r141 58 81 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.15 $Y=0 $X2=1.165
+ $Y2=0
r142 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r143 54 58 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r144 50 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r145 50 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r146 46 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.37 $Y=0.085
+ $X2=6.37 $Y2=0
r147 46 48 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=6.37 $Y=0.085
+ $X2=6.37 $Y2=0.4
r148 45 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.595 $Y=0 $X2=5.43
+ $Y2=0
r149 44 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.205 $Y=0 $X2=6.37
+ $Y2=0
r150 44 45 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.205 $Y=0
+ $X2=5.595 $Y2=0
r151 40 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.43 $Y=0.085
+ $X2=5.43 $Y2=0
r152 40 42 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.43 $Y=0.085
+ $X2=5.43 $Y2=0.4
r153 39 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.655 $Y=0 $X2=4.49
+ $Y2=0
r154 38 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.265 $Y=0 $X2=5.43
+ $Y2=0
r155 38 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.265 $Y=0
+ $X2=4.655 $Y2=0
r156 34 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=0.085
+ $X2=4.49 $Y2=0
r157 34 36 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.49 $Y=0.085
+ $X2=4.49 $Y2=0.4
r158 33 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.55
+ $Y2=0
r159 32 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.325 $Y=0 $X2=4.49
+ $Y2=0
r160 32 33 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.325 $Y=0
+ $X2=3.715 $Y2=0
r161 28 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0
r162 28 30 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0.4
r163 27 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.61
+ $Y2=0
r164 26 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.55
+ $Y2=0
r165 26 27 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.385 $Y=0
+ $X2=2.775 $Y2=0
r166 22 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0
r167 22 24 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0.4
r168 7 105 91 $w=1.7e-07 $l=6.01872e-07 $layer=licon1_NDIFF $count=2 $X=7.125
+ $Y=0.235 $X2=7.65 $Y2=0.4
r169 6 48 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=6.185
+ $Y=0.235 $X2=6.37 $Y2=0.4
r170 5 42 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=5.245
+ $Y=0.235 $X2=5.43 $Y2=0.4
r171 4 36 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.235 $X2=4.49 $Y2=0.4
r172 3 30 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.4
r173 2 24 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.4
r174 1 83 91 $w=1.7e-07 $l=5.41249e-07 $layer=licon1_NDIFF $count=2 $X=1.205
+ $Y=0.235 $X2=1.67 $Y2=0.4
.ends

