# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__xnor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xnor3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.58000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.075000 1.075000 9.535000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.735900 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.155000 0.995000 8.375000 1.445000 ;
        RECT 8.155000 1.445000 8.785000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.425400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.245000 1.075000 3.860000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 0.375000 0.925000 0.995000 ;
        RECT 0.625000 0.995000 1.860000 1.325000 ;
        RECT 0.625000 1.325000 1.005000 2.425000 ;
        RECT 1.565000 0.350000 1.875000 0.925000 ;
        RECT 1.565000 0.925000 1.860000 0.995000 ;
        RECT 1.565000 1.325000 1.860000 1.440000 ;
        RECT 1.565000 1.440000 1.895000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.770000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.580000 0.085000 ;
      RECT  0.000000  2.635000 10.580000 2.805000 ;
      RECT  0.285000  0.085000  0.455000 0.735000 ;
      RECT  0.285000  1.490000  0.455000 2.635000 ;
      RECT  1.225000  0.085000  1.395000 0.735000 ;
      RECT  1.225000  1.495000  1.395000 2.635000 ;
      RECT  2.030000  0.995000  2.285000 1.325000 ;
      RECT  2.045000  0.085000  2.345000 0.525000 ;
      RECT  2.060000  0.695000  2.735000 0.865000 ;
      RECT  2.060000  0.865000  2.285000 0.995000 ;
      RECT  2.065000  1.325000  2.285000 1.875000 ;
      RECT  2.065000  1.875000  2.850000 2.045000 ;
      RECT  2.065000  2.215000  2.450000 2.635000 ;
      RECT  2.515000  0.255000  4.185000 0.425000 ;
      RECT  2.515000  0.425000  2.735000 0.695000 ;
      RECT  2.515000  1.535000  4.200000 1.705000 ;
      RECT  2.630000  2.045000  2.850000 2.235000 ;
      RECT  2.630000  2.235000  4.200000 2.405000 ;
      RECT  2.905000  0.595000  3.075000 1.535000 ;
      RECT  3.190000  1.895000  5.890000 2.065000 ;
      RECT  3.375000  0.625000  4.695000 0.795000 ;
      RECT  3.375000  0.795000  3.755000 0.905000 ;
      RECT  3.700000  0.425000  4.185000 0.455000 ;
      RECT  4.030000  0.995000  4.355000 1.325000 ;
      RECT  4.030000  1.325000  4.200000 1.535000 ;
      RECT  4.405000  0.285000  5.035000 0.455000 ;
      RECT  4.420000  1.525000  4.805000 1.695000 ;
      RECT  4.525000  0.795000  4.695000 1.375000 ;
      RECT  4.525000  1.375000  4.805000 1.525000 ;
      RECT  4.865000  0.455000  5.035000 1.035000 ;
      RECT  4.865000  1.035000  5.145000 1.205000 ;
      RECT  4.955000  2.235000  5.285000 2.635000 ;
      RECT  4.975000  1.205000  5.145000 1.895000 ;
      RECT  5.205000  0.085000  5.375000 0.865000 ;
      RECT  5.375000  1.445000  5.895000 1.715000 ;
      RECT  5.605000  0.415000  5.895000 1.445000 ;
      RECT  5.720000  2.065000  5.890000 2.275000 ;
      RECT  5.720000  2.275000  9.015000 2.445000 ;
      RECT  6.075000  0.265000  6.520000 0.485000 ;
      RECT  6.075000  0.485000  6.245000 2.105000 ;
      RECT  6.415000  0.655000  6.875000 0.825000 ;
      RECT  6.415000  0.825000  6.585000 2.275000 ;
      RECT  6.705000  0.320000  6.875000 0.655000 ;
      RECT  6.815000  1.445000  7.645000 1.615000 ;
      RECT  6.815000  1.615000  7.230000 2.045000 ;
      RECT  6.830000  0.995000  7.255000 1.270000 ;
      RECT  7.045000  0.630000  7.255000 0.995000 ;
      RECT  7.475000  0.255000  8.670000 0.425000 ;
      RECT  7.475000  0.425000  7.645000 1.445000 ;
      RECT  7.815000  0.595000  7.985000 1.935000 ;
      RECT  7.815000  1.935000 10.325000 2.105000 ;
      RECT  8.155000  0.425000  8.670000 0.465000 ;
      RECT  8.545000  0.730000  8.750000 0.945000 ;
      RECT  8.545000  0.945000  8.855000 1.275000 ;
      RECT  9.005000  1.495000  9.875000 1.705000 ;
      RECT  9.045000  0.295000  9.335000 0.735000 ;
      RECT  9.045000  0.735000  9.875000 0.750000 ;
      RECT  9.085000  0.750000  9.875000 0.905000 ;
      RECT  9.425000  2.275000  9.810000 2.635000 ;
      RECT  9.555000  0.085000  9.725000 0.565000 ;
      RECT  9.705000  0.905000  9.875000 0.995000 ;
      RECT  9.705000  0.995000  9.985000 1.325000 ;
      RECT  9.705000  1.325000  9.875000 1.495000 ;
      RECT  9.790000  1.875000 10.325000 1.935000 ;
      RECT 10.025000  0.255000 10.325000 0.585000 ;
      RECT 10.030000  2.105000 10.325000 2.465000 ;
      RECT 10.155000  0.585000 10.325000 1.875000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.635000  1.445000  4.805000 1.615000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.605000  0.765000  5.775000 0.935000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.075000  0.425000  6.245000 0.595000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.085000  0.765000  7.255000 0.935000 ;
      RECT  7.085000  1.445000  7.255000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.565000  0.765000  8.735000 0.935000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.075000  0.425000  9.245000 0.595000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
    LAYER met1 ;
      RECT 4.575000 1.415000 4.865000 1.460000 ;
      RECT 4.575000 1.460000 7.315000 1.600000 ;
      RECT 4.575000 1.600000 4.865000 1.645000 ;
      RECT 5.545000 0.735000 5.835000 0.780000 ;
      RECT 5.545000 0.780000 8.795000 0.920000 ;
      RECT 5.545000 0.920000 5.835000 0.965000 ;
      RECT 6.015000 0.395000 6.315000 0.440000 ;
      RECT 6.015000 0.440000 9.305000 0.580000 ;
      RECT 6.015000 0.580000 6.315000 0.625000 ;
      RECT 7.025000 0.735000 7.315000 0.780000 ;
      RECT 7.025000 0.920000 7.315000 0.965000 ;
      RECT 7.025000 1.415000 7.315000 1.460000 ;
      RECT 7.025000 1.600000 7.315000 1.645000 ;
      RECT 8.505000 0.735000 8.795000 0.780000 ;
      RECT 8.505000 0.920000 8.795000 0.965000 ;
      RECT 9.015000 0.395000 9.305000 0.440000 ;
      RECT 9.015000 0.580000 9.305000 0.625000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xnor3_4
END LIBRARY
