* File: sky130_fd_sc_hdll__and4b_1.spice
* Created: Wed Sep  2 08:23:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and4b_1.pex.spice"
.subckt sky130_fd_sc_hdll__and4b_1  VNB VPB A_N B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_N_M1008_g N_A_27_47#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1302 PD=1.36 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 A_307_47# N_A_27_47#_M1011_g N_A_213_413#_M1011_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1000 A_379_47# N_B_M1000_g A_307_47# VNB NSHORT L=0.15 W=0.42 AD=0.105
+ AS=0.0441 PD=0.92 PS=0.63 NRD=55.704 NRS=14.28 M=1 R=2.8 SA=75000.5 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1002 A_509_47# N_C_M1002_g A_379_47# VNB NSHORT L=0.15 W=0.42 AD=0.07455
+ AS=0.105 PD=0.775 PS=0.92 NRD=34.992 NRS=55.704 M=1 R=2.8 SA=75001.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_D_M1005_g A_509_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0914579 AS=0.07455 PD=0.812523 PS=0.775 NRD=0 NRS=34.992 M=1 R=2.8
+ SA=75001.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_X_M1003_d N_A_213_413#_M1003_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.141542 PD=1.82 PS=1.25748 NRD=0 NRS=20.304 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_A_N_M1001_g N_A_27_47#_M1001_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.063 AS=0.1134 PD=0.72 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90003.2 A=0.0756 P=1.2 MULT=1
MM1006 N_A_213_413#_M1006_d N_A_27_47#_M1006_g N_VPWR_M1001_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0903 AS=0.063 PD=0.85 PS=0.72 NRD=37.5088 NRS=7.0329 M=1 R=2.33333
+ SA=90000.7 SB=90002.7 A=0.0756 P=1.2 MULT=1
MM1004 N_VPWR_M1004_d N_B_M1004_g N_A_213_413#_M1006_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.1428 AS=0.0903 PD=1.1 PS=0.85 NRD=2.3443 NRS=32.8202 M=1 R=2.33333
+ SA=90001.3 SB=90002.1 A=0.0756 P=1.2 MULT=1
MM1009 N_A_213_413#_M1009_d N_C_M1009_g N_VPWR_M1004_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.06825 AS=0.1428 PD=0.745 PS=1.1 NRD=18.7544 NRS=2.3443 M=1 R=2.33333
+ SA=90002.1 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_D_M1010_g N_A_213_413#_M1009_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0887028 AS=0.06825 PD=0.801549 PS=0.745 NRD=21.0987 NRS=2.3443 M=1
+ R=2.33333 SA=90002.6 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1007 N_X_M1007_d N_A_213_413#_M1007_g N_VPWR_M1010_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.211197 PD=2.54 PS=1.90845 NRD=0.9653 NRS=5.8903 M=1 R=5.55556
+ SA=90001.4 SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hdll__and4b_1.pxi.spice"
*
.ends
*
*
