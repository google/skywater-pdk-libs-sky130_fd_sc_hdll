* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nand2_16 A B VGND VNB VPB VPWR Y
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X26 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X31 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X34 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X36 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X37 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X38 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X40 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X41 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X42 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X43 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X44 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X45 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X46 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X47 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X48 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X49 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X50 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X51 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X52 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X53 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X54 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X55 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X56 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X57 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X58 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X59 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X60 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X61 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X62 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X63 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
