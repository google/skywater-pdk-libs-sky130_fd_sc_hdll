* File: sky130_fd_sc_hdll__nand4b_1.pex.spice
* Created: Wed Sep  2 08:38:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND4B_1%A_N 1 3 4 6 7 15
r27 11 15 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.51 $Y=1.16
+ $X2=0.685 $Y2=1.16
r28 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r29 7 15 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.69 $Y=1.16 $X2=0.685
+ $Y2=1.16
r30 4 10 45.964 $w=3.43e-07 $l=2.91548e-07 $layer=POLY_cond $X=0.62 $Y=1.41
+ $X2=0.53 $Y2=1.16
r31 4 6 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.62 $Y=1.41 $X2=0.62
+ $Y2=1.695
r32 1 10 38.7084 $w=3.43e-07 $l=1.92678e-07 $layer=POLY_cond $X=0.59 $Y=0.995
+ $X2=0.53 $Y2=1.16
r33 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.59 $Y=0.995 $X2=0.59
+ $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_1%D 1 3 4 6 7 14
r31 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.095
+ $Y=1.16 $X2=1.095 $Y2=1.16
r32 7 14 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=1.15 $Y=1.16
+ $X2=1.095 $Y2=1.16
r33 4 10 38.7084 $w=3.43e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.18 $Y=0.995
+ $X2=1.12 $Y2=1.16
r34 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.18 $Y=0.995 $X2=1.18
+ $Y2=0.56
r35 1 10 45.964 $w=3.43e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.155 $Y=1.41
+ $X2=1.12 $Y2=1.16
r36 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.155 $Y=1.41
+ $X2=1.155 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_1%C 1 3 4 6 7 13
c35 7 0 2.79153e-20 $X=1.525 $Y=1.105
r36 7 13 0.115094 $w=5.3e-07 $l=5e-09 $layer=LI1_cond $X=1.61 $Y=1.045 $X2=1.605
+ $Y2=1.045
r37 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.655
+ $Y=1.16 $X2=1.655 $Y2=1.16
r38 4 10 51.486 $w=2.55e-07 $l=2.64575e-07 $layer=POLY_cond $X=1.625 $Y=1.41
+ $X2=1.655 $Y2=1.16
r39 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.625 $Y=1.41
+ $X2=1.625 $Y2=1.985
r40 1 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.595 $Y=0.995
+ $X2=1.655 $Y2=1.16
r41 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.595 $Y=0.995
+ $X2=1.595 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_1%B 1 3 4 6 7 13
c36 7 0 2.75894e-20 $X=1.985 $Y=1.105
r37 7 13 0.106793 $w=5.58e-07 $l=5e-09 $layer=LI1_cond $X=2.07 $Y=1.045
+ $X2=2.065 $Y2=1.045
r38 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.16 $X2=2.14 $Y2=1.16
r39 4 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.105 $Y=1.41
+ $X2=2.14 $Y2=1.16
r40 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.105 $Y=1.41
+ $X2=2.105 $Y2=1.985
r41 1 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.08 $Y=0.995
+ $X2=2.14 $Y2=1.16
r42 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.08 $Y=0.995 $X2=2.08
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_1%A_40_93# 1 2 7 9 10 12 14 15 17 20 25 29
+ 31 38
c81 20 0 2.79153e-20 $X=2.497 $Y=0.995
r82 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.62
+ $Y=1.16 $X2=2.62 $Y2=1.16
r83 35 38 4.29547 $w=3.28e-07 $l=1.23e-07 $layer=LI1_cond $X=2.497 $Y=1.16
+ $X2=2.62 $Y2=1.16
r84 31 33 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.285 $Y=0.51
+ $X2=1.285 $Y2=0.74
r85 26 29 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=0.17 $Y=1.76
+ $X2=0.385 $Y2=1.76
r86 24 25 7.96465 $w=3.78e-07 $l=1.45e-07 $layer=LI1_cond $X=0.325 $Y=0.635
+ $X2=0.47 $Y2=0.635
r87 21 24 4.70075 $w=3.78e-07 $l=1.55e-07 $layer=LI1_cond $X=0.17 $Y=0.635
+ $X2=0.325 $Y2=0.635
r88 20 35 3.54104 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=2.497 $Y=0.995
+ $X2=2.497 $Y2=1.16
r89 19 20 21.6408 $w=2.03e-07 $l=4e-07 $layer=LI1_cond $X=2.497 $Y=0.595
+ $X2=2.497 $Y2=0.995
r90 18 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=0.51
+ $X2=1.285 $Y2=0.51
r91 17 19 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=2.395 $Y=0.51
+ $X2=2.497 $Y2=0.595
r92 17 18 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=2.395 $Y=0.51
+ $X2=1.37 $Y2=0.51
r93 15 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.74
+ $X2=1.285 $Y2=0.74
r94 15 25 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.2 $Y=0.74 $X2=0.47
+ $Y2=0.74
r95 14 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=1.595
+ $X2=0.17 $Y2=1.76
r96 13 21 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=0.635
r97 13 14 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=1.595
r98 10 39 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.585 $Y=1.41
+ $X2=2.62 $Y2=1.16
r99 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.585 $Y=1.41
+ $X2=2.585 $Y2=1.985
r100 7 39 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.56 $Y=0.995
+ $X2=2.62 $Y2=1.16
r101 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.56 $Y=0.995
+ $X2=2.56 $Y2=0.56
r102 2 29 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.26
+ $Y=1.485 $X2=0.385 $Y2=1.76
r103 1 24 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.2
+ $Y=0.465 $X2=0.325 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_1%VPWR 1 2 3 12 18 20 22 25 26 28 29 30 39
+ 45
r44 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 42 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r46 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r47 39 44 3.70618 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.875 $Y=2.72
+ $X2=3.047 $Y2=2.72
r48 39 41 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.875 $Y=2.72
+ $X2=2.53 $Y2=2.72
r49 38 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r50 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r51 34 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r52 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r53 30 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r54 28 37 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.725 $Y=2.72
+ $X2=1.61 $Y2=2.72
r55 28 29 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=1.725 $Y=2.72
+ $X2=1.862 $Y2=2.72
r56 27 41 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2 $Y=2.72 $X2=2.53
+ $Y2=2.72
r57 27 29 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=2 $Y=2.72 $X2=1.862
+ $Y2=2.72
r58 25 33 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.755 $Y=2.72
+ $X2=0.69 $Y2=2.72
r59 25 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.755 $Y=2.72
+ $X2=0.88 $Y2=2.72
r60 24 37 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.005 $Y=2.72
+ $X2=1.61 $Y2=2.72
r61 24 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.005 $Y=2.72
+ $X2=0.88 $Y2=2.72
r62 20 44 3.23214 $w=2.15e-07 $l=1.12916e-07 $layer=LI1_cond $X=2.982 $Y=2.635
+ $X2=3.047 $Y2=2.72
r63 20 22 34.0373 $w=2.13e-07 $l=6.35e-07 $layer=LI1_cond $X=2.982 $Y=2.635
+ $X2=2.982 $Y2=2
r64 16 29 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.862 $Y=2.635
+ $X2=1.862 $Y2=2.72
r65 16 18 26.611 $w=2.73e-07 $l=6.35e-07 $layer=LI1_cond $X=1.862 $Y=2.635
+ $X2=1.862 $Y2=2
r66 12 15 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.88 $Y=1.66
+ $X2=0.88 $Y2=2
r67 10 26 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=2.635
+ $X2=0.88 $Y2=2.72
r68 10 15 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.88 $Y=2.635
+ $X2=0.88 $Y2=2
r69 3 22 300 $w=1.7e-07 $l=6.41872e-07 $layer=licon1_PDIFF $count=2 $X=2.675
+ $Y=1.485 $X2=2.96 $Y2=2
r70 2 18 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.715
+ $Y=1.485 $X2=1.86 $Y2=2
r71 1 15 300 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=2 $X=0.71
+ $Y=1.485 $X2=0.92 $Y2=2
r72 1 12 600 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_PDIFF $count=1 $X=0.71
+ $Y=1.485 $X2=0.92 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_1%Y 1 2 3 10 12 14 18 20 23 27 29 30 33
c50 23 0 2.75894e-20 $X=3.005 $Y=1.495
r51 30 33 3.36129 $w=3.58e-07 $l=1.05e-07 $layer=LI1_cond $X=2.955 $Y=0.51
+ $X2=2.955 $Y2=0.405
r52 28 30 4.64178 $w=3.58e-07 $l=1.45e-07 $layer=LI1_cond $X=2.955 $Y=0.655
+ $X2=2.955 $Y2=0.51
r53 28 29 6.67067 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=2.955 $Y=0.655
+ $X2=2.955 $Y2=0.835
r54 23 29 29.2543 $w=2.58e-07 $l=6.6e-07 $layer=LI1_cond $X=3.005 $Y=1.495
+ $X2=3.005 $Y2=0.835
r55 21 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=1.58
+ $X2=2.34 $Y2=1.58
r56 20 23 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.875 $Y=1.58
+ $X2=3.005 $Y2=1.495
r57 20 21 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.875 $Y=1.58
+ $X2=2.505 $Y2=1.58
r58 16 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=1.665
+ $X2=2.34 $Y2=1.58
r59 16 18 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=2.34 $Y=1.665
+ $X2=2.34 $Y2=2.335
r60 15 25 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.555 $Y=1.58
+ $X2=1.365 $Y2=1.58
r61 14 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=1.58
+ $X2=2.34 $Y2=1.58
r62 14 15 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.175 $Y=1.58
+ $X2=1.555 $Y2=1.58
r63 10 25 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=1.665
+ $X2=1.365 $Y2=1.58
r64 10 12 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.365 $Y=1.665
+ $X2=1.365 $Y2=2.34
r65 3 27 400 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=2.195
+ $Y=1.485 $X2=2.34 $Y2=1.655
r66 3 18 400 $w=1.7e-07 $l=9.19647e-07 $layer=licon1_PDIFF $count=1 $X=2.195
+ $Y=1.485 $X2=2.34 $Y2=2.335
r67 2 25 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.245
+ $Y=1.485 $X2=1.39 $Y2=1.66
r68 2 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.245
+ $Y=1.485 $X2=1.39 $Y2=2.34
r69 1 33 91 $w=1.7e-07 $l=3.80624e-07 $layer=licon1_NDIFF $count=2 $X=2.635
+ $Y=0.235 $X2=2.94 $Y2=0.405
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_1%VGND 1 8 10 17 18 21
r35 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r36 17 18 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r37 15 18 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r38 15 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r39 14 17 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r40 14 15 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r41 12 21 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=0.847
+ $Y2=0
r42 12 14 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=1.15
+ $Y2=0
r43 10 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r44 6 21 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.847 $Y=0.085
+ $X2=0.847 $Y2=0
r45 6 8 9.31427 $w=3.63e-07 $l=2.95e-07 $layer=LI1_cond $X=0.847 $Y=0.085
+ $X2=0.847 $Y2=0.38
r46 1 8 182 $w=1.7e-07 $l=2.38747e-07 $layer=licon1_NDIFF $count=1 $X=0.665
+ $Y=0.465 $X2=0.865 $Y2=0.38
.ends

