* File: sky130_fd_sc_hdll__a21o_1.pex.spice
* Created: Thu Aug 27 18:52:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A21O_1%A_81_21# 1 2 7 9 10 12 16 18 19 20 22 24 32
c56 18 0 1.18052e-19 $X=1.515 $Y=0.735
r57 31 32 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.48 $Y=1.202
+ $X2=0.505 $Y2=1.202
r58 24 26 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=0.635
+ $X2=1.665 $Y2=0.55
r59 20 22 3.62806 $w=2.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=1.725
+ $X2=1.23 $Y2=1.81
r60 18 24 7.17723 $w=2e-07 $l=1.93649e-07 $layer=LI1_cond $X=1.515 $Y=0.735
+ $X2=1.665 $Y2=0.635
r61 18 19 34.9364 $w=1.98e-07 $l=6.3e-07 $layer=LI1_cond $X=1.515 $Y=0.735
+ $X2=0.885 $Y2=0.735
r62 17 32 31.6932 $w=3.65e-07 $l=2.4e-07 $layer=POLY_cond $X=0.745 $Y=1.202
+ $X2=0.505 $Y2=1.202
r63 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.745
+ $Y=1.16 $X2=0.745 $Y2=1.16
r64 14 20 26.9776 $w=2.18e-07 $l=5.15e-07 $layer=LI1_cond $X=0.715 $Y=1.615
+ $X2=1.23 $Y2=1.615
r65 14 16 11.6939 $w=3.38e-07 $l=3.45e-07 $layer=LI1_cond $X=0.715 $Y=1.505
+ $X2=0.715 $Y2=1.16
r66 13 19 7.42997 $w=2e-07 $l=2.14243e-07 $layer=LI1_cond $X=0.715 $Y=0.835
+ $X2=0.885 $Y2=0.735
r67 13 16 11.016 $w=3.38e-07 $l=3.25e-07 $layer=LI1_cond $X=0.715 $Y=0.835
+ $X2=0.715 $Y2=1.16
r68 10 32 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.41
+ $X2=0.505 $Y2=1.202
r69 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.41
+ $X2=0.505 $Y2=1.985
r70 7 31 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.48 $Y=0.995
+ $X2=0.48 $Y2=1.202
r71 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.48 $Y=0.995 $X2=0.48
+ $Y2=0.56
r72 2 22 300 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_PDIFF $count=2 $X=1.135
+ $Y=1.485 $X2=1.26 $Y2=1.81
r73 1 26 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.73 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_1%B1 1 3 4 6 7 11 13
r29 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.445
+ $Y=1.16 $X2=1.445 $Y2=1.16
r30 7 11 9.10802 $w=3.08e-07 $l=2.45e-07 $layer=LI1_cond $X=1.2 $Y=1.17
+ $X2=1.445 $Y2=1.17
r31 7 13 1.85878 $w=3.08e-07 $l=5e-08 $layer=LI1_cond $X=1.2 $Y=1.17 $X2=1.15
+ $Y2=1.17
r32 4 10 38.9672 $w=2.67e-07 $l=1.96074e-07 $layer=POLY_cond $X=1.52 $Y=0.995
+ $X2=1.452 $Y2=1.16
r33 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.52 $Y=0.995 $X2=1.52
+ $Y2=0.56
r34 1 10 50.2707 $w=2.67e-07 $l=2.70647e-07 $layer=POLY_cond $X=1.495 $Y=1.41
+ $X2=1.452 $Y2=1.16
r35 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.495 $Y=1.41
+ $X2=1.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_1%A1 1 3 4 6 7 8 9 25
c38 1 0 1.18052e-19 $X=1.98 $Y=1.41
r39 15 25 4.64695 $w=3.08e-07 $l=1.25e-07 $layer=LI1_cond $X=1.945 $Y=1.17
+ $X2=2.07 $Y2=1.17
r40 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.945
+ $Y=1.16 $X2=1.945 $Y2=1.16
r41 9 25 1.11527 $w=3.08e-07 $l=3e-08 $layer=LI1_cond $X=2.1 $Y=1.17 $X2=2.07
+ $Y2=1.17
r42 9 16 2.48709 $w=2.3e-07 $l=1.55e-07 $layer=LI1_cond $X=2.1 $Y=1.17 $X2=2.1
+ $Y2=1.015
r43 8 16 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.1 $Y=0.85 $X2=2.1
+ $Y2=1.015
r44 7 8 17.0361 $w=2.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.1 $Y=0.51 $X2=2.1
+ $Y2=0.85
r45 4 14 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.005 $Y=0.995
+ $X2=1.945 $Y2=1.16
r46 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.005 $Y=0.995
+ $X2=2.005 $Y2=0.56
r47 1 14 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.98 $Y=1.41
+ $X2=1.945 $Y2=1.16
r48 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.98 $Y=1.41 $X2=1.98
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_1%A2 1 3 4 6 7 15
r20 7 15 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=2.495 $Y=1.16 $X2=2.545
+ $Y2=1.16
r21 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.495
+ $Y=1.16 $X2=2.495 $Y2=1.16
r22 4 10 46.8511 $w=3.19e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.46 $Y=1.41
+ $X2=2.535 $Y2=1.16
r23 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.46 $Y=1.41 $X2=2.46
+ $Y2=1.985
r24 1 10 38.5462 $w=3.19e-07 $l=2.09105e-07 $layer=POLY_cond $X=2.435 $Y=0.995
+ $X2=2.535 $Y2=1.16
r25 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.435 $Y=0.995
+ $X2=2.435 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_1%X 1 2 7 8 9 10 11 12
r13 11 12 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.225 $Y=1.87
+ $X2=0.225 $Y2=2.21
r14 11 30 4.43247 $w=2.58e-07 $l=1e-07 $layer=LI1_cond $X=0.225 $Y=1.87
+ $X2=0.225 $Y2=1.77
r15 10 30 10.6379 $w=2.58e-07 $l=2.4e-07 $layer=LI1_cond $X=0.225 $Y=1.53
+ $X2=0.225 $Y2=1.77
r16 9 10 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.225 $Y=1.19
+ $X2=0.225 $Y2=1.53
r17 8 9 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.225 $Y=0.85
+ $X2=0.225 $Y2=1.19
r18 7 8 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.225 $Y=0.51
+ $X2=0.225 $Y2=0.85
r19 2 30 300 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_PDIFF $count=2 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=1.77
r20 1 7 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.235 $X2=0.27 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_1%VPWR 1 2 9 13 15 17 22 29 30 33 36
r42 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r43 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r44 30 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r45 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r46 27 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.385 $Y=2.72
+ $X2=2.195 $Y2=2.72
r47 27 29 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.385 $Y=2.72
+ $X2=2.99 $Y2=2.72
r48 26 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r49 26 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r51 23 33 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.915 $Y=2.72
+ $X2=0.72 $Y2=2.72
r52 23 25 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.915 $Y=2.72
+ $X2=1.15 $Y2=2.72
r53 22 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=2.195 $Y2=2.72
r54 22 25 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=1.15 $Y2=2.72
r55 17 33 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.72 $Y2=2.72
r56 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.23 $Y2=2.72
r57 15 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r58 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r59 11 36 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=2.635
+ $X2=2.195 $Y2=2.72
r60 11 13 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=2.195 $Y=2.635
+ $X2=2.195 $Y2=2.02
r61 7 33 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=2.635 $X2=0.72
+ $Y2=2.72
r62 7 9 18.7641 $w=3.88e-07 $l=6.35e-07 $layer=LI1_cond $X=0.72 $Y=2.635
+ $X2=0.72 $Y2=2
r63 2 13 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=2.07
+ $Y=1.485 $X2=2.22 $Y2=2.02
r64 1 9 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.485 $X2=0.74 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_1%A_317_297# 1 2 9 11 12 15
r19 13 15 3.7676 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=1.745
+ $X2=2.735 $Y2=1.83
r20 11 13 6.83069 $w=2.4e-07 $l=1.80278e-07 $layer=LI1_cond $X=2.605 $Y=1.625
+ $X2=2.735 $Y2=1.745
r21 11 12 37.4544 $w=2.38e-07 $l=7.8e-07 $layer=LI1_cond $X=2.605 $Y=1.625
+ $X2=1.825 $Y2=1.625
r22 7 12 6.82051 $w=2.4e-07 $l=1.67929e-07 $layer=LI1_cond $X=1.71 $Y=1.745
+ $X2=1.825 $Y2=1.625
r23 7 9 4.25903 $w=2.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.745 $X2=1.71
+ $Y2=1.83
r24 2 15 300 $w=1.7e-07 $l=4.13249e-07 $layer=licon1_PDIFF $count=2 $X=2.55
+ $Y=1.485 $X2=2.7 $Y2=1.83
r25 1 9 300 $w=1.7e-07 $l=4.11157e-07 $layer=licon1_PDIFF $count=2 $X=1.585
+ $Y=1.485 $X2=1.73 $Y2=1.83
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_1%VGND 1 2 11 14 15 16 26 27 30 38
r41 37 38 9.76796 $w=5.38e-07 $l=1.65e-07 $layer=LI1_cond $X=1.17 $Y=0.185
+ $X2=1.335 $Y2=0.185
r42 34 37 0.442992 $w=5.38e-07 $l=2e-08 $layer=LI1_cond $X=1.15 $Y=0.185
+ $X2=1.17 $Y2=0.185
r43 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r44 31 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r45 30 34 10.1888 $w=5.38e-07 $l=4.6e-07 $layer=LI1_cond $X=0.69 $Y=0.185
+ $X2=1.15 $Y2=0.185
r46 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r47 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r48 24 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r49 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r50 21 24 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r51 21 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r52 20 23 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r53 20 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.335
+ $Y2=0
r54 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r55 16 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r56 14 23 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.575 $Y=0 $X2=2.53
+ $Y2=0
r57 14 15 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.575 $Y=0 $X2=2.72
+ $Y2=0
r58 13 26 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.99
+ $Y2=0
r59 13 15 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.72
+ $Y2=0
r60 9 15 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.72 $Y=0.085
+ $X2=2.72 $Y2=0
r61 9 11 17.684 $w=2.88e-07 $l=4.45e-07 $layer=LI1_cond $X=2.72 $Y=0.085
+ $X2=2.72 $Y2=0.53
r62 2 11 182 $w=1.7e-07 $l=3.78253e-07 $layer=licon1_NDIFF $count=1 $X=2.51
+ $Y=0.235 $X2=2.7 $Y2=0.53
r63 1 37 91 $w=1.7e-07 $l=6.74611e-07 $layer=licon1_NDIFF $count=2 $X=0.555
+ $Y=0.235 $X2=1.17 $Y2=0.36
.ends

