* File: sky130_fd_sc_hdll__nor3_2.pxi.spice
* Created: Wed Sep  2 08:40:21 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR3_2%A N_A_c_53_n N_A_M1005_g N_A_c_57_n N_A_M1000_g
+ N_A_c_58_n N_A_M1008_g N_A_c_54_n N_A_M1011_g A A N_A_c_56_n A
+ PM_SKY130_FD_SC_HDLL__NOR3_2%A
x_PM_SKY130_FD_SC_HDLL__NOR3_2%B N_B_c_90_n N_B_M1006_g N_B_c_94_n N_B_M1002_g
+ N_B_c_95_n N_B_M1004_g N_B_c_91_n N_B_M1010_g B B N_B_c_93_n B
+ PM_SKY130_FD_SC_HDLL__NOR3_2%B
x_PM_SKY130_FD_SC_HDLL__NOR3_2%C N_C_c_132_n N_C_M1001_g N_C_c_136_n N_C_M1003_g
+ N_C_c_137_n N_C_M1007_g N_C_c_133_n N_C_M1009_g N_C_c_156_p C C N_C_c_134_n
+ N_C_c_135_n PM_SKY130_FD_SC_HDLL__NOR3_2%C
x_PM_SKY130_FD_SC_HDLL__NOR3_2%A_27_297# N_A_27_297#_M1000_s N_A_27_297#_M1008_s
+ N_A_27_297#_M1004_d N_A_27_297#_c_175_n N_A_27_297#_c_199_p
+ N_A_27_297#_c_176_n N_A_27_297#_c_195_p N_A_27_297#_c_177_n
+ N_A_27_297#_c_178_n N_A_27_297#_c_179_n PM_SKY130_FD_SC_HDLL__NOR3_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__NOR3_2%VPWR N_VPWR_M1000_d N_VPWR_c_211_n VPWR
+ N_VPWR_c_212_n N_VPWR_c_210_n N_VPWR_c_214_n PM_SKY130_FD_SC_HDLL__NOR3_2%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR3_2%A_309_297# N_A_309_297#_M1002_s
+ N_A_309_297#_M1003_d N_A_309_297#_M1007_d N_A_309_297#_c_260_n
+ N_A_309_297#_c_250_n N_A_309_297#_c_270_n N_A_309_297#_c_253_n
+ N_A_309_297#_c_251_n N_A_309_297#_c_279_p N_A_309_297#_c_274_n
+ PM_SKY130_FD_SC_HDLL__NOR3_2%A_309_297#
x_PM_SKY130_FD_SC_HDLL__NOR3_2%Y N_Y_M1005_d N_Y_M1006_s N_Y_M1001_s N_Y_M1003_s
+ N_Y_c_288_n N_Y_c_281_n N_Y_c_282_n N_Y_c_294_n N_Y_c_283_n N_Y_c_306_n
+ N_Y_c_284_n N_Y_c_285_n Y N_Y_c_324_n Y PM_SKY130_FD_SC_HDLL__NOR3_2%Y
x_PM_SKY130_FD_SC_HDLL__NOR3_2%VGND N_VGND_M1005_s N_VGND_M1011_s N_VGND_M1010_d
+ N_VGND_M1001_d N_VGND_M1009_d N_VGND_c_350_n N_VGND_c_351_n N_VGND_c_352_n
+ N_VGND_c_353_n N_VGND_c_354_n N_VGND_c_355_n VGND N_VGND_c_356_n
+ N_VGND_c_357_n N_VGND_c_358_n N_VGND_c_359_n N_VGND_c_360_n
+ PM_SKY130_FD_SC_HDLL__NOR3_2%VGND
cc_1 VNB N_A_c_53_n 0.0222857f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_54_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_3 VNB A 0.0161137f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_4 VNB N_A_c_56_n 0.0440201f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_5 VNB N_B_c_90_n 0.0169338f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_6 VNB N_B_c_91_n 0.0224149f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_7 VNB B 0.0103571f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_8 VNB N_B_c_93_n 0.0421799f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_9 VNB N_C_c_132_n 0.0223802f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_10 VNB N_C_c_133_n 0.020726f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_11 VNB N_C_c_134_n 0.0462418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_C_c_135_n 0.00885357f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_13 VNB N_VPWR_c_210_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_14 VNB N_Y_c_281_n 0.00355899f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.202
cc_15 VNB N_Y_c_282_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_16 VNB N_Y_c_283_n 0.0187564f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.202
cc_17 VNB N_Y_c_284_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Y_c_285_n 0.0140207f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB Y 0.0200326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_350_n 0.0103581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_351_n 0.0349588f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_22 VNB N_VGND_c_352_n 0.0199314f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_23 VNB N_VGND_c_353_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.18
cc_24 VNB N_VGND_c_354_n 0.0139264f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.18
cc_25 VNB N_VGND_c_355_n 0.0187017f $X=-0.19 $Y=-0.24 $X2=0.745 $Y2=1.18
cc_26 VNB N_VGND_c_356_n 0.0193093f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_357_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_358_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_359_n 0.0318808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_360_n 0.220593f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VPB N_A_c_57_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_32 VPB N_A_c_58_n 0.0161064f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_33 VPB N_A_c_56_n 0.022695f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_34 VPB N_B_c_94_n 0.0161064f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_35 VPB N_B_c_95_n 0.0194161f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_36 VPB N_B_c_93_n 0.0204291f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_37 VPB N_C_c_136_n 0.0190998f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_38 VPB N_C_c_137_n 0.0194429f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_39 VPB N_C_c_134_n 0.0233271f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_C_c_135_n 0.0108596f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.19
cc_41 VPB N_A_27_297#_c_175_n 0.00371848f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_42 VPB N_A_27_297#_c_176_n 0.0020765f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_43 VPB N_A_27_297#_c_177_n 0.00199216f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_44 VPB N_A_27_297#_c_178_n 0.00322557f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.19
cc_45 VPB N_A_27_297#_c_179_n 0.00255575f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_211_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.985
cc_47 VPB N_VPWR_c_212_n 0.0816898f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.202
cc_48 VPB N_VPWR_c_210_n 0.0563046f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_49 VPB N_VPWR_c_214_n 0.0244347f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_50 VPB N_A_309_297#_c_250_n 0.0134708f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_51 VPB N_A_309_297#_c_251_n 0.00692367f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_52 VPB Y 0.0235511f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 N_A_c_54_n N_B_c_90_n 0.024264f $X=1.01 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_54 N_A_c_58_n N_B_c_94_n 0.00985632f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_55 A B 0.0152605f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_56 N_A_c_56_n B 0.0018186f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_57 N_A_c_56_n N_B_c_93_n 0.024264f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_58 A N_A_27_297#_c_175_n 0.021852f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_59 N_A_c_57_n N_A_27_297#_c_176_n 0.0158351f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_60 N_A_c_58_n N_A_27_297#_c_176_n 0.016363f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_61 A N_A_27_297#_c_176_n 0.0431894f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_62 N_A_c_56_n N_A_27_297#_c_176_n 0.00794509f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_63 N_A_c_57_n N_VPWR_c_211_n 0.00300743f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_64 N_A_c_58_n N_VPWR_c_211_n 0.00300743f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_65 N_A_c_58_n N_VPWR_c_212_n 0.00702461f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_66 N_A_c_57_n N_VPWR_c_210_n 0.0133387f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_67 N_A_c_58_n N_VPWR_c_210_n 0.0124344f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_68 N_A_c_57_n N_VPWR_c_214_n 0.00702461f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_69 N_A_c_53_n N_Y_c_288_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_70 N_A_c_54_n N_Y_c_281_n 0.0114598f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_71 A N_Y_c_281_n 0.00695775f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_72 N_A_c_53_n N_Y_c_282_n 0.00269085f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_73 A N_Y_c_282_n 0.030835f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A_c_56_n N_Y_c_282_n 0.00486271f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_75 N_A_c_54_n N_Y_c_294_n 5.32212e-19 $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_76 N_A_c_53_n N_VGND_c_351_n 0.00496762f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_77 A N_VGND_c_351_n 0.019624f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_78 N_A_c_53_n N_VGND_c_352_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_79 N_A_c_54_n N_VGND_c_352_n 0.00437852f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_80 N_A_c_54_n N_VGND_c_353_n 0.00268723f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A_c_53_n N_VGND_c_360_n 0.0107167f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A_c_54_n N_VGND_c_360_n 0.00615622f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_83 B N_C_c_134_n 6.28004e-19 $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_84 N_B_c_95_n N_C_c_135_n 0.00172372f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_85 B N_C_c_135_n 0.0189349f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_86 N_B_c_93_n N_C_c_135_n 0.00496642f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_87 N_B_c_94_n N_A_27_297#_c_177_n 0.0156202f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_88 N_B_c_95_n N_A_27_297#_c_177_n 0.0130803f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_89 B N_A_27_297#_c_177_n 0.0487774f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_90 N_B_c_93_n N_A_27_297#_c_177_n 0.00789593f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_91 B N_A_27_297#_c_178_n 0.00942636f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_92 B N_A_27_297#_c_179_n 0.0205419f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_93 N_B_c_94_n N_VPWR_c_212_n 0.00702461f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_94 N_B_c_95_n N_VPWR_c_212_n 0.00429453f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_95 N_B_c_94_n N_VPWR_c_210_n 0.0126324f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_96 N_B_c_95_n N_VPWR_c_210_n 0.00739666f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_97 N_B_c_95_n N_A_309_297#_c_250_n 0.0136098f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_98 N_B_c_95_n N_A_309_297#_c_253_n 0.00394323f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_99 N_B_c_90_n N_Y_c_281_n 0.00865686f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_100 B N_Y_c_281_n 0.0174927f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_101 N_B_c_90_n N_Y_c_294_n 0.00644736f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_102 N_B_c_91_n N_Y_c_283_n 0.01289f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_103 B N_Y_c_283_n 0.0310163f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_104 N_B_c_90_n N_Y_c_284_n 0.00119564f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_105 B N_Y_c_284_n 0.030835f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_106 N_B_c_93_n N_Y_c_284_n 0.00486271f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_107 N_B_c_90_n N_VGND_c_353_n 0.00268723f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_108 N_B_c_90_n N_VGND_c_358_n 0.00423334f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_109 N_B_c_91_n N_VGND_c_358_n 0.00437852f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_110 N_B_c_91_n N_VGND_c_359_n 0.00483063f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_111 N_B_c_90_n N_VGND_c_360_n 0.00598581f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_112 N_B_c_91_n N_VGND_c_360_n 0.00745263f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_113 N_C_c_136_n N_A_27_297#_c_179_n 0.00415386f $X=3.03 $Y=1.41 $X2=0 $Y2=0
cc_114 N_C_c_135_n N_A_27_297#_c_179_n 0.0152278f $X=2.69 $Y=1.18 $X2=0 $Y2=0
cc_115 N_C_c_136_n N_VPWR_c_212_n 0.00429453f $X=3.03 $Y=1.41 $X2=0 $Y2=0
cc_116 N_C_c_137_n N_VPWR_c_212_n 0.00429453f $X=3.5 $Y=1.41 $X2=0 $Y2=0
cc_117 N_C_c_136_n N_VPWR_c_210_n 0.00734734f $X=3.03 $Y=1.41 $X2=0 $Y2=0
cc_118 N_C_c_137_n N_VPWR_c_210_n 0.00708599f $X=3.5 $Y=1.41 $X2=0 $Y2=0
cc_119 N_C_c_135_n N_A_309_297#_M1003_d 0.00364872f $X=2.69 $Y=1.18 $X2=0 $Y2=0
cc_120 N_C_c_135_n N_A_309_297#_c_250_n 0.00823266f $X=2.69 $Y=1.18 $X2=0 $Y2=0
cc_121 N_C_c_135_n N_A_309_297#_c_253_n 0.0152506f $X=2.69 $Y=1.18 $X2=0 $Y2=0
cc_122 N_C_c_136_n N_A_309_297#_c_251_n 0.0143578f $X=3.03 $Y=1.41 $X2=0 $Y2=0
cc_123 N_C_c_137_n N_A_309_297#_c_251_n 0.01161f $X=3.5 $Y=1.41 $X2=0 $Y2=0
cc_124 N_C_c_132_n N_Y_c_283_n 0.0108632f $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_125 N_C_c_156_p N_Y_c_283_n 0.0267838f $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_126 N_C_c_135_n N_Y_c_283_n 0.0406302f $X=2.69 $Y=1.18 $X2=0 $Y2=0
cc_127 N_C_c_132_n N_Y_c_306_n 0.0112055f $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_128 N_C_c_132_n N_Y_c_285_n 0.00133045f $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_129 N_C_c_133_n N_Y_c_285_n 0.0115202f $X=3.525 $Y=0.995 $X2=0 $Y2=0
cc_130 N_C_c_134_n N_Y_c_285_n 0.00491863f $X=3.5 $Y=1.202 $X2=0 $Y2=0
cc_131 N_C_c_132_n Y 4.90655e-19 $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_132 N_C_c_136_n Y 0.00102406f $X=3.03 $Y=1.41 $X2=0 $Y2=0
cc_133 N_C_c_137_n Y 0.0163943f $X=3.5 $Y=1.41 $X2=0 $Y2=0
cc_134 N_C_c_133_n Y 0.00473468f $X=3.525 $Y=0.995 $X2=0 $Y2=0
cc_135 N_C_c_156_p Y 0.0258404f $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_136 N_C_c_134_n Y 0.0292604f $X=3.5 $Y=1.202 $X2=0 $Y2=0
cc_137 N_C_c_135_n Y 0.0122233f $X=2.69 $Y=1.18 $X2=0 $Y2=0
cc_138 N_C_c_133_n N_VGND_c_355_n 0.0045387f $X=3.525 $Y=0.995 $X2=0 $Y2=0
cc_139 N_C_c_132_n N_VGND_c_356_n 0.0042235f $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_140 N_C_c_133_n N_VGND_c_356_n 0.00437852f $X=3.525 $Y=0.995 $X2=0 $Y2=0
cc_141 N_C_c_132_n N_VGND_c_359_n 0.00483063f $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_142 N_C_c_132_n N_VGND_c_360_n 0.00729686f $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_143 N_C_c_133_n N_VGND_c_360_n 0.00719616f $X=3.525 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_27_297#_c_176_n N_VPWR_M1000_d 0.00187091f $X=1.095 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_145 N_A_27_297#_c_176_n N_VPWR_c_211_n 0.0143191f $X=1.095 $Y=1.54 $X2=0
+ $Y2=0
cc_146 N_A_27_297#_c_195_p N_VPWR_c_212_n 0.0149311f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_147 N_A_27_297#_M1000_s N_VPWR_c_210_n 0.00358889f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_148 N_A_27_297#_M1008_s N_VPWR_c_210_n 0.00370124f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_149 N_A_27_297#_M1004_d N_VPWR_c_210_n 0.00234744f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_150 N_A_27_297#_c_199_p N_VPWR_c_210_n 0.00974347f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_151 N_A_27_297#_c_195_p N_VPWR_c_210_n 0.00955092f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_152 N_A_27_297#_c_199_p N_VPWR_c_214_n 0.0165369f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_153 N_A_27_297#_c_177_n N_A_309_297#_M1002_s 0.00187091f $X=2.035 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_154 N_A_27_297#_c_177_n N_A_309_297#_c_260_n 0.0143018f $X=2.035 $Y=1.54
+ $X2=0 $Y2=0
cc_155 N_A_27_297#_M1004_d N_A_309_297#_c_250_n 0.0065032f $X=2.015 $Y=1.485
+ $X2=0 $Y2=0
cc_156 N_A_27_297#_c_177_n N_A_309_297#_c_250_n 0.00385532f $X=2.035 $Y=1.54
+ $X2=0 $Y2=0
cc_157 N_A_27_297#_c_179_n N_A_309_297#_c_250_n 0.0153739f $X=2.16 $Y=1.62 $X2=0
+ $Y2=0
cc_158 N_A_27_297#_c_179_n N_A_309_297#_c_253_n 0.0125002f $X=2.16 $Y=1.62 $X2=0
+ $Y2=0
cc_159 N_A_27_297#_c_176_n N_Y_c_281_n 0.00217122f $X=1.095 $Y=1.54 $X2=0 $Y2=0
cc_160 N_A_27_297#_c_178_n N_Y_c_281_n 0.00524452f $X=1.22 $Y=1.62 $X2=0 $Y2=0
cc_161 N_VPWR_c_210_n N_A_309_297#_M1002_s 0.00297222f $X=3.91 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_162 N_VPWR_c_210_n N_A_309_297#_M1003_d 0.00217523f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_163 N_VPWR_c_210_n N_A_309_297#_M1007_d 0.00217519f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_164 N_VPWR_c_212_n N_A_309_297#_c_250_n 0.0545557f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_165 N_VPWR_c_210_n N_A_309_297#_c_250_n 0.0324382f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_166 N_VPWR_c_212_n N_A_309_297#_c_270_n 0.0149886f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_167 N_VPWR_c_210_n N_A_309_297#_c_270_n 0.00962421f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_168 N_VPWR_c_212_n N_A_309_297#_c_251_n 0.0549564f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_169 N_VPWR_c_210_n N_A_309_297#_c_251_n 0.0335386f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_170 N_VPWR_c_212_n N_A_309_297#_c_274_n 0.0134651f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_171 N_VPWR_c_210_n N_A_309_297#_c_274_n 0.00808434f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_172 N_VPWR_c_210_n N_Y_M1003_s 0.00232895f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_173 N_A_309_297#_c_251_n N_Y_M1003_s 0.00345323f $X=3.61 $Y=2.38 $X2=0 $Y2=0
cc_174 N_A_309_297#_M1007_d Y 0.00288792f $X=3.59 $Y=1.485 $X2=0 $Y2=0
cc_175 N_A_309_297#_c_251_n Y 0.00388117f $X=3.61 $Y=2.38 $X2=0 $Y2=0
cc_176 N_A_309_297#_c_279_p Y 0.0172271f $X=3.735 $Y=1.96 $X2=0 $Y2=0
cc_177 N_A_309_297#_c_251_n N_Y_c_324_n 0.0128011f $X=3.61 $Y=2.38 $X2=0 $Y2=0
cc_178 N_Y_c_281_n N_VGND_M1011_s 0.00162089f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_179 N_Y_c_283_n N_VGND_M1010_d 0.00281828f $X=3.05 $Y=0.815 $X2=0 $Y2=0
cc_180 N_Y_c_283_n N_VGND_M1001_d 0.00281828f $X=3.05 $Y=0.815 $X2=0 $Y2=0
cc_181 N_Y_c_285_n N_VGND_M1009_d 0.0028133f $X=3.737 $Y=0.905 $X2=0 $Y2=0
cc_182 N_Y_c_282_n N_VGND_c_351_n 0.00835456f $X=0.915 $Y=0.815 $X2=0 $Y2=0
cc_183 N_Y_c_288_n N_VGND_c_352_n 0.0231806f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_184 N_Y_c_281_n N_VGND_c_352_n 0.00254521f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_185 N_Y_c_281_n N_VGND_c_353_n 0.0122559f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_186 N_Y_c_285_n N_VGND_c_354_n 8.44018e-19 $X=3.737 $Y=0.905 $X2=0 $Y2=0
cc_187 N_Y_c_285_n N_VGND_c_355_n 0.0223917f $X=3.737 $Y=0.905 $X2=0 $Y2=0
cc_188 N_Y_c_283_n N_VGND_c_356_n 0.00455335f $X=3.05 $Y=0.815 $X2=0 $Y2=0
cc_189 N_Y_c_306_n N_VGND_c_356_n 0.0227209f $X=3.265 $Y=0.39 $X2=0 $Y2=0
cc_190 N_Y_c_281_n N_VGND_c_358_n 0.00198695f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_191 N_Y_c_294_n N_VGND_c_358_n 0.0231806f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_192 N_Y_c_283_n N_VGND_c_358_n 0.00254521f $X=3.05 $Y=0.815 $X2=0 $Y2=0
cc_193 N_Y_c_283_n N_VGND_c_359_n 0.0629774f $X=3.05 $Y=0.815 $X2=0 $Y2=0
cc_194 N_Y_M1005_d N_VGND_c_360_n 0.00304143f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_195 N_Y_M1006_s N_VGND_c_360_n 0.00304143f $X=1.505 $Y=0.235 $X2=0 $Y2=0
cc_196 N_Y_M1001_s N_VGND_c_360_n 0.00305443f $X=3.08 $Y=0.235 $X2=0 $Y2=0
cc_197 N_Y_c_288_n N_VGND_c_360_n 0.0143352f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_198 N_Y_c_281_n N_VGND_c_360_n 0.0094839f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_199 N_Y_c_294_n N_VGND_c_360_n 0.0143352f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_200 N_Y_c_283_n N_VGND_c_360_n 0.0169329f $X=3.05 $Y=0.815 $X2=0 $Y2=0
cc_201 N_Y_c_306_n N_VGND_c_360_n 0.0142163f $X=3.265 $Y=0.39 $X2=0 $Y2=0
cc_202 N_Y_c_285_n N_VGND_c_360_n 0.00259547f $X=3.737 $Y=0.905 $X2=0 $Y2=0
