* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
X0 a_27_410# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_335_297# a_224_297# a_425_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_335_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 X a_335_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND D_N a_224_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_335_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 VGND a_224_297# a_335_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_335_297# a_27_410# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_625_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 a_27_410# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X10 VGND a_335_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_531_297# B a_625_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 VPWR D_N a_224_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X13 VGND B a_335_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 X a_335_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 X a_335_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 VGND a_335_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VPWR a_335_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 X a_335_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_425_297# a_27_410# a_531_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
