* File: sky130_fd_sc_hdll__o221ai_4.spice
* Created: Wed Sep  2 08:45:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o221ai_4.pex.spice"
.subckt sky130_fd_sc_hdll__o221ai_4  VNB VPB C1 B1 B2 A1 A2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2	A2
* A1	A1
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1006 N_Y_M1006_d N_C1_M1006_g N_A_27_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.2145 PD=0.97 PS=1.96 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.3
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1016 N_Y_M1006_d N_C1_M1016_g N_A_27_47#_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1020 N_Y_M1020_d N_C1_M1020_g N_A_27_47#_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1031 N_Y_M1020_d N_C1_M1031_g N_A_27_47#_M1031_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.169 PD=0.97 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1021 N_A_27_47#_M1021_d N_B1_M1021_g N_A_511_47#_M1021_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.2015 PD=0.97 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75007.3 A=0.0975 P=1.6 MULT=1
MM1023 N_A_27_47#_M1021_d N_B1_M1023_g N_A_511_47#_M1023_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75006.8 A=0.0975 P=1.6 MULT=1
MM1033 N_A_27_47#_M1033_d N_B1_M1033_g N_A_511_47#_M1023_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.2 SB=75006.4 A=0.0975 P=1.6 MULT=1
MM1007 N_A_511_47#_M1007_d N_B2_M1007_g N_A_27_47#_M1033_d VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75006 A=0.0975 P=1.6 MULT=1
MM1027 N_A_511_47#_M1007_d N_B2_M1027_g N_A_27_47#_M1027_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75002.1 SB=75005.5 A=0.0975 P=1.6 MULT=1
MM1029 N_A_511_47#_M1029_d N_B2_M1029_g N_A_27_47#_M1027_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75002.5 SB=75005 A=0.0975 P=1.6 MULT=1
MM1039 N_A_511_47#_M1029_d N_B2_M1039_g N_A_27_47#_M1039_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75003.1 SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1037 N_A_27_47#_M1039_s N_B1_M1037_g N_A_511_47#_M1037_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.13 PD=0.97 PS=1.05 NRD=8.304 NRS=13.836 M=1 R=4.33333
+ SA=75003.5 SB=75004 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A1_M1009_g N_A_511_47#_M1037_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.13 PD=0.92 PS=1.05 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.1
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1004 N_A_511_47#_M1004_d N_A2_M1004_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75004.5
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1017 N_A_511_47#_M1004_d N_A2_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75005
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1019 N_A_511_47#_M1019_d N_A2_M1019_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75005.4
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1036 N_A_511_47#_M1019_d N_A2_M1036_g N_VGND_M1036_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75006
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1036_s N_A1_M1011_g N_A_511_47#_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75006.4
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1014_d N_A1_M1014_g N_A_511_47#_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75006.8
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1032 N_VGND_M1014_d N_A1_M1032_g N_A_511_47#_M1032_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.2015 PD=0.97 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75007.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_Y_M1000_d N_C1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90009.7 A=0.18 P=2.36 MULT=1
MM1008 N_Y_M1000_d N_C1_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.7
+ SB=90009.3 A=0.18 P=2.36 MULT=1
MM1012 N_Y_M1012_d N_C1_M1012_g N_VPWR_M1008_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.1
+ SB=90008.8 A=0.18 P=2.36 MULT=1
MM1024 N_Y_M1012_d N_C1_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.405 PD=1.29 PS=1.81 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.6
+ SB=90008.3 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1024_s N_B1_M1013_g N_A_601_297#_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.405 AS=0.145 PD=1.81 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.6 SB=90007.3 A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1018_d N_B1_M1018_g N_A_601_297#_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.1 SB=90006.9 A=0.18 P=2.36 MULT=1
MM1028 N_VPWR_M1018_d N_B1_M1028_g N_A_601_297#_M1028_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90006.4 A=0.18 P=2.36 MULT=1
MM1001 N_A_601_297#_M1028_s N_B2_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90004
+ SB=90005.9 A=0.18 P=2.36 MULT=1
MM1010 N_A_601_297#_M1010_d N_B2_M1010_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.5 SB=90005.5 A=0.18 P=2.36 MULT=1
MM1025 N_A_601_297#_M1010_d N_B2_M1025_g N_Y_M1025_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.9 SB=90005 A=0.18 P=2.36 MULT=1
MM1030 N_A_601_297#_M1030_d N_B2_M1030_g N_Y_M1025_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.4 SB=90004.5 A=0.18 P=2.36 MULT=1
MM1034 N_VPWR_M1034_d N_B1_M1034_g N_A_601_297#_M1030_d VPB PHIGHVT L=0.18 W=1
+ AD=0.185 AS=0.145 PD=1.37 PS=1.29 NRD=8.8453 NRS=0.9653 M=1 R=5.55556
+ SA=90005.9 SB=90004.1 A=0.18 P=2.36 MULT=1
MM1003 N_A_1369_297#_M1003_d N_A1_M1003_g N_VPWR_M1034_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.185 PD=1.29 PS=1.37 NRD=0.9653 NRS=8.8453 M=1 R=5.55556
+ SA=90006.4 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1002 N_Y_M1002_d N_A2_M1002_g N_A_1369_297#_M1003_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90006.9 SB=90003 A=0.18 P=2.36 MULT=1
MM1005 N_Y_M1002_d N_A2_M1005_g N_A_1369_297#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90007.4 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1015 N_Y_M1015_d N_A2_M1015_g N_A_1369_297#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90007.8 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1038 N_Y_M1015_d N_A2_M1038_g N_A_1369_297#_M1038_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90008.3 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1022 N_A_1369_297#_M1038_s N_A1_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90008.8 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1026 N_A_1369_297#_M1026_d N_A1_M1026_g N_VPWR_M1022_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90009.3 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1035 N_A_1369_297#_M1026_d N_A1_M1035_g N_VPWR_M1035_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.305 PD=1.29 PS=2.61 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90009.7 SB=90000.2 A=0.18 P=2.36 MULT=1
DX40_noxref VNB VPB NWDIODE A=17.5908 P=25.13
pX41_noxref noxref_15 B1 B1 PROBETYPE=1
pX42_noxref noxref_16 B2 B2 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o221ai_4.pxi.spice"
*
.ends
*
*
