* File: sky130_fd_sc_hdll__or4_1.pxi.spice
* Created: Wed Sep  2 08:49:12 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR4_1%D N_D_c_61_n N_D_M1003_g N_D_M1000_g D D
+ N_D_c_60_n PM_SKY130_FD_SC_HDLL__OR4_1%D
x_PM_SKY130_FD_SC_HDLL__OR4_1%C N_C_c_87_n N_C_M1009_g N_C_M1005_g C C C C
+ PM_SKY130_FD_SC_HDLL__OR4_1%C
x_PM_SKY130_FD_SC_HDLL__OR4_1%B N_B_c_126_n N_B_c_127_n N_B_c_129_n N_B_c_130_n
+ N_B_M1006_g N_B_M1007_g N_B_c_128_n B B B N_B_c_132_n B B
+ PM_SKY130_FD_SC_HDLL__OR4_1%B
x_PM_SKY130_FD_SC_HDLL__OR4_1%A N_A_c_168_n N_A_M1004_g N_A_M1002_g A
+ N_A_c_170_n A PM_SKY130_FD_SC_HDLL__OR4_1%A
x_PM_SKY130_FD_SC_HDLL__OR4_1%A_27_297# N_A_27_297#_M1000_d N_A_27_297#_M1007_d
+ N_A_27_297#_M1003_s N_A_27_297#_c_208_n N_A_27_297#_M1008_g
+ N_A_27_297#_c_209_n N_A_27_297#_M1001_g N_A_27_297#_c_217_n
+ N_A_27_297#_c_230_n N_A_27_297#_c_210_n N_A_27_297#_c_211_n
+ N_A_27_297#_c_289_p N_A_27_297#_c_212_n N_A_27_297#_c_244_n
+ N_A_27_297#_c_218_n N_A_27_297#_c_219_n N_A_27_297#_c_213_n
+ N_A_27_297#_c_220_n N_A_27_297#_c_214_n N_A_27_297#_c_215_n
+ PM_SKY130_FD_SC_HDLL__OR4_1%A_27_297#
x_PM_SKY130_FD_SC_HDLL__OR4_1%VPWR N_VPWR_M1004_d N_VPWR_c_312_n N_VPWR_c_313_n
+ N_VPWR_c_314_n VPWR N_VPWR_c_315_n N_VPWR_c_311_n
+ PM_SKY130_FD_SC_HDLL__OR4_1%VPWR
x_PM_SKY130_FD_SC_HDLL__OR4_1%X N_X_M1001_d N_X_M1008_d N_X_c_335_n N_X_c_337_n
+ N_X_c_336_n X PM_SKY130_FD_SC_HDLL__OR4_1%X
x_PM_SKY130_FD_SC_HDLL__OR4_1%VGND N_VGND_M1000_s N_VGND_M1005_d N_VGND_M1002_d
+ N_VGND_c_354_n N_VGND_c_355_n N_VGND_c_356_n VGND N_VGND_c_357_n
+ N_VGND_c_358_n N_VGND_c_359_n N_VGND_c_360_n N_VGND_c_361_n N_VGND_c_362_n
+ PM_SKY130_FD_SC_HDLL__OR4_1%VGND
cc_1 VNB N_D_M1000_g 0.0338621f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_2 VNB D 0.0267048f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_3 VNB N_D_c_60_n 0.0387829f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_C_c_87_n 0.0211609f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_C_M1005_g 0.0263621f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_6 VNB C 0.00587769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_B_c_126_n 0.00672106f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_8 VNB N_B_c_127_n 0.0217657f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.695
cc_9 VNB N_B_c_128_n 0.0143238f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_c_168_n 0.0195868f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_11 VNB N_A_M1002_g 0.0285024f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_12 VNB N_A_c_170_n 0.00455736f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.202
cc_13 VNB N_A_27_297#_c_208_n 0.0242606f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_297#_c_209_n 0.0211873f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_15 VNB N_A_27_297#_c_210_n 0.00370552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_297#_c_211_n 0.0032469f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_297#_c_212_n 0.00154854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_297#_c_213_n 0.00155735f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_297#_c_214_n 0.00264294f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_297#_c_215_n 0.00196069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_311_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_X_c_335_n 0.0137322f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.202
cc_23 VNB N_X_c_336_n 0.0252742f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_24 VNB N_VGND_c_354_n 0.0115524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_355_n 0.0193841f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.202
cc_26 VNB N_VGND_c_356_n 8.49086e-19 $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_27 VNB N_VGND_c_357_n 0.0164754f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.16
cc_28 VNB N_VGND_c_358_n 0.0129653f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_359_n 0.0258474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_360_n 0.192674f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_361_n 0.00544933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_362_n 0.0102719f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VPB N_D_c_61_n 0.0213218f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_34 VPB D 0.00359125f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_35 VPB N_D_c_60_n 0.0178492f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_36 VPB N_C_c_87_n 0.0240375f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_37 VPB C 0.0018628f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_B_c_129_n 0.00563909f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.695
cc_39 VPB N_B_c_130_n 0.0497412f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_40 VPB N_B_M1006_g 0.0107365f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.475
cc_41 VPB N_B_c_132_n 0.0521007f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_c_168_n 0.0274047f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_43 VPB N_A_c_170_n 0.00326435f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.202
cc_44 VPB N_A_27_297#_c_208_n 0.0312736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_297#_c_217_n 0.00597646f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_46 VPB N_A_27_297#_c_218_n 0.00156472f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_27_297#_c_219_n 0.021096f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_27_297#_c_220_n 0.00210247f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_312_n 0.0116412f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.475
cc_50 VPB N_VPWR_c_313_n 0.0540731f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_51 VPB N_VPWR_c_314_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_315_n 0.0258752f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_311_n 0.0665821f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_X_c_337_n 0.0051537f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_55 VPB N_X_c_336_n 0.00928216f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_56 VPB X 0.0321952f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_57 N_D_c_61_n N_C_c_87_n 0.0216385f $X=0.495 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_58 D N_C_c_87_n 2.56827e-19 $X=0.15 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_59 N_D_c_60_n N_C_c_87_n 0.0236968f $X=0.495 $Y=1.202 $X2=-0.19 $Y2=-0.24
cc_60 N_D_M1000_g N_C_M1005_g 0.0191324f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_61 N_D_c_61_n C 0.00392215f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_62 D C 0.0230021f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_63 N_D_c_60_n C 0.00564283f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_64 N_D_c_61_n N_B_c_132_n 0.00528936f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_65 N_D_c_61_n N_A_27_297#_c_217_n 0.0140535f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_66 D N_A_27_297#_c_217_n 9.67991e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_67 N_D_M1000_g N_A_27_297#_c_211_n 0.00384738f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_68 D N_A_27_297#_c_211_n 0.00494723f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_69 N_D_c_61_n N_A_27_297#_c_219_n 0.00661664f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_70 D N_A_27_297#_c_219_n 0.0243773f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_71 N_D_c_60_n N_A_27_297#_c_219_n 0.00192889f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_72 N_D_M1000_g N_VGND_c_355_n 0.00426752f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_73 D N_VGND_c_355_n 0.0271923f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_74 N_D_c_60_n N_VGND_c_355_n 0.00130319f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_75 N_D_M1000_g N_VGND_c_356_n 5.72193e-19 $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_76 N_D_M1000_g N_VGND_c_357_n 0.00555245f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_77 D N_VGND_c_357_n 2.15148e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_78 N_D_M1000_g N_VGND_c_360_n 0.0113233f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_79 D N_VGND_c_360_n 0.00195847f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_80 N_C_M1005_g N_B_c_126_n 0.020096f $X=1.05 $Y=0.475 $X2=-0.19 $Y2=-0.24
cc_81 N_C_c_87_n N_B_c_127_n 0.020096f $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_82 C N_B_c_127_n 0.00761675f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_83 C N_B_c_129_n 0.00303888f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_84 N_C_c_87_n N_B_M1006_g 0.0348558f $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_85 C N_B_M1006_g 0.00416637f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_86 N_C_M1005_g N_B_c_128_n 0.0137426f $X=1.05 $Y=0.475 $X2=0 $Y2=0
cc_87 N_C_c_87_n N_B_c_132_n 0.00527095f $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_88 C N_A_c_168_n 9.45363e-19 $X=1.17 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_89 N_C_c_87_n N_A_c_170_n 2.10621e-19 $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_90 C N_A_c_170_n 0.0273602f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_91 N_C_c_87_n N_A_27_297#_c_217_n 0.0110624f $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_92 C N_A_27_297#_c_217_n 0.0411859f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_93 N_C_M1005_g N_A_27_297#_c_230_n 0.00520782f $X=1.05 $Y=0.475 $X2=0 $Y2=0
cc_94 N_C_c_87_n N_A_27_297#_c_210_n 0.00308093f $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_95 N_C_M1005_g N_A_27_297#_c_210_n 0.0110002f $X=1.05 $Y=0.475 $X2=0 $Y2=0
cc_96 C N_A_27_297#_c_210_n 0.040618f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_97 N_C_c_87_n N_A_27_297#_c_211_n 9.23324e-19 $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_98 C N_A_27_297#_c_211_n 0.0152593f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_99 N_C_c_87_n N_A_27_297#_c_219_n 9.15255e-19 $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_100 C N_A_27_297#_c_219_n 0.00730153f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_101 C N_A_27_297#_c_220_n 0.00596189f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_102 C A_117_297# 0.00421255f $X=1.17 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_103 C A_223_297# 0.00139712f $X=1.17 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_104 N_C_M1005_g N_VGND_c_356_n 0.0101314f $X=1.05 $Y=0.475 $X2=0 $Y2=0
cc_105 N_C_M1005_g N_VGND_c_357_n 0.00187556f $X=1.05 $Y=0.475 $X2=0 $Y2=0
cc_106 N_C_M1005_g N_VGND_c_360_n 0.00271727f $X=1.05 $Y=0.475 $X2=0 $Y2=0
cc_107 N_B_c_127_n N_A_c_168_n 0.0171853f $X=1.445 $Y=1.31 $X2=-0.19 $Y2=-0.24
cc_108 N_B_c_129_n N_A_c_168_n 0.00358094f $X=1.445 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_109 N_B_M1006_g N_A_c_168_n 0.0202457f $X=1.445 $Y=1.695 $X2=-0.19 $Y2=-0.24
cc_110 N_B_c_132_n N_A_c_168_n 6.66635e-19 $X=1.48 $Y=2.31 $X2=-0.19 $Y2=-0.24
cc_111 N_B_c_128_n N_A_M1002_g 0.0166388f $X=1.445 $Y=0.76 $X2=0 $Y2=0
cc_112 N_B_c_127_n N_A_c_170_n 0.00834593f $X=1.445 $Y=1.31 $X2=0 $Y2=0
cc_113 N_B_c_129_n N_A_c_170_n 7.53623e-19 $X=1.445 $Y=1.41 $X2=0 $Y2=0
cc_114 N_B_c_130_n N_A_27_297#_c_217_n 7.17844e-19 $X=1.445 $Y=2.035 $X2=0 $Y2=0
cc_115 N_B_M1006_g N_A_27_297#_c_217_n 0.0161318f $X=1.445 $Y=1.695 $X2=0 $Y2=0
cc_116 N_B_c_132_n N_A_27_297#_c_217_n 0.0923574f $X=1.48 $Y=2.31 $X2=0 $Y2=0
cc_117 N_B_c_126_n N_A_27_297#_c_210_n 0.0114865f $X=1.445 $Y=0.86 $X2=0 $Y2=0
cc_118 N_B_c_128_n N_A_27_297#_c_210_n 0.00713678f $X=1.445 $Y=0.76 $X2=0 $Y2=0
cc_119 N_B_c_132_n N_A_27_297#_c_244_n 0.00163296f $X=1.48 $Y=2.31 $X2=0 $Y2=0
cc_120 N_B_c_132_n N_A_27_297#_c_219_n 0.0261176f $X=1.48 $Y=2.31 $X2=0 $Y2=0
cc_121 N_B_M1006_g N_A_27_297#_c_220_n 0.00517026f $X=1.445 $Y=1.695 $X2=0 $Y2=0
cc_122 N_B_c_132_n N_A_27_297#_c_220_n 0.0138065f $X=1.48 $Y=2.31 $X2=0 $Y2=0
cc_123 N_B_c_130_n N_VPWR_c_312_n 0.00506259f $X=1.445 $Y=2.035 $X2=0 $Y2=0
cc_124 N_B_c_132_n N_VPWR_c_312_n 0.0210036f $X=1.48 $Y=2.31 $X2=0 $Y2=0
cc_125 N_B_c_130_n N_VPWR_c_313_n 0.00687133f $X=1.445 $Y=2.035 $X2=0 $Y2=0
cc_126 N_B_c_132_n N_VPWR_c_313_n 0.0911288f $X=1.48 $Y=2.31 $X2=0 $Y2=0
cc_127 N_B_c_130_n N_VPWR_c_311_n 0.00939765f $X=1.445 $Y=2.035 $X2=0 $Y2=0
cc_128 N_B_c_132_n N_VPWR_c_311_n 0.0658875f $X=1.48 $Y=2.31 $X2=0 $Y2=0
cc_129 N_B_c_128_n N_VGND_c_356_n 0.00720367f $X=1.445 $Y=0.76 $X2=0 $Y2=0
cc_130 N_B_c_128_n N_VGND_c_358_n 0.00322006f $X=1.445 $Y=0.76 $X2=0 $Y2=0
cc_131 N_B_c_128_n N_VGND_c_360_n 0.00408297f $X=1.445 $Y=0.76 $X2=0 $Y2=0
cc_132 N_B_c_128_n N_VGND_c_362_n 5.53035e-19 $X=1.445 $Y=0.76 $X2=0 $Y2=0
cc_133 N_A_c_168_n N_A_27_297#_c_208_n 0.0346242f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_c_170_n N_A_27_297#_c_208_n 0.00106108f $X=1.93 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_M1002_g N_A_27_297#_c_209_n 0.0178481f $X=1.99 $Y=0.475 $X2=0 $Y2=0
cc_136 N_A_c_170_n N_A_27_297#_c_217_n 0.00407647f $X=1.93 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_c_170_n N_A_27_297#_c_210_n 0.00931915f $X=1.93 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_c_168_n N_A_27_297#_c_212_n 0.00240831f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_M1002_g N_A_27_297#_c_212_n 0.0117073f $X=1.99 $Y=0.475 $X2=0 $Y2=0
cc_140 N_A_c_170_n N_A_27_297#_c_212_n 0.0205685f $X=1.93 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A_c_168_n N_A_27_297#_c_244_n 0.0155871f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_c_170_n N_A_27_297#_c_244_n 0.016167f $X=1.93 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_c_168_n N_A_27_297#_c_218_n 0.00173315f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_168_n N_A_27_297#_c_213_n 4.61771e-19 $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_c_170_n N_A_27_297#_c_213_n 0.0146461f $X=1.93 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A_c_168_n N_A_27_297#_c_220_n 0.0025153f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_c_170_n N_A_27_297#_c_220_n 0.0135338f $X=1.93 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_c_168_n N_A_27_297#_c_214_n 0.00458419f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_c_170_n N_A_27_297#_c_214_n 0.0283407f $X=1.93 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A_M1002_g N_A_27_297#_c_215_n 0.00177765f $X=1.99 $Y=0.475 $X2=0 $Y2=0
cc_151 N_A_c_168_n N_VPWR_c_312_n 0.00342204f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_c_168_n N_VPWR_c_313_n 0.00351268f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_c_168_n N_VPWR_c_311_n 0.00445321f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_M1002_g N_VGND_c_356_n 5.02092e-19 $X=1.99 $Y=0.475 $X2=0 $Y2=0
cc_155 N_A_M1002_g N_VGND_c_358_n 0.00188229f $X=1.99 $Y=0.475 $X2=0 $Y2=0
cc_156 N_A_M1002_g N_VGND_c_360_n 0.00270076f $X=1.99 $Y=0.475 $X2=0 $Y2=0
cc_157 N_A_M1002_g N_VGND_c_362_n 0.01011f $X=1.99 $Y=0.475 $X2=0 $Y2=0
cc_158 N_A_27_297#_c_217_n A_117_297# 0.00291425f $X=1.66 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_159 N_A_27_297#_c_217_n A_223_297# 0.00134267f $X=1.66 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_160 N_A_27_297#_c_217_n A_307_297# 0.00146656f $X=1.66 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_161 N_A_27_297#_c_220_n A_307_297# 0.0056502f $X=1.745 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_162 N_A_27_297#_c_244_n N_VPWR_M1004_d 0.00563715f $X=2.265 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_163 N_A_27_297#_c_208_n N_VPWR_c_312_n 0.00499543f $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_164 N_A_27_297#_c_244_n N_VPWR_c_312_n 0.0204259f $X=2.265 $Y=1.58 $X2=0
+ $Y2=0
cc_165 N_A_27_297#_c_220_n N_VPWR_c_312_n 0.00457307f $X=1.745 $Y=1.58 $X2=0
+ $Y2=0
cc_166 N_A_27_297#_c_208_n N_VPWR_c_315_n 0.00702461f $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_167 N_A_27_297#_c_208_n N_VPWR_c_311_n 0.0148715f $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_168 N_A_27_297#_c_209_n N_X_c_335_n 0.00961493f $X=2.53 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_27_297#_c_208_n N_X_c_337_n 0.0233895f $X=2.505 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_27_297#_c_244_n N_X_c_337_n 0.00747506f $X=2.265 $Y=1.58 $X2=0 $Y2=0
cc_171 N_A_27_297#_c_208_n N_X_c_336_n 0.00162368f $X=2.505 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A_27_297#_c_209_n N_X_c_336_n 0.0127645f $X=2.53 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A_27_297#_c_218_n N_X_c_336_n 0.00560514f $X=2.35 $Y=1.495 $X2=0 $Y2=0
cc_174 N_A_27_297#_c_214_n N_X_c_336_n 0.0143335f $X=2.47 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_27_297#_c_215_n N_X_c_336_n 0.00506543f $X=2.41 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_27_297#_c_210_n N_VGND_M1005_d 0.00160115f $X=1.645 $Y=0.74 $X2=0
+ $Y2=0
cc_177 N_A_27_297#_c_212_n N_VGND_M1002_d 0.00670822f $X=2.265 $Y=0.74 $X2=0
+ $Y2=0
cc_178 N_A_27_297#_c_215_n N_VGND_M1002_d 6.98847e-19 $X=2.41 $Y=0.995 $X2=0
+ $Y2=0
cc_179 N_A_27_297#_c_230_n N_VGND_c_356_n 0.0118543f $X=0.76 $Y=0.47 $X2=0 $Y2=0
cc_180 N_A_27_297#_c_210_n N_VGND_c_356_n 0.0196541f $X=1.645 $Y=0.74 $X2=0
+ $Y2=0
cc_181 N_A_27_297#_c_289_p N_VGND_c_356_n 0.0110177f $X=1.73 $Y=0.47 $X2=0 $Y2=0
cc_182 N_A_27_297#_c_230_n N_VGND_c_357_n 0.00876148f $X=0.76 $Y=0.47 $X2=0
+ $Y2=0
cc_183 N_A_27_297#_c_210_n N_VGND_c_357_n 0.00282959f $X=1.645 $Y=0.74 $X2=0
+ $Y2=0
cc_184 N_A_27_297#_c_210_n N_VGND_c_358_n 0.00310196f $X=1.645 $Y=0.74 $X2=0
+ $Y2=0
cc_185 N_A_27_297#_c_289_p N_VGND_c_358_n 0.00876148f $X=1.73 $Y=0.47 $X2=0
+ $Y2=0
cc_186 N_A_27_297#_c_212_n N_VGND_c_358_n 0.00232988f $X=2.265 $Y=0.74 $X2=0
+ $Y2=0
cc_187 N_A_27_297#_c_209_n N_VGND_c_359_n 0.00585385f $X=2.53 $Y=0.995 $X2=0
+ $Y2=0
cc_188 N_A_27_297#_c_209_n N_VGND_c_360_n 0.0123583f $X=2.53 $Y=0.995 $X2=0
+ $Y2=0
cc_189 N_A_27_297#_c_230_n N_VGND_c_360_n 0.00625722f $X=0.76 $Y=0.47 $X2=0
+ $Y2=0
cc_190 N_A_27_297#_c_210_n N_VGND_c_360_n 0.0123925f $X=1.645 $Y=0.74 $X2=0
+ $Y2=0
cc_191 N_A_27_297#_c_289_p N_VGND_c_360_n 0.00625722f $X=1.73 $Y=0.47 $X2=0
+ $Y2=0
cc_192 N_A_27_297#_c_212_n N_VGND_c_360_n 0.00689417f $X=2.265 $Y=0.74 $X2=0
+ $Y2=0
cc_193 N_A_27_297#_c_208_n N_VGND_c_362_n 2.73815e-19 $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_194 N_A_27_297#_c_209_n N_VGND_c_362_n 0.00498808f $X=2.53 $Y=0.995 $X2=0
+ $Y2=0
cc_195 N_A_27_297#_c_289_p N_VGND_c_362_n 0.0135697f $X=1.73 $Y=0.47 $X2=0 $Y2=0
cc_196 N_A_27_297#_c_212_n N_VGND_c_362_n 0.0278587f $X=2.265 $Y=0.74 $X2=0
+ $Y2=0
cc_197 N_VPWR_c_311_n N_X_M1008_d 0.0108199f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_198 N_VPWR_c_315_n X 0.0189133f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_199 N_VPWR_c_311_n X 0.0103212f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_200 N_X_c_335_n N_VGND_c_359_n 0.00886414f $X=2.99 $Y=0.587 $X2=0 $Y2=0
cc_201 N_X_M1001_d N_VGND_c_360_n 0.010552f $X=2.605 $Y=0.235 $X2=0 $Y2=0
cc_202 N_X_c_335_n N_VGND_c_360_n 0.00924648f $X=2.99 $Y=0.587 $X2=0 $Y2=0
