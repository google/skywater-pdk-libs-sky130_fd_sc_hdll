* File: sky130_fd_sc_hdll__nor4b_2.pex.spice
* Created: Wed Sep  2 08:41:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR4B_2%A 1 3 4 6 7 9 10 12 13 14 15 24 29
c43 24 0 1.30114e-19 $X=0.965 $Y=1.202
r44 24 25 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r45 22 24 43.1263 $w=3.8e-07 $l=3.4e-07 $layer=POLY_cond $X=0.625 $Y=1.202
+ $X2=0.965 $Y2=1.202
r46 22 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.625
+ $Y=1.16 $X2=0.625 $Y2=1.16
r47 20 22 16.4895 $w=3.8e-07 $l=1.3e-07 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.625 $Y2=1.202
r48 19 20 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r49 14 15 22.974 $w=2.08e-07 $l=4.35e-07 $layer=LI1_cond $X=0.725 $Y=1.18
+ $X2=1.16 $Y2=1.18
r50 14 29 5.28139 $w=2.08e-07 $l=1e-07 $layer=LI1_cond $X=0.725 $Y=1.18
+ $X2=0.625 $Y2=1.18
r51 13 29 20.5974 $w=2.08e-07 $l=3.9e-07 $layer=LI1_cond $X=0.235 $Y=1.18
+ $X2=0.625 $Y2=1.18
r52 10 25 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r53 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r54 7 24 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r55 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r56 4 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r57 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r58 1 19 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.202
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_2%B 1 3 4 6 7 9 10 12 13 14 15 24 29
c40 15 0 1.30114e-19 $X=2.445 $Y=1.105
r41 24 25 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=1.93 $Y2=1.202
r42 22 24 21.5632 $w=3.8e-07 $l=1.7e-07 $layer=POLY_cond $X=1.735 $Y=1.202
+ $X2=1.905 $Y2=1.202
r43 22 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.735
+ $Y=1.16 $X2=1.735 $Y2=1.16
r44 20 22 38.0526 $w=3.8e-07 $l=3e-07 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.735 $Y2=1.202
r45 19 20 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.202
+ $X2=1.435 $Y2=1.202
r46 14 15 24.0303 $w=2.08e-07 $l=4.55e-07 $layer=LI1_cond $X=2.075 $Y=1.18
+ $X2=2.53 $Y2=1.18
r47 14 29 21.6537 $w=2.08e-07 $l=4.1e-07 $layer=LI1_cond $X=2.075 $Y=1.18
+ $X2=1.665 $Y2=1.18
r48 13 29 1.84848 $w=2.08e-07 $l=3.5e-08 $layer=LI1_cond $X=1.63 $Y=1.18
+ $X2=1.665 $Y2=1.18
r49 10 25 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r50 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r51 7 24 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r52 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r53 4 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r54 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r55 1 19 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.202
r56 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995 $X2=1.41
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_2%C 1 3 4 6 7 9 10 12 13 14 22 25
r46 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.4 $Y=1.202
+ $X2=3.425 $Y2=1.202
r47 20 22 21.5632 $w=3.8e-07 $l=1.7e-07 $layer=POLY_cond $X=3.23 $Y=1.202
+ $X2=3.4 $Y2=1.202
r48 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.23
+ $Y=1.16 $X2=3.23 $Y2=1.16
r49 18 20 38.0526 $w=3.8e-07 $l=3e-07 $layer=POLY_cond $X=2.93 $Y=1.202 $X2=3.23
+ $Y2=1.202
r50 17 18 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=2.905 $Y=1.202
+ $X2=2.93 $Y2=1.202
r51 14 21 11.8831 $w=2.08e-07 $l=2.25e-07 $layer=LI1_cond $X=3.455 $Y=1.18
+ $X2=3.23 $Y2=1.18
r52 13 21 12.4113 $w=2.08e-07 $l=2.35e-07 $layer=LI1_cond $X=2.995 $Y=1.18
+ $X2=3.23 $Y2=1.18
r53 13 25 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=2.995 $Y=1.18
+ $X2=2.99 $Y2=1.18
r54 10 23 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.425 $Y=0.995
+ $X2=3.425 $Y2=1.202
r55 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.425 $Y=0.995
+ $X2=3.425 $Y2=0.56
r56 7 22 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.4 $Y=1.41 $X2=3.4
+ $Y2=1.202
r57 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.4 $Y=1.41 $X2=3.4
+ $Y2=1.985
r58 4 18 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.93 $Y=1.41
+ $X2=2.93 $Y2=1.202
r59 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.93 $Y=1.41 $X2=2.93
+ $Y2=1.985
r60 1 17 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.905 $Y=0.995
+ $X2=2.905 $Y2=1.202
r61 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.905 $Y=0.995
+ $X2=2.905 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_2%A_754_21# 1 2 7 9 10 12 13 15 16 18 19 25
+ 29 30 34 38 39
r71 38 39 11.2584 $w=3.53e-07 $l=2.5e-07 $layer=LI1_cond $X=5.042 $Y=2.285
+ $X2=5.042 $Y2=2.035
r72 34 36 11.0961 $w=3.53e-07 $l=2.45e-07 $layer=LI1_cond $X=5.042 $Y=0.66
+ $X2=5.042 $Y2=0.905
r73 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.885
+ $Y=1.16 $X2=4.885 $Y2=1.16
r74 26 29 0.716491 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=4.95 $Y=1.245
+ $X2=4.885 $Y2=1.16
r75 26 39 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.95 $Y=1.245
+ $X2=4.95 $Y2=2.035
r76 25 29 0.716491 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=4.95 $Y=1.075
+ $X2=4.885 $Y2=1.16
r77 25 36 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.95 $Y=1.075
+ $X2=4.95 $Y2=0.905
r78 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.315 $Y=1.202
+ $X2=4.34 $Y2=1.202
r79 21 22 56.4447 $w=3.8e-07 $l=4.45e-07 $layer=POLY_cond $X=3.87 $Y=1.202
+ $X2=4.315 $Y2=1.202
r80 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.845 $Y=1.202
+ $X2=3.87 $Y2=1.202
r81 19 30 77.8133 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=4.44 $Y=1.16
+ $X2=4.885 $Y2=1.16
r82 19 23 13.6483 $w=3.8e-07 $l=1.19164e-07 $layer=POLY_cond $X=4.44 $Y=1.16
+ $X2=4.34 $Y2=1.202
r83 16 23 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.34 $Y=1.41
+ $X2=4.34 $Y2=1.202
r84 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.34 $Y=1.41
+ $X2=4.34 $Y2=1.985
r85 13 22 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.315 $Y=0.995
+ $X2=4.315 $Y2=1.202
r86 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.315 $Y=0.995
+ $X2=4.315 $Y2=0.56
r87 10 21 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.87 $Y=1.41
+ $X2=3.87 $Y2=1.202
r88 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.87 $Y=1.41
+ $X2=3.87 $Y2=1.985
r89 7 20 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.845 $Y=0.995
+ $X2=3.845 $Y2=1.202
r90 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.845 $Y=0.995
+ $X2=3.845 $Y2=0.56
r91 2 38 600 $w=1.7e-07 $l=2.755e-07 $layer=licon1_PDIFF $count=1 $X=4.97
+ $Y=2.065 $X2=5.095 $Y2=2.285
r92 1 34 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=4.97
+ $Y=0.465 $X2=5.095 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_2%D_N 3 5 6 8 9 12 14 15 16 21 23
r33 15 16 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.75 $Y=1.53
+ $X2=5.75 $Y2=1.87
r34 15 23 10.4574 $w=2.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.75 $Y=1.53
+ $X2=5.75 $Y2=1.285
r35 14 23 3.04322 $w=2.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.75 $Y=1.18
+ $X2=5.75 $Y2=1.285
r36 12 22 37.7763 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=5.392 $Y=1.16
+ $X2=5.392 $Y2=1.325
r37 12 21 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=5.392 $Y=1.16
+ $X2=5.392 $Y2=0.995
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.37
+ $Y=1.16 $X2=5.37 $Y2=1.16
r39 9 14 3.91272 $w=2.1e-07 $l=1.35e-07 $layer=LI1_cond $X=5.615 $Y=1.18
+ $X2=5.75 $Y2=1.18
r40 9 11 12.9394 $w=2.08e-07 $l=2.45e-07 $layer=LI1_cond $X=5.615 $Y=1.18
+ $X2=5.37 $Y2=1.18
r41 6 8 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.33 $Y=1.99 $X2=5.33
+ $Y2=2.275
r42 5 6 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=5.33 $Y=1.89 $X2=5.33
+ $Y2=1.99
r43 5 22 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=5.33 $Y=1.89 $X2=5.33
+ $Y2=1.325
r44 3 21 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.305 $Y=0.675
+ $X2=5.305 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_2%A_27_297# 1 2 3 12 16 17 20 22 26 29
r45 24 26 0.151637 $w=3.78e-07 $l=5e-09 $layer=LI1_cond $X=2.115 $Y=1.625
+ $X2=2.115 $Y2=1.63
r46 23 29 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.325 $Y=1.54
+ $X2=1.2 $Y2=1.54
r47 22 24 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=1.925 $Y=1.54
+ $X2=2.115 $Y2=1.625
r48 22 23 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.925 $Y=1.54
+ $X2=1.325 $Y2=1.54
r49 18 29 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=1.625
+ $X2=1.2 $Y2=1.54
r50 18 20 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.2 $Y=1.625 $X2=1.2
+ $Y2=2.3
r51 16 29 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.075 $Y=1.54
+ $X2=1.2 $Y2=1.54
r52 16 17 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.075 $Y=1.54
+ $X2=0.425 $Y2=1.54
r53 12 14 23.0489 $w=3.38e-07 $l=6.8e-07 $layer=LI1_cond $X=0.255 $Y=1.63
+ $X2=0.255 $Y2=2.31
r54 10 17 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.255 $Y=1.625
+ $X2=0.425 $Y2=1.54
r55 10 12 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=0.255 $Y=1.625
+ $X2=0.255 $Y2=1.63
r56 3 26 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.63
r57 2 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.62
r58 2 20 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.3
r59 1 14 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.31
r60 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_2%VPWR 1 2 11 15 18 19 20 30 31 34
r58 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r59 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r60 28 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r61 27 28 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r62 25 28 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=1.15 $Y=2.72 $X2=5.29
+ $Y2=2.72
r63 25 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r64 24 27 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=5.29 $Y2=2.72
r65 24 25 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r66 22 34 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=0.75 $Y2=2.72
r67 22 24 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=1.15 $Y2=2.72
r68 20 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 18 27 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.44 $Y=2.72 $X2=5.29
+ $Y2=2.72
r70 18 19 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.44 $Y=2.72
+ $X2=5.565 $Y2=2.72
r71 17 30 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=5.69 $Y=2.72 $X2=5.75
+ $Y2=2.72
r72 17 19 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.69 $Y=2.72
+ $X2=5.565 $Y2=2.72
r73 13 19 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=2.635
+ $X2=5.565 $Y2=2.72
r74 13 15 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.565 $Y=2.635
+ $X2=5.565 $Y2=2.3
r75 9 34 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r76 9 11 35.6493 $w=2.08e-07 $l=6.75e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=1.96
r77 2 15 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=5.42
+ $Y=2.065 $X2=5.565 $Y2=2.3
r78 1 11 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_2%A_305_297# 1 2 9 11 12 15
r21 13 15 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=3.185 $Y=2.295
+ $X2=3.185 $Y2=1.96
r22 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.08 $Y=2.38
+ $X2=3.185 $Y2=2.295
r23 11 12 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=3.08 $Y=2.38
+ $X2=1.755 $Y2=2.38
r24 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.65 $Y=2.295
+ $X2=1.755 $Y2=2.38
r25 7 9 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=1.65 $Y=2.295
+ $X2=1.65 $Y2=1.96
r26 2 15 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.02
+ $Y=1.485 $X2=3.165 $Y2=1.96
r27 1 9 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_2%A_514_297# 1 2 3 12 14 15 16 17 18 22
r43 20 22 15.7579 $w=2.43e-07 $l=3.35e-07 $layer=LI1_cond $X=4.572 $Y=2.295
+ $X2=4.572 $Y2=1.96
r44 19 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.76 $Y=2.38
+ $X2=3.635 $Y2=2.38
r45 18 20 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=4.45 $Y=2.38
+ $X2=4.572 $Y2=2.295
r46 18 19 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.45 $Y=2.38 $X2=3.76
+ $Y2=2.38
r47 17 27 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=2.295
+ $X2=3.635 $Y2=2.38
r48 16 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=1.625
+ $X2=3.635 $Y2=1.54
r49 16 17 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=3.635 $Y=1.625
+ $X2=3.635 $Y2=2.295
r50 14 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.51 $Y=1.54
+ $X2=3.635 $Y2=1.54
r51 14 15 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.51 $Y=1.54
+ $X2=2.86 $Y2=1.54
r52 10 15 8.24022 $w=1.7e-07 $l=2.31633e-07 $layer=LI1_cond $X=2.667 $Y=1.625
+ $X2=2.86 $Y2=1.54
r53 10 12 0.149668 $w=3.83e-07 $l=5e-09 $layer=LI1_cond $X=2.667 $Y=1.625
+ $X2=2.667 $Y2=1.63
r54 3 22 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.43
+ $Y=1.485 $X2=4.575 $Y2=1.96
r55 2 27 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.49
+ $Y=1.485 $X2=3.635 $Y2=2.3
r56 2 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.49
+ $Y=1.485 $X2=3.635 $Y2=1.62
r57 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.57
+ $Y=1.485 $X2=2.695 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_2%Y 1 2 3 4 5 18 20 21 24 26 30 32 36 41 42
+ 43 44 45 46 54
r93 45 54 2.43459 $w=4.51e-07 $l=9e-08 $layer=LI1_cond $X=4.235 $Y=1.53
+ $X2=4.235 $Y2=1.62
r94 45 46 9.19734 $w=4.51e-07 $l=3.4e-07 $layer=LI1_cond $X=4.235 $Y=1.53
+ $X2=4.235 $Y2=1.19
r95 41 46 6.78104 $w=4.51e-07 $l=1.45069e-07 $layer=LI1_cond $X=4.167 $Y=1.075
+ $X2=4.235 $Y2=1.19
r96 40 44 3.39178 $w=2.92e-07 $l=1.26214e-07 $layer=LI1_cond $X=4.167 $Y=0.905
+ $X2=4.08 $Y2=0.815
r97 40 41 9.19734 $w=2.03e-07 $l=1.7e-07 $layer=LI1_cond $X=4.167 $Y=0.905
+ $X2=4.167 $Y2=1.075
r98 34 44 3.39178 $w=2.92e-07 $l=9e-08 $layer=LI1_cond $X=4.08 $Y=0.725 $X2=4.08
+ $Y2=0.815
r99 34 36 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.08 $Y=0.725
+ $X2=4.08 $Y2=0.39
r100 33 43 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.33 $Y=0.815
+ $X2=3.14 $Y2=0.815
r101 32 44 3.13665 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.89 $Y=0.815
+ $X2=4.08 $Y2=0.815
r102 32 33 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.89 $Y=0.815
+ $X2=3.33 $Y2=0.815
r103 28 43 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=3.14 $Y=0.725 $X2=3.14
+ $Y2=0.815
r104 28 30 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.14 $Y=0.725
+ $X2=3.14 $Y2=0.39
r105 27 42 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=0.815
+ $X2=1.645 $Y2=0.815
r106 26 43 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.95 $Y=0.815
+ $X2=3.14 $Y2=0.815
r107 26 27 68.702 $w=1.78e-07 $l=1.115e-06 $layer=LI1_cond $X=2.95 $Y=0.815
+ $X2=1.835 $Y2=0.815
r108 22 42 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=1.645 $Y=0.725
+ $X2=1.645 $Y2=0.815
r109 22 24 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.645 $Y=0.725
+ $X2=1.645 $Y2=0.39
r110 20 42 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=0.815
+ $X2=1.645 $Y2=0.815
r111 20 21 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.455 $Y=0.815
+ $X2=0.895 $Y2=0.815
r112 16 21 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=0.705 $Y=0.725
+ $X2=0.895 $Y2=0.815
r113 16 18 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.705 $Y=0.725
+ $X2=0.705 $Y2=0.39
r114 5 54 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.96
+ $Y=1.485 $X2=4.105 $Y2=1.62
r115 4 36 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.92
+ $Y=0.235 $X2=4.105 $Y2=0.39
r116 3 30 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=2.98
+ $Y=0.235 $X2=3.165 $Y2=0.39
r117 2 24 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.39
r118 1 18 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_2%VGND 1 2 3 4 5 6 7 22 24 26 30 36 40 44 47
+ 48 50 51 53 54 55 68 69 75 80 88
r87 87 88 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=0.235
+ $X2=2.78 $Y2=0.235
r88 84 87 3.08364 $w=6.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=0.235
+ $X2=2.695 $Y2=0.235
r89 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r90 82 84 7.2886 $w=6.38e-07 $l=3.9e-07 $layer=LI1_cond $X=2.14 $Y=0.235
+ $X2=2.53 $Y2=0.235
r91 79 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r92 78 82 1.30821 $w=6.38e-07 $l=7e-08 $layer=LI1_cond $X=2.07 $Y=0.235 $X2=2.14
+ $Y2=0.235
r93 78 80 7.61355 $w=6.38e-07 $l=1.5e-08 $layer=LI1_cond $X=2.07 $Y=0.235
+ $X2=2.055 $Y2=0.235
r94 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r95 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r96 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r97 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r98 66 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r99 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r100 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r101 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r102 60 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r103 60 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r104 59 88 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=2.78
+ $Y2=0
r105 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r106 55 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r107 55 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r108 53 65 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.44 $Y=0 $X2=5.29
+ $Y2=0
r109 53 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.44 $Y=0 $X2=5.565
+ $Y2=0
r110 52 68 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=5.69 $Y=0 $X2=5.75
+ $Y2=0
r111 52 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.69 $Y=0 $X2=5.565
+ $Y2=0
r112 50 62 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.49 $Y=0 $X2=4.37
+ $Y2=0
r113 50 51 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=4.49 $Y=0 $X2=4.592
+ $Y2=0
r114 49 65 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=4.695 $Y=0
+ $X2=5.29 $Y2=0
r115 49 51 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=4.695 $Y=0
+ $X2=4.592 $Y2=0
r116 47 59 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.55 $Y=0 $X2=3.45
+ $Y2=0
r117 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=0 $X2=3.635
+ $Y2=0
r118 46 62 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=4.37
+ $Y2=0
r119 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.635
+ $Y2=0
r120 42 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=0.085
+ $X2=5.565 $Y2=0
r121 42 44 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=5.565 $Y=0.085
+ $X2=5.565 $Y2=0.66
r122 38 51 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.592 $Y=0.085
+ $X2=4.592 $Y2=0
r123 38 40 16.5011 $w=2.03e-07 $l=3.05e-07 $layer=LI1_cond $X=4.592 $Y=0.085
+ $X2=4.592 $Y2=0.39
r124 34 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=0.085
+ $X2=3.635 $Y2=0
r125 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.635 $Y=0.085
+ $X2=3.635 $Y2=0.39
r126 33 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.2
+ $Y2=0
r127 33 80 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=2.055 $Y2=0
r128 28 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.085 $X2=1.2
+ $Y2=0
r129 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0.39
r130 27 72 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r131 26 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.2
+ $Y2=0
r132 26 27 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=0.345 $Y2=0
r133 22 72 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.172 $Y2=0
r134 22 24 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.215 $Y2=0.39
r135 7 44 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=5.38
+ $Y=0.465 $X2=5.565 $Y2=0.66
r136 6 40 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.39
+ $Y=0.235 $X2=4.575 $Y2=0.39
r137 5 36 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.5
+ $Y=0.235 $X2=3.635 $Y2=0.39
r138 4 87 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.57
+ $Y=0.235 $X2=2.695 $Y2=0.39
r139 3 82 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.39
r140 2 30 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.39
r141 1 24 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

