* File: sky130_fd_sc_hdll__nand3b_2.pex.spice
* Created: Thu Aug 27 19:14:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND3B_2%A_N 3 6 7 9 10 13 20
r33 14 20 5.54545 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=0.595 $Y=1.175
+ $X2=0.695 $Y2=1.175
r34 13 16 36.6246 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=1.16
+ $X2=0.587 $Y2=1.325
r35 13 15 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=1.16
+ $X2=0.587 $Y2=0.995
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.595
+ $Y=1.16 $X2=0.595 $Y2=1.16
r37 10 20 2.77273 $w=1.98e-07 $l=5e-08 $layer=LI1_cond $X=0.745 $Y=1.175
+ $X2=0.695 $Y2=1.175
r38 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r39 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.89 $X2=0.495
+ $Y2=1.99
r40 6 16 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.495 $Y=1.89
+ $X2=0.495 $Y2=1.325
r41 3 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.445
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_2%C 3 5 7 8 10 13 15 16 24 27
c46 24 0 1.32669e-19 $X=1.56 $Y=1.217
r47 24 25 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=1.56 $Y=1.217
+ $X2=1.585 $Y2=1.217
r48 22 24 33.5118 $w=3.38e-07 $l=2.35e-07 $layer=POLY_cond $X=1.325 $Y=1.217
+ $X2=1.56 $Y2=1.217
r49 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.16 $X2=1.325 $Y2=1.16
r50 20 22 33.5118 $w=3.38e-07 $l=2.35e-07 $layer=POLY_cond $X=1.09 $Y=1.217
+ $X2=1.325 $Y2=1.217
r51 19 20 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=1.065 $Y=1.217
+ $X2=1.09 $Y2=1.217
r52 16 23 24.4 $w=1.98e-07 $l=4.4e-07 $layer=LI1_cond $X=1.765 $Y=1.175
+ $X2=1.325 $Y2=1.175
r53 15 23 6.65455 $w=1.98e-07 $l=1.2e-07 $layer=LI1_cond $X=1.205 $Y=1.175
+ $X2=1.325 $Y2=1.175
r54 15 27 2.77273 $w=1.98e-07 $l=5e-08 $layer=LI1_cond $X=1.205 $Y=1.175
+ $X2=1.155 $Y2=1.175
r55 11 25 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.585 $Y=1.025
+ $X2=1.585 $Y2=1.217
r56 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.585 $Y=1.025
+ $X2=1.585 $Y2=0.56
r57 8 24 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.56 $Y=1.41
+ $X2=1.56 $Y2=1.217
r58 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.56 $Y=1.41
+ $X2=1.56 $Y2=1.985
r59 5 20 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.09 $Y=1.41
+ $X2=1.09 $Y2=1.217
r60 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.09 $Y=1.41 $X2=1.09
+ $Y2=1.985
r61 1 19 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.065 $Y=1.025
+ $X2=1.065 $Y2=1.217
r62 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.065 $Y=1.025
+ $X2=1.065 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_2%B 1 3 4 6 9 13 15 19 20 21 22 30
c45 22 0 1.32669e-19 $X=3.23 $Y=1.105
c46 13 0 3.57174e-19 $X=3.095 $Y=0.56
r47 21 22 32.7182 $w=1.98e-07 $l=5.9e-07 $layer=LI1_cond $X=2.725 $Y=1.175
+ $X2=3.315 $Y2=1.175
r48 21 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.725
+ $Y=1.16 $X2=2.725 $Y2=1.16
r49 20 21 24.9545 $w=1.98e-07 $l=4.5e-07 $layer=LI1_cond $X=2.275 $Y=1.175
+ $X2=2.725 $Y2=1.175
r50 20 30 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=2.275 $Y=1.175
+ $X2=2.27 $Y2=1.175
r51 19 27 65.5412 $w=2.7e-07 $l=2.95e-07 $layer=POLY_cond $X=3.02 $Y=1.16
+ $X2=2.725 $Y2=1.16
r52 17 18 18.3131 $w=3.29e-07 $l=1.25e-07 $layer=POLY_cond $X=2.5 $Y=1.217
+ $X2=2.625 $Y2=1.217
r53 16 17 68.8571 $w=3.29e-07 $l=4.7e-07 $layer=POLY_cond $X=2.03 $Y=1.217
+ $X2=2.5 $Y2=1.217
r54 15 27 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=2.7 $Y=1.16
+ $X2=2.725 $Y2=1.16
r55 15 18 12.6805 $w=3.29e-07 $l=9.94987e-08 $layer=POLY_cond $X=2.7 $Y=1.16
+ $X2=2.625 $Y2=1.217
r56 11 19 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.095 $Y=1.025
+ $X2=3.02 $Y2=1.16
r57 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.095 $Y=1.025
+ $X2=3.095 $Y2=0.56
r58 7 18 21.1507 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.625 $Y=1.025
+ $X2=2.625 $Y2=1.217
r59 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.625 $Y=1.025
+ $X2=2.625 $Y2=0.56
r60 4 17 16.8611 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.5 $Y=1.41 $X2=2.5
+ $Y2=1.217
r61 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.5 $Y=1.41 $X2=2.5
+ $Y2=1.985
r62 1 16 16.8611 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.03 $Y=1.41
+ $X2=2.03 $Y2=1.217
r63 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.03 $Y=1.41 $X2=2.03
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_2%A_27_47# 1 2 9 11 13 14 16 19 22 25 29 33
+ 36 38 39 44
c86 29 0 9.80354e-20 $X=3.835 $Y=1.16
c87 9 0 1.52405e-19 $X=3.515 $Y=0.56
r88 44 45 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=4.01 $Y=1.217
+ $X2=4.035 $Y2=1.217
r89 41 42 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=3.515 $Y=1.217
+ $X2=3.54 $Y2=1.217
r90 38 39 10.9812 $w=3.18e-07 $l=2.35e-07 $layer=LI1_cond $X=0.25 $Y=2.3
+ $X2=0.25 $Y2=2.065
r91 33 35 10.9812 $w=3.18e-07 $l=2.35e-07 $layer=LI1_cond $X=0.25 $Y=0.42
+ $X2=0.25 $Y2=0.655
r92 30 44 24.9556 $w=3.38e-07 $l=1.75e-07 $layer=POLY_cond $X=3.835 $Y=1.217
+ $X2=4.01 $Y2=1.217
r93 30 42 42.068 $w=3.38e-07 $l=2.95e-07 $layer=POLY_cond $X=3.835 $Y=1.217
+ $X2=3.54 $Y2=1.217
r94 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.835
+ $Y=1.16 $X2=3.835 $Y2=1.16
r95 27 29 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.835 $Y=1.445
+ $X2=3.835 $Y2=1.16
r96 26 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.53
+ $X2=0.175 $Y2=1.53
r97 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.67 $Y=1.53
+ $X2=3.835 $Y2=1.445
r98 25 26 222.471 $w=1.68e-07 $l=3.41e-06 $layer=LI1_cond $X=3.67 $Y=1.53
+ $X2=0.26 $Y2=1.53
r99 23 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.175 $Y=1.615
+ $X2=0.175 $Y2=1.53
r100 23 39 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.175 $Y=1.615
+ $X2=0.175 $Y2=2.065
r101 22 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.175 $Y=1.445
+ $X2=0.175 $Y2=1.53
r102 22 35 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.175 $Y=1.445
+ $X2=0.175 $Y2=0.655
r103 17 45 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.035 $Y=1.025
+ $X2=4.035 $Y2=1.217
r104 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.035 $Y=1.025
+ $X2=4.035 $Y2=0.56
r105 14 44 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.01 $Y=1.41
+ $X2=4.01 $Y2=1.217
r106 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.01 $Y=1.41
+ $X2=4.01 $Y2=1.985
r107 11 42 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.54 $Y=1.41
+ $X2=3.54 $Y2=1.217
r108 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.54 $Y=1.41
+ $X2=3.54 $Y2=1.985
r109 7 41 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.515 $Y=1.025
+ $X2=3.515 $Y2=1.217
r110 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.515 $Y=1.025
+ $X2=3.515 $Y2=0.56
r111 2 38 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
r112 1 33 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_2%VPWR 1 2 3 4 5 20 24 28 32 34 36 39 40 42
+ 43 45 46 47 59 64 68
r78 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r79 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r80 62 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r81 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r82 59 67 4.30612 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=4.16 $Y=2.72 $X2=4.38
+ $Y2=2.72
r83 59 61 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.16 $Y=2.72
+ $X2=3.91 $Y2=2.72
r84 58 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r85 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r86 55 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r87 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r88 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r89 52 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r90 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r91 49 64 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.94 $Y=2.72
+ $X2=0.785 $Y2=2.72
r92 49 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.94 $Y=2.72
+ $X2=1.61 $Y2=2.72
r93 47 65 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r94 45 57 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.09 $Y=2.72 $X2=2.99
+ $Y2=2.72
r95 45 46 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.09 $Y=2.72 $X2=3.24
+ $Y2=2.72
r96 44 61 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.39 $Y=2.72
+ $X2=3.91 $Y2=2.72
r97 44 46 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.39 $Y=2.72 $X2=3.24
+ $Y2=2.72
r98 42 54 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.65 $Y=2.72
+ $X2=2.53 $Y2=2.72
r99 42 43 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.65 $Y=2.72
+ $X2=2.775 $Y2=2.72
r100 41 57 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.9 $Y=2.72 $X2=2.99
+ $Y2=2.72
r101 41 43 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.9 $Y=2.72
+ $X2=2.775 $Y2=2.72
r102 39 51 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.71 $Y=2.72 $X2=1.61
+ $Y2=2.72
r103 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=2.72
+ $X2=1.795 $Y2=2.72
r104 38 54 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.88 $Y=2.72
+ $X2=2.53 $Y2=2.72
r105 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.88 $Y=2.72
+ $X2=1.795 $Y2=2.72
r106 34 67 3.13172 $w=2.9e-07 $l=1.16619e-07 $layer=LI1_cond $X=4.305 $Y=2.635
+ $X2=4.38 $Y2=2.72
r107 34 36 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=4.305 $Y=2.635
+ $X2=4.305 $Y2=2.34
r108 30 46 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.24 $Y=2.635
+ $X2=3.24 $Y2=2.72
r109 30 32 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=3.24 $Y=2.635
+ $X2=3.24 $Y2=2.34
r110 26 43 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=2.635
+ $X2=2.775 $Y2=2.72
r111 26 28 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.775 $Y=2.635
+ $X2=2.775 $Y2=2.34
r112 22 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=2.635
+ $X2=1.795 $Y2=2.72
r113 22 24 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.795 $Y=2.635
+ $X2=1.795 $Y2=2.34
r114 18 64 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=2.635
+ $X2=0.785 $Y2=2.72
r115 18 20 23.6065 $w=3.08e-07 $l=6.35e-07 $layer=LI1_cond $X=0.785 $Y=2.635
+ $X2=0.785 $Y2=2
r116 5 36 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.1
+ $Y=1.485 $X2=4.245 $Y2=2.34
r117 4 32 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=3.18
+ $Y=1.485 $X2=3.305 $Y2=2.34
r118 3 28 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.59
+ $Y=1.485 $X2=2.735 $Y2=2.34
r119 2 24 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=1.485 $X2=1.795 $Y2=2.34
r120 1 20 300 $w=1.7e-07 $l=2.40312e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=2.065 $X2=0.795 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_2%Y 1 2 3 4 15 19 21 27 30 32 34 37 38
r75 37 38 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=4.37 $Y=1.19
+ $X2=4.37 $Y2=1.53
r76 36 38 12.2447 $w=2.38e-07 $l=2.55e-07 $layer=LI1_cond $X=4.37 $Y=1.785
+ $X2=4.37 $Y2=1.53
r77 35 37 13.6853 $w=2.38e-07 $l=2.85e-07 $layer=LI1_cond $X=4.37 $Y=0.905
+ $X2=4.37 $Y2=1.19
r78 28 34 7.27225 $w=1.95e-07 $l=1.5e-07 $layer=LI1_cond $X=3.86 $Y=1.895
+ $X2=3.71 $Y2=1.895
r79 27 36 6.83327 $w=2.2e-07 $l=1.66132e-07 $layer=LI1_cond $X=4.25 $Y=1.895
+ $X2=4.37 $Y2=1.785
r80 27 28 20.4297 $w=2.18e-07 $l=3.9e-07 $layer=LI1_cond $X=4.25 $Y=1.895
+ $X2=3.86 $Y2=1.895
r81 21 35 6.84722 $w=2.7e-07 $l=1.8554e-07 $layer=LI1_cond $X=4.25 $Y=0.77
+ $X2=4.37 $Y2=0.905
r82 21 23 20.2745 $w=2.68e-07 $l=4.75e-07 $layer=LI1_cond $X=4.25 $Y=0.77
+ $X2=3.775 $Y2=0.77
r83 20 32 8.63406 $w=1.95e-07 $l=2.02114e-07 $layer=LI1_cond $X=2.43 $Y=1.87
+ $X2=2.24 $Y2=1.895
r84 19 34 7.27225 $w=1.95e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.56 $Y=1.87
+ $X2=3.71 $Y2=1.895
r85 19 20 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=3.56 $Y=1.87
+ $X2=2.43 $Y2=1.87
r86 16 30 4.72888 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.49 $Y=1.895 $X2=1.3
+ $Y2=1.895
r87 15 32 8.63406 $w=1.95e-07 $l=1.9e-07 $layer=LI1_cond $X=2.05 $Y=1.895
+ $X2=2.24 $Y2=1.895
r88 15 16 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=2.05 $Y=1.895
+ $X2=1.49 $Y2=1.895
r89 4 34 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.63
+ $Y=1.485 $X2=3.775 $Y2=1.96
r90 3 32 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.12
+ $Y=1.485 $X2=2.265 $Y2=2
r91 2 30 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.18
+ $Y=1.485 $X2=1.325 $Y2=2
r92 1 23 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=3.59
+ $Y=0.235 $X2=3.775 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_2%VGND 1 2 11 15 18 19 20 30 31 34 37
r56 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r57 30 31 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r58 28 31 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=4.37
+ $Y2=0
r59 27 30 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=4.37
+ $Y2=0
r60 27 28 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r61 25 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r62 25 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r63 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r64 22 34 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.94 $Y=0 $X2=0.785
+ $Y2=0
r65 22 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.94 $Y=0 $X2=1.61
+ $Y2=0
r66 20 35 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r67 20 37 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r68 18 24 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.71 $Y=0 $X2=1.61
+ $Y2=0
r69 18 19 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.71 $Y=0 $X2=1.835
+ $Y2=0
r70 17 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.96 $Y=0 $X2=2.07
+ $Y2=0
r71 17 19 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.96 $Y=0 $X2=1.835
+ $Y2=0
r72 13 19 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.835 $Y=0.085
+ $X2=1.835 $Y2=0
r73 13 15 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.835 $Y=0.085
+ $X2=1.835 $Y2=0.38
r74 9 34 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0
r75 9 11 10.9668 $w=3.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0.38
r76 2 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.66
+ $Y=0.235 $X2=1.795 $Y2=0.38
r77 1 11 91 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.795 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_2%A_228_47# 1 2 9 12 13 15 17
c31 15 0 1.91459e-19 $X=2.835 $Y=0.72
r32 13 17 6.78806 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.335 $Y=0.77
+ $X2=2.2 $Y2=0.77
r33 13 15 21.3415 $w=2.68e-07 $l=5e-07 $layer=LI1_cond $X=2.335 $Y=0.77
+ $X2=2.835 $Y2=0.77
r34 12 17 41.445 $w=1.88e-07 $l=7.1e-07 $layer=LI1_cond $X=1.49 $Y=0.81 $X2=2.2
+ $Y2=0.81
r35 7 12 7.85115 $w=1.9e-07 $l=2.32702e-07 $layer=LI1_cond $X=1.3 $Y=0.715
+ $X2=1.49 $Y2=0.81
r36 7 9 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.3 $Y=0.715 $X2=1.3
+ $Y2=0.38
r37 2 15 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.235 $X2=2.835 $Y2=0.72
r38 1 9 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=1.14
+ $Y=0.235 $X2=1.325 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_2%A_448_47# 1 2 3 10 16 20 23
c28 16 0 3.18121e-19 $X=3.305 $Y=0.72
r29 18 23 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.39 $Y=0.36 $X2=3.305
+ $Y2=0.36
r30 18 20 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=3.39 $Y=0.36
+ $X2=4.245 $Y2=0.36
r31 14 23 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.305 $Y=0.465
+ $X2=3.305 $Y2=0.36
r32 14 16 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.305 $Y=0.465
+ $X2=3.305 $Y2=0.72
r33 10 23 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=0.36 $X2=3.305
+ $Y2=0.36
r34 10 12 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=3.22 $Y=0.36
+ $X2=2.365 $Y2=0.36
r35 3 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.11
+ $Y=0.235 $X2=4.245 $Y2=0.38
r36 2 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.17
+ $Y=0.235 $X2=3.305 $Y2=0.38
r37 2 16 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.17
+ $Y=0.235 $X2=3.305 $Y2=0.72
r38 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.24
+ $Y=0.235 $X2=2.365 $Y2=0.38
.ends

