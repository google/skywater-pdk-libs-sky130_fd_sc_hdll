* File: sky130_fd_sc_hdll__diode_6.spice
* Created: Thu Aug 27 19:05:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__diode_6.pex.spice"
.subckt sky130_fd_sc_hdll__diode_6  VNB VPB DIODE VGND VPWR
* 
* DIODE	DIODE
* VPB	VPB
* VNB	VNB
D0_noxref VNB N_DIODE_D0_noxref_neg NDIODE  AREA=2.2032 PJ=7.9 M=1
+ AHFTEMPPERIM=7.9
DX1_noxref VNB VPB NWDIODE A=3.9228 P=11.02
*
.include "sky130_fd_sc_hdll__diode_6.pxi.spice"
*
.ends
*
*
