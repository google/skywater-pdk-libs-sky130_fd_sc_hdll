* File: sky130_fd_sc_hdll__o21a_2.pex.spice
* Created: Thu Aug 27 19:18:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O21A_2%A_79_21# 1 2 7 9 10 12 13 15 16 18 20 22 23
+ 24 25 26 29 31 33 36 44
r73 43 44 3.22193 $w=3.74e-07 $l=2.5e-08 $layer=POLY_cond $X=0.945 $Y=1.202
+ $X2=0.97 $Y2=1.202
r74 42 43 57.9947 $w=3.74e-07 $l=4.5e-07 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.945 $Y2=1.202
r75 41 42 3.22193 $w=3.74e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r76 37 44 14.1765 $w=3.74e-07 $l=1.1e-07 $layer=POLY_cond $X=1.08 $Y=1.202
+ $X2=0.97 $Y2=1.202
r77 36 38 8.67109 $w=3.58e-07 $l=1.7e-07 $layer=LI1_cond $X=1.175 $Y=1.16
+ $X2=1.175 $Y2=1.33
r78 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.08
+ $Y=1.16 $X2=1.08 $Y2=1.16
r79 31 40 3.15253 $w=2.6e-07 $l=1.1e-07 $layer=LI1_cond $X=2.245 $Y=2.005
+ $X2=2.245 $Y2=1.895
r80 31 33 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=2.245 $Y=2.005
+ $X2=2.245 $Y2=2.3
r81 27 29 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.73 $Y=0.635
+ $X2=1.73 $Y2=0.385
r82 25 40 3.72571 $w=2.2e-07 $l=1.3e-07 $layer=LI1_cond $X=2.115 $Y=1.895
+ $X2=2.245 $Y2=1.895
r83 25 26 39.8117 $w=2.18e-07 $l=7.6e-07 $layer=LI1_cond $X=2.115 $Y=1.895
+ $X2=1.355 $Y2=1.895
r84 23 27 7.31195 $w=2.05e-07 $l=2.09893e-07 $layer=LI1_cond $X=1.565 $Y=0.737
+ $X2=1.73 $Y2=0.635
r85 23 24 11.3614 $w=2.03e-07 $l=2.1e-07 $layer=LI1_cond $X=1.565 $Y=0.737
+ $X2=1.355 $Y2=0.737
r86 22 26 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.27 $Y=1.785
+ $X2=1.355 $Y2=1.895
r87 22 38 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.27 $Y=1.785
+ $X2=1.27 $Y2=1.33
r88 20 36 0.320123 $w=3.58e-07 $l=1e-08 $layer=LI1_cond $X=1.175 $Y=1.15
+ $X2=1.175 $Y2=1.16
r89 19 24 7.50588 $w=2.05e-07 $l=2.25699e-07 $layer=LI1_cond $X=1.175 $Y=0.84
+ $X2=1.355 $Y2=0.737
r90 19 20 9.92381 $w=3.58e-07 $l=3.1e-07 $layer=LI1_cond $X=1.175 $Y=0.84
+ $X2=1.175 $Y2=1.15
r91 16 44 19.8678 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.97 $Y=1.41
+ $X2=0.97 $Y2=1.202
r92 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.97 $Y=1.41
+ $X2=0.97 $Y2=1.985
r93 13 43 24.2268 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.945 $Y=0.995
+ $X2=0.945 $Y2=1.202
r94 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.945 $Y=0.995
+ $X2=0.945 $Y2=0.56
r95 10 42 19.8678 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r96 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r97 7 41 24.2268 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.202
r98 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
r99 2 40 600 $w=1.7e-07 $l=5.04455e-07 $layer=licon1_PDIFF $count=1 $X=2.06
+ $Y=1.485 $X2=2.21 $Y2=1.92
r100 2 33 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=2.06
+ $Y=1.485 $X2=2.21 $Y2=2.3
r101 1 29 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=1.605
+ $Y=0.235 $X2=1.73 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_2%B1 1 3 4 6 7 11
r29 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.79
+ $Y=1.16 $X2=1.79 $Y2=1.16
r30 7 11 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.74 $Y=1.53 $X2=1.74
+ $Y2=1.16
r31 4 10 39.4698 $w=3.94e-07 $l=2.27255e-07 $layer=POLY_cond $X=1.995 $Y=0.995
+ $X2=1.847 $Y2=1.16
r32 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.995 $Y=0.995
+ $X2=1.995 $Y2=0.56
r33 1 10 44.9511 $w=3.94e-07 $l=3.05369e-07 $layer=POLY_cond $X=1.97 $Y=1.41
+ $X2=1.847 $Y2=1.16
r34 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.97 $Y=1.41 $X2=1.97
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_2%A2 1 3 4 6 7 13
r36 12 13 19.6963 $w=2.73e-07 $l=4.7e-07 $layer=LI1_cond $X=2.937 $Y=1.4
+ $X2=2.937 $Y2=1.87
r37 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.485
+ $Y=1.16 $X2=2.485 $Y2=1.16
r38 7 12 7.02845 $w=3.75e-07 $l=2.47184e-07 $layer=LI1_cond $X=2.8 $Y=1.212
+ $X2=2.937 $Y2=1.4
r39 7 9 9.68052 $w=3.73e-07 $l=3.15e-07 $layer=LI1_cond $X=2.8 $Y=1.212
+ $X2=2.485 $Y2=1.212
r40 4 10 48.651 $w=2.87e-07 $l=2.76134e-07 $layer=POLY_cond $X=2.45 $Y=1.41
+ $X2=2.505 $Y2=1.16
r41 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.45 $Y=1.41 $X2=2.45
+ $Y2=1.985
r42 1 10 38.6443 $w=2.87e-07 $l=2.0106e-07 $layer=POLY_cond $X=2.425 $Y=0.995
+ $X2=2.505 $Y2=1.16
r43 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.425 $Y=0.995
+ $X2=2.425 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_2%A1 1 3 4 6 7 10
r29 10 12 33.7665 $w=3.64e-07 $l=2.55e-07 $layer=POLY_cond $X=3.13 $Y=1.202
+ $X2=3.385 $Y2=1.202
r30 9 10 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=3.105 $Y=1.202
+ $X2=3.13 $Y2=1.202
r31 7 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.385
+ $Y=1.16 $X2=3.385 $Y2=1.16
r32 4 10 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.13 $Y=1.41
+ $X2=3.13 $Y2=1.202
r33 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.13 $Y=1.41 $X2=3.13
+ $Y2=1.985
r34 1 9 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.105 $Y=0.995
+ $X2=3.105 $Y2=1.202
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.105 $Y=0.995
+ $X2=3.105 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_2%VPWR 1 2 3 10 12 14 16 18 25 39 42 45
r46 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r47 41 42 10.2865 $w=6.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.73 $Y=2.495
+ $X2=1.895 $Y2=2.495
r48 37 41 2.31499 $w=6.18e-07 $l=1.2e-07 $layer=LI1_cond $X=1.61 $Y=2.495
+ $X2=1.73 $Y2=2.495
r49 37 39 18.9677 $w=6.18e-07 $l=6.15e-07 $layer=LI1_cond $X=1.61 $Y=2.495
+ $X2=0.995 $Y2=2.495
r50 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r51 32 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r52 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r54 29 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r55 28 31 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r56 28 42 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=1.895 $Y2=2.72
r57 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 25 44 4.25865 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=3.245 $Y=2.72
+ $X2=3.462 $Y2=2.72
r59 25 31 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.245 $Y=2.72
+ $X2=2.99 $Y2=2.72
r60 24 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r61 23 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=0.995 $Y2=2.72
r62 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r63 21 34 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r64 21 23 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 18 24 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r66 18 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r67 14 44 3.14002 $w=2.85e-07 $l=1.16619e-07 $layer=LI1_cond $X=3.387 $Y=2.635
+ $X2=3.462 $Y2=2.72
r68 14 16 32.1471 $w=2.83e-07 $l=7.95e-07 $layer=LI1_cond $X=3.387 $Y=2.635
+ $X2=3.387 $Y2=1.84
r69 10 34 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r70 10 12 37.059 $w=2.53e-07 $l=8.2e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=1.815
r71 3 16 300 $w=1.7e-07 $l=4.23409e-07 $layer=licon1_PDIFF $count=2 $X=3.22
+ $Y=1.485 $X2=3.37 $Y2=1.84
r72 2 41 300 $w=1.7e-07 $l=1.14187e-06 $layer=licon1_PDIFF $count=2 $X=1.06
+ $Y=1.485 $X2=1.73 $Y2=2.34
r73 1 12 300 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.815
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_2%X 1 2 7 10
r16 10 13 54.3016 $w=2.93e-07 $l=1.39e-06 $layer=LI1_cond $X=0.677 $Y=0.42
+ $X2=0.677 $Y2=1.81
r17 7 13 15.6263 $w=2.93e-07 $l=4e-07 $layer=LI1_cond $X=0.677 $Y=2.21 $X2=0.677
+ $Y2=1.81
r18 2 13 300 $w=1.7e-07 $l=3.90832e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.81
r19 1 10 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_2%VGND 1 2 3 10 12 14 16 21 28 29 36 43
r50 43 46 8.41685 $w=5.38e-07 $l=3.8e-07 $layer=LI1_cond $X=2.765 $Y=0 $X2=2.765
+ $Y2=0.38
r51 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r52 36 39 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.185
+ $Y2=0.38
r53 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r54 29 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r55 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r56 26 43 7.6426 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=3.035 $Y=0 $X2=2.765
+ $Y2=0
r57 26 28 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.035 $Y=0 $X2=3.45
+ $Y2=0
r58 25 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r59 25 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r60 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r61 22 36 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.185
+ $Y2=0
r62 22 24 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.61
+ $Y2=0
r63 21 43 7.6426 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=2.495 $Y=0 $X2=2.765
+ $Y2=0
r64 21 24 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.495 $Y=0 $X2=1.61
+ $Y2=0
r65 20 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r66 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r67 17 32 3.93736 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r68 17 19 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r69 16 36 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=1.185
+ $Y2=0
r70 16 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=0.69
+ $Y2=0
r71 14 20 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r72 14 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r73 10 32 3.14078 $w=2.4e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.172 $Y2=0
r74 10 12 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.225 $Y2=0.38
r75 3 46 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.5
+ $Y=0.235 $X2=2.71 $Y2=0.38
r76 2 39 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.235 $X2=1.21 $Y2=0.38
r77 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_2%A_414_47# 1 2 7 10 15
r19 10 12 3.69697 $w=2.08e-07 $l=7e-08 $layer=LI1_cond $X=2.22 $Y=0.66 $X2=2.22
+ $Y2=0.73
r20 8 12 1.31963 $w=1.9e-07 $l=1.05e-07 $layer=LI1_cond $X=2.325 $Y=0.73
+ $X2=2.22 $Y2=0.73
r21 7 15 2.93349 $w=2.73e-07 $l=7e-08 $layer=LI1_cond $X=3.392 $Y=0.73 $X2=3.392
+ $Y2=0.66
r22 7 8 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=3.255 $Y=0.73
+ $X2=2.325 $Y2=0.73
r23 2 15 182 $w=1.7e-07 $l=5.11248e-07 $layer=licon1_NDIFF $count=1 $X=3.18
+ $Y=0.235 $X2=3.37 $Y2=0.66
r24 1 10 182 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.235 $X2=2.21 $Y2=0.66
.ends

