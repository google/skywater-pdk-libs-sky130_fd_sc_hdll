* File: sky130_fd_sc_hdll__inv_1.spice
* Created: Wed Sep  2 08:32:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__inv_1.pex.spice"
.subckt sky130_fd_sc_hdll__inv_1  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.2015 PD=1.82 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1001 N_Y_M1001_d N_A_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.27 PD=2.54 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX2_noxref VNB VPB NWDIODE A=2.8248 P=6.73
*
.include "sky130_fd_sc_hdll__inv_1.pxi.spice"
*
.ends
*
*
