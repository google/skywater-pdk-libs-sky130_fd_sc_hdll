# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__o2bb2ai_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.675000 1.445000 ;
        RECT 0.090000 1.445000 2.145000 1.615000 ;
        RECT 1.765000 1.075000 2.145000 1.445000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.845000 1.075000 1.500000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.650000 1.075000 4.040000 1.445000 ;
        RECT 3.650000 1.445000 5.460000 1.615000 ;
        RECT 5.130000 1.075000 5.460000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.260000 1.075000 4.900000 1.275000 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  0.788000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.895000 0.645000 3.275000 1.075000 ;
        RECT 2.895000 1.075000 3.465000 1.785000 ;
        RECT 2.895000 1.785000 4.680000 1.955000 ;
        RECT 2.895000 1.955000 3.235000 2.465000 ;
        RECT 4.430000 1.955000 4.680000 2.125000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.150000  1.795000 0.400000 2.635000 ;
      RECT 0.195000  0.085000 0.365000 0.895000 ;
      RECT 0.535000  0.305000 1.855000 0.475000 ;
      RECT 0.535000  0.475000 0.835000 0.895000 ;
      RECT 0.625000  1.785000 2.485000 1.965000 ;
      RECT 0.625000  1.965000 0.875000 2.465000 ;
      RECT 1.005000  0.645000 1.385000 0.725000 ;
      RECT 1.005000  0.725000 2.485000 0.905000 ;
      RECT 1.095000  2.135000 1.345000 2.635000 ;
      RECT 2.035000  0.085000 2.205000 0.555000 ;
      RECT 2.035000  2.135000 2.725000 2.635000 ;
      RECT 2.315000  0.905000 2.485000 0.995000 ;
      RECT 2.315000  0.995000 2.725000 1.325000 ;
      RECT 2.315000  1.325000 2.485000 1.785000 ;
      RECT 2.475000  0.255000 3.780000 0.475000 ;
      RECT 2.475000  0.475000 2.725000 0.555000 ;
      RECT 3.455000  2.125000 3.740000 2.635000 ;
      RECT 3.495000  0.475000 3.780000 0.735000 ;
      RECT 3.495000  0.735000 5.660000 0.905000 ;
      RECT 3.960000  2.125000 4.210000 2.295000 ;
      RECT 3.960000  2.295000 5.150000 2.465000 ;
      RECT 4.000000  0.085000 4.170000 0.555000 ;
      RECT 4.340000  0.255000 4.720000 0.725000 ;
      RECT 4.340000  0.725000 5.660000 0.735000 ;
      RECT 4.900000  1.785000 5.150000 2.295000 ;
      RECT 4.940000  0.085000 5.110000 0.555000 ;
      RECT 5.280000  0.255000 5.660000 0.725000 ;
      RECT 5.415000  1.795000 5.620000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o2bb2ai_2
