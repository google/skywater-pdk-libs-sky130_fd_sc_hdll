* File: sky130_fd_sc_hdll__muxb16to1_2.pex.spice
* Created: Wed Sep  2 08:35:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[0] 3 7 11 15 17 27 29
c51 15 0 5.84221e-22 $X=0.965 $Y=1.985
r52 28 29 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.16
+ $X2=0.965 $Y2=1.16
r53 26 28 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=0.75 $Y=1.16 $X2=0.94
+ $Y2=1.16
r54 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.16 $X2=0.75 $Y2=1.16
r55 24 26 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=0.52 $Y=1.16 $X2=0.75
+ $Y2=1.16
r56 23 24 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r57 21 27 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.41 $Y=1.19
+ $X2=0.75 $Y2=1.19
r58 20 23 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=0.41 $Y=1.16
+ $X2=0.495 $Y2=1.16
r59 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r60 17 21 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.23 $Y=1.19
+ $X2=0.41 $Y2=1.19
r61 13 29 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=0.965 $Y=1.295
+ $X2=0.965 $Y2=1.16
r62 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.965 $Y=1.295
+ $X2=0.965 $Y2=1.985
r63 9 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.94 $Y=1.025
+ $X2=0.94 $Y2=1.16
r64 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.94 $Y=1.025
+ $X2=0.94 $Y2=0.56
r65 5 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=1.16
r66 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=0.56
r67 1 23 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=1.16
r68 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[8] 3 7 11 15 17 27 29
c52 15 0 5.84221e-22 $X=0.965 $Y=3.455
r53 28 29 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=4.28
+ $X2=0.965 $Y2=4.28
r54 26 28 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=0.75 $Y=4.28 $X2=0.94
+ $Y2=4.28
r55 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=4.28 $X2=0.75 $Y2=4.28
r56 24 26 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=0.52 $Y=4.28 $X2=0.75
+ $Y2=4.28
r57 23 24 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=4.28
+ $X2=0.52 $Y2=4.28
r58 21 27 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.41 $Y=4.25
+ $X2=0.75 $Y2=4.25
r59 20 23 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=0.41 $Y=4.28
+ $X2=0.495 $Y2=4.28
r60 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=4.28 $X2=0.41 $Y2=4.28
r61 17 21 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.23 $Y=4.25
+ $X2=0.41 $Y2=4.25
r62 13 29 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=0.965 $Y=4.145
+ $X2=0.965 $Y2=4.28
r63 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.965 $Y=4.145
+ $X2=0.965 $Y2=3.455
r64 9 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.94 $Y=4.415
+ $X2=0.94 $Y2=4.28
r65 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.94 $Y=4.415
+ $X2=0.94 $Y2=4.88
r66 5 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.52 $Y=4.415
+ $X2=0.52 $Y2=4.28
r67 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.52 $Y=4.415
+ $X2=0.52 $Y2=4.88
r68 1 23 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=0.495 $Y=4.145
+ $X2=0.495 $Y2=4.28
r69 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.495 $Y=4.145
+ $X2=0.495 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_278_265# 1 2 9 11 12 15 17 18 21 28
+ 32
c84 15 0 8.59607e-20 $X=1.96 $Y=2.075
c85 9 0 2.06539e-19 $X=1.49 $Y=2.075
r86 26 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=2.43 $Y=1.42
+ $X2=2.715 $Y2=1.63
r87 25 32 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=2.265 $Y=1.34
+ $X2=1.96 $Y2=1.34
r88 24 26 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=1.42
+ $X2=2.43 $Y2=1.42
r89 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.265
+ $Y=1.34 $X2=2.265 $Y2=1.34
r90 21 28 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.715 $Y=2.31
+ $X2=2.715 $Y2=1.635
r91 18 26 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.43 $Y=1.205
+ $X2=2.43 $Y2=1.42
r92 17 31 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=2.43 $Y=0.755
+ $X2=2.8 $Y2=0.457
r93 17 18 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.43 $Y=0.755
+ $X2=2.43 $Y2=1.205
r94 13 32 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=1.96 $Y=1.475
+ $X2=1.96 $Y2=1.34
r95 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=1.96 $Y=1.475 $X2=1.96
+ $Y2=2.075
r96 11 32 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=1.87 $Y=1.4
+ $X2=1.96 $Y2=1.34
r97 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.87 $Y=1.4 $X2=1.58
+ $Y2=1.4
r98 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.49 $Y=1.475
+ $X2=1.58 $Y2=1.4
r99 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=1.49 $Y=1.475 $X2=1.49
+ $Y2=2.075
r100 2 28 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.59
+ $Y=1.485 $X2=2.715 $Y2=1.63
r101 2 21 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=2.59
+ $Y=1.485 $X2=2.715 $Y2=2.31
r102 1 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=2.675
+ $Y=0.235 $X2=2.8 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_278_793# 1 2 9 11 12 15 18 19 21 32
c79 15 0 8.62217e-20 $X=1.96 $Y=3.365
c80 9 0 1.91829e-19 $X=1.49 $Y=3.365
r81 25 32 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=2.265 $Y=4.1
+ $X2=1.96 $Y2=4.1
r82 24 26 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=4.02
+ $X2=2.43 $Y2=4.02
r83 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.265
+ $Y=4.1 $X2=2.265 $Y2=4.1
r84 19 26 13.4767 $w=2.58e-07 $l=3.77492e-07 $layer=LI1_cond $X=2.715 $Y=3.805
+ $X2=2.43 $Y2=4.02
r85 19 21 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.715 $Y=3.805
+ $X2=2.715 $Y2=3.13
r86 18 31 16.1792 $w=2.79e-07 $l=4.9678e-07 $layer=LI1_cond $X=2.43 $Y=4.685
+ $X2=2.8 $Y2=4.982
r87 17 26 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.43 $Y=4.235
+ $X2=2.43 $Y2=4.02
r88 17 18 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.43 $Y=4.235
+ $X2=2.43 $Y2=4.685
r89 13 32 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=1.96 $Y=3.965
+ $X2=1.96 $Y2=4.1
r90 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=1.96 $Y=3.965 $X2=1.96
+ $Y2=3.365
r91 11 32 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=1.87 $Y=4.04
+ $X2=1.96 $Y2=4.1
r92 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.87 $Y=4.04
+ $X2=1.58 $Y2=4.04
r93 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.49 $Y=3.965
+ $X2=1.58 $Y2=4.04
r94 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=1.49 $Y=3.965 $X2=1.49
+ $Y2=3.365
r95 2 19 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.59
+ $Y=2.955 $X2=2.715 $Y2=3.81
r96 2 21 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=2.59
+ $Y=2.955 $X2=2.715 $Y2=3.13
r97 1 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=2.675
+ $Y=4.685 $X2=2.8 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[0] 1 3 4 5 6 8 9 12 13 14 15 17 18
+ 20 21 22
r66 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=2.955 $Y=0.92
+ $X2=2.955 $Y2=1.16
r67 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.955
+ $Y=1.16 $X2=2.955 $Y2=1.16
r68 18 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=3.01 $Y=0.845
+ $X2=2.955 $Y2=0.92
r69 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.01 $Y=0.845
+ $X2=3.01 $Y2=0.495
r70 15 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=2.95 $Y=1.41
+ $X2=2.955 $Y2=1.16
r71 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.95 $Y=1.41
+ $X2=2.95 $Y2=1.985
r72 13 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.82 $Y=0.92
+ $X2=2.955 $Y2=0.92
r73 13 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.82 $Y=0.92
+ $X2=2.44 $Y2=0.92
r74 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.365 $Y=0.845
+ $X2=2.44 $Y2=0.92
r75 11 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.365 $Y=0.255
+ $X2=2.365 $Y2=0.845
r76 10 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.955 $Y=0.18
+ $X2=1.88 $Y2=0.18
r77 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.29 $Y=0.18
+ $X2=2.365 $Y2=0.255
r78 9 10 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.29 $Y=0.18
+ $X2=1.955 $Y2=0.18
r79 6 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.88 $Y=0.255
+ $X2=1.88 $Y2=0.18
r80 6 8 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.88 $Y=0.255 $X2=1.88
+ $Y2=0.605
r81 4 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.805 $Y=0.18
+ $X2=1.88 $Y2=0.18
r82 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.805 $Y=0.18
+ $X2=1.535 $Y2=0.18
r83 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.46 $Y=0.255
+ $X2=1.535 $Y2=0.18
r84 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.46 $Y=0.255 $X2=1.46
+ $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[8] 1 3 4 5 6 8 9 12 13 14 15 17 18
+ 20 21 22
r66 25 27 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=2.955 $Y=4.28
+ $X2=2.955 $Y2=4.52
r67 22 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.955
+ $Y=4.28 $X2=2.955 $Y2=4.28
r68 18 27 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=3.01 $Y=4.595
+ $X2=2.955 $Y2=4.52
r69 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.01 $Y=4.595
+ $X2=3.01 $Y2=4.945
r70 15 25 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=2.95 $Y=4.03
+ $X2=2.955 $Y2=4.28
r71 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.95 $Y=4.03
+ $X2=2.95 $Y2=3.455
r72 13 27 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.82 $Y=4.52
+ $X2=2.955 $Y2=4.52
r73 13 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.82 $Y=4.52
+ $X2=2.44 $Y2=4.52
r74 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.365 $Y=4.595
+ $X2=2.44 $Y2=4.52
r75 11 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.365 $Y=4.595
+ $X2=2.365 $Y2=5.185
r76 10 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.955 $Y=5.26
+ $X2=1.88 $Y2=5.26
r77 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.29 $Y=5.26
+ $X2=2.365 $Y2=5.185
r78 9 10 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.29 $Y=5.26
+ $X2=1.955 $Y2=5.26
r79 6 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.88 $Y=5.185
+ $X2=1.88 $Y2=5.26
r80 6 8 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.88 $Y=5.185 $X2=1.88
+ $Y2=4.835
r81 4 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.805 $Y=5.26
+ $X2=1.88 $Y2=5.26
r82 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.805 $Y=5.26
+ $X2=1.535 $Y2=5.26
r83 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.46 $Y=5.185
+ $X2=1.535 $Y2=5.26
r84 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.46 $Y=5.185 $X2=1.46
+ $Y2=4.835
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[1] 1 3 4 6 7 10 11 12 13 15 16 18 20
+ 21 22
r63 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=3.485 $Y=0.92
+ $X2=3.485 $Y2=1.16
r64 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.485
+ $Y=1.16 $X2=3.485 $Y2=1.16
r65 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.98 $Y=0.255
+ $X2=4.98 $Y2=0.605
r66 17 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.635 $Y=0.18
+ $X2=4.56 $Y2=0.18
r67 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.905 $Y=0.18
+ $X2=4.98 $Y2=0.255
r68 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.905 $Y=0.18
+ $X2=4.635 $Y2=0.18
r69 13 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.56 $Y=0.255
+ $X2=4.56 $Y2=0.18
r70 13 15 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.56 $Y=0.255
+ $X2=4.56 $Y2=0.605
r71 11 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.485 $Y=0.18
+ $X2=4.56 $Y2=0.18
r72 11 12 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=4.485 $Y=0.18
+ $X2=4.15 $Y2=0.18
r73 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.075 $Y=0.255
+ $X2=4.15 $Y2=0.18
r74 9 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=4.075 $Y=0.255
+ $X2=4.075 $Y2=0.845
r75 8 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.62 $Y=0.92
+ $X2=3.485 $Y2=0.92
r76 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4 $Y=0.92
+ $X2=4.075 $Y2=0.845
r77 7 8 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=4 $Y=0.92 $X2=3.62
+ $Y2=0.92
r78 4 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=3.49 $Y=1.41
+ $X2=3.485 $Y2=1.16
r79 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.49 $Y=1.41 $X2=3.49
+ $Y2=1.985
r80 1 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=3.43 $Y=0.845
+ $X2=3.485 $Y2=0.92
r81 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.43 $Y=0.845 $X2=3.43
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[9] 1 3 4 6 7 10 11 12 13 15 16 18 20
+ 21 22
r66 25 27 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=3.485 $Y=4.28
+ $X2=3.485 $Y2=4.52
r67 22 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.485
+ $Y=4.28 $X2=3.485 $Y2=4.28
r68 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.98 $Y=5.185
+ $X2=4.98 $Y2=4.835
r69 17 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.635 $Y=5.26
+ $X2=4.56 $Y2=5.26
r70 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.905 $Y=5.26
+ $X2=4.98 $Y2=5.185
r71 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.905 $Y=5.26
+ $X2=4.635 $Y2=5.26
r72 13 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.56 $Y=5.185
+ $X2=4.56 $Y2=5.26
r73 13 15 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.56 $Y=5.185
+ $X2=4.56 $Y2=4.835
r74 11 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.485 $Y=5.26
+ $X2=4.56 $Y2=5.26
r75 11 12 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=4.485 $Y=5.26
+ $X2=4.15 $Y2=5.26
r76 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.075 $Y=5.185
+ $X2=4.15 $Y2=5.26
r77 9 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=4.075 $Y=4.595
+ $X2=4.075 $Y2=5.185
r78 8 27 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.62 $Y=4.52
+ $X2=3.485 $Y2=4.52
r79 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4 $Y=4.52
+ $X2=4.075 $Y2=4.595
r80 7 8 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=4 $Y=4.52 $X2=3.62
+ $Y2=4.52
r81 4 25 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=3.49 $Y=4.03
+ $X2=3.485 $Y2=4.28
r82 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.49 $Y=4.03 $X2=3.49
+ $Y2=3.455
r83 1 27 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=3.43 $Y=4.595
+ $X2=3.485 $Y2=4.52
r84 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.43 $Y=4.595 $X2=3.43
+ $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_701_47# 1 2 9 11 12 15 19 22 24 28
c81 15 0 2.06539e-19 $X=4.95 $Y=2.075
c82 11 0 1.93373e-19 $X=4.86 $Y=1.4
c83 9 0 8.59607e-20 $X=4.48 $Y=2.075
r84 31 33 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=4.175 $Y=1.34
+ $X2=4.48 $Y2=1.34
r85 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.175
+ $Y=1.34 $X2=4.175 $Y2=1.34
r86 28 30 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.01 $Y=1.42
+ $X2=4.175 $Y2=1.42
r87 27 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=3.725 $Y=1.63
+ $X2=4.01 $Y2=1.42
r88 22 28 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=4.01 $Y=1.205
+ $X2=4.01 $Y2=1.42
r89 21 24 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=4.01 $Y=0.755
+ $X2=3.64 $Y2=0.457
r90 21 22 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.01 $Y=0.755
+ $X2=4.01 $Y2=1.205
r91 19 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.725 $Y=2.31
+ $X2=3.725 $Y2=1.635
r92 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=4.95 $Y=1.475 $X2=4.95
+ $Y2=2.075
r93 12 33 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=4.57 $Y=1.4
+ $X2=4.48 $Y2=1.34
r94 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.86 $Y=1.4
+ $X2=4.95 $Y2=1.475
r95 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.86 $Y=1.4 $X2=4.57
+ $Y2=1.4
r96 7 33 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=4.48 $Y=1.475
+ $X2=4.48 $Y2=1.34
r97 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=4.48 $Y=1.475 $X2=4.48
+ $Y2=2.075
r98 2 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=1.485 $X2=3.725 $Y2=1.63
r99 2 19 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=1.485 $X2=3.725 $Y2=2.31
r100 1 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=3.505
+ $Y=0.235 $X2=3.64 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_701_937# 1 2 9 11 12 15 19 22 24 28
c81 15 0 1.91829e-19 $X=4.95 $Y=3.365
c82 11 0 1.93373e-19 $X=4.86 $Y=4.04
c83 9 0 8.62217e-20 $X=4.48 $Y=3.365
r84 31 33 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=4.175 $Y=4.1
+ $X2=4.48 $Y2=4.1
r85 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.175
+ $Y=4.1 $X2=4.175 $Y2=4.1
r86 28 30 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.01 $Y=4.02
+ $X2=4.175 $Y2=4.02
r87 22 24 16.1792 $w=2.79e-07 $l=4.9678e-07 $layer=LI1_cond $X=4.01 $Y=4.685
+ $X2=3.64 $Y2=4.982
r88 21 28 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=4.01 $Y=4.235
+ $X2=4.01 $Y2=4.02
r89 21 22 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.01 $Y=4.235
+ $X2=4.01 $Y2=4.685
r90 17 28 13.4767 $w=2.58e-07 $l=3.77492e-07 $layer=LI1_cond $X=3.725 $Y=3.805
+ $X2=4.01 $Y2=4.02
r91 17 19 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.725 $Y=3.805
+ $X2=3.725 $Y2=3.13
r92 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=4.95 $Y=3.965 $X2=4.95
+ $Y2=3.365
r93 12 33 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=4.57 $Y=4.04
+ $X2=4.48 $Y2=4.1
r94 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.86 $Y=4.04
+ $X2=4.95 $Y2=3.965
r95 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.86 $Y=4.04
+ $X2=4.57 $Y2=4.04
r96 7 33 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=4.48 $Y=3.965
+ $X2=4.48 $Y2=4.1
r97 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=4.48 $Y=3.965 $X2=4.48
+ $Y2=3.365
r98 2 17 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=2.955 $X2=3.725 $Y2=3.81
r99 2 19 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=2.955 $X2=3.725 $Y2=3.13
r100 1 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=3.505
+ $Y=4.685 $X2=3.64 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[1] 3 7 11 15 17 28
c57 17 0 1.17966e-19 $X=6.21 $Y=1.19
c58 15 0 1.17966e-19 $X=5.945 $Y=1.985
c59 3 0 5.84221e-22 $X=5.475 $Y=1.985
r60 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.03
+ $Y=1.16 $X2=6.03 $Y2=1.16
r61 26 28 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=5.945 $Y=1.16
+ $X2=6.03 $Y2=1.16
r62 25 26 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.92 $Y=1.16
+ $X2=5.945 $Y2=1.16
r63 24 29 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.69 $Y=1.19
+ $X2=6.03 $Y2=1.19
r64 23 25 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=5.69 $Y=1.16 $X2=5.92
+ $Y2=1.16
r65 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.69
+ $Y=1.16 $X2=5.69 $Y2=1.16
r66 21 23 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=5.5 $Y=1.16 $X2=5.69
+ $Y2=1.16
r67 19 21 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.475 $Y=1.16
+ $X2=5.5 $Y2=1.16
r68 17 29 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.21 $Y=1.19
+ $X2=6.03 $Y2=1.19
r69 13 26 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.945 $Y=1.295
+ $X2=5.945 $Y2=1.16
r70 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=5.945 $Y=1.295
+ $X2=5.945 $Y2=1.985
r71 9 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.92 $Y=1.025
+ $X2=5.92 $Y2=1.16
r72 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.92 $Y=1.025
+ $X2=5.92 $Y2=0.56
r73 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.5 $Y=1.025 $X2=5.5
+ $Y2=1.16
r74 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.5 $Y=1.025 $X2=5.5
+ $Y2=0.56
r75 1 19 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.475 $Y=1.295
+ $X2=5.475 $Y2=1.16
r76 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=5.475 $Y=1.295
+ $X2=5.475 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[9] 3 7 11 15 17 28
c57 17 0 1.17966e-19 $X=6.21 $Y=4.25
c58 15 0 1.17966e-19 $X=5.945 $Y=3.455
c59 3 0 5.84221e-22 $X=5.475 $Y=3.455
r60 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.03
+ $Y=4.28 $X2=6.03 $Y2=4.28
r61 26 28 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=5.945 $Y=4.28
+ $X2=6.03 $Y2=4.28
r62 25 26 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.92 $Y=4.28
+ $X2=5.945 $Y2=4.28
r63 24 29 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.69 $Y=4.25
+ $X2=6.03 $Y2=4.25
r64 23 25 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=5.69 $Y=4.28 $X2=5.92
+ $Y2=4.28
r65 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.69
+ $Y=4.28 $X2=5.69 $Y2=4.28
r66 21 23 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=5.5 $Y=4.28 $X2=5.69
+ $Y2=4.28
r67 19 21 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.475 $Y=4.28
+ $X2=5.5 $Y2=4.28
r68 17 29 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.21 $Y=4.25
+ $X2=6.03 $Y2=4.25
r69 13 26 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.945 $Y=4.145
+ $X2=5.945 $Y2=4.28
r70 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=5.945 $Y=4.145
+ $X2=5.945 $Y2=3.455
r71 9 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.92 $Y=4.415
+ $X2=5.92 $Y2=4.28
r72 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.92 $Y=4.415
+ $X2=5.92 $Y2=4.88
r73 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.5 $Y=4.415 $X2=5.5
+ $Y2=4.28
r74 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.5 $Y=4.415 $X2=5.5
+ $Y2=4.88
r75 1 19 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.475 $Y=4.145
+ $X2=5.475 $Y2=4.28
r76 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=5.475 $Y=4.145
+ $X2=5.475 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[2] 3 7 11 15 17 27 29
c58 27 0 1.17966e-19 $X=7.19 $Y=1.16
c59 15 0 5.84221e-22 $X=7.405 $Y=1.985
c60 3 0 1.17966e-19 $X=6.935 $Y=1.985
r61 28 29 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=7.38 $Y=1.16
+ $X2=7.405 $Y2=1.16
r62 26 28 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=7.19 $Y=1.16 $X2=7.38
+ $Y2=1.16
r63 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.19
+ $Y=1.16 $X2=7.19 $Y2=1.16
r64 24 26 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=6.96 $Y=1.16 $X2=7.19
+ $Y2=1.16
r65 23 24 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=6.935 $Y=1.16
+ $X2=6.96 $Y2=1.16
r66 21 27 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.85 $Y=1.19
+ $X2=7.19 $Y2=1.19
r67 20 23 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=6.85 $Y=1.16
+ $X2=6.935 $Y2=1.16
r68 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.85
+ $Y=1.16 $X2=6.85 $Y2=1.16
r69 17 21 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.67 $Y=1.19
+ $X2=6.85 $Y2=1.19
r70 13 29 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=7.405 $Y=1.295
+ $X2=7.405 $Y2=1.16
r71 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=7.405 $Y=1.295
+ $X2=7.405 $Y2=1.985
r72 9 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.38 $Y=1.025
+ $X2=7.38 $Y2=1.16
r73 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.38 $Y=1.025
+ $X2=7.38 $Y2=0.56
r74 5 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.96 $Y=1.025
+ $X2=6.96 $Y2=1.16
r75 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.96 $Y=1.025
+ $X2=6.96 $Y2=0.56
r76 1 23 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=6.935 $Y=1.295
+ $X2=6.935 $Y2=1.16
r77 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=6.935 $Y=1.295
+ $X2=6.935 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[10] 3 7 11 15 17 27 29
c59 27 0 1.17966e-19 $X=7.19 $Y=4.28
c60 15 0 5.84221e-22 $X=7.405 $Y=3.455
c61 3 0 1.17966e-19 $X=6.935 $Y=3.455
r62 28 29 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=7.38 $Y=4.28
+ $X2=7.405 $Y2=4.28
r63 26 28 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=7.19 $Y=4.28 $X2=7.38
+ $Y2=4.28
r64 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.19
+ $Y=4.28 $X2=7.19 $Y2=4.28
r65 24 26 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=6.96 $Y=4.28 $X2=7.19
+ $Y2=4.28
r66 23 24 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=6.935 $Y=4.28
+ $X2=6.96 $Y2=4.28
r67 21 27 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.85 $Y=4.25
+ $X2=7.19 $Y2=4.25
r68 20 23 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=6.85 $Y=4.28
+ $X2=6.935 $Y2=4.28
r69 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.85
+ $Y=4.28 $X2=6.85 $Y2=4.28
r70 17 21 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.67 $Y=4.25
+ $X2=6.85 $Y2=4.25
r71 13 29 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=7.405 $Y=4.145
+ $X2=7.405 $Y2=4.28
r72 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=7.405 $Y=4.145
+ $X2=7.405 $Y2=3.455
r73 9 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.38 $Y=4.415
+ $X2=7.38 $Y2=4.28
r74 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.38 $Y=4.415
+ $X2=7.38 $Y2=4.88
r75 5 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.96 $Y=4.415
+ $X2=6.96 $Y2=4.28
r76 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.96 $Y=4.415
+ $X2=6.96 $Y2=4.88
r77 1 23 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=6.935 $Y=4.145
+ $X2=6.935 $Y2=4.28
r78 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=6.935 $Y=4.145
+ $X2=6.935 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1566_265# 1 2 9 11 12 15 17 18 21 28
+ 32
c85 15 0 8.59607e-20 $X=8.4 $Y=2.075
c86 12 0 1.93373e-19 $X=8.02 $Y=1.4
c87 9 0 2.06539e-19 $X=7.93 $Y=2.075
r88 26 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=8.87 $Y=1.42
+ $X2=9.155 $Y2=1.63
r89 25 32 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=8.705 $Y=1.34
+ $X2=8.4 $Y2=1.34
r90 24 26 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=8.705 $Y=1.42
+ $X2=8.87 $Y2=1.42
r91 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.705
+ $Y=1.34 $X2=8.705 $Y2=1.34
r92 21 28 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=9.155 $Y=2.31
+ $X2=9.155 $Y2=1.635
r93 18 26 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=8.87 $Y=1.205
+ $X2=8.87 $Y2=1.42
r94 17 31 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=8.87 $Y=0.755
+ $X2=9.24 $Y2=0.457
r95 17 18 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.87 $Y=0.755
+ $X2=8.87 $Y2=1.205
r96 13 32 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=8.4 $Y=1.475
+ $X2=8.4 $Y2=1.34
r97 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=8.4 $Y=1.475 $X2=8.4
+ $Y2=2.075
r98 11 32 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=8.31 $Y=1.4
+ $X2=8.4 $Y2=1.34
r99 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.31 $Y=1.4 $X2=8.02
+ $Y2=1.4
r100 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=7.93 $Y=1.475
+ $X2=8.02 $Y2=1.4
r101 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=7.93 $Y=1.475 $X2=7.93
+ $Y2=2.075
r102 2 28 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=9.03
+ $Y=1.485 $X2=9.155 $Y2=1.63
r103 2 21 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=9.03
+ $Y=1.485 $X2=9.155 $Y2=2.31
r104 1 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=9.115
+ $Y=0.235 $X2=9.24 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1566_793# 1 2 9 11 12 15 18 19 21 32
c80 15 0 8.62217e-20 $X=8.4 $Y=3.365
c81 12 0 1.93373e-19 $X=8.02 $Y=4.04
c82 9 0 1.91829e-19 $X=7.93 $Y=3.365
r83 25 32 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=8.705 $Y=4.1
+ $X2=8.4 $Y2=4.1
r84 24 26 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=8.705 $Y=4.02
+ $X2=8.87 $Y2=4.02
r85 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.705
+ $Y=4.1 $X2=8.705 $Y2=4.1
r86 19 26 13.4767 $w=2.58e-07 $l=3.77492e-07 $layer=LI1_cond $X=9.155 $Y=3.805
+ $X2=8.87 $Y2=4.02
r87 19 21 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=9.155 $Y=3.805
+ $X2=9.155 $Y2=3.13
r88 18 31 16.1792 $w=2.79e-07 $l=4.9678e-07 $layer=LI1_cond $X=8.87 $Y=4.685
+ $X2=9.24 $Y2=4.982
r89 17 26 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=8.87 $Y=4.235
+ $X2=8.87 $Y2=4.02
r90 17 18 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.87 $Y=4.235
+ $X2=8.87 $Y2=4.685
r91 13 32 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=8.4 $Y=3.965
+ $X2=8.4 $Y2=4.1
r92 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=8.4 $Y=3.965 $X2=8.4
+ $Y2=3.365
r93 11 32 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=8.31 $Y=4.04
+ $X2=8.4 $Y2=4.1
r94 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.31 $Y=4.04
+ $X2=8.02 $Y2=4.04
r95 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=7.93 $Y=3.965
+ $X2=8.02 $Y2=4.04
r96 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=7.93 $Y=3.965 $X2=7.93
+ $Y2=3.365
r97 2 19 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=9.03
+ $Y=2.955 $X2=9.155 $Y2=3.81
r98 2 21 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=9.03
+ $Y=2.955 $X2=9.155 $Y2=3.13
r99 1 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=9.115
+ $Y=4.685 $X2=9.24 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[2] 1 3 4 5 6 8 9 12 13 14 15 17 18
+ 20 21 22
r66 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=9.395 $Y=0.92
+ $X2=9.395 $Y2=1.16
r67 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.395
+ $Y=1.16 $X2=9.395 $Y2=1.16
r68 18 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=9.45 $Y=0.845
+ $X2=9.395 $Y2=0.92
r69 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.45 $Y=0.845
+ $X2=9.45 $Y2=0.495
r70 15 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=9.39 $Y=1.41
+ $X2=9.395 $Y2=1.16
r71 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.39 $Y=1.41
+ $X2=9.39 $Y2=1.985
r72 13 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.26 $Y=0.92
+ $X2=9.395 $Y2=0.92
r73 13 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=9.26 $Y=0.92
+ $X2=8.88 $Y2=0.92
r74 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.805 $Y=0.845
+ $X2=8.88 $Y2=0.92
r75 11 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=8.805 $Y=0.255
+ $X2=8.805 $Y2=0.845
r76 10 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.395 $Y=0.18
+ $X2=8.32 $Y2=0.18
r77 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.73 $Y=0.18
+ $X2=8.805 $Y2=0.255
r78 9 10 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=8.73 $Y=0.18
+ $X2=8.395 $Y2=0.18
r79 6 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.32 $Y=0.255
+ $X2=8.32 $Y2=0.18
r80 6 8 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=8.32 $Y=0.255 $X2=8.32
+ $Y2=0.605
r81 4 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.245 $Y=0.18
+ $X2=8.32 $Y2=0.18
r82 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.245 $Y=0.18
+ $X2=7.975 $Y2=0.18
r83 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.9 $Y=0.255
+ $X2=7.975 $Y2=0.18
r84 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=7.9 $Y=0.255 $X2=7.9
+ $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[10] 1 3 4 5 6 8 9 12 13 14 15 17 18
+ 20 21 22
r66 25 27 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=9.395 $Y=4.28
+ $X2=9.395 $Y2=4.52
r67 22 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.395
+ $Y=4.28 $X2=9.395 $Y2=4.28
r68 18 27 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=9.45 $Y=4.595
+ $X2=9.395 $Y2=4.52
r69 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.45 $Y=4.595
+ $X2=9.45 $Y2=4.945
r70 15 25 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=9.39 $Y=4.03
+ $X2=9.395 $Y2=4.28
r71 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.39 $Y=4.03
+ $X2=9.39 $Y2=3.455
r72 13 27 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.26 $Y=4.52
+ $X2=9.395 $Y2=4.52
r73 13 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=9.26 $Y=4.52
+ $X2=8.88 $Y2=4.52
r74 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.805 $Y=4.595
+ $X2=8.88 $Y2=4.52
r75 11 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=8.805 $Y=4.595
+ $X2=8.805 $Y2=5.185
r76 10 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.395 $Y=5.26
+ $X2=8.32 $Y2=5.26
r77 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.73 $Y=5.26
+ $X2=8.805 $Y2=5.185
r78 9 10 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=8.73 $Y=5.26
+ $X2=8.395 $Y2=5.26
r79 6 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.32 $Y=5.185
+ $X2=8.32 $Y2=5.26
r80 6 8 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=8.32 $Y=5.185 $X2=8.32
+ $Y2=4.835
r81 4 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.245 $Y=5.26
+ $X2=8.32 $Y2=5.26
r82 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.245 $Y=5.26
+ $X2=7.975 $Y2=5.26
r83 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.9 $Y=5.185
+ $X2=7.975 $Y2=5.26
r84 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=7.9 $Y=5.185 $X2=7.9
+ $Y2=4.835
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[3] 1 3 4 6 7 10 11 12 13 15 16 18 20
+ 21 22
r63 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=9.925 $Y=0.92
+ $X2=9.925 $Y2=1.16
r64 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.925
+ $Y=1.16 $X2=9.925 $Y2=1.16
r65 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=11.42 $Y=0.255
+ $X2=11.42 $Y2=0.605
r66 17 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.075 $Y=0.18
+ $X2=11 $Y2=0.18
r67 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.345 $Y=0.18
+ $X2=11.42 $Y2=0.255
r68 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=11.345 $Y=0.18
+ $X2=11.075 $Y2=0.18
r69 13 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11 $Y=0.255 $X2=11
+ $Y2=0.18
r70 13 15 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=11 $Y=0.255 $X2=11
+ $Y2=0.605
r71 11 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.925 $Y=0.18
+ $X2=11 $Y2=0.18
r72 11 12 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.925 $Y=0.18
+ $X2=10.59 $Y2=0.18
r73 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.515 $Y=0.255
+ $X2=10.59 $Y2=0.18
r74 9 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=10.515 $Y=0.255
+ $X2=10.515 $Y2=0.845
r75 8 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.06 $Y=0.92
+ $X2=9.925 $Y2=0.92
r76 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.44 $Y=0.92
+ $X2=10.515 $Y2=0.845
r77 7 8 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=10.44 $Y=0.92
+ $X2=10.06 $Y2=0.92
r78 4 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=9.93 $Y=1.41
+ $X2=9.925 $Y2=1.16
r79 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.93 $Y=1.41 $X2=9.93
+ $Y2=1.985
r80 1 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=9.87 $Y=0.845
+ $X2=9.925 $Y2=0.92
r81 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.87 $Y=0.845 $X2=9.87
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[11] 1 3 4 6 7 10 11 12 13 15 16 18
+ 20 21 22
r66 25 27 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=9.925 $Y=4.28
+ $X2=9.925 $Y2=4.52
r67 22 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.925
+ $Y=4.28 $X2=9.925 $Y2=4.28
r68 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=11.42 $Y=5.185
+ $X2=11.42 $Y2=4.835
r69 17 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.075 $Y=5.26
+ $X2=11 $Y2=5.26
r70 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.345 $Y=5.26
+ $X2=11.42 $Y2=5.185
r71 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=11.345 $Y=5.26
+ $X2=11.075 $Y2=5.26
r72 13 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11 $Y=5.185 $X2=11
+ $Y2=5.26
r73 13 15 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=11 $Y=5.185 $X2=11
+ $Y2=4.835
r74 11 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.925 $Y=5.26
+ $X2=11 $Y2=5.26
r75 11 12 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.925 $Y=5.26
+ $X2=10.59 $Y2=5.26
r76 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.515 $Y=5.185
+ $X2=10.59 $Y2=5.26
r77 9 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=10.515 $Y=4.595
+ $X2=10.515 $Y2=5.185
r78 8 27 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.06 $Y=4.52
+ $X2=9.925 $Y2=4.52
r79 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.44 $Y=4.52
+ $X2=10.515 $Y2=4.595
r80 7 8 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=10.44 $Y=4.52
+ $X2=10.06 $Y2=4.52
r81 4 25 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=9.93 $Y=4.03
+ $X2=9.925 $Y2=4.28
r82 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.93 $Y=4.03 $X2=9.93
+ $Y2=3.455
r83 1 27 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=9.87 $Y=4.595
+ $X2=9.925 $Y2=4.52
r84 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.87 $Y=4.595 $X2=9.87
+ $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1989_47# 1 2 9 11 12 15 19 22 24 28
c81 15 0 2.06539e-19 $X=11.39 $Y=2.075
c82 11 0 1.93373e-19 $X=11.3 $Y=1.4
c83 9 0 8.59607e-20 $X=10.92 $Y=2.075
r84 31 33 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=10.615 $Y=1.34
+ $X2=10.92 $Y2=1.34
r85 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.615
+ $Y=1.34 $X2=10.615 $Y2=1.34
r86 28 30 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=10.45 $Y=1.42
+ $X2=10.615 $Y2=1.42
r87 27 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=10.165 $Y=1.63
+ $X2=10.45 $Y2=1.42
r88 22 28 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=10.45 $Y=1.205
+ $X2=10.45 $Y2=1.42
r89 21 24 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=10.45 $Y=0.755
+ $X2=10.08 $Y2=0.457
r90 21 22 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=10.45 $Y=0.755
+ $X2=10.45 $Y2=1.205
r91 19 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=10.165 $Y=2.31
+ $X2=10.165 $Y2=1.635
r92 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=11.39 $Y=1.475
+ $X2=11.39 $Y2=2.075
r93 12 33 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=11.01 $Y=1.4
+ $X2=10.92 $Y2=1.34
r94 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=11.3 $Y=1.4
+ $X2=11.39 $Y2=1.475
r95 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=11.3 $Y=1.4
+ $X2=11.01 $Y2=1.4
r96 7 33 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=10.92 $Y=1.475
+ $X2=10.92 $Y2=1.34
r97 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=10.92 $Y=1.475 $X2=10.92
+ $Y2=2.075
r98 2 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.02
+ $Y=1.485 $X2=10.165 $Y2=1.63
r99 2 19 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=10.02
+ $Y=1.485 $X2=10.165 $Y2=2.31
r100 1 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=9.945
+ $Y=0.235 $X2=10.08 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1989_937# 1 2 9 11 12 15 19 22 24 28
c81 15 0 1.91829e-19 $X=11.39 $Y=3.365
c82 11 0 1.93373e-19 $X=11.3 $Y=4.04
c83 9 0 8.62217e-20 $X=10.92 $Y=3.365
r84 31 33 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=10.615 $Y=4.1
+ $X2=10.92 $Y2=4.1
r85 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.615
+ $Y=4.1 $X2=10.615 $Y2=4.1
r86 28 30 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=10.45 $Y=4.02
+ $X2=10.615 $Y2=4.02
r87 22 24 16.1792 $w=2.79e-07 $l=4.9678e-07 $layer=LI1_cond $X=10.45 $Y=4.685
+ $X2=10.08 $Y2=4.982
r88 21 28 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=10.45 $Y=4.235
+ $X2=10.45 $Y2=4.02
r89 21 22 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=10.45 $Y=4.235
+ $X2=10.45 $Y2=4.685
r90 17 28 13.4767 $w=2.58e-07 $l=3.77492e-07 $layer=LI1_cond $X=10.165 $Y=3.805
+ $X2=10.45 $Y2=4.02
r91 17 19 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=10.165 $Y=3.805
+ $X2=10.165 $Y2=3.13
r92 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=11.39 $Y=3.965
+ $X2=11.39 $Y2=3.365
r93 12 33 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=11.01 $Y=4.04
+ $X2=10.92 $Y2=4.1
r94 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=11.3 $Y=4.04
+ $X2=11.39 $Y2=3.965
r95 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=11.3 $Y=4.04
+ $X2=11.01 $Y2=4.04
r96 7 33 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=10.92 $Y=3.965
+ $X2=10.92 $Y2=4.1
r97 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=10.92 $Y=3.965 $X2=10.92
+ $Y2=3.365
r98 2 17 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.02
+ $Y=2.955 $X2=10.165 $Y2=3.81
r99 2 19 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=10.02
+ $Y=2.955 $X2=10.165 $Y2=3.13
r100 1 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=9.945
+ $Y=4.685 $X2=10.08 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[3] 3 7 11 15 17 28
c57 17 0 1.17966e-19 $X=12.65 $Y=1.19
c58 15 0 1.17966e-19 $X=12.385 $Y=1.985
c59 3 0 5.84221e-22 $X=11.915 $Y=1.985
r60 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.47
+ $Y=1.16 $X2=12.47 $Y2=1.16
r61 26 28 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=12.385 $Y=1.16
+ $X2=12.47 $Y2=1.16
r62 25 26 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=12.36 $Y=1.16
+ $X2=12.385 $Y2=1.16
r63 24 29 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=12.13 $Y=1.19
+ $X2=12.47 $Y2=1.19
r64 23 25 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=12.13 $Y=1.16 $X2=12.36
+ $Y2=1.16
r65 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.13
+ $Y=1.16 $X2=12.13 $Y2=1.16
r66 21 23 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=11.94 $Y=1.16
+ $X2=12.13 $Y2=1.16
r67 19 21 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=11.915 $Y=1.16
+ $X2=11.94 $Y2=1.16
r68 17 29 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=12.65 $Y=1.19
+ $X2=12.47 $Y2=1.19
r69 13 26 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=12.385 $Y=1.295
+ $X2=12.385 $Y2=1.16
r70 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=12.385 $Y=1.295
+ $X2=12.385 $Y2=1.985
r71 9 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=12.36 $Y=1.025
+ $X2=12.36 $Y2=1.16
r72 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=12.36 $Y=1.025
+ $X2=12.36 $Y2=0.56
r73 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.94 $Y=1.025
+ $X2=11.94 $Y2=1.16
r74 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.94 $Y=1.025
+ $X2=11.94 $Y2=0.56
r75 1 19 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=11.915 $Y=1.295
+ $X2=11.915 $Y2=1.16
r76 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=11.915 $Y=1.295
+ $X2=11.915 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[11] 3 7 11 15 17 28
c57 17 0 1.17966e-19 $X=12.65 $Y=4.25
c58 15 0 1.17966e-19 $X=12.385 $Y=3.455
c59 3 0 5.84221e-22 $X=11.915 $Y=3.455
r60 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.47
+ $Y=4.28 $X2=12.47 $Y2=4.28
r61 26 28 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=12.385 $Y=4.28
+ $X2=12.47 $Y2=4.28
r62 25 26 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=12.36 $Y=4.28
+ $X2=12.385 $Y2=4.28
r63 24 29 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=12.13 $Y=4.25
+ $X2=12.47 $Y2=4.25
r64 23 25 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=12.13 $Y=4.28 $X2=12.36
+ $Y2=4.28
r65 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.13
+ $Y=4.28 $X2=12.13 $Y2=4.28
r66 21 23 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=11.94 $Y=4.28
+ $X2=12.13 $Y2=4.28
r67 19 21 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=11.915 $Y=4.28
+ $X2=11.94 $Y2=4.28
r68 17 29 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=12.65 $Y=4.25
+ $X2=12.47 $Y2=4.25
r69 13 26 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=12.385 $Y=4.145
+ $X2=12.385 $Y2=4.28
r70 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=12.385 $Y=4.145
+ $X2=12.385 $Y2=3.455
r71 9 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=12.36 $Y=4.415
+ $X2=12.36 $Y2=4.28
r72 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=12.36 $Y=4.415
+ $X2=12.36 $Y2=4.88
r73 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.94 $Y=4.415
+ $X2=11.94 $Y2=4.28
r74 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.94 $Y=4.415
+ $X2=11.94 $Y2=4.88
r75 1 19 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=11.915 $Y=4.145
+ $X2=11.915 $Y2=4.28
r76 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=11.915 $Y=4.145
+ $X2=11.915 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[4] 3 7 11 15 17 27 29
c58 27 0 1.17966e-19 $X=13.63 $Y=1.16
c59 15 0 5.84221e-22 $X=13.845 $Y=1.985
c60 3 0 1.17966e-19 $X=13.375 $Y=1.985
r61 28 29 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=13.82 $Y=1.16
+ $X2=13.845 $Y2=1.16
r62 26 28 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=13.63 $Y=1.16
+ $X2=13.82 $Y2=1.16
r63 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.63
+ $Y=1.16 $X2=13.63 $Y2=1.16
r64 24 26 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=13.4 $Y=1.16 $X2=13.63
+ $Y2=1.16
r65 23 24 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=13.375 $Y=1.16
+ $X2=13.4 $Y2=1.16
r66 21 27 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=13.29 $Y=1.19
+ $X2=13.63 $Y2=1.19
r67 20 23 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=13.29 $Y=1.16
+ $X2=13.375 $Y2=1.16
r68 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.29
+ $Y=1.16 $X2=13.29 $Y2=1.16
r69 17 21 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=13.11 $Y=1.19
+ $X2=13.29 $Y2=1.19
r70 13 29 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=13.845 $Y=1.295
+ $X2=13.845 $Y2=1.16
r71 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=13.845 $Y=1.295
+ $X2=13.845 $Y2=1.985
r72 9 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.82 $Y=1.025
+ $X2=13.82 $Y2=1.16
r73 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=13.82 $Y=1.025
+ $X2=13.82 $Y2=0.56
r74 5 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.4 $Y=1.025
+ $X2=13.4 $Y2=1.16
r75 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=13.4 $Y=1.025
+ $X2=13.4 $Y2=0.56
r76 1 23 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=13.375 $Y=1.295
+ $X2=13.375 $Y2=1.16
r77 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=13.375 $Y=1.295
+ $X2=13.375 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[12] 3 7 11 15 17 27 29
c59 27 0 1.17966e-19 $X=13.63 $Y=4.28
c60 15 0 5.84221e-22 $X=13.845 $Y=3.455
c61 3 0 1.17966e-19 $X=13.375 $Y=3.455
r62 28 29 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=13.82 $Y=4.28
+ $X2=13.845 $Y2=4.28
r63 26 28 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=13.63 $Y=4.28
+ $X2=13.82 $Y2=4.28
r64 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.63
+ $Y=4.28 $X2=13.63 $Y2=4.28
r65 24 26 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=13.4 $Y=4.28 $X2=13.63
+ $Y2=4.28
r66 23 24 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=13.375 $Y=4.28
+ $X2=13.4 $Y2=4.28
r67 21 27 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=13.29 $Y=4.25
+ $X2=13.63 $Y2=4.25
r68 20 23 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=13.29 $Y=4.28
+ $X2=13.375 $Y2=4.28
r69 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.29
+ $Y=4.28 $X2=13.29 $Y2=4.28
r70 17 21 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=13.11 $Y=4.25
+ $X2=13.29 $Y2=4.25
r71 13 29 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=13.845 $Y=4.145
+ $X2=13.845 $Y2=4.28
r72 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=13.845 $Y=4.145
+ $X2=13.845 $Y2=3.455
r73 9 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.82 $Y=4.415
+ $X2=13.82 $Y2=4.28
r74 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=13.82 $Y=4.415
+ $X2=13.82 $Y2=4.88
r75 5 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.4 $Y=4.415
+ $X2=13.4 $Y2=4.28
r76 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=13.4 $Y=4.415
+ $X2=13.4 $Y2=4.88
r77 1 23 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=13.375 $Y=4.145
+ $X2=13.375 $Y2=4.28
r78 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=13.375 $Y=4.145
+ $X2=13.375 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2854_265# 1 2 9 11 12 15 17 18 21 28
+ 32
c85 15 0 8.59607e-20 $X=14.84 $Y=2.075
c86 12 0 1.93373e-19 $X=14.46 $Y=1.4
c87 9 0 2.06539e-19 $X=14.37 $Y=2.075
r88 26 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=15.31 $Y=1.42
+ $X2=15.595 $Y2=1.63
r89 25 32 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=15.145 $Y=1.34
+ $X2=14.84 $Y2=1.34
r90 24 26 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=15.145 $Y=1.42
+ $X2=15.31 $Y2=1.42
r91 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.145
+ $Y=1.34 $X2=15.145 $Y2=1.34
r92 21 28 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=15.595 $Y=2.31
+ $X2=15.595 $Y2=1.635
r93 18 26 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=15.31 $Y=1.205
+ $X2=15.31 $Y2=1.42
r94 17 31 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=15.31 $Y=0.755
+ $X2=15.68 $Y2=0.457
r95 17 18 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=15.31 $Y=0.755
+ $X2=15.31 $Y2=1.205
r96 13 32 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=14.84 $Y=1.475
+ $X2=14.84 $Y2=1.34
r97 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=14.84 $Y=1.475
+ $X2=14.84 $Y2=2.075
r98 11 32 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=14.75 $Y=1.4
+ $X2=14.84 $Y2=1.34
r99 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=14.75 $Y=1.4
+ $X2=14.46 $Y2=1.4
r100 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=14.37 $Y=1.475
+ $X2=14.46 $Y2=1.4
r101 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=14.37 $Y=1.475
+ $X2=14.37 $Y2=2.075
r102 2 28 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=15.47
+ $Y=1.485 $X2=15.595 $Y2=1.63
r103 2 21 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=15.47
+ $Y=1.485 $X2=15.595 $Y2=2.31
r104 1 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=15.555
+ $Y=0.235 $X2=15.68 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2854_793# 1 2 9 11 12 15 18 19 21 32
c80 15 0 8.62217e-20 $X=14.84 $Y=3.365
c81 12 0 1.93373e-19 $X=14.46 $Y=4.04
c82 9 0 1.91829e-19 $X=14.37 $Y=3.365
r83 25 32 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=15.145 $Y=4.1
+ $X2=14.84 $Y2=4.1
r84 24 26 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=15.145 $Y=4.02
+ $X2=15.31 $Y2=4.02
r85 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.145
+ $Y=4.1 $X2=15.145 $Y2=4.1
r86 19 26 13.4767 $w=2.58e-07 $l=3.77492e-07 $layer=LI1_cond $X=15.595 $Y=3.805
+ $X2=15.31 $Y2=4.02
r87 19 21 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=15.595 $Y=3.805
+ $X2=15.595 $Y2=3.13
r88 18 31 16.1792 $w=2.79e-07 $l=4.9678e-07 $layer=LI1_cond $X=15.31 $Y=4.685
+ $X2=15.68 $Y2=4.982
r89 17 26 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=15.31 $Y=4.235
+ $X2=15.31 $Y2=4.02
r90 17 18 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=15.31 $Y=4.235
+ $X2=15.31 $Y2=4.685
r91 13 32 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=14.84 $Y=3.965
+ $X2=14.84 $Y2=4.1
r92 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=14.84 $Y=3.965
+ $X2=14.84 $Y2=3.365
r93 11 32 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=14.75 $Y=4.04
+ $X2=14.84 $Y2=4.1
r94 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=14.75 $Y=4.04
+ $X2=14.46 $Y2=4.04
r95 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=14.37 $Y=3.965
+ $X2=14.46 $Y2=4.04
r96 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=14.37 $Y=3.965 $X2=14.37
+ $Y2=3.365
r97 2 19 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=15.47
+ $Y=2.955 $X2=15.595 $Y2=3.81
r98 2 21 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=15.47
+ $Y=2.955 $X2=15.595 $Y2=3.13
r99 1 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=15.555
+ $Y=4.685 $X2=15.68 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[4] 1 3 4 5 6 8 9 12 13 14 15 17 18
+ 20 21 22
r66 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=15.835 $Y=0.92
+ $X2=15.835 $Y2=1.16
r67 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.835
+ $Y=1.16 $X2=15.835 $Y2=1.16
r68 18 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=15.89 $Y=0.845
+ $X2=15.835 $Y2=0.92
r69 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=15.89 $Y=0.845
+ $X2=15.89 $Y2=0.495
r70 15 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=15.83 $Y=1.41
+ $X2=15.835 $Y2=1.16
r71 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.83 $Y=1.41
+ $X2=15.83 $Y2=1.985
r72 13 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=15.7 $Y=0.92
+ $X2=15.835 $Y2=0.92
r73 13 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=15.7 $Y=0.92
+ $X2=15.32 $Y2=0.92
r74 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.245 $Y=0.845
+ $X2=15.32 $Y2=0.92
r75 11 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=15.245 $Y=0.255
+ $X2=15.245 $Y2=0.845
r76 10 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.835 $Y=0.18
+ $X2=14.76 $Y2=0.18
r77 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.17 $Y=0.18
+ $X2=15.245 $Y2=0.255
r78 9 10 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=15.17 $Y=0.18
+ $X2=14.835 $Y2=0.18
r79 6 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.76 $Y=0.255
+ $X2=14.76 $Y2=0.18
r80 6 8 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=14.76 $Y=0.255
+ $X2=14.76 $Y2=0.605
r81 4 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.685 $Y=0.18
+ $X2=14.76 $Y2=0.18
r82 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=14.685 $Y=0.18
+ $X2=14.415 $Y2=0.18
r83 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=14.34 $Y=0.255
+ $X2=14.415 $Y2=0.18
r84 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=14.34 $Y=0.255
+ $X2=14.34 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[12] 1 3 4 5 6 8 9 12 13 14 15 17 18
+ 20 21 22
r66 25 27 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=15.835 $Y=4.28
+ $X2=15.835 $Y2=4.52
r67 22 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.835
+ $Y=4.28 $X2=15.835 $Y2=4.28
r68 18 27 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=15.89 $Y=4.595
+ $X2=15.835 $Y2=4.52
r69 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=15.89 $Y=4.595
+ $X2=15.89 $Y2=4.945
r70 15 25 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=15.83 $Y=4.03
+ $X2=15.835 $Y2=4.28
r71 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.83 $Y=4.03
+ $X2=15.83 $Y2=3.455
r72 13 27 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=15.7 $Y=4.52
+ $X2=15.835 $Y2=4.52
r73 13 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=15.7 $Y=4.52
+ $X2=15.32 $Y2=4.52
r74 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.245 $Y=4.595
+ $X2=15.32 $Y2=4.52
r75 11 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=15.245 $Y=4.595
+ $X2=15.245 $Y2=5.185
r76 10 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.835 $Y=5.26
+ $X2=14.76 $Y2=5.26
r77 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.17 $Y=5.26
+ $X2=15.245 $Y2=5.185
r78 9 10 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=15.17 $Y=5.26
+ $X2=14.835 $Y2=5.26
r79 6 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.76 $Y=5.185
+ $X2=14.76 $Y2=5.26
r80 6 8 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=14.76 $Y=5.185
+ $X2=14.76 $Y2=4.835
r81 4 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.685 $Y=5.26
+ $X2=14.76 $Y2=5.26
r82 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=14.685 $Y=5.26
+ $X2=14.415 $Y2=5.26
r83 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=14.34 $Y=5.185
+ $X2=14.415 $Y2=5.26
r84 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=14.34 $Y=5.185
+ $X2=14.34 $Y2=4.835
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[5] 1 3 4 6 7 10 11 12 13 15 16 18 20
+ 21 22
r63 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=16.365 $Y=0.92
+ $X2=16.365 $Y2=1.16
r64 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.365
+ $Y=1.16 $X2=16.365 $Y2=1.16
r65 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=17.86 $Y=0.255
+ $X2=17.86 $Y2=0.605
r66 17 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.515 $Y=0.18
+ $X2=17.44 $Y2=0.18
r67 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=17.785 $Y=0.18
+ $X2=17.86 $Y2=0.255
r68 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=17.785 $Y=0.18
+ $X2=17.515 $Y2=0.18
r69 13 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.44 $Y=0.255
+ $X2=17.44 $Y2=0.18
r70 13 15 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=17.44 $Y=0.255
+ $X2=17.44 $Y2=0.605
r71 11 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.365 $Y=0.18
+ $X2=17.44 $Y2=0.18
r72 11 12 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=17.365 $Y=0.18
+ $X2=17.03 $Y2=0.18
r73 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=16.955 $Y=0.255
+ $X2=17.03 $Y2=0.18
r74 9 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=16.955 $Y=0.255
+ $X2=16.955 $Y2=0.845
r75 8 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=16.5 $Y=0.92
+ $X2=16.365 $Y2=0.92
r76 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=16.88 $Y=0.92
+ $X2=16.955 $Y2=0.845
r77 7 8 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=16.88 $Y=0.92 $X2=16.5
+ $Y2=0.92
r78 4 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=16.37 $Y=1.41
+ $X2=16.365 $Y2=1.16
r79 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=16.37 $Y=1.41
+ $X2=16.37 $Y2=1.985
r80 1 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=16.31 $Y=0.845
+ $X2=16.365 $Y2=0.92
r81 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=16.31 $Y=0.845
+ $X2=16.31 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[13] 1 3 4 6 7 10 11 12 13 15 16 18
+ 20 21 22
r66 25 27 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=16.365 $Y=4.28
+ $X2=16.365 $Y2=4.52
r67 22 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.365
+ $Y=4.28 $X2=16.365 $Y2=4.28
r68 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=17.86 $Y=5.185
+ $X2=17.86 $Y2=4.835
r69 17 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.515 $Y=5.26
+ $X2=17.44 $Y2=5.26
r70 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=17.785 $Y=5.26
+ $X2=17.86 $Y2=5.185
r71 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=17.785 $Y=5.26
+ $X2=17.515 $Y2=5.26
r72 13 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.44 $Y=5.185
+ $X2=17.44 $Y2=5.26
r73 13 15 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=17.44 $Y=5.185
+ $X2=17.44 $Y2=4.835
r74 11 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.365 $Y=5.26
+ $X2=17.44 $Y2=5.26
r75 11 12 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=17.365 $Y=5.26
+ $X2=17.03 $Y2=5.26
r76 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=16.955 $Y=5.185
+ $X2=17.03 $Y2=5.26
r77 9 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=16.955 $Y=4.595
+ $X2=16.955 $Y2=5.185
r78 8 27 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=16.5 $Y=4.52
+ $X2=16.365 $Y2=4.52
r79 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=16.88 $Y=4.52
+ $X2=16.955 $Y2=4.595
r80 7 8 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=16.88 $Y=4.52 $X2=16.5
+ $Y2=4.52
r81 4 25 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=16.37 $Y=4.03
+ $X2=16.365 $Y2=4.28
r82 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=16.37 $Y=4.03
+ $X2=16.37 $Y2=3.455
r83 1 27 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=16.31 $Y=4.595
+ $X2=16.365 $Y2=4.52
r84 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=16.31 $Y=4.595
+ $X2=16.31 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3277_47# 1 2 9 11 12 15 19 22 24 28
c81 15 0 2.06539e-19 $X=17.83 $Y=2.075
c82 11 0 1.93373e-19 $X=17.74 $Y=1.4
c83 9 0 8.59607e-20 $X=17.36 $Y=2.075
r84 31 33 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=17.055 $Y=1.34
+ $X2=17.36 $Y2=1.34
r85 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.055
+ $Y=1.34 $X2=17.055 $Y2=1.34
r86 28 30 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=16.89 $Y=1.42
+ $X2=17.055 $Y2=1.42
r87 27 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=16.605 $Y=1.63
+ $X2=16.89 $Y2=1.42
r88 22 28 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=16.89 $Y=1.205
+ $X2=16.89 $Y2=1.42
r89 21 24 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=16.89 $Y=0.755
+ $X2=16.52 $Y2=0.457
r90 21 22 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=16.89 $Y=0.755
+ $X2=16.89 $Y2=1.205
r91 19 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=16.605 $Y=2.31
+ $X2=16.605 $Y2=1.635
r92 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=17.83 $Y=1.475
+ $X2=17.83 $Y2=2.075
r93 12 33 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=17.45 $Y=1.4
+ $X2=17.36 $Y2=1.34
r94 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=17.74 $Y=1.4
+ $X2=17.83 $Y2=1.475
r95 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=17.74 $Y=1.4
+ $X2=17.45 $Y2=1.4
r96 7 33 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=17.36 $Y=1.475
+ $X2=17.36 $Y2=1.34
r97 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=17.36 $Y=1.475 $X2=17.36
+ $Y2=2.075
r98 2 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=16.46
+ $Y=1.485 $X2=16.605 $Y2=1.63
r99 2 19 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=16.46
+ $Y=1.485 $X2=16.605 $Y2=2.31
r100 1 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=16.385
+ $Y=0.235 $X2=16.52 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3277_937# 1 2 9 11 12 15 19 22 24 28
c81 15 0 1.91829e-19 $X=17.83 $Y=3.365
c82 11 0 1.93373e-19 $X=17.74 $Y=4.04
c83 9 0 8.62217e-20 $X=17.36 $Y=3.365
r84 31 33 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=17.055 $Y=4.1
+ $X2=17.36 $Y2=4.1
r85 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.055
+ $Y=4.1 $X2=17.055 $Y2=4.1
r86 28 30 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=16.89 $Y=4.02
+ $X2=17.055 $Y2=4.02
r87 22 24 16.1792 $w=2.79e-07 $l=4.9678e-07 $layer=LI1_cond $X=16.89 $Y=4.685
+ $X2=16.52 $Y2=4.982
r88 21 28 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=16.89 $Y=4.235
+ $X2=16.89 $Y2=4.02
r89 21 22 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=16.89 $Y=4.235
+ $X2=16.89 $Y2=4.685
r90 17 28 13.4767 $w=2.58e-07 $l=3.77492e-07 $layer=LI1_cond $X=16.605 $Y=3.805
+ $X2=16.89 $Y2=4.02
r91 17 19 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=16.605 $Y=3.805
+ $X2=16.605 $Y2=3.13
r92 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=17.83 $Y=3.965
+ $X2=17.83 $Y2=3.365
r93 12 33 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=17.45 $Y=4.04
+ $X2=17.36 $Y2=4.1
r94 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=17.74 $Y=4.04
+ $X2=17.83 $Y2=3.965
r95 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=17.74 $Y=4.04
+ $X2=17.45 $Y2=4.04
r96 7 33 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=17.36 $Y=3.965
+ $X2=17.36 $Y2=4.1
r97 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=17.36 $Y=3.965 $X2=17.36
+ $Y2=3.365
r98 2 17 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=16.46
+ $Y=2.955 $X2=16.605 $Y2=3.81
r99 2 19 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=16.46
+ $Y=2.955 $X2=16.605 $Y2=3.13
r100 1 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=16.385
+ $Y=4.685 $X2=16.52 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[5] 3 7 11 15 17 28
c57 17 0 1.17966e-19 $X=19.09 $Y=1.19
c58 15 0 1.17966e-19 $X=18.825 $Y=1.985
c59 3 0 5.84221e-22 $X=18.355 $Y=1.985
r60 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=18.91
+ $Y=1.16 $X2=18.91 $Y2=1.16
r61 26 28 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=18.825 $Y=1.16
+ $X2=18.91 $Y2=1.16
r62 25 26 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=18.8 $Y=1.16
+ $X2=18.825 $Y2=1.16
r63 24 29 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=18.57 $Y=1.19
+ $X2=18.91 $Y2=1.19
r64 23 25 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=18.57 $Y=1.16 $X2=18.8
+ $Y2=1.16
r65 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=18.57
+ $Y=1.16 $X2=18.57 $Y2=1.16
r66 21 23 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=18.38 $Y=1.16
+ $X2=18.57 $Y2=1.16
r67 19 21 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=18.355 $Y=1.16
+ $X2=18.38 $Y2=1.16
r68 17 29 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=19.09 $Y=1.19
+ $X2=18.91 $Y2=1.19
r69 13 26 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=18.825 $Y=1.295
+ $X2=18.825 $Y2=1.16
r70 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=18.825 $Y=1.295
+ $X2=18.825 $Y2=1.985
r71 9 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=18.8 $Y=1.025
+ $X2=18.8 $Y2=1.16
r72 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=18.8 $Y=1.025
+ $X2=18.8 $Y2=0.56
r73 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=18.38 $Y=1.025
+ $X2=18.38 $Y2=1.16
r74 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=18.38 $Y=1.025
+ $X2=18.38 $Y2=0.56
r75 1 19 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=18.355 $Y=1.295
+ $X2=18.355 $Y2=1.16
r76 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=18.355 $Y=1.295
+ $X2=18.355 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[13] 3 7 11 15 17 28
c57 17 0 1.17966e-19 $X=19.09 $Y=4.25
c58 15 0 1.17966e-19 $X=18.825 $Y=3.455
c59 3 0 5.84221e-22 $X=18.355 $Y=3.455
r60 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=18.91
+ $Y=4.28 $X2=18.91 $Y2=4.28
r61 26 28 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=18.825 $Y=4.28
+ $X2=18.91 $Y2=4.28
r62 25 26 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=18.8 $Y=4.28
+ $X2=18.825 $Y2=4.28
r63 24 29 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=18.57 $Y=4.25
+ $X2=18.91 $Y2=4.25
r64 23 25 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=18.57 $Y=4.28 $X2=18.8
+ $Y2=4.28
r65 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=18.57
+ $Y=4.28 $X2=18.57 $Y2=4.28
r66 21 23 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=18.38 $Y=4.28
+ $X2=18.57 $Y2=4.28
r67 19 21 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=18.355 $Y=4.28
+ $X2=18.38 $Y2=4.28
r68 17 29 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=19.09 $Y=4.25
+ $X2=18.91 $Y2=4.25
r69 13 26 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=18.825 $Y=4.145
+ $X2=18.825 $Y2=4.28
r70 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=18.825 $Y=4.145
+ $X2=18.825 $Y2=3.455
r71 9 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=18.8 $Y=4.415
+ $X2=18.8 $Y2=4.28
r72 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=18.8 $Y=4.415
+ $X2=18.8 $Y2=4.88
r73 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=18.38 $Y=4.415
+ $X2=18.38 $Y2=4.28
r74 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=18.38 $Y=4.415
+ $X2=18.38 $Y2=4.88
r75 1 19 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=18.355 $Y=4.145
+ $X2=18.355 $Y2=4.28
r76 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=18.355 $Y=4.145
+ $X2=18.355 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[6] 3 7 11 15 17 27 29
c58 27 0 1.17966e-19 $X=20.07 $Y=1.16
c59 15 0 5.84221e-22 $X=20.285 $Y=1.985
c60 3 0 1.17966e-19 $X=19.815 $Y=1.985
r61 28 29 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=20.26 $Y=1.16
+ $X2=20.285 $Y2=1.16
r62 26 28 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=20.07 $Y=1.16
+ $X2=20.26 $Y2=1.16
r63 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=20.07
+ $Y=1.16 $X2=20.07 $Y2=1.16
r64 24 26 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=19.84 $Y=1.16 $X2=20.07
+ $Y2=1.16
r65 23 24 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=19.815 $Y=1.16
+ $X2=19.84 $Y2=1.16
r66 21 27 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=19.73 $Y=1.19
+ $X2=20.07 $Y2=1.19
r67 20 23 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=19.73 $Y=1.16
+ $X2=19.815 $Y2=1.16
r68 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=19.73
+ $Y=1.16 $X2=19.73 $Y2=1.16
r69 17 21 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=19.55 $Y=1.19
+ $X2=19.73 $Y2=1.19
r70 13 29 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=20.285 $Y=1.295
+ $X2=20.285 $Y2=1.16
r71 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=20.285 $Y=1.295
+ $X2=20.285 $Y2=1.985
r72 9 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=20.26 $Y=1.025
+ $X2=20.26 $Y2=1.16
r73 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=20.26 $Y=1.025
+ $X2=20.26 $Y2=0.56
r74 5 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=19.84 $Y=1.025
+ $X2=19.84 $Y2=1.16
r75 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=19.84 $Y=1.025
+ $X2=19.84 $Y2=0.56
r76 1 23 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=19.815 $Y=1.295
+ $X2=19.815 $Y2=1.16
r77 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=19.815 $Y=1.295
+ $X2=19.815 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[14] 3 7 11 15 17 27 29
c59 27 0 1.17966e-19 $X=20.07 $Y=4.28
c60 15 0 5.84221e-22 $X=20.285 $Y=3.455
c61 3 0 1.17966e-19 $X=19.815 $Y=3.455
r62 28 29 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=20.26 $Y=4.28
+ $X2=20.285 $Y2=4.28
r63 26 28 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=20.07 $Y=4.28
+ $X2=20.26 $Y2=4.28
r64 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=20.07
+ $Y=4.28 $X2=20.07 $Y2=4.28
r65 24 26 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=19.84 $Y=4.28 $X2=20.07
+ $Y2=4.28
r66 23 24 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=19.815 $Y=4.28
+ $X2=19.84 $Y2=4.28
r67 21 27 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=19.73 $Y=4.25
+ $X2=20.07 $Y2=4.25
r68 20 23 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=19.73 $Y=4.28
+ $X2=19.815 $Y2=4.28
r69 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=19.73
+ $Y=4.28 $X2=19.73 $Y2=4.28
r70 17 21 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=19.55 $Y=4.25
+ $X2=19.73 $Y2=4.25
r71 13 29 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=20.285 $Y=4.145
+ $X2=20.285 $Y2=4.28
r72 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=20.285 $Y=4.145
+ $X2=20.285 $Y2=3.455
r73 9 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=20.26 $Y=4.415
+ $X2=20.26 $Y2=4.28
r74 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=20.26 $Y=4.415
+ $X2=20.26 $Y2=4.88
r75 5 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=19.84 $Y=4.415
+ $X2=19.84 $Y2=4.28
r76 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=19.84 $Y=4.415
+ $X2=19.84 $Y2=4.88
r77 1 23 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=19.815 $Y=4.145
+ $X2=19.815 $Y2=4.28
r78 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=19.815 $Y=4.145
+ $X2=19.815 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4142_265# 1 2 9 11 12 15 17 18 21 28
+ 32
c85 15 0 8.59607e-20 $X=21.28 $Y=2.075
c86 12 0 1.93373e-19 $X=20.9 $Y=1.4
c87 9 0 2.06539e-19 $X=20.81 $Y=2.075
r88 26 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=21.75 $Y=1.42
+ $X2=22.035 $Y2=1.63
r89 25 32 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=21.585 $Y=1.34
+ $X2=21.28 $Y2=1.34
r90 24 26 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=21.585 $Y=1.42
+ $X2=21.75 $Y2=1.42
r91 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=21.585
+ $Y=1.34 $X2=21.585 $Y2=1.34
r92 21 28 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=22.035 $Y=2.31
+ $X2=22.035 $Y2=1.635
r93 18 26 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=21.75 $Y=1.205
+ $X2=21.75 $Y2=1.42
r94 17 31 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=21.75 $Y=0.755
+ $X2=22.12 $Y2=0.457
r95 17 18 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=21.75 $Y=0.755
+ $X2=21.75 $Y2=1.205
r96 13 32 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=21.28 $Y=1.475
+ $X2=21.28 $Y2=1.34
r97 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=21.28 $Y=1.475
+ $X2=21.28 $Y2=2.075
r98 11 32 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=21.19 $Y=1.4
+ $X2=21.28 $Y2=1.34
r99 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=21.19 $Y=1.4
+ $X2=20.9 $Y2=1.4
r100 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=20.81 $Y=1.475
+ $X2=20.9 $Y2=1.4
r101 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=20.81 $Y=1.475
+ $X2=20.81 $Y2=2.075
r102 2 28 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=21.91
+ $Y=1.485 $X2=22.035 $Y2=1.63
r103 2 21 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=21.91
+ $Y=1.485 $X2=22.035 $Y2=2.31
r104 1 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=21.995
+ $Y=0.235 $X2=22.12 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4142_793# 1 2 9 11 12 15 18 19 21 32
c80 15 0 8.62217e-20 $X=21.28 $Y=3.365
c81 12 0 1.93373e-19 $X=20.9 $Y=4.04
c82 9 0 1.91829e-19 $X=20.81 $Y=3.365
r83 25 32 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=21.585 $Y=4.1
+ $X2=21.28 $Y2=4.1
r84 24 26 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=21.585 $Y=4.02
+ $X2=21.75 $Y2=4.02
r85 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=21.585
+ $Y=4.1 $X2=21.585 $Y2=4.1
r86 19 26 13.4767 $w=2.58e-07 $l=3.77492e-07 $layer=LI1_cond $X=22.035 $Y=3.805
+ $X2=21.75 $Y2=4.02
r87 19 21 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=22.035 $Y=3.805
+ $X2=22.035 $Y2=3.13
r88 18 31 16.1792 $w=2.79e-07 $l=4.9678e-07 $layer=LI1_cond $X=21.75 $Y=4.685
+ $X2=22.12 $Y2=4.982
r89 17 26 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=21.75 $Y=4.235
+ $X2=21.75 $Y2=4.02
r90 17 18 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=21.75 $Y=4.235
+ $X2=21.75 $Y2=4.685
r91 13 32 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=21.28 $Y=3.965
+ $X2=21.28 $Y2=4.1
r92 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=21.28 $Y=3.965
+ $X2=21.28 $Y2=3.365
r93 11 32 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=21.19 $Y=4.04
+ $X2=21.28 $Y2=4.1
r94 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=21.19 $Y=4.04
+ $X2=20.9 $Y2=4.04
r95 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=20.81 $Y=3.965
+ $X2=20.9 $Y2=4.04
r96 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=20.81 $Y=3.965 $X2=20.81
+ $Y2=3.365
r97 2 19 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=21.91
+ $Y=2.955 $X2=22.035 $Y2=3.81
r98 2 21 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=21.91
+ $Y=2.955 $X2=22.035 $Y2=3.13
r99 1 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=21.995
+ $Y=4.685 $X2=22.12 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[6] 1 3 4 5 6 8 9 12 13 14 15 17 18
+ 20 21 22
r66 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=22.275 $Y=0.92
+ $X2=22.275 $Y2=1.16
r67 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=22.275
+ $Y=1.16 $X2=22.275 $Y2=1.16
r68 18 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=22.33 $Y=0.845
+ $X2=22.275 $Y2=0.92
r69 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=22.33 $Y=0.845
+ $X2=22.33 $Y2=0.495
r70 15 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=22.27 $Y=1.41
+ $X2=22.275 $Y2=1.16
r71 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=22.27 $Y=1.41
+ $X2=22.27 $Y2=1.985
r72 13 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=22.14 $Y=0.92
+ $X2=22.275 $Y2=0.92
r73 13 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=22.14 $Y=0.92
+ $X2=21.76 $Y2=0.92
r74 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=21.685 $Y=0.845
+ $X2=21.76 $Y2=0.92
r75 11 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=21.685 $Y=0.255
+ $X2=21.685 $Y2=0.845
r76 10 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.275 $Y=0.18
+ $X2=21.2 $Y2=0.18
r77 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=21.61 $Y=0.18
+ $X2=21.685 $Y2=0.255
r78 9 10 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=21.61 $Y=0.18
+ $X2=21.275 $Y2=0.18
r79 6 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.2 $Y=0.255
+ $X2=21.2 $Y2=0.18
r80 6 8 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=21.2 $Y=0.255 $X2=21.2
+ $Y2=0.605
r81 4 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.125 $Y=0.18
+ $X2=21.2 $Y2=0.18
r82 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=21.125 $Y=0.18
+ $X2=20.855 $Y2=0.18
r83 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=20.78 $Y=0.255
+ $X2=20.855 $Y2=0.18
r84 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=20.78 $Y=0.255
+ $X2=20.78 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[14] 1 3 4 5 6 8 9 12 13 14 15 17 18
+ 20 21 22
r66 25 27 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=22.275 $Y=4.28
+ $X2=22.275 $Y2=4.52
r67 22 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=22.275
+ $Y=4.28 $X2=22.275 $Y2=4.28
r68 18 27 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=22.33 $Y=4.595
+ $X2=22.275 $Y2=4.52
r69 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=22.33 $Y=4.595
+ $X2=22.33 $Y2=4.945
r70 15 25 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=22.27 $Y=4.03
+ $X2=22.275 $Y2=4.28
r71 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=22.27 $Y=4.03
+ $X2=22.27 $Y2=3.455
r72 13 27 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=22.14 $Y=4.52
+ $X2=22.275 $Y2=4.52
r73 13 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=22.14 $Y=4.52
+ $X2=21.76 $Y2=4.52
r74 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=21.685 $Y=4.595
+ $X2=21.76 $Y2=4.52
r75 11 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=21.685 $Y=4.595
+ $X2=21.685 $Y2=5.185
r76 10 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.275 $Y=5.26
+ $X2=21.2 $Y2=5.26
r77 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=21.61 $Y=5.26
+ $X2=21.685 $Y2=5.185
r78 9 10 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=21.61 $Y=5.26
+ $X2=21.275 $Y2=5.26
r79 6 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.2 $Y=5.185
+ $X2=21.2 $Y2=5.26
r80 6 8 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=21.2 $Y=5.185 $X2=21.2
+ $Y2=4.835
r81 4 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.125 $Y=5.26
+ $X2=21.2 $Y2=5.26
r82 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=21.125 $Y=5.26
+ $X2=20.855 $Y2=5.26
r83 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=20.78 $Y=5.185
+ $X2=20.855 $Y2=5.26
r84 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=20.78 $Y=5.185
+ $X2=20.78 $Y2=4.835
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[7] 1 3 4 6 7 10 11 12 13 15 16 18 20
+ 21 22
r63 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=22.805 $Y=0.92
+ $X2=22.805 $Y2=1.16
r64 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=22.805
+ $Y=1.16 $X2=22.805 $Y2=1.16
r65 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=24.3 $Y=0.255
+ $X2=24.3 $Y2=0.605
r66 17 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=23.955 $Y=0.18
+ $X2=23.88 $Y2=0.18
r67 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=24.225 $Y=0.18
+ $X2=24.3 $Y2=0.255
r68 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=24.225 $Y=0.18
+ $X2=23.955 $Y2=0.18
r69 13 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=23.88 $Y=0.255
+ $X2=23.88 $Y2=0.18
r70 13 15 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=23.88 $Y=0.255
+ $X2=23.88 $Y2=0.605
r71 11 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=23.805 $Y=0.18
+ $X2=23.88 $Y2=0.18
r72 11 12 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=23.805 $Y=0.18
+ $X2=23.47 $Y2=0.18
r73 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=23.395 $Y=0.255
+ $X2=23.47 $Y2=0.18
r74 9 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=23.395 $Y=0.255
+ $X2=23.395 $Y2=0.845
r75 8 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=22.94 $Y=0.92
+ $X2=22.805 $Y2=0.92
r76 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=23.32 $Y=0.92
+ $X2=23.395 $Y2=0.845
r77 7 8 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=23.32 $Y=0.92
+ $X2=22.94 $Y2=0.92
r78 4 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=22.81 $Y=1.41
+ $X2=22.805 $Y2=1.16
r79 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=22.81 $Y=1.41
+ $X2=22.81 $Y2=1.985
r80 1 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=22.75 $Y=0.845
+ $X2=22.805 $Y2=0.92
r81 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=22.75 $Y=0.845
+ $X2=22.75 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[15] 1 3 4 6 7 10 11 12 13 15 16 18
+ 20 21 22
r66 25 27 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=22.805 $Y=4.28
+ $X2=22.805 $Y2=4.52
r67 22 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=22.805
+ $Y=4.28 $X2=22.805 $Y2=4.28
r68 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=24.3 $Y=5.185
+ $X2=24.3 $Y2=4.835
r69 17 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=23.955 $Y=5.26
+ $X2=23.88 $Y2=5.26
r70 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=24.225 $Y=5.26
+ $X2=24.3 $Y2=5.185
r71 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=24.225 $Y=5.26
+ $X2=23.955 $Y2=5.26
r72 13 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=23.88 $Y=5.185
+ $X2=23.88 $Y2=5.26
r73 13 15 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=23.88 $Y=5.185
+ $X2=23.88 $Y2=4.835
r74 11 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=23.805 $Y=5.26
+ $X2=23.88 $Y2=5.26
r75 11 12 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=23.805 $Y=5.26
+ $X2=23.47 $Y2=5.26
r76 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=23.395 $Y=5.185
+ $X2=23.47 $Y2=5.26
r77 9 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=23.395 $Y=4.595
+ $X2=23.395 $Y2=5.185
r78 8 27 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=22.94 $Y=4.52
+ $X2=22.805 $Y2=4.52
r79 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=23.32 $Y=4.52
+ $X2=23.395 $Y2=4.595
r80 7 8 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=23.32 $Y=4.52
+ $X2=22.94 $Y2=4.52
r81 4 25 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=22.81 $Y=4.03
+ $X2=22.805 $Y2=4.28
r82 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=22.81 $Y=4.03
+ $X2=22.81 $Y2=3.455
r83 1 27 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=22.75 $Y=4.595
+ $X2=22.805 $Y2=4.52
r84 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=22.75 $Y=4.595
+ $X2=22.75 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4565_47# 1 2 9 11 12 15 19 22 24 28
c80 15 0 2.06539e-19 $X=24.27 $Y=2.075
c81 9 0 8.59607e-20 $X=23.8 $Y=2.075
r82 31 33 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=23.495 $Y=1.34
+ $X2=23.8 $Y2=1.34
r83 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=23.495
+ $Y=1.34 $X2=23.495 $Y2=1.34
r84 28 30 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=23.33 $Y=1.42
+ $X2=23.495 $Y2=1.42
r85 27 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=23.045 $Y=1.63
+ $X2=23.33 $Y2=1.42
r86 22 28 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=23.33 $Y=1.205
+ $X2=23.33 $Y2=1.42
r87 21 24 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=23.33 $Y=0.755
+ $X2=22.96 $Y2=0.457
r88 21 22 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=23.33 $Y=0.755
+ $X2=23.33 $Y2=1.205
r89 19 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=23.045 $Y=2.31
+ $X2=23.045 $Y2=1.635
r90 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=24.27 $Y=1.475
+ $X2=24.27 $Y2=2.075
r91 12 33 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=23.89 $Y=1.4
+ $X2=23.8 $Y2=1.34
r92 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=24.18 $Y=1.4
+ $X2=24.27 $Y2=1.475
r93 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=24.18 $Y=1.4
+ $X2=23.89 $Y2=1.4
r94 7 33 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=23.8 $Y=1.475
+ $X2=23.8 $Y2=1.34
r95 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=23.8 $Y=1.475 $X2=23.8
+ $Y2=2.075
r96 2 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=22.9
+ $Y=1.485 $X2=23.045 $Y2=1.63
r97 2 19 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=22.9
+ $Y=1.485 $X2=23.045 $Y2=2.31
r98 1 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=22.825
+ $Y=0.235 $X2=22.96 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4565_937# 1 2 9 11 12 15 19 22 24 28
c80 15 0 1.91829e-19 $X=24.27 $Y=3.365
c81 9 0 8.62217e-20 $X=23.8 $Y=3.365
r82 31 33 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=23.495 $Y=4.1
+ $X2=23.8 $Y2=4.1
r83 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=23.495
+ $Y=4.1 $X2=23.495 $Y2=4.1
r84 28 30 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=23.33 $Y=4.02
+ $X2=23.495 $Y2=4.02
r85 22 24 16.1792 $w=2.79e-07 $l=4.9678e-07 $layer=LI1_cond $X=23.33 $Y=4.685
+ $X2=22.96 $Y2=4.982
r86 21 28 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=23.33 $Y=4.235
+ $X2=23.33 $Y2=4.02
r87 21 22 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=23.33 $Y=4.235
+ $X2=23.33 $Y2=4.685
r88 17 28 13.4767 $w=2.58e-07 $l=3.77492e-07 $layer=LI1_cond $X=23.045 $Y=3.805
+ $X2=23.33 $Y2=4.02
r89 17 19 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=23.045 $Y=3.805
+ $X2=23.045 $Y2=3.13
r90 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=24.27 $Y=3.965
+ $X2=24.27 $Y2=3.365
r91 12 33 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=23.89 $Y=4.04
+ $X2=23.8 $Y2=4.1
r92 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=24.18 $Y=4.04
+ $X2=24.27 $Y2=3.965
r93 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=24.18 $Y=4.04
+ $X2=23.89 $Y2=4.04
r94 7 33 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=23.8 $Y=3.965
+ $X2=23.8 $Y2=4.1
r95 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=23.8 $Y=3.965 $X2=23.8
+ $Y2=3.365
r96 2 17 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=22.9
+ $Y=2.955 $X2=23.045 $Y2=3.81
r97 2 19 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=22.9
+ $Y=2.955 $X2=23.045 $Y2=3.13
r98 1 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=22.825
+ $Y=4.685 $X2=22.96 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[7] 3 7 11 15 17 28
c50 3 0 5.84221e-22 $X=24.795 $Y=1.985
r51 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=25.35
+ $Y=1.16 $X2=25.35 $Y2=1.16
r52 26 28 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=25.265 $Y=1.16
+ $X2=25.35 $Y2=1.16
r53 25 26 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=25.24 $Y=1.16
+ $X2=25.265 $Y2=1.16
r54 24 29 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=25.01 $Y=1.19
+ $X2=25.35 $Y2=1.19
r55 23 25 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=25.01 $Y=1.16 $X2=25.24
+ $Y2=1.16
r56 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=25.01
+ $Y=1.16 $X2=25.01 $Y2=1.16
r57 21 23 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=24.82 $Y=1.16
+ $X2=25.01 $Y2=1.16
r58 19 21 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=24.795 $Y=1.16
+ $X2=24.82 $Y2=1.16
r59 17 29 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=25.53 $Y=1.19
+ $X2=25.35 $Y2=1.19
r60 13 26 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=25.265 $Y=1.295
+ $X2=25.265 $Y2=1.16
r61 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=25.265 $Y=1.295
+ $X2=25.265 $Y2=1.985
r62 9 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=25.24 $Y=1.025
+ $X2=25.24 $Y2=1.16
r63 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=25.24 $Y=1.025
+ $X2=25.24 $Y2=0.56
r64 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=24.82 $Y=1.025
+ $X2=24.82 $Y2=1.16
r65 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=24.82 $Y=1.025
+ $X2=24.82 $Y2=0.56
r66 1 19 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=24.795 $Y=1.295
+ $X2=24.795 $Y2=1.16
r67 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=24.795 $Y=1.295
+ $X2=24.795 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[15] 3 7 11 15 17 28
c50 3 0 5.84221e-22 $X=24.795 $Y=3.455
r51 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=25.35
+ $Y=4.28 $X2=25.35 $Y2=4.28
r52 26 28 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=25.265 $Y=4.28
+ $X2=25.35 $Y2=4.28
r53 25 26 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=25.24 $Y=4.28
+ $X2=25.265 $Y2=4.28
r54 24 29 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=25.01 $Y=4.25
+ $X2=25.35 $Y2=4.25
r55 23 25 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=25.01 $Y=4.28 $X2=25.24
+ $Y2=4.28
r56 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=25.01
+ $Y=4.28 $X2=25.01 $Y2=4.28
r57 21 23 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=24.82 $Y=4.28
+ $X2=25.01 $Y2=4.28
r58 19 21 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=24.795 $Y=4.28
+ $X2=24.82 $Y2=4.28
r59 17 29 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=25.53 $Y=4.25
+ $X2=25.35 $Y2=4.25
r60 13 26 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=25.265 $Y=4.145
+ $X2=25.265 $Y2=4.28
r61 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=25.265 $Y=4.145
+ $X2=25.265 $Y2=3.455
r62 9 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=25.24 $Y=4.415
+ $X2=25.24 $Y2=4.28
r63 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=25.24 $Y=4.415
+ $X2=25.24 $Y2=4.88
r64 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=24.82 $Y=4.415
+ $X2=24.82 $Y2=4.28
r65 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=24.82 $Y=4.415
+ $X2=24.82 $Y2=4.88
r66 1 19 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=24.795 $Y=4.145
+ $X2=24.795 $Y2=4.28
r67 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=24.795 $Y=4.145
+ $X2=24.795 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_27_297# 1 2 3 10 12 23 24 25 26 29
+ 33 35 36 39 42 46
c78 25 0 2.60796e-19 $X=2.05 $Y=2.225
c79 24 0 1.97849e-19 $X=0.405 $Y=2.225
c80 23 0 1.02092e-19 $X=1.055 $Y=2.225
r81 36 42 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.195 $Y=2.225
+ $X2=2.195 $Y2=1.81
r82 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.195 $Y=2.225
+ $X2=2.195 $Y2=2.225
r83 33 39 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.2 $Y=2.225
+ $X2=1.2 $Y2=1.78
r84 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.225 $X2=1.2
+ $Y2=2.225
r85 29 46 0.642024 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.26 $Y=2.225
+ $X2=0.26 $Y2=2.21
r86 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=2.225
+ $X2=0.26 $Y2=2.225
r87 26 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.225
+ $X2=1.2 $Y2=2.225
r88 25 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.05 $Y=2.225
+ $X2=2.195 $Y2=2.225
r89 25 26 0.872523 $w=1.4e-07 $l=7.05e-07 $layer=MET1_cond $X=2.05 $Y=2.225
+ $X2=1.345 $Y2=2.225
r90 24 28 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.405 $Y=2.225
+ $X2=0.26 $Y2=2.225
r91 23 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.055 $Y=2.225
+ $X2=1.2 $Y2=2.225
r92 23 24 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=1.055 $Y=2.225
+ $X2=0.405 $Y2=2.225
r93 16 39 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.665
+ $X2=1.2 $Y2=1.78
r94 13 15 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.395 $Y=1.58
+ $X2=0.245 $Y2=1.58
r95 12 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.115 $Y=1.58
+ $X2=1.2 $Y2=1.665
r96 12 13 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.115 $Y=1.58
+ $X2=0.395 $Y2=1.58
r97 10 15 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=1.665
+ $X2=0.245 $Y2=1.58
r98 10 46 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=0.245 $Y=1.665
+ $X2=0.245 $Y2=2.21
r99 3 42 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=2.05
+ $Y=1.665 $X2=2.195 $Y2=1.81
r100 2 39 300 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.78
r101 1 29 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r102 1 15 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_27_591# 1 2 3 13 14 15 17 23 25 26
+ 27 28 35 37 43
c76 27 0 2.13961e-19 $X=2.05 $Y=3.215
c77 26 0 1.97849e-19 $X=0.405 $Y=3.215
c78 25 0 1.02092e-19 $X=1.055 $Y=3.215
r79 43 45 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.26 $Y=3.1 $X2=0.26
+ $Y2=3.23
r80 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.195 $Y=3.215
+ $X2=2.195 $Y2=3.215
r81 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.215 $X2=1.2
+ $Y2=3.215
r82 30 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=3.215
+ $X2=0.26 $Y2=3.215
r83 28 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=3.215
+ $X2=1.2 $Y2=3.215
r84 27 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.05 $Y=3.215
+ $X2=2.195 $Y2=3.215
r85 27 28 0.872523 $w=1.4e-07 $l=7.05e-07 $layer=MET1_cond $X=2.05 $Y=3.215
+ $X2=1.345 $Y2=3.215
r86 26 30 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.405 $Y=3.215
+ $X2=0.26 $Y2=3.215
r87 25 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.055 $Y=3.215
+ $X2=1.2 $Y2=3.215
r88 25 26 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=1.055 $Y=3.215
+ $X2=0.405 $Y2=3.215
r89 23 38 5.02353 $w=1.7e-07 $l=7e-08 $layer=LI1_cond $X=2.195 $Y=3.145
+ $X2=2.195 $Y2=3.215
r90 21 35 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.2 $Y=3.775 $X2=1.2
+ $Y2=3.215
r91 19 35 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=1.2 $Y=3.145 $X2=1.2
+ $Y2=3.215
r92 17 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=3.06 $X2=1.2
+ $Y2=3.145
r93 14 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.115 $Y=3.86
+ $X2=1.2 $Y2=3.775
r94 14 15 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.115 $Y=3.86
+ $X2=0.395 $Y2=3.86
r95 13 45 8.0671 $w=2.98e-07 $l=2.1e-07 $layer=LI1_cond $X=0.245 $Y=3.44
+ $X2=0.245 $Y2=3.23
r96 11 15 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=0.245 $Y=3.775
+ $X2=0.395 $Y2=3.86
r97 11 13 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=0.245 $Y=3.775
+ $X2=0.245 $Y2=3.44
r98 3 23 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=2.05
+ $Y=2.955 $X2=2.195 $Y2=3.14
r99 2 17 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=2.955 $X2=1.2 $Y2=3.14
r100 1 43 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.955 $X2=0.26 $Y2=3.1
r101 1 13 300 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.955 $X2=0.26 $Y2=3.44
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 18 19 20 21 22 23 24 76 80 83 89 96 100 104 108 111 117 124 128 132
+ 136 139 145 152 156 160 164 167 173 180 184 186 190 194 195 197 201 205 209
+ 213 214 216 220 224 228 232 233 235 239 243 247 251 252 254 258 261 262 263
+ 264 265 266 267 268 277 284 298 301 306 313 327 330 335 342 356 359 364 371
+ 385 388 395 399 402 405 408 411 414 417 420
c956 395 0 3.95698e-19 $X=25.53 $Y=2.72
c957 388 0 2.52313e-19 $X=24.865 $Y=2.72
c958 385 0 1.70179e-19 $X=23.69 $Y=2.72
c959 371 0 2.52313e-19 $X=20.47 $Y=2.72
c960 364 0 7.91396e-19 $X=19.915 $Y=2.72
c961 359 0 2.52313e-19 $X=18.425 $Y=2.72
c962 356 0 1.70179e-19 $X=17.25 $Y=2.72
c963 342 0 2.52313e-19 $X=14.03 $Y=2.72
c964 335 0 7.91396e-19 $X=13.475 $Y=2.72
c965 330 0 2.52313e-19 $X=11.985 $Y=2.72
c966 327 0 1.70179e-19 $X=10.81 $Y=2.72
c967 313 0 2.52313e-19 $X=7.59 $Y=2.72
c968 306 0 7.91396e-19 $X=7.035 $Y=2.72
c969 301 0 2.52313e-19 $X=5.545 $Y=2.72
c970 298 0 1.70179e-19 $X=4.37 $Y=2.72
c971 284 0 2.52313e-19 $X=1.15 $Y=2.72
c972 277 0 3.95698e-19 $X=0.595 $Y=2.72
c973 251 0 1.70179e-19 $X=22.375 $Y=2.72
c974 232 0 1.70179e-19 $X=15.935 $Y=2.72
c975 213 0 1.70179e-19 $X=9.495 $Y=2.72
c976 194 0 1.70179e-19 $X=3.055 $Y=2.72
c977 24 0 1.01508e-19 $X=24.885 $Y=2.955
c978 23 0 1.01508e-19 $X=24.885 $Y=1.485
c979 20 0 8.08707e-20 $X=19.905 $Y=2.955
c980 19 0 8.08707e-20 $X=19.905 $Y=1.485
c981 18 0 8.08707e-20 $X=18.445 $Y=2.955
c982 17 0 8.08707e-20 $X=18.445 $Y=1.485
c983 14 0 8.08707e-20 $X=13.465 $Y=2.955
c984 13 0 8.08707e-20 $X=13.465 $Y=1.485
c985 12 0 8.08707e-20 $X=12.005 $Y=2.955
c986 11 0 8.08707e-20 $X=12.005 $Y=1.485
c987 8 0 8.08707e-20 $X=7.025 $Y=2.955
c988 7 0 8.08707e-20 $X=7.025 $Y=1.485
c989 6 0 8.08707e-20 $X=5.565 $Y=2.955
c990 5 0 8.08707e-20 $X=5.565 $Y=1.485
c991 2 0 1.01508e-19 $X=0.585 $Y=2.955
c992 1 0 1.01508e-19 $X=0.585 $Y=1.485
r993 420 421 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.07 $Y=2.72
+ $X2=25.07 $Y2=2.72
r994 417 418 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=20.01 $Y=2.72
+ $X2=20.01 $Y2=2.72
r995 414 415 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.63 $Y=2.72
+ $X2=18.63 $Y2=2.72
r996 411 412 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=2.72
+ $X2=13.57 $Y2=2.72
r997 408 409 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r998 405 406 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r999 402 403 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r1000 399 400 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r1001 393 420 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=25.165 $Y=2.72
+ $X2=25.015 $Y2=2.72
r1002 393 395 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=25.165 $Y=2.72
+ $X2=25.53 $Y2=2.72
r1003 391 421 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=24.61 $Y=2.72
+ $X2=25.07 $Y2=2.72
r1004 390 391 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.61 $Y=2.72
+ $X2=24.61 $Y2=2.72
r1005 388 420 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=24.865 $Y=2.72
+ $X2=25.015 $Y2=2.72
r1006 388 390 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=24.865 $Y=2.72
+ $X2=24.61 $Y2=2.72
r1007 386 391 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=23.69 $Y=2.72
+ $X2=24.61 $Y2=2.72
r1008 385 386 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=23.69 $Y=2.72
+ $X2=23.69 $Y2=2.72
r1009 383 386 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=22.77 $Y=2.72
+ $X2=23.69 $Y2=2.72
r1010 382 385 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=22.77 $Y=2.72
+ $X2=23.69 $Y2=2.72
r1011 382 383 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=22.77 $Y=2.72
+ $X2=22.77 $Y2=2.72
r1012 380 383 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=22.31 $Y=2.72
+ $X2=22.77 $Y2=2.72
r1013 379 380 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=22.31 $Y=2.72
+ $X2=22.31 $Y2=2.72
r1014 376 380 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=21.39 $Y=2.72
+ $X2=22.31 $Y2=2.72
r1015 375 379 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=21.39 $Y=2.72
+ $X2=22.31 $Y2=2.72
r1016 375 376 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=21.39 $Y=2.72
+ $X2=21.39 $Y2=2.72
r1017 372 376 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=20.47 $Y=2.72
+ $X2=21.39 $Y2=2.72
r1018 372 418 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=20.47 $Y=2.72
+ $X2=20.01 $Y2=2.72
r1019 371 372 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=20.47 $Y=2.72
+ $X2=20.47 $Y2=2.72
r1020 369 417 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=20.215 $Y=2.72
+ $X2=20.065 $Y2=2.72
r1021 369 371 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=20.215 $Y=2.72
+ $X2=20.47 $Y2=2.72
r1022 365 414 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=18.725 $Y=2.72
+ $X2=18.575 $Y2=2.72
r1023 365 367 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=18.725 $Y=2.72
+ $X2=19.55 $Y2=2.72
r1024 364 417 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=19.915 $Y=2.72
+ $X2=20.065 $Y2=2.72
r1025 364 367 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=19.915 $Y=2.72
+ $X2=19.55 $Y2=2.72
r1026 362 415 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=18.17 $Y=2.72
+ $X2=18.63 $Y2=2.72
r1027 361 362 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.17 $Y=2.72
+ $X2=18.17 $Y2=2.72
r1028 359 414 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=18.425 $Y=2.72
+ $X2=18.575 $Y2=2.72
r1029 359 361 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=18.425 $Y=2.72
+ $X2=18.17 $Y2=2.72
r1030 357 362 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=17.25 $Y=2.72
+ $X2=18.17 $Y2=2.72
r1031 356 357 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=17.25 $Y=2.72
+ $X2=17.25 $Y2=2.72
r1032 354 357 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=16.33 $Y=2.72
+ $X2=17.25 $Y2=2.72
r1033 353 356 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=16.33 $Y=2.72
+ $X2=17.25 $Y2=2.72
r1034 353 354 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.33 $Y=2.72
+ $X2=16.33 $Y2=2.72
r1035 351 354 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.87 $Y=2.72
+ $X2=16.33 $Y2=2.72
r1036 350 351 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.87 $Y=2.72
+ $X2=15.87 $Y2=2.72
r1037 347 351 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=14.95 $Y=2.72
+ $X2=15.87 $Y2=2.72
r1038 346 350 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=14.95 $Y=2.72
+ $X2=15.87 $Y2=2.72
r1039 346 347 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.95 $Y=2.72
+ $X2=14.95 $Y2=2.72
r1040 343 347 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=14.03 $Y=2.72
+ $X2=14.95 $Y2=2.72
r1041 343 412 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.03 $Y=2.72
+ $X2=13.57 $Y2=2.72
r1042 342 343 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=2.72
+ $X2=14.03 $Y2=2.72
r1043 340 411 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=13.775 $Y=2.72
+ $X2=13.625 $Y2=2.72
r1044 340 342 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=13.775 $Y=2.72
+ $X2=14.03 $Y2=2.72
r1045 336 408 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=12.285 $Y=2.72
+ $X2=12.135 $Y2=2.72
r1046 336 338 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=12.285 $Y=2.72
+ $X2=13.11 $Y2=2.72
r1047 335 411 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=13.475 $Y=2.72
+ $X2=13.625 $Y2=2.72
r1048 335 338 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=13.475 $Y=2.72
+ $X2=13.11 $Y2=2.72
r1049 333 409 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=12.19 $Y2=2.72
r1050 332 333 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r1051 330 408 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=11.985 $Y=2.72
+ $X2=12.135 $Y2=2.72
r1052 330 332 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.985 $Y=2.72
+ $X2=11.73 $Y2=2.72
r1053 328 333 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.73 $Y2=2.72
r1054 327 328 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r1055 325 328 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.81 $Y2=2.72
r1056 324 327 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=9.89 $Y=2.72
+ $X2=10.81 $Y2=2.72
r1057 324 325 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r1058 322 325 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=9.89 $Y2=2.72
r1059 321 322 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r1060 318 322 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r1061 317 321 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r1062 317 318 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r1063 314 318 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r1064 314 406 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r1065 313 314 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r1066 311 405 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=7.335 $Y=2.72
+ $X2=7.185 $Y2=2.72
r1067 311 313 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.335 $Y=2.72
+ $X2=7.59 $Y2=2.72
r1068 307 402 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.845 $Y=2.72
+ $X2=5.695 $Y2=2.72
r1069 307 309 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=5.845 $Y=2.72
+ $X2=6.67 $Y2=2.72
r1070 306 405 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=7.035 $Y=2.72
+ $X2=7.185 $Y2=2.72
r1071 306 309 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.035 $Y=2.72
+ $X2=6.67 $Y2=2.72
r1072 304 403 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r1073 303 304 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r1074 301 402 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.545 $Y=2.72
+ $X2=5.695 $Y2=2.72
r1075 301 303 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.545 $Y=2.72
+ $X2=5.29 $Y2=2.72
r1076 299 304 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r1077 298 299 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r1078 296 299 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r1079 295 298 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r1080 295 296 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r1081 293 296 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r1082 292 293 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r1083 289 293 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r1084 288 292 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r1085 288 289 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r1086 285 289 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r1087 285 400 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r1088 284 285 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r1089 282 399 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.745 $Y2=2.72
r1090 282 284 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r1091 277 399 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.745 $Y2=2.72
r1092 277 279 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r1093 268 421 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.53 $Y=2.72
+ $X2=25.07 $Y2=2.72
r1094 268 395 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.53 $Y=2.72
+ $X2=25.53 $Y2=2.72
r1095 267 418 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.55 $Y=2.72
+ $X2=20.01 $Y2=2.72
r1096 267 367 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=19.55 $Y=2.72
+ $X2=19.55 $Y2=2.72
r1097 266 267 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.09 $Y=2.72
+ $X2=19.55 $Y2=2.72
r1098 266 415 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.09 $Y=2.72
+ $X2=18.63 $Y2=2.72
r1099 265 412 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=2.72
+ $X2=13.57 $Y2=2.72
r1100 265 338 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r1101 264 265 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=13.11 $Y2=2.72
r1102 264 409 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=12.19 $Y2=2.72
r1103 263 406 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r1104 263 309 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r1105 262 263 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r1106 262 403 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r1107 261 400 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r1108 261 279 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r1109 258 259 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=25.03 $Y=3.5
+ $X2=25.03 $Y2=3.335
r1110 254 256 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=25.03 $Y=1.94
+ $X2=25.03 $Y2=2.105
r1111 251 379 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=22.375 $Y=2.72
+ $X2=22.31 $Y2=2.72
r1112 251 252 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=22.375 $Y=2.72
+ $X2=22.54 $Y2=2.72
r1113 250 382 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=22.705 $Y=2.72
+ $X2=22.77 $Y2=2.72
r1114 250 252 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=22.705 $Y=2.72
+ $X2=22.54 $Y2=2.72
r1115 247 248 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=20.05 $Y=3.5
+ $X2=20.05 $Y2=3.335
r1116 243 245 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=20.05 $Y=1.94
+ $X2=20.05 $Y2=2.105
r1117 239 240 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=18.59 $Y=3.5
+ $X2=18.59 $Y2=3.335
r1118 235 237 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=18.59 $Y=1.94
+ $X2=18.59 $Y2=2.105
r1119 232 350 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=15.935 $Y=2.72
+ $X2=15.87 $Y2=2.72
r1120 232 233 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.935 $Y=2.72
+ $X2=16.1 $Y2=2.72
r1121 231 353 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=16.265 $Y=2.72
+ $X2=16.33 $Y2=2.72
r1122 231 233 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.265 $Y=2.72
+ $X2=16.1 $Y2=2.72
r1123 228 229 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=13.61 $Y=3.5
+ $X2=13.61 $Y2=3.335
r1124 224 226 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=13.61 $Y=1.94
+ $X2=13.61 $Y2=2.105
r1125 220 221 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.15 $Y=3.5
+ $X2=12.15 $Y2=3.335
r1126 216 218 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.15 $Y=1.94
+ $X2=12.15 $Y2=2.105
r1127 213 321 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=9.495 $Y=2.72
+ $X2=9.43 $Y2=2.72
r1128 213 214 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.495 $Y=2.72
+ $X2=9.66 $Y2=2.72
r1129 212 324 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=9.825 $Y=2.72
+ $X2=9.89 $Y2=2.72
r1130 212 214 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.825 $Y=2.72
+ $X2=9.66 $Y2=2.72
r1131 209 210 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.17 $Y=3.5
+ $X2=7.17 $Y2=3.335
r1132 205 207 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.17 $Y=1.94
+ $X2=7.17 $Y2=2.105
r1133 201 202 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.71 $Y=3.5
+ $X2=5.71 $Y2=3.335
r1134 197 199 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.71 $Y=1.94
+ $X2=5.71 $Y2=2.105
r1135 194 292 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.055 $Y=2.72
+ $X2=2.99 $Y2=2.72
r1136 194 195 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.055 $Y=2.72
+ $X2=3.22 $Y2=2.72
r1137 193 295 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.385 $Y=2.72
+ $X2=3.45 $Y2=2.72
r1138 193 195 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=2.72
+ $X2=3.22 $Y2=2.72
r1139 190 191 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=3.5
+ $X2=0.73 $Y2=3.335
r1140 186 188 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=1.94
+ $X2=0.73 $Y2=2.105
r1141 184 259 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=25.015 $Y=3.1
+ $X2=25.015 $Y2=3.335
r1142 181 420 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=25.015 $Y=2.805
+ $X2=25.015 $Y2=2.72
r1143 181 184 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=25.015 $Y=2.805
+ $X2=25.015 $Y2=3.1
r1144 180 256 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=25.015 $Y=2.34
+ $X2=25.015 $Y2=2.105
r1145 178 420 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=25.015 $Y=2.635
+ $X2=25.015 $Y2=2.72
r1146 178 180 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=25.015 $Y=2.635
+ $X2=25.015 $Y2=2.34
r1147 173 175 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=22.54 $Y=3.13
+ $X2=22.54 $Y2=3.81
r1148 171 252 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=22.54 $Y=2.805
+ $X2=22.54 $Y2=2.72
r1149 171 173 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=22.54 $Y=2.805
+ $X2=22.54 $Y2=3.13
r1150 167 170 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=22.54 $Y=1.63
+ $X2=22.54 $Y2=2.31
r1151 165 252 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=22.54 $Y=2.635
+ $X2=22.54 $Y2=2.72
r1152 165 170 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=22.54 $Y=2.635
+ $X2=22.54 $Y2=2.31
r1153 164 248 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=20.065 $Y=3.1
+ $X2=20.065 $Y2=3.335
r1154 161 417 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=20.065 $Y=2.805
+ $X2=20.065 $Y2=2.72
r1155 161 164 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=20.065 $Y=2.805
+ $X2=20.065 $Y2=3.1
r1156 160 245 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=20.065 $Y=2.34
+ $X2=20.065 $Y2=2.105
r1157 158 417 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=20.065 $Y=2.635
+ $X2=20.065 $Y2=2.72
r1158 158 160 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=20.065 $Y=2.635
+ $X2=20.065 $Y2=2.34
r1159 156 240 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=18.575 $Y=3.1
+ $X2=18.575 $Y2=3.335
r1160 153 414 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.575 $Y=2.805
+ $X2=18.575 $Y2=2.72
r1161 153 156 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=18.575 $Y=2.805
+ $X2=18.575 $Y2=3.1
r1162 152 237 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=18.575 $Y=2.34
+ $X2=18.575 $Y2=2.105
r1163 150 414 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.575 $Y=2.635
+ $X2=18.575 $Y2=2.72
r1164 150 152 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=18.575 $Y=2.635
+ $X2=18.575 $Y2=2.34
r1165 145 147 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=16.1 $Y=3.13
+ $X2=16.1 $Y2=3.81
r1166 143 233 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=16.1 $Y=2.805
+ $X2=16.1 $Y2=2.72
r1167 143 145 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=16.1 $Y=2.805
+ $X2=16.1 $Y2=3.13
r1168 139 142 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=16.1 $Y=1.63
+ $X2=16.1 $Y2=2.31
r1169 137 233 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=16.1 $Y=2.635
+ $X2=16.1 $Y2=2.72
r1170 137 142 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=16.1 $Y=2.635
+ $X2=16.1 $Y2=2.31
r1171 136 229 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=13.625 $Y=3.1
+ $X2=13.625 $Y2=3.335
r1172 133 411 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.625 $Y=2.805
+ $X2=13.625 $Y2=2.72
r1173 133 136 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=13.625 $Y=2.805
+ $X2=13.625 $Y2=3.1
r1174 132 226 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=13.625 $Y=2.34
+ $X2=13.625 $Y2=2.105
r1175 130 411 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.625 $Y=2.635
+ $X2=13.625 $Y2=2.72
r1176 130 132 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=13.625 $Y=2.635
+ $X2=13.625 $Y2=2.34
r1177 128 221 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=12.135 $Y=3.1
+ $X2=12.135 $Y2=3.335
r1178 125 408 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.135 $Y=2.805
+ $X2=12.135 $Y2=2.72
r1179 125 128 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=12.135 $Y=2.805
+ $X2=12.135 $Y2=3.1
r1180 124 218 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=12.135 $Y=2.34
+ $X2=12.135 $Y2=2.105
r1181 122 408 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.135 $Y=2.635
+ $X2=12.135 $Y2=2.72
r1182 122 124 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=12.135 $Y=2.635
+ $X2=12.135 $Y2=2.34
r1183 117 119 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.66 $Y=3.13
+ $X2=9.66 $Y2=3.81
r1184 115 214 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.66 $Y=2.805
+ $X2=9.66 $Y2=2.72
r1185 115 117 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=9.66 $Y=2.805
+ $X2=9.66 $Y2=3.13
r1186 111 114 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.66 $Y=1.63
+ $X2=9.66 $Y2=2.31
r1187 109 214 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.66 $Y=2.635
+ $X2=9.66 $Y2=2.72
r1188 109 114 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=9.66 $Y=2.635
+ $X2=9.66 $Y2=2.31
r1189 108 210 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=7.185 $Y=3.1
+ $X2=7.185 $Y2=3.335
r1190 105 405 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.185 $Y=2.805
+ $X2=7.185 $Y2=2.72
r1191 105 108 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=7.185 $Y=2.805
+ $X2=7.185 $Y2=3.1
r1192 104 207 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=7.185 $Y=2.34
+ $X2=7.185 $Y2=2.105
r1193 102 405 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.185 $Y=2.635
+ $X2=7.185 $Y2=2.72
r1194 102 104 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=7.185 $Y=2.635
+ $X2=7.185 $Y2=2.34
r1195 100 202 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=5.695 $Y=3.1
+ $X2=5.695 $Y2=3.335
r1196 97 402 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.695 $Y=2.805
+ $X2=5.695 $Y2=2.72
r1197 97 100 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=5.695 $Y=2.805
+ $X2=5.695 $Y2=3.1
r1198 96 199 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=5.695 $Y=2.34
+ $X2=5.695 $Y2=2.105
r1199 94 402 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.695 $Y=2.635
+ $X2=5.695 $Y2=2.72
r1200 94 96 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=5.695 $Y=2.635
+ $X2=5.695 $Y2=2.34
r1201 89 91 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.22 $Y=3.13
+ $X2=3.22 $Y2=3.81
r1202 87 195 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=2.805
+ $X2=3.22 $Y2=2.72
r1203 87 89 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.22 $Y=2.805
+ $X2=3.22 $Y2=3.13
r1204 83 86 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.22 $Y=1.63
+ $X2=3.22 $Y2=2.31
r1205 81 195 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=2.635
+ $X2=3.22 $Y2=2.72
r1206 81 86 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.22 $Y=2.635
+ $X2=3.22 $Y2=2.31
r1207 80 191 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=0.745 $Y=3.1
+ $X2=0.745 $Y2=3.335
r1208 77 399 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=2.805
+ $X2=0.745 $Y2=2.72
r1209 77 80 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.745 $Y=2.805
+ $X2=0.745 $Y2=3.1
r1210 76 188 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=0.745 $Y=2.34
+ $X2=0.745 $Y2=2.105
r1211 74 399 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=2.635
+ $X2=0.745 $Y2=2.72
r1212 74 76 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.745 $Y=2.635
+ $X2=0.745 $Y2=2.34
r1213 24 258 600 $w=1.7e-07 $l=6.13229e-07 $layer=licon1_PDIFF $count=1
+ $X=24.885 $Y=2.955 $X2=25.03 $Y2=3.5
r1214 24 184 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1
+ $X=24.885 $Y=2.955 $X2=25.03 $Y2=3.1
r1215 23 254 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1
+ $X=24.885 $Y=1.485 $X2=25.03 $Y2=1.94
r1216 23 180 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1
+ $X=24.885 $Y=1.485 $X2=25.03 $Y2=2.34
r1217 22 175 400 $w=1.7e-07 $l=9.40705e-07 $layer=licon1_PDIFF $count=1 $X=22.36
+ $Y=2.955 $X2=22.54 $Y2=3.81
r1218 22 173 400 $w=1.7e-07 $l=2.52785e-07 $layer=licon1_PDIFF $count=1 $X=22.36
+ $Y=2.955 $X2=22.54 $Y2=3.13
r1219 21 170 400 $w=1.7e-07 $l=9.10563e-07 $layer=licon1_PDIFF $count=1 $X=22.36
+ $Y=1.485 $X2=22.54 $Y2=2.31
r1220 21 167 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=22.36
+ $Y=1.485 $X2=22.54 $Y2=1.63
r1221 20 247 600 $w=1.7e-07 $l=6.13229e-07 $layer=licon1_PDIFF $count=1
+ $X=19.905 $Y=2.955 $X2=20.05 $Y2=3.5
r1222 20 164 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1
+ $X=19.905 $Y=2.955 $X2=20.05 $Y2=3.1
r1223 19 243 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1
+ $X=19.905 $Y=1.485 $X2=20.05 $Y2=1.94
r1224 19 160 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1
+ $X=19.905 $Y=1.485 $X2=20.05 $Y2=2.34
r1225 18 239 600 $w=1.7e-07 $l=6.13229e-07 $layer=licon1_PDIFF $count=1
+ $X=18.445 $Y=2.955 $X2=18.59 $Y2=3.5
r1226 18 156 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1
+ $X=18.445 $Y=2.955 $X2=18.59 $Y2=3.1
r1227 17 235 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1
+ $X=18.445 $Y=1.485 $X2=18.59 $Y2=1.94
r1228 17 152 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1
+ $X=18.445 $Y=1.485 $X2=18.59 $Y2=2.34
r1229 16 147 400 $w=1.7e-07 $l=9.40705e-07 $layer=licon1_PDIFF $count=1 $X=15.92
+ $Y=2.955 $X2=16.1 $Y2=3.81
r1230 16 145 400 $w=1.7e-07 $l=2.52785e-07 $layer=licon1_PDIFF $count=1 $X=15.92
+ $Y=2.955 $X2=16.1 $Y2=3.13
r1231 15 142 400 $w=1.7e-07 $l=9.10563e-07 $layer=licon1_PDIFF $count=1 $X=15.92
+ $Y=1.485 $X2=16.1 $Y2=2.31
r1232 15 139 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=15.92
+ $Y=1.485 $X2=16.1 $Y2=1.63
r1233 14 228 600 $w=1.7e-07 $l=6.13229e-07 $layer=licon1_PDIFF $count=1
+ $X=13.465 $Y=2.955 $X2=13.61 $Y2=3.5
r1234 14 136 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1
+ $X=13.465 $Y=2.955 $X2=13.61 $Y2=3.1
r1235 13 224 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1
+ $X=13.465 $Y=1.485 $X2=13.61 $Y2=1.94
r1236 13 132 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1
+ $X=13.465 $Y=1.485 $X2=13.61 $Y2=2.34
r1237 12 220 600 $w=1.7e-07 $l=6.13229e-07 $layer=licon1_PDIFF $count=1
+ $X=12.005 $Y=2.955 $X2=12.15 $Y2=3.5
r1238 12 128 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1
+ $X=12.005 $Y=2.955 $X2=12.15 $Y2=3.1
r1239 11 216 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1
+ $X=12.005 $Y=1.485 $X2=12.15 $Y2=1.94
r1240 11 124 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1
+ $X=12.005 $Y=1.485 $X2=12.15 $Y2=2.34
r1241 10 119 400 $w=1.7e-07 $l=9.40705e-07 $layer=licon1_PDIFF $count=1 $X=9.48
+ $Y=2.955 $X2=9.66 $Y2=3.81
r1242 10 117 400 $w=1.7e-07 $l=2.52785e-07 $layer=licon1_PDIFF $count=1 $X=9.48
+ $Y=2.955 $X2=9.66 $Y2=3.13
r1243 9 114 400 $w=1.7e-07 $l=9.10563e-07 $layer=licon1_PDIFF $count=1 $X=9.48
+ $Y=1.485 $X2=9.66 $Y2=2.31
r1244 9 111 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=9.48
+ $Y=1.485 $X2=9.66 $Y2=1.63
r1245 8 209 600 $w=1.7e-07 $l=6.13229e-07 $layer=licon1_PDIFF $count=1 $X=7.025
+ $Y=2.955 $X2=7.17 $Y2=3.5
r1246 8 108 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.025
+ $Y=2.955 $X2=7.17 $Y2=3.1
r1247 7 205 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=7.025
+ $Y=1.485 $X2=7.17 $Y2=1.94
r1248 7 104 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.025
+ $Y=1.485 $X2=7.17 $Y2=2.34
r1249 6 201 600 $w=1.7e-07 $l=6.13229e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=2.955 $X2=5.71 $Y2=3.5
r1250 6 100 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=2.955 $X2=5.71 $Y2=3.1
r1251 5 197 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=1.485 $X2=5.71 $Y2=1.94
r1252 5 96 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=1.485 $X2=5.71 $Y2=2.34
r1253 4 91 400 $w=1.7e-07 $l=9.40705e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=2.955 $X2=3.22 $Y2=3.81
r1254 4 89 400 $w=1.7e-07 $l=2.52785e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=2.955 $X2=3.22 $Y2=3.13
r1255 3 86 400 $w=1.7e-07 $l=9.10563e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=1.485 $X2=3.22 $Y2=2.31
r1256 3 83 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=1.485 $X2=3.22 $Y2=1.63
r1257 2 190 600 $w=1.7e-07 $l=6.13229e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.955 $X2=0.73 $Y2=3.5
r1258 2 80 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.955 $X2=0.73 $Y2=3.1
r1259 1 186 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.94
r1260 1 76 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%Z 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
+ 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 102 108 114 120 126 132 138
+ 144 146 149 152 155 158 161 164 167 170 173 176 179 182 185 188 191 193 194
+ 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213
+ 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232
+ 233 234 235 236 254 256 260 261 266 268 272 273 278 280 284 285 290 292 296
+ 297 302 304 308 309 314 316 320 321 326 328 332 333 338 340 344 345
c1216 344 0 5.38286e-20 $X=24.035 $Y=3.42
c1217 338 0 5.38286e-20 $X=24.15 $Y=1.87
c1218 332 0 5.38286e-20 $X=21.045 $Y=3.42
c1219 326 0 5.38286e-20 $X=20.93 $Y=1.87
c1220 320 0 5.38286e-20 $X=17.595 $Y=3.42
c1221 314 0 5.38286e-20 $X=17.71 $Y=1.87
c1222 308 0 5.38286e-20 $X=14.605 $Y=3.42
c1223 302 0 5.38286e-20 $X=14.49 $Y=1.87
c1224 296 0 5.38286e-20 $X=11.155 $Y=3.42
c1225 290 0 5.38286e-20 $X=11.27 $Y=1.87
c1226 284 0 5.38286e-20 $X=8.165 $Y=3.42
c1227 278 0 5.38286e-20 $X=8.05 $Y=1.87
c1228 272 0 5.38286e-20 $X=4.715 $Y=3.42
c1229 266 0 5.38286e-20 $X=4.83 $Y=1.87
c1230 260 0 5.38286e-20 $X=1.725 $Y=3.42
c1231 254 0 5.38286e-20 $X=1.61 $Y=1.87
c1232 215 0 8.64527e-19 $X=20.785 $Y=3.57
c1233 213 0 8.64527e-19 $X=20.785 $Y=1.87
c1234 207 0 8.64527e-19 $X=14.345 $Y=3.57
c1235 205 0 8.64527e-19 $X=14.345 $Y=1.87
c1236 199 0 8.64527e-19 $X=7.905 $Y=3.57
c1237 197 0 8.64527e-19 $X=7.905 $Y=1.87
r1238 344 348 11.465 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=24.08 $Y=3.42
+ $X2=24.08 $Y2=3.685
r1239 344 345 7.17683 $w=4.28e-07 $l=1.05e-07 $layer=LI1_cond $X=24.08 $Y=3.42
+ $X2=24.08 $Y2=3.315
r1240 342 345 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=24.09 $Y=2.125
+ $X2=24.09 $Y2=3.315
r1241 338 342 11.197 $w=4.28e-07 $l=2.55e-07 $layer=LI1_cond $X=24.08 $Y=1.87
+ $X2=24.08 $Y2=2.125
r1242 338 340 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=24.08 $Y=1.87
+ $X2=24.08 $Y2=1.755
r1243 332 336 11.465 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=21 $Y=3.42
+ $X2=21 $Y2=3.685
r1244 332 333 7.17683 $w=4.28e-07 $l=1.05e-07 $layer=LI1_cond $X=21 $Y=3.42
+ $X2=21 $Y2=3.315
r1245 330 333 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=20.99 $Y=2.125
+ $X2=20.99 $Y2=3.315
r1246 326 330 11.197 $w=4.28e-07 $l=2.55e-07 $layer=LI1_cond $X=21 $Y=1.87
+ $X2=21 $Y2=2.125
r1247 326 328 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=21 $Y=1.87
+ $X2=21 $Y2=1.755
r1248 320 324 11.465 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=17.64 $Y=3.42
+ $X2=17.64 $Y2=3.685
r1249 320 321 7.17683 $w=4.28e-07 $l=1.05e-07 $layer=LI1_cond $X=17.64 $Y=3.42
+ $X2=17.64 $Y2=3.315
r1250 318 321 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=17.65 $Y=2.125
+ $X2=17.65 $Y2=3.315
r1251 314 318 11.197 $w=4.28e-07 $l=2.55e-07 $layer=LI1_cond $X=17.64 $Y=1.87
+ $X2=17.64 $Y2=2.125
r1252 314 316 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=17.64 $Y=1.87
+ $X2=17.64 $Y2=1.755
r1253 308 312 11.465 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=14.56 $Y=3.42
+ $X2=14.56 $Y2=3.685
r1254 308 309 7.17683 $w=4.28e-07 $l=1.05e-07 $layer=LI1_cond $X=14.56 $Y=3.42
+ $X2=14.56 $Y2=3.315
r1255 306 309 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=14.55 $Y=2.125
+ $X2=14.55 $Y2=3.315
r1256 302 306 11.197 $w=4.28e-07 $l=2.55e-07 $layer=LI1_cond $X=14.56 $Y=1.87
+ $X2=14.56 $Y2=2.125
r1257 302 304 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=14.56 $Y=1.87
+ $X2=14.56 $Y2=1.755
r1258 296 300 11.465 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=11.2 $Y=3.42
+ $X2=11.2 $Y2=3.685
r1259 296 297 7.17683 $w=4.28e-07 $l=1.05e-07 $layer=LI1_cond $X=11.2 $Y=3.42
+ $X2=11.2 $Y2=3.315
r1260 294 297 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=11.21 $Y=2.125
+ $X2=11.21 $Y2=3.315
r1261 290 294 11.197 $w=4.28e-07 $l=2.55e-07 $layer=LI1_cond $X=11.2 $Y=1.87
+ $X2=11.2 $Y2=2.125
r1262 290 292 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=11.2 $Y=1.87
+ $X2=11.2 $Y2=1.755
r1263 284 288 11.465 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=8.12 $Y=3.42
+ $X2=8.12 $Y2=3.685
r1264 284 285 7.17683 $w=4.28e-07 $l=1.05e-07 $layer=LI1_cond $X=8.12 $Y=3.42
+ $X2=8.12 $Y2=3.315
r1265 282 285 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=8.11 $Y=2.125
+ $X2=8.11 $Y2=3.315
r1266 278 282 11.197 $w=4.28e-07 $l=2.55e-07 $layer=LI1_cond $X=8.12 $Y=1.87
+ $X2=8.12 $Y2=2.125
r1267 278 280 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=8.12 $Y=1.87
+ $X2=8.12 $Y2=1.755
r1268 272 276 11.465 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=4.76 $Y=3.42
+ $X2=4.76 $Y2=3.685
r1269 272 273 7.17683 $w=4.28e-07 $l=1.05e-07 $layer=LI1_cond $X=4.76 $Y=3.42
+ $X2=4.76 $Y2=3.315
r1270 270 273 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=4.77 $Y=2.125
+ $X2=4.77 $Y2=3.315
r1271 266 270 11.197 $w=4.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.76 $Y=1.87
+ $X2=4.76 $Y2=2.125
r1272 266 268 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.76 $Y=1.87
+ $X2=4.76 $Y2=1.755
r1273 260 264 11.465 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.68 $Y=3.42
+ $X2=1.68 $Y2=3.685
r1274 260 261 7.17683 $w=4.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.68 $Y=3.42
+ $X2=1.68 $Y2=3.315
r1275 258 261 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=1.67 $Y=2.125
+ $X2=1.67 $Y2=3.315
r1276 254 258 11.197 $w=4.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=1.87
+ $X2=1.68 $Y2=2.125
r1277 254 256 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.87
+ $X2=1.68 $Y2=1.755
r1278 236 344 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.15 $Y=3.57
+ $X2=24.15 $Y2=3.57
r1279 235 338 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.15 $Y=1.87
+ $X2=24.15 $Y2=1.87
r1280 234 332 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=20.93 $Y=3.57
+ $X2=20.93 $Y2=3.57
r1281 233 326 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=20.93 $Y=1.87
+ $X2=20.93 $Y2=1.87
r1282 232 320 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.71 $Y=3.57
+ $X2=17.71 $Y2=3.57
r1283 231 314 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.71 $Y=1.87
+ $X2=17.71 $Y2=1.87
r1284 230 308 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.49 $Y=3.57
+ $X2=14.49 $Y2=3.57
r1285 229 302 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.49 $Y=1.87
+ $X2=14.49 $Y2=1.87
r1286 228 296 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=3.57
+ $X2=11.27 $Y2=3.57
r1287 227 290 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=1.87
+ $X2=11.27 $Y2=1.87
r1288 226 284 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=3.57
+ $X2=8.05 $Y2=3.57
r1289 225 278 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=1.87
+ $X2=8.05 $Y2=1.87
r1290 224 272 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=3.57
+ $X2=4.83 $Y2=3.57
r1291 223 266 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=1.87
+ $X2=4.83 $Y2=1.87
r1292 222 260 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=3.57
+ $X2=1.61 $Y2=3.57
r1293 221 254 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=1.87
+ $X2=1.61 $Y2=1.87
r1294 220 234 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.075 $Y=3.57
+ $X2=20.93 $Y2=3.57
r1295 219 236 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=24.005 $Y=3.57
+ $X2=24.15 $Y2=3.57
r1296 219 220 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=24.005 $Y=3.57
+ $X2=21.075 $Y2=3.57
r1297 218 233 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.075 $Y=1.87
+ $X2=20.93 $Y2=1.87
r1298 217 235 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=24.005 $Y=1.87
+ $X2=24.15 $Y2=1.87
r1299 217 218 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=24.005 $Y=1.87
+ $X2=21.075 $Y2=1.87
r1300 216 232 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.855 $Y=3.57
+ $X2=17.71 $Y2=3.57
r1301 215 234 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=20.785 $Y=3.57
+ $X2=20.93 $Y2=3.57
r1302 215 216 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=20.785 $Y=3.57
+ $X2=17.855 $Y2=3.57
r1303 214 231 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.855 $Y=1.87
+ $X2=17.71 $Y2=1.87
r1304 213 233 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=20.785 $Y=1.87
+ $X2=20.93 $Y2=1.87
r1305 213 214 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=20.785 $Y=1.87
+ $X2=17.855 $Y2=1.87
r1306 212 230 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.635 $Y=3.57
+ $X2=14.49 $Y2=3.57
r1307 211 232 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.565 $Y=3.57
+ $X2=17.71 $Y2=3.57
r1308 211 212 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=17.565 $Y=3.57
+ $X2=14.635 $Y2=3.57
r1309 210 229 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.635 $Y=1.87
+ $X2=14.49 $Y2=1.87
r1310 209 231 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.565 $Y=1.87
+ $X2=17.71 $Y2=1.87
r1311 209 210 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=17.565 $Y=1.87
+ $X2=14.635 $Y2=1.87
r1312 208 228 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.415 $Y=3.57
+ $X2=11.27 $Y2=3.57
r1313 207 230 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.345 $Y=3.57
+ $X2=14.49 $Y2=3.57
r1314 207 208 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=14.345 $Y=3.57
+ $X2=11.415 $Y2=3.57
r1315 206 227 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.415 $Y=1.87
+ $X2=11.27 $Y2=1.87
r1316 205 229 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.345 $Y=1.87
+ $X2=14.49 $Y2=1.87
r1317 205 206 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=14.345 $Y=1.87
+ $X2=11.415 $Y2=1.87
r1318 204 226 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.195 $Y=3.57
+ $X2=8.05 $Y2=3.57
r1319 203 228 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.125 $Y=3.57
+ $X2=11.27 $Y2=3.57
r1320 203 204 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=11.125 $Y=3.57
+ $X2=8.195 $Y2=3.57
r1321 202 225 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.195 $Y=1.87
+ $X2=8.05 $Y2=1.87
r1322 201 227 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.125 $Y=1.87
+ $X2=11.27 $Y2=1.87
r1323 201 202 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=11.125 $Y=1.87
+ $X2=8.195 $Y2=1.87
r1324 200 224 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.975 $Y=3.57
+ $X2=4.83 $Y2=3.57
r1325 199 226 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.905 $Y=3.57
+ $X2=8.05 $Y2=3.57
r1326 199 200 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=7.905 $Y=3.57
+ $X2=4.975 $Y2=3.57
r1327 198 223 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.975 $Y=1.87
+ $X2=4.83 $Y2=1.87
r1328 197 225 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.905 $Y=1.87
+ $X2=8.05 $Y2=1.87
r1329 197 198 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=7.905 $Y=1.87
+ $X2=4.975 $Y2=1.87
r1330 196 222 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.755 $Y=3.57
+ $X2=1.61 $Y2=3.57
r1331 195 224 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.685 $Y=3.57
+ $X2=4.83 $Y2=3.57
r1332 195 196 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=4.685 $Y=3.57
+ $X2=1.755 $Y2=3.57
r1333 194 221 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.755 $Y=1.87
+ $X2=1.61 $Y2=1.87
r1334 193 223 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.685 $Y=1.87
+ $X2=4.83 $Y2=1.87
r1335 193 194 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=4.685 $Y=1.87
+ $X2=1.755 $Y2=1.87
r1336 144 191 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=24.09 $Y=4.555
+ $X2=24.09 $Y2=4.76
r1337 144 348 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=24.09 $Y=4.555
+ $X2=24.09 $Y2=3.685
r1338 139 188 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=24.09 $Y=0.885
+ $X2=24.09 $Y2=0.68
r1339 139 340 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=24.09 $Y=0.885
+ $X2=24.09 $Y2=1.755
r1340 138 185 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=20.99 $Y=4.555
+ $X2=20.99 $Y2=4.76
r1341 138 336 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=20.99 $Y=4.555
+ $X2=20.99 $Y2=3.685
r1342 133 182 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=20.99 $Y=0.885
+ $X2=20.99 $Y2=0.68
r1343 133 328 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=20.99 $Y=0.885
+ $X2=20.99 $Y2=1.755
r1344 132 179 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=17.65 $Y=4.555
+ $X2=17.65 $Y2=4.76
r1345 132 324 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=17.65 $Y=4.555
+ $X2=17.65 $Y2=3.685
r1346 127 176 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=17.65 $Y=0.885
+ $X2=17.65 $Y2=0.68
r1347 127 316 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=17.65 $Y=0.885
+ $X2=17.65 $Y2=1.755
r1348 126 173 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=14.55 $Y=4.555
+ $X2=14.55 $Y2=4.76
r1349 126 312 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=14.55 $Y=4.555
+ $X2=14.55 $Y2=3.685
r1350 121 170 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=14.55 $Y=0.885
+ $X2=14.55 $Y2=0.68
r1351 121 304 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=14.55 $Y=0.885
+ $X2=14.55 $Y2=1.755
r1352 120 167 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=11.21 $Y=4.555
+ $X2=11.21 $Y2=4.76
r1353 120 300 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=11.21 $Y=4.555
+ $X2=11.21 $Y2=3.685
r1354 115 164 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=11.21 $Y=0.885
+ $X2=11.21 $Y2=0.68
r1355 115 292 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=11.21 $Y=0.885
+ $X2=11.21 $Y2=1.755
r1356 114 161 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=8.11 $Y=4.555
+ $X2=8.11 $Y2=4.76
r1357 114 288 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=8.11 $Y=4.555
+ $X2=8.11 $Y2=3.685
r1358 109 158 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=8.11 $Y=0.885
+ $X2=8.11 $Y2=0.68
r1359 109 280 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=8.11 $Y=0.885
+ $X2=8.11 $Y2=1.755
r1360 108 155 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=4.77 $Y=4.555
+ $X2=4.77 $Y2=4.76
r1361 108 276 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=4.77 $Y=4.555
+ $X2=4.77 $Y2=3.685
r1362 103 152 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=4.77 $Y=0.885
+ $X2=4.77 $Y2=0.68
r1363 103 268 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=4.77 $Y=0.885
+ $X2=4.77 $Y2=1.755
r1364 102 149 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.67 $Y=4.555
+ $X2=1.67 $Y2=4.76
r1365 102 264 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=1.67 $Y=4.555
+ $X2=1.67 $Y2=3.685
r1366 97 146 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.67 $Y=0.885
+ $X2=1.67 $Y2=0.68
r1367 97 256 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=1.67 $Y=0.885
+ $X2=1.67 $Y2=1.755
r1368 32 344 600 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=1 $X=23.89
+ $Y=2.955 $X2=24.035 $Y2=3.42
r1369 31 338 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=23.89
+ $Y=1.665 $X2=24.035 $Y2=2.02
r1370 30 332 600 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=1 $X=20.9
+ $Y=2.955 $X2=21.045 $Y2=3.42
r1371 29 326 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=20.9
+ $Y=1.665 $X2=21.045 $Y2=2.02
r1372 28 320 600 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=1 $X=17.45
+ $Y=2.955 $X2=17.595 $Y2=3.42
r1373 27 314 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=17.45
+ $Y=1.665 $X2=17.595 $Y2=2.02
r1374 26 308 600 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=1 $X=14.46
+ $Y=2.955 $X2=14.605 $Y2=3.42
r1375 25 302 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=14.46
+ $Y=1.665 $X2=14.605 $Y2=2.02
r1376 24 296 600 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=1 $X=11.01
+ $Y=2.955 $X2=11.155 $Y2=3.42
r1377 23 290 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=11.01
+ $Y=1.665 $X2=11.155 $Y2=2.02
r1378 22 284 600 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=1 $X=8.02
+ $Y=2.955 $X2=8.165 $Y2=3.42
r1379 21 278 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=8.02
+ $Y=1.665 $X2=8.165 $Y2=2.02
r1380 20 272 600 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=1 $X=4.57
+ $Y=2.955 $X2=4.715 $Y2=3.42
r1381 19 266 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=4.57
+ $Y=1.665 $X2=4.715 $Y2=2.02
r1382 18 260 600 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=2.955 $X2=1.725 $Y2=3.42
r1383 17 254 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.665 $X2=1.725 $Y2=2.02
r1384 16 191 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1
+ $X=23.955 $Y=4.575 $X2=24.09 $Y2=4.76
r1385 15 188 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=23.955
+ $Y=0.345 $X2=24.09 $Y2=0.68
r1386 14 185 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1
+ $X=20.855 $Y=4.575 $X2=20.99 $Y2=4.76
r1387 13 182 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=20.855
+ $Y=0.345 $X2=20.99 $Y2=0.68
r1388 12 179 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1
+ $X=17.515 $Y=4.575 $X2=17.65 $Y2=4.76
r1389 11 176 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=17.515
+ $Y=0.345 $X2=17.65 $Y2=0.68
r1390 10 173 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1
+ $X=14.415 $Y=4.575 $X2=14.55 $Y2=4.76
r1391 9 170 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=14.415
+ $Y=0.345 $X2=14.55 $Y2=0.68
r1392 8 167 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=11.075
+ $Y=4.575 $X2=11.21 $Y2=4.76
r1393 7 164 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=11.075
+ $Y=0.345 $X2=11.21 $Y2=0.68
r1394 6 161 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=7.975
+ $Y=4.575 $X2=8.11 $Y2=4.76
r1395 5 158 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=7.975
+ $Y=0.345 $X2=8.11 $Y2=0.68
r1396 4 155 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.635
+ $Y=4.575 $X2=4.77 $Y2=4.76
r1397 3 152 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=4.635
+ $Y=0.345 $X2=4.77 $Y2=0.68
r1398 2 149 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=4.575 $X2=1.67 $Y2=4.76
r1399 1 146 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.345 $X2=1.67 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_824_333# 1 2 3 10 11 12 23 24 25 26
+ 29 33 35 36 39 43 46
c96 36 0 1.37732e-19 $X=6.18 $Y=2.225
c97 35 0 1.97849e-19 $X=6.18 $Y=2.225
c98 25 0 8.14549e-20 $X=6.035 $Y=2.225
c99 23 0 2.60796e-19 $X=5.095 $Y=2.225
c100 3 0 1.01158e-19 $X=6.035 $Y=1.485
r101 36 46 0.642024 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.18 $Y=2.225
+ $X2=6.18 $Y2=2.21
r102 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.18 $Y=2.225
+ $X2=6.18 $Y2=2.225
r103 33 43 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=5.24 $Y=2.225
+ $X2=5.24 $Y2=1.78
r104 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.24 $Y=2.225
+ $X2=5.24 $Y2=2.225
r105 29 39 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.245 $Y=2.225
+ $X2=4.245 $Y2=1.81
r106 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.245 $Y=2.225
+ $X2=4.245 $Y2=2.225
r107 26 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.385 $Y=2.225
+ $X2=5.24 $Y2=2.225
r108 25 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.035 $Y=2.225
+ $X2=6.18 $Y2=2.225
r109 25 26 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=6.035 $Y=2.225
+ $X2=5.385 $Y2=2.225
r110 24 28 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.39 $Y=2.225
+ $X2=4.245 $Y2=2.225
r111 23 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.095 $Y=2.225
+ $X2=5.24 $Y2=2.225
r112 23 24 0.872523 $w=1.4e-07 $l=7.05e-07 $layer=MET1_cond $X=5.095 $Y=2.225
+ $X2=4.39 $Y2=2.225
r113 20 43 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=5.24 $Y=1.665
+ $X2=5.24 $Y2=1.78
r114 12 22 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.195 $Y=1.665
+ $X2=6.195 $Y2=1.58
r115 12 46 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=6.195 $Y=1.665
+ $X2=6.195 $Y2=2.21
r116 11 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.325 $Y=1.58
+ $X2=5.24 $Y2=1.665
r117 10 22 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.045 $Y=1.58
+ $X2=6.195 $Y2=1.58
r118 10 11 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.045 $Y=1.58
+ $X2=5.325 $Y2=1.58
r119 3 36 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.035
+ $Y=1.485 $X2=6.18 $Y2=2.34
r120 3 22 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=6.035
+ $Y=1.485 $X2=6.18 $Y2=1.66
r121 2 43 300 $w=1.7e-07 $l=2.50998e-07 $layer=licon1_PDIFF $count=2 $X=5.04
+ $Y=1.665 $X2=5.24 $Y2=1.78
r122 1 39 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=4.12
+ $Y=1.665 $X2=4.245 $Y2=1.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_824_591# 1 2 3 10 11 15 17 20 25 26
+ 27 28 35 37 43
c91 43 0 1.37732e-19 $X=6.18 $Y=3.1
c92 37 0 1.97849e-19 $X=6.18 $Y=3.215
c93 27 0 8.14549e-20 $X=6.035 $Y=3.215
c94 25 0 2.13961e-19 $X=5.095 $Y=3.215
c95 3 0 1.01158e-19 $X=6.035 $Y=2.955
r96 43 45 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=6.18 $Y=3.1 $X2=6.18
+ $Y2=3.23
r97 37 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.18 $Y=3.215
+ $X2=6.18 $Y2=3.215
r98 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.24 $Y=3.215
+ $X2=5.24 $Y2=3.215
r99 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.245 $Y=3.215
+ $X2=4.245 $Y2=3.215
r100 28 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.385 $Y=3.215
+ $X2=5.24 $Y2=3.215
r101 27 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.035 $Y=3.215
+ $X2=6.18 $Y2=3.215
r102 27 28 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=6.035 $Y=3.215
+ $X2=5.385 $Y2=3.215
r103 26 30 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.39 $Y=3.215
+ $X2=4.245 $Y2=3.215
r104 25 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.095 $Y=3.215
+ $X2=5.24 $Y2=3.215
r105 25 26 0.872523 $w=1.4e-07 $l=7.05e-07 $layer=MET1_cond $X=5.095 $Y=3.215
+ $X2=4.39 $Y2=3.215
r106 24 35 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.24 $Y=3.775
+ $X2=5.24 $Y2=3.215
r107 22 35 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=5.24 $Y=3.145
+ $X2=5.24 $Y2=3.215
r108 20 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.24 $Y=3.06
+ $X2=5.24 $Y2=3.145
r109 17 31 5.02353 $w=1.7e-07 $l=7e-08 $layer=LI1_cond $X=4.245 $Y=3.145
+ $X2=4.245 $Y2=3.215
r110 15 45 8.0671 $w=2.98e-07 $l=2.1e-07 $layer=LI1_cond $X=6.195 $Y=3.44
+ $X2=6.195 $Y2=3.23
r111 13 15 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=6.195 $Y=3.775
+ $X2=6.195 $Y2=3.44
r112 11 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.325 $Y=3.86
+ $X2=5.24 $Y2=3.775
r113 10 13 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=6.045 $Y=3.86
+ $X2=6.195 $Y2=3.775
r114 10 11 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.045 $Y=3.86
+ $X2=5.325 $Y2=3.86
r115 3 43 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.035
+ $Y=2.955 $X2=6.18 $Y2=3.1
r116 3 15 300 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=2 $X=6.035
+ $Y=2.955 $X2=6.18 $Y2=3.44
r117 2 20 300 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_PDIFF $count=2 $X=5.04
+ $Y=2.955 $X2=5.24 $Y2=3.14
r118 1 17 300 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_PDIFF $count=2 $X=4.12
+ $Y=2.955 $X2=4.245 $Y2=3.14
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1315_297# 1 2 3 10 12 23 24 25 26 29
+ 33 35 36 39 42 46
c94 29 0 1.37732e-19 $X=6.7 $Y=2.225
c95 25 0 2.60796e-19 $X=8.49 $Y=2.225
c96 24 0 1.97849e-19 $X=6.845 $Y=2.225
c97 23 0 8.14549e-20 $X=7.495 $Y=2.225
c98 1 0 1.01158e-19 $X=6.575 $Y=1.485
r99 36 42 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.635 $Y=2.225
+ $X2=8.635 $Y2=1.81
r100 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.635 $Y=2.225
+ $X2=8.635 $Y2=2.225
r101 33 39 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=7.64 $Y=2.225
+ $X2=7.64 $Y2=1.78
r102 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.64 $Y=2.225
+ $X2=7.64 $Y2=2.225
r103 29 46 0.642024 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.7 $Y=2.225
+ $X2=6.7 $Y2=2.21
r104 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.7 $Y=2.225
+ $X2=6.7 $Y2=2.225
r105 26 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.785 $Y=2.225
+ $X2=7.64 $Y2=2.225
r106 25 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.49 $Y=2.225
+ $X2=8.635 $Y2=2.225
r107 25 26 0.872523 $w=1.4e-07 $l=7.05e-07 $layer=MET1_cond $X=8.49 $Y=2.225
+ $X2=7.785 $Y2=2.225
r108 24 28 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.845 $Y=2.225
+ $X2=6.7 $Y2=2.225
r109 23 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.495 $Y=2.225
+ $X2=7.64 $Y2=2.225
r110 23 24 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=7.495 $Y=2.225
+ $X2=6.845 $Y2=2.225
r111 16 39 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.64 $Y=1.665
+ $X2=7.64 $Y2=1.78
r112 13 15 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.835 $Y=1.58
+ $X2=6.685 $Y2=1.58
r113 12 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.555 $Y=1.58
+ $X2=7.64 $Y2=1.665
r114 12 13 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=7.555 $Y=1.58
+ $X2=6.835 $Y2=1.58
r115 10 15 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.685 $Y=1.665
+ $X2=6.685 $Y2=1.58
r116 10 46 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=6.685 $Y=1.665
+ $X2=6.685 $Y2=2.21
r117 3 42 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=8.49
+ $Y=1.665 $X2=8.635 $Y2=1.81
r118 2 39 300 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=2 $X=7.495
+ $Y=1.485 $X2=7.64 $Y2=1.78
r119 1 29 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=6.575
+ $Y=1.485 $X2=6.7 $Y2=2.34
r120 1 15 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=6.575
+ $Y=1.485 $X2=6.7 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1315_591# 1 2 3 13 14 15 17 23 25 26
+ 27 28 35 37 43
c92 43 0 1.37732e-19 $X=6.7 $Y=3.1
c93 27 0 2.13961e-19 $X=8.49 $Y=3.215
c94 26 0 1.97849e-19 $X=6.845 $Y=3.215
c95 25 0 8.14549e-20 $X=7.495 $Y=3.215
c96 1 0 1.01158e-19 $X=6.575 $Y=2.955
r97 43 45 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=6.7 $Y=3.1 $X2=6.7
+ $Y2=3.23
r98 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.635 $Y=3.215
+ $X2=8.635 $Y2=3.215
r99 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.64 $Y=3.215
+ $X2=7.64 $Y2=3.215
r100 30 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.7 $Y=3.215
+ $X2=6.7 $Y2=3.215
r101 28 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.785 $Y=3.215
+ $X2=7.64 $Y2=3.215
r102 27 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.49 $Y=3.215
+ $X2=8.635 $Y2=3.215
r103 27 28 0.872523 $w=1.4e-07 $l=7.05e-07 $layer=MET1_cond $X=8.49 $Y=3.215
+ $X2=7.785 $Y2=3.215
r104 26 30 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.845 $Y=3.215
+ $X2=6.7 $Y2=3.215
r105 25 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.495 $Y=3.215
+ $X2=7.64 $Y2=3.215
r106 25 26 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=7.495 $Y=3.215
+ $X2=6.845 $Y2=3.215
r107 23 38 5.02353 $w=1.7e-07 $l=7e-08 $layer=LI1_cond $X=8.635 $Y=3.145
+ $X2=8.635 $Y2=3.215
r108 21 35 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.64 $Y=3.775
+ $X2=7.64 $Y2=3.215
r109 19 35 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=7.64 $Y=3.145
+ $X2=7.64 $Y2=3.215
r110 17 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.64 $Y=3.06
+ $X2=7.64 $Y2=3.145
r111 14 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.555 $Y=3.86
+ $X2=7.64 $Y2=3.775
r112 14 15 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=7.555 $Y=3.86
+ $X2=6.835 $Y2=3.86
r113 13 45 8.0671 $w=2.98e-07 $l=2.1e-07 $layer=LI1_cond $X=6.685 $Y=3.44
+ $X2=6.685 $Y2=3.23
r114 11 15 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=6.685 $Y=3.775
+ $X2=6.835 $Y2=3.86
r115 11 13 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=6.685 $Y=3.775
+ $X2=6.685 $Y2=3.44
r116 3 23 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=8.49
+ $Y=2.955 $X2=8.635 $Y2=3.14
r117 2 17 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=7.495
+ $Y=2.955 $X2=7.64 $Y2=3.14
r118 1 43 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=6.575
+ $Y=2.955 $X2=6.7 $Y2=3.1
r119 1 13 300 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_PDIFF $count=2 $X=6.575
+ $Y=2.955 $X2=6.7 $Y2=3.44
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2112_333# 1 2 3 10 11 12 23 24 25 26
+ 29 33 35 36 39 43 46
c96 36 0 1.37732e-19 $X=12.62 $Y=2.225
c97 35 0 1.97849e-19 $X=12.62 $Y=2.225
c98 25 0 8.14549e-20 $X=12.475 $Y=2.225
c99 23 0 2.60796e-19 $X=11.535 $Y=2.225
c100 3 0 1.01158e-19 $X=12.475 $Y=1.485
r101 36 46 0.642024 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=12.62 $Y=2.225
+ $X2=12.62 $Y2=2.21
r102 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.62 $Y=2.225
+ $X2=12.62 $Y2=2.225
r103 33 43 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=11.68 $Y=2.225
+ $X2=11.68 $Y2=1.78
r104 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.68 $Y=2.225
+ $X2=11.68 $Y2=2.225
r105 29 39 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=10.685 $Y=2.225
+ $X2=10.685 $Y2=1.81
r106 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.685 $Y=2.225
+ $X2=10.685 $Y2=2.225
r107 26 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.825 $Y=2.225
+ $X2=11.68 $Y2=2.225
r108 25 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.475 $Y=2.225
+ $X2=12.62 $Y2=2.225
r109 25 26 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=12.475 $Y=2.225
+ $X2=11.825 $Y2=2.225
r110 24 28 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.83 $Y=2.225
+ $X2=10.685 $Y2=2.225
r111 23 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.535 $Y=2.225
+ $X2=11.68 $Y2=2.225
r112 23 24 0.872523 $w=1.4e-07 $l=7.05e-07 $layer=MET1_cond $X=11.535 $Y=2.225
+ $X2=10.83 $Y2=2.225
r113 20 43 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=11.68 $Y=1.665
+ $X2=11.68 $Y2=1.78
r114 12 22 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.635 $Y=1.665
+ $X2=12.635 $Y2=1.58
r115 12 46 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=12.635 $Y=1.665
+ $X2=12.635 $Y2=2.21
r116 11 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.765 $Y=1.58
+ $X2=11.68 $Y2=1.665
r117 10 22 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=12.485 $Y=1.58
+ $X2=12.635 $Y2=1.58
r118 10 11 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=12.485 $Y=1.58
+ $X2=11.765 $Y2=1.58
r119 3 36 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=12.475
+ $Y=1.485 $X2=12.62 $Y2=2.34
r120 3 22 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=12.475
+ $Y=1.485 $X2=12.62 $Y2=1.66
r121 2 43 300 $w=1.7e-07 $l=2.50998e-07 $layer=licon1_PDIFF $count=2 $X=11.48
+ $Y=1.665 $X2=11.68 $Y2=1.78
r122 1 39 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=10.56
+ $Y=1.665 $X2=10.685 $Y2=1.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2112_591# 1 2 3 10 11 15 17 20 25 26
+ 27 28 35 37 43
c91 43 0 1.37732e-19 $X=12.62 $Y=3.1
c92 37 0 1.97849e-19 $X=12.62 $Y=3.215
c93 27 0 8.14549e-20 $X=12.475 $Y=3.215
c94 25 0 2.13961e-19 $X=11.535 $Y=3.215
c95 3 0 1.01158e-19 $X=12.475 $Y=2.955
r96 43 45 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=12.62 $Y=3.1
+ $X2=12.62 $Y2=3.23
r97 37 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.62 $Y=3.215
+ $X2=12.62 $Y2=3.215
r98 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.68 $Y=3.215
+ $X2=11.68 $Y2=3.215
r99 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.685 $Y=3.215
+ $X2=10.685 $Y2=3.215
r100 28 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.825 $Y=3.215
+ $X2=11.68 $Y2=3.215
r101 27 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.475 $Y=3.215
+ $X2=12.62 $Y2=3.215
r102 27 28 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=12.475 $Y=3.215
+ $X2=11.825 $Y2=3.215
r103 26 30 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.83 $Y=3.215
+ $X2=10.685 $Y2=3.215
r104 25 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.535 $Y=3.215
+ $X2=11.68 $Y2=3.215
r105 25 26 0.872523 $w=1.4e-07 $l=7.05e-07 $layer=MET1_cond $X=11.535 $Y=3.215
+ $X2=10.83 $Y2=3.215
r106 24 35 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=11.68 $Y=3.775
+ $X2=11.68 $Y2=3.215
r107 22 35 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=11.68 $Y=3.145
+ $X2=11.68 $Y2=3.215
r108 20 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.68 $Y=3.06
+ $X2=11.68 $Y2=3.145
r109 17 31 5.02353 $w=1.7e-07 $l=7e-08 $layer=LI1_cond $X=10.685 $Y=3.145
+ $X2=10.685 $Y2=3.215
r110 15 45 8.0671 $w=2.98e-07 $l=2.1e-07 $layer=LI1_cond $X=12.635 $Y=3.44
+ $X2=12.635 $Y2=3.23
r111 13 15 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=12.635 $Y=3.775
+ $X2=12.635 $Y2=3.44
r112 11 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.765 $Y=3.86
+ $X2=11.68 $Y2=3.775
r113 10 13 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=12.485 $Y=3.86
+ $X2=12.635 $Y2=3.775
r114 10 11 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=12.485 $Y=3.86
+ $X2=11.765 $Y2=3.86
r115 3 43 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=12.475
+ $Y=2.955 $X2=12.62 $Y2=3.1
r116 3 15 300 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=2 $X=12.475
+ $Y=2.955 $X2=12.62 $Y2=3.44
r117 2 20 300 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_PDIFF $count=2 $X=11.48
+ $Y=2.955 $X2=11.68 $Y2=3.14
r118 1 17 300 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_PDIFF $count=2 $X=10.56
+ $Y=2.955 $X2=10.685 $Y2=3.14
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2603_297# 1 2 3 10 12 23 24 25 26 29
+ 33 35 36 39 42 46
c94 29 0 1.37732e-19 $X=13.14 $Y=2.225
c95 25 0 2.60796e-19 $X=14.93 $Y=2.225
c96 24 0 1.97849e-19 $X=13.285 $Y=2.225
c97 23 0 8.14549e-20 $X=13.935 $Y=2.225
c98 1 0 1.01158e-19 $X=13.015 $Y=1.485
r99 36 42 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=15.075 $Y=2.225
+ $X2=15.075 $Y2=1.81
r100 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.075 $Y=2.225
+ $X2=15.075 $Y2=2.225
r101 33 39 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=14.08 $Y=2.225
+ $X2=14.08 $Y2=1.78
r102 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.08 $Y=2.225
+ $X2=14.08 $Y2=2.225
r103 29 46 0.642024 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=13.14 $Y=2.225
+ $X2=13.14 $Y2=2.21
r104 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.14 $Y=2.225
+ $X2=13.14 $Y2=2.225
r105 26 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.225 $Y=2.225
+ $X2=14.08 $Y2=2.225
r106 25 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.93 $Y=2.225
+ $X2=15.075 $Y2=2.225
r107 25 26 0.872523 $w=1.4e-07 $l=7.05e-07 $layer=MET1_cond $X=14.93 $Y=2.225
+ $X2=14.225 $Y2=2.225
r108 24 28 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.285 $Y=2.225
+ $X2=13.14 $Y2=2.225
r109 23 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.935 $Y=2.225
+ $X2=14.08 $Y2=2.225
r110 23 24 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=13.935 $Y=2.225
+ $X2=13.285 $Y2=2.225
r111 16 39 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=14.08 $Y=1.665
+ $X2=14.08 $Y2=1.78
r112 13 15 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=13.275 $Y=1.58
+ $X2=13.125 $Y2=1.58
r113 12 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.995 $Y=1.58
+ $X2=14.08 $Y2=1.665
r114 12 13 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=13.995 $Y=1.58
+ $X2=13.275 $Y2=1.58
r115 10 15 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.125 $Y=1.665
+ $X2=13.125 $Y2=1.58
r116 10 46 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=13.125 $Y=1.665
+ $X2=13.125 $Y2=2.21
r117 3 42 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=14.93
+ $Y=1.665 $X2=15.075 $Y2=1.81
r118 2 39 300 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=2 $X=13.935
+ $Y=1.485 $X2=14.08 $Y2=1.78
r119 1 29 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=13.015
+ $Y=1.485 $X2=13.14 $Y2=2.34
r120 1 15 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=13.015
+ $Y=1.485 $X2=13.14 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2603_591# 1 2 3 13 14 15 17 23 25 26
+ 27 28 35 37 43
c92 43 0 1.37732e-19 $X=13.14 $Y=3.1
c93 27 0 2.13961e-19 $X=14.93 $Y=3.215
c94 26 0 1.97849e-19 $X=13.285 $Y=3.215
c95 25 0 8.14549e-20 $X=13.935 $Y=3.215
c96 1 0 1.01158e-19 $X=13.015 $Y=2.955
r97 43 45 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=13.14 $Y=3.1
+ $X2=13.14 $Y2=3.23
r98 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.075 $Y=3.215
+ $X2=15.075 $Y2=3.215
r99 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.08 $Y=3.215
+ $X2=14.08 $Y2=3.215
r100 30 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.14 $Y=3.215
+ $X2=13.14 $Y2=3.215
r101 28 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.225 $Y=3.215
+ $X2=14.08 $Y2=3.215
r102 27 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.93 $Y=3.215
+ $X2=15.075 $Y2=3.215
r103 27 28 0.872523 $w=1.4e-07 $l=7.05e-07 $layer=MET1_cond $X=14.93 $Y=3.215
+ $X2=14.225 $Y2=3.215
r104 26 30 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.285 $Y=3.215
+ $X2=13.14 $Y2=3.215
r105 25 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.935 $Y=3.215
+ $X2=14.08 $Y2=3.215
r106 25 26 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=13.935 $Y=3.215
+ $X2=13.285 $Y2=3.215
r107 23 38 5.02353 $w=1.7e-07 $l=7e-08 $layer=LI1_cond $X=15.075 $Y=3.145
+ $X2=15.075 $Y2=3.215
r108 21 35 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=14.08 $Y=3.775
+ $X2=14.08 $Y2=3.215
r109 19 35 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=14.08 $Y=3.145
+ $X2=14.08 $Y2=3.215
r110 17 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.08 $Y=3.06
+ $X2=14.08 $Y2=3.145
r111 14 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.995 $Y=3.86
+ $X2=14.08 $Y2=3.775
r112 14 15 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=13.995 $Y=3.86
+ $X2=13.275 $Y2=3.86
r113 13 45 8.0671 $w=2.98e-07 $l=2.1e-07 $layer=LI1_cond $X=13.125 $Y=3.44
+ $X2=13.125 $Y2=3.23
r114 11 15 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=13.125 $Y=3.775
+ $X2=13.275 $Y2=3.86
r115 11 13 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=13.125 $Y=3.775
+ $X2=13.125 $Y2=3.44
r116 3 23 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=14.93
+ $Y=2.955 $X2=15.075 $Y2=3.14
r117 2 17 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=13.935
+ $Y=2.955 $X2=14.08 $Y2=3.14
r118 1 43 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=13.015
+ $Y=2.955 $X2=13.14 $Y2=3.1
r119 1 13 300 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_PDIFF $count=2 $X=13.015
+ $Y=2.955 $X2=13.14 $Y2=3.44
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3400_333# 1 2 3 10 11 12 23 24 25 26
+ 29 33 35 36 39 43 46
c96 36 0 1.37732e-19 $X=19.06 $Y=2.225
c97 35 0 1.97849e-19 $X=19.06 $Y=2.225
c98 25 0 8.14549e-20 $X=18.915 $Y=2.225
c99 23 0 2.60796e-19 $X=17.975 $Y=2.225
c100 3 0 1.01158e-19 $X=18.915 $Y=1.485
r101 36 46 0.642024 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=19.06 $Y=2.225
+ $X2=19.06 $Y2=2.21
r102 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=19.06 $Y=2.225
+ $X2=19.06 $Y2=2.225
r103 33 43 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=18.12 $Y=2.225
+ $X2=18.12 $Y2=1.78
r104 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.12 $Y=2.225
+ $X2=18.12 $Y2=2.225
r105 29 39 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=17.125 $Y=2.225
+ $X2=17.125 $Y2=1.81
r106 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.125 $Y=2.225
+ $X2=17.125 $Y2=2.225
r107 26 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=18.265 $Y=2.225
+ $X2=18.12 $Y2=2.225
r108 25 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=18.915 $Y=2.225
+ $X2=19.06 $Y2=2.225
r109 25 26 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=18.915 $Y=2.225
+ $X2=18.265 $Y2=2.225
r110 24 28 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.27 $Y=2.225
+ $X2=17.125 $Y2=2.225
r111 23 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.975 $Y=2.225
+ $X2=18.12 $Y2=2.225
r112 23 24 0.872523 $w=1.4e-07 $l=7.05e-07 $layer=MET1_cond $X=17.975 $Y=2.225
+ $X2=17.27 $Y2=2.225
r113 20 43 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=18.12 $Y=1.665
+ $X2=18.12 $Y2=1.78
r114 12 22 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=19.075 $Y=1.665
+ $X2=19.075 $Y2=1.58
r115 12 46 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=19.075 $Y=1.665
+ $X2=19.075 $Y2=2.21
r116 11 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=18.205 $Y=1.58
+ $X2=18.12 $Y2=1.665
r117 10 22 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=18.925 $Y=1.58
+ $X2=19.075 $Y2=1.58
r118 10 11 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=18.925 $Y=1.58
+ $X2=18.205 $Y2=1.58
r119 3 36 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=18.915
+ $Y=1.485 $X2=19.06 $Y2=2.34
r120 3 22 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=18.915
+ $Y=1.485 $X2=19.06 $Y2=1.66
r121 2 43 300 $w=1.7e-07 $l=2.50998e-07 $layer=licon1_PDIFF $count=2 $X=17.92
+ $Y=1.665 $X2=18.12 $Y2=1.78
r122 1 39 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=17
+ $Y=1.665 $X2=17.125 $Y2=1.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3400_591# 1 2 3 10 11 15 17 20 25 26
+ 27 28 35 37 43
c91 43 0 1.37732e-19 $X=19.06 $Y=3.1
c92 37 0 1.97849e-19 $X=19.06 $Y=3.215
c93 27 0 8.14549e-20 $X=18.915 $Y=3.215
c94 25 0 2.13961e-19 $X=17.975 $Y=3.215
c95 3 0 1.01158e-19 $X=18.915 $Y=2.955
r96 43 45 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=19.06 $Y=3.1
+ $X2=19.06 $Y2=3.23
r97 37 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=19.06 $Y=3.215
+ $X2=19.06 $Y2=3.215
r98 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.12 $Y=3.215
+ $X2=18.12 $Y2=3.215
r99 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.125 $Y=3.215
+ $X2=17.125 $Y2=3.215
r100 28 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=18.265 $Y=3.215
+ $X2=18.12 $Y2=3.215
r101 27 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=18.915 $Y=3.215
+ $X2=19.06 $Y2=3.215
r102 27 28 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=18.915 $Y=3.215
+ $X2=18.265 $Y2=3.215
r103 26 30 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.27 $Y=3.215
+ $X2=17.125 $Y2=3.215
r104 25 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.975 $Y=3.215
+ $X2=18.12 $Y2=3.215
r105 25 26 0.872523 $w=1.4e-07 $l=7.05e-07 $layer=MET1_cond $X=17.975 $Y=3.215
+ $X2=17.27 $Y2=3.215
r106 24 35 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=18.12 $Y=3.775
+ $X2=18.12 $Y2=3.215
r107 22 35 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=18.12 $Y=3.145
+ $X2=18.12 $Y2=3.215
r108 20 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=18.12 $Y=3.06
+ $X2=18.12 $Y2=3.145
r109 17 31 5.02353 $w=1.7e-07 $l=7e-08 $layer=LI1_cond $X=17.125 $Y=3.145
+ $X2=17.125 $Y2=3.215
r110 15 45 8.0671 $w=2.98e-07 $l=2.1e-07 $layer=LI1_cond $X=19.075 $Y=3.44
+ $X2=19.075 $Y2=3.23
r111 13 15 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=19.075 $Y=3.775
+ $X2=19.075 $Y2=3.44
r112 11 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=18.205 $Y=3.86
+ $X2=18.12 $Y2=3.775
r113 10 13 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=18.925 $Y=3.86
+ $X2=19.075 $Y2=3.775
r114 10 11 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=18.925 $Y=3.86
+ $X2=18.205 $Y2=3.86
r115 3 43 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=18.915
+ $Y=2.955 $X2=19.06 $Y2=3.1
r116 3 15 300 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=2 $X=18.915
+ $Y=2.955 $X2=19.06 $Y2=3.44
r117 2 20 300 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_PDIFF $count=2 $X=17.92
+ $Y=2.955 $X2=18.12 $Y2=3.14
r118 1 17 300 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_PDIFF $count=2 $X=17
+ $Y=2.955 $X2=17.125 $Y2=3.14
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3891_297# 1 2 3 10 12 23 24 25 26 29
+ 33 35 36 39 42 46
c94 29 0 1.37732e-19 $X=19.58 $Y=2.225
c95 25 0 2.60796e-19 $X=21.37 $Y=2.225
c96 24 0 1.97849e-19 $X=19.725 $Y=2.225
c97 23 0 8.14549e-20 $X=20.375 $Y=2.225
c98 1 0 1.01158e-19 $X=19.455 $Y=1.485
r99 36 42 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=21.515 $Y=2.225
+ $X2=21.515 $Y2=1.81
r100 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=21.515 $Y=2.225
+ $X2=21.515 $Y2=2.225
r101 33 39 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=20.52 $Y=2.225
+ $X2=20.52 $Y2=1.78
r102 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=20.52 $Y=2.225
+ $X2=20.52 $Y2=2.225
r103 29 46 0.642024 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=19.58 $Y=2.225
+ $X2=19.58 $Y2=2.21
r104 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=19.58 $Y=2.225
+ $X2=19.58 $Y2=2.225
r105 26 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=20.665 $Y=2.225
+ $X2=20.52 $Y2=2.225
r106 25 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.37 $Y=2.225
+ $X2=21.515 $Y2=2.225
r107 25 26 0.872523 $w=1.4e-07 $l=7.05e-07 $layer=MET1_cond $X=21.37 $Y=2.225
+ $X2=20.665 $Y2=2.225
r108 24 28 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=19.725 $Y=2.225
+ $X2=19.58 $Y2=2.225
r109 23 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=20.375 $Y=2.225
+ $X2=20.52 $Y2=2.225
r110 23 24 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=20.375 $Y=2.225
+ $X2=19.725 $Y2=2.225
r111 16 39 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=20.52 $Y=1.665
+ $X2=20.52 $Y2=1.78
r112 13 15 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=19.715 $Y=1.58
+ $X2=19.565 $Y2=1.58
r113 12 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=20.435 $Y=1.58
+ $X2=20.52 $Y2=1.665
r114 12 13 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=20.435 $Y=1.58
+ $X2=19.715 $Y2=1.58
r115 10 15 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=19.565 $Y=1.665
+ $X2=19.565 $Y2=1.58
r116 10 46 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=19.565 $Y=1.665
+ $X2=19.565 $Y2=2.21
r117 3 42 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=21.37
+ $Y=1.665 $X2=21.515 $Y2=1.81
r118 2 39 300 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=2 $X=20.375
+ $Y=1.485 $X2=20.52 $Y2=1.78
r119 1 29 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=19.455
+ $Y=1.485 $X2=19.58 $Y2=2.34
r120 1 15 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=19.455
+ $Y=1.485 $X2=19.58 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3891_591# 1 2 3 13 14 15 17 23 25 26
+ 27 28 35 37 43
c92 43 0 1.37732e-19 $X=19.58 $Y=3.1
c93 27 0 2.13961e-19 $X=21.37 $Y=3.215
c94 26 0 1.97849e-19 $X=19.725 $Y=3.215
c95 25 0 8.14549e-20 $X=20.375 $Y=3.215
c96 1 0 1.01158e-19 $X=19.455 $Y=2.955
r97 43 45 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=19.58 $Y=3.1
+ $X2=19.58 $Y2=3.23
r98 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=21.515 $Y=3.215
+ $X2=21.515 $Y2=3.215
r99 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=20.52 $Y=3.215
+ $X2=20.52 $Y2=3.215
r100 30 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=19.58 $Y=3.215
+ $X2=19.58 $Y2=3.215
r101 28 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=20.665 $Y=3.215
+ $X2=20.52 $Y2=3.215
r102 27 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.37 $Y=3.215
+ $X2=21.515 $Y2=3.215
r103 27 28 0.872523 $w=1.4e-07 $l=7.05e-07 $layer=MET1_cond $X=21.37 $Y=3.215
+ $X2=20.665 $Y2=3.215
r104 26 30 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=19.725 $Y=3.215
+ $X2=19.58 $Y2=3.215
r105 25 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=20.375 $Y=3.215
+ $X2=20.52 $Y2=3.215
r106 25 26 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=20.375 $Y=3.215
+ $X2=19.725 $Y2=3.215
r107 23 38 5.02353 $w=1.7e-07 $l=7e-08 $layer=LI1_cond $X=21.515 $Y=3.145
+ $X2=21.515 $Y2=3.215
r108 21 35 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=20.52 $Y=3.775
+ $X2=20.52 $Y2=3.215
r109 19 35 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=20.52 $Y=3.145
+ $X2=20.52 $Y2=3.215
r110 17 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=20.52 $Y=3.06
+ $X2=20.52 $Y2=3.145
r111 14 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=20.435 $Y=3.86
+ $X2=20.52 $Y2=3.775
r112 14 15 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=20.435 $Y=3.86
+ $X2=19.715 $Y2=3.86
r113 13 45 8.0671 $w=2.98e-07 $l=2.1e-07 $layer=LI1_cond $X=19.565 $Y=3.44
+ $X2=19.565 $Y2=3.23
r114 11 15 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=19.565 $Y=3.775
+ $X2=19.715 $Y2=3.86
r115 11 13 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=19.565 $Y=3.775
+ $X2=19.565 $Y2=3.44
r116 3 23 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=21.37
+ $Y=2.955 $X2=21.515 $Y2=3.14
r117 2 17 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=20.375
+ $Y=2.955 $X2=20.52 $Y2=3.14
r118 1 43 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=19.455
+ $Y=2.955 $X2=19.58 $Y2=3.1
r119 1 13 300 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_PDIFF $count=2 $X=19.455
+ $Y=2.955 $X2=19.58 $Y2=3.44
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4688_333# 1 2 3 10 11 12 23 24 25 26
+ 29 33 35 36 39 43 46
c80 35 0 1.97849e-19 $X=25.5 $Y=2.225
c81 25 0 1.02092e-19 $X=25.355 $Y=2.225
c82 23 0 2.60796e-19 $X=24.415 $Y=2.225
r83 36 46 0.642024 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=25.5 $Y=2.225
+ $X2=25.5 $Y2=2.21
r84 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.5 $Y=2.225
+ $X2=25.5 $Y2=2.225
r85 33 43 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=24.56 $Y=2.225
+ $X2=24.56 $Y2=1.78
r86 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.56 $Y=2.225
+ $X2=24.56 $Y2=2.225
r87 29 39 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=23.565 $Y=2.225
+ $X2=23.565 $Y2=1.81
r88 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=23.565 $Y=2.225
+ $X2=23.565 $Y2=2.225
r89 26 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=24.705 $Y=2.225
+ $X2=24.56 $Y2=2.225
r90 25 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=25.355 $Y=2.225
+ $X2=25.5 $Y2=2.225
r91 25 26 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=25.355 $Y=2.225
+ $X2=24.705 $Y2=2.225
r92 24 28 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=23.71 $Y=2.225
+ $X2=23.565 $Y2=2.225
r93 23 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=24.415 $Y=2.225
+ $X2=24.56 $Y2=2.225
r94 23 24 0.872523 $w=1.4e-07 $l=7.05e-07 $layer=MET1_cond $X=24.415 $Y=2.225
+ $X2=23.71 $Y2=2.225
r95 20 43 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=24.56 $Y=1.665
+ $X2=24.56 $Y2=1.78
r96 12 22 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=25.515 $Y=1.665
+ $X2=25.515 $Y2=1.58
r97 12 46 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=25.515 $Y=1.665
+ $X2=25.515 $Y2=2.21
r98 11 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=24.645 $Y=1.58
+ $X2=24.56 $Y2=1.665
r99 10 22 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=25.365 $Y=1.58
+ $X2=25.515 $Y2=1.58
r100 10 11 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=25.365 $Y=1.58
+ $X2=24.645 $Y2=1.58
r101 3 36 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=25.355
+ $Y=1.485 $X2=25.5 $Y2=2.34
r102 3 22 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=25.355
+ $Y=1.485 $X2=25.5 $Y2=1.66
r103 2 43 300 $w=1.7e-07 $l=2.50998e-07 $layer=licon1_PDIFF $count=2 $X=24.36
+ $Y=1.665 $X2=24.56 $Y2=1.78
r104 1 39 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=23.44
+ $Y=1.665 $X2=23.565 $Y2=1.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4688_591# 1 2 3 10 11 15 17 20 25 26
+ 27 28 35 37 43
c75 37 0 1.97849e-19 $X=25.5 $Y=3.215
c76 27 0 1.02092e-19 $X=25.355 $Y=3.215
c77 25 0 2.13961e-19 $X=24.415 $Y=3.215
r78 43 45 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=25.5 $Y=3.1 $X2=25.5
+ $Y2=3.23
r79 37 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.5 $Y=3.215
+ $X2=25.5 $Y2=3.215
r80 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.56 $Y=3.215
+ $X2=24.56 $Y2=3.215
r81 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=23.565 $Y=3.215
+ $X2=23.565 $Y2=3.215
r82 28 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=24.705 $Y=3.215
+ $X2=24.56 $Y2=3.215
r83 27 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=25.355 $Y=3.215
+ $X2=25.5 $Y2=3.215
r84 27 28 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=25.355 $Y=3.215
+ $X2=24.705 $Y2=3.215
r85 26 30 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=23.71 $Y=3.215
+ $X2=23.565 $Y2=3.215
r86 25 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=24.415 $Y=3.215
+ $X2=24.56 $Y2=3.215
r87 25 26 0.872523 $w=1.4e-07 $l=7.05e-07 $layer=MET1_cond $X=24.415 $Y=3.215
+ $X2=23.71 $Y2=3.215
r88 24 35 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=24.56 $Y=3.775
+ $X2=24.56 $Y2=3.215
r89 22 35 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=24.56 $Y=3.145
+ $X2=24.56 $Y2=3.215
r90 20 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=24.56 $Y=3.06
+ $X2=24.56 $Y2=3.145
r91 17 31 5.02353 $w=1.7e-07 $l=7e-08 $layer=LI1_cond $X=23.565 $Y=3.145
+ $X2=23.565 $Y2=3.215
r92 15 45 8.0671 $w=2.98e-07 $l=2.1e-07 $layer=LI1_cond $X=25.515 $Y=3.44
+ $X2=25.515 $Y2=3.23
r93 13 15 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=25.515 $Y=3.775
+ $X2=25.515 $Y2=3.44
r94 11 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=24.645 $Y=3.86
+ $X2=24.56 $Y2=3.775
r95 10 13 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=25.365 $Y=3.86
+ $X2=25.515 $Y2=3.775
r96 10 11 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=25.365 $Y=3.86
+ $X2=24.645 $Y2=3.86
r97 3 43 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=25.355
+ $Y=2.955 $X2=25.5 $Y2=3.1
r98 3 15 300 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=2 $X=25.355
+ $Y=2.955 $X2=25.5 $Y2=3.44
r99 2 20 300 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_PDIFF $count=2 $X=24.36
+ $Y=2.955 $X2=24.56 $Y2=3.14
r100 1 17 300 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_PDIFF $count=2 $X=23.44
+ $Y=2.955 $X2=23.565 $Y2=3.14
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_27_47# 1 2 3 12 14 15 16 18 22
c42 16 0 1.81988e-19 $X=1.182 $Y=0.425
r43 20 22 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.09 $Y=0.425
+ $X2=2.09 $Y2=0.605
r44 19 25 4.85887 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.335 $Y=0.34
+ $X2=1.182 $Y2=0.34
r45 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.005 $Y=0.34
+ $X2=2.09 $Y2=0.425
r46 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=0.34
+ $X2=1.335 $Y2=0.34
r47 16 25 2.69937 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.182 $Y=0.425
+ $X2=1.182 $Y2=0.34
r48 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=1.182 $Y=0.425
+ $X2=1.182 $Y2=0.715
r49 14 17 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=1.03 $Y=0.8
+ $X2=1.182 $Y2=0.715
r50 14 15 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.03 $Y=0.8
+ $X2=0.475 $Y2=0.8
r51 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.31 $Y=0.715
+ $X2=0.475 $Y2=0.8
r52 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.31 $Y=0.715
+ $X2=0.31 $Y2=0.38
r53 3 22 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.345 $X2=2.09 $Y2=0.605
r54 2 25 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.235 $X2=1.175 $Y2=0.42
r55 1 12 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.31 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_27_911# 1 2 3 12 14 16 17 20 23
c43 17 0 1.81988e-19 $X=1.335 $Y=5.1
r44 18 20 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.09 $Y=5.015
+ $X2=2.09 $Y2=4.835
r45 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.005 $Y=5.1
+ $X2=2.09 $Y2=5.015
r46 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=5.1
+ $X2=1.335 $Y2=5.1
r47 15 17 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.182 $Y=5.015
+ $X2=1.335 $Y2=5.1
r48 14 25 2.86504 $w=3.05e-07 $l=1.05e-07 $layer=LI1_cond $X=1.182 $Y=4.725
+ $X2=1.182 $Y2=4.62
r49 14 15 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=1.182 $Y=4.725
+ $X2=1.182 $Y2=5.015
r50 13 23 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.475 $Y=4.64
+ $X2=0.31 $Y2=4.64
r51 12 25 4.6932 $w=1.7e-07 $l=1.61691e-07 $layer=LI1_cond $X=1.03 $Y=4.64
+ $X2=1.182 $Y2=4.62
r52 12 13 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.03 $Y=4.64
+ $X2=0.475 $Y2=4.64
r53 3 20 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=4.575 $X2=2.09 $Y2=4.835
r54 2 25 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=4.555 $X2=1.175 $Y2=4.68
r55 1 23 91 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=4.555 $X2=0.31 $Y2=4.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 18 19 20 21 22 23 24 79 83 87 91 95 99 101 103 107 111 115 119 123
+ 127 129 131 135 139 143 147 151 155 157 159 163 167 171 175 179 183 186 187
+ 189 190 192 193 195 196 198 199 201 202 204 205 207 208 210 211 213 214 215
+ 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 261 268 289 296
+ 317 324 358 362 366 369 372 375 378 381 384 387 390 393 396 399 402 405
r562 405 406 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.01 $Y=5.44
+ $X2=20.01 $Y2=5.44
r563 402 403 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.01 $Y=0
+ $X2=20.01 $Y2=0
r564 399 400 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=18.63 $Y=5.44
+ $X2=18.63 $Y2=5.44
r565 396 397 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=18.63 $Y=0
+ $X2=18.63 $Y2=0
r566 393 394 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.57 $Y=5.44
+ $X2=13.57 $Y2=5.44
r567 390 391 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r568 387 388 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.19 $Y=5.44
+ $X2=12.19 $Y2=5.44
r569 384 385 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r570 381 382 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=5.44
+ $X2=7.13 $Y2=5.44
r571 378 379 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r572 375 376 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=5.44
+ $X2=5.75 $Y2=5.44
r573 372 373 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r574 369 370 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=5.44
+ $X2=0.69 $Y2=5.44
r575 366 367 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r576 355 356 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=24.61 $Y=5.44
+ $X2=24.61 $Y2=5.44
r577 353 356 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=22.77 $Y=5.44
+ $X2=24.61 $Y2=5.44
r578 352 355 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=22.77 $Y=5.44
+ $X2=24.61 $Y2=5.44
r579 352 353 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=22.77 $Y=5.44
+ $X2=22.77 $Y2=5.44
r580 349 350 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=24.61 $Y=0
+ $X2=24.61 $Y2=0
r581 347 350 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=22.77 $Y=0
+ $X2=24.61 $Y2=0
r582 346 349 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=22.77 $Y=0
+ $X2=24.61 $Y2=0
r583 346 347 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=22.77 $Y=0
+ $X2=22.77 $Y2=0
r584 344 353 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=22.31 $Y=5.44
+ $X2=22.77 $Y2=5.44
r585 343 344 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=22.31 $Y=5.44
+ $X2=22.31 $Y2=5.44
r586 341 344 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=20.47 $Y=5.44
+ $X2=22.31 $Y2=5.44
r587 341 406 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=20.47 $Y=5.44
+ $X2=20.01 $Y2=5.44
r588 340 343 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=20.47 $Y=5.44
+ $X2=22.31 $Y2=5.44
r589 340 341 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=20.47 $Y=5.44
+ $X2=20.47 $Y2=5.44
r590 338 405 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=20.18 $Y=5.44
+ $X2=20.072 $Y2=5.44
r591 338 340 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=20.18 $Y=5.44
+ $X2=20.47 $Y2=5.44
r592 337 347 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=22.31 $Y=0
+ $X2=22.77 $Y2=0
r593 336 337 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=22.31 $Y=0
+ $X2=22.31 $Y2=0
r594 334 337 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=20.47 $Y=0
+ $X2=22.31 $Y2=0
r595 334 403 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=20.47 $Y=0
+ $X2=20.01 $Y2=0
r596 333 336 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=20.47 $Y=0
+ $X2=22.31 $Y2=0
r597 333 334 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=20.47 $Y=0
+ $X2=20.47 $Y2=0
r598 331 402 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=20.18 $Y=0
+ $X2=20.072 $Y2=0
r599 331 333 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=20.18 $Y=0
+ $X2=20.47 $Y2=0
r600 330 400 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=18.17 $Y=5.44
+ $X2=18.63 $Y2=5.44
r601 329 330 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=18.17 $Y=5.44
+ $X2=18.17 $Y2=5.44
r602 327 330 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=16.33 $Y=5.44
+ $X2=18.17 $Y2=5.44
r603 326 329 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=16.33 $Y=5.44
+ $X2=18.17 $Y2=5.44
r604 326 327 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=16.33 $Y=5.44
+ $X2=16.33 $Y2=5.44
r605 324 399 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=18.46 $Y=5.44
+ $X2=18.567 $Y2=5.44
r606 324 329 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=18.46 $Y=5.44
+ $X2=18.17 $Y2=5.44
r607 323 397 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=18.17 $Y=0
+ $X2=18.63 $Y2=0
r608 322 323 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=18.17 $Y=0
+ $X2=18.17 $Y2=0
r609 320 323 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=16.33 $Y=0
+ $X2=18.17 $Y2=0
r610 319 322 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=16.33 $Y=0
+ $X2=18.17 $Y2=0
r611 319 320 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=16.33 $Y=0
+ $X2=16.33 $Y2=0
r612 317 396 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=18.46 $Y=0
+ $X2=18.567 $Y2=0
r613 317 322 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=18.46 $Y=0
+ $X2=18.17 $Y2=0
r614 316 327 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.87 $Y=5.44
+ $X2=16.33 $Y2=5.44
r615 315 316 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=15.87 $Y=5.44
+ $X2=15.87 $Y2=5.44
r616 313 316 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=14.03 $Y=5.44
+ $X2=15.87 $Y2=5.44
r617 313 394 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.03 $Y=5.44
+ $X2=13.57 $Y2=5.44
r618 312 315 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=14.03 $Y=5.44
+ $X2=15.87 $Y2=5.44
r619 312 313 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=14.03 $Y=5.44
+ $X2=14.03 $Y2=5.44
r620 310 393 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=13.74 $Y=5.44
+ $X2=13.632 $Y2=5.44
r621 310 312 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=13.74 $Y=5.44
+ $X2=14.03 $Y2=5.44
r622 309 320 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.87 $Y=0
+ $X2=16.33 $Y2=0
r623 308 309 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=15.87 $Y=0
+ $X2=15.87 $Y2=0
r624 306 309 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=14.03 $Y=0
+ $X2=15.87 $Y2=0
r625 306 391 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.03 $Y=0
+ $X2=13.57 $Y2=0
r626 305 308 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=14.03 $Y=0
+ $X2=15.87 $Y2=0
r627 305 306 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=14.03 $Y=0
+ $X2=14.03 $Y2=0
r628 303 390 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=13.74 $Y=0
+ $X2=13.632 $Y2=0
r629 303 305 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=13.74 $Y=0
+ $X2=14.03 $Y2=0
r630 302 388 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=5.44
+ $X2=12.19 $Y2=5.44
r631 301 302 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.73 $Y=5.44
+ $X2=11.73 $Y2=5.44
r632 299 302 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=9.89 $Y=5.44
+ $X2=11.73 $Y2=5.44
r633 298 301 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=9.89 $Y=5.44
+ $X2=11.73 $Y2=5.44
r634 298 299 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.89 $Y=5.44
+ $X2=9.89 $Y2=5.44
r635 296 387 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=12.02 $Y=5.44
+ $X2=12.127 $Y2=5.44
r636 296 301 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=12.02 $Y=5.44
+ $X2=11.73 $Y2=5.44
r637 295 385 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.19 $Y2=0
r638 294 295 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r639 292 295 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=11.73 $Y2=0
r640 291 294 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=9.89 $Y=0
+ $X2=11.73 $Y2=0
r641 291 292 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r642 289 384 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=12.02 $Y=0
+ $X2=12.127 $Y2=0
r643 289 294 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=12.02 $Y=0
+ $X2=11.73 $Y2=0
r644 288 299 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=5.44
+ $X2=9.89 $Y2=5.44
r645 287 288 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.43 $Y=5.44
+ $X2=9.43 $Y2=5.44
r646 285 288 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=7.59 $Y=5.44
+ $X2=9.43 $Y2=5.44
r647 285 382 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=5.44
+ $X2=7.13 $Y2=5.44
r648 284 287 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=7.59 $Y=5.44
+ $X2=9.43 $Y2=5.44
r649 284 285 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.59 $Y=5.44
+ $X2=7.59 $Y2=5.44
r650 282 381 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=7.3 $Y=5.44
+ $X2=7.192 $Y2=5.44
r651 282 284 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.3 $Y=5.44
+ $X2=7.59 $Y2=5.44
r652 281 292 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=9.89 $Y2=0
r653 280 281 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r654 278 281 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=9.43 $Y2=0
r655 278 379 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=7.13 $Y2=0
r656 277 280 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=7.59 $Y=0
+ $X2=9.43 $Y2=0
r657 277 278 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r658 275 378 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=7.3 $Y=0
+ $X2=7.192 $Y2=0
r659 275 277 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.3 $Y=0 $X2=7.59
+ $Y2=0
r660 274 376 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=5.44
+ $X2=5.75 $Y2=5.44
r661 273 274 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.29 $Y=5.44
+ $X2=5.29 $Y2=5.44
r662 271 274 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.45 $Y=5.44
+ $X2=5.29 $Y2=5.44
r663 270 273 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=3.45 $Y=5.44
+ $X2=5.29 $Y2=5.44
r664 270 271 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=5.44
+ $X2=3.45 $Y2=5.44
r665 268 375 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=5.58 $Y=5.44
+ $X2=5.687 $Y2=5.44
r666 268 273 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.58 $Y=5.44
+ $X2=5.29 $Y2=5.44
r667 267 373 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=5.75 $Y2=0
r668 266 267 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r669 264 267 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=5.29 $Y2=0
r670 263 266 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=3.45 $Y=0
+ $X2=5.29 $Y2=0
r671 263 264 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r672 261 372 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=5.58 $Y=0
+ $X2=5.687 $Y2=0
r673 261 266 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.58 $Y=0
+ $X2=5.29 $Y2=0
r674 260 271 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=5.44
+ $X2=3.45 $Y2=5.44
r675 259 260 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=5.44
+ $X2=2.99 $Y2=5.44
r676 257 260 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=5.44
+ $X2=2.99 $Y2=5.44
r677 257 370 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=5.44
+ $X2=0.69 $Y2=5.44
r678 256 259 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=5.44
+ $X2=2.99 $Y2=5.44
r679 256 257 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=5.44
+ $X2=1.15 $Y2=5.44
r680 254 369 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=0.86 $Y=5.44
+ $X2=0.752 $Y2=5.44
r681 254 256 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.86 $Y=5.44
+ $X2=1.15 $Y2=5.44
r682 253 264 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.45 $Y2=0
r683 252 253 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r684 250 253 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.99 $Y2=0
r685 250 367 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r686 249 252 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=0
+ $X2=2.99 $Y2=0
r687 249 250 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r688 247 366 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=0.86 $Y=0
+ $X2=0.752 $Y2=0
r689 247 249 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.86 $Y=0
+ $X2=1.15 $Y2=0
r690 230 356 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=25.53 $Y=5.44
+ $X2=24.61 $Y2=5.44
r691 230 362 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=25.53 $Y=5.44
+ $X2=25.53 $Y2=5.44
r692 229 350 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=25.53 $Y=0
+ $X2=24.61 $Y2=0
r693 229 358 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=25.53 $Y=0
+ $X2=25.53 $Y2=0
r694 228 406 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.55 $Y=5.44
+ $X2=20.01 $Y2=5.44
r695 227 403 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.55 $Y=0
+ $X2=20.01 $Y2=0
r696 226 228 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.09 $Y=5.44
+ $X2=19.55 $Y2=5.44
r697 226 400 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.09 $Y=5.44
+ $X2=18.63 $Y2=5.44
r698 225 227 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.09 $Y=0
+ $X2=19.55 $Y2=0
r699 225 397 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.09 $Y=0
+ $X2=18.63 $Y2=0
r700 224 394 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=5.44
+ $X2=13.57 $Y2=5.44
r701 223 391 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=0
+ $X2=13.57 $Y2=0
r702 222 224 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=5.44
+ $X2=13.11 $Y2=5.44
r703 222 388 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=5.44
+ $X2=12.19 $Y2=5.44
r704 221 223 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.11 $Y2=0
r705 221 385 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=12.19 $Y2=0
r706 220 382 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=5.44
+ $X2=7.13 $Y2=5.44
r707 219 379 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r708 218 220 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=5.44
+ $X2=6.67 $Y2=5.44
r709 218 376 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=5.44
+ $X2=5.75 $Y2=5.44
r710 217 219 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=6.67 $Y2=0
r711 217 373 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=5.75 $Y2=0
r712 216 370 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=5.44
+ $X2=0.69 $Y2=5.44
r713 215 367 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r714 213 355 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=24.9 $Y=5.44
+ $X2=24.61 $Y2=5.44
r715 213 214 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=24.9 $Y=5.44
+ $X2=25.007 $Y2=5.44
r716 212 362 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=25.115 $Y=5.44
+ $X2=25.53 $Y2=5.44
r717 212 214 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=25.115 $Y=5.44
+ $X2=25.007 $Y2=5.44
r718 210 349 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=24.9 $Y=0
+ $X2=24.61 $Y2=0
r719 210 211 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=24.9 $Y=0
+ $X2=25.007 $Y2=0
r720 209 358 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=25.115 $Y=0
+ $X2=25.53 $Y2=0
r721 209 211 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=25.115 $Y=0
+ $X2=25.007 $Y2=0
r722 207 343 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=22.415 $Y=5.44
+ $X2=22.31 $Y2=5.44
r723 207 208 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=22.415 $Y=5.44
+ $X2=22.54 $Y2=5.44
r724 206 352 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=22.665 $Y=5.44
+ $X2=22.77 $Y2=5.44
r725 206 208 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=22.665 $Y=5.44
+ $X2=22.54 $Y2=5.44
r726 204 336 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=22.415 $Y=0
+ $X2=22.31 $Y2=0
r727 204 205 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=22.415 $Y=0
+ $X2=22.54 $Y2=0
r728 203 346 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=22.665 $Y=0
+ $X2=22.77 $Y2=0
r729 203 205 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=22.665 $Y=0
+ $X2=22.54 $Y2=0
r730 201 315 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=15.975 $Y=5.44
+ $X2=15.87 $Y2=5.44
r731 201 202 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.975 $Y=5.44
+ $X2=16.1 $Y2=5.44
r732 200 326 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=16.225 $Y=5.44
+ $X2=16.33 $Y2=5.44
r733 200 202 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.225 $Y=5.44
+ $X2=16.1 $Y2=5.44
r734 198 308 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=15.975 $Y=0
+ $X2=15.87 $Y2=0
r735 198 199 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.975 $Y=0
+ $X2=16.1 $Y2=0
r736 197 319 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=16.225 $Y=0
+ $X2=16.33 $Y2=0
r737 197 199 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.225 $Y=0
+ $X2=16.1 $Y2=0
r738 195 287 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=9.535 $Y=5.44
+ $X2=9.43 $Y2=5.44
r739 195 196 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.535 $Y=5.44
+ $X2=9.66 $Y2=5.44
r740 194 298 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=9.785 $Y=5.44
+ $X2=9.89 $Y2=5.44
r741 194 196 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.785 $Y=5.44
+ $X2=9.66 $Y2=5.44
r742 192 280 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=9.535 $Y=0
+ $X2=9.43 $Y2=0
r743 192 193 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.535 $Y=0
+ $X2=9.66 $Y2=0
r744 191 291 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=9.785 $Y=0
+ $X2=9.89 $Y2=0
r745 191 193 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.785 $Y=0
+ $X2=9.66 $Y2=0
r746 189 259 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.095 $Y=5.44
+ $X2=2.99 $Y2=5.44
r747 189 190 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.095 $Y=5.44
+ $X2=3.22 $Y2=5.44
r748 188 270 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.345 $Y=5.44
+ $X2=3.45 $Y2=5.44
r749 188 190 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.345 $Y=5.44
+ $X2=3.22 $Y2=5.44
r750 186 252 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.095 $Y=0
+ $X2=2.99 $Y2=0
r751 186 187 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.095 $Y=0
+ $X2=3.22 $Y2=0
r752 185 263 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.345 $Y=0
+ $X2=3.45 $Y2=0
r753 185 187 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.345 $Y=0
+ $X2=3.22 $Y2=0
r754 181 214 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=25.007 $Y=5.355
+ $X2=25.007 $Y2=5.44
r755 181 183 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=25.007 $Y=5.355
+ $X2=25.007 $Y2=5.06
r756 177 211 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=25.007 $Y=0.085
+ $X2=25.007 $Y2=0
r757 177 179 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=25.007 $Y=0.085
+ $X2=25.007 $Y2=0.38
r758 173 208 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=22.54 $Y=5.355
+ $X2=22.54 $Y2=5.44
r759 173 175 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=22.54 $Y=5.355
+ $X2=22.54 $Y2=4.945
r760 169 205 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=22.54 $Y=0.085
+ $X2=22.54 $Y2=0
r761 169 171 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=22.54 $Y=0.085
+ $X2=22.54 $Y2=0.495
r762 165 405 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=20.072 $Y=5.355
+ $X2=20.072 $Y2=5.44
r763 165 167 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=20.072 $Y=5.355
+ $X2=20.072 $Y2=5.06
r764 161 402 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=20.072 $Y=0.085
+ $X2=20.072 $Y2=0
r765 161 163 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=20.072 $Y=0.085
+ $X2=20.072 $Y2=0.38
r766 160 399 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=18.675 $Y=5.44
+ $X2=18.567 $Y2=5.44
r767 159 405 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=19.965 $Y=5.44
+ $X2=20.072 $Y2=5.44
r768 159 160 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=19.965 $Y=5.44
+ $X2=18.675 $Y2=5.44
r769 158 396 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=18.675 $Y=0
+ $X2=18.567 $Y2=0
r770 157 402 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=19.965 $Y=0
+ $X2=20.072 $Y2=0
r771 157 158 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=19.965 $Y=0
+ $X2=18.675 $Y2=0
r772 153 399 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=18.567 $Y=5.355
+ $X2=18.567 $Y2=5.44
r773 153 155 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=18.567 $Y=5.355
+ $X2=18.567 $Y2=5.06
r774 149 396 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=18.567 $Y=0.085
+ $X2=18.567 $Y2=0
r775 149 151 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=18.567 $Y=0.085
+ $X2=18.567 $Y2=0.38
r776 145 202 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.1 $Y=5.355
+ $X2=16.1 $Y2=5.44
r777 145 147 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=16.1 $Y=5.355
+ $X2=16.1 $Y2=4.945
r778 141 199 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.1 $Y=0.085
+ $X2=16.1 $Y2=0
r779 141 143 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=16.1 $Y=0.085
+ $X2=16.1 $Y2=0.495
r780 137 393 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=13.632 $Y=5.355
+ $X2=13.632 $Y2=5.44
r781 137 139 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=13.632 $Y=5.355
+ $X2=13.632 $Y2=5.06
r782 133 390 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=13.632 $Y=0.085
+ $X2=13.632 $Y2=0
r783 133 135 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=13.632 $Y=0.085
+ $X2=13.632 $Y2=0.38
r784 132 387 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=12.235 $Y=5.44
+ $X2=12.127 $Y2=5.44
r785 131 393 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=13.525 $Y=5.44
+ $X2=13.632 $Y2=5.44
r786 131 132 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=13.525 $Y=5.44
+ $X2=12.235 $Y2=5.44
r787 130 384 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=12.235 $Y=0
+ $X2=12.127 $Y2=0
r788 129 390 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=13.525 $Y=0
+ $X2=13.632 $Y2=0
r789 129 130 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=13.525 $Y=0
+ $X2=12.235 $Y2=0
r790 125 387 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=12.127 $Y=5.355
+ $X2=12.127 $Y2=5.44
r791 125 127 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=12.127 $Y=5.355
+ $X2=12.127 $Y2=5.06
r792 121 384 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=12.127 $Y=0.085
+ $X2=12.127 $Y2=0
r793 121 123 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=12.127 $Y=0.085
+ $X2=12.127 $Y2=0.38
r794 117 196 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.66 $Y=5.355
+ $X2=9.66 $Y2=5.44
r795 117 119 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=9.66 $Y=5.355
+ $X2=9.66 $Y2=4.945
r796 113 193 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.66 $Y=0.085
+ $X2=9.66 $Y2=0
r797 113 115 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=9.66 $Y=0.085
+ $X2=9.66 $Y2=0.495
r798 109 381 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=7.192 $Y=5.355
+ $X2=7.192 $Y2=5.44
r799 109 111 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=7.192 $Y=5.355
+ $X2=7.192 $Y2=5.06
r800 105 378 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=7.192 $Y=0.085
+ $X2=7.192 $Y2=0
r801 105 107 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=7.192 $Y=0.085
+ $X2=7.192 $Y2=0.38
r802 104 375 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=5.795 $Y=5.44
+ $X2=5.687 $Y2=5.44
r803 103 381 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=7.085 $Y=5.44
+ $X2=7.192 $Y2=5.44
r804 103 104 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=7.085 $Y=5.44
+ $X2=5.795 $Y2=5.44
r805 102 372 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=5.795 $Y=0
+ $X2=5.687 $Y2=0
r806 101 378 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=7.085 $Y=0
+ $X2=7.192 $Y2=0
r807 101 102 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=7.085 $Y=0
+ $X2=5.795 $Y2=0
r808 97 375 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.687 $Y=5.355
+ $X2=5.687 $Y2=5.44
r809 97 99 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=5.687 $Y=5.355
+ $X2=5.687 $Y2=5.06
r810 93 372 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.687 $Y=0.085
+ $X2=5.687 $Y2=0
r811 93 95 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=5.687 $Y=0.085
+ $X2=5.687 $Y2=0.38
r812 89 190 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=5.355
+ $X2=3.22 $Y2=5.44
r813 89 91 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=3.22 $Y=5.355
+ $X2=3.22 $Y2=4.945
r814 85 187 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=0.085
+ $X2=3.22 $Y2=0
r815 85 87 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=3.22 $Y=0.085
+ $X2=3.22 $Y2=0.495
r816 81 369 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.752 $Y=5.355
+ $X2=0.752 $Y2=5.44
r817 81 83 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=0.752 $Y=5.355
+ $X2=0.752 $Y2=5.06
r818 77 366 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.752 $Y=0.085
+ $X2=0.752 $Y2=0
r819 77 79 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=0.752 $Y=0.085
+ $X2=0.752 $Y2=0.38
r820 24 183 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=24.895
+ $Y=4.555 $X2=25.03 $Y2=5.06
r821 23 179 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=24.895
+ $Y=0.235 $X2=25.03 $Y2=0.38
r822 22 175 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=22.405
+ $Y=4.685 $X2=22.54 $Y2=4.945
r823 21 171 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=22.405
+ $Y=0.235 $X2=22.54 $Y2=0.495
r824 20 167 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=19.915
+ $Y=4.555 $X2=20.05 $Y2=5.06
r825 19 163 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=19.915
+ $Y=0.235 $X2=20.05 $Y2=0.38
r826 18 155 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=18.455
+ $Y=4.555 $X2=18.59 $Y2=5.06
r827 17 151 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=18.455
+ $Y=0.235 $X2=18.59 $Y2=0.38
r828 16 147 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=15.965
+ $Y=4.685 $X2=16.1 $Y2=4.945
r829 15 143 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=15.965
+ $Y=0.235 $X2=16.1 $Y2=0.495
r830 14 139 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=13.475
+ $Y=4.555 $X2=13.61 $Y2=5.06
r831 13 135 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=13.475
+ $Y=0.235 $X2=13.61 $Y2=0.38
r832 12 127 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=12.015
+ $Y=4.555 $X2=12.15 $Y2=5.06
r833 11 123 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=12.015
+ $Y=0.235 $X2=12.15 $Y2=0.38
r834 10 119 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=9.525
+ $Y=4.685 $X2=9.66 $Y2=4.945
r835 9 115 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=9.525
+ $Y=0.235 $X2=9.66 $Y2=0.495
r836 8 111 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=7.035
+ $Y=4.555 $X2=7.17 $Y2=5.06
r837 7 107 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.035
+ $Y=0.235 $X2=7.17 $Y2=0.38
r838 6 99 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=5.575
+ $Y=4.555 $X2=5.71 $Y2=5.06
r839 5 95 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.575
+ $Y=0.235 $X2=5.71 $Y2=0.38
r840 4 91 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=3.085
+ $Y=4.685 $X2=3.22 $Y2=4.945
r841 3 87 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=3.085
+ $Y=0.235 $X2=3.22 $Y2=0.495
r842 2 83 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=4.555 $X2=0.73 $Y2=5.06
r843 1 79 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_845_69# 1 2 3 12 14 15 16 18 19 22
c48 16 0 1.81988e-19 $X=5.257 $Y=0.425
r49 20 22 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.13 $Y=0.715
+ $X2=6.13 $Y2=0.38
r50 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.965 $Y=0.8
+ $X2=6.13 $Y2=0.715
r51 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=5.965 $Y=0.8
+ $X2=5.41 $Y2=0.8
r52 17 19 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=5.257 $Y=0.715
+ $X2=5.41 $Y2=0.8
r53 16 25 2.71076 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.257 $Y=0.425
+ $X2=5.257 $Y2=0.34
r54 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=5.257 $Y=0.425
+ $X2=5.257 $Y2=0.715
r55 14 25 4.84748 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.105 $Y=0.34
+ $X2=5.257 $Y2=0.34
r56 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.105 $Y=0.34
+ $X2=4.435 $Y2=0.34
r57 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.35 $Y=0.425
+ $X2=4.435 $Y2=0.34
r58 10 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.35 $Y=0.425
+ $X2=4.35 $Y2=0.605
r59 3 22 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.995
+ $Y=0.235 $X2=6.13 $Y2=0.38
r60 2 25 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=5.055
+ $Y=0.345 $X2=5.265 $Y2=0.42
r61 1 12 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=4.225
+ $Y=0.345 $X2=4.35 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_845_915# 1 2 3 12 14 15 16 18 25
r47 19 23 4.70351 $w=1.7e-07 $l=1.62693e-07 $layer=LI1_cond $X=5.41 $Y=4.64
+ $X2=5.257 $Y2=4.62
r48 18 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.965 $Y=4.64
+ $X2=6.13 $Y2=4.64
r49 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=5.965 $Y=4.64
+ $X2=5.41 $Y2=4.64
r50 16 23 2.85473 $w=3.05e-07 $l=1.05e-07 $layer=LI1_cond $X=5.257 $Y=4.725
+ $X2=5.257 $Y2=4.62
r51 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=5.257 $Y=4.725
+ $X2=5.257 $Y2=5.015
r52 14 17 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=5.105 $Y=5.1
+ $X2=5.257 $Y2=5.015
r53 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.105 $Y=5.1
+ $X2=4.435 $Y2=5.1
r54 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.35 $Y=5.015
+ $X2=4.435 $Y2=5.1
r55 10 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.35 $Y=5.015
+ $X2=4.35 $Y2=4.835
r56 3 25 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=5.995
+ $Y=4.555 $X2=6.13 $Y2=4.72
r57 2 23 91 $w=1.7e-07 $l=2.57196e-07 $layer=licon1_NDIFF $count=2 $X=5.055
+ $Y=4.575 $X2=5.265 $Y2=4.68
r58 1 12 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=4.225
+ $Y=4.575 $X2=4.35 $Y2=4.835
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1315_47# 1 2 3 12 14 15 16 18 22
c44 16 0 1.81988e-19 $X=7.622 $Y=0.425
r45 20 22 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.53 $Y=0.425
+ $X2=8.53 $Y2=0.605
r46 19 25 4.85887 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.775 $Y=0.34
+ $X2=7.622 $Y2=0.34
r47 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.445 $Y=0.34
+ $X2=8.53 $Y2=0.425
r48 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.445 $Y=0.34
+ $X2=7.775 $Y2=0.34
r49 16 25 2.69937 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.622 $Y=0.425
+ $X2=7.622 $Y2=0.34
r50 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=7.622 $Y=0.425
+ $X2=7.622 $Y2=0.715
r51 14 17 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=7.47 $Y=0.8
+ $X2=7.622 $Y2=0.715
r52 14 15 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=7.47 $Y=0.8
+ $X2=6.915 $Y2=0.8
r53 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.75 $Y=0.715
+ $X2=6.915 $Y2=0.8
r54 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.75 $Y=0.715
+ $X2=6.75 $Y2=0.38
r55 3 22 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=8.395
+ $Y=0.345 $X2=8.53 $Y2=0.605
r56 2 25 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=7.455
+ $Y=0.235 $X2=7.615 $Y2=0.42
r57 1 12 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=6.575
+ $Y=0.235 $X2=6.75 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1315_911# 1 2 3 12 14 16 17 20 23
c44 17 0 1.81988e-19 $X=7.775 $Y=5.1
r45 18 20 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.53 $Y=5.015
+ $X2=8.53 $Y2=4.835
r46 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.445 $Y=5.1
+ $X2=8.53 $Y2=5.015
r47 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.445 $Y=5.1
+ $X2=7.775 $Y2=5.1
r48 15 17 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=7.622 $Y=5.015
+ $X2=7.775 $Y2=5.1
r49 14 25 2.86504 $w=3.05e-07 $l=1.05e-07 $layer=LI1_cond $X=7.622 $Y=4.725
+ $X2=7.622 $Y2=4.62
r50 14 15 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=7.622 $Y=4.725
+ $X2=7.622 $Y2=5.015
r51 13 23 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.915 $Y=4.64
+ $X2=6.75 $Y2=4.64
r52 12 25 4.6932 $w=1.7e-07 $l=1.61691e-07 $layer=LI1_cond $X=7.47 $Y=4.64
+ $X2=7.622 $Y2=4.62
r53 12 13 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=7.47 $Y=4.64
+ $X2=6.915 $Y2=4.64
r54 3 20 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=8.395
+ $Y=4.575 $X2=8.53 $Y2=4.835
r55 2 25 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=7.455
+ $Y=4.555 $X2=7.615 $Y2=4.68
r56 1 23 91 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_NDIFF $count=2 $X=6.575
+ $Y=4.555 $X2=6.75 $Y2=4.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2133_69# 1 2 3 12 14 15 16 18 19 22
c48 16 0 1.81988e-19 $X=11.697 $Y=0.425
r49 20 22 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=12.57 $Y=0.715
+ $X2=12.57 $Y2=0.38
r50 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.405 $Y=0.8
+ $X2=12.57 $Y2=0.715
r51 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=12.405 $Y=0.8
+ $X2=11.85 $Y2=0.8
r52 17 19 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=11.697 $Y=0.715
+ $X2=11.85 $Y2=0.8
r53 16 25 2.71076 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=11.697 $Y=0.425
+ $X2=11.697 $Y2=0.34
r54 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=11.697 $Y=0.425
+ $X2=11.697 $Y2=0.715
r55 14 25 4.84748 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=11.545 $Y=0.34
+ $X2=11.697 $Y2=0.34
r56 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.545 $Y=0.34
+ $X2=10.875 $Y2=0.34
r57 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.79 $Y=0.425
+ $X2=10.875 $Y2=0.34
r58 10 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=10.79 $Y=0.425
+ $X2=10.79 $Y2=0.605
r59 3 22 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=12.435
+ $Y=0.235 $X2=12.57 $Y2=0.38
r60 2 25 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=11.495
+ $Y=0.345 $X2=11.705 $Y2=0.42
r61 1 12 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=10.665
+ $Y=0.345 $X2=10.79 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2133_915# 1 2 3 12 14 15 16 18 25
r47 19 23 4.70351 $w=1.7e-07 $l=1.62693e-07 $layer=LI1_cond $X=11.85 $Y=4.64
+ $X2=11.697 $Y2=4.62
r48 18 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.405 $Y=4.64
+ $X2=12.57 $Y2=4.64
r49 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=12.405 $Y=4.64
+ $X2=11.85 $Y2=4.64
r50 16 23 2.85473 $w=3.05e-07 $l=1.05e-07 $layer=LI1_cond $X=11.697 $Y=4.725
+ $X2=11.697 $Y2=4.62
r51 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=11.697 $Y=4.725
+ $X2=11.697 $Y2=5.015
r52 14 17 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=11.545 $Y=5.1
+ $X2=11.697 $Y2=5.015
r53 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.545 $Y=5.1
+ $X2=10.875 $Y2=5.1
r54 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.79 $Y=5.015
+ $X2=10.875 $Y2=5.1
r55 10 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=10.79 $Y=5.015
+ $X2=10.79 $Y2=4.835
r56 3 25 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=12.435
+ $Y=4.555 $X2=12.57 $Y2=4.72
r57 2 23 91 $w=1.7e-07 $l=2.57196e-07 $layer=licon1_NDIFF $count=2 $X=11.495
+ $Y=4.575 $X2=11.705 $Y2=4.68
r58 1 12 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=10.665
+ $Y=4.575 $X2=10.79 $Y2=4.835
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2603_47# 1 2 3 12 14 15 16 18 22
c44 16 0 1.81988e-19 $X=14.062 $Y=0.425
r45 20 22 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=14.97 $Y=0.425
+ $X2=14.97 $Y2=0.605
r46 19 25 4.85887 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=14.215 $Y=0.34
+ $X2=14.062 $Y2=0.34
r47 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.885 $Y=0.34
+ $X2=14.97 $Y2=0.425
r48 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=14.885 $Y=0.34
+ $X2=14.215 $Y2=0.34
r49 16 25 2.69937 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=14.062 $Y=0.425
+ $X2=14.062 $Y2=0.34
r50 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=14.062 $Y=0.425
+ $X2=14.062 $Y2=0.715
r51 14 17 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=13.91 $Y=0.8
+ $X2=14.062 $Y2=0.715
r52 14 15 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=13.91 $Y=0.8
+ $X2=13.355 $Y2=0.8
r53 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.19 $Y=0.715
+ $X2=13.355 $Y2=0.8
r54 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=13.19 $Y=0.715
+ $X2=13.19 $Y2=0.38
r55 3 22 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=14.835
+ $Y=0.345 $X2=14.97 $Y2=0.605
r56 2 25 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=13.895
+ $Y=0.235 $X2=14.055 $Y2=0.42
r57 1 12 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=13.015
+ $Y=0.235 $X2=13.19 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2603_911# 1 2 3 12 14 16 17 20 23
c44 17 0 1.81988e-19 $X=14.215 $Y=5.1
r45 18 20 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=14.97 $Y=5.015
+ $X2=14.97 $Y2=4.835
r46 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.885 $Y=5.1
+ $X2=14.97 $Y2=5.015
r47 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=14.885 $Y=5.1
+ $X2=14.215 $Y2=5.1
r48 15 17 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=14.062 $Y=5.015
+ $X2=14.215 $Y2=5.1
r49 14 25 2.86504 $w=3.05e-07 $l=1.05e-07 $layer=LI1_cond $X=14.062 $Y=4.725
+ $X2=14.062 $Y2=4.62
r50 14 15 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=14.062 $Y=4.725
+ $X2=14.062 $Y2=5.015
r51 13 23 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.355 $Y=4.64
+ $X2=13.19 $Y2=4.64
r52 12 25 4.6932 $w=1.7e-07 $l=1.61691e-07 $layer=LI1_cond $X=13.91 $Y=4.64
+ $X2=14.062 $Y2=4.62
r53 12 13 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=13.91 $Y=4.64
+ $X2=13.355 $Y2=4.64
r54 3 20 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=14.835
+ $Y=4.575 $X2=14.97 $Y2=4.835
r55 2 25 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=13.895
+ $Y=4.555 $X2=14.055 $Y2=4.68
r56 1 23 91 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_NDIFF $count=2 $X=13.015
+ $Y=4.555 $X2=13.19 $Y2=4.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3421_69# 1 2 3 12 14 15 16 18 19 22
c48 16 0 1.81988e-19 $X=18.137 $Y=0.425
r49 20 22 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=19.01 $Y=0.715
+ $X2=19.01 $Y2=0.38
r50 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=18.845 $Y=0.8
+ $X2=19.01 $Y2=0.715
r51 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=18.845 $Y=0.8
+ $X2=18.29 $Y2=0.8
r52 17 19 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=18.137 $Y=0.715
+ $X2=18.29 $Y2=0.8
r53 16 25 2.71076 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=18.137 $Y=0.425
+ $X2=18.137 $Y2=0.34
r54 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=18.137 $Y=0.425
+ $X2=18.137 $Y2=0.715
r55 14 25 4.84748 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=17.985 $Y=0.34
+ $X2=18.137 $Y2=0.34
r56 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=17.985 $Y=0.34
+ $X2=17.315 $Y2=0.34
r57 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=17.23 $Y=0.425
+ $X2=17.315 $Y2=0.34
r58 10 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=17.23 $Y=0.425
+ $X2=17.23 $Y2=0.605
r59 3 22 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=18.875
+ $Y=0.235 $X2=19.01 $Y2=0.38
r60 2 25 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=17.935
+ $Y=0.345 $X2=18.145 $Y2=0.42
r61 1 12 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=17.105
+ $Y=0.345 $X2=17.23 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3421_915# 1 2 3 12 14 15 16 18 25
r47 19 23 4.70351 $w=1.7e-07 $l=1.62693e-07 $layer=LI1_cond $X=18.29 $Y=4.64
+ $X2=18.137 $Y2=4.62
r48 18 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.845 $Y=4.64
+ $X2=19.01 $Y2=4.64
r49 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=18.845 $Y=4.64
+ $X2=18.29 $Y2=4.64
r50 16 23 2.85473 $w=3.05e-07 $l=1.05e-07 $layer=LI1_cond $X=18.137 $Y=4.725
+ $X2=18.137 $Y2=4.62
r51 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=18.137 $Y=4.725
+ $X2=18.137 $Y2=5.015
r52 14 17 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=17.985 $Y=5.1
+ $X2=18.137 $Y2=5.015
r53 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=17.985 $Y=5.1
+ $X2=17.315 $Y2=5.1
r54 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=17.23 $Y=5.015
+ $X2=17.315 $Y2=5.1
r55 10 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=17.23 $Y=5.015
+ $X2=17.23 $Y2=4.835
r56 3 25 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=18.875
+ $Y=4.555 $X2=19.01 $Y2=4.72
r57 2 23 91 $w=1.7e-07 $l=2.57196e-07 $layer=licon1_NDIFF $count=2 $X=17.935
+ $Y=4.575 $X2=18.145 $Y2=4.68
r58 1 12 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=17.105
+ $Y=4.575 $X2=17.23 $Y2=4.835
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3891_47# 1 2 3 12 14 15 16 18 22
c44 16 0 1.81988e-19 $X=20.502 $Y=0.425
r45 20 22 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=21.41 $Y=0.425
+ $X2=21.41 $Y2=0.605
r46 19 25 4.85887 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=20.655 $Y=0.34
+ $X2=20.502 $Y2=0.34
r47 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=21.325 $Y=0.34
+ $X2=21.41 $Y2=0.425
r48 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=21.325 $Y=0.34
+ $X2=20.655 $Y2=0.34
r49 16 25 2.69937 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=20.502 $Y=0.425
+ $X2=20.502 $Y2=0.34
r50 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=20.502 $Y=0.425
+ $X2=20.502 $Y2=0.715
r51 14 17 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=20.35 $Y=0.8
+ $X2=20.502 $Y2=0.715
r52 14 15 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=20.35 $Y=0.8
+ $X2=19.795 $Y2=0.8
r53 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=19.63 $Y=0.715
+ $X2=19.795 $Y2=0.8
r54 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=19.63 $Y=0.715
+ $X2=19.63 $Y2=0.38
r55 3 22 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=21.275
+ $Y=0.345 $X2=21.41 $Y2=0.605
r56 2 25 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=20.335
+ $Y=0.235 $X2=20.495 $Y2=0.42
r57 1 12 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=19.455
+ $Y=0.235 $X2=19.63 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3891_911# 1 2 3 12 14 16 17 20 23
c44 17 0 1.81988e-19 $X=20.655 $Y=5.1
r45 18 20 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=21.41 $Y=5.015
+ $X2=21.41 $Y2=4.835
r46 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=21.325 $Y=5.1
+ $X2=21.41 $Y2=5.015
r47 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=21.325 $Y=5.1
+ $X2=20.655 $Y2=5.1
r48 15 17 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=20.502 $Y=5.015
+ $X2=20.655 $Y2=5.1
r49 14 25 2.86504 $w=3.05e-07 $l=1.05e-07 $layer=LI1_cond $X=20.502 $Y=4.725
+ $X2=20.502 $Y2=4.62
r50 14 15 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=20.502 $Y=4.725
+ $X2=20.502 $Y2=5.015
r51 13 23 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=19.795 $Y=4.64
+ $X2=19.63 $Y2=4.64
r52 12 25 4.6932 $w=1.7e-07 $l=1.61691e-07 $layer=LI1_cond $X=20.35 $Y=4.64
+ $X2=20.502 $Y2=4.62
r53 12 13 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=20.35 $Y=4.64
+ $X2=19.795 $Y2=4.64
r54 3 20 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=21.275
+ $Y=4.575 $X2=21.41 $Y2=4.835
r55 2 25 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=20.335
+ $Y=4.555 $X2=20.495 $Y2=4.68
r56 1 23 91 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_NDIFF $count=2 $X=19.455
+ $Y=4.555 $X2=19.63 $Y2=4.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4709_69# 1 2 3 12 14 15 16 18 19 22
c46 16 0 1.81988e-19 $X=24.577 $Y=0.425
r47 20 22 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=25.45 $Y=0.715
+ $X2=25.45 $Y2=0.38
r48 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=25.285 $Y=0.8
+ $X2=25.45 $Y2=0.715
r49 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=25.285 $Y=0.8
+ $X2=24.73 $Y2=0.8
r50 17 19 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=24.577 $Y=0.715
+ $X2=24.73 $Y2=0.8
r51 16 25 2.71076 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=24.577 $Y=0.425
+ $X2=24.577 $Y2=0.34
r52 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=24.577 $Y=0.425
+ $X2=24.577 $Y2=0.715
r53 14 25 4.84748 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=24.425 $Y=0.34
+ $X2=24.577 $Y2=0.34
r54 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=24.425 $Y=0.34
+ $X2=23.755 $Y2=0.34
r55 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=23.67 $Y=0.425
+ $X2=23.755 $Y2=0.34
r56 10 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=23.67 $Y=0.425
+ $X2=23.67 $Y2=0.605
r57 3 22 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=25.315
+ $Y=0.235 $X2=25.45 $Y2=0.38
r58 2 25 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=24.375
+ $Y=0.345 $X2=24.585 $Y2=0.42
r59 1 12 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=23.545
+ $Y=0.345 $X2=23.67 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4709_915# 1 2 3 12 14 15 16 18 25
r46 19 23 4.70351 $w=1.7e-07 $l=1.62693e-07 $layer=LI1_cond $X=24.73 $Y=4.64
+ $X2=24.577 $Y2=4.62
r47 18 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=25.285 $Y=4.64
+ $X2=25.45 $Y2=4.64
r48 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=25.285 $Y=4.64
+ $X2=24.73 $Y2=4.64
r49 16 23 2.85473 $w=3.05e-07 $l=1.05e-07 $layer=LI1_cond $X=24.577 $Y=4.725
+ $X2=24.577 $Y2=4.62
r50 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=24.577 $Y=4.725
+ $X2=24.577 $Y2=5.015
r51 14 17 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=24.425 $Y=5.1
+ $X2=24.577 $Y2=5.015
r52 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=24.425 $Y=5.1
+ $X2=23.755 $Y2=5.1
r53 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=23.67 $Y=5.015
+ $X2=23.755 $Y2=5.1
r54 10 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=23.67 $Y=5.015
+ $X2=23.67 $Y2=4.835
r55 3 25 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=25.315
+ $Y=4.555 $X2=25.45 $Y2=4.72
r56 2 23 91 $w=1.7e-07 $l=2.57196e-07 $layer=licon1_NDIFF $count=2 $X=24.375
+ $Y=4.575 $X2=24.585 $Y2=4.68
r57 1 12 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=23.545
+ $Y=4.575 $X2=23.67 $Y2=4.835
.ends

