* File: sky130_fd_sc_hdll__isobufsrc_8.pxi.spice
* Created: Wed Sep  2 08:34:01 2020
* 
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%A N_A_c_137_n N_A_M1001_g N_A_c_132_n
+ N_A_M1018_g N_A_c_138_n N_A_M1014_g N_A_c_133_n N_A_M1027_g A N_A_c_135_n
+ N_A_c_136_n PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%A
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%A_117_297# N_A_117_297#_M1018_s
+ N_A_117_297#_M1001_s N_A_117_297#_c_177_n N_A_117_297#_M1006_g
+ N_A_117_297#_c_187_n N_A_117_297#_M1000_g N_A_117_297#_c_178_n
+ N_A_117_297#_M1008_g N_A_117_297#_c_188_n N_A_117_297#_M1002_g
+ N_A_117_297#_c_179_n N_A_117_297#_M1011_g N_A_117_297#_c_189_n
+ N_A_117_297#_M1004_g N_A_117_297#_c_180_n N_A_117_297#_M1019_g
+ N_A_117_297#_c_190_n N_A_117_297#_M1005_g N_A_117_297#_c_181_n
+ N_A_117_297#_M1020_g N_A_117_297#_c_191_n N_A_117_297#_M1015_g
+ N_A_117_297#_c_182_n N_A_117_297#_M1026_g N_A_117_297#_c_192_n
+ N_A_117_297#_M1017_g N_A_117_297#_c_183_n N_A_117_297#_M1029_g
+ N_A_117_297#_c_193_n N_A_117_297#_M1023_g N_A_117_297#_c_194_n
+ N_A_117_297#_M1031_g N_A_117_297#_c_184_n N_A_117_297#_M1032_g
+ N_A_117_297#_c_199_n N_A_117_297#_c_201_n N_A_117_297#_c_185_n
+ N_A_117_297#_c_195_n N_A_117_297#_c_196_n N_A_117_297#_c_212_n
+ N_A_117_297#_c_186_n PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%A_117_297#
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%SLEEP N_SLEEP_c_351_n N_SLEEP_M1009_g
+ N_SLEEP_c_360_n N_SLEEP_M1003_g N_SLEEP_c_352_n N_SLEEP_M1010_g
+ N_SLEEP_c_361_n N_SLEEP_M1007_g N_SLEEP_c_353_n N_SLEEP_M1012_g
+ N_SLEEP_c_362_n N_SLEEP_M1016_g N_SLEEP_c_354_n N_SLEEP_M1013_g
+ N_SLEEP_c_363_n N_SLEEP_M1021_g N_SLEEP_c_355_n N_SLEEP_M1022_g
+ N_SLEEP_c_364_n N_SLEEP_M1025_g N_SLEEP_c_356_n N_SLEEP_M1024_g
+ N_SLEEP_c_365_n N_SLEEP_M1028_g N_SLEEP_c_357_n N_SLEEP_M1030_g
+ N_SLEEP_c_366_n N_SLEEP_M1034_g N_SLEEP_c_367_n N_SLEEP_M1035_g
+ N_SLEEP_c_358_n N_SLEEP_M1033_g SLEEP N_SLEEP_c_371_n N_SLEEP_c_359_n SLEEP
+ PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%SLEEP
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%VPWR N_VPWR_M1001_d N_VPWR_M1014_d
+ N_VPWR_M1000_d N_VPWR_M1004_d N_VPWR_M1015_d N_VPWR_M1023_d N_VPWR_c_491_n
+ N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_494_n N_VPWR_c_495_n N_VPWR_c_496_n
+ N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_500_n N_VPWR_c_501_n
+ N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n N_VPWR_c_506_n
+ N_VPWR_c_507_n VPWR N_VPWR_c_508_n N_VPWR_c_490_n
+ PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%VPWR
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%A_345_297# N_A_345_297#_M1000_s
+ N_A_345_297#_M1002_s N_A_345_297#_M1005_s N_A_345_297#_M1017_s
+ N_A_345_297#_M1031_s N_A_345_297#_M1007_d N_A_345_297#_M1021_d
+ N_A_345_297#_M1028_d N_A_345_297#_M1035_d N_A_345_297#_c_614_n
+ N_A_345_297#_c_615_n N_A_345_297#_c_616_n N_A_345_297#_c_672_n
+ N_A_345_297#_c_617_n N_A_345_297#_c_676_n N_A_345_297#_c_618_n
+ N_A_345_297#_c_680_n N_A_345_297#_c_619_n N_A_345_297#_c_620_n
+ N_A_345_297#_c_684_n N_A_345_297#_c_649_n N_A_345_297#_c_707_p
+ N_A_345_297#_c_651_n N_A_345_297#_c_711_p N_A_345_297#_c_653_n
+ N_A_345_297#_c_714_p N_A_345_297#_c_655_n N_A_345_297#_c_717_p
+ N_A_345_297#_c_621_n N_A_345_297#_c_622_n N_A_345_297#_c_623_n
+ N_A_345_297#_c_694_n N_A_345_297#_c_696_n N_A_345_297#_c_698_n
+ PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%A_345_297#
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%X N_X_M1006_d N_X_M1011_d N_X_M1020_d
+ N_X_M1029_d N_X_M1009_d N_X_M1012_d N_X_M1022_d N_X_M1030_d N_X_M1003_s
+ N_X_M1016_s N_X_M1025_s N_X_M1034_s N_X_c_741_n N_X_c_718_n N_X_c_719_n
+ N_X_c_752_n N_X_c_720_n N_X_c_760_n N_X_c_721_n N_X_c_768_n N_X_c_722_n
+ N_X_c_772_n N_X_c_859_n N_X_c_734_n N_X_c_735_n N_X_c_723_n N_X_c_800_n
+ N_X_c_863_n N_X_c_736_n N_X_c_724_n N_X_c_812_n N_X_c_866_n N_X_c_737_n
+ N_X_c_725_n N_X_c_869_n N_X_c_726_n N_X_c_727_n N_X_c_728_n N_X_c_729_n
+ N_X_c_730_n N_X_c_738_n N_X_c_731_n N_X_c_739_n N_X_c_732_n X
+ PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%X
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%VGND N_VGND_M1018_d N_VGND_M1027_d
+ N_VGND_M1008_s N_VGND_M1019_s N_VGND_M1026_s N_VGND_M1032_s N_VGND_M1010_s
+ N_VGND_M1013_s N_VGND_M1024_s N_VGND_M1033_s N_VGND_c_940_n N_VGND_c_941_n
+ N_VGND_c_942_n N_VGND_c_943_n N_VGND_c_944_n N_VGND_c_945_n N_VGND_c_946_n
+ N_VGND_c_947_n N_VGND_c_948_n N_VGND_c_949_n N_VGND_c_950_n N_VGND_c_951_n
+ N_VGND_c_952_n N_VGND_c_953_n N_VGND_c_954_n N_VGND_c_955_n N_VGND_c_956_n
+ N_VGND_c_957_n N_VGND_c_958_n N_VGND_c_959_n N_VGND_c_960_n N_VGND_c_961_n
+ N_VGND_c_962_n N_VGND_c_963_n N_VGND_c_964_n N_VGND_c_965_n N_VGND_c_966_n
+ VGND N_VGND_c_967_n N_VGND_c_968_n N_VGND_c_969_n N_VGND_c_970_n
+ PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%VGND
cc_1 VNB N_A_c_132_n 0.019708f $X=-0.19 $Y=-0.24 $X2=0.81 $Y2=0.995
cc_2 VNB N_A_c_133_n 0.0189049f $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=0.995
cc_3 VNB A 0.0409628f $X=-0.19 $Y=-0.24 $X2=0.115 $Y2=1.105
cc_4 VNB N_A_c_135_n 0.0102908f $X=-0.19 $Y=-0.24 $X2=0.29 $Y2=1.16
cc_5 VNB N_A_c_136_n 0.081451f $X=-0.19 $Y=-0.24 $X2=1.015 $Y2=1.202
cc_6 VNB N_A_117_297#_c_177_n 0.0192774f $X=-0.19 $Y=-0.24 $X2=1.015 $Y2=1.41
cc_7 VNB N_A_117_297#_c_178_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_117_297#_c_179_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.29 $Y2=1.16
cc_9 VNB N_A_117_297#_c_180_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_117_297#_c_181_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_117_297#_c_182_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_117_297#_c_183_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_117_297#_c_184_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_117_297#_c_185_n 0.0255745f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_117_297#_c_186_n 0.15153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_SLEEP_c_351_n 0.0164943f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_17 VNB N_SLEEP_c_352_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=1.015 $Y2=1.41
cc_18 VNB N_SLEEP_c_353_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_SLEEP_c_354_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.29 $Y2=1.16
cc_20 VNB N_SLEEP_c_355_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_SLEEP_c_356_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_SLEEP_c_357_n 0.0171931f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_SLEEP_c_358_n 0.0203186f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_SLEEP_c_359_n 0.1537f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_490_n 0.402575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_X_c_718_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_719_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_X_c_720_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_X_c_721_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_X_c_722_n 0.0043236f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_X_c_723_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_X_c_724_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_X_c_725_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_X_c_726_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_X_c_727_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_X_c_728_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_X_c_729_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_X_c_730_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_X_c_731_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_X_c_732_n 0.0108369f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB X 0.0181686f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_940_n 0.00708452f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_941_n 0.0119006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_942_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_943_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_944_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_945_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_946_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_947_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_948_n 0.00467908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_949_n 0.0100782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_950_n 0.0183426f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_951_n 0.015432f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_952_n 0.00422832f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_953_n 0.0198149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_954_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_955_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_956_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_957_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_958_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_959_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_960_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_961_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_962_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_963_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_964_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_965_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_966_n 0.00323927f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_967_n 0.019881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_968_n 0.0192963f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_969_n 0.0098064f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_970_n 0.450337f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VPB N_A_c_137_n 0.0205299f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_74 VPB N_A_c_138_n 0.0203504f $X=-0.19 $Y=1.305 $X2=1.015 $Y2=1.41
cc_75 VPB N_A_c_136_n 0.04377f $X=-0.19 $Y=1.305 $X2=1.015 $Y2=1.202
cc_76 VPB N_A_117_297#_c_187_n 0.0203443f $X=-0.19 $Y=1.305 $X2=1.28 $Y2=0.995
cc_77 VPB N_A_117_297#_c_188_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_117_297#_c_189_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.015 $Y2=1.202
cc_79 VPB N_A_117_297#_c_190_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_117_297#_c_191_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_117_297#_c_192_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_117_297#_c_193_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_117_297#_c_194_n 0.0161059f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_117_297#_c_195_n 0.00134342f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_117_297#_c_196_n 0.00124937f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_117_297#_c_186_n 0.0992988f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_SLEEP_c_360_n 0.0164196f $X=-0.19 $Y=1.305 $X2=0.81 $Y2=0.995
cc_88 VPB N_SLEEP_c_361_n 0.0158911f $X=-0.19 $Y=1.305 $X2=1.28 $Y2=0.995
cc_89 VPB N_SLEEP_c_362_n 0.0158911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_SLEEP_c_363_n 0.0158911f $X=-0.19 $Y=1.305 $X2=1.015 $Y2=1.202
cc_91 VPB N_SLEEP_c_364_n 0.0158911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_SLEEP_c_365_n 0.0158911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_SLEEP_c_366_n 0.0158911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_SLEEP_c_367_n 0.0192434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_SLEEP_c_359_n 0.0978077f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_491_n 0.0103907f $X=-0.19 $Y=1.305 $X2=0.29 $Y2=1.16
cc_97 VPB N_VPWR_c_492_n 0.0434765f $X=-0.19 $Y=1.305 $X2=0.81 $Y2=1.202
cc_98 VPB N_VPWR_c_493_n 0.0172172f $X=-0.19 $Y=1.305 $X2=0.29 $Y2=1.175
cc_99 VPB N_VPWR_c_494_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_495_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_496_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_497_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_498_n 0.0217449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_499_n 0.00564836f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_500_n 0.0209703f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_501_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_502_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_503_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_504_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_505_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_506_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_507_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_508_n 0.102558f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_490_n 0.0565044f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_345_297#_c_614_n 0.00522845f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_345_297#_c_615_n 0.00826138f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_345_297#_c_616_n 0.00196986f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_345_297#_c_617_n 0.00194026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_345_297#_c_618_n 0.00194026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_345_297#_c_619_n 0.00196986f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_345_297#_c_620_n 0.00410164f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_345_297#_c_621_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_345_297#_c_622_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_345_297#_c_623_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_X_c_734_n 0.00192677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_X_c_735_n 0.00188018f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_X_c_736_n 0.00192677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_X_c_737_n 0.00192677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_X_c_738_n 0.0014926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_X_c_739_n 0.0014926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB X 0.017754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 N_A_c_133_n N_A_117_297#_c_177_n 0.00524218f $X=1.28 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_c_137_n N_A_117_297#_c_199_n 0.0120954f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_c_138_n N_A_117_297#_c_199_n 0.00995304f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_c_132_n N_A_117_297#_c_201_n 0.0095611f $X=0.81 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_c_133_n N_A_117_297#_c_201_n 0.0134441f $X=1.28 $Y=0.995 $X2=0 $Y2=0
cc_137 A N_A_117_297#_c_201_n 0.00504935f $X=0.115 $Y=1.105 $X2=0 $Y2=0
cc_138 N_A_c_136_n N_A_117_297#_c_201_n 0.0105872f $X=1.015 $Y=1.202 $X2=0 $Y2=0
cc_139 N_A_c_136_n N_A_117_297#_c_185_n 0.0127213f $X=1.015 $Y=1.202 $X2=0 $Y2=0
cc_140 N_A_c_137_n N_A_117_297#_c_195_n 0.00514095f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_c_138_n N_A_117_297#_c_195_n 0.00306149f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_c_136_n N_A_117_297#_c_195_n 0.00464693f $X=1.015 $Y=1.202 $X2=0
+ $Y2=0
cc_143 N_A_c_137_n N_A_117_297#_c_196_n 0.00102919f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_138_n N_A_117_297#_c_196_n 0.00220819f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_c_136_n N_A_117_297#_c_196_n 0.0155462f $X=1.015 $Y=1.202 $X2=0 $Y2=0
cc_146 N_A_c_135_n N_A_117_297#_c_212_n 0.0144402f $X=0.29 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_c_136_n N_A_117_297#_c_212_n 0.033704f $X=1.015 $Y=1.202 $X2=0 $Y2=0
cc_148 N_A_c_136_n N_A_117_297#_c_186_n 0.00524218f $X=1.015 $Y=1.202 $X2=0
+ $Y2=0
cc_149 N_A_c_137_n N_VPWR_c_492_n 0.00833409f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_c_135_n N_VPWR_c_492_n 0.0180017f $X=0.29 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_c_136_n N_VPWR_c_492_n 0.00462085f $X=1.015 $Y=1.202 $X2=0 $Y2=0
cc_152 N_A_c_138_n N_VPWR_c_493_n 0.00947717f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_c_136_n N_VPWR_c_493_n 0.0053981f $X=1.015 $Y=1.202 $X2=0 $Y2=0
cc_154 N_A_c_137_n N_VPWR_c_498_n 0.00597712f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_c_138_n N_VPWR_c_498_n 0.00673617f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_c_137_n N_VPWR_c_490_n 0.0110282f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_c_138_n N_VPWR_c_490_n 0.0132483f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_c_132_n N_VGND_c_940_n 0.00484352f $X=0.81 $Y=0.995 $X2=0 $Y2=0
cc_159 A N_VGND_c_940_n 0.0493999f $X=0.115 $Y=1.105 $X2=0 $Y2=0
cc_160 N_A_c_135_n N_VGND_c_940_n 0.001559f $X=0.29 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A_c_136_n N_VGND_c_940_n 0.00740052f $X=1.015 $Y=1.202 $X2=0 $Y2=0
cc_162 N_A_c_133_n N_VGND_c_941_n 0.00642784f $X=1.28 $Y=0.995 $X2=0 $Y2=0
cc_163 A N_VGND_c_951_n 0.0163465f $X=0.115 $Y=1.105 $X2=0 $Y2=0
cc_164 N_A_c_132_n N_VGND_c_967_n 0.00571722f $X=0.81 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_c_133_n N_VGND_c_967_n 0.00541359f $X=1.28 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A_c_132_n N_VGND_c_970_n 0.0116441f $X=0.81 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_c_133_n N_VGND_c_970_n 0.0104346f $X=1.28 $Y=0.995 $X2=0 $Y2=0
cc_168 A N_VGND_c_970_n 0.00878068f $X=0.115 $Y=1.105 $X2=0 $Y2=0
cc_169 N_A_117_297#_c_184_n N_SLEEP_c_351_n 0.0244381f $X=5.42 $Y=0.995
+ $X2=-0.19 $Y2=-0.24
cc_170 N_A_117_297#_c_194_n N_SLEEP_c_360_n 0.00966468f $X=5.395 $Y=1.41 $X2=0
+ $Y2=0
cc_171 N_A_117_297#_c_185_n N_SLEEP_c_371_n 0.0124677f $X=5.26 $Y=1.16 $X2=0
+ $Y2=0
cc_172 N_A_117_297#_c_186_n N_SLEEP_c_371_n 2.30564e-19 $X=5.395 $Y=1.202 $X2=0
+ $Y2=0
cc_173 N_A_117_297#_c_185_n N_SLEEP_c_359_n 0.00185127f $X=5.26 $Y=1.16 $X2=0
+ $Y2=0
cc_174 N_A_117_297#_c_186_n N_SLEEP_c_359_n 0.0244381f $X=5.395 $Y=1.202 $X2=0
+ $Y2=0
cc_175 N_A_117_297#_c_195_n N_VPWR_c_492_n 0.0775881f $X=0.73 $Y=1.62 $X2=0
+ $Y2=0
cc_176 N_A_117_297#_c_187_n N_VPWR_c_493_n 0.00371652f $X=2.105 $Y=1.41 $X2=0
+ $Y2=0
cc_177 N_A_117_297#_c_185_n N_VPWR_c_493_n 0.0186935f $X=5.26 $Y=1.16 $X2=0
+ $Y2=0
cc_178 N_A_117_297#_c_195_n N_VPWR_c_493_n 0.0650428f $X=0.73 $Y=1.62 $X2=0
+ $Y2=0
cc_179 N_A_117_297#_c_212_n N_VPWR_c_493_n 0.006109f $X=0.98 $Y=1.175 $X2=0
+ $Y2=0
cc_180 N_A_117_297#_c_187_n N_VPWR_c_494_n 0.00300743f $X=2.105 $Y=1.41 $X2=0
+ $Y2=0
cc_181 N_A_117_297#_c_188_n N_VPWR_c_494_n 0.00300743f $X=2.575 $Y=1.41 $X2=0
+ $Y2=0
cc_182 N_A_117_297#_c_189_n N_VPWR_c_495_n 0.00300743f $X=3.045 $Y=1.41 $X2=0
+ $Y2=0
cc_183 N_A_117_297#_c_190_n N_VPWR_c_495_n 0.00300743f $X=3.515 $Y=1.41 $X2=0
+ $Y2=0
cc_184 N_A_117_297#_c_191_n N_VPWR_c_496_n 0.00300743f $X=3.985 $Y=1.41 $X2=0
+ $Y2=0
cc_185 N_A_117_297#_c_192_n N_VPWR_c_496_n 0.00300743f $X=4.455 $Y=1.41 $X2=0
+ $Y2=0
cc_186 N_A_117_297#_c_193_n N_VPWR_c_497_n 0.00300743f $X=4.925 $Y=1.41 $X2=0
+ $Y2=0
cc_187 N_A_117_297#_c_194_n N_VPWR_c_497_n 0.00300743f $X=5.395 $Y=1.41 $X2=0
+ $Y2=0
cc_188 N_A_117_297#_c_199_n N_VPWR_c_498_n 0.0258718f $X=0.73 $Y=2.3 $X2=0 $Y2=0
cc_189 N_A_117_297#_c_187_n N_VPWR_c_500_n 0.00702461f $X=2.105 $Y=1.41 $X2=0
+ $Y2=0
cc_190 N_A_117_297#_c_188_n N_VPWR_c_502_n 0.00702461f $X=2.575 $Y=1.41 $X2=0
+ $Y2=0
cc_191 N_A_117_297#_c_189_n N_VPWR_c_502_n 0.00702461f $X=3.045 $Y=1.41 $X2=0
+ $Y2=0
cc_192 N_A_117_297#_c_190_n N_VPWR_c_504_n 0.00702461f $X=3.515 $Y=1.41 $X2=0
+ $Y2=0
cc_193 N_A_117_297#_c_191_n N_VPWR_c_504_n 0.00702461f $X=3.985 $Y=1.41 $X2=0
+ $Y2=0
cc_194 N_A_117_297#_c_192_n N_VPWR_c_506_n 0.00702461f $X=4.455 $Y=1.41 $X2=0
+ $Y2=0
cc_195 N_A_117_297#_c_193_n N_VPWR_c_506_n 0.00702461f $X=4.925 $Y=1.41 $X2=0
+ $Y2=0
cc_196 N_A_117_297#_c_194_n N_VPWR_c_508_n 0.00702461f $X=5.395 $Y=1.41 $X2=0
+ $Y2=0
cc_197 N_A_117_297#_M1001_s N_VPWR_c_490_n 0.0027141f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_198 N_A_117_297#_c_187_n N_VPWR_c_490_n 0.0136915f $X=2.105 $Y=1.41 $X2=0
+ $Y2=0
cc_199 N_A_117_297#_c_188_n N_VPWR_c_490_n 0.0124092f $X=2.575 $Y=1.41 $X2=0
+ $Y2=0
cc_200 N_A_117_297#_c_189_n N_VPWR_c_490_n 0.0124092f $X=3.045 $Y=1.41 $X2=0
+ $Y2=0
cc_201 N_A_117_297#_c_190_n N_VPWR_c_490_n 0.0124092f $X=3.515 $Y=1.41 $X2=0
+ $Y2=0
cc_202 N_A_117_297#_c_191_n N_VPWR_c_490_n 0.0124092f $X=3.985 $Y=1.41 $X2=0
+ $Y2=0
cc_203 N_A_117_297#_c_192_n N_VPWR_c_490_n 0.0124092f $X=4.455 $Y=1.41 $X2=0
+ $Y2=0
cc_204 N_A_117_297#_c_193_n N_VPWR_c_490_n 0.0124092f $X=4.925 $Y=1.41 $X2=0
+ $Y2=0
cc_205 N_A_117_297#_c_194_n N_VPWR_c_490_n 0.0124344f $X=5.395 $Y=1.41 $X2=0
+ $Y2=0
cc_206 N_A_117_297#_c_199_n N_VPWR_c_490_n 0.0159357f $X=0.73 $Y=2.3 $X2=0 $Y2=0
cc_207 N_A_117_297#_c_185_n N_A_345_297#_c_614_n 0.0274221f $X=5.26 $Y=1.16
+ $X2=0 $Y2=0
cc_208 N_A_117_297#_c_187_n N_A_345_297#_c_616_n 0.0172483f $X=2.105 $Y=1.41
+ $X2=0 $Y2=0
cc_209 N_A_117_297#_c_188_n N_A_345_297#_c_616_n 0.0170128f $X=2.575 $Y=1.41
+ $X2=0 $Y2=0
cc_210 N_A_117_297#_c_185_n N_A_345_297#_c_616_n 0.0495443f $X=5.26 $Y=1.16
+ $X2=0 $Y2=0
cc_211 N_A_117_297#_c_186_n N_A_345_297#_c_616_n 0.00841423f $X=5.395 $Y=1.202
+ $X2=0 $Y2=0
cc_212 N_A_117_297#_c_189_n N_A_345_297#_c_617_n 0.0170128f $X=3.045 $Y=1.41
+ $X2=0 $Y2=0
cc_213 N_A_117_297#_c_190_n N_A_345_297#_c_617_n 0.0170128f $X=3.515 $Y=1.41
+ $X2=0 $Y2=0
cc_214 N_A_117_297#_c_185_n N_A_345_297#_c_617_n 0.0495054f $X=5.26 $Y=1.16
+ $X2=0 $Y2=0
cc_215 N_A_117_297#_c_186_n N_A_345_297#_c_617_n 0.00868907f $X=5.395 $Y=1.202
+ $X2=0 $Y2=0
cc_216 N_A_117_297#_c_191_n N_A_345_297#_c_618_n 0.0170128f $X=3.985 $Y=1.41
+ $X2=0 $Y2=0
cc_217 N_A_117_297#_c_192_n N_A_345_297#_c_618_n 0.0170128f $X=4.455 $Y=1.41
+ $X2=0 $Y2=0
cc_218 N_A_117_297#_c_185_n N_A_345_297#_c_618_n 0.0495054f $X=5.26 $Y=1.16
+ $X2=0 $Y2=0
cc_219 N_A_117_297#_c_186_n N_A_345_297#_c_618_n 0.00868907f $X=5.395 $Y=1.202
+ $X2=0 $Y2=0
cc_220 N_A_117_297#_c_193_n N_A_345_297#_c_619_n 0.0170128f $X=4.925 $Y=1.41
+ $X2=0 $Y2=0
cc_221 N_A_117_297#_c_194_n N_A_345_297#_c_619_n 0.0169521f $X=5.395 $Y=1.41
+ $X2=0 $Y2=0
cc_222 N_A_117_297#_c_185_n N_A_345_297#_c_619_n 0.0495443f $X=5.26 $Y=1.16
+ $X2=0 $Y2=0
cc_223 N_A_117_297#_c_186_n N_A_345_297#_c_619_n 0.0082085f $X=5.395 $Y=1.202
+ $X2=0 $Y2=0
cc_224 N_A_117_297#_c_185_n N_A_345_297#_c_620_n 0.00128541f $X=5.26 $Y=1.16
+ $X2=0 $Y2=0
cc_225 N_A_117_297#_c_185_n N_A_345_297#_c_621_n 0.0204509f $X=5.26 $Y=1.16
+ $X2=0 $Y2=0
cc_226 N_A_117_297#_c_186_n N_A_345_297#_c_621_n 0.00656533f $X=5.395 $Y=1.202
+ $X2=0 $Y2=0
cc_227 N_A_117_297#_c_185_n N_A_345_297#_c_622_n 0.0204509f $X=5.26 $Y=1.16
+ $X2=0 $Y2=0
cc_228 N_A_117_297#_c_186_n N_A_345_297#_c_622_n 0.00656533f $X=5.395 $Y=1.202
+ $X2=0 $Y2=0
cc_229 N_A_117_297#_c_185_n N_A_345_297#_c_623_n 0.0204509f $X=5.26 $Y=1.16
+ $X2=0 $Y2=0
cc_230 N_A_117_297#_c_186_n N_A_345_297#_c_623_n 0.00656533f $X=5.395 $Y=1.202
+ $X2=0 $Y2=0
cc_231 N_A_117_297#_c_177_n N_X_c_741_n 0.00539651f $X=2.08 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_117_297#_c_178_n N_X_c_741_n 0.00686626f $X=2.55 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_117_297#_c_179_n N_X_c_741_n 5.45498e-19 $X=3.02 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A_117_297#_c_178_n N_X_c_718_n 0.00901745f $X=2.55 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A_117_297#_c_179_n N_X_c_718_n 0.00901745f $X=3.02 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A_117_297#_c_185_n N_X_c_718_n 0.0398926f $X=5.26 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A_117_297#_c_186_n N_X_c_718_n 0.00345541f $X=5.395 $Y=1.202 $X2=0
+ $Y2=0
cc_238 N_A_117_297#_c_177_n N_X_c_719_n 0.00266157f $X=2.08 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A_117_297#_c_178_n N_X_c_719_n 0.00116636f $X=2.55 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A_117_297#_c_185_n N_X_c_719_n 0.0307014f $X=5.26 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A_117_297#_c_186_n N_X_c_719_n 0.00358305f $X=5.395 $Y=1.202 $X2=0
+ $Y2=0
cc_242 N_A_117_297#_c_178_n N_X_c_752_n 5.24597e-19 $X=2.55 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A_117_297#_c_179_n N_X_c_752_n 0.00651696f $X=3.02 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_117_297#_c_180_n N_X_c_752_n 0.00686626f $X=3.49 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A_117_297#_c_181_n N_X_c_752_n 5.45498e-19 $X=3.96 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_117_297#_c_180_n N_X_c_720_n 0.00901745f $X=3.49 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A_117_297#_c_181_n N_X_c_720_n 0.00901745f $X=3.96 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A_117_297#_c_185_n N_X_c_720_n 0.0398926f $X=5.26 $Y=1.16 $X2=0 $Y2=0
cc_249 N_A_117_297#_c_186_n N_X_c_720_n 0.00345541f $X=5.395 $Y=1.202 $X2=0
+ $Y2=0
cc_250 N_A_117_297#_c_180_n N_X_c_760_n 5.24597e-19 $X=3.49 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A_117_297#_c_181_n N_X_c_760_n 0.00651696f $X=3.96 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A_117_297#_c_182_n N_X_c_760_n 0.00686626f $X=4.43 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A_117_297#_c_183_n N_X_c_760_n 5.45498e-19 $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A_117_297#_c_182_n N_X_c_721_n 0.00901745f $X=4.43 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A_117_297#_c_183_n N_X_c_721_n 0.00901745f $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_256 N_A_117_297#_c_185_n N_X_c_721_n 0.0398926f $X=5.26 $Y=1.16 $X2=0 $Y2=0
cc_257 N_A_117_297#_c_186_n N_X_c_721_n 0.00345541f $X=5.395 $Y=1.202 $X2=0
+ $Y2=0
cc_258 N_A_117_297#_c_182_n N_X_c_768_n 5.24597e-19 $X=4.43 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A_117_297#_c_183_n N_X_c_768_n 0.00651696f $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_260 N_A_117_297#_c_184_n N_X_c_722_n 0.0106151f $X=5.42 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A_117_297#_c_185_n N_X_c_722_n 0.0137232f $X=5.26 $Y=1.16 $X2=0 $Y2=0
cc_262 N_A_117_297#_c_184_n N_X_c_772_n 5.32212e-19 $X=5.42 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A_117_297#_c_179_n N_X_c_726_n 0.00116636f $X=3.02 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A_117_297#_c_180_n N_X_c_726_n 0.00116636f $X=3.49 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A_117_297#_c_185_n N_X_c_726_n 0.0307014f $X=5.26 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A_117_297#_c_186_n N_X_c_726_n 0.00358305f $X=5.395 $Y=1.202 $X2=0
+ $Y2=0
cc_267 N_A_117_297#_c_181_n N_X_c_727_n 0.00116636f $X=3.96 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A_117_297#_c_182_n N_X_c_727_n 0.00116636f $X=4.43 $Y=0.995 $X2=0 $Y2=0
cc_269 N_A_117_297#_c_185_n N_X_c_727_n 0.0307014f $X=5.26 $Y=1.16 $X2=0 $Y2=0
cc_270 N_A_117_297#_c_186_n N_X_c_727_n 0.00358305f $X=5.395 $Y=1.202 $X2=0
+ $Y2=0
cc_271 N_A_117_297#_c_183_n N_X_c_728_n 0.00119564f $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A_117_297#_c_185_n N_X_c_728_n 0.030835f $X=5.26 $Y=1.16 $X2=0 $Y2=0
cc_273 N_A_117_297#_c_186_n N_X_c_728_n 0.00486271f $X=5.395 $Y=1.202 $X2=0
+ $Y2=0
cc_274 N_A_117_297#_c_201_n N_VGND_c_940_n 0.0246884f $X=1.04 $Y=0.39 $X2=0
+ $Y2=0
cc_275 N_A_117_297#_c_195_n N_VGND_c_940_n 0.00726615f $X=0.73 $Y=1.62 $X2=0
+ $Y2=0
cc_276 N_A_117_297#_c_177_n N_VGND_c_941_n 0.00373705f $X=2.08 $Y=0.995 $X2=0
+ $Y2=0
cc_277 N_A_117_297#_c_201_n N_VGND_c_941_n 0.0446925f $X=1.04 $Y=0.39 $X2=0
+ $Y2=0
cc_278 N_A_117_297#_c_185_n N_VGND_c_941_n 0.0435327f $X=5.26 $Y=1.16 $X2=0
+ $Y2=0
cc_279 N_A_117_297#_c_178_n N_VGND_c_942_n 0.00379224f $X=2.55 $Y=0.995 $X2=0
+ $Y2=0
cc_280 N_A_117_297#_c_179_n N_VGND_c_942_n 0.00276126f $X=3.02 $Y=0.995 $X2=0
+ $Y2=0
cc_281 N_A_117_297#_c_180_n N_VGND_c_943_n 0.00379224f $X=3.49 $Y=0.995 $X2=0
+ $Y2=0
cc_282 N_A_117_297#_c_181_n N_VGND_c_943_n 0.00276126f $X=3.96 $Y=0.995 $X2=0
+ $Y2=0
cc_283 N_A_117_297#_c_182_n N_VGND_c_944_n 0.00379224f $X=4.43 $Y=0.995 $X2=0
+ $Y2=0
cc_284 N_A_117_297#_c_183_n N_VGND_c_944_n 0.00276126f $X=4.9 $Y=0.995 $X2=0
+ $Y2=0
cc_285 N_A_117_297#_c_184_n N_VGND_c_945_n 0.00268723f $X=5.42 $Y=0.995 $X2=0
+ $Y2=0
cc_286 N_A_117_297#_c_177_n N_VGND_c_953_n 0.00541359f $X=2.08 $Y=0.995 $X2=0
+ $Y2=0
cc_287 N_A_117_297#_c_178_n N_VGND_c_953_n 0.00423334f $X=2.55 $Y=0.995 $X2=0
+ $Y2=0
cc_288 N_A_117_297#_c_179_n N_VGND_c_955_n 0.00423334f $X=3.02 $Y=0.995 $X2=0
+ $Y2=0
cc_289 N_A_117_297#_c_180_n N_VGND_c_955_n 0.00423334f $X=3.49 $Y=0.995 $X2=0
+ $Y2=0
cc_290 N_A_117_297#_c_181_n N_VGND_c_957_n 0.00423334f $X=3.96 $Y=0.995 $X2=0
+ $Y2=0
cc_291 N_A_117_297#_c_182_n N_VGND_c_957_n 0.00423334f $X=4.43 $Y=0.995 $X2=0
+ $Y2=0
cc_292 N_A_117_297#_c_183_n N_VGND_c_959_n 0.00423334f $X=4.9 $Y=0.995 $X2=0
+ $Y2=0
cc_293 N_A_117_297#_c_184_n N_VGND_c_959_n 0.00437852f $X=5.42 $Y=0.995 $X2=0
+ $Y2=0
cc_294 N_A_117_297#_c_201_n N_VGND_c_967_n 0.0210564f $X=1.04 $Y=0.39 $X2=0
+ $Y2=0
cc_295 N_A_117_297#_M1018_s N_VGND_c_970_n 0.0025535f $X=0.885 $Y=0.235 $X2=0
+ $Y2=0
cc_296 N_A_117_297#_c_177_n N_VGND_c_970_n 0.0103342f $X=2.08 $Y=0.995 $X2=0
+ $Y2=0
cc_297 N_A_117_297#_c_178_n N_VGND_c_970_n 0.006093f $X=2.55 $Y=0.995 $X2=0
+ $Y2=0
cc_298 N_A_117_297#_c_179_n N_VGND_c_970_n 0.00597024f $X=3.02 $Y=0.995 $X2=0
+ $Y2=0
cc_299 N_A_117_297#_c_180_n N_VGND_c_970_n 0.006093f $X=3.49 $Y=0.995 $X2=0
+ $Y2=0
cc_300 N_A_117_297#_c_181_n N_VGND_c_970_n 0.00597024f $X=3.96 $Y=0.995 $X2=0
+ $Y2=0
cc_301 N_A_117_297#_c_182_n N_VGND_c_970_n 0.006093f $X=4.43 $Y=0.995 $X2=0
+ $Y2=0
cc_302 N_A_117_297#_c_183_n N_VGND_c_970_n 0.00608558f $X=4.9 $Y=0.995 $X2=0
+ $Y2=0
cc_303 N_A_117_297#_c_184_n N_VGND_c_970_n 0.00615622f $X=5.42 $Y=0.995 $X2=0
+ $Y2=0
cc_304 N_A_117_297#_c_201_n N_VGND_c_970_n 0.0134685f $X=1.04 $Y=0.39 $X2=0
+ $Y2=0
cc_305 N_SLEEP_c_360_n N_VPWR_c_508_n 0.00429453f $X=5.865 $Y=1.41 $X2=0 $Y2=0
cc_306 N_SLEEP_c_361_n N_VPWR_c_508_n 0.00429453f $X=6.335 $Y=1.41 $X2=0 $Y2=0
cc_307 N_SLEEP_c_362_n N_VPWR_c_508_n 0.00429453f $X=6.805 $Y=1.41 $X2=0 $Y2=0
cc_308 N_SLEEP_c_363_n N_VPWR_c_508_n 0.00429453f $X=7.275 $Y=1.41 $X2=0 $Y2=0
cc_309 N_SLEEP_c_364_n N_VPWR_c_508_n 0.00429453f $X=7.745 $Y=1.41 $X2=0 $Y2=0
cc_310 N_SLEEP_c_365_n N_VPWR_c_508_n 0.00429453f $X=8.215 $Y=1.41 $X2=0 $Y2=0
cc_311 N_SLEEP_c_366_n N_VPWR_c_508_n 0.00429453f $X=8.685 $Y=1.41 $X2=0 $Y2=0
cc_312 N_SLEEP_c_367_n N_VPWR_c_508_n 0.00429453f $X=9.155 $Y=1.41 $X2=0 $Y2=0
cc_313 N_SLEEP_c_360_n N_VPWR_c_490_n 0.00609021f $X=5.865 $Y=1.41 $X2=0 $Y2=0
cc_314 N_SLEEP_c_361_n N_VPWR_c_490_n 0.00606499f $X=6.335 $Y=1.41 $X2=0 $Y2=0
cc_315 N_SLEEP_c_362_n N_VPWR_c_490_n 0.00606499f $X=6.805 $Y=1.41 $X2=0 $Y2=0
cc_316 N_SLEEP_c_363_n N_VPWR_c_490_n 0.00606499f $X=7.275 $Y=1.41 $X2=0 $Y2=0
cc_317 N_SLEEP_c_364_n N_VPWR_c_490_n 0.00606499f $X=7.745 $Y=1.41 $X2=0 $Y2=0
cc_318 N_SLEEP_c_365_n N_VPWR_c_490_n 0.00606499f $X=8.215 $Y=1.41 $X2=0 $Y2=0
cc_319 N_SLEEP_c_366_n N_VPWR_c_490_n 0.00606499f $X=8.685 $Y=1.41 $X2=0 $Y2=0
cc_320 N_SLEEP_c_367_n N_VPWR_c_490_n 0.00698562f $X=9.155 $Y=1.41 $X2=0 $Y2=0
cc_321 N_SLEEP_c_360_n N_A_345_297#_c_620_n 2.98195e-19 $X=5.865 $Y=1.41 $X2=0
+ $Y2=0
cc_322 N_SLEEP_c_360_n N_A_345_297#_c_649_n 0.0143578f $X=5.865 $Y=1.41 $X2=0
+ $Y2=0
cc_323 N_SLEEP_c_361_n N_A_345_297#_c_649_n 0.0143578f $X=6.335 $Y=1.41 $X2=0
+ $Y2=0
cc_324 N_SLEEP_c_362_n N_A_345_297#_c_651_n 0.0143578f $X=6.805 $Y=1.41 $X2=0
+ $Y2=0
cc_325 N_SLEEP_c_363_n N_A_345_297#_c_651_n 0.0143578f $X=7.275 $Y=1.41 $X2=0
+ $Y2=0
cc_326 N_SLEEP_c_364_n N_A_345_297#_c_653_n 0.0143578f $X=7.745 $Y=1.41 $X2=0
+ $Y2=0
cc_327 N_SLEEP_c_365_n N_A_345_297#_c_653_n 0.0143578f $X=8.215 $Y=1.41 $X2=0
+ $Y2=0
cc_328 N_SLEEP_c_366_n N_A_345_297#_c_655_n 0.0143578f $X=8.685 $Y=1.41 $X2=0
+ $Y2=0
cc_329 N_SLEEP_c_367_n N_A_345_297#_c_655_n 0.0143578f $X=9.155 $Y=1.41 $X2=0
+ $Y2=0
cc_330 N_SLEEP_c_351_n N_X_c_722_n 0.00940242f $X=5.84 $Y=0.995 $X2=0 $Y2=0
cc_331 N_SLEEP_c_371_n N_X_c_722_n 0.00651491f $X=8.645 $Y=1.16 $X2=0 $Y2=0
cc_332 N_SLEEP_c_351_n N_X_c_772_n 0.00644736f $X=5.84 $Y=0.995 $X2=0 $Y2=0
cc_333 N_SLEEP_c_352_n N_X_c_772_n 0.00686626f $X=6.31 $Y=0.995 $X2=0 $Y2=0
cc_334 N_SLEEP_c_353_n N_X_c_772_n 5.45498e-19 $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_335 N_SLEEP_c_361_n N_X_c_734_n 0.015669f $X=6.335 $Y=1.41 $X2=0 $Y2=0
cc_336 N_SLEEP_c_362_n N_X_c_734_n 0.0157513f $X=6.805 $Y=1.41 $X2=0 $Y2=0
cc_337 N_SLEEP_c_371_n N_X_c_734_n 0.0485189f $X=8.645 $Y=1.16 $X2=0 $Y2=0
cc_338 N_SLEEP_c_359_n N_X_c_734_n 0.00875187f $X=9.155 $Y=1.202 $X2=0 $Y2=0
cc_339 N_SLEEP_c_360_n N_X_c_735_n 6.32035e-19 $X=5.865 $Y=1.41 $X2=0 $Y2=0
cc_340 N_SLEEP_c_371_n N_X_c_735_n 0.020385f $X=8.645 $Y=1.16 $X2=0 $Y2=0
cc_341 N_SLEEP_c_359_n N_X_c_735_n 0.00663436f $X=9.155 $Y=1.202 $X2=0 $Y2=0
cc_342 N_SLEEP_c_352_n N_X_c_723_n 0.00901745f $X=6.31 $Y=0.995 $X2=0 $Y2=0
cc_343 N_SLEEP_c_353_n N_X_c_723_n 0.00901745f $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_344 N_SLEEP_c_371_n N_X_c_723_n 0.0397461f $X=8.645 $Y=1.16 $X2=0 $Y2=0
cc_345 N_SLEEP_c_359_n N_X_c_723_n 0.00345541f $X=9.155 $Y=1.202 $X2=0 $Y2=0
cc_346 N_SLEEP_c_352_n N_X_c_800_n 5.24597e-19 $X=6.31 $Y=0.995 $X2=0 $Y2=0
cc_347 N_SLEEP_c_353_n N_X_c_800_n 0.00651696f $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_348 N_SLEEP_c_354_n N_X_c_800_n 0.00686626f $X=7.25 $Y=0.995 $X2=0 $Y2=0
cc_349 N_SLEEP_c_355_n N_X_c_800_n 5.45498e-19 $X=7.72 $Y=0.995 $X2=0 $Y2=0
cc_350 N_SLEEP_c_363_n N_X_c_736_n 0.0157513f $X=7.275 $Y=1.41 $X2=0 $Y2=0
cc_351 N_SLEEP_c_364_n N_X_c_736_n 0.0157513f $X=7.745 $Y=1.41 $X2=0 $Y2=0
cc_352 N_SLEEP_c_371_n N_X_c_736_n 0.0485189f $X=8.645 $Y=1.16 $X2=0 $Y2=0
cc_353 N_SLEEP_c_359_n N_X_c_736_n 0.00875187f $X=9.155 $Y=1.202 $X2=0 $Y2=0
cc_354 N_SLEEP_c_354_n N_X_c_724_n 0.00901745f $X=7.25 $Y=0.995 $X2=0 $Y2=0
cc_355 N_SLEEP_c_355_n N_X_c_724_n 0.00901745f $X=7.72 $Y=0.995 $X2=0 $Y2=0
cc_356 N_SLEEP_c_371_n N_X_c_724_n 0.0397461f $X=8.645 $Y=1.16 $X2=0 $Y2=0
cc_357 N_SLEEP_c_359_n N_X_c_724_n 0.00345541f $X=9.155 $Y=1.202 $X2=0 $Y2=0
cc_358 N_SLEEP_c_354_n N_X_c_812_n 5.24597e-19 $X=7.25 $Y=0.995 $X2=0 $Y2=0
cc_359 N_SLEEP_c_355_n N_X_c_812_n 0.00651696f $X=7.72 $Y=0.995 $X2=0 $Y2=0
cc_360 N_SLEEP_c_356_n N_X_c_812_n 0.00686352f $X=8.19 $Y=0.995 $X2=0 $Y2=0
cc_361 N_SLEEP_c_357_n N_X_c_812_n 5.45311e-19 $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_362 N_SLEEP_c_365_n N_X_c_737_n 0.0157513f $X=8.215 $Y=1.41 $X2=0 $Y2=0
cc_363 N_SLEEP_c_366_n N_X_c_737_n 0.0157513f $X=8.685 $Y=1.41 $X2=0 $Y2=0
cc_364 N_SLEEP_c_371_n N_X_c_737_n 0.0485189f $X=8.645 $Y=1.16 $X2=0 $Y2=0
cc_365 N_SLEEP_c_359_n N_X_c_737_n 0.00875187f $X=9.155 $Y=1.202 $X2=0 $Y2=0
cc_366 N_SLEEP_c_356_n N_X_c_725_n 0.00901745f $X=8.19 $Y=0.995 $X2=0 $Y2=0
cc_367 N_SLEEP_c_357_n N_X_c_725_n 0.00901745f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_368 N_SLEEP_c_371_n N_X_c_725_n 0.0397461f $X=8.645 $Y=1.16 $X2=0 $Y2=0
cc_369 N_SLEEP_c_359_n N_X_c_725_n 0.00345541f $X=9.155 $Y=1.202 $X2=0 $Y2=0
cc_370 N_SLEEP_c_351_n N_X_c_729_n 0.00116636f $X=5.84 $Y=0.995 $X2=0 $Y2=0
cc_371 N_SLEEP_c_352_n N_X_c_729_n 0.00116636f $X=6.31 $Y=0.995 $X2=0 $Y2=0
cc_372 N_SLEEP_c_371_n N_X_c_729_n 0.0306016f $X=8.645 $Y=1.16 $X2=0 $Y2=0
cc_373 N_SLEEP_c_359_n N_X_c_729_n 0.00358305f $X=9.155 $Y=1.202 $X2=0 $Y2=0
cc_374 N_SLEEP_c_353_n N_X_c_730_n 0.00116636f $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_375 N_SLEEP_c_354_n N_X_c_730_n 0.00116636f $X=7.25 $Y=0.995 $X2=0 $Y2=0
cc_376 N_SLEEP_c_371_n N_X_c_730_n 0.0306016f $X=8.645 $Y=1.16 $X2=0 $Y2=0
cc_377 N_SLEEP_c_359_n N_X_c_730_n 0.00358305f $X=9.155 $Y=1.202 $X2=0 $Y2=0
cc_378 N_SLEEP_c_371_n N_X_c_738_n 0.020385f $X=8.645 $Y=1.16 $X2=0 $Y2=0
cc_379 N_SLEEP_c_359_n N_X_c_738_n 0.00663436f $X=9.155 $Y=1.202 $X2=0 $Y2=0
cc_380 N_SLEEP_c_355_n N_X_c_731_n 0.00116636f $X=7.72 $Y=0.995 $X2=0 $Y2=0
cc_381 N_SLEEP_c_356_n N_X_c_731_n 0.00116636f $X=8.19 $Y=0.995 $X2=0 $Y2=0
cc_382 N_SLEEP_c_371_n N_X_c_731_n 0.0306016f $X=8.645 $Y=1.16 $X2=0 $Y2=0
cc_383 N_SLEEP_c_359_n N_X_c_731_n 0.00358305f $X=9.155 $Y=1.202 $X2=0 $Y2=0
cc_384 N_SLEEP_c_371_n N_X_c_739_n 0.020385f $X=8.645 $Y=1.16 $X2=0 $Y2=0
cc_385 N_SLEEP_c_359_n N_X_c_739_n 0.00663436f $X=9.155 $Y=1.202 $X2=0 $Y2=0
cc_386 N_SLEEP_c_356_n N_X_c_732_n 5.25778e-19 $X=8.19 $Y=0.995 $X2=0 $Y2=0
cc_387 N_SLEEP_c_357_n N_X_c_732_n 0.00777632f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_388 N_SLEEP_c_358_n N_X_c_732_n 0.0102332f $X=9.18 $Y=0.995 $X2=0 $Y2=0
cc_389 N_SLEEP_c_371_n N_X_c_732_n 0.0140822f $X=8.645 $Y=1.16 $X2=0 $Y2=0
cc_390 N_SLEEP_c_359_n N_X_c_732_n 0.0056758f $X=9.155 $Y=1.202 $X2=0 $Y2=0
cc_391 N_SLEEP_c_357_n X 8.93496e-19 $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_392 N_SLEEP_c_367_n X 0.0177539f $X=9.155 $Y=1.41 $X2=0 $Y2=0
cc_393 N_SLEEP_c_358_n X 0.00401352f $X=9.18 $Y=0.995 $X2=0 $Y2=0
cc_394 N_SLEEP_c_371_n X 0.0232619f $X=8.645 $Y=1.16 $X2=0 $Y2=0
cc_395 N_SLEEP_c_359_n X 0.0357067f $X=9.155 $Y=1.202 $X2=0 $Y2=0
cc_396 N_SLEEP_c_351_n N_VGND_c_945_n 0.00268723f $X=5.84 $Y=0.995 $X2=0 $Y2=0
cc_397 N_SLEEP_c_352_n N_VGND_c_946_n 0.00379224f $X=6.31 $Y=0.995 $X2=0 $Y2=0
cc_398 N_SLEEP_c_353_n N_VGND_c_946_n 0.00276126f $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_399 N_SLEEP_c_354_n N_VGND_c_947_n 0.00379224f $X=7.25 $Y=0.995 $X2=0 $Y2=0
cc_400 N_SLEEP_c_355_n N_VGND_c_947_n 0.00276126f $X=7.72 $Y=0.995 $X2=0 $Y2=0
cc_401 N_SLEEP_c_356_n N_VGND_c_948_n 0.00379224f $X=8.19 $Y=0.995 $X2=0 $Y2=0
cc_402 N_SLEEP_c_357_n N_VGND_c_948_n 0.00276126f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_403 N_SLEEP_c_358_n N_VGND_c_950_n 0.00451776f $X=9.18 $Y=0.995 $X2=0 $Y2=0
cc_404 N_SLEEP_c_351_n N_VGND_c_961_n 0.00423334f $X=5.84 $Y=0.995 $X2=0 $Y2=0
cc_405 N_SLEEP_c_352_n N_VGND_c_961_n 0.00423334f $X=6.31 $Y=0.995 $X2=0 $Y2=0
cc_406 N_SLEEP_c_353_n N_VGND_c_963_n 0.00423334f $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_407 N_SLEEP_c_354_n N_VGND_c_963_n 0.00423334f $X=7.25 $Y=0.995 $X2=0 $Y2=0
cc_408 N_SLEEP_c_355_n N_VGND_c_965_n 0.00423334f $X=7.72 $Y=0.995 $X2=0 $Y2=0
cc_409 N_SLEEP_c_356_n N_VGND_c_965_n 0.00423334f $X=8.19 $Y=0.995 $X2=0 $Y2=0
cc_410 N_SLEEP_c_357_n N_VGND_c_968_n 0.00421816f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_411 N_SLEEP_c_358_n N_VGND_c_968_n 0.00437716f $X=9.18 $Y=0.995 $X2=0 $Y2=0
cc_412 N_SLEEP_c_351_n N_VGND_c_970_n 0.00587047f $X=5.84 $Y=0.995 $X2=0 $Y2=0
cc_413 N_SLEEP_c_352_n N_VGND_c_970_n 0.006093f $X=6.31 $Y=0.995 $X2=0 $Y2=0
cc_414 N_SLEEP_c_353_n N_VGND_c_970_n 0.00597024f $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_415 N_SLEEP_c_354_n N_VGND_c_970_n 0.006093f $X=7.25 $Y=0.995 $X2=0 $Y2=0
cc_416 N_SLEEP_c_355_n N_VGND_c_970_n 0.00597024f $X=7.72 $Y=0.995 $X2=0 $Y2=0
cc_417 N_SLEEP_c_356_n N_VGND_c_970_n 0.006093f $X=8.19 $Y=0.995 $X2=0 $Y2=0
cc_418 N_SLEEP_c_357_n N_VGND_c_970_n 0.00609466f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_419 N_SLEEP_c_358_n N_VGND_c_970_n 0.00709025f $X=9.18 $Y=0.995 $X2=0 $Y2=0
cc_420 N_VPWR_c_490_n N_A_345_297#_M1000_s 0.00303344f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_421 N_VPWR_c_490_n N_A_345_297#_M1002_s 0.00370124f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_490_n N_A_345_297#_M1005_s 0.00370124f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_423 N_VPWR_c_490_n N_A_345_297#_M1017_s 0.00370124f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_490_n N_A_345_297#_M1031_s 0.00297222f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_490_n N_A_345_297#_M1007_d 0.00231264f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_490_n N_A_345_297#_M1021_d 0.00231264f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_490_n N_A_345_297#_M1028_d 0.00231264f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_490_n N_A_345_297#_M1035_d 0.00260432f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_493_n N_A_345_297#_c_614_n 0.0156204f $X=1.25 $Y=1.64 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_493_n N_A_345_297#_c_615_n 0.0558737f $X=1.25 $Y=1.64 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_500_n N_A_345_297#_c_615_n 0.0211751f $X=2.215 $Y=2.72 $X2=0
+ $Y2=0
cc_432 N_VPWR_c_490_n N_A_345_297#_c_615_n 0.0122467f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_433 N_VPWR_M1000_d N_A_345_297#_c_616_n 0.00188315f $X=2.195 $Y=1.485 $X2=0
+ $Y2=0
cc_434 N_VPWR_c_494_n N_A_345_297#_c_616_n 0.0145257f $X=2.34 $Y=2 $X2=0 $Y2=0
cc_435 N_VPWR_c_502_n N_A_345_297#_c_672_n 0.0149311f $X=3.155 $Y=2.72 $X2=0
+ $Y2=0
cc_436 N_VPWR_c_490_n N_A_345_297#_c_672_n 0.00955092f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_437 N_VPWR_M1004_d N_A_345_297#_c_617_n 0.00188315f $X=3.135 $Y=1.485 $X2=0
+ $Y2=0
cc_438 N_VPWR_c_495_n N_A_345_297#_c_617_n 0.0145257f $X=3.28 $Y=2 $X2=0 $Y2=0
cc_439 N_VPWR_c_504_n N_A_345_297#_c_676_n 0.0149311f $X=4.095 $Y=2.72 $X2=0
+ $Y2=0
cc_440 N_VPWR_c_490_n N_A_345_297#_c_676_n 0.00955092f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_441 N_VPWR_M1015_d N_A_345_297#_c_618_n 0.00188315f $X=4.075 $Y=1.485 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_496_n N_A_345_297#_c_618_n 0.0145257f $X=4.22 $Y=2 $X2=0 $Y2=0
cc_443 N_VPWR_c_506_n N_A_345_297#_c_680_n 0.0149311f $X=5.035 $Y=2.72 $X2=0
+ $Y2=0
cc_444 N_VPWR_c_490_n N_A_345_297#_c_680_n 0.00955092f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_445 N_VPWR_M1023_d N_A_345_297#_c_619_n 0.00188315f $X=5.015 $Y=1.485 $X2=0
+ $Y2=0
cc_446 N_VPWR_c_497_n N_A_345_297#_c_619_n 0.0145257f $X=5.16 $Y=2 $X2=0 $Y2=0
cc_447 N_VPWR_c_508_n N_A_345_297#_c_684_n 0.015002f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_448 N_VPWR_c_490_n N_A_345_297#_c_684_n 0.00962794f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_449 N_VPWR_c_508_n N_A_345_297#_c_649_n 0.0386815f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_450 N_VPWR_c_490_n N_A_345_297#_c_649_n 0.0239144f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_451 N_VPWR_c_508_n N_A_345_297#_c_651_n 0.0386815f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_452 N_VPWR_c_490_n N_A_345_297#_c_651_n 0.0239144f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_453 N_VPWR_c_508_n N_A_345_297#_c_653_n 0.0386815f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_454 N_VPWR_c_490_n N_A_345_297#_c_653_n 0.0239144f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_455 N_VPWR_c_508_n N_A_345_297#_c_655_n 0.0549726f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_456 N_VPWR_c_490_n N_A_345_297#_c_655_n 0.0335424f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_457 N_VPWR_c_508_n N_A_345_297#_c_694_n 0.015002f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_458 N_VPWR_c_490_n N_A_345_297#_c_694_n 0.00962794f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_459 N_VPWR_c_508_n N_A_345_297#_c_696_n 0.015002f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_460 N_VPWR_c_490_n N_A_345_297#_c_696_n 0.00962794f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_461 N_VPWR_c_508_n N_A_345_297#_c_698_n 0.015002f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_462 N_VPWR_c_490_n N_A_345_297#_c_698_n 0.00962794f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_490_n N_X_M1003_s 0.00232895f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_464 N_VPWR_c_490_n N_X_M1016_s 0.00232895f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_465 N_VPWR_c_490_n N_X_M1025_s 0.00232895f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_466 N_VPWR_c_490_n N_X_M1034_s 0.00232895f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_467 N_A_345_297#_c_649_n N_X_M1003_s 0.00352392f $X=6.445 $Y=2.38 $X2=0 $Y2=0
cc_468 N_A_345_297#_c_651_n N_X_M1016_s 0.00352392f $X=7.385 $Y=2.38 $X2=0 $Y2=0
cc_469 N_A_345_297#_c_653_n N_X_M1025_s 0.00352392f $X=8.325 $Y=2.38 $X2=0 $Y2=0
cc_470 N_A_345_297#_c_655_n N_X_M1034_s 0.00352392f $X=9.265 $Y=2.38 $X2=0 $Y2=0
cc_471 N_A_345_297#_c_620_n N_X_c_722_n 0.0088033f $X=5.63 $Y=1.665 $X2=0 $Y2=0
cc_472 N_A_345_297#_c_649_n N_X_c_859_n 0.0134104f $X=6.445 $Y=2.38 $X2=0 $Y2=0
cc_473 N_A_345_297#_M1007_d N_X_c_734_n 0.00187091f $X=6.425 $Y=1.485 $X2=0
+ $Y2=0
cc_474 N_A_345_297#_c_707_p N_X_c_734_n 0.0143191f $X=6.57 $Y=1.96 $X2=0 $Y2=0
cc_475 N_A_345_297#_c_620_n N_X_c_735_n 0.00226124f $X=5.63 $Y=1.665 $X2=0 $Y2=0
cc_476 N_A_345_297#_c_651_n N_X_c_863_n 0.0134104f $X=7.385 $Y=2.38 $X2=0 $Y2=0
cc_477 N_A_345_297#_M1021_d N_X_c_736_n 0.00187091f $X=7.365 $Y=1.485 $X2=0
+ $Y2=0
cc_478 N_A_345_297#_c_711_p N_X_c_736_n 0.0143191f $X=7.51 $Y=1.96 $X2=0 $Y2=0
cc_479 N_A_345_297#_c_653_n N_X_c_866_n 0.0134104f $X=8.325 $Y=2.38 $X2=0 $Y2=0
cc_480 N_A_345_297#_M1028_d N_X_c_737_n 0.00187091f $X=8.305 $Y=1.485 $X2=0
+ $Y2=0
cc_481 N_A_345_297#_c_714_p N_X_c_737_n 0.0143191f $X=8.45 $Y=1.96 $X2=0 $Y2=0
cc_482 N_A_345_297#_c_655_n N_X_c_869_n 0.0134104f $X=9.265 $Y=2.38 $X2=0 $Y2=0
cc_483 N_A_345_297#_M1035_d X 0.0035037f $X=9.245 $Y=1.485 $X2=0 $Y2=0
cc_484 N_A_345_297#_c_717_p X 0.0191143f $X=9.39 $Y=1.96 $X2=0 $Y2=0
cc_485 N_X_c_718_n N_VGND_M1008_s 0.00251047f $X=3.065 $Y=0.815 $X2=0 $Y2=0
cc_486 N_X_c_720_n N_VGND_M1019_s 0.00251047f $X=4.005 $Y=0.815 $X2=0 $Y2=0
cc_487 N_X_c_721_n N_VGND_M1026_s 0.00251047f $X=4.945 $Y=0.815 $X2=0 $Y2=0
cc_488 N_X_c_722_n N_VGND_M1032_s 0.00162089f $X=5.885 $Y=0.815 $X2=0 $Y2=0
cc_489 N_X_c_723_n N_VGND_M1010_s 0.00251047f $X=6.825 $Y=0.815 $X2=0 $Y2=0
cc_490 N_X_c_724_n N_VGND_M1013_s 0.00251047f $X=7.765 $Y=0.815 $X2=0 $Y2=0
cc_491 N_X_c_725_n N_VGND_M1024_s 0.00251047f $X=8.705 $Y=0.815 $X2=0 $Y2=0
cc_492 N_X_c_732_n N_VGND_M1033_s 0.00290026f $X=8.92 $Y=0.39 $X2=0 $Y2=0
cc_493 N_X_c_719_n N_VGND_c_941_n 0.00843013f $X=2.505 $Y=0.815 $X2=0 $Y2=0
cc_494 N_X_c_741_n N_VGND_c_942_n 0.0183628f $X=2.34 $Y=0.39 $X2=0 $Y2=0
cc_495 N_X_c_718_n N_VGND_c_942_n 0.0127273f $X=3.065 $Y=0.815 $X2=0 $Y2=0
cc_496 N_X_c_752_n N_VGND_c_943_n 0.0183628f $X=3.28 $Y=0.39 $X2=0 $Y2=0
cc_497 N_X_c_720_n N_VGND_c_943_n 0.0127273f $X=4.005 $Y=0.815 $X2=0 $Y2=0
cc_498 N_X_c_760_n N_VGND_c_944_n 0.0183628f $X=4.22 $Y=0.39 $X2=0 $Y2=0
cc_499 N_X_c_721_n N_VGND_c_944_n 0.0127273f $X=4.945 $Y=0.815 $X2=0 $Y2=0
cc_500 N_X_c_722_n N_VGND_c_945_n 0.0122559f $X=5.885 $Y=0.815 $X2=0 $Y2=0
cc_501 N_X_c_772_n N_VGND_c_946_n 0.0183628f $X=6.1 $Y=0.39 $X2=0 $Y2=0
cc_502 N_X_c_723_n N_VGND_c_946_n 0.0127273f $X=6.825 $Y=0.815 $X2=0 $Y2=0
cc_503 N_X_c_800_n N_VGND_c_947_n 0.0183628f $X=7.04 $Y=0.39 $X2=0 $Y2=0
cc_504 N_X_c_724_n N_VGND_c_947_n 0.0127273f $X=7.765 $Y=0.815 $X2=0 $Y2=0
cc_505 N_X_c_812_n N_VGND_c_948_n 0.0183628f $X=7.98 $Y=0.39 $X2=0 $Y2=0
cc_506 N_X_c_725_n N_VGND_c_948_n 0.0127273f $X=8.705 $Y=0.815 $X2=0 $Y2=0
cc_507 N_X_c_732_n N_VGND_c_950_n 0.0220486f $X=8.92 $Y=0.39 $X2=0 $Y2=0
cc_508 N_X_c_741_n N_VGND_c_953_n 0.0223596f $X=2.34 $Y=0.39 $X2=0 $Y2=0
cc_509 N_X_c_718_n N_VGND_c_953_n 0.00266636f $X=3.065 $Y=0.815 $X2=0 $Y2=0
cc_510 N_X_c_718_n N_VGND_c_955_n 0.00198695f $X=3.065 $Y=0.815 $X2=0 $Y2=0
cc_511 N_X_c_752_n N_VGND_c_955_n 0.0223596f $X=3.28 $Y=0.39 $X2=0 $Y2=0
cc_512 N_X_c_720_n N_VGND_c_955_n 0.00266636f $X=4.005 $Y=0.815 $X2=0 $Y2=0
cc_513 N_X_c_720_n N_VGND_c_957_n 0.00198695f $X=4.005 $Y=0.815 $X2=0 $Y2=0
cc_514 N_X_c_760_n N_VGND_c_957_n 0.0223596f $X=4.22 $Y=0.39 $X2=0 $Y2=0
cc_515 N_X_c_721_n N_VGND_c_957_n 0.00266636f $X=4.945 $Y=0.815 $X2=0 $Y2=0
cc_516 N_X_c_721_n N_VGND_c_959_n 0.00198695f $X=4.945 $Y=0.815 $X2=0 $Y2=0
cc_517 N_X_c_768_n N_VGND_c_959_n 0.0231806f $X=5.16 $Y=0.39 $X2=0 $Y2=0
cc_518 N_X_c_722_n N_VGND_c_959_n 0.00254521f $X=5.885 $Y=0.815 $X2=0 $Y2=0
cc_519 N_X_c_722_n N_VGND_c_961_n 0.00198695f $X=5.885 $Y=0.815 $X2=0 $Y2=0
cc_520 N_X_c_772_n N_VGND_c_961_n 0.0223596f $X=6.1 $Y=0.39 $X2=0 $Y2=0
cc_521 N_X_c_723_n N_VGND_c_961_n 0.00266636f $X=6.825 $Y=0.815 $X2=0 $Y2=0
cc_522 N_X_c_723_n N_VGND_c_963_n 0.00198695f $X=6.825 $Y=0.815 $X2=0 $Y2=0
cc_523 N_X_c_800_n N_VGND_c_963_n 0.0223596f $X=7.04 $Y=0.39 $X2=0 $Y2=0
cc_524 N_X_c_724_n N_VGND_c_963_n 0.00266636f $X=7.765 $Y=0.815 $X2=0 $Y2=0
cc_525 N_X_c_724_n N_VGND_c_965_n 0.00198695f $X=7.765 $Y=0.815 $X2=0 $Y2=0
cc_526 N_X_c_812_n N_VGND_c_965_n 0.0223596f $X=7.98 $Y=0.39 $X2=0 $Y2=0
cc_527 N_X_c_725_n N_VGND_c_965_n 0.00266636f $X=8.705 $Y=0.815 $X2=0 $Y2=0
cc_528 N_X_c_725_n N_VGND_c_968_n 0.00198695f $X=8.705 $Y=0.815 $X2=0 $Y2=0
cc_529 N_X_c_732_n N_VGND_c_968_n 0.0260268f $X=8.92 $Y=0.39 $X2=0 $Y2=0
cc_530 N_X_M1006_d N_VGND_c_970_n 0.0025535f $X=2.155 $Y=0.235 $X2=0 $Y2=0
cc_531 N_X_M1011_d N_VGND_c_970_n 0.0025535f $X=3.095 $Y=0.235 $X2=0 $Y2=0
cc_532 N_X_M1020_d N_VGND_c_970_n 0.0025535f $X=4.035 $Y=0.235 $X2=0 $Y2=0
cc_533 N_X_M1029_d N_VGND_c_970_n 0.00304143f $X=4.975 $Y=0.235 $X2=0 $Y2=0
cc_534 N_X_M1009_d N_VGND_c_970_n 0.0025535f $X=5.915 $Y=0.235 $X2=0 $Y2=0
cc_535 N_X_M1012_d N_VGND_c_970_n 0.0025535f $X=6.855 $Y=0.235 $X2=0 $Y2=0
cc_536 N_X_M1022_d N_VGND_c_970_n 0.0025535f $X=7.795 $Y=0.235 $X2=0 $Y2=0
cc_537 N_X_M1030_d N_VGND_c_970_n 0.00304917f $X=8.735 $Y=0.235 $X2=0 $Y2=0
cc_538 N_X_c_741_n N_VGND_c_970_n 0.0141302f $X=2.34 $Y=0.39 $X2=0 $Y2=0
cc_539 N_X_c_718_n N_VGND_c_970_n 0.00972452f $X=3.065 $Y=0.815 $X2=0 $Y2=0
cc_540 N_X_c_752_n N_VGND_c_970_n 0.0141302f $X=3.28 $Y=0.39 $X2=0 $Y2=0
cc_541 N_X_c_720_n N_VGND_c_970_n 0.00972452f $X=4.005 $Y=0.815 $X2=0 $Y2=0
cc_542 N_X_c_760_n N_VGND_c_970_n 0.0141302f $X=4.22 $Y=0.39 $X2=0 $Y2=0
cc_543 N_X_c_721_n N_VGND_c_970_n 0.00972452f $X=4.945 $Y=0.815 $X2=0 $Y2=0
cc_544 N_X_c_768_n N_VGND_c_970_n 0.0143352f $X=5.16 $Y=0.39 $X2=0 $Y2=0
cc_545 N_X_c_722_n N_VGND_c_970_n 0.0094839f $X=5.885 $Y=0.815 $X2=0 $Y2=0
cc_546 N_X_c_772_n N_VGND_c_970_n 0.0141302f $X=6.1 $Y=0.39 $X2=0 $Y2=0
cc_547 N_X_c_723_n N_VGND_c_970_n 0.00972452f $X=6.825 $Y=0.815 $X2=0 $Y2=0
cc_548 N_X_c_800_n N_VGND_c_970_n 0.0141302f $X=7.04 $Y=0.39 $X2=0 $Y2=0
cc_549 N_X_c_724_n N_VGND_c_970_n 0.00972452f $X=7.765 $Y=0.815 $X2=0 $Y2=0
cc_550 N_X_c_812_n N_VGND_c_970_n 0.0141302f $X=7.98 $Y=0.39 $X2=0 $Y2=0
cc_551 N_X_c_725_n N_VGND_c_970_n 0.00972452f $X=8.705 $Y=0.815 $X2=0 $Y2=0
cc_552 N_X_c_732_n N_VGND_c_970_n 0.020863f $X=8.92 $Y=0.39 $X2=0 $Y2=0
