* File: sky130_fd_sc_hdll__inputiso0p_1.spice
* Created: Thu Aug 27 19:08:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__inputiso0p_1.pex.spice"
.subckt sky130_fd_sc_hdll__inputiso0p_1  VNB VPB SLEEP A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* SLEEP	SLEEP
* VPB	VPB
* VNB	VNB
MM1005 N_A_27_413#_M1005_d N_SLEEP_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.1302 PD=1.36 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 A_307_47# N_A_27_413#_M1007_g N_A_211_413#_M1007_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_M1000_g A_307_47# VNB NSHORT L=0.15 W=0.42 AD=0.113636
+ AS=0.0441 PD=0.92243 PS=0.63 NRD=57.132 NRS=14.28 M=1 R=2.8 SA=75000.5
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1003 N_X_M1003_d N_A_211_413#_M1003_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.175864 PD=1.82 PS=1.42757 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.9 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_SLEEP_M1001_g N_A_27_413#_M1001_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0609 AS=0.1134 PD=0.71 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90002.2 A=0.0756 P=1.2 MULT=1
MM1006 N_A_211_413#_M1006_d N_A_27_413#_M1006_g N_VPWR_M1001_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.0651 AS=0.0609 PD=0.73 PS=0.71 NRD=7.0329 NRS=2.3443 M=1
+ R=2.33333 SA=90000.6 SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_A_211_413#_M1006_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.148331 AS=0.0651 PD=1.08549 PS=0.73 NRD=25.7873 NRS=7.0329 M=1 R=2.33333
+ SA=90001.1 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1004 N_X_M1004_d N_A_211_413#_M1004_g N_VPWR_M1002_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.353169 PD=2.54 PS=2.58451 NRD=0.9653 NRS=98.4803 M=1 R=5.55556
+ SA=90001 SB=90000.2 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.778 P=10.41
pX9_noxref noxref_11 A A PROBETYPE=1
*
.include "sky130_fd_sc_hdll__inputiso0p_1.pxi.spice"
*
.ends
*
*
