* File: sky130_fd_sc_hdll__clkbuf_2.pex.spice
* Created: Wed Sep  2 08:25:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_2%A 1 3 6 8 9
c29 6 0 5.61802e-20 $X=0.525 $Y=0.445
r30 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.16 $X2=0.53 $Y2=1.16
r31 9 14 0.843251 $w=4.08e-07 $l=3e-08 $layer=LI1_cond $X=0.63 $Y=1.19 $X2=0.63
+ $Y2=1.16
r32 8 14 8.71359 $w=4.08e-07 $l=3.1e-07 $layer=LI1_cond $X=0.63 $Y=0.85 $X2=0.63
+ $Y2=1.16
r33 4 13 41.6009 $w=3.62e-07 $l=1.87483e-07 $layer=POLY_cond $X=0.525 $Y=0.975
+ $X2=0.53 $Y2=1.16
r34 4 6 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.525 $Y=0.975
+ $X2=0.525 $Y2=0.445
r35 1 13 45.4695 $w=3.62e-07 $l=2.64575e-07 $layer=POLY_cond $X=0.5 $Y=1.41
+ $X2=0.53 $Y2=1.16
r36 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_2%A_27_47# 1 2 7 9 10 12 13 15 16 18 20 23
+ 25 29 35 37 41
c63 41 0 1.25119e-19 $X=1.495 $Y=1.077
c64 29 0 7.49684e-20 $X=1.1 $Y=1.16
r65 41 42 1.83131 $w=6.58e-07 $l=2.5e-08 $layer=POLY_cond $X=1.495 $Y=1.077
+ $X2=1.52 $Y2=1.077
r66 38 39 1.83131 $w=6.58e-07 $l=2.5e-08 $layer=POLY_cond $X=1 $Y=1.077
+ $X2=1.025 $Y2=1.077
r67 32 35 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.17 $Y=0.42 $X2=0.26
+ $Y2=0.42
r68 30 41 28.9347 $w=6.58e-07 $l=3.95e-07 $layer=POLY_cond $X=1.1 $Y=1.077
+ $X2=1.495 $Y2=1.077
r69 30 39 5.49392 $w=6.58e-07 $l=7.5e-08 $layer=POLY_cond $X=1.1 $Y=1.077
+ $X2=1.025 $Y2=1.077
r70 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.1
+ $Y=1.16 $X2=1.1 $Y2=1.16
r71 27 29 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=1.165 $Y=1.495
+ $X2=1.165 $Y2=1.16
r72 26 37 2.28545 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.355 $Y=1.58
+ $X2=0.22 $Y2=1.58
r73 25 27 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.015 $Y=1.58
+ $X2=1.165 $Y2=1.495
r74 25 26 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.015 $Y=1.58
+ $X2=0.355 $Y2=1.58
r75 21 37 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.22 $Y=1.665
+ $X2=0.22 $Y2=1.58
r76 21 23 3.41465 $w=2.68e-07 $l=8e-08 $layer=LI1_cond $X=0.22 $Y=1.665 $X2=0.22
+ $Y2=1.745
r77 20 37 4.14756 $w=2.2e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.17 $Y=1.495
+ $X2=0.22 $Y2=1.58
r78 19 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.17 $Y2=0.42
r79 19 20 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.17 $Y2=1.495
r80 16 42 38.4816 $w=1.5e-07 $l=3.32e-07 $layer=POLY_cond $X=1.52 $Y=0.745
+ $X2=1.52 $Y2=1.077
r81 16 18 96.4 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=1.52 $Y=0.745 $X2=1.52
+ $Y2=0.445
r82 13 41 33.7549 $w=1.8e-07 $l=3.33e-07 $layer=POLY_cond $X=1.495 $Y=1.41
+ $X2=1.495 $Y2=1.077
r83 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.495 $Y=1.41
+ $X2=1.495 $Y2=1.985
r84 10 39 33.7549 $w=1.8e-07 $l=3.33e-07 $layer=POLY_cond $X=1.025 $Y=1.41
+ $X2=1.025 $Y2=1.077
r85 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.025 $Y=1.41
+ $X2=1.025 $Y2=1.985
r86 7 38 38.4816 $w=1.5e-07 $l=3.32e-07 $layer=POLY_cond $X=1 $Y=0.745 $X2=1
+ $Y2=1.077
r87 7 9 96.4 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=1 $Y=0.745 $X2=1 $Y2=0.445
r88 2 23 300 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.745
r89 1 35 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_2%VPWR 1 2 9 13 15 17 22 29 30 33 36
r33 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r34 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r35 30 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r36 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r37 27 36 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.9 $Y=2.72
+ $X2=1.707 $Y2=2.72
r38 27 29 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.9 $Y=2.72 $X2=2.07
+ $Y2=2.72
r39 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r40 26 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r41 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r42 23 33 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.905 $Y=2.72
+ $X2=0.715 $Y2=2.72
r43 23 25 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.905 $Y=2.72
+ $X2=1.15 $Y2=2.72
r44 22 36 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=1.515 $Y=2.72
+ $X2=1.707 $Y2=2.72
r45 22 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.515 $Y=2.72
+ $X2=1.15 $Y2=2.72
r46 17 33 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.715 $Y2=2.72
r47 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.23 $Y2=2.72
r48 15 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r49 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r50 11 36 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.707 $Y=2.635
+ $X2=1.707 $Y2=2.72
r51 11 13 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=1.707 $Y=2.635
+ $X2=1.707 $Y2=2.295
r52 7 33 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=2.635
+ $X2=0.715 $Y2=2.72
r53 7 9 21.0776 $w=3.78e-07 $l=6.95e-07 $layer=LI1_cond $X=0.715 $Y=2.635
+ $X2=0.715 $Y2=1.94
r54 2 13 600 $w=1.7e-07 $l=8.79517e-07 $layer=licon1_PDIFF $count=1 $X=1.585
+ $Y=1.485 $X2=1.73 $Y2=2.295
r55 1 9 300 $w=1.7e-07 $l=5.24667e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=1.485 $X2=0.74 $Y2=1.94
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_2%X 1 2 9 13 15 16 17 18 28 46
c40 15 0 5.61802e-20 $X=1.675 $Y=0.765
c41 2 0 7.49684e-20 $X=1.115 $Y=1.485
r42 43 46 22.6888 $w=1.73e-07 $l=3.58e-07 $layer=LI1_cond $X=1.252 $Y=1.942
+ $X2=1.61 $Y2=1.942
r43 26 46 4.43636 $w=1.73e-07 $l=7e-08 $layer=LI1_cond $X=1.68 $Y=1.942 $X2=1.61
+ $Y2=1.942
r44 25 28 0.738746 $w=3.88e-07 $l=2.5e-08 $layer=LI1_cond $X=1.68 $Y=0.825
+ $X2=1.68 $Y2=0.85
r45 18 26 5.07013 $w=1.73e-07 $l=8e-08 $layer=LI1_cond $X=1.76 $Y=1.942 $X2=1.68
+ $Y2=1.942
r46 18 26 1.03424 $w=3.88e-07 $l=3.5e-08 $layer=LI1_cond $X=1.68 $Y=1.82
+ $X2=1.68 $Y2=1.855
r47 17 18 8.56945 $w=3.88e-07 $l=2.9e-07 $layer=LI1_cond $X=1.68 $Y=1.53
+ $X2=1.68 $Y2=1.82
r48 16 17 10.0469 $w=3.88e-07 $l=3.4e-07 $layer=LI1_cond $X=1.68 $Y=1.19
+ $X2=1.68 $Y2=1.53
r49 15 25 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.76 $Y=0.74 $X2=1.68
+ $Y2=0.74
r50 15 16 9.16044 $w=3.88e-07 $l=3.1e-07 $layer=LI1_cond $X=1.68 $Y=0.88
+ $X2=1.68 $Y2=1.19
r51 15 28 0.886495 $w=3.88e-07 $l=3e-08 $layer=LI1_cond $X=1.68 $Y=0.88 $X2=1.68
+ $Y2=0.85
r52 11 43 0.409621 $w=1.85e-07 $l=8.8e-08 $layer=LI1_cond $X=1.252 $Y=2.03
+ $X2=1.252 $Y2=1.942
r53 11 13 14.3882 $w=1.83e-07 $l=2.4e-07 $layer=LI1_cond $X=1.252 $Y=2.03
+ $X2=1.252 $Y2=2.27
r54 7 25 28.5754 $w=1.68e-07 $l=4.38e-07 $layer=LI1_cond $X=1.242 $Y=0.74
+ $X2=1.68 $Y2=0.74
r55 7 9 12.714 $w=2.03e-07 $l=2.35e-07 $layer=LI1_cond $X=1.242 $Y=0.655
+ $X2=1.242 $Y2=0.42
r56 2 13 600 $w=1.7e-07 $l=8.5443e-07 $layer=licon1_PDIFF $count=1 $X=1.115
+ $Y=1.485 $X2=1.26 $Y2=2.27
r57 1 9 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_2%VGND 1 2 9 13 15 17 22 29 30 33 36
c32 22 0 1.25119e-19 $X=1.515 $Y=0
r33 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r34 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r35 30 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r36 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r37 27 36 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.9 $Y=0 $X2=1.707
+ $Y2=0
r38 27 29 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.9 $Y=0 $X2=2.07
+ $Y2=0
r39 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r40 26 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r41 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r42 23 33 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.742
+ $Y2=0
r43 23 25 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=1.15
+ $Y2=0
r44 22 36 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=1.515 $Y=0 $X2=1.707
+ $Y2=0
r45 22 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.515 $Y=0 $X2=1.15
+ $Y2=0
r46 17 33 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.742
+ $Y2=0
r47 17 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.23
+ $Y2=0
r48 15 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r49 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r50 11 36 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.707 $Y=0.085
+ $X2=1.707 $Y2=0
r51 11 13 9.42908 $w=3.83e-07 $l=3.15e-07 $layer=LI1_cond $X=1.707 $Y=0.085
+ $X2=1.707 $Y2=0.4
r52 7 33 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.742 $Y=0.085
+ $X2=0.742 $Y2=0
r53 7 9 13.2007 $w=2.73e-07 $l=3.15e-07 $layer=LI1_cond $X=0.742 $Y=0.085
+ $X2=0.742 $Y2=0.4
r54 2 13 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.73 $Y2=0.4
r55 1 9 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.235 $X2=0.74 $Y2=0.4
.ends

