* NGSPICE file created from sky130_fd_sc_hdll__tapvpwrvgnd_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__tapvpwrvgnd_1 VGND VPWR
.ends

