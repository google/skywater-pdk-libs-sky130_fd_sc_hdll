* NGSPICE file created from sky130_fd_sc_hdll__nor2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__nor2_2 A B VGND VNB VPB VPWR Y
M1000 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=8.5e+11p ps=7.7e+06u
M1001 a_27_297# B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1002 Y B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A VGND VNB nshort w=650000u l=150000u
+  ad=4.81e+11p pd=4.08e+06u as=6.0125e+11p ps=5.75e+06u
M1004 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

