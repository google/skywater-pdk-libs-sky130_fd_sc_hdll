* File: sky130_fd_sc_hdll__nand2_8.pex.spice
* Created: Wed Sep  2 08:37:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND2_8%B 3 5 7 10 12 14 17 19 21 24 26 28 31 33
+ 35 38 40 42 45 47 49 50 52 55 57 58 59 60 61 62 88 89 94 97 100 103 106 109
c164 88 0 1.83863e-19 $X=3.55 $Y=1.16
c165 55 0 8.09502e-20 $X=3.81 $Y=0.56
r166 89 90 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=3.785 $Y=1.217
+ $X2=3.81 $Y2=1.217
r167 88 109 29.073 $w=2.18e-07 $l=5.55e-07 $layer=LI1_cond $X=3.55 $Y=1.185
+ $X2=2.995 $Y2=1.185
r168 87 89 35.177 $w=3.22e-07 $l=2.35e-07 $layer=POLY_cond $X=3.55 $Y=1.217
+ $X2=3.785 $Y2=1.217
r169 87 88 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=3.55
+ $Y=1.16 $X2=3.55 $Y2=1.16
r170 85 87 35.177 $w=3.22e-07 $l=2.35e-07 $layer=POLY_cond $X=3.315 $Y=1.217
+ $X2=3.55 $Y2=1.217
r171 84 85 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.217
+ $X2=3.315 $Y2=1.217
r172 83 84 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=2.845 $Y=1.217
+ $X2=3.29 $Y2=1.217
r173 82 83 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.217
+ $X2=2.845 $Y2=1.217
r174 81 82 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=2.375 $Y=1.217
+ $X2=2.82 $Y2=1.217
r175 80 81 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.217
+ $X2=2.375 $Y2=1.217
r176 79 80 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=1.905 $Y=1.217
+ $X2=2.35 $Y2=1.217
r177 78 79 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=1.88 $Y=1.217
+ $X2=1.905 $Y2=1.217
r178 77 78 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=1.435 $Y=1.217
+ $X2=1.88 $Y2=1.217
r179 76 77 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.217
+ $X2=1.435 $Y2=1.217
r180 75 76 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=0.965 $Y=1.217
+ $X2=1.41 $Y2=1.217
r181 74 75 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.217
+ $X2=0.965 $Y2=1.217
r182 72 74 32.1832 $w=3.22e-07 $l=2.15e-07 $layer=POLY_cond $X=0.725 $Y=1.217
+ $X2=0.94 $Y2=1.217
r183 72 94 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=0.725
+ $Y=1.16 $X2=0.725 $Y2=1.16
r184 70 72 34.4286 $w=3.22e-07 $l=2.3e-07 $layer=POLY_cond $X=0.495 $Y=1.217
+ $X2=0.725 $Y2=1.217
r185 69 70 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.217
+ $X2=0.495 $Y2=1.217
r186 62 109 0.261919 $w=2.18e-07 $l=5e-09 $layer=LI1_cond $X=2.99 $Y=1.185
+ $X2=2.995 $Y2=1.185
r187 62 106 23.8346 $w=2.18e-07 $l=4.55e-07 $layer=LI1_cond $X=2.99 $Y=1.185
+ $X2=2.535 $Y2=1.185
r188 61 106 0.261919 $w=2.18e-07 $l=5e-09 $layer=LI1_cond $X=2.53 $Y=1.185
+ $X2=2.535 $Y2=1.185
r189 61 103 23.8346 $w=2.18e-07 $l=4.55e-07 $layer=LI1_cond $X=2.53 $Y=1.185
+ $X2=2.075 $Y2=1.185
r190 60 103 0.261919 $w=2.18e-07 $l=5e-09 $layer=LI1_cond $X=2.07 $Y=1.185
+ $X2=2.075 $Y2=1.185
r191 60 100 23.8346 $w=2.18e-07 $l=4.55e-07 $layer=LI1_cond $X=2.07 $Y=1.185
+ $X2=1.615 $Y2=1.185
r192 59 100 0.261919 $w=2.18e-07 $l=5e-09 $layer=LI1_cond $X=1.61 $Y=1.185
+ $X2=1.615 $Y2=1.185
r193 59 97 23.8346 $w=2.18e-07 $l=4.55e-07 $layer=LI1_cond $X=1.61 $Y=1.185
+ $X2=1.155 $Y2=1.185
r194 58 97 0.261919 $w=2.18e-07 $l=5e-09 $layer=LI1_cond $X=1.15 $Y=1.185
+ $X2=1.155 $Y2=1.185
r195 58 94 23.8346 $w=2.18e-07 $l=4.55e-07 $layer=LI1_cond $X=1.15 $Y=1.185
+ $X2=0.695 $Y2=1.185
r196 57 94 0.261919 $w=2.18e-07 $l=5e-09 $layer=LI1_cond $X=0.69 $Y=1.185
+ $X2=0.695 $Y2=1.185
r197 53 90 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.81 $Y=1.025
+ $X2=3.81 $Y2=1.217
r198 53 55 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.81 $Y=1.025
+ $X2=3.81 $Y2=0.56
r199 50 89 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.217
r200 50 52 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r201 47 85 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.217
r202 47 49 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r203 43 84 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=1.217
r204 43 45 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=0.56
r205 40 83 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.217
r206 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r207 36 82 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.82 $Y=1.025
+ $X2=2.82 $Y2=1.217
r208 36 38 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.82 $Y=1.025
+ $X2=2.82 $Y2=0.56
r209 33 81 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.217
r210 33 35 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r211 29 80 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=1.217
r212 29 31 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=0.56
r213 26 79 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.217
r214 26 28 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r215 22 78 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.88 $Y=1.025
+ $X2=1.88 $Y2=1.217
r216 22 24 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.88 $Y=1.025
+ $X2=1.88 $Y2=0.56
r217 19 77 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.217
r218 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r219 15 76 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=1.217
r220 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=0.56
r221 12 75 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.217
r222 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r223 8 74 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.94 $Y=1.025
+ $X2=0.94 $Y2=1.217
r224 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.94 $Y=1.025
+ $X2=0.94 $Y2=0.56
r225 5 70 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.217
r226 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r227 1 69 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=1.217
r228 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_8%A 3 5 7 10 12 14 17 19 21 24 26 28 31 33
+ 35 38 40 42 45 47 49 50 52 55 57 58 59 60 61 84 87 92 96 99 102
c132 87 0 1.83863e-19 $X=7.545 $Y=1.217
c133 3 0 1.56255e-19 $X=4.23 $Y=0.56
r134 87 88 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=7.545 $Y=1.217
+ $X2=7.57 $Y2=1.217
r135 86 87 70.354 $w=3.22e-07 $l=4.7e-07 $layer=POLY_cond $X=7.075 $Y=1.217
+ $X2=7.545 $Y2=1.217
r136 85 86 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=7.05 $Y=1.217
+ $X2=7.075 $Y2=1.217
r137 83 85 31.4348 $w=3.22e-07 $l=2.1e-07 $layer=POLY_cond $X=6.84 $Y=1.217
+ $X2=7.05 $Y2=1.217
r138 83 84 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=6.84
+ $Y=1.16 $X2=6.84 $Y2=1.16
r139 81 83 35.177 $w=3.22e-07 $l=2.35e-07 $layer=POLY_cond $X=6.605 $Y=1.217
+ $X2=6.84 $Y2=1.217
r140 80 81 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=6.58 $Y=1.217
+ $X2=6.605 $Y2=1.217
r141 79 80 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=6.135 $Y=1.217
+ $X2=6.58 $Y2=1.217
r142 78 79 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=6.11 $Y=1.217
+ $X2=6.135 $Y2=1.217
r143 77 78 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=5.665 $Y=1.217
+ $X2=6.11 $Y2=1.217
r144 76 77 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=5.64 $Y=1.217
+ $X2=5.665 $Y2=1.217
r145 75 76 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=5.195 $Y=1.217
+ $X2=5.64 $Y2=1.217
r146 74 75 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=5.17 $Y=1.217
+ $X2=5.195 $Y2=1.217
r147 73 92 6.93182 $w=1.98e-07 $l=1.25e-07 $layer=LI1_cond $X=4.96 $Y=1.175
+ $X2=4.835 $Y2=1.175
r148 72 74 31.4348 $w=3.22e-07 $l=2.1e-07 $layer=POLY_cond $X=4.96 $Y=1.217
+ $X2=5.17 $Y2=1.217
r149 72 73 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.96
+ $Y=1.16 $X2=4.96 $Y2=1.16
r150 70 72 35.177 $w=3.22e-07 $l=2.35e-07 $layer=POLY_cond $X=4.725 $Y=1.217
+ $X2=4.96 $Y2=1.217
r151 69 70 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=4.7 $Y=1.217
+ $X2=4.725 $Y2=1.217
r152 68 69 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=4.255 $Y=1.217
+ $X2=4.7 $Y2=1.217
r153 67 68 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=4.23 $Y=1.217
+ $X2=4.255 $Y2=1.217
r154 61 84 9.42727 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=6.67 $Y=1.175
+ $X2=6.84 $Y2=1.175
r155 61 102 25.2318 $w=1.98e-07 $l=4.55e-07 $layer=LI1_cond $X=6.67 $Y=1.175
+ $X2=6.215 $Y2=1.175
r156 60 102 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=6.21 $Y=1.175
+ $X2=6.215 $Y2=1.175
r157 60 99 25.2318 $w=1.98e-07 $l=4.55e-07 $layer=LI1_cond $X=6.21 $Y=1.175
+ $X2=5.755 $Y2=1.175
r158 59 99 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=5.75 $Y=1.175
+ $X2=5.755 $Y2=1.175
r159 59 96 25.2318 $w=1.98e-07 $l=4.55e-07 $layer=LI1_cond $X=5.75 $Y=1.175
+ $X2=5.295 $Y2=1.175
r160 58 96 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=5.29 $Y=1.175
+ $X2=5.295 $Y2=1.175
r161 58 73 18.3 $w=1.98e-07 $l=3.3e-07 $layer=LI1_cond $X=5.29 $Y=1.175 $X2=4.96
+ $Y2=1.175
r162 57 92 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=4.83 $Y=1.175
+ $X2=4.835 $Y2=1.175
r163 53 88 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.57 $Y=1.025
+ $X2=7.57 $Y2=1.217
r164 53 55 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.57 $Y=1.025
+ $X2=7.57 $Y2=0.56
r165 50 87 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.217
r166 50 52 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.985
r167 47 86 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.217
r168 47 49 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.985
r169 43 85 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.05 $Y=1.025
+ $X2=7.05 $Y2=1.217
r170 43 45 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.05 $Y=1.025
+ $X2=7.05 $Y2=0.56
r171 40 81 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.217
r172 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.985
r173 36 80 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.58 $Y=1.025
+ $X2=6.58 $Y2=1.217
r174 36 38 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.58 $Y=1.025
+ $X2=6.58 $Y2=0.56
r175 33 79 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.217
r176 33 35 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.985
r177 29 78 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.11 $Y=1.025
+ $X2=6.11 $Y2=1.217
r178 29 31 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.11 $Y=1.025
+ $X2=6.11 $Y2=0.56
r179 26 77 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.217
r180 26 28 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.985
r181 22 76 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.64 $Y=1.025
+ $X2=5.64 $Y2=1.217
r182 22 24 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.64 $Y=1.025
+ $X2=5.64 $Y2=0.56
r183 19 75 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.217
r184 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.985
r185 15 74 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.17 $Y=1.025
+ $X2=5.17 $Y2=1.217
r186 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.17 $Y=1.025
+ $X2=5.17 $Y2=0.56
r187 12 70 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.217
r188 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.985
r189 8 69 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.7 $Y=1.025
+ $X2=4.7 $Y2=1.217
r190 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.7 $Y=1.025
+ $X2=4.7 $Y2=0.56
r191 5 68 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.217
r192 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.985
r193 1 67 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.23 $Y=1.025
+ $X2=4.23 $Y2=1.217
r194 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.23 $Y=1.025
+ $X2=4.23 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_8%VPWR 1 2 3 4 5 6 7 8 9 28 30 34 38 40 44
+ 48 52 56 60 64 66 68 73 74 76 77 79 80 82 83 85 86 87 105 113 116 120
r136 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r137 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r138 114 117 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r139 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r140 108 120 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r141 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r142 105 119 4.76767 $w=1.7e-07 $l=2.82e-07 $layer=LI1_cond $X=7.715 $Y=2.72
+ $X2=7.997 $Y2=2.72
r143 105 107 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.715 $Y=2.72
+ $X2=7.59 $Y2=2.72
r144 104 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r145 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r146 101 104 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r147 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r148 98 101 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r149 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r150 95 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r151 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r152 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r153 92 117 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r154 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r155 89 116 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.14 $Y2=2.72
r156 89 91 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.99 $Y2=2.72
r157 87 114 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r158 87 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r159 85 103 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.755 $Y=2.72
+ $X2=6.67 $Y2=2.72
r160 85 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.755 $Y=2.72
+ $X2=6.84 $Y2=2.72
r161 84 107 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=6.925 $Y=2.72
+ $X2=7.59 $Y2=2.72
r162 84 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.925 $Y=2.72
+ $X2=6.84 $Y2=2.72
r163 82 100 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.815 $Y=2.72
+ $X2=5.75 $Y2=2.72
r164 82 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.815 $Y=2.72
+ $X2=5.9 $Y2=2.72
r165 81 103 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=5.985 $Y=2.72
+ $X2=6.67 $Y2=2.72
r166 81 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.985 $Y=2.72
+ $X2=5.9 $Y2=2.72
r167 79 97 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.875 $Y=2.72
+ $X2=4.83 $Y2=2.72
r168 79 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.875 $Y=2.72
+ $X2=4.96 $Y2=2.72
r169 78 100 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=5.045 $Y=2.72
+ $X2=5.75 $Y2=2.72
r170 78 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=2.72
+ $X2=4.96 $Y2=2.72
r171 76 94 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.935 $Y=2.72
+ $X2=3.91 $Y2=2.72
r172 76 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=2.72
+ $X2=4.02 $Y2=2.72
r173 75 97 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=4.105 $Y=2.72
+ $X2=4.83 $Y2=2.72
r174 75 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=2.72
+ $X2=4.02 $Y2=2.72
r175 73 91 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.995 $Y=2.72
+ $X2=2.99 $Y2=2.72
r176 73 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=2.72
+ $X2=3.08 $Y2=2.72
r177 72 94 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3.165 $Y=2.72
+ $X2=3.91 $Y2=2.72
r178 72 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=2.72
+ $X2=3.08 $Y2=2.72
r179 68 71 22.075 $w=3.53e-07 $l=6.8e-07 $layer=LI1_cond $X=7.892 $Y=1.66
+ $X2=7.892 $Y2=2.34
r180 66 119 3.21226 $w=3.55e-07 $l=1.41244e-07 $layer=LI1_cond $X=7.892 $Y=2.635
+ $X2=7.997 $Y2=2.72
r181 66 71 9.57664 $w=3.53e-07 $l=2.95e-07 $layer=LI1_cond $X=7.892 $Y=2.635
+ $X2=7.892 $Y2=2.34
r182 62 86 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=2.635
+ $X2=6.84 $Y2=2.72
r183 62 64 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.84 $Y=2.635
+ $X2=6.84 $Y2=2
r184 58 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=2.635 $X2=5.9
+ $Y2=2.72
r185 58 60 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.9 $Y=2.635
+ $X2=5.9 $Y2=2
r186 54 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=2.72
r187 54 56 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=2
r188 50 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=2.72
r189 50 52 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=2
r190 46 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2.72
r191 46 48 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2
r192 42 116 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.72
r193 42 44 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2
r194 41 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=1.2 $Y2=2.72
r195 40 116 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=2.14 $Y2=2.72
r196 40 41 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=1.285 $Y2=2.72
r197 36 113 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.72
r198 36 38 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r199 35 110 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r200 34 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=1.2 $Y2=2.72
r201 34 35 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=0.345 $Y2=2.72
r202 30 33 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.34
r203 28 110 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r204 28 33 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.34
r205 9 71 400 $w=1.7e-07 $l=9.69794e-07 $layer=licon1_PDIFF $count=1 $X=7.635
+ $Y=1.485 $X2=7.88 $Y2=2.34
r206 9 68 400 $w=1.7e-07 $l=3.2078e-07 $layer=licon1_PDIFF $count=1 $X=7.635
+ $Y=1.485 $X2=7.88 $Y2=1.66
r207 8 64 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.695
+ $Y=1.485 $X2=6.84 $Y2=2
r208 7 60 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.755
+ $Y=1.485 $X2=5.9 $Y2=2
r209 6 56 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=2
r210 5 52 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=2
r211 4 48 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2
r212 3 44 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r213 2 38 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r214 1 33 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r215 1 30 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_8%Y 1 2 3 4 5 6 7 8 9 10 11 12 37 39 41 45
+ 47 51 53 57 59 61 62 65 67 73 74 77 79 83 85 89 91 92 96 98 100 104 106 108
+ 111
c208 91 0 1.21485e-19 $X=7.35 $Y=0.905
c209 61 0 8.09502e-20 $X=4.422 $Y=0.905
r210 118 120 0.978731 $w=5.36e-07 $l=4.3e-08 $layer=LI1_cond $X=4.422 $Y=1.37
+ $X2=4.465 $Y2=1.37
r211 111 118 1.18358 $w=5.36e-07 $l=5.2e-08 $layer=LI1_cond $X=4.37 $Y=1.37
+ $X2=4.422 $Y2=1.37
r212 92 108 3.48797 $w=3.15e-07 $l=1.28452e-07 $layer=LI1_cond $X=7.35 $Y=1.465
+ $X2=7.285 $Y2=1.565
r213 91 110 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=7.35 $Y=0.905
+ $X2=7.35 $Y2=0.78
r214 91 92 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=7.35 $Y=0.905
+ $X2=7.35 $Y2=1.465
r215 87 108 3.48797 $w=3.15e-07 $l=1e-07 $layer=LI1_cond $X=7.285 $Y=1.665
+ $X2=7.285 $Y2=1.565
r216 87 89 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=7.285 $Y=1.665
+ $X2=7.285 $Y2=2.34
r217 86 106 8.48182 $w=2e-07 $l=1.9e-07 $layer=LI1_cond $X=6.535 $Y=1.565
+ $X2=6.345 $Y2=1.565
r218 85 108 3.01902 $w=2e-07 $l=1.9e-07 $layer=LI1_cond $X=7.095 $Y=1.565
+ $X2=7.285 $Y2=1.565
r219 85 86 31.0545 $w=1.98e-07 $l=5.6e-07 $layer=LI1_cond $X=7.095 $Y=1.565
+ $X2=6.535 $Y2=1.565
r220 81 106 0.829748 $w=3.8e-07 $l=1e-07 $layer=LI1_cond $X=6.345 $Y=1.665
+ $X2=6.345 $Y2=1.565
r221 81 83 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=6.345 $Y=1.665
+ $X2=6.345 $Y2=2.34
r222 80 104 8.48182 $w=2e-07 $l=1.9e-07 $layer=LI1_cond $X=5.595 $Y=1.565
+ $X2=5.405 $Y2=1.565
r223 79 106 8.48182 $w=2e-07 $l=1.9e-07 $layer=LI1_cond $X=6.155 $Y=1.565
+ $X2=6.345 $Y2=1.565
r224 79 80 31.0545 $w=1.98e-07 $l=5.6e-07 $layer=LI1_cond $X=6.155 $Y=1.565
+ $X2=5.595 $Y2=1.565
r225 75 104 0.829748 $w=3.8e-07 $l=1e-07 $layer=LI1_cond $X=5.405 $Y=1.665
+ $X2=5.405 $Y2=1.565
r226 75 77 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=5.405 $Y=1.665
+ $X2=5.405 $Y2=2.34
r227 74 120 9.34666 $w=5.36e-07 $l=2.73998e-07 $layer=LI1_cond $X=4.655 $Y=1.565
+ $X2=4.465 $Y2=1.37
r228 73 104 8.48182 $w=2e-07 $l=1.9e-07 $layer=LI1_cond $X=5.215 $Y=1.565
+ $X2=5.405 $Y2=1.565
r229 73 74 31.0545 $w=1.98e-07 $l=5.6e-07 $layer=LI1_cond $X=5.215 $Y=1.565
+ $X2=4.655 $Y2=1.565
r230 70 72 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=5.43 $Y=0.78
+ $X2=6.37 $Y2=0.78
r231 68 102 3.72825 $w=2.5e-07 $l=1.48e-07 $layer=LI1_cond $X=4.57 $Y=0.78
+ $X2=4.422 $Y2=0.78
r232 68 70 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=4.57 $Y=0.78
+ $X2=5.43 $Y2=0.78
r233 67 110 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=7.225 $Y=0.78
+ $X2=7.35 $Y2=0.78
r234 67 72 39.4136 $w=2.48e-07 $l=8.55e-07 $layer=LI1_cond $X=7.225 $Y=0.78
+ $X2=6.37 $Y2=0.78
r235 63 120 2.7522 $w=3.8e-07 $l=2.95e-07 $layer=LI1_cond $X=4.465 $Y=1.665
+ $X2=4.465 $Y2=1.37
r236 63 65 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=4.465 $Y=1.665
+ $X2=4.465 $Y2=2.34
r237 62 118 4.2441 $w=2.95e-07 $l=2.95e-07 $layer=LI1_cond $X=4.422 $Y=1.075
+ $X2=4.422 $Y2=1.37
r238 61 102 3.14886 $w=2.95e-07 $l=1.25e-07 $layer=LI1_cond $X=4.422 $Y=0.905
+ $X2=4.422 $Y2=0.78
r239 61 62 6.6412 $w=2.93e-07 $l=1.7e-07 $layer=LI1_cond $X=4.422 $Y=0.905
+ $X2=4.422 $Y2=1.075
r240 60 100 8.48182 $w=2e-07 $l=1.9e-07 $layer=LI1_cond $X=3.715 $Y=1.565
+ $X2=3.525 $Y2=1.565
r241 59 111 12.5332 $w=5.36e-07 $l=4.16233e-07 $layer=LI1_cond $X=4.04 $Y=1.565
+ $X2=4.37 $Y2=1.37
r242 59 60 18.0227 $w=1.98e-07 $l=3.25e-07 $layer=LI1_cond $X=4.04 $Y=1.565
+ $X2=3.715 $Y2=1.565
r243 55 100 0.829748 $w=3.8e-07 $l=1e-07 $layer=LI1_cond $X=3.525 $Y=1.665
+ $X2=3.525 $Y2=1.565
r244 55 57 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=3.525 $Y=1.665
+ $X2=3.525 $Y2=2.34
r245 54 98 8.48182 $w=2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=1.565
+ $X2=2.585 $Y2=1.565
r246 53 100 8.48182 $w=2e-07 $l=1.9e-07 $layer=LI1_cond $X=3.335 $Y=1.565
+ $X2=3.525 $Y2=1.565
r247 53 54 31.0545 $w=1.98e-07 $l=5.6e-07 $layer=LI1_cond $X=3.335 $Y=1.565
+ $X2=2.775 $Y2=1.565
r248 49 98 0.829748 $w=3.8e-07 $l=1e-07 $layer=LI1_cond $X=2.585 $Y=1.665
+ $X2=2.585 $Y2=1.565
r249 49 51 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=2.585 $Y=1.665
+ $X2=2.585 $Y2=2.34
r250 48 96 8.48182 $w=2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=1.565
+ $X2=1.645 $Y2=1.565
r251 47 98 8.48182 $w=2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=1.565
+ $X2=2.585 $Y2=1.565
r252 47 48 31.0545 $w=1.98e-07 $l=5.6e-07 $layer=LI1_cond $X=2.395 $Y=1.565
+ $X2=1.835 $Y2=1.565
r253 43 96 0.829748 $w=3.8e-07 $l=1e-07 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.645 $Y2=1.565
r254 43 45 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.645 $Y2=2.34
r255 42 94 5.04956 $w=2e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=1.565
+ $X2=0.705 $Y2=1.565
r256 41 96 8.48182 $w=2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=1.565
+ $X2=1.645 $Y2=1.565
r257 41 42 31.0545 $w=1.98e-07 $l=5.6e-07 $layer=LI1_cond $X=1.455 $Y=1.565
+ $X2=0.895 $Y2=1.565
r258 37 94 2.65766 $w=3.8e-07 $l=1e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=1.565
r259 37 39 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=2.34
r260 12 108 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=7.165
+ $Y=1.485 $X2=7.31 $Y2=1.66
r261 12 89 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.165
+ $Y=1.485 $X2=7.31 $Y2=2.34
r262 11 106 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=6.225
+ $Y=1.485 $X2=6.37 $Y2=1.66
r263 11 83 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.225
+ $Y=1.485 $X2=6.37 $Y2=2.34
r264 10 104 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=1.66
r265 10 77 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=2.34
r266 9 120 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=1.66
r267 9 65 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=2.34
r268 8 100 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.66
r269 8 57 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2.34
r270 7 98 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.66
r271 7 51 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.34
r272 6 96 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r273 6 45 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
r274 5 94 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r275 5 39 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r276 4 110 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=7.125
+ $Y=0.235 $X2=7.31 $Y2=0.74
r277 3 72 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=6.185
+ $Y=0.235 $X2=6.37 $Y2=0.74
r278 2 70 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=5.245
+ $Y=0.235 $X2=5.43 $Y2=0.74
r279 1 102 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.235 $X2=4.49 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_8%A_27_47# 1 2 3 4 5 6 7 8 9 30 32 33 36 38
+ 42 44 48 50 52 53 54 62 64 66 67 68
c135 53 0 1.56255e-19 $X=3.955 $Y=0.735
r136 62 74 2.79446 $w=3.75e-07 $l=1.15e-07 $layer=LI1_cond $X=7.882 $Y=0.485
+ $X2=7.882 $Y2=0.37
r137 62 64 7.83661 $w=3.73e-07 $l=2.55e-07 $layer=LI1_cond $X=7.882 $Y=0.485
+ $X2=7.882 $Y2=0.74
r138 59 61 47.0998 $w=2.28e-07 $l=9.4e-07 $layer=LI1_cond $X=5.9 $Y=0.37
+ $X2=6.84 $Y2=0.37
r139 57 59 47.0998 $w=2.28e-07 $l=9.4e-07 $layer=LI1_cond $X=4.96 $Y=0.37
+ $X2=5.9 $Y2=0.37
r140 55 70 3.94658 $w=2.3e-07 $l=1.5e-07 $layer=LI1_cond $X=4.105 $Y=0.37
+ $X2=3.955 $Y2=0.37
r141 55 57 42.8408 $w=2.28e-07 $l=8.55e-07 $layer=LI1_cond $X=4.105 $Y=0.37
+ $X2=4.96 $Y2=0.37
r142 54 74 4.54403 $w=2.3e-07 $l=1.87e-07 $layer=LI1_cond $X=7.695 $Y=0.37
+ $X2=7.882 $Y2=0.37
r143 54 61 42.8408 $w=2.28e-07 $l=8.55e-07 $layer=LI1_cond $X=7.695 $Y=0.37
+ $X2=6.84 $Y2=0.37
r144 53 72 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.955 $Y=0.735
+ $X2=3.955 $Y2=0.82
r145 52 70 3.02571 $w=3e-07 $l=1.15e-07 $layer=LI1_cond $X=3.955 $Y=0.485
+ $X2=3.955 $Y2=0.37
r146 52 53 9.60369 $w=2.98e-07 $l=2.5e-07 $layer=LI1_cond $X=3.955 $Y=0.485
+ $X2=3.955 $Y2=0.735
r147 51 68 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.245 $Y=0.82
+ $X2=3.055 $Y2=0.82
r148 50 72 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.805 $Y=0.82
+ $X2=3.955 $Y2=0.82
r149 50 51 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.805 $Y=0.82
+ $X2=3.245 $Y2=0.82
r150 46 68 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=0.735
+ $X2=3.055 $Y2=0.82
r151 46 48 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.055 $Y=0.735
+ $X2=3.055 $Y2=0.4
r152 45 67 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.305 $Y=0.82
+ $X2=2.115 $Y2=0.82
r153 44 68 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.865 $Y=0.82
+ $X2=3.055 $Y2=0.82
r154 44 45 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.865 $Y=0.82
+ $X2=2.305 $Y2=0.82
r155 40 67 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.115 $Y=0.735
+ $X2=2.115 $Y2=0.82
r156 40 42 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.115 $Y=0.735
+ $X2=2.115 $Y2=0.4
r157 39 66 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.365 $Y=0.82
+ $X2=1.175 $Y2=0.82
r158 38 67 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.925 $Y=0.82
+ $X2=2.115 $Y2=0.82
r159 38 39 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.925 $Y=0.82
+ $X2=1.365 $Y2=0.82
r160 34 66 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=0.735
+ $X2=1.175 $Y2=0.82
r161 34 36 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.175 $Y=0.735
+ $X2=1.175 $Y2=0.4
r162 32 66 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.985 $Y=0.82
+ $X2=1.175 $Y2=0.82
r163 32 33 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.985 $Y=0.82
+ $X2=0.425 $Y2=0.82
r164 28 33 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.425 $Y2=0.82
r165 28 30 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.257 $Y2=0.4
r166 9 74 182 $w=1.7e-07 $l=3.06594e-07 $layer=licon1_NDIFF $count=1 $X=7.645
+ $Y=0.235 $X2=7.88 $Y2=0.4
r167 9 64 182 $w=1.7e-07 $l=6.1131e-07 $layer=licon1_NDIFF $count=1 $X=7.645
+ $Y=0.235 $X2=7.88 $Y2=0.74
r168 8 61 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=6.655
+ $Y=0.235 $X2=6.84 $Y2=0.4
r169 7 59 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=5.715
+ $Y=0.235 $X2=5.9 $Y2=0.4
r170 6 57 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.235 $X2=4.96 $Y2=0.4
r171 5 72 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.235 $X2=4.02 $Y2=0.74
r172 5 70 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.235 $X2=4.02 $Y2=0.4
r173 4 48 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.4
r174 3 42 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=1.955
+ $Y=0.235 $X2=2.14 $Y2=0.4
r175 2 36 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.4
r176 1 30 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_8%VGND 1 2 3 4 17 19 23 25 29 33 36 37 38 48
+ 49 52 55 58
r106 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r107 56 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r108 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r109 53 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r110 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r111 48 49 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r112 46 49 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=3.91 $Y=0 $X2=8.05
+ $Y2=0
r113 45 48 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=8.05
+ $Y2=0
r114 45 46 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r115 43 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r116 43 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r117 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r118 40 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.61
+ $Y2=0
r119 40 42 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.695 $Y=0
+ $X2=3.45 $Y2=0
r120 38 53 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r121 36 42 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.465 $Y=0 $X2=3.45
+ $Y2=0
r122 36 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.465 $Y=0 $X2=3.55
+ $Y2=0
r123 35 45 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.635 $Y=0
+ $X2=3.91 $Y2=0
r124 35 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.55
+ $Y2=0
r125 31 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0
r126 31 33 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0.4
r127 27 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0
r128 27 29 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0.4
r129 26 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=0 $X2=1.67
+ $Y2=0
r130 25 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=0 $X2=2.61
+ $Y2=0
r131 25 26 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.525 $Y=0
+ $X2=1.755 $Y2=0
r132 21 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0
r133 21 23 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0.4
r134 20 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.73
+ $Y2=0
r135 19 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=0 $X2=1.67
+ $Y2=0
r136 19 20 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.585 $Y=0
+ $X2=0.815 $Y2=0
r137 15 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r138 15 17 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.4
r139 4 33 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.4
r140 3 29 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.4
r141 2 23 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.4
r142 1 17 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.4
.ends

