* File: sky130_fd_sc_hdll__a21o_2.pex.spice
* Created: Wed Sep  2 08:17:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A21O_2%A_80_21# 1 2 7 9 11 12 14 15 17 19 20 22 23
+ 27 29 30 31 32 37 40
c73 11 0 8.49032e-20 $X=0.5 $Y=1.31
r74 35 37 13.7177 $w=1.88e-07 $l=2.35e-07 $layer=LI1_cond $X=2.145 $Y=0.655
+ $X2=2.145 $Y2=0.42
r75 31 40 4.46303 $w=2.3e-07 $l=1.82e-07 $layer=LI1_cond $X=1.675 $Y=1.805
+ $X2=1.857 $Y2=1.805
r76 31 32 12.276 $w=2.28e-07 $l=2.45e-07 $layer=LI1_cond $X=1.675 $Y=1.805
+ $X2=1.43 $Y2=1.805
r77 29 35 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.05 $Y=0.74
+ $X2=2.145 $Y2=0.655
r78 29 30 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.05 $Y=0.74
+ $X2=1.43 $Y2=0.74
r79 28 41 16.2472 $w=2.67e-07 $l=9e-08 $layer=POLY_cond $X=1.072 $Y=1.16
+ $X2=1.072 $Y2=1.07
r80 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.08
+ $Y=1.16 $X2=1.08 $Y2=1.16
r81 25 32 7.69484 $w=2.3e-07 $l=2.69433e-07 $layer=LI1_cond $X=1.212 $Y=1.69
+ $X2=1.43 $Y2=1.805
r82 25 27 14.0413 $w=4.33e-07 $l=5.3e-07 $layer=LI1_cond $X=1.212 $Y=1.69
+ $X2=1.212 $Y2=1.16
r83 24 30 8.67519 $w=1.7e-07 $l=2.5701e-07 $layer=LI1_cond $X=1.212 $Y=0.825
+ $X2=1.43 $Y2=0.74
r84 24 27 8.87514 $w=4.33e-07 $l=3.35e-07 $layer=LI1_cond $X=1.212 $Y=0.825
+ $X2=1.212 $Y2=1.16
r85 20 41 22.72 $w=2.67e-07 $l=8.30662e-08 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=1.072 $Y2=1.07
r86 20 22 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=1.055 $Y2=0.56
r87 17 28 50.2707 $w=2.67e-07 $l=2.70185e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.072 $Y2=1.16
r88 17 19 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.03 $Y2=1.985
r89 16 23 7.5188 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=0.6 $Y=1.07 $X2=0.5
+ $Y2=1.07
r90 15 41 16.2448 $w=1.5e-07 $l=1.42e-07 $layer=POLY_cond $X=0.93 $Y=1.07
+ $X2=1.072 $Y2=1.07
r91 15 16 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.93 $Y=1.07 $X2=0.6
+ $Y2=1.07
r92 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.985
r93 11 12 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.5 $Y=1.31 $X2=0.5
+ $Y2=1.41
r94 10 23 17.9196 $w=1.75e-07 $l=7.5e-08 $layer=POLY_cond $X=0.5 $Y=1.145
+ $X2=0.5 $Y2=1.07
r95 10 11 54.7102 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.145 $X2=0.5
+ $Y2=1.31
r96 7 23 17.9196 $w=1.75e-07 $l=8.66025e-08 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.5 $Y2=1.07
r97 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=0.56
r98 2 40 300 $w=1.7e-07 $l=4.53211e-07 $layer=licon1_PDIFF $count=2 $X=1.715
+ $Y=1.485 $X2=1.84 $Y2=1.88
r99 1 37 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.02
+ $Y=0.235 $X2=2.155 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_2%B1 1 3 4 6 7
r27 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.055
+ $Y=1.16 $X2=2.055 $Y2=1.16
r28 4 10 46.5183 $w=3.27e-07 $l=2.87228e-07 $layer=POLY_cond $X=2.13 $Y=1.41
+ $X2=2.05 $Y2=1.16
r29 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.13 $Y=1.41 $X2=2.13
+ $Y2=1.985
r30 1 10 38.5818 $w=3.27e-07 $l=2.11069e-07 $layer=POLY_cond $X=1.945 $Y=0.995
+ $X2=2.05 $Y2=1.16
r31 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.945 $Y=0.995
+ $X2=1.945 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_2%A1 1 3 4 6 7 8
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.645
+ $Y=1.16 $X2=2.645 $Y2=1.16
r37 8 13 11.1643 $w=3.18e-07 $l=3.1e-07 $layer=LI1_cond $X=2.57 $Y=0.85 $X2=2.57
+ $Y2=1.16
r38 7 8 12.2447 $w=3.18e-07 $l=3.4e-07 $layer=LI1_cond $X=2.57 $Y=0.51 $X2=2.57
+ $Y2=0.85
r39 4 12 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.61 $Y=1.41
+ $X2=2.645 $Y2=1.16
r40 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.61 $Y=1.41 $X2=2.61
+ $Y2=1.985
r41 1 12 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.585 $Y=0.995
+ $X2=2.645 $Y2=1.16
r42 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.585 $Y=0.995
+ $X2=2.585 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_2%A2 1 3 4 6 7 15
r26 11 15 2.49616 $w=5.73e-07 $l=1.2e-07 $layer=LI1_cond $X=3.245 $Y=1.037
+ $X2=3.365 $Y2=1.037
r27 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.245
+ $Y=1.16 $X2=3.245 $Y2=1.16
r28 7 15 0.624041 $w=5.73e-07 $l=3e-08 $layer=LI1_cond $X=3.395 $Y=1.037
+ $X2=3.365 $Y2=1.037
r29 4 10 46.6797 $w=3.23e-07 $l=2.8592e-07 $layer=POLY_cond $X=3.125 $Y=1.41
+ $X2=3.202 $Y2=1.16
r30 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.125 $Y=1.41
+ $X2=3.125 $Y2=1.985
r31 1 10 38.5615 $w=3.23e-07 $l=2.09893e-07 $layer=POLY_cond $X=3.1 $Y=0.995
+ $X2=3.202 $Y2=1.16
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.1 $Y=0.995 $X2=3.1
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_2%VPWR 1 2 3 10 12 16 19 20 21 23 36 37 43
r50 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r51 43 46 10.1844 $w=4.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.27 $Y=2.34
+ $X2=1.27 $Y2=2.72
r52 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r53 34 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r54 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r55 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r56 31 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r57 30 33 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r58 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r59 28 46 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=1.485 $Y=2.72
+ $X2=1.27 $Y2=2.72
r60 28 30 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.485 $Y=2.72
+ $X2=1.61 $Y2=2.72
r61 27 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r62 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r63 24 40 4.31056 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=2.72
+ $X2=0.187 $Y2=2.72
r64 24 26 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.375 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 23 46 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=1.055 $Y=2.72
+ $X2=1.27 $Y2=2.72
r66 23 26 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.055 $Y=2.72
+ $X2=0.69 $Y2=2.72
r67 21 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r68 21 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r69 19 33 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.705 $Y=2.72
+ $X2=2.53 $Y2=2.72
r70 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.705 $Y=2.72
+ $X2=2.87 $Y2=2.72
r71 18 36 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.035 $Y=2.72
+ $X2=3.45 $Y2=2.72
r72 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=2.72
+ $X2=2.87 $Y2=2.72
r73 14 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=2.635
+ $X2=2.87 $Y2=2.72
r74 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.87 $Y=2.635
+ $X2=2.87 $Y2=2.34
r75 10 40 3.04949 $w=2.8e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.235 $Y=2.635
+ $X2=0.187 $Y2=2.72
r76 10 12 32.5154 $w=2.78e-07 $l=7.9e-07 $layer=LI1_cond $X=0.235 $Y=2.635
+ $X2=0.235 $Y2=1.845
r77 3 16 600 $w=1.7e-07 $l=9.36149e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.485 $X2=2.87 $Y2=2.34
r78 2 43 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.485 $X2=1.27 $Y2=2.34
r79 1 12 300 $w=1.7e-07 $l=4.17852e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.845
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_2%X 1 2 7 10
r20 10 13 57.8279 $w=2.78e-07 $l=1.405e-06 $layer=LI1_cond $X=0.685 $Y=0.42
+ $X2=0.685 $Y2=1.825
r21 7 13 15.8461 $w=2.78e-07 $l=3.85e-07 $layer=LI1_cond $X=0.685 $Y=2.21
+ $X2=0.685 $Y2=1.825
r22 2 13 300 $w=1.7e-07 $l=4.08167e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=1.485 $X2=0.74 $Y2=1.825
r23 1 10 182 $w=1.7e-07 $l=2.66927e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.74 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_2%A_444_297# 1 2 7 9 11 13 15
r16 13 20 3.77276 $w=2.2e-07 $l=1.33e-07 $layer=LI1_cond $X=3.365 $Y=1.935
+ $X2=3.365 $Y2=1.802
r17 13 15 19.1201 $w=2.18e-07 $l=3.65e-07 $layer=LI1_cond $X=3.365 $Y=1.935
+ $X2=3.365 $Y2=2.3
r18 12 18 3.15837 $w=2.65e-07 $l=1.13e-07 $layer=LI1_cond $X=2.485 $Y=1.802
+ $X2=2.372 $Y2=1.802
r19 11 20 3.12033 $w=2.65e-07 $l=1.1e-07 $layer=LI1_cond $X=3.255 $Y=1.802
+ $X2=3.365 $Y2=1.802
r20 11 12 33.4861 $w=2.63e-07 $l=7.7e-07 $layer=LI1_cond $X=3.255 $Y=1.802
+ $X2=2.485 $Y2=1.802
r21 7 18 3.71737 $w=2.25e-07 $l=1.33e-07 $layer=LI1_cond $X=2.372 $Y=1.935
+ $X2=2.372 $Y2=1.802
r22 7 9 18.6952 $w=2.23e-07 $l=3.65e-07 $layer=LI1_cond $X=2.372 $Y=1.935
+ $X2=2.372 $Y2=2.3
r23 2 20 600 $w=1.7e-07 $l=4.31451e-07 $layer=licon1_PDIFF $count=1 $X=3.215
+ $Y=1.485 $X2=3.36 $Y2=1.85
r24 2 15 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.215
+ $Y=1.485 $X2=3.36 $Y2=2.3
r25 1 18 600 $w=1.7e-07 $l=4.33561e-07 $layer=licon1_PDIFF $count=1 $X=2.22
+ $Y=1.485 $X2=2.37 $Y2=1.85
r26 1 9 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=2.22
+ $Y=1.485 $X2=2.37 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_2%VGND 1 2 3 10 12 14 16 18 20 25 35 42
r47 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r48 35 38 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=1.465 $Y=0 $X2=1.465
+ $Y2=0.36
r49 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r50 29 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r51 29 36 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.99 $Y=0 $X2=1.61
+ $Y2=0
r52 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r53 26 35 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.655 $Y=0 $X2=1.465
+ $Y2=0
r54 26 28 87.0963 $w=1.68e-07 $l=1.335e-06 $layer=LI1_cond $X=1.655 $Y=0
+ $X2=2.99 $Y2=0
r55 25 41 5.12538 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=3.155 $Y=0 $X2=3.417
+ $Y2=0
r56 25 28 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=0 $X2=2.99
+ $Y2=0
r57 24 36 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r58 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r59 21 31 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r60 21 23 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=1.15
+ $Y2=0
r61 20 35 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.275 $Y=0 $X2=1.465
+ $Y2=0
r62 20 23 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.275 $Y=0 $X2=1.15
+ $Y2=0
r63 18 24 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r64 18 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r65 14 41 3.07131 $w=3.8e-07 $l=1.15521e-07 $layer=LI1_cond $X=3.345 $Y=0.085
+ $X2=3.417 $Y2=0
r66 14 16 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=3.345 $Y=0.085
+ $X2=3.345 $Y2=0.38
r67 10 31 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r68 10 12 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r69 3 16 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.175
+ $Y=0.235 $X2=3.36 $Y2=0.38
r70 2 38 182 $w=1.7e-07 $l=4.17852e-07 $layer=licon1_NDIFF $count=1 $X=1.13
+ $Y=0.235 $X2=1.49 $Y2=0.36
r71 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

