* File: sky130_fd_sc_hdll__clkmux2_4.spice
* Created: Wed Sep  2 08:27:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__clkmux2_4.pex.spice"
.subckt sky130_fd_sc_hdll__clkmux2_4  VNB VPB S A1 A0 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A0	A0
* A1	A1
* S	S
* VPB	VPB
* VNB	VNB
MM1003 N_X_M1003_d N_A_79_199#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75004.3 A=0.078 P=1.34 MULT=1
MM1008 N_X_M1003_d N_A_79_199#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0962 PD=0.79 PS=0.89 NRD=0 NRS=8.076 M=1 R=3.46667 SA=75000.6
+ SB=75003.9 A=0.078 P=1.34 MULT=1
MM1011 N_X_M1011_d N_A_79_199#_M1011_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0962 PD=0.79 PS=0.89 NRD=0 NRS=12.684 M=1 R=3.46667 SA=75001.1
+ SB=75003.4 A=0.078 P=1.34 MULT=1
MM1014 N_X_M1011_d N_A_79_199#_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.139183 PD=0.79 PS=1.1617 NRD=0 NRS=5.76 M=1 R=3.46667
+ SA=75001.5 SB=75003 A=0.078 P=1.34 MULT=1
MM1016 A_525_47# N_S_M1016_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.42 AD=0.0714
+ AS=0.112417 PD=0.76 PS=0.938298 NRD=32.856 NRS=64.284 M=1 R=2.8 SA=75002.2
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1005 N_A_79_199#_M1005_d N_A1_M1005_g A_525_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.10605 AS=0.0714 PD=0.925 PS=0.76 NRD=45.708 NRS=32.856 M=1 R=2.8
+ SA=75002.7 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1009 A_754_47# N_A0_M1009_g N_A_79_199#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.17955 AS=0.10605 PD=1.275 PS=0.925 NRD=106.428 NRS=18.564 M=1 R=2.8
+ SA=75003.4 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_925_21#_M1001_g A_754_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0993702 AS=0.17955 PD=0.884681 PS=1.275 NRD=27.132 NRS=106.428 M=1 R=2.8
+ SA=75004.4 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1002 N_A_925_21#_M1002_d N_S_M1002_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.12303 PD=1.56 PS=1.09532 NRD=0 NRS=21.912 M=1 R=3.46667
+ SA=75004.1 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1000 N_VPWR_M1000_d N_A_79_199#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90004.8 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A_79_199#_M1004_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90004.3 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1004_d N_A_79_199#_M1010_g N_X_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90003.9 A=0.18 P=2.36 MULT=1
MM1015 N_VPWR_M1015_d N_A_79_199#_M1015_g N_X_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.222784 AS=0.145 PD=1.48454 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90003.4 A=0.18 P=2.36 MULT=1
MM1012 A_523_309# N_S_M1012_g N_VPWR_M1015_d VPB PHIGHVT L=0.18 W=0.94
+ AD=0.18565 AS=0.209416 PD=1.335 PS=1.39546 NRD=29.8455 NRS=32.4656 M=1
+ R=5.22222 SA=90002.2 SB=90003 A=0.1692 P=2.24 MULT=1
MM1013 N_A_79_199#_M1013_d N_A0_M1013_g A_523_309# VPB PHIGHVT L=0.18 W=0.94
+ AD=0.47235 AS=0.18565 PD=1.945 PS=1.335 NRD=1.0441 NRS=29.8455 M=1 R=5.22222
+ SA=90002.8 SB=90002.4 A=0.1692 P=2.24 MULT=1
MM1007 A_875_309# N_A1_M1007_g N_A_79_199#_M1013_d VPB PHIGHVT L=0.18 W=0.94
+ AD=0.1222 AS=0.47235 PD=1.2 PS=1.945 NRD=15.7009 NRS=1.0441 M=1 R=5.22222
+ SA=90004 SB=90001.2 A=0.1692 P=2.24 MULT=1
MM1017 N_VPWR_M1017_d N_A_925_21#_M1017_g A_875_309# VPB PHIGHVT L=0.18 W=0.94
+ AD=0.1833 AS=0.1222 PD=1.33 PS=1.2 NRD=19.897 NRS=15.7009 M=1 R=5.22222
+ SA=90004.4 SB=90000.8 A=0.1692 P=2.24 MULT=1
MM1006 N_A_925_21#_M1006_d N_S_M1006_g N_VPWR_M1017_d VPB PHIGHVT L=0.18 W=0.94
+ AD=0.2726 AS=0.1833 PD=2.46 PS=1.33 NRD=1.0441 NRS=3.1323 M=1 R=5.22222
+ SA=90005 SB=90000.2 A=0.1692 P=2.24 MULT=1
DX18_noxref VNB VPB NWDIODE A=10.2078 P=15.93
c_47 VNB 0 1.9931e-19 $X=1.8 $Y=-0.085
*
.include "sky130_fd_sc_hdll__clkmux2_4.pxi.spice"
*
.ends
*
*
