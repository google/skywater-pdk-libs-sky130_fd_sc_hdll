* File: sky130_fd_sc_hdll__nand4_1.spice
* Created: Wed Sep  2 08:38:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nand4_1.pex.spice"
.subckt sky130_fd_sc_hdll__nand4_1  VNB VPB D C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1006 A_119_47# N_D_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.2015 PD=0.97 PS=1.92 NRD=19.38 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1001 A_213_47# N_C_M1001_g A_119_47# VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.104 PD=0.92 PS=0.97 NRD=14.76 NRS=19.38 M=1 R=4.33333 SA=75000.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1003 A_297_47# N_B_M1003_g A_213_47# VNB NSHORT L=0.15 W=0.65 AD=0.1235
+ AS=0.08775 PD=1.03 PS=0.92 NRD=24.912 NRS=14.76 M=1 R=4.33333 SA=75001.1
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g A_297_47# VNB NSHORT L=0.15 W=0.65 AD=0.2275
+ AS=0.1235 PD=2 PS=1.03 NRD=8.304 NRS=24.912 M=1 R=4.33333 SA=75001.7
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_D_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_C_M1000_g N_Y_M1004_d VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.6
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1007 N_Y_M1007_d N_B_M1007_g N_VPWR_M1000_d VPB PHIGHVT L=0.18 W=1 AD=0.175
+ AS=0.145 PD=1.35 PS=1.29 NRD=6.8753 NRS=0.9653 M=1 R=5.55556 SA=90001.1
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g N_Y_M1007_d VPB PHIGHVT L=0.18 W=1 AD=0.31
+ AS=0.175 PD=2.62 PS=1.35 NRD=0.9653 NRS=6.8753 M=1 R=5.55556 SA=90001.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
pX9_noxref noxref_13 B B PROBETYPE=1
c_293 A_297_47# 0 1.19981e-19 $X=1.485 $Y=0.235
*
.include "sky130_fd_sc_hdll__nand4_1.pxi.spice"
*
.ends
*
*
