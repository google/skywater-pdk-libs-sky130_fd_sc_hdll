* File: sky130_fd_sc_hdll__clkinvlp_4.spice
* Created: Thu Aug 27 19:03:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__clkinvlp_4.pex.spice"
.subckt sky130_fd_sc_hdll__clkinvlp_4  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_M1003_g A_110_47# VNB NSHORT L=0.15 W=0.55 AD=0.14575
+ AS=0.05775 PD=1.63 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75000.2
+ SB=75001.3 A=0.0825 P=1.4 MULT=1
MM1001 A_110_47# N_A_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75000.5 SB=75001
+ A=0.0825 P=1.4 MULT=1
MM1005 A_268_47# N_A_M1005_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75001 SB=75000.5
+ A=0.0825 P=1.4 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g A_268_47# VNB NSHORT L=0.15 W=0.55 AD=0.143
+ AS=0.05775 PD=1.62 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75001.3
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.25 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002 A=0.25 P=2.5
+ MULT=1
MM1002 N_Y_M1000_d N_A_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.25 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25 P=2.5
+ MULT=1
MM1006 N_Y_M1006_d N_A_M1006_g N_VPWR_M1002_s VPB PHIGHVT L=0.25 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25 P=2.5
+ MULT=1
MM1007 N_Y_M1006_d N_A_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.25 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125000 A=0.25 P=2.5
+ MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hdll__clkinvlp_4.pxi.spice"
*
.ends
*
*
