* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__xor2_4 A B VGND VNB VPB VPWR X
X0 a_886_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_886_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_886_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_886_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 X B a_886_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_886_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_886_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 a_886_47# B X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 X B a_886_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR A a_886_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 VPWR B a_886_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 X a_112_47# a_886_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 VPWR A a_886_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_886_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 VGND A a_886_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 VGND A a_886_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X32 a_886_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 X a_112_47# a_886_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X35 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X36 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 a_886_47# B X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X38 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X39 VPWR B a_886_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
