* File: sky130_fd_sc_hdll__nor4b_4.pex.spice
* Created: Wed Sep  2 08:41:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR4B_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39 44
r75 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=1.93 $Y2=1.202
r76 37 39 22.6747 $w=3.72e-07 $l=1.75e-07 $layer=POLY_cond $X=1.73 $Y=1.202
+ $X2=1.905 $Y2=1.202
r77 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.73
+ $Y=1.16 $X2=1.73 $Y2=1.16
r78 35 37 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.73 $Y2=1.202
r79 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.202
+ $X2=1.435 $Y2=1.202
r80 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=1.41 $Y2=1.202
r81 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.202
+ $X2=0.965 $Y2=1.202
r82 31 44 30.368 $w=2.08e-07 $l=5.75e-07 $layer=LI1_cond $X=0.56 $Y=1.18
+ $X2=1.135 $Y2=1.18
r83 30 32 49.2366 $w=3.72e-07 $l=3.8e-07 $layer=POLY_cond $X=0.56 $Y=1.202
+ $X2=0.94 $Y2=1.202
r84 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.56
+ $Y=1.16 $X2=0.56 $Y2=1.16
r85 28 30 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.56 $Y2=1.202
r86 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r87 25 38 26.1429 $w=2.08e-07 $l=4.95e-07 $layer=LI1_cond $X=1.235 $Y=1.18
+ $X2=1.73 $Y2=1.18
r88 25 44 5.28139 $w=2.08e-07 $l=1e-07 $layer=LI1_cond $X=1.235 $Y=1.18
+ $X2=1.135 $Y2=1.18
r89 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r90 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r91 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r92 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r93 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r94 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r95 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.202
r96 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=0.56
r97 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r98 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r99 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=1.202
r100 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=0.56
r101 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r102 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r103 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.202
r104 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_4%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39 44
r77 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.785 $Y=1.202
+ $X2=3.81 $Y2=1.202
r78 37 39 22.6747 $w=3.72e-07 $l=1.75e-07 $layer=POLY_cond $X=3.61 $Y=1.202
+ $X2=3.785 $Y2=1.202
r79 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.61
+ $Y=1.16 $X2=3.61 $Y2=1.16
r80 35 37 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=3.315 $Y=1.202
+ $X2=3.61 $Y2=1.202
r81 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.202
+ $X2=3.315 $Y2=1.202
r82 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=3.29 $Y2=1.202
r83 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.845 $Y2=1.202
r84 31 44 28.2554 $w=2.08e-07 $l=5.35e-07 $layer=LI1_cond $X=2.44 $Y=1.18
+ $X2=2.975 $Y2=1.18
r85 30 32 49.2366 $w=3.72e-07 $l=3.8e-07 $layer=POLY_cond $X=2.44 $Y=1.202
+ $X2=2.82 $Y2=1.202
r86 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.44
+ $Y=1.16 $X2=2.44 $Y2=1.16
r87 28 30 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.44 $Y2=1.202
r88 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.202
+ $X2=2.375 $Y2=1.202
r89 25 38 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=3.275 $Y=1.18
+ $X2=3.61 $Y2=1.18
r90 25 44 15.8442 $w=2.08e-07 $l=3e-07 $layer=LI1_cond $X=3.275 $Y=1.18
+ $X2=2.975 $Y2=1.18
r91 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=1.202
r92 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=0.56
r93 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.202
r94 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r95 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.202
r96 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r97 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=1.202
r98 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=0.56
r99 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r100 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r101 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=1.202
r102 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=0.56
r103 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r104 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r105 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.202
r106 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_4%C 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39 45
r78 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.185 $Y=1.202
+ $X2=6.21 $Y2=1.202
r79 38 45 38.026 $w=2.08e-07 $l=7.2e-07 $layer=LI1_cond $X=6.01 $Y=1.18 $X2=5.29
+ $Y2=1.18
r80 37 39 22.6747 $w=3.72e-07 $l=1.75e-07 $layer=POLY_cond $X=6.01 $Y=1.202
+ $X2=6.185 $Y2=1.202
r81 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.01
+ $Y=1.16 $X2=6.01 $Y2=1.16
r82 35 37 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=5.715 $Y=1.202
+ $X2=6.01 $Y2=1.202
r83 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.69 $Y=1.202
+ $X2=5.715 $Y2=1.202
r84 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=5.245 $Y=1.202
+ $X2=5.69 $Y2=1.202
r85 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.22 $Y=1.202
+ $X2=5.245 $Y2=1.202
r86 30 32 49.2366 $w=3.72e-07 $l=3.8e-07 $layer=POLY_cond $X=4.84 $Y=1.202
+ $X2=5.22 $Y2=1.202
r87 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.84
+ $Y=1.16 $X2=4.84 $Y2=1.16
r88 28 30 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=4.775 $Y=1.202
+ $X2=4.84 $Y2=1.202
r89 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.75 $Y=1.202
+ $X2=4.775 $Y2=1.202
r90 25 45 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=5.285 $Y=1.18
+ $X2=5.29 $Y2=1.18
r91 25 31 23.5022 $w=2.08e-07 $l=4.45e-07 $layer=LI1_cond $X=5.285 $Y=1.18
+ $X2=4.84 $Y2=1.18
r92 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.21 $Y=0.995
+ $X2=6.21 $Y2=1.202
r93 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.21 $Y=0.995
+ $X2=6.21 $Y2=0.56
r94 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.202
r95 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.985
r96 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.202
r97 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.985
r98 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=1.202
r99 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=0.56
r100 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.202
r101 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.985
r102 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.22 $Y=0.995
+ $X2=5.22 $Y2=1.202
r103 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.22 $Y=0.995
+ $X2=5.22 $Y2=0.56
r104 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.202
r105 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
r106 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.75 $Y=0.995
+ $X2=4.75 $Y2=1.202
r107 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.75 $Y=0.995
+ $X2=4.75 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_4%A_1311_21# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 31 37 39 40 41 42 44 48 57 58 59
r118 69 70 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.04 $Y=1.202
+ $X2=8.065 $Y2=1.202
r119 66 67 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.57 $Y=1.202
+ $X2=7.595 $Y2=1.202
r120 65 66 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=7.125 $Y=1.202
+ $X2=7.57 $Y2=1.202
r121 64 65 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.1 $Y=1.202
+ $X2=7.125 $Y2=1.202
r122 63 64 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=6.655 $Y=1.202
+ $X2=7.1 $Y2=1.202
r123 62 63 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.63 $Y=1.202
+ $X2=6.655 $Y2=1.202
r124 59 70 13.6879 $w=3.72e-07 $l=1.19164e-07 $layer=POLY_cond $X=8.165 $Y=1.16
+ $X2=8.065 $Y2=1.202
r125 58 59 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=8.355 $Y=1.16
+ $X2=8.165 $Y2=1.16
r126 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.355
+ $Y=1.16 $X2=8.355 $Y2=1.16
r127 48 50 23.3929 $w=3.33e-07 $l=6.8e-07 $layer=LI1_cond $X=8.817 $Y=1.63
+ $X2=8.817 $Y2=2.31
r128 46 48 0.172006 $w=3.33e-07 $l=5e-09 $layer=LI1_cond $X=8.817 $Y=1.625
+ $X2=8.817 $Y2=1.63
r129 42 52 28.8364 $w=1.68e-07 $l=4.42e-07 $layer=LI1_cond $X=8.797 $Y=0.82
+ $X2=8.355 $Y2=0.82
r130 42 44 10.6025 $w=3.73e-07 $l=3.45e-07 $layer=LI1_cond $X=8.797 $Y=0.735
+ $X2=8.797 $Y2=0.39
r131 40 46 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=8.65 $Y=1.54
+ $X2=8.817 $Y2=1.625
r132 40 41 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=8.65 $Y=1.54
+ $X2=8.44 $Y2=1.54
r133 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.355 $Y=1.455
+ $X2=8.44 $Y2=1.54
r134 38 57 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=8.355 $Y=1.285
+ $X2=8.355 $Y2=1.18
r135 38 39 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.355 $Y=1.285
+ $X2=8.355 $Y2=1.455
r136 37 57 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=8.355 $Y=1.075
+ $X2=8.355 $Y2=1.18
r137 36 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.355 $Y=0.905
+ $X2=8.355 $Y2=0.82
r138 36 37 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.355 $Y=0.905
+ $X2=8.355 $Y2=1.075
r139 34 69 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.015 $Y=1.202
+ $X2=8.04 $Y2=1.202
r140 34 67 54.4194 $w=3.72e-07 $l=4.2e-07 $layer=POLY_cond $X=8.015 $Y=1.202
+ $X2=7.595 $Y2=1.202
r141 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.015
+ $Y=1.16 $X2=8.015 $Y2=1.16
r142 31 57 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=8.27 $Y=1.18
+ $X2=8.355 $Y2=1.18
r143 31 33 13.4675 $w=2.08e-07 $l=2.55e-07 $layer=LI1_cond $X=8.27 $Y=1.18
+ $X2=8.015 $Y2=1.18
r144 28 70 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.065 $Y=1.41
+ $X2=8.065 $Y2=1.202
r145 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.065 $Y=1.41
+ $X2=8.065 $Y2=1.985
r146 25 69 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.04 $Y=0.995
+ $X2=8.04 $Y2=1.202
r147 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.04 $Y=0.995
+ $X2=8.04 $Y2=0.56
r148 22 67 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.595 $Y=1.41
+ $X2=7.595 $Y2=1.202
r149 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.595 $Y=1.41
+ $X2=7.595 $Y2=1.985
r150 19 66 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.57 $Y=0.995
+ $X2=7.57 $Y2=1.202
r151 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.57 $Y=0.995
+ $X2=7.57 $Y2=0.56
r152 16 65 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.202
r153 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.985
r154 13 64 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.1 $Y=0.995
+ $X2=7.1 $Y2=1.202
r155 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.1 $Y=0.995
+ $X2=7.1 $Y2=0.56
r156 10 63 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.202
r157 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.985
r158 7 62 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=1.202
r159 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=0.56
r160 2 50 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=8.695
+ $Y=1.485 $X2=8.82 $Y2=2.31
r161 2 48 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=8.695
+ $Y=1.485 $X2=8.82 $Y2=1.63
r162 1 44 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=8.695
+ $Y=0.235 $X2=8.82 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_4%D_N 1 3 4 6 7 14
r27 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.245
+ $Y=1.16 $X2=9.245 $Y2=1.16
r28 7 14 6.33766 $w=2.08e-07 $l=1.2e-07 $layer=LI1_cond $X=9.365 $Y=1.18
+ $X2=9.245 $Y2=1.18
r29 4 10 44.8713 $w=4.02e-07 $l=3.07002e-07 $layer=POLY_cond $X=9.055 $Y=1.41
+ $X2=9.182 $Y2=1.16
r30 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.055 $Y=1.41
+ $X2=9.055 $Y2=1.985
r31 1 10 39.6247 $w=4.02e-07 $l=2.28703e-07 $layer=POLY_cond $X=9.03 $Y=0.995
+ $X2=9.182 $Y2=1.16
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.03 $Y=0.995 $X2=9.03
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_4%A_27_297# 1 2 3 4 5 18 22 23 26 28 30 31
+ 32 36 38 42 45 50
r66 40 42 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.02 $Y=2.295
+ $X2=4.02 $Y2=1.96
r67 39 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.205 $Y=2.38
+ $X2=3.08 $Y2=2.38
r68 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.895 $Y=2.38
+ $X2=4.02 $Y2=2.295
r69 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.895 $Y=2.38
+ $X2=3.205 $Y2=2.38
r70 34 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.295
+ $X2=3.08 $Y2=2.38
r71 34 36 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.08 $Y=2.295
+ $X2=3.08 $Y2=1.96
r72 33 49 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.265 $Y=2.38
+ $X2=2.14 $Y2=2.38
r73 32 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.955 $Y=2.38
+ $X2=3.08 $Y2=2.38
r74 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.955 $Y=2.38
+ $X2=2.265 $Y2=2.38
r75 31 49 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.295
+ $X2=2.14 $Y2=2.38
r76 30 47 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=1.625
+ $X2=2.14 $Y2=1.54
r77 30 31 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=2.14 $Y=1.625
+ $X2=2.14 $Y2=2.295
r78 29 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.325 $Y=1.54
+ $X2=1.2 $Y2=1.54
r79 28 47 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.015 $Y=1.54
+ $X2=2.14 $Y2=1.54
r80 28 29 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.015 $Y=1.54
+ $X2=1.325 $Y2=1.54
r81 24 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=1.625
+ $X2=1.2 $Y2=1.54
r82 24 26 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.2 $Y=1.625 $X2=1.2
+ $Y2=2.3
r83 22 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.075 $Y=1.54
+ $X2=1.2 $Y2=1.54
r84 22 23 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.075 $Y=1.54
+ $X2=0.425 $Y2=1.54
r85 18 20 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.63
+ $X2=0.26 $Y2=2.31
r86 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.425 $Y2=1.54
r87 16 18 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.26 $Y2=1.63
r88 5 42 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=1.96
r89 4 36 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=1.96
r90 3 49 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2.3
r91 3 47 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.62
r92 2 45 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.62
r93 2 26 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.3
r94 1 20 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.31
r95 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_4%VPWR 1 2 3 14 16 20 22 24 28 30 39 42 46
r104 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r105 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r106 40 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r107 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r108 37 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.43 $Y2=2.72
r109 36 37 1.1625 $w=1.7e-07 $l=1.36e-06 $layer=mcon $count=8 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r110 34 37 1.96334 $w=4.8e-07 $l=6.9e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=8.97 $Y2=2.72
r111 34 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r112 33 36 450.16 $w=1.68e-07 $l=6.9e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=8.97 $Y2=2.72
r113 33 34 1.1625 $w=1.7e-07 $l=1.36e-06 $layer=mcon $count=8 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r114 31 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.795 $Y=2.72
+ $X2=1.67 $Y2=2.72
r115 31 33 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.795 $Y=2.72
+ $X2=2.07 $Y2=2.72
r116 30 45 3.75722 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=9.205 $Y=2.72
+ $X2=9.432 $Y2=2.72
r117 30 36 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.205 $Y=2.72
+ $X2=8.97 $Y2=2.72
r118 28 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r119 24 27 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.32 $Y=1.63
+ $X2=9.32 $Y2=2.31
r120 22 45 3.26067 $w=2.3e-07 $l=1.4854e-07 $layer=LI1_cond $X=9.32 $Y=2.635
+ $X2=9.432 $Y2=2.72
r121 22 27 16.2845 $w=2.28e-07 $l=3.25e-07 $layer=LI1_cond $X=9.32 $Y=2.635
+ $X2=9.32 $Y2=2.31
r122 18 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.72
r123 18 20 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=1.96
r124 17 39 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=0.75 $Y2=2.72
r125 16 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.545 $Y=2.72
+ $X2=1.67 $Y2=2.72
r126 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.545 $Y=2.72
+ $X2=0.855 $Y2=2.72
r127 12 39 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r128 12 14 35.6493 $w=2.08e-07 $l=6.75e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=1.96
r129 3 27 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=9.145
+ $Y=1.485 $X2=9.29 $Y2=2.31
r130 3 24 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=9.145
+ $Y=1.485 $X2=9.29 $Y2=1.63
r131 2 20 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.96
r132 1 14 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_4%A_493_297# 1 2 3 4 15 19 23 28 30 32 34
r60 24 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.135 $Y=1.54
+ $X2=5.01 $Y2=1.54
r61 23 34 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.825 $Y=1.54
+ $X2=5.95 $Y2=1.54
r62 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.825 $Y=1.54
+ $X2=5.135 $Y2=1.54
r63 20 30 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.675 $Y=1.54
+ $X2=3.55 $Y2=1.54
r64 19 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.885 $Y=1.54
+ $X2=5.01 $Y2=1.54
r65 19 20 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=4.885 $Y=1.54
+ $X2=3.675 $Y2=1.54
r66 16 28 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.735 $Y=1.54
+ $X2=2.61 $Y2=1.54
r67 15 30 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.425 $Y=1.54
+ $X2=3.55 $Y2=1.54
r68 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.425 $Y=1.54
+ $X2=2.735 $Y2=1.54
r69 4 34 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=1.62
r70 3 32 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=1.62
r71 2 30 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.62
r72 1 28 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_4%A_883_297# 1 2 3 4 5 18 20 21 24 26 30 32
+ 36 38 42 44 46 47
r65 40 42 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=8.3 $Y=2.295
+ $X2=8.3 $Y2=1.96
r66 39 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.485 $Y=2.38
+ $X2=7.36 $Y2=2.38
r67 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.175 $Y=2.38
+ $X2=8.3 $Y2=2.295
r68 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.175 $Y=2.38
+ $X2=7.485 $Y2=2.38
r69 34 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=2.295
+ $X2=7.36 $Y2=2.38
r70 34 36 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=7.36 $Y=2.295
+ $X2=7.36 $Y2=1.96
r71 33 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.545 $Y=2.38
+ $X2=6.42 $Y2=2.38
r72 32 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.235 $Y=2.38
+ $X2=7.36 $Y2=2.38
r73 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.235 $Y=2.38
+ $X2=6.545 $Y2=2.38
r74 28 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=2.295
+ $X2=6.42 $Y2=2.38
r75 28 30 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=6.42 $Y=2.295
+ $X2=6.42 $Y2=1.62
r76 27 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.605 $Y=2.38
+ $X2=5.48 $Y2=2.38
r77 26 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.295 $Y=2.38
+ $X2=6.42 $Y2=2.38
r78 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.295 $Y=2.38
+ $X2=5.605 $Y2=2.38
r79 22 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=2.295
+ $X2=5.48 $Y2=2.38
r80 22 24 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.48 $Y=2.295
+ $X2=5.48 $Y2=1.96
r81 20 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.355 $Y=2.38
+ $X2=5.48 $Y2=2.38
r82 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.355 $Y=2.38
+ $X2=4.665 $Y2=2.38
r83 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.54 $Y=2.295
+ $X2=4.665 $Y2=2.38
r84 16 18 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.54 $Y=2.295
+ $X2=4.54 $Y2=1.96
r85 5 42 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=8.155
+ $Y=1.485 $X2=8.3 $Y2=1.96
r86 4 36 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=7.215
+ $Y=1.485 $X2=7.36 $Y2=1.96
r87 3 46 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=6.275
+ $Y=1.485 $X2=6.42 $Y2=2.3
r88 3 30 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.275
+ $Y=1.485 $X2=6.42 $Y2=1.62
r89 2 24 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=1.96
r90 1 18 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=4.415
+ $Y=1.485 $X2=4.54 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_4%Y 1 2 3 4 5 6 7 8 9 10 33 35 36 39 41 45
+ 47 51 53 57 59 63 65 69 72 73 75 79 83 84 85 86 87 88 91 93 94
c196 91 0 1.85425e-19 $X=6.89 $Y=1.62
r197 89 94 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=6.89 $Y=1.625
+ $X2=6.89 $Y2=1.87
r198 89 91 2.61584 $w=3.67e-07 $l=1.53734e-07 $layer=LI1_cond $X=6.89 $Y=1.625
+ $X2=7.007 $Y2=1.54
r199 77 79 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.805 $Y=0.725
+ $X2=7.805 $Y2=0.39
r200 76 91 4.2195 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=7.25 $Y=1.54
+ $X2=7.007 $Y2=1.54
r201 75 93 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.705 $Y=1.54
+ $X2=7.83 $Y2=1.54
r202 75 76 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=7.705 $Y=1.54
+ $X2=7.25 $Y2=1.54
r203 74 88 6.0485 $w=1.8e-07 $l=2.88e-07 $layer=LI1_cond $X=7.25 $Y=0.815
+ $X2=6.962 $Y2=0.815
r204 73 77 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=7.615 $Y=0.815
+ $X2=7.805 $Y2=0.725
r205 73 74 22.4899 $w=1.78e-07 $l=3.65e-07 $layer=LI1_cond $X=7.615 $Y=0.815
+ $X2=7.25 $Y2=0.815
r206 72 91 2.61584 $w=3.67e-07 $l=8.5e-08 $layer=LI1_cond $X=7.007 $Y=1.455
+ $X2=7.007 $Y2=1.54
r207 71 88 0.865627 $w=4.85e-07 $l=1.10227e-07 $layer=LI1_cond $X=7.007 $Y=0.905
+ $X2=6.962 $Y2=0.815
r208 71 72 13.5638 $w=4.83e-07 $l=5.5e-07 $layer=LI1_cond $X=7.007 $Y=0.905
+ $X2=7.007 $Y2=1.455
r209 67 88 0.865627 $w=3.8e-07 $l=1.34681e-07 $layer=LI1_cond $X=6.865 $Y=0.725
+ $X2=6.962 $Y2=0.815
r210 67 69 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.865 $Y=0.725
+ $X2=6.865 $Y2=0.39
r211 66 87 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.115 $Y=0.815
+ $X2=5.925 $Y2=0.815
r212 65 88 6.0485 $w=1.8e-07 $l=2.87e-07 $layer=LI1_cond $X=6.675 $Y=0.815
+ $X2=6.962 $Y2=0.815
r213 65 66 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=6.675 $Y=0.815
+ $X2=6.115 $Y2=0.815
r214 61 87 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=5.925 $Y=0.725
+ $X2=5.925 $Y2=0.815
r215 61 63 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.925 $Y=0.725
+ $X2=5.925 $Y2=0.39
r216 60 86 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.175 $Y=0.815
+ $X2=4.985 $Y2=0.815
r217 59 87 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.735 $Y=0.815
+ $X2=5.925 $Y2=0.815
r218 59 60 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=5.735 $Y=0.815
+ $X2=5.175 $Y2=0.815
r219 55 86 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=4.985 $Y=0.725
+ $X2=4.985 $Y2=0.815
r220 55 57 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.985 $Y=0.725
+ $X2=4.985 $Y2=0.39
r221 54 85 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.715 $Y=0.815
+ $X2=3.525 $Y2=0.815
r222 53 86 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.795 $Y=0.815
+ $X2=4.985 $Y2=0.815
r223 53 54 66.5455 $w=1.78e-07 $l=1.08e-06 $layer=LI1_cond $X=4.795 $Y=0.815
+ $X2=3.715 $Y2=0.815
r224 49 85 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=3.525 $Y=0.725
+ $X2=3.525 $Y2=0.815
r225 49 51 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.525 $Y=0.725
+ $X2=3.525 $Y2=0.39
r226 48 84 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=0.815
+ $X2=2.585 $Y2=0.815
r227 47 85 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.335 $Y=0.815
+ $X2=3.525 $Y2=0.815
r228 47 48 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.335 $Y=0.815
+ $X2=2.775 $Y2=0.815
r229 43 84 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=2.585 $Y=0.725
+ $X2=2.585 $Y2=0.815
r230 43 45 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.585 $Y=0.725
+ $X2=2.585 $Y2=0.39
r231 42 83 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=0.815
+ $X2=1.645 $Y2=0.815
r232 41 84 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=0.815
+ $X2=2.585 $Y2=0.815
r233 41 42 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=2.395 $Y=0.815
+ $X2=1.835 $Y2=0.815
r234 37 83 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=1.645 $Y=0.725
+ $X2=1.645 $Y2=0.815
r235 37 39 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.645 $Y=0.725
+ $X2=1.645 $Y2=0.39
r236 35 83 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=0.815
+ $X2=1.645 $Y2=0.815
r237 35 36 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.455 $Y=0.815
+ $X2=0.895 $Y2=0.815
r238 31 36 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=0.705 $Y=0.725
+ $X2=0.895 $Y2=0.815
r239 31 33 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.705 $Y=0.725
+ $X2=0.705 $Y2=0.39
r240 10 93 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=7.685
+ $Y=1.485 $X2=7.83 $Y2=1.62
r241 9 91 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=1.62
r242 8 79 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=7.645
+ $Y=0.235 $X2=7.83 $Y2=0.39
r243 7 69 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=6.705
+ $Y=0.235 $X2=6.89 $Y2=0.39
r244 6 63 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=5.765
+ $Y=0.235 $X2=5.95 $Y2=0.39
r245 5 57 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.825
+ $Y=0.235 $X2=5.01 $Y2=0.39
r246 4 51 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.39
r247 3 45 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.39
r248 2 39 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.39
r249 1 33 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_4%VGND 1 2 3 4 5 6 7 8 9 10 31 33 35 39 41
+ 45 49 53 57 61 65 67 69 72 73 75 76 78 79 81 82 84 85 86 109 117 120 125 128
+ 131
r164 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r165 127 128 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=0.235
+ $X2=4.625 $Y2=0.235
r166 123 127 3.17708 $w=6.38e-07 $l=1.7e-07 $layer=LI1_cond $X=4.37 $Y=0.235
+ $X2=4.54 $Y2=0.235
r167 123 125 15.4628 $w=6.38e-07 $l=4.35e-07 $layer=LI1_cond $X=4.37 $Y=0.235
+ $X2=3.935 $Y2=0.235
r168 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r169 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r170 118 121 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.07 $Y2=0
r171 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r172 112 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.43 $Y2=0
r173 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r174 109 130 3.75722 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=9.205 $Y=0
+ $X2=9.432 $Y2=0
r175 109 111 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.205 $Y=0
+ $X2=8.97 $Y2=0
r176 108 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.97 $Y2=0
r177 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r178 105 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r179 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r180 102 105 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.13 $Y2=0
r181 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r182 99 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.21 $Y2=0
r183 99 124 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=4.37 $Y2=0
r184 98 128 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=5.29 $Y=0
+ $X2=4.625 $Y2=0
r185 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r186 95 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.37 $Y2=0
r187 94 125 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.91 $Y=0
+ $X2=3.935 $Y2=0
r188 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r189 91 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r190 91 121 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=2.07 $Y2=0
r191 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r192 88 120 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=0 $X2=2.14
+ $Y2=0
r193 88 90 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.225 $Y=0
+ $X2=2.99 $Y2=0
r194 86 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=1.15 $Y2=0
r195 86 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r196 84 107 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.215 $Y=0
+ $X2=8.05 $Y2=0
r197 84 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.215 $Y=0 $X2=8.3
+ $Y2=0
r198 83 111 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=8.385 $Y=0
+ $X2=8.97 $Y2=0
r199 83 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.385 $Y=0 $X2=8.3
+ $Y2=0
r200 81 104 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.275 $Y=0
+ $X2=7.13 $Y2=0
r201 81 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.275 $Y=0 $X2=7.36
+ $Y2=0
r202 80 107 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=7.445 $Y=0
+ $X2=8.05 $Y2=0
r203 80 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.445 $Y=0 $X2=7.36
+ $Y2=0
r204 78 101 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.335 $Y=0
+ $X2=6.21 $Y2=0
r205 78 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.335 $Y=0 $X2=6.42
+ $Y2=0
r206 77 104 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=6.505 $Y=0
+ $X2=7.13 $Y2=0
r207 77 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.505 $Y=0 $X2=6.42
+ $Y2=0
r208 75 98 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=5.395 $Y=0
+ $X2=5.29 $Y2=0
r209 75 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=0 $X2=5.48
+ $Y2=0
r210 74 101 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=5.565 $Y=0
+ $X2=6.21 $Y2=0
r211 74 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=0 $X2=5.48
+ $Y2=0
r212 72 90 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.995 $Y=0 $X2=2.99
+ $Y2=0
r213 72 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=0 $X2=3.08
+ $Y2=0
r214 71 94 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3.165 $Y=0
+ $X2=3.91 $Y2=0
r215 71 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=0 $X2=3.08
+ $Y2=0
r216 67 130 3.26067 $w=2.3e-07 $l=1.4854e-07 $layer=LI1_cond $X=9.32 $Y=0.085
+ $X2=9.432 $Y2=0
r217 67 69 15.2824 $w=2.28e-07 $l=3.05e-07 $layer=LI1_cond $X=9.32 $Y=0.085
+ $X2=9.32 $Y2=0.39
r218 63 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.3 $Y=0.085 $X2=8.3
+ $Y2=0
r219 63 65 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.3 $Y=0.085
+ $X2=8.3 $Y2=0.39
r220 59 82 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0
r221 59 61 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0.39
r222 55 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0
r223 55 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0.39
r224 51 76 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0
r225 51 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.39
r226 47 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0
r227 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.39
r228 43 120 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0
r229 43 45 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0.39
r230 42 117 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.2
+ $Y2=0
r231 41 120 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0 $X2=2.14
+ $Y2=0
r232 41 42 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=0
+ $X2=1.285 $Y2=0
r233 37 117 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0
r234 37 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0.39
r235 36 114 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r236 35 117 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.2
+ $Y2=0
r237 35 36 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=0.345 $Y2=0
r238 31 114 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r239 31 33 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.39
r240 10 69 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=9.105
+ $Y=0.235 $X2=9.29 $Y2=0.39
r241 9 65 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=8.115
+ $Y=0.235 $X2=8.3 $Y2=0.39
r242 8 61 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=7.175
+ $Y=0.235 $X2=7.36 $Y2=0.39
r243 7 57 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.285
+ $Y=0.235 $X2=6.42 $Y2=0.39
r244 6 53 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=5.295
+ $Y=0.235 $X2=5.48 $Y2=0.39
r245 5 127 91 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_NDIFF $count=2 $X=3.885
+ $Y=0.235 $X2=4.54 $Y2=0.39
r246 4 49 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.39
r247 3 45 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.39
r248 2 39 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.39
r249 1 33 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

