* File: sky130_fd_sc_hdll__o211a_1.spice
* Created: Wed Sep  2 08:42:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o211a_1.pex.spice"
.subckt sky130_fd_sc_hdll__o211a_1  VNB VPB A1 A2 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_79_21#_M1008_g N_X_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.169 PD=1.92 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A1_M1009_g N_A_225_47#_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.121875 AS=0.169 PD=1.025 PS=1.82 NRD=13.836 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1000 N_A_225_47#_M1000_d N_A2_M1000_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.15925 AS=0.121875 PD=1.14 PS=1.025 NRD=8.304 NRS=3.684 M=1 R=4.33333
+ SA=75000.7 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1003 A_540_47# N_B1_M1003_g N_A_225_47#_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.15925 PD=1.21 PS=1.14 NRD=41.532 NRS=30.456 M=1 R=4.33333
+ SA=75001.3 SB=75001 A=0.0975 P=1.6 MULT=1
MM1006 N_A_79_21#_M1006_d N_C1_M1006_g A_540_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.2275 AS=0.182 PD=2 PS=1.21 NRD=15.684 NRS=41.532 M=1 R=4.33333 SA=75002.1
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_A_79_21#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.27 PD=2.54 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1007 A_315_297# N_A1_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1 AD=0.1725
+ AS=0.27 PD=1.345 PS=2.54 NRD=23.1278 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90002.1 A=0.18 P=2.36 MULT=1
MM1005 N_A_79_21#_M1005_d N_A2_M1005_g A_315_297# VPB PHIGHVT L=0.18 W=1 AD=0.23
+ AS=0.1725 PD=1.46 PS=1.345 NRD=11.8003 NRS=23.1278 M=1 R=5.55556 SA=90000.7
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_B1_M1002_g N_A_79_21#_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.265 AS=0.23 PD=1.53 PS=1.46 NRD=8.8453 NRS=23.6203 M=1 R=5.55556
+ SA=90001.3 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1001 N_A_79_21#_M1001_d N_C1_M1001_g N_VPWR_M1002_d VPB PHIGHVT L=0.18 W=1
+ AD=0.31 AS=0.265 PD=2.62 PS=1.53 NRD=8.8453 NRS=40.3653 M=1 R=5.55556
+ SA=90002.1 SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hdll__o211a_1.pxi.spice"
*
.ends
*
*
