* File: sky130_fd_sc_hdll__einvn_2.pxi.spice
* Created: Thu Aug 27 19:07:28 2020
* 
x_PM_SKY130_FD_SC_HDLL__EINVN_2%TE_B N_TE_B_c_60_n N_TE_B_c_64_n N_TE_B_c_65_n
+ N_TE_B_M1001_g N_TE_B_M1004_g N_TE_B_c_66_n N_TE_B_c_67_n N_TE_B_M1000_g
+ N_TE_B_c_68_n N_TE_B_c_69_n N_TE_B_M1002_g N_TE_B_c_70_n TE_B
+ PM_SKY130_FD_SC_HDLL__EINVN_2%TE_B
x_PM_SKY130_FD_SC_HDLL__EINVN_2%A_27_47# N_A_27_47#_M1004_s N_A_27_47#_M1001_s
+ N_A_27_47#_c_109_n N_A_27_47#_M1005_g N_A_27_47#_c_110_n N_A_27_47#_c_111_n
+ N_A_27_47#_c_112_n N_A_27_47#_M1006_g N_A_27_47#_c_113_n N_A_27_47#_c_118_n
+ N_A_27_47#_c_114_n N_A_27_47#_c_115_n N_A_27_47#_c_116_n N_A_27_47#_c_117_n
+ PM_SKY130_FD_SC_HDLL__EINVN_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__EINVN_2%A N_A_M1003_g N_A_c_181_n N_A_M1007_g
+ N_A_c_178_n N_A_M1008_g N_A_c_182_n N_A_M1009_g A N_A_c_179_n A
+ PM_SKY130_FD_SC_HDLL__EINVN_2%A
x_PM_SKY130_FD_SC_HDLL__EINVN_2%VPWR N_VPWR_M1001_d N_VPWR_M1002_d
+ N_VPWR_c_225_n N_VPWR_c_226_n N_VPWR_c_227_n N_VPWR_c_228_n N_VPWR_c_229_n
+ VPWR N_VPWR_c_230_n N_VPWR_c_231_n N_VPWR_c_224_n N_VPWR_c_233_n
+ PM_SKY130_FD_SC_HDLL__EINVN_2%VPWR
x_PM_SKY130_FD_SC_HDLL__EINVN_2%A_222_309# N_A_222_309#_M1000_s
+ N_A_222_309#_M1007_s N_A_222_309#_c_281_n N_A_222_309#_c_279_n
+ N_A_222_309#_c_295_n N_A_222_309#_c_280_n
+ PM_SKY130_FD_SC_HDLL__EINVN_2%A_222_309#
x_PM_SKY130_FD_SC_HDLL__EINVN_2%Z N_Z_M1003_s N_Z_M1007_d N_Z_M1009_d Z Z Z Z Z
+ Z Z N_Z_c_325_n Z N_Z_c_322_n Z Z PM_SKY130_FD_SC_HDLL__EINVN_2%Z
x_PM_SKY130_FD_SC_HDLL__EINVN_2%VGND N_VGND_M1004_d N_VGND_M1005_s
+ N_VGND_c_363_n N_VGND_c_364_n N_VGND_c_365_n VGND N_VGND_c_366_n
+ N_VGND_c_367_n N_VGND_c_368_n N_VGND_c_369_n N_VGND_c_370_n
+ PM_SKY130_FD_SC_HDLL__EINVN_2%VGND
x_PM_SKY130_FD_SC_HDLL__EINVN_2%A_234_47# N_A_234_47#_M1005_d
+ N_A_234_47#_M1006_d N_A_234_47#_M1008_d N_A_234_47#_c_415_n
+ N_A_234_47#_c_423_n N_A_234_47#_c_411_n N_A_234_47#_c_447_n
+ N_A_234_47#_c_412_n N_A_234_47#_c_413_n
+ PM_SKY130_FD_SC_HDLL__EINVN_2%A_234_47#
cc_1 VNB N_TE_B_c_60_n 0.0430855f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.47
cc_2 VNB N_TE_B_M1004_g 0.0427154f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_3 VNB TE_B 0.0133203f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_27_47#_c_109_n 0.0176859f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_5 VNB N_A_27_47#_c_110_n 0.00920612f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=1.395
cc_6 VNB N_A_27_47#_c_111_n 0.00910466f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.395
cc_7 VNB N_A_27_47#_c_112_n 0.0151136f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=1.47
cc_8 VNB N_A_27_47#_c_113_n 0.0155207f $X=-0.19 $Y=-0.24 $X2=1.49 $Y2=1.47
cc_9 VNB N_A_27_47#_c_114_n 0.0011226f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_10 VNB N_A_27_47#_c_115_n 0.0193981f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_11 VNB N_A_27_47#_c_116_n 0.022058f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_117_n 0.0230217f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_M1003_g 0.0188584f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.77
cc_14 VNB N_A_c_178_n 0.0224229f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_15 VNB N_A_c_179_n 0.0626808f $X=-0.19 $Y=-0.24 $X2=1.49 $Y2=2.015
cc_16 VNB A 0.0159091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VPWR_c_224_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Z_c_322_n 0.00152249f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_363_n 0.00553967f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_364_n 0.0174316f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.395
cc_21 VNB N_VGND_c_365_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=1.4 $Y2=1.395
cc_22 VNB N_VGND_c_366_n 0.0143218f $X=-0.19 $Y=-0.24 $X2=1.49 $Y2=2.015
cc_23 VNB N_VGND_c_367_n 0.0432272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_368_n 0.214539f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_369_n 0.00573782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_370_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_234_47#_c_411_n 0.00772857f $X=-0.19 $Y=-0.24 $X2=1.49 $Y2=2.015
cc_28 VNB N_A_234_47#_c_412_n 0.0141396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_234_47#_c_413_n 0.0088592f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_30 VPB N_TE_B_c_60_n 0.0193621f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.47
cc_31 VPB N_TE_B_c_64_n 0.0145983f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.67
cc_32 VPB N_TE_B_c_65_n 0.0263165f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_33 VPB N_TE_B_c_66_n 0.0192593f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=1.395
cc_34 VPB N_TE_B_c_67_n 0.0161657f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.47
cc_35 VPB N_TE_B_c_68_n 0.0291206f $X=-0.19 $Y=1.305 $X2=1.4 $Y2=1.395
cc_36 VPB N_TE_B_c_69_n 0.0181916f $X=-0.19 $Y=1.305 $X2=1.49 $Y2=1.47
cc_37 VPB N_TE_B_c_70_n 0.00737735f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.395
cc_38 VPB TE_B 0.0054315f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_39 VPB N_A_27_47#_c_118_n 0.0305614f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_40 VPB N_A_27_47#_c_114_n 0.0140749f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_41 VPB N_A_27_47#_c_117_n 0.00992428f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_c_181_n 0.0184286f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.165
cc_43 VPB N_A_c_182_n 0.0200807f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.395
cc_44 VPB N_A_c_179_n 0.0226943f $X=-0.19 $Y=1.305 $X2=1.49 $Y2=2.015
cc_45 VPB N_VPWR_c_225_n 4.0558e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_226_n 0.00410146f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.395
cc_47 VPB N_VPWR_c_227_n 0.0134677f $X=-0.19 $Y=1.305 $X2=1.4 $Y2=1.395
cc_48 VPB N_VPWR_c_228_n 0.0158318f $X=-0.19 $Y=1.305 $X2=1.49 $Y2=1.47
cc_49 VPB N_VPWR_c_229_n 0.00476476f $X=-0.19 $Y=1.305 $X2=1.49 $Y2=2.015
cc_50 VPB N_VPWR_c_230_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_51 VPB N_VPWR_c_231_n 0.032042f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_224_n 0.0470377f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_233_n 0.00570037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_222_309#_c_279_n 0.00697965f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.395
cc_55 VPB N_A_222_309#_c_280_n 0.00996977f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.395
cc_56 VPB Z 0.016935f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=2.015
cc_57 VPB Z 0.0363333f $X=-0.19 $Y=1.305 $X2=1.4 $Y2=1.395
cc_58 VPB N_Z_c_325_n 0.0105741f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_59 VPB N_Z_c_322_n 0.00328219f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 N_TE_B_c_68_n N_A_27_47#_c_111_n 0.00714934f $X=1.4 $Y=1.395 $X2=0 $Y2=0
cc_61 N_TE_B_M1004_g N_A_27_47#_c_113_n 0.00440201f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_62 N_TE_B_c_65_n N_A_27_47#_c_118_n 0.0123666f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_63 N_TE_B_c_60_n N_A_27_47#_c_114_n 0.0113076f $X=0.495 $Y=1.47 $X2=0 $Y2=0
cc_64 N_TE_B_c_64_n N_A_27_47#_c_114_n 0.0165034f $X=0.495 $Y=1.67 $X2=0 $Y2=0
cc_65 N_TE_B_c_65_n N_A_27_47#_c_114_n 0.00914214f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_66 N_TE_B_c_66_n N_A_27_47#_c_114_n 0.0160355f $X=0.93 $Y=1.395 $X2=0 $Y2=0
cc_67 N_TE_B_c_67_n N_A_27_47#_c_114_n 0.00667189f $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_68 N_TE_B_c_70_n N_A_27_47#_c_114_n 0.00687677f $X=1.02 $Y=1.395 $X2=0 $Y2=0
cc_69 TE_B N_A_27_47#_c_114_n 0.0276632f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_70 N_TE_B_c_60_n N_A_27_47#_c_115_n 0.0202305f $X=0.495 $Y=1.47 $X2=0 $Y2=0
cc_71 N_TE_B_M1004_g N_A_27_47#_c_115_n 0.0262746f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_72 TE_B N_A_27_47#_c_115_n 0.042038f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_73 N_TE_B_c_70_n N_A_27_47#_c_116_n 0.0206866f $X=1.02 $Y=1.395 $X2=0 $Y2=0
cc_74 N_TE_B_c_68_n N_A_27_47#_c_117_n 3.89238e-19 $X=1.4 $Y=1.395 $X2=0 $Y2=0
cc_75 N_TE_B_c_65_n N_VPWR_c_225_n 0.0165036f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_76 N_TE_B_c_67_n N_VPWR_c_225_n 0.0108784f $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_77 N_TE_B_c_69_n N_VPWR_c_225_n 5.83063e-19 $X=1.49 $Y=1.47 $X2=0 $Y2=0
cc_78 N_TE_B_c_67_n N_VPWR_c_226_n 5.96983e-19 $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_79 N_TE_B_c_69_n N_VPWR_c_226_n 0.0110177f $X=1.49 $Y=1.47 $X2=0 $Y2=0
cc_80 N_TE_B_c_67_n N_VPWR_c_227_n 0.00642146f $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_81 N_TE_B_c_69_n N_VPWR_c_227_n 0.00311027f $X=1.49 $Y=1.47 $X2=0 $Y2=0
cc_82 N_TE_B_c_65_n N_VPWR_c_230_n 0.00427505f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_83 N_TE_B_c_65_n N_VPWR_c_224_n 0.00835414f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_84 N_TE_B_c_67_n N_VPWR_c_224_n 0.0107862f $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_85 N_TE_B_c_69_n N_VPWR_c_224_n 0.00374038f $X=1.49 $Y=1.47 $X2=0 $Y2=0
cc_86 N_TE_B_c_67_n N_A_222_309#_c_281_n 0.00136916f $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_87 N_TE_B_c_68_n N_A_222_309#_c_281_n 2.12311e-19 $X=1.4 $Y=1.395 $X2=0 $Y2=0
cc_88 N_TE_B_c_69_n N_A_222_309#_c_281_n 0.00393677f $X=1.49 $Y=1.47 $X2=0 $Y2=0
cc_89 N_TE_B_c_67_n N_A_222_309#_c_280_n 0.00802954f $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_90 N_TE_B_c_68_n N_A_222_309#_c_280_n 0.00813048f $X=1.4 $Y=1.395 $X2=0 $Y2=0
cc_91 N_TE_B_c_69_n N_A_222_309#_c_280_n 0.0297722f $X=1.49 $Y=1.47 $X2=0 $Y2=0
cc_92 N_TE_B_c_69_n N_Z_c_325_n 8.84519e-19 $X=1.49 $Y=1.47 $X2=0 $Y2=0
cc_93 N_TE_B_M1004_g N_VGND_c_363_n 0.0126377f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_94 N_TE_B_M1004_g N_VGND_c_366_n 0.00198948f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_95 N_TE_B_M1004_g N_VGND_c_368_n 0.00369246f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_96 N_TE_B_M1004_g N_A_234_47#_c_413_n 0.00417016f $X=0.52 $Y=0.445 $X2=0
+ $Y2=0
cc_97 N_A_27_47#_c_112_n N_A_M1003_g 0.0189987f $X=1.975 $Y=0.96 $X2=0 $Y2=0
cc_98 N_A_27_47#_c_116_n N_A_M1003_g 0.0024483f $X=1.935 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_27_47#_c_117_n N_A_M1003_g 0.0108025f $X=1.935 $Y=1.035 $X2=0 $Y2=0
cc_100 N_A_27_47#_c_114_n N_VPWR_M1001_d 0.00326699f $X=0.72 $Y=1.555 $X2=-0.19
+ $Y2=-0.24
cc_101 N_A_27_47#_c_118_n N_VPWR_c_225_n 0.0443303f $X=0.26 $Y=2.165 $X2=0 $Y2=0
cc_102 N_A_27_47#_c_114_n N_VPWR_c_225_n 0.0271869f $X=0.72 $Y=1.555 $X2=0 $Y2=0
cc_103 N_A_27_47#_c_118_n N_VPWR_c_230_n 0.0182101f $X=0.26 $Y=2.165 $X2=0 $Y2=0
cc_104 N_A_27_47#_M1001_s N_VPWR_c_224_n 0.00430086f $X=0.135 $Y=1.845 $X2=0
+ $Y2=0
cc_105 N_A_27_47#_c_118_n N_VPWR_c_224_n 0.00993603f $X=0.26 $Y=2.165 $X2=0
+ $Y2=0
cc_106 N_A_27_47#_c_116_n N_A_222_309#_c_279_n 0.00679059f $X=1.935 $Y=1.16
+ $X2=0 $Y2=0
cc_107 N_A_27_47#_c_117_n N_A_222_309#_c_279_n 0.00285081f $X=1.935 $Y=1.035
+ $X2=0 $Y2=0
cc_108 N_A_27_47#_c_111_n N_A_222_309#_c_280_n 0.00118695f $X=1.63 $Y=1.035
+ $X2=0 $Y2=0
cc_109 N_A_27_47#_c_114_n N_A_222_309#_c_280_n 0.019261f $X=0.72 $Y=1.555 $X2=0
+ $Y2=0
cc_110 N_A_27_47#_c_116_n N_A_222_309#_c_280_n 0.0629552f $X=1.935 $Y=1.16 $X2=0
+ $Y2=0
cc_111 N_A_27_47#_c_117_n N_A_222_309#_c_280_n 0.0035639f $X=1.935 $Y=1.035
+ $X2=0 $Y2=0
cc_112 N_A_27_47#_c_116_n N_Z_c_325_n 0.00281867f $X=1.935 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_27_47#_c_112_n N_Z_c_322_n 0.00104132f $X=1.975 $Y=0.96 $X2=0 $Y2=0
cc_114 N_A_27_47#_c_116_n N_Z_c_322_n 0.0169441f $X=1.935 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_27_47#_c_117_n N_Z_c_322_n 6.96903e-19 $X=1.935 $Y=1.035 $X2=0 $Y2=0
cc_116 N_A_27_47#_c_115_n N_VGND_M1004_d 0.00277784f $X=0.945 $Y=1.135 $X2=-0.19
+ $Y2=-0.24
cc_117 N_A_27_47#_c_109_n N_VGND_c_363_n 0.0025078f $X=1.555 $Y=0.96 $X2=0 $Y2=0
cc_118 N_A_27_47#_c_113_n N_VGND_c_363_n 0.0177195f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_119 N_A_27_47#_c_115_n N_VGND_c_363_n 0.028875f $X=0.945 $Y=1.135 $X2=0 $Y2=0
cc_120 N_A_27_47#_c_109_n N_VGND_c_364_n 0.00341689f $X=1.555 $Y=0.96 $X2=0
+ $Y2=0
cc_121 N_A_27_47#_c_109_n N_VGND_c_365_n 0.00886746f $X=1.555 $Y=0.96 $X2=0
+ $Y2=0
cc_122 N_A_27_47#_c_112_n N_VGND_c_365_n 0.00811151f $X=1.975 $Y=0.96 $X2=0
+ $Y2=0
cc_123 N_A_27_47#_c_113_n N_VGND_c_366_n 0.0179755f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_115_n N_VGND_c_366_n 0.00279825f $X=0.945 $Y=1.135 $X2=0
+ $Y2=0
cc_125 N_A_27_47#_c_112_n N_VGND_c_367_n 0.00341689f $X=1.975 $Y=0.96 $X2=0
+ $Y2=0
cc_126 N_A_27_47#_M1004_s N_VGND_c_368_n 0.00292082f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_127 N_A_27_47#_c_109_n N_VGND_c_368_n 0.00540327f $X=1.555 $Y=0.96 $X2=0
+ $Y2=0
cc_128 N_A_27_47#_c_112_n N_VGND_c_368_n 0.00434166f $X=1.975 $Y=0.96 $X2=0
+ $Y2=0
cc_129 N_A_27_47#_c_113_n N_VGND_c_368_n 0.00989054f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_130 N_A_27_47#_c_115_n N_VGND_c_368_n 0.00625509f $X=0.945 $Y=1.135 $X2=0
+ $Y2=0
cc_131 N_A_27_47#_c_109_n N_A_234_47#_c_415_n 0.00940897f $X=1.555 $Y=0.96 $X2=0
+ $Y2=0
cc_132 N_A_27_47#_c_110_n N_A_234_47#_c_415_n 0.00181329f $X=1.8 $Y=1.035 $X2=0
+ $Y2=0
cc_133 N_A_27_47#_c_112_n N_A_234_47#_c_415_n 0.0102743f $X=1.975 $Y=0.96 $X2=0
+ $Y2=0
cc_134 N_A_27_47#_c_116_n N_A_234_47#_c_415_n 0.0505724f $X=1.935 $Y=1.16 $X2=0
+ $Y2=0
cc_135 N_A_27_47#_c_109_n N_A_234_47#_c_413_n 0.00977934f $X=1.555 $Y=0.96 $X2=0
+ $Y2=0
cc_136 N_A_27_47#_c_115_n N_A_234_47#_c_413_n 0.0156018f $X=0.945 $Y=1.135 $X2=0
+ $Y2=0
cc_137 N_A_27_47#_c_116_n N_A_234_47#_c_413_n 0.0268006f $X=1.935 $Y=1.16 $X2=0
+ $Y2=0
cc_138 N_A_c_181_n N_VPWR_c_229_n 0.0150535f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_c_182_n N_VPWR_c_229_n 0.00115985f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_c_181_n N_VPWR_c_231_n 0.00452725f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_c_182_n N_VPWR_c_231_n 0.00597712f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_c_181_n N_VPWR_c_224_n 0.00516686f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_c_182_n N_VPWR_c_224_n 0.0112863f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_181_n N_A_222_309#_c_279_n 0.0172938f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_c_182_n N_A_222_309#_c_279_n 0.0017602f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_c_181_n N_A_222_309#_c_295_n 0.00406869f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_c_182_n N_A_222_309#_c_295_n 0.00106439f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_c_181_n N_A_222_309#_c_280_n 0.00414624f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_c_181_n Z 0.0110655f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_c_182_n Z 0.0208407f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_c_179_n Z 0.0103429f $X=3.015 $Y=1.202 $X2=0 $Y2=0
cc_152 A Z 0.0415496f $X=3.295 $Y=1.19 $X2=0 $Y2=0
cc_153 N_A_c_181_n Z 0.00102085f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_c_182_n Z 0.0156233f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_M1003_g N_Z_c_322_n 0.0133333f $X=2.52 $Y=0.56 $X2=0 $Y2=0
cc_156 N_A_c_181_n N_Z_c_322_n 0.0019019f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_c_178_n N_Z_c_322_n 0.00725869f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A_c_182_n N_Z_c_322_n 9.12153e-19 $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_c_179_n N_Z_c_322_n 0.0333456f $X=3.015 $Y=1.202 $X2=0 $Y2=0
cc_160 A N_Z_c_322_n 0.0156722f $X=3.295 $Y=1.19 $X2=0 $Y2=0
cc_161 N_A_M1003_g N_VGND_c_365_n 0.00110206f $X=2.52 $Y=0.56 $X2=0 $Y2=0
cc_162 N_A_M1003_g N_VGND_c_367_n 0.00357877f $X=2.52 $Y=0.56 $X2=0 $Y2=0
cc_163 N_A_c_178_n N_VGND_c_367_n 0.00357877f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_M1003_g N_VGND_c_368_n 0.00570228f $X=2.52 $Y=0.56 $X2=0 $Y2=0
cc_165 N_A_c_178_n N_VGND_c_368_n 0.00654724f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A_M1003_g N_A_234_47#_c_415_n 0.00128808f $X=2.52 $Y=0.56 $X2=0 $Y2=0
cc_167 N_A_M1003_g N_A_234_47#_c_423_n 0.00407416f $X=2.52 $Y=0.56 $X2=0 $Y2=0
cc_168 N_A_M1003_g N_A_234_47#_c_411_n 0.0102043f $X=2.52 $Y=0.56 $X2=0 $Y2=0
cc_169 N_A_c_178_n N_A_234_47#_c_411_n 0.0135444f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_c_179_n N_A_234_47#_c_411_n 0.00223016f $X=3.015 $Y=1.202 $X2=0 $Y2=0
cc_171 A N_A_234_47#_c_411_n 0.00347749f $X=3.295 $Y=1.19 $X2=0 $Y2=0
cc_172 N_A_c_178_n N_A_234_47#_c_412_n 0.00484527f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A_c_179_n N_A_234_47#_c_412_n 0.00279554f $X=3.015 $Y=1.202 $X2=0 $Y2=0
cc_174 A N_A_234_47#_c_412_n 0.0142244f $X=3.295 $Y=1.19 $X2=0 $Y2=0
cc_175 N_VPWR_c_224_n N_A_222_309#_M1000_s 0.00462612f $X=3.45 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_176 N_VPWR_c_224_n N_A_222_309#_M1007_s 0.00465719f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_177 N_VPWR_c_225_n N_A_222_309#_c_281_n 0.0230841f $X=0.755 $Y=2.02 $X2=0
+ $Y2=0
cc_178 N_VPWR_c_226_n N_A_222_309#_c_281_n 0.016427f $X=1.785 $Y=2.53 $X2=0
+ $Y2=0
cc_179 N_VPWR_c_227_n N_A_222_309#_c_281_n 0.0113299f $X=1.51 $Y=2.53 $X2=0
+ $Y2=0
cc_180 N_VPWR_c_224_n N_A_222_309#_c_281_n 0.00637602f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_181 N_VPWR_c_228_n N_A_222_309#_c_279_n 0.0340519f $X=2.2 $Y=2.53 $X2=0 $Y2=0
cc_182 N_VPWR_c_231_n N_A_222_309#_c_279_n 0.0032312f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_183 N_VPWR_c_224_n N_A_222_309#_c_279_n 0.00546504f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_184 N_VPWR_c_229_n N_A_222_309#_c_295_n 0.013449f $X=2.475 $Y=2.53 $X2=0
+ $Y2=0
cc_185 N_VPWR_c_231_n N_A_222_309#_c_295_n 0.0117062f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_186 N_VPWR_c_224_n N_A_222_309#_c_295_n 0.00644886f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_187 N_VPWR_M1002_d N_A_222_309#_c_280_n 0.00490108f $X=1.58 $Y=1.545 $X2=0
+ $Y2=0
cc_188 N_VPWR_c_225_n N_A_222_309#_c_280_n 0.0128103f $X=0.755 $Y=2.02 $X2=0
+ $Y2=0
cc_189 N_VPWR_c_226_n N_A_222_309#_c_280_n 0.0340519f $X=1.785 $Y=2.53 $X2=0
+ $Y2=0
cc_190 N_VPWR_c_227_n N_A_222_309#_c_280_n 0.00259877f $X=1.51 $Y=2.53 $X2=0
+ $Y2=0
cc_191 N_VPWR_c_224_n N_A_222_309#_c_280_n 0.00912831f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_192 N_VPWR_c_228_n N_Z_M1007_d 8.06578e-19 $X=2.2 $Y=2.53 $X2=0 $Y2=0
cc_193 N_VPWR_c_229_n N_Z_M1007_d 0.00313808f $X=2.475 $Y=2.53 $X2=0 $Y2=0
cc_194 N_VPWR_c_224_n N_Z_M1009_d 0.0021832f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_195 N_VPWR_c_231_n Z 0.0331047f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_196 N_VPWR_c_224_n Z 0.0188633f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_197 N_A_222_309#_c_279_n N_Z_M1007_d 0.00623747f $X=2.695 $Y=1.975 $X2=0
+ $Y2=0
cc_198 N_A_222_309#_M1007_s Z 0.00182874f $X=2.635 $Y=1.485 $X2=0 $Y2=0
cc_199 N_A_222_309#_c_279_n Z 0.014061f $X=2.695 $Y=1.975 $X2=0 $Y2=0
cc_200 N_A_222_309#_c_279_n Z 0.0187115f $X=2.695 $Y=1.975 $X2=0 $Y2=0
cc_201 N_A_222_309#_c_295_n Z 0.0289569f $X=2.78 $Y=2.265 $X2=0 $Y2=0
cc_202 N_A_222_309#_c_279_n N_Z_c_325_n 0.0322407f $X=2.695 $Y=1.975 $X2=0 $Y2=0
cc_203 N_A_222_309#_c_280_n N_Z_c_325_n 0.0193624f $X=1.925 $Y=1.765 $X2=0 $Y2=0
cc_204 N_Z_M1003_s N_VGND_c_368_n 0.00256987f $X=2.595 $Y=0.235 $X2=0 $Y2=0
cc_205 N_Z_c_325_n N_A_234_47#_c_415_n 0.0029497f $X=2.445 $Y=1.57 $X2=0 $Y2=0
cc_206 N_Z_c_322_n N_A_234_47#_c_415_n 0.0138372f $X=2.73 $Y=0.76 $X2=0 $Y2=0
cc_207 N_Z_c_322_n N_A_234_47#_c_423_n 0.0043353f $X=2.73 $Y=0.76 $X2=0 $Y2=0
cc_208 N_Z_M1003_s N_A_234_47#_c_411_n 0.00498317f $X=2.595 $Y=0.235 $X2=0 $Y2=0
cc_209 N_Z_c_322_n N_A_234_47#_c_411_n 0.0229345f $X=2.73 $Y=0.76 $X2=0 $Y2=0
cc_210 N_Z_c_322_n N_A_234_47#_c_412_n 0.00842979f $X=2.73 $Y=0.76 $X2=0 $Y2=0
cc_211 N_VGND_c_368_n N_A_234_47#_M1005_d 0.0028969f $X=3.45 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_212 N_VGND_c_368_n N_A_234_47#_M1006_d 0.00336888f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_213 N_VGND_c_368_n N_A_234_47#_M1008_d 0.00251122f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_214 N_VGND_M1005_s N_A_234_47#_c_415_n 0.00304947f $X=1.63 $Y=0.235 $X2=0
+ $Y2=0
cc_215 N_VGND_c_364_n N_A_234_47#_c_415_n 0.00310196f $X=1.6 $Y=0 $X2=0 $Y2=0
cc_216 N_VGND_c_365_n N_A_234_47#_c_415_n 0.0160613f $X=1.765 $Y=0.36 $X2=0
+ $Y2=0
cc_217 N_VGND_c_367_n N_A_234_47#_c_415_n 0.00232396f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_218 N_VGND_c_368_n N_A_234_47#_c_415_n 0.0111001f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_219 N_VGND_c_367_n N_A_234_47#_c_411_n 0.0684056f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_220 N_VGND_c_368_n N_A_234_47#_c_411_n 0.0422894f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_221 N_VGND_c_367_n N_A_234_47#_c_447_n 0.0115639f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_222 N_VGND_c_368_n N_A_234_47#_c_447_n 0.00651702f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_223 N_VGND_c_363_n N_A_234_47#_c_413_n 0.0192911f $X=0.73 $Y=0.38 $X2=0 $Y2=0
cc_224 N_VGND_c_364_n N_A_234_47#_c_413_n 0.0218666f $X=1.6 $Y=0 $X2=0 $Y2=0
cc_225 N_VGND_c_365_n N_A_234_47#_c_413_n 0.0145922f $X=1.765 $Y=0.36 $X2=0
+ $Y2=0
cc_226 N_VGND_c_368_n N_A_234_47#_c_413_n 0.011999f $X=3.45 $Y=0 $X2=0 $Y2=0
