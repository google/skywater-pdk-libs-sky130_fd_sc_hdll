* File: sky130_fd_sc_hdll__a31o_2.spice
* Created: Wed Sep  2 08:19:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a31o_2.pex.spice"
.subckt sky130_fd_sc_hdll__a31o_2  VNB VPB A3 A2 A1 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_79_21#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A_79_21#_M1009_g N_X_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1011 A_307_47# N_A3_M1011_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.104 PD=0.92 PS=0.97 NRD=14.76 NRS=8.304 M=1 R=4.33333 SA=75001.2
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1010 A_391_47# N_A2_M1010_g A_307_47# VNB NSHORT L=0.15 W=0.65 AD=0.1235
+ AS=0.08775 PD=1.03 PS=0.92 NRD=24.912 NRS=14.76 M=1 R=4.33333 SA=75001.6
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1002 N_A_79_21#_M1002_d N_A1_M1002_g A_391_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.1235 PD=1.17 PS=1.03 NRD=45.228 NRS=24.912 M=1 R=4.33333
+ SA=75002.1 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_B1_M1003_g N_A_79_21#_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.169 PD=1.82 PS=1.17 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_79_21#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.7 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A_79_21#_M1005_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1008 N_A_305_297#_M1008_d N_A3_M1008_g N_VPWR_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A2_M1006_g N_A_305_297#_M1008_d VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.145 PD=1.35 PS=1.29 NRD=8.8453 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1004 N_A_305_297#_M1004_d N_A1_M1004_g N_VPWR_M1006_d VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=12.7853 NRS=4.9053 M=1 R=5.55556
+ SA=90002.1 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1007 N_A_79_21#_M1007_d N_B1_M1007_g N_A_305_297#_M1004_d VPB PHIGHVT L=0.18
+ W=1 AD=0.33 AS=0.175 PD=2.66 PS=1.35 NRD=12.7853 NRS=0.9653 M=1 R=5.55556
+ SA=90002.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hdll__a31o_2.pxi.spice"
*
.ends
*
*
