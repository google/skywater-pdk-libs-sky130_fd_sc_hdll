* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
X0 a_615_93# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_511_93# C a_615_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND a_339_93# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR C a_339_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X4 a_339_93# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X5 VPWR B_N a_225_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X6 a_339_93# a_27_47# a_425_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_425_93# a_225_413# a_511_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_27_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_339_93# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_27_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X11 VPWR a_27_47# a_339_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X12 a_339_93# a_225_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X13 VGND B_N a_225_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
