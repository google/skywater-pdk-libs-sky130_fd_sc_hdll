* File: sky130_fd_sc_hdll__and4_2.pex.spice
* Created: Thu Aug 27 18:58:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND4_2%A 2 3 5 8 10 11 12 13 23
r35 22 23 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r36 19 22 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.495 $Y2=1.16
r37 12 13 18.3947 $w=2.03e-07 $l=3.4e-07 $layer=LI1_cond $X=0.227 $Y=1.53
+ $X2=0.227 $Y2=1.87
r38 11 12 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.227 $Y=1.16
+ $X2=0.227 $Y2=1.53
r39 11 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r40 10 11 16.7716 $w=2.03e-07 $l=3.1e-07 $layer=LI1_cond $X=0.227 $Y=0.85
+ $X2=0.227 $Y2=1.16
r41 6 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.16
r42 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r43 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r44 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.89 $X2=0.495
+ $Y2=1.99
r45 1 22 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r46 1 2 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_2%B 3 6 7 9 10 11 15
r38 15 18 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.16 $X2=1
+ $Y2=1.325
r39 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.16 $X2=1
+ $Y2=0.995
r40 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.16
+ $X2=1 $Y2=1.16
r41 11 16 9.40151 $w=3.78e-07 $l=3.1e-07 $layer=LI1_cond $X=1.045 $Y=0.85
+ $X2=1.045 $Y2=1.16
r42 10 11 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=1.045 $Y=0.51
+ $X2=1.045 $Y2=0.85
r43 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.965 $Y=1.99
+ $X2=0.965 $Y2=2.275
r44 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.89 $X2=0.965
+ $Y2=1.99
r45 6 18 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.965 $Y=1.89
+ $X2=0.965 $Y2=1.325
r46 3 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.94 $Y=0.445
+ $X2=0.94 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_2%C 3 6 7 9 10 11 12 17
c38 17 0 1.0356e-19 $X=1.49 $Y=1.16
r39 17 20 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=1.16
+ $X2=1.49 $Y2=1.325
r40 17 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=1.16
+ $X2=1.49 $Y2=0.995
r41 12 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.49
+ $Y=1.16 $X2=1.49 $Y2=1.16
r42 11 12 11.9086 $w=2.98e-07 $l=3.1e-07 $layer=LI1_cond $X=1.555 $Y=0.85
+ $X2=1.555 $Y2=1.16
r43 10 11 13.061 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=1.555 $Y=0.51
+ $X2=1.555 $Y2=0.85
r44 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.455 $Y=1.99
+ $X2=1.455 $Y2=2.275
r45 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.455 $Y=1.89 $X2=1.455
+ $Y2=1.99
r46 6 20 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=1.455 $Y=1.89
+ $X2=1.455 $Y2=1.325
r47 3 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.43 $Y=0.445
+ $X2=1.43 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_2%D 3 6 7 9 10 11 15
r42 15 18 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.97 $Y=1.16
+ $X2=1.97 $Y2=1.325
r43 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.97 $Y=1.16
+ $X2=1.97 $Y2=0.995
r44 11 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.97
+ $Y=1.16 $X2=1.97 $Y2=1.16
r45 10 11 13.2318 $w=2.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.02 $Y=0.85
+ $X2=2.02 $Y2=1.16
r46 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.935 $Y=1.99
+ $X2=1.935 $Y2=2.275
r47 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.935 $Y=1.89 $X2=1.935
+ $Y2=1.99
r48 6 18 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=1.935 $Y=1.89
+ $X2=1.935 $Y2=1.325
r49 3 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.91 $Y=0.445
+ $X2=1.91 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_2%A_27_47# 1 2 3 10 12 13 15 16 18 19 21 23
+ 26 28 29 32 34 38 44 49 52
c102 52 0 1.89144e-19 $X=3.135 $Y=1.202
c103 28 0 1.0356e-19 $X=1.57 $Y=1.58
r104 52 53 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=3.135 $Y=1.202
+ $X2=3.16 $Y2=1.202
r105 51 52 68.4879 $w=3.73e-07 $l=5.3e-07 $layer=POLY_cond $X=2.605 $Y=1.202
+ $X2=3.135 $Y2=1.202
r106 46 48 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.585 $Y=1.58
+ $X2=0.73 $Y2=1.58
r107 42 44 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.26 $Y=0.42
+ $X2=0.585 $Y2=0.42
r108 39 51 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=2.58 $Y=1.202
+ $X2=2.605 $Y2=1.202
r109 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.58
+ $Y=1.16 $X2=2.58 $Y2=1.16
r110 36 38 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.58 $Y=1.495
+ $X2=2.58 $Y2=1.16
r111 35 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.82 $Y=1.58
+ $X2=1.695 $Y2=1.58
r112 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.495 $Y=1.58
+ $X2=2.58 $Y2=1.495
r113 34 35 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.495 $Y=1.58
+ $X2=1.82 $Y2=1.58
r114 30 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=1.58
r115 30 32 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=2.3
r116 29 48 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=1.58
+ $X2=0.73 $Y2=1.58
r117 28 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.57 $Y=1.58
+ $X2=1.695 $Y2=1.58
r118 28 29 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.57 $Y=1.58
+ $X2=0.815 $Y2=1.58
r119 24 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=1.58
r120 24 26 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=2.3
r121 23 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.585 $Y=1.495
+ $X2=0.585 $Y2=1.58
r122 22 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0.585
+ $X2=0.585 $Y2=0.42
r123 22 23 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=0.585 $Y=0.585
+ $X2=0.585 $Y2=1.495
r124 19 53 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.16 $Y=0.995
+ $X2=3.16 $Y2=1.202
r125 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.16 $Y=0.995
+ $X2=3.16 $Y2=0.56
r126 16 52 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.135 $Y=1.41
+ $X2=3.135 $Y2=1.202
r127 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.135 $Y=1.41
+ $X2=3.135 $Y2=1.985
r128 13 51 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.605 $Y=1.41
+ $X2=2.605 $Y2=1.202
r129 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.605 $Y=1.41
+ $X2=2.605 $Y2=1.985
r130 10 39 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.58 $Y=0.995
+ $X2=2.58 $Y2=1.202
r131 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.58 $Y=0.995
+ $X2=2.58 $Y2=0.56
r132 3 32 600 $w=1.7e-07 $l=3.00791e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=2.065 $X2=1.695 $Y2=2.3
r133 2 26 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.065 $X2=0.73 $Y2=2.3
r134 1 42 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_2%VPWR 1 2 3 4 13 15 19 23 25 27 30 31 32 34
+ 43 51 55
r54 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r55 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r56 46 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r57 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r58 43 54 4.64351 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=3.245 $Y=2.72
+ $X2=3.462 $Y2=2.72
r59 43 45 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.245 $Y=2.72
+ $X2=2.99 $Y2=2.72
r60 42 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r61 42 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r62 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r63 39 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.2 $Y2=2.72
r64 39 41 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=2.07 $Y2=2.72
r65 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r66 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r67 35 48 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r68 35 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=1.2 $Y2=2.72
r70 34 37 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=0.69 $Y2=2.72
r71 32 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r72 32 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r73 30 41 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.165 $Y=2.72
+ $X2=2.07 $Y2=2.72
r74 30 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.165 $Y=2.72
+ $X2=2.29 $Y2=2.72
r75 29 45 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.415 $Y=2.72
+ $X2=2.99 $Y2=2.72
r76 29 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.415 $Y=2.72
+ $X2=2.29 $Y2=2.72
r77 25 54 3.03861 $w=3.2e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.405 $Y=2.635
+ $X2=3.462 $Y2=2.72
r78 25 27 22.8688 $w=3.18e-07 $l=6.35e-07 $layer=LI1_cond $X=3.405 $Y=2.635
+ $X2=3.405 $Y2=2
r79 21 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=2.635
+ $X2=2.29 $Y2=2.72
r80 21 23 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=2.29 $Y=2.635
+ $X2=2.29 $Y2=2
r81 17 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.72
r82 17 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.34
r83 13 48 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r84 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r85 4 27 300 $w=1.7e-07 $l=5.96112e-07 $layer=licon1_PDIFF $count=2 $X=3.225
+ $Y=1.485 $X2=3.4 $Y2=2
r86 3 23 300 $w=1.7e-07 $l=3.35932e-07 $layer=licon1_PDIFF $count=2 $X=2.025
+ $Y=2.065 $X2=2.33 $Y2=2
r87 2 19 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=2.065 $X2=1.2 $Y2=2.34
r88 1 15 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_2%X 1 2 7 8 9 10 11 12 24 32 39
r25 39 40 3.51978 $w=4.48e-07 $l=3.5e-08 $layer=LI1_cond $X=2.85 $Y=1.87
+ $X2=2.85 $Y2=1.835
r26 24 37 2.16083 $w=2.38e-07 $l=4.5e-08 $layer=LI1_cond $X=2.955 $Y=0.85
+ $X2=2.955 $Y2=0.805
r27 12 43 5.5817 $w=4.48e-07 $l=2.1e-07 $layer=LI1_cond $X=2.85 $Y=2.21 $X2=2.85
+ $Y2=2
r28 11 43 2.79085 $w=4.48e-07 $l=1.05e-07 $layer=LI1_cond $X=2.85 $Y=1.895
+ $X2=2.85 $Y2=2
r29 11 39 0.664488 $w=4.48e-07 $l=2.5e-08 $layer=LI1_cond $X=2.85 $Y=1.895
+ $X2=2.85 $Y2=1.87
r30 11 40 1.20046 $w=2.38e-07 $l=2.5e-08 $layer=LI1_cond $X=2.955 $Y=1.81
+ $X2=2.955 $Y2=1.835
r31 10 11 13.4452 $w=2.38e-07 $l=2.8e-07 $layer=LI1_cond $X=2.955 $Y=1.53
+ $X2=2.955 $Y2=1.81
r32 9 10 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.955 $Y=1.19
+ $X2=2.955 $Y2=1.53
r33 8 37 3.12109 $w=4.48e-07 $l=2e-08 $layer=LI1_cond $X=2.85 $Y=0.785 $X2=2.85
+ $Y2=0.805
r34 8 9 15.3659 $w=2.38e-07 $l=3.2e-07 $layer=LI1_cond $X=2.955 $Y=0.87
+ $X2=2.955 $Y2=1.19
r35 8 24 0.960369 $w=2.38e-07 $l=2e-08 $layer=LI1_cond $X=2.955 $Y=0.87
+ $X2=2.955 $Y2=0.85
r36 7 8 7.30937 $w=4.48e-07 $l=2.75e-07 $layer=LI1_cond $X=2.85 $Y=0.51 $X2=2.85
+ $Y2=0.785
r37 7 32 3.45534 $w=4.48e-07 $l=1.3e-07 $layer=LI1_cond $X=2.85 $Y=0.51 $X2=2.85
+ $Y2=0.38
r38 2 43 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.695
+ $Y=1.485 $X2=2.84 $Y2=2
r39 1 32 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=2.655
+ $Y=0.235 $X2=2.84 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_2%VGND 1 2 9 11 13 16 17 18 27 33
c41 9 0 1.89144e-19 $X=2.37 $Y=0.385
r42 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r43 30 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r44 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r45 27 32 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=3.245 $Y=0 $X2=3.462
+ $Y2=0
r46 27 29 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.245 $Y=0 $X2=2.99
+ $Y2=0
r47 26 30 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r48 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r49 21 25 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r50 18 26 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r51 18 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r52 16 25 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.07
+ $Y2=0
r53 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.37
+ $Y2=0
r54 15 29 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.99
+ $Y2=0
r55 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.37
+ $Y2=0
r56 11 32 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=3.41 $Y=0.085
+ $X2=3.462 $Y2=0
r57 11 13 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.41 $Y=0.085 $X2=3.41
+ $Y2=0.385
r58 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.37 $Y=0.085 $X2=2.37
+ $Y2=0
r59 7 9 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.37 $Y=0.085 $X2=2.37
+ $Y2=0.385
r60 2 13 91 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_NDIFF $count=2 $X=3.235
+ $Y=0.235 $X2=3.41 $Y2=0.385
r61 1 9 182 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_NDIFF $count=1 $X=1.985
+ $Y=0.235 $X2=2.37 $Y2=0.385
.ends

