* NGSPICE file created from sky130_fd_sc_hdll__xor2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__xor2_4 A B VGND VNB VPB VPWR X
M1000 a_27_297# B a_112_47# VPB phighvt w=1e+06u l=180000u
+  ad=1.425e+12p pd=1.285e+07u as=5.8e+11p ps=5.16e+06u
M1001 VPWR A a_886_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.74e+12p pd=1.548e+07u as=1.9868e+12p ps=1.798e+07u
M1002 X B a_886_47# VNB nshort w=650000u l=150000u
+  ad=8.97e+11p pd=7.96e+06u as=9.295e+11p ps=9.36e+06u
M1003 a_112_47# A VGND VNB nshort w=650000u l=150000u
+  ad=8.645e+11p pd=7.86e+06u as=1.97925e+12p ps=1.909e+07u
M1004 a_886_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_112_47# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_886_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A a_886_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR B a_886_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_112_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B a_112_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A a_886_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A a_112_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_886_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_886_297# a_112_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.6245e+11p ps=7.74e+06u
M1017 X B a_886_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_886_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_112_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_886_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_886_47# B X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_297# B a_112_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X a_112_47# a_886_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_112_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND B a_112_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR B a_886_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 X a_112_47# a_886_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_112_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND A a_112_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND A a_886_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_112_47# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_886_297# a_112_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_886_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 X a_112_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_886_47# B X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND a_112_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_112_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

