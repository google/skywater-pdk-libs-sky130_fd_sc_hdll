* File: sky130_fd_sc_hdll__a21boi_2.pex.spice
* Created: Wed Sep  2 08:16:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A21BOI_2%B1_N 2 3 5 8 10 11 13 14 17
c35 14 0 1.59155e-19 $X=0.23 $Y=0.85
r36 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.34
+ $Y=0.93 $X2=0.34 $Y2=0.93
r37 14 18 3.0228 $w=3.03e-07 $l=8e-08 $layer=LI1_cond $X=0.272 $Y=0.85 $X2=0.272
+ $Y2=0.93
r38 12 17 38.3419 $w=4.25e-07 $l=2.93e-07 $layer=POLY_cond $X=0.387 $Y=1.223
+ $X2=0.387 $Y2=0.93
r39 12 13 43.4286 $w=4.25e-07 $l=2.12e-07 $layer=POLY_cond $X=0.387 $Y=1.223
+ $X2=0.387 $Y2=1.435
r40 11 17 6.54299 $w=4.25e-07 $l=5e-08 $layer=POLY_cond $X=0.387 $Y=0.88
+ $X2=0.387 $Y2=0.93
r41 10 11 44.3146 $w=4.25e-07 $l=1.5e-07 $layer=POLY_cond $X=0.49 $Y=0.73
+ $X2=0.49 $Y2=0.88
r42 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.73 $Y=0.445 $X2=0.73
+ $Y2=0.73
r43 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.5 $Y=1.815 $X2=0.5
+ $Y2=2.1
r44 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.5 $Y=1.715 $X2=0.5
+ $Y2=1.815
r45 2 13 92.8416 $w=2e-07 $l=2.8e-07 $layer=POLY_cond $X=0.5 $Y=1.715 $X2=0.5
+ $Y2=1.435
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_2%A_61_47# 1 2 7 9 10 12 13 15 18 20 23 25
+ 30 33 37 40
c72 23 0 1.57088e-19 $X=2.015 $Y=1.202
c73 20 0 1.59155e-19 $X=1.445 $Y=1.16
r74 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.19
+ $Y=1.16 $X2=1.19 $Y2=1.16
r75 35 40 0.711257 $w=2.15e-07 $l=9e-08 $layer=LI1_cond $X=0.825 $Y=1.177
+ $X2=0.735 $Y2=1.177
r76 35 37 19.5647 $w=2.13e-07 $l=3.65e-07 $layer=LI1_cond $X=0.825 $Y=1.177
+ $X2=1.19 $Y2=1.177
r77 31 40 5.97344 $w=1.8e-07 $l=1.08e-07 $layer=LI1_cond $X=0.735 $Y=1.285
+ $X2=0.735 $Y2=1.177
r78 31 33 50.2172 $w=1.78e-07 $l=8.15e-07 $layer=LI1_cond $X=0.735 $Y=1.285
+ $X2=0.735 $Y2=2.1
r79 30 40 5.97344 $w=1.8e-07 $l=1.07e-07 $layer=LI1_cond $X=0.735 $Y=1.07
+ $X2=0.735 $Y2=1.177
r80 29 30 33.2727 $w=1.78e-07 $l=5.4e-07 $layer=LI1_cond $X=0.735 $Y=0.53
+ $X2=0.735 $Y2=1.07
r81 25 29 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.645 $Y=0.445
+ $X2=0.735 $Y2=0.53
r82 25 27 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.645 $Y=0.445
+ $X2=0.43 $Y2=0.445
r83 23 24 3.36592 $w=3.58e-07 $l=2.5e-08 $layer=POLY_cond $X=2.015 $Y=1.202
+ $X2=2.04 $Y2=1.202
r84 22 23 59.9134 $w=3.58e-07 $l=4.45e-07 $layer=POLY_cond $X=1.57 $Y=1.202
+ $X2=2.015 $Y2=1.202
r85 21 22 3.36592 $w=3.58e-07 $l=2.5e-08 $layer=POLY_cond $X=1.545 $Y=1.202
+ $X2=1.57 $Y2=1.202
r86 20 38 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=1.445 $Y=1.16
+ $X2=1.19 $Y2=1.16
r87 20 21 13.8405 $w=3.58e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.445 $Y=1.16
+ $X2=1.545 $Y2=1.202
r88 16 24 23.1716 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=2.04 $Y=1.015
+ $X2=2.04 $Y2=1.202
r89 16 18 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.04 $Y=1.015
+ $X2=2.04 $Y2=0.56
r90 13 23 18.8375 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.015 $Y=1.41
+ $X2=2.015 $Y2=1.202
r91 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.015 $Y=1.41
+ $X2=2.015 $Y2=1.985
r92 10 22 23.1716 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.57 $Y=0.995
+ $X2=1.57 $Y2=1.202
r93 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.57 $Y=0.995
+ $X2=1.57 $Y2=0.56
r94 7 21 18.8375 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.545 $Y=1.41
+ $X2=1.545 $Y2=1.202
r95 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.545 $Y=1.41
+ $X2=1.545 $Y2=1.985
r96 2 33 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.89 $X2=0.74 $Y2=2.1
r97 1 27 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.305
+ $Y=0.235 $X2=0.43 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_2%A2 1 3 4 6 7 9 10 12 14 15 16 18 22 28 29
c81 28 0 1.17192e-19 $X=3.95 $Y=1.16
c82 14 0 2.32029e-19 $X=2.487 $Y=1.495
c83 10 0 8.70193e-20 $X=3.915 $Y=1.41
r84 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.16 $X2=3.95 $Y2=1.16
r85 22 29 2.63916 $w=3.5e-07 $l=9e-08 $layer=LI1_cond $X=3.91 $Y=1.585 $X2=3.91
+ $Y2=1.495
r86 22 29 0.823174 $w=3.48e-07 $l=2.5e-08 $layer=LI1_cond $X=3.91 $Y=1.47
+ $X2=3.91 $Y2=1.495
r87 22 28 10.2074 $w=3.48e-07 $l=3.1e-07 $layer=LI1_cond $X=3.91 $Y=1.47
+ $X2=3.91 $Y2=1.16
r88 18 21 2.57783 $w=3.78e-07 $l=8.5e-08 $layer=LI1_cond $X=2.485 $Y=1.16
+ $X2=2.485 $Y2=1.245
r89 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.46
+ $Y=1.16 $X2=2.46 $Y2=1.16
r90 15 22 5.13171 $w=1.8e-07 $l=1.75e-07 $layer=LI1_cond $X=3.735 $Y=1.585
+ $X2=3.91 $Y2=1.585
r91 15 16 65.3131 $w=1.78e-07 $l=1.06e-06 $layer=LI1_cond $X=3.735 $Y=1.585
+ $X2=2.675 $Y2=1.585
r92 14 16 7.97274 $w=1.8e-07 $l=2.28613e-07 $layer=LI1_cond $X=2.487 $Y=1.495
+ $X2=2.675 $Y2=1.585
r93 14 21 7.68295 $w=3.73e-07 $l=2.5e-07 $layer=LI1_cond $X=2.487 $Y=1.495
+ $X2=2.487 $Y2=1.245
r94 10 27 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.915 $Y=1.41
+ $X2=3.95 $Y2=1.16
r95 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.915 $Y=1.41
+ $X2=3.915 $Y2=1.985
r96 7 27 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.89 $Y=0.995
+ $X2=3.95 $Y2=1.16
r97 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.89 $Y=0.995 $X2=3.89
+ $Y2=0.56
r98 4 19 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.485 $Y2=1.16
r99 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.57 $Y=0.995 $X2=2.57
+ $Y2=0.56
r100 1 19 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=2.485 $Y=1.41
+ $X2=2.485 $Y2=1.16
r101 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.485 $Y=1.41
+ $X2=2.485 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_2%A1 1 3 4 6 7 9 10 12 13 20 23
r47 20 21 3.19629 $w=3.77e-07 $l=2.5e-08 $layer=POLY_cond $X=3.41 $Y=1.202
+ $X2=3.435 $Y2=1.202
r48 18 20 3.83554 $w=3.77e-07 $l=3e-08 $layer=POLY_cond $X=3.38 $Y=1.202
+ $X2=3.41 $Y2=1.202
r49 16 18 54.3369 $w=3.77e-07 $l=4.25e-07 $layer=POLY_cond $X=2.955 $Y=1.202
+ $X2=3.38 $Y2=1.202
r50 15 16 3.19629 $w=3.77e-07 $l=2.5e-08 $layer=POLY_cond $X=2.93 $Y=1.202
+ $X2=2.955 $Y2=1.202
r51 13 23 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.315 $Y=1.16
+ $X2=3.015 $Y2=1.16
r52 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.38
+ $Y=1.16 $X2=3.38 $Y2=1.16
r53 10 21 20.0566 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.435 $Y=1.41
+ $X2=3.435 $Y2=1.202
r54 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.435 $Y=1.41
+ $X2=3.435 $Y2=1.985
r55 7 20 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=1.202
r56 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.41 $Y=0.995 $X2=3.41
+ $Y2=0.56
r57 4 16 20.0566 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.955 $Y=1.41
+ $X2=2.955 $Y2=1.202
r58 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.955 $Y=1.41
+ $X2=2.955 $Y2=1.985
r59 1 15 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.93 $Y=0.995
+ $X2=2.93 $Y2=1.202
r60 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.93 $Y=0.995 $X2=2.93
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_2%VPWR 1 2 3 10 12 16 19 20 22 25 28 41 42
c67 3 0 1.17192e-19 $X=3.525 $Y=1.485
c68 2 0 1.16442e-19 $X=2.575 $Y=1.485
r69 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r70 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r71 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r72 36 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r73 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r74 33 36 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r75 32 35 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r76 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r77 30 45 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r78 30 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r79 28 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r80 28 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r81 26 41 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.84 $Y=2.72
+ $X2=4.37 $Y2=2.72
r82 25 38 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=3.46 $Y=2.72 $X2=3.45
+ $Y2=2.72
r83 24 26 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.65 $Y=2.72 $X2=3.84
+ $Y2=2.72
r84 24 25 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.65 $Y=2.72 $X2=3.46
+ $Y2=2.72
r85 22 24 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.65 $Y=2.36
+ $X2=3.65 $Y2=2.72
r86 19 35 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.635 $Y=2.72
+ $X2=2.53 $Y2=2.72
r87 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=2.72
+ $X2=2.72 $Y2=2.72
r88 18 38 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=2.805 $Y=2.72
+ $X2=3.45 $Y2=2.72
r89 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.805 $Y=2.72
+ $X2=2.72 $Y2=2.72
r90 14 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.72 $Y=2.635
+ $X2=2.72 $Y2=2.72
r91 14 16 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.72 $Y=2.635
+ $X2=2.72 $Y2=2.36
r92 10 45 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r93 10 12 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.165
r94 3 22 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=3.525
+ $Y=1.485 $X2=3.675 $Y2=2.36
r95 2 16 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=2.575
+ $Y=1.485 $X2=2.72 $Y2=2.36
r96 1 12 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.89 $X2=0.26 $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_2%A_228_297# 1 2 3 4 15 17 18 19 20 21 25
+ 27 29 31 36
c65 29 0 8.70193e-20 $X=4.19 $Y=2.105
c66 2 0 1.15587e-19 $X=2.105 $Y=1.485
r67 29 38 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=4.19 $Y=2.105
+ $X2=4.19 $Y2=1.98
r68 29 31 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=4.19 $Y=2.105
+ $X2=4.19 $Y2=2.3
r69 28 36 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.28 $Y=1.98 $X2=3.195
+ $Y2=1.98
r70 27 38 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=4.06 $Y=1.98 $X2=4.19
+ $Y2=1.98
r71 27 28 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=4.06 $Y=1.98
+ $X2=3.28 $Y2=1.98
r72 23 36 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.195 $Y=2.105
+ $X2=3.195 $Y2=1.98
r73 23 25 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.195 $Y=2.105
+ $X2=3.195 $Y2=2.3
r74 22 34 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.415 $Y=1.94
+ $X2=2.225 $Y2=1.94
r75 21 36 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=3.11 $Y=1.94
+ $X2=3.195 $Y2=1.98
r76 21 22 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.11 $Y=1.94
+ $X2=2.415 $Y2=1.94
r77 19 34 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.025
+ $X2=2.225 $Y2=1.94
r78 19 20 7.88514 $w=3.78e-07 $l=2.6e-07 $layer=LI1_cond $X=2.225 $Y=2.025
+ $X2=2.225 $Y2=2.285
r79 17 20 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=2.035 $Y=2.375
+ $X2=2.225 $Y2=2.285
r80 17 18 42.2071 $w=1.78e-07 $l=6.85e-07 $layer=LI1_cond $X=2.035 $Y=2.375
+ $X2=1.35 $Y2=2.375
r81 13 18 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=1.225 $Y=2.285
+ $X2=1.35 $Y2=2.375
r82 13 15 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=1.225 $Y=2.285
+ $X2=1.225 $Y2=1.96
r83 4 38 600 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.485 $X2=4.155 $Y2=1.96
r84 4 31 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.485 $X2=4.155 $Y2=2.3
r85 3 36 600 $w=1.7e-07 $l=5.24667e-07 $layer=licon1_PDIFF $count=1 $X=3.045
+ $Y=1.485 $X2=3.195 $Y2=1.94
r86 3 25 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=3.045
+ $Y=1.485 $X2=3.195 $Y2=2.3
r87 2 34 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=2.105
+ $Y=1.485 $X2=2.25 $Y2=2.02
r88 1 15 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=1.14
+ $Y=1.485 $X2=1.265 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_2%Y 1 2 3 12 14 18 20 24 27
c48 14 0 1.57088e-19 $X=2.98 $Y=0.7
r49 24 27 3.00637 $w=3.43e-07 $l=9e-08 $layer=LI1_cond $X=1.697 $Y=0.51
+ $X2=1.697 $Y2=0.42
r50 20 22 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=3.17 $Y=0.36
+ $X2=3.17 $Y2=0.7
r51 16 24 3.50744 $w=3.43e-07 $l=1.05e-07 $layer=LI1_cond $X=1.697 $Y=0.615
+ $X2=1.697 $Y2=0.51
r52 16 18 2.79095 $w=3.42e-07 $l=8.5e-08 $layer=LI1_cond $X=1.697 $Y=0.615
+ $X2=1.697 $Y2=0.7
r53 15 18 3.95098 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=1.87 $Y=0.7
+ $X2=1.697 $Y2=0.7
r54 14 22 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.98 $Y=0.7 $X2=3.17
+ $Y2=0.7
r55 14 15 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=2.98 $Y=0.7
+ $X2=1.87 $Y2=0.7
r56 10 18 2.79095 $w=3.42e-07 $l=8.59942e-08 $layer=LI1_cond $X=1.695 $Y=0.785
+ $X2=1.697 $Y2=0.7
r57 10 12 27.9637 $w=3.38e-07 $l=8.25e-07 $layer=LI1_cond $X=1.695 $Y=0.785
+ $X2=1.695 $Y2=1.61
r58 3 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.635
+ $Y=1.485 $X2=1.78 $Y2=1.61
r59 2 20 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=3.005
+ $Y=0.235 $X2=3.195 $Y2=0.36
r60 1 27 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.645
+ $Y=0.235 $X2=1.78 $Y2=0.42
r61 1 18 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=1.645
+ $Y=0.235 $X2=1.78 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_2%VGND 1 2 3 12 16 18 20 23 24 25 27 36 44
+ 48
r56 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r57 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r58 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r59 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r60 39 42 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r61 38 41 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r62 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r63 36 47 4.56115 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=3.99 $Y=0 $X2=4.295
+ $Y2=0
r64 36 41 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.99 $Y=0 $X2=3.91
+ $Y2=0
r65 35 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r66 35 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r67 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r68 32 44 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.325 $Y=0 $X2=1.205
+ $Y2=0
r69 32 34 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=1.325 $Y=0 $X2=2.07
+ $Y2=0
r70 27 44 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.085 $Y=0 $X2=1.205
+ $Y2=0
r71 27 29 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=1.085 $Y=0 $X2=0.23
+ $Y2=0
r72 25 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r73 25 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r74 23 34 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.14 $Y=0 $X2=2.07
+ $Y2=0
r75 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.14 $Y=0 $X2=2.305
+ $Y2=0
r76 22 38 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.53
+ $Y2=0
r77 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.305
+ $Y2=0
r78 18 47 3.29001 $w=3.4e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.16 $Y=0.085
+ $X2=4.295 $Y2=0
r79 18 20 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=4.16 $Y=0.085
+ $X2=4.16 $Y2=0.36
r80 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=0.085
+ $X2=2.305 $Y2=0
r81 14 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.305 $Y=0.085
+ $X2=2.305 $Y2=0.36
r82 10 44 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.085
+ $X2=1.205 $Y2=0
r83 10 12 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=1.205 $Y=0.085
+ $X2=1.205 $Y2=0.38
r84 3 20 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=3.965
+ $Y=0.235 $X2=4.155 $Y2=0.36
r85 2 16 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=2.115
+ $Y=0.235 $X2=2.305 $Y2=0.36
r86 1 12 91 $w=1.7e-07 $l=4.66905e-07 $layer=licon1_NDIFF $count=2 $X=0.805
+ $Y=0.235 $X2=1.205 $Y2=0.38
.ends

