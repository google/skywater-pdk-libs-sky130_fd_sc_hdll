* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__bufinv_8 A VGND VNB VPB VPWR Y
X0 VPWR a_225_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_225_47# a_117_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND a_225_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_117_297# a_225_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 a_225_47# a_117_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 Y a_225_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 Y a_225_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 Y a_225_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y a_225_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Y a_225_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 Y a_225_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND a_117_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 Y a_225_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 VPWR a_225_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 VGND A a_117_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR a_225_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_225_47# a_117_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VGND a_225_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VGND a_225_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VPWR a_225_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 Y a_225_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 a_225_47# a_117_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VGND a_225_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
