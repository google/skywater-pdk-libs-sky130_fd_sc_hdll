* File: sky130_fd_sc_hdll__nor4bb_4.pxi.spice
* Created: Thu Aug 27 19:18:03 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR4BB_4%C_N N_C_N_c_155_n N_C_N_M1002_g N_C_N_c_152_n
+ N_C_N_M1006_g C_N N_C_N_c_154_n C_N PM_SKY130_FD_SC_HDLL__NOR4BB_4%C_N
x_PM_SKY130_FD_SC_HDLL__NOR4BB_4%D_N N_D_N_c_178_n N_D_N_M1003_g N_D_N_c_181_n
+ N_D_N_M1026_g D_N N_D_N_c_180_n D_N PM_SKY130_FD_SC_HDLL__NOR4BB_4%D_N
x_PM_SKY130_FD_SC_HDLL__NOR4BB_4%A_207_47# N_A_207_47#_M1003_d
+ N_A_207_47#_M1026_d N_A_207_47#_c_218_n N_A_207_47#_M1007_g
+ N_A_207_47#_c_230_n N_A_207_47#_M1000_g N_A_207_47#_c_219_n
+ N_A_207_47#_M1019_g N_A_207_47#_c_231_n N_A_207_47#_M1010_g
+ N_A_207_47#_c_220_n N_A_207_47#_M1027_g N_A_207_47#_c_232_n
+ N_A_207_47#_M1016_g N_A_207_47#_c_233_n N_A_207_47#_M1029_g
+ N_A_207_47#_c_221_n N_A_207_47#_M1028_g N_A_207_47#_c_222_n
+ N_A_207_47#_c_234_n N_A_207_47#_c_223_n N_A_207_47#_c_224_n
+ N_A_207_47#_c_225_n N_A_207_47#_c_226_n N_A_207_47#_c_227_n
+ N_A_207_47#_c_228_n N_A_207_47#_c_229_n
+ PM_SKY130_FD_SC_HDLL__NOR4BB_4%A_207_47#
x_PM_SKY130_FD_SC_HDLL__NOR4BB_4%A_27_297# N_A_27_297#_M1006_s
+ N_A_27_297#_M1002_s N_A_27_297#_c_342_n N_A_27_297#_M1004_g
+ N_A_27_297#_c_353_n N_A_27_297#_M1013_g N_A_27_297#_c_343_n
+ N_A_27_297#_M1005_g N_A_27_297#_c_354_n N_A_27_297#_M1018_g
+ N_A_27_297#_c_344_n N_A_27_297#_M1012_g N_A_27_297#_c_355_n
+ N_A_27_297#_M1024_g N_A_27_297#_c_356_n N_A_27_297#_M1035_g
+ N_A_27_297#_c_345_n N_A_27_297#_M1015_g N_A_27_297#_c_346_n
+ N_A_27_297#_c_357_n N_A_27_297#_c_347_n N_A_27_297#_c_348_n
+ N_A_27_297#_c_349_n N_A_27_297#_c_359_n N_A_27_297#_c_360_n
+ N_A_27_297#_c_350_n N_A_27_297#_c_351_n N_A_27_297#_c_361_n
+ N_A_27_297#_c_352_n PM_SKY130_FD_SC_HDLL__NOR4BB_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__NOR4BB_4%B N_B_c_491_n N_B_M1009_g N_B_c_497_n
+ N_B_M1001_g N_B_c_492_n N_B_M1014_g N_B_c_498_n N_B_M1011_g N_B_c_493_n
+ N_B_M1031_g N_B_c_499_n N_B_M1017_g N_B_c_500_n N_B_M1022_g N_B_c_494_n
+ N_B_M1033_g B N_B_c_495_n N_B_c_496_n B PM_SKY130_FD_SC_HDLL__NOR4BB_4%B
x_PM_SKY130_FD_SC_HDLL__NOR4BB_4%A N_A_c_568_n N_A_M1008_g N_A_c_574_n
+ N_A_M1020_g N_A_c_569_n N_A_M1021_g N_A_c_575_n N_A_M1025_g N_A_c_570_n
+ N_A_M1023_g N_A_c_576_n N_A_M1030_g N_A_c_577_n N_A_M1032_g N_A_c_571_n
+ N_A_M1034_g A N_A_c_572_n N_A_c_573_n A PM_SKY130_FD_SC_HDLL__NOR4BB_4%A
x_PM_SKY130_FD_SC_HDLL__NOR4BB_4%VPWR N_VPWR_M1002_d N_VPWR_M1020_d
+ N_VPWR_M1030_d N_VPWR_c_638_n N_VPWR_c_639_n N_VPWR_c_640_n N_VPWR_c_641_n
+ N_VPWR_c_642_n N_VPWR_c_643_n N_VPWR_c_644_n VPWR N_VPWR_c_645_n
+ N_VPWR_c_646_n N_VPWR_c_637_n N_VPWR_c_648_n
+ PM_SKY130_FD_SC_HDLL__NOR4BB_4%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR4BB_4%A_331_297# N_A_331_297#_M1000_s
+ N_A_331_297#_M1010_s N_A_331_297#_M1029_s N_A_331_297#_M1018_s
+ N_A_331_297#_M1035_s N_A_331_297#_c_743_n N_A_331_297#_c_758_n
+ N_A_331_297#_c_782_p N_A_331_297#_c_744_n N_A_331_297#_c_745_n
+ N_A_331_297#_c_762_n N_A_331_297#_c_773_n
+ PM_SKY130_FD_SC_HDLL__NOR4BB_4%A_331_297#
x_PM_SKY130_FD_SC_HDLL__NOR4BB_4%Y N_Y_M1007_s N_Y_M1027_s N_Y_M1004_d
+ N_Y_M1012_d N_Y_M1009_d N_Y_M1031_d N_Y_M1008_d N_Y_M1023_d N_Y_M1000_d
+ N_Y_M1016_d N_Y_c_808_n N_Y_c_791_n N_Y_c_792_n N_Y_c_822_n N_Y_c_793_n
+ N_Y_c_794_n N_Y_c_829_n N_Y_c_795_n N_Y_c_858_n N_Y_c_796_n N_Y_c_874_n
+ N_Y_c_797_n N_Y_c_881_n N_Y_c_798_n N_Y_c_885_n N_Y_c_799_n N_Y_c_903_n
+ N_Y_c_800_n N_Y_c_807_n N_Y_c_801_n N_Y_c_802_n N_Y_c_803_n N_Y_c_804_n
+ N_Y_c_805_n Y Y PM_SKY130_FD_SC_HDLL__NOR4BB_4%Y
x_PM_SKY130_FD_SC_HDLL__NOR4BB_4%A_797_297# N_A_797_297#_M1013_d
+ N_A_797_297#_M1024_d N_A_797_297#_M1001_s N_A_797_297#_M1017_s
+ N_A_797_297#_c_983_n N_A_797_297#_c_984_n N_A_797_297#_c_985_n
+ N_A_797_297#_c_986_n N_A_797_297#_c_987_n N_A_797_297#_c_988_n
+ N_A_797_297#_c_989_n PM_SKY130_FD_SC_HDLL__NOR4BB_4%A_797_297#
x_PM_SKY130_FD_SC_HDLL__NOR4BB_4%A_1187_297# N_A_1187_297#_M1001_d
+ N_A_1187_297#_M1011_d N_A_1187_297#_M1022_d N_A_1187_297#_M1025_s
+ N_A_1187_297#_M1032_s N_A_1187_297#_c_1044_n N_A_1187_297#_c_1052_n
+ N_A_1187_297#_c_1045_n N_A_1187_297#_c_1102_n N_A_1187_297#_c_1054_n
+ N_A_1187_297#_c_1046_n N_A_1187_297#_c_1079_n N_A_1187_297#_c_1047_n
+ N_A_1187_297#_c_1083_n N_A_1187_297#_c_1048_n N_A_1187_297#_c_1049_n
+ N_A_1187_297#_c_1050_n N_A_1187_297#_c_1089_n N_A_1187_297#_c_1051_n
+ PM_SKY130_FD_SC_HDLL__NOR4BB_4%A_1187_297#
x_PM_SKY130_FD_SC_HDLL__NOR4BB_4%VGND N_VGND_M1006_d N_VGND_M1007_d
+ N_VGND_M1019_d N_VGND_M1028_d N_VGND_M1005_s N_VGND_M1015_s N_VGND_M1014_s
+ N_VGND_M1033_s N_VGND_M1021_s N_VGND_M1034_s N_VGND_c_1107_n N_VGND_c_1108_n
+ N_VGND_c_1109_n N_VGND_c_1110_n N_VGND_c_1111_n N_VGND_c_1112_n
+ N_VGND_c_1113_n N_VGND_c_1114_n N_VGND_c_1115_n N_VGND_c_1116_n
+ N_VGND_c_1117_n N_VGND_c_1118_n N_VGND_c_1119_n N_VGND_c_1120_n
+ N_VGND_c_1121_n N_VGND_c_1122_n N_VGND_c_1123_n N_VGND_c_1124_n
+ N_VGND_c_1125_n N_VGND_c_1126_n N_VGND_c_1127_n N_VGND_c_1128_n
+ N_VGND_c_1129_n N_VGND_c_1130_n VGND N_VGND_c_1131_n N_VGND_c_1132_n
+ N_VGND_c_1133_n N_VGND_c_1134_n N_VGND_c_1135_n VGND
+ PM_SKY130_FD_SC_HDLL__NOR4BB_4%VGND
cc_1 VNB N_C_N_c_152_n 0.0218983f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_2 VNB C_N 0.00888669f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_C_N_c_154_n 0.0397621f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_4 VNB N_D_N_c_178_n 0.0201641f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_5 VNB D_N 0.0017601f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_6 VNB N_D_N_c_180_n 0.0375609f $X=-0.19 $Y=-0.24 $X2=0.28 $Y2=1.16
cc_7 VNB N_A_207_47#_c_218_n 0.0196746f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_8 VNB N_A_207_47#_c_219_n 0.0167613f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.202
cc_9 VNB N_A_207_47#_c_220_n 0.0171746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_207_47#_c_221_n 0.0165308f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_207_47#_c_222_n 0.0059198f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_207_47#_c_223_n 0.0082966f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_207_47#_c_224_n 0.00237058f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_207_47#_c_225_n 0.00460374f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_207_47#_c_226_n 0.00129226f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_207_47#_c_227_n 0.00655567f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_207_47#_c_228_n 0.00210943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_207_47#_c_229_n 0.0773793f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_297#_c_342_n 0.0164668f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_20 VNB N_A_27_297#_c_343_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.202
cc_21 VNB N_A_27_297#_c_344_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_297#_c_345_n 0.0224149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_297#_c_346_n 0.0189957f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_297#_c_347_n 9.49372e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_297#_c_348_n 0.00982927f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_297#_c_349_n 0.00754719f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_297#_c_350_n 0.00268481f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_27_297#_c_351_n 0.0022324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_27_297#_c_352_n 0.0799867f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_B_c_491_n 0.021971f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_31 VNB N_B_c_492_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_32 VNB N_B_c_493_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.202
cc_33 VNB N_B_c_494_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_B_c_495_n 0.0159176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_B_c_496_n 0.0801694f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_c_568_n 0.0164943f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_37 VNB N_A_c_569_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_38 VNB N_A_c_570_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.202
cc_39 VNB N_A_c_571_n 0.0223809f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_c_572_n 0.0184554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_c_573_n 0.0801694f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VPWR_c_637_n 0.421552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_Y_c_791_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_Y_c_792_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_Y_c_793_n 9.16142e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_Y_c_794_n 0.00578238f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_Y_c_795_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_Y_c_796_n 0.00921701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_Y_c_797_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_Y_c_798_n 0.00447396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_Y_c_799_n 0.00528609f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_Y_c_800_n 0.00212267f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_Y_c_801_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_Y_c_802_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_Y_c_803_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_Y_c_804_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_Y_c_805_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1107_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1108_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1109_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1110_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1111_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1112_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1113_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1114_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1115_n 0.0109994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1116_n 0.0335222f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1117_n 0.022483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1118_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1119_n 0.0198149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1120_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1121_n 0.0192905f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1122_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1123_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1124_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1125_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1126_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1127_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1128_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1129_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1130_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1131_n 0.0201171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1132_n 0.0223506f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1133_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1134_n 0.0208752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1135_n 0.470539f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VPB N_C_N_c_155_n 0.0207484f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_88 VPB C_N 0.00503237f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_89 VPB N_C_N_c_154_n 0.0168807f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_90 VPB N_D_N_c_181_n 0.0195915f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_91 VPB D_N 2.38784e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_92 VPB N_D_N_c_180_n 0.0156566f $X=-0.19 $Y=1.305 $X2=0.28 $Y2=1.16
cc_93 VPB N_A_207_47#_c_230_n 0.0189193f $X=-0.19 $Y=1.305 $X2=0.28 $Y2=1.16
cc_94 VPB N_A_207_47#_c_231_n 0.015551f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_207_47#_c_232_n 0.015551f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_207_47#_c_233_n 0.0160334f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_207_47#_c_234_n 0.00716661f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_207_47#_c_226_n 0.0055574f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_207_47#_c_229_n 0.0453205f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_27_297#_c_353_n 0.0159278f $X=-0.19 $Y=1.305 $X2=0.28 $Y2=1.16
cc_101 VPB N_A_27_297#_c_354_n 0.015972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_27_297#_c_355_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_27_297#_c_356_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_27_297#_c_357_n 0.0165958f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_27_297#_c_349_n 0.00353117f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_27_297#_c_359_n 0.00813339f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_27_297#_c_360_n 0.00114801f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_27_297#_c_361_n 0.0223622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_27_297#_c_352_n 0.0495373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_B_c_497_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_111 VPB N_B_c_498_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.28 $Y2=1.16
cc_112 VPB N_B_c_499_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_B_c_500_n 0.0164231f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_B_c_496_n 0.0492916f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_c_574_n 0.0161064f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_116 VPB N_A_c_575_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.28 $Y2=1.16
cc_117 VPB N_A_c_576_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_c_577_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_c_573_n 0.048391f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_638_n 4.89699e-19 $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_121 VPB N_VPWR_c_639_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_640_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_641_n 0.169989f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_642_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_643_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_644_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_645_n 0.0147956f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_646_n 0.0197239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_637_n 0.0578601f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_648_n 0.00502902f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_331_297#_c_743_n 0.00492884f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_331_297#_c_744_n 0.00166712f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_331_297#_c_745_n 0.00452881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_Y_c_793_n 8.39856e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_Y_c_807_n 0.00497668f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_797_297#_c_983_n 0.00193318f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_137 VPB N_A_797_297#_c_984_n 0.0181179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_797_297#_c_985_n 0.00193318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_797_297#_c_986_n 0.00148765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_797_297#_c_987_n 0.00149756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_797_297#_c_988_n 0.00149756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_797_297#_c_989_n 0.00174485f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_1187_297#_c_1044_n 0.00518462f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_1187_297#_c_1045_n 0.0019907f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_1187_297#_c_1046_n 0.00416269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_1187_297#_c_1047_n 0.00201678f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_1187_297#_c_1048_n 0.00196267f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_1187_297#_c_1049_n 0.010274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_1187_297#_c_1050_n 0.0327764f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_1187_297#_c_1051_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 N_C_N_c_152_n N_D_N_c_178_n 0.0206501f $X=0.54 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_152 N_C_N_c_155_n N_D_N_c_181_n 0.033124f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_153 N_C_N_c_154_n N_D_N_c_180_n 0.0206501f $X=0.515 $Y=1.202 $X2=0 $Y2=0
cc_154 N_C_N_c_152_n N_A_207_47#_c_222_n 5.41954e-19 $X=0.54 $Y=0.995 $X2=0
+ $Y2=0
cc_155 N_C_N_c_152_n N_A_27_297#_c_347_n 0.0119068f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_156 N_C_N_c_154_n N_A_27_297#_c_347_n 6.70277e-19 $X=0.515 $Y=1.202 $X2=0
+ $Y2=0
cc_157 C_N N_A_27_297#_c_348_n 0.0268296f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_158 N_C_N_c_154_n N_A_27_297#_c_348_n 0.00773312f $X=0.515 $Y=1.202 $X2=0
+ $Y2=0
cc_159 N_C_N_c_155_n N_A_27_297#_c_349_n 0.00299893f $X=0.515 $Y=1.41 $X2=0
+ $Y2=0
cc_160 N_C_N_c_152_n N_A_27_297#_c_349_n 0.00802928f $X=0.54 $Y=0.995 $X2=0
+ $Y2=0
cc_161 C_N N_A_27_297#_c_349_n 0.0179248f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_162 N_C_N_c_155_n N_A_27_297#_c_361_n 0.022051f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_163 C_N N_A_27_297#_c_361_n 0.0254007f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_164 N_C_N_c_154_n N_A_27_297#_c_361_n 0.00173959f $X=0.515 $Y=1.202 $X2=0
+ $Y2=0
cc_165 N_C_N_c_155_n N_VPWR_c_638_n 0.0115795f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_166 N_C_N_c_155_n N_VPWR_c_645_n 0.00315243f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_167 N_C_N_c_155_n N_VPWR_c_637_n 0.00471211f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_168 N_C_N_c_152_n N_VGND_c_1107_n 0.00268723f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_169 N_C_N_c_152_n N_VGND_c_1132_n 0.00437852f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_170 N_C_N_c_152_n N_VGND_c_1135_n 0.00692883f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_171 N_D_N_c_178_n N_A_207_47#_c_222_n 0.00655146f $X=0.96 $Y=0.995 $X2=0
+ $Y2=0
cc_172 N_D_N_c_181_n N_A_207_47#_c_234_n 0.00435012f $X=0.985 $Y=1.41 $X2=0
+ $Y2=0
cc_173 D_N N_A_207_47#_c_234_n 0.0220686f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_174 N_D_N_c_180_n N_A_207_47#_c_234_n 0.00643511f $X=0.985 $Y=1.202 $X2=0
+ $Y2=0
cc_175 D_N N_A_207_47#_c_223_n 7.38065e-19 $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_176 N_D_N_c_178_n N_A_207_47#_c_224_n 0.00264289f $X=0.96 $Y=0.995 $X2=0
+ $Y2=0
cc_177 D_N N_A_207_47#_c_224_n 0.031193f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_178 N_D_N_c_180_n N_A_207_47#_c_224_n 0.00914167f $X=0.985 $Y=1.202 $X2=0
+ $Y2=0
cc_179 N_D_N_c_178_n N_A_207_47#_c_225_n 0.00209138f $X=0.96 $Y=0.995 $X2=0
+ $Y2=0
cc_180 N_D_N_c_180_n N_A_207_47#_c_225_n 0.00195033f $X=0.985 $Y=1.202 $X2=0
+ $Y2=0
cc_181 N_D_N_c_181_n N_A_207_47#_c_226_n 0.00246835f $X=0.985 $Y=1.41 $X2=0
+ $Y2=0
cc_182 D_N N_A_207_47#_c_226_n 0.0063378f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_183 N_D_N_c_180_n N_A_207_47#_c_226_n 0.00246283f $X=0.985 $Y=1.202 $X2=0
+ $Y2=0
cc_184 D_N N_A_207_47#_c_228_n 0.0151968f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_185 N_D_N_c_180_n N_A_207_47#_c_228_n 7.69385e-19 $X=0.985 $Y=1.202 $X2=0
+ $Y2=0
cc_186 D_N N_A_207_47#_c_229_n 4.45324e-19 $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_187 N_D_N_c_180_n N_A_207_47#_c_229_n 0.00576083f $X=0.985 $Y=1.202 $X2=0
+ $Y2=0
cc_188 N_D_N_c_178_n N_A_27_297#_c_347_n 7.36469e-19 $X=0.96 $Y=0.995 $X2=0
+ $Y2=0
cc_189 N_D_N_c_178_n N_A_27_297#_c_349_n 0.00836752f $X=0.96 $Y=0.995 $X2=0
+ $Y2=0
cc_190 N_D_N_c_181_n N_A_27_297#_c_349_n 0.00299893f $X=0.985 $Y=1.41 $X2=0
+ $Y2=0
cc_191 D_N N_A_27_297#_c_349_n 0.0189691f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_192 N_D_N_c_181_n N_A_27_297#_c_359_n 0.0188628f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_193 N_D_N_c_181_n N_A_27_297#_c_361_n 0.0068236f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_194 N_D_N_c_181_n N_VPWR_c_638_n 0.016743f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_195 N_D_N_c_181_n N_VPWR_c_641_n 0.00458874f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_196 N_D_N_c_181_n N_VPWR_c_637_n 0.00661886f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_197 N_D_N_c_181_n N_A_331_297#_c_743_n 0.00704772f $X=0.985 $Y=1.41 $X2=0
+ $Y2=0
cc_198 N_D_N_c_178_n N_VGND_c_1107_n 0.00268723f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_199 N_D_N_c_178_n N_VGND_c_1108_n 0.0016715f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_200 N_D_N_c_178_n N_VGND_c_1117_n 0.00541359f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_201 N_D_N_c_178_n N_VGND_c_1135_n 0.0108548f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_207_47#_c_221_n N_A_27_297#_c_342_n 0.0229083f $X=3.45 $Y=0.995 $X2=0
+ $Y2=0
cc_203 N_A_207_47#_c_233_n N_A_27_297#_c_353_n 0.0345562f $X=3.425 $Y=1.41 $X2=0
+ $Y2=0
cc_204 N_A_207_47#_c_224_n N_A_27_297#_c_347_n 0.00719342f $X=1.385 $Y=0.82
+ $X2=0 $Y2=0
cc_205 N_A_207_47#_c_224_n N_A_27_297#_c_349_n 7.61274e-19 $X=1.385 $Y=0.82
+ $X2=0 $Y2=0
cc_206 N_A_207_47#_M1026_d N_A_27_297#_c_359_n 0.00751209f $X=1.075 $Y=1.485
+ $X2=0 $Y2=0
cc_207 N_A_207_47#_c_230_n N_A_27_297#_c_359_n 0.0141027f $X=2.015 $Y=1.41 $X2=0
+ $Y2=0
cc_208 N_A_207_47#_c_231_n N_A_27_297#_c_359_n 0.0118884f $X=2.485 $Y=1.41 $X2=0
+ $Y2=0
cc_209 N_A_207_47#_c_232_n N_A_27_297#_c_359_n 0.0118884f $X=2.955 $Y=1.41 $X2=0
+ $Y2=0
cc_210 N_A_207_47#_c_233_n N_A_27_297#_c_359_n 0.0142709f $X=3.425 $Y=1.41 $X2=0
+ $Y2=0
cc_211 N_A_207_47#_c_234_n N_A_27_297#_c_359_n 0.0506754f $X=1.565 $Y=1.62 $X2=0
+ $Y2=0
cc_212 N_A_207_47#_c_227_n N_A_27_297#_c_359_n 0.00497139f $X=2.88 $Y=1.16 $X2=0
+ $Y2=0
cc_213 N_A_207_47#_c_229_n N_A_27_297#_c_359_n 3.28191e-19 $X=3.425 $Y=1.202
+ $X2=0 $Y2=0
cc_214 N_A_207_47#_c_233_n N_A_27_297#_c_360_n 0.00566158f $X=3.425 $Y=1.41
+ $X2=0 $Y2=0
cc_215 N_A_207_47#_c_229_n N_A_27_297#_c_360_n 8.9079e-19 $X=3.425 $Y=1.202
+ $X2=0 $Y2=0
cc_216 N_A_207_47#_c_229_n N_A_27_297#_c_350_n 0.00193165f $X=3.425 $Y=1.202
+ $X2=0 $Y2=0
cc_217 N_A_207_47#_c_234_n N_A_27_297#_c_361_n 0.0146837f $X=1.565 $Y=1.62 $X2=0
+ $Y2=0
cc_218 N_A_207_47#_c_229_n N_A_27_297#_c_352_n 0.0229083f $X=3.425 $Y=1.202
+ $X2=0 $Y2=0
cc_219 N_A_207_47#_c_230_n N_VPWR_c_641_n 0.00429453f $X=2.015 $Y=1.41 $X2=0
+ $Y2=0
cc_220 N_A_207_47#_c_231_n N_VPWR_c_641_n 0.00429453f $X=2.485 $Y=1.41 $X2=0
+ $Y2=0
cc_221 N_A_207_47#_c_232_n N_VPWR_c_641_n 0.00429453f $X=2.955 $Y=1.41 $X2=0
+ $Y2=0
cc_222 N_A_207_47#_c_233_n N_VPWR_c_641_n 0.00429453f $X=3.425 $Y=1.41 $X2=0
+ $Y2=0
cc_223 N_A_207_47#_M1026_d N_VPWR_c_637_n 0.00357409f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_224 N_A_207_47#_c_230_n N_VPWR_c_637_n 0.00734734f $X=2.015 $Y=1.41 $X2=0
+ $Y2=0
cc_225 N_A_207_47#_c_231_n N_VPWR_c_637_n 0.00606499f $X=2.485 $Y=1.41 $X2=0
+ $Y2=0
cc_226 N_A_207_47#_c_232_n N_VPWR_c_637_n 0.00606499f $X=2.955 $Y=1.41 $X2=0
+ $Y2=0
cc_227 N_A_207_47#_c_233_n N_VPWR_c_637_n 0.00609021f $X=3.425 $Y=1.41 $X2=0
+ $Y2=0
cc_228 N_A_207_47#_c_234_n N_A_331_297#_M1000_s 0.003221f $X=1.565 $Y=1.62
+ $X2=-0.19 $Y2=-0.24
cc_229 N_A_207_47#_c_226_n N_A_331_297#_M1000_s 6.57336e-19 $X=1.65 $Y=1.535
+ $X2=-0.19 $Y2=-0.24
cc_230 N_A_207_47#_c_230_n N_A_331_297#_c_743_n 0.0112654f $X=2.015 $Y=1.41
+ $X2=0 $Y2=0
cc_231 N_A_207_47#_c_231_n N_A_331_297#_c_743_n 0.0112654f $X=2.485 $Y=1.41
+ $X2=0 $Y2=0
cc_232 N_A_207_47#_c_232_n N_A_331_297#_c_743_n 0.0112654f $X=2.955 $Y=1.41
+ $X2=0 $Y2=0
cc_233 N_A_207_47#_c_233_n N_A_331_297#_c_743_n 0.0112515f $X=3.425 $Y=1.41
+ $X2=0 $Y2=0
cc_234 N_A_207_47#_c_218_n N_Y_c_808_n 0.00730874f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A_207_47#_c_219_n N_Y_c_808_n 0.00686626f $X=2.46 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A_207_47#_c_220_n N_Y_c_808_n 5.45498e-19 $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A_207_47#_c_222_n N_Y_c_808_n 0.00495038f $X=1.22 $Y=0.39 $X2=0 $Y2=0
cc_238 N_A_207_47#_c_219_n N_Y_c_791_n 0.00901745f $X=2.46 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A_207_47#_c_220_n N_Y_c_791_n 0.00901745f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A_207_47#_c_227_n N_Y_c_791_n 0.0392656f $X=2.88 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A_207_47#_c_229_n N_Y_c_791_n 0.00345541f $X=3.425 $Y=1.202 $X2=0 $Y2=0
cc_242 N_A_207_47#_c_218_n N_Y_c_792_n 0.00334463f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A_207_47#_c_219_n N_Y_c_792_n 0.00116636f $X=2.46 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_207_47#_c_222_n N_Y_c_792_n 2.87375e-19 $X=1.22 $Y=0.39 $X2=0 $Y2=0
cc_245 N_A_207_47#_c_223_n N_Y_c_792_n 0.00961296f $X=1.565 $Y=0.82 $X2=0 $Y2=0
cc_246 N_A_207_47#_c_227_n N_Y_c_792_n 0.030274f $X=2.88 $Y=1.16 $X2=0 $Y2=0
cc_247 N_A_207_47#_c_229_n N_Y_c_792_n 0.00358305f $X=3.425 $Y=1.202 $X2=0 $Y2=0
cc_248 N_A_207_47#_c_219_n N_Y_c_822_n 5.24597e-19 $X=2.46 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A_207_47#_c_220_n N_Y_c_822_n 0.00651696f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A_207_47#_c_220_n N_Y_c_793_n 0.00172173f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A_207_47#_c_221_n N_Y_c_793_n 0.00246161f $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A_207_47#_c_227_n N_Y_c_793_n 0.0127974f $X=2.88 $Y=1.16 $X2=0 $Y2=0
cc_253 N_A_207_47#_c_229_n N_Y_c_793_n 0.0234004f $X=3.425 $Y=1.202 $X2=0 $Y2=0
cc_254 N_A_207_47#_c_221_n N_Y_c_794_n 0.00969879f $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A_207_47#_c_221_n N_Y_c_829_n 5.32212e-19 $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_256 N_A_207_47#_c_220_n N_Y_c_800_n 0.00119564f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_257 N_A_207_47#_c_221_n N_Y_c_800_n 0.00277851f $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_258 N_A_207_47#_c_227_n N_Y_c_800_n 0.00951185f $X=2.88 $Y=1.16 $X2=0 $Y2=0
cc_259 N_A_207_47#_c_229_n N_Y_c_800_n 0.00530543f $X=3.425 $Y=1.202 $X2=0 $Y2=0
cc_260 N_A_207_47#_c_230_n N_Y_c_807_n 0.01166f $X=2.015 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A_207_47#_c_231_n N_Y_c_807_n 0.0142715f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A_207_47#_c_232_n N_Y_c_807_n 0.0142715f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A_207_47#_c_233_n N_Y_c_807_n 0.00725439f $X=3.425 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A_207_47#_c_234_n N_Y_c_807_n 0.0127689f $X=1.565 $Y=1.62 $X2=0 $Y2=0
cc_265 N_A_207_47#_c_226_n N_Y_c_807_n 0.00815109f $X=1.65 $Y=1.535 $X2=0 $Y2=0
cc_266 N_A_207_47#_c_227_n N_Y_c_807_n 0.0841619f $X=2.88 $Y=1.16 $X2=0 $Y2=0
cc_267 N_A_207_47#_c_229_n N_Y_c_807_n 0.0224318f $X=3.425 $Y=1.202 $X2=0 $Y2=0
cc_268 N_A_207_47#_c_223_n N_VGND_M1007_d 0.00356387f $X=1.565 $Y=0.82 $X2=0
+ $Y2=0
cc_269 N_A_207_47#_c_218_n N_VGND_c_1108_n 0.00438629f $X=1.99 $Y=0.995 $X2=0
+ $Y2=0
cc_270 N_A_207_47#_c_222_n N_VGND_c_1108_n 0.01542f $X=1.22 $Y=0.39 $X2=0 $Y2=0
cc_271 N_A_207_47#_c_223_n N_VGND_c_1108_n 0.00321628f $X=1.565 $Y=0.82 $X2=0
+ $Y2=0
cc_272 N_A_207_47#_c_227_n N_VGND_c_1108_n 0.00460552f $X=2.88 $Y=1.16 $X2=0
+ $Y2=0
cc_273 N_A_207_47#_c_219_n N_VGND_c_1109_n 0.00379224f $X=2.46 $Y=0.995 $X2=0
+ $Y2=0
cc_274 N_A_207_47#_c_220_n N_VGND_c_1109_n 0.00276126f $X=2.93 $Y=0.995 $X2=0
+ $Y2=0
cc_275 N_A_207_47#_c_221_n N_VGND_c_1110_n 0.00268723f $X=3.45 $Y=0.995 $X2=0
+ $Y2=0
cc_276 N_A_207_47#_c_222_n N_VGND_c_1117_n 0.0244796f $X=1.22 $Y=0.39 $X2=0
+ $Y2=0
cc_277 N_A_207_47#_c_223_n N_VGND_c_1117_n 0.00480319f $X=1.565 $Y=0.82 $X2=0
+ $Y2=0
cc_278 N_A_207_47#_c_218_n N_VGND_c_1119_n 0.00541359f $X=1.99 $Y=0.995 $X2=0
+ $Y2=0
cc_279 N_A_207_47#_c_219_n N_VGND_c_1119_n 0.00423334f $X=2.46 $Y=0.995 $X2=0
+ $Y2=0
cc_280 N_A_207_47#_c_220_n N_VGND_c_1121_n 0.00423334f $X=2.93 $Y=0.995 $X2=0
+ $Y2=0
cc_281 N_A_207_47#_c_221_n N_VGND_c_1121_n 0.00437798f $X=3.45 $Y=0.995 $X2=0
+ $Y2=0
cc_282 N_A_207_47#_M1003_d N_VGND_c_1135_n 0.00250309f $X=1.035 $Y=0.235 $X2=0
+ $Y2=0
cc_283 N_A_207_47#_c_218_n N_VGND_c_1135_n 0.0109546f $X=1.99 $Y=0.995 $X2=0
+ $Y2=0
cc_284 N_A_207_47#_c_219_n N_VGND_c_1135_n 0.006093f $X=2.46 $Y=0.995 $X2=0
+ $Y2=0
cc_285 N_A_207_47#_c_220_n N_VGND_c_1135_n 0.00608558f $X=2.93 $Y=0.995 $X2=0
+ $Y2=0
cc_286 N_A_207_47#_c_221_n N_VGND_c_1135_n 0.00615524f $X=3.45 $Y=0.995 $X2=0
+ $Y2=0
cc_287 N_A_207_47#_c_222_n N_VGND_c_1135_n 0.0143352f $X=1.22 $Y=0.39 $X2=0
+ $Y2=0
cc_288 N_A_207_47#_c_223_n N_VGND_c_1135_n 0.00855541f $X=1.565 $Y=0.82 $X2=0
+ $Y2=0
cc_289 N_A_27_297#_c_351_n N_B_c_495_n 0.0140827f $X=5.19 $Y=1.16 $X2=0 $Y2=0
cc_290 N_A_27_297#_c_352_n N_B_c_495_n 0.00155889f $X=5.305 $Y=1.202 $X2=0 $Y2=0
cc_291 N_A_27_297#_c_349_n N_VPWR_M1002_d 0.00170744f $X=0.75 $Y=1.535 $X2=-0.19
+ $Y2=-0.24
cc_292 N_A_27_297#_c_361_n N_VPWR_M1002_d 0.00628473f $X=0.835 $Y=1.79 $X2=-0.19
+ $Y2=-0.24
cc_293 N_A_27_297#_c_357_n N_VPWR_c_638_n 0.0193679f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_294 N_A_27_297#_c_361_n N_VPWR_c_638_n 0.0211498f $X=0.835 $Y=1.79 $X2=0
+ $Y2=0
cc_295 N_A_27_297#_c_353_n N_VPWR_c_641_n 0.00429453f $X=3.895 $Y=1.41 $X2=0
+ $Y2=0
cc_296 N_A_27_297#_c_354_n N_VPWR_c_641_n 0.00429453f $X=4.365 $Y=1.41 $X2=0
+ $Y2=0
cc_297 N_A_27_297#_c_355_n N_VPWR_c_641_n 0.00429453f $X=4.835 $Y=1.41 $X2=0
+ $Y2=0
cc_298 N_A_27_297#_c_356_n N_VPWR_c_641_n 0.00429453f $X=5.305 $Y=1.41 $X2=0
+ $Y2=0
cc_299 N_A_27_297#_c_359_n N_VPWR_c_641_n 0.0108294f $X=3.655 $Y=1.96 $X2=0
+ $Y2=0
cc_300 N_A_27_297#_c_357_n N_VPWR_c_645_n 0.0189422f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_301 N_A_27_297#_c_361_n N_VPWR_c_645_n 0.00234071f $X=0.835 $Y=1.79 $X2=0
+ $Y2=0
cc_302 N_A_27_297#_M1002_s N_VPWR_c_637_n 0.00259298f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_303 N_A_27_297#_c_353_n N_VPWR_c_637_n 0.00609021f $X=3.895 $Y=1.41 $X2=0
+ $Y2=0
cc_304 N_A_27_297#_c_354_n N_VPWR_c_637_n 0.00606499f $X=4.365 $Y=1.41 $X2=0
+ $Y2=0
cc_305 N_A_27_297#_c_355_n N_VPWR_c_637_n 0.00606499f $X=4.835 $Y=1.41 $X2=0
+ $Y2=0
cc_306 N_A_27_297#_c_356_n N_VPWR_c_637_n 0.00734734f $X=5.305 $Y=1.41 $X2=0
+ $Y2=0
cc_307 N_A_27_297#_c_357_n N_VPWR_c_637_n 0.0105763f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_308 N_A_27_297#_c_359_n N_VPWR_c_637_n 0.0219165f $X=3.655 $Y=1.96 $X2=0
+ $Y2=0
cc_309 N_A_27_297#_c_361_n N_VPWR_c_637_n 0.00603004f $X=0.835 $Y=1.79 $X2=0
+ $Y2=0
cc_310 N_A_27_297#_c_359_n N_A_331_297#_M1000_s 0.00659249f $X=3.655 $Y=1.96
+ $X2=-0.19 $Y2=-0.24
cc_311 N_A_27_297#_c_359_n N_A_331_297#_M1010_s 0.00350871f $X=3.655 $Y=1.96
+ $X2=0 $Y2=0
cc_312 N_A_27_297#_c_359_n N_A_331_297#_M1029_s 0.00496372f $X=3.655 $Y=1.96
+ $X2=0 $Y2=0
cc_313 N_A_27_297#_c_360_n N_A_331_297#_M1029_s 0.00392753f $X=3.74 $Y=1.875
+ $X2=0 $Y2=0
cc_314 N_A_27_297#_c_359_n N_A_331_297#_c_743_n 0.118574f $X=3.655 $Y=1.96 $X2=0
+ $Y2=0
cc_315 N_A_27_297#_c_353_n N_A_331_297#_c_758_n 0.0129846f $X=3.895 $Y=1.41
+ $X2=0 $Y2=0
cc_316 N_A_27_297#_c_354_n N_A_331_297#_c_758_n 0.01161f $X=4.365 $Y=1.41 $X2=0
+ $Y2=0
cc_317 N_A_27_297#_c_355_n N_A_331_297#_c_744_n 0.01161f $X=4.835 $Y=1.41 $X2=0
+ $Y2=0
cc_318 N_A_27_297#_c_356_n N_A_331_297#_c_744_n 0.01161f $X=5.305 $Y=1.41 $X2=0
+ $Y2=0
cc_319 N_A_27_297#_c_353_n N_A_331_297#_c_762_n 0.002273f $X=3.895 $Y=1.41 $X2=0
+ $Y2=0
cc_320 N_A_27_297#_c_354_n N_A_331_297#_c_762_n 2.34252e-19 $X=4.365 $Y=1.41
+ $X2=0 $Y2=0
cc_321 N_A_27_297#_c_359_n N_Y_M1000_d 0.00350871f $X=3.655 $Y=1.96 $X2=0 $Y2=0
cc_322 N_A_27_297#_c_359_n N_Y_M1016_d 0.00349883f $X=3.655 $Y=1.96 $X2=0 $Y2=0
cc_323 N_A_27_297#_c_342_n N_Y_c_793_n 9.68601e-19 $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_324 N_A_27_297#_c_360_n N_Y_c_793_n 0.00758122f $X=3.74 $Y=1.875 $X2=0 $Y2=0
cc_325 N_A_27_297#_c_350_n N_Y_c_793_n 0.0139762f $X=3.825 $Y=1.18 $X2=0 $Y2=0
cc_326 N_A_27_297#_c_352_n N_Y_c_793_n 3.02604e-19 $X=5.305 $Y=1.202 $X2=0 $Y2=0
cc_327 N_A_27_297#_c_342_n N_Y_c_794_n 0.00865562f $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_328 N_A_27_297#_c_350_n N_Y_c_794_n 0.014165f $X=3.825 $Y=1.18 $X2=0 $Y2=0
cc_329 N_A_27_297#_c_351_n N_Y_c_794_n 0.00615875f $X=5.19 $Y=1.16 $X2=0 $Y2=0
cc_330 N_A_27_297#_c_342_n N_Y_c_829_n 0.00644736f $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_331 N_A_27_297#_c_343_n N_Y_c_829_n 0.00686626f $X=4.34 $Y=0.995 $X2=0 $Y2=0
cc_332 N_A_27_297#_c_344_n N_Y_c_829_n 5.45498e-19 $X=4.81 $Y=0.995 $X2=0 $Y2=0
cc_333 N_A_27_297#_c_343_n N_Y_c_795_n 0.00901745f $X=4.34 $Y=0.995 $X2=0 $Y2=0
cc_334 N_A_27_297#_c_344_n N_Y_c_795_n 0.00901745f $X=4.81 $Y=0.995 $X2=0 $Y2=0
cc_335 N_A_27_297#_c_351_n N_Y_c_795_n 0.0398926f $X=5.19 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A_27_297#_c_352_n N_Y_c_795_n 0.00345541f $X=5.305 $Y=1.202 $X2=0 $Y2=0
cc_337 N_A_27_297#_c_343_n N_Y_c_858_n 5.24597e-19 $X=4.34 $Y=0.995 $X2=0 $Y2=0
cc_338 N_A_27_297#_c_344_n N_Y_c_858_n 0.00651696f $X=4.81 $Y=0.995 $X2=0 $Y2=0
cc_339 N_A_27_297#_c_345_n N_Y_c_796_n 0.01289f $X=5.33 $Y=0.995 $X2=0 $Y2=0
cc_340 N_A_27_297#_c_351_n N_Y_c_796_n 0.0118017f $X=5.19 $Y=1.16 $X2=0 $Y2=0
cc_341 N_A_27_297#_c_353_n N_Y_c_807_n 2.61756e-19 $X=3.895 $Y=1.41 $X2=0 $Y2=0
cc_342 N_A_27_297#_c_359_n N_Y_c_807_n 0.0845095f $X=3.655 $Y=1.96 $X2=0 $Y2=0
cc_343 N_A_27_297#_c_360_n N_Y_c_807_n 0.0187595f $X=3.74 $Y=1.875 $X2=0 $Y2=0
cc_344 N_A_27_297#_c_342_n N_Y_c_801_n 0.00116636f $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_345 N_A_27_297#_c_343_n N_Y_c_801_n 0.00116636f $X=4.34 $Y=0.995 $X2=0 $Y2=0
cc_346 N_A_27_297#_c_351_n N_Y_c_801_n 0.0307014f $X=5.19 $Y=1.16 $X2=0 $Y2=0
cc_347 N_A_27_297#_c_352_n N_Y_c_801_n 0.00358305f $X=5.305 $Y=1.202 $X2=0 $Y2=0
cc_348 N_A_27_297#_c_344_n N_Y_c_802_n 0.00119564f $X=4.81 $Y=0.995 $X2=0 $Y2=0
cc_349 N_A_27_297#_c_351_n N_Y_c_802_n 0.030835f $X=5.19 $Y=1.16 $X2=0 $Y2=0
cc_350 N_A_27_297#_c_352_n N_Y_c_802_n 0.00486271f $X=5.305 $Y=1.202 $X2=0 $Y2=0
cc_351 N_A_27_297#_c_354_n N_A_797_297#_c_983_n 0.0127983f $X=4.365 $Y=1.41
+ $X2=0 $Y2=0
cc_352 N_A_27_297#_c_355_n N_A_797_297#_c_983_n 0.0128365f $X=4.835 $Y=1.41
+ $X2=0 $Y2=0
cc_353 N_A_27_297#_c_351_n N_A_797_297#_c_983_n 0.0486996f $X=5.19 $Y=1.16 $X2=0
+ $Y2=0
cc_354 N_A_27_297#_c_352_n N_A_797_297#_c_983_n 0.00864922f $X=5.305 $Y=1.202
+ $X2=0 $Y2=0
cc_355 N_A_27_297#_c_356_n N_A_797_297#_c_984_n 0.0148794f $X=5.305 $Y=1.41
+ $X2=0 $Y2=0
cc_356 N_A_27_297#_c_351_n N_A_797_297#_c_984_n 0.0145434f $X=5.19 $Y=1.16 $X2=0
+ $Y2=0
cc_357 N_A_27_297#_c_352_n N_A_797_297#_c_984_n 8.84531e-19 $X=5.305 $Y=1.202
+ $X2=0 $Y2=0
cc_358 N_A_27_297#_c_353_n N_A_797_297#_c_986_n 9.55966e-19 $X=3.895 $Y=1.41
+ $X2=0 $Y2=0
cc_359 N_A_27_297#_c_359_n N_A_797_297#_c_986_n 0.0111041f $X=3.655 $Y=1.96
+ $X2=0 $Y2=0
cc_360 N_A_27_297#_c_360_n N_A_797_297#_c_986_n 0.0256374f $X=3.74 $Y=1.875
+ $X2=0 $Y2=0
cc_361 N_A_27_297#_c_351_n N_A_797_297#_c_986_n 0.0171572f $X=5.19 $Y=1.16 $X2=0
+ $Y2=0
cc_362 N_A_27_297#_c_352_n N_A_797_297#_c_986_n 0.00545262f $X=5.305 $Y=1.202
+ $X2=0 $Y2=0
cc_363 N_A_27_297#_c_351_n N_A_797_297#_c_987_n 0.0204252f $X=5.19 $Y=1.16 $X2=0
+ $Y2=0
cc_364 N_A_27_297#_c_352_n N_A_797_297#_c_987_n 0.00634604f $X=5.305 $Y=1.202
+ $X2=0 $Y2=0
cc_365 N_A_27_297#_c_347_n N_VGND_M1006_d 0.00195f $X=0.665 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_366 N_A_27_297#_c_347_n N_VGND_c_1107_n 0.0134908f $X=0.665 $Y=0.81 $X2=0
+ $Y2=0
cc_367 N_A_27_297#_c_342_n N_VGND_c_1110_n 0.00268723f $X=3.87 $Y=0.995 $X2=0
+ $Y2=0
cc_368 N_A_27_297#_c_343_n N_VGND_c_1111_n 0.00379224f $X=4.34 $Y=0.995 $X2=0
+ $Y2=0
cc_369 N_A_27_297#_c_344_n N_VGND_c_1111_n 0.00276126f $X=4.81 $Y=0.995 $X2=0
+ $Y2=0
cc_370 N_A_27_297#_c_342_n N_VGND_c_1123_n 0.00423334f $X=3.87 $Y=0.995 $X2=0
+ $Y2=0
cc_371 N_A_27_297#_c_343_n N_VGND_c_1123_n 0.00423334f $X=4.34 $Y=0.995 $X2=0
+ $Y2=0
cc_372 N_A_27_297#_c_346_n N_VGND_c_1132_n 0.0238935f $X=0.28 $Y=0.39 $X2=0
+ $Y2=0
cc_373 N_A_27_297#_c_347_n N_VGND_c_1132_n 0.00253779f $X=0.665 $Y=0.81 $X2=0
+ $Y2=0
cc_374 N_A_27_297#_c_344_n N_VGND_c_1133_n 0.00423334f $X=4.81 $Y=0.995 $X2=0
+ $Y2=0
cc_375 N_A_27_297#_c_345_n N_VGND_c_1133_n 0.00437852f $X=5.33 $Y=0.995 $X2=0
+ $Y2=0
cc_376 N_A_27_297#_c_345_n N_VGND_c_1134_n 0.00481673f $X=5.33 $Y=0.995 $X2=0
+ $Y2=0
cc_377 N_A_27_297#_M1006_s N_VGND_c_1135_n 0.00271249f $X=0.14 $Y=0.235 $X2=0
+ $Y2=0
cc_378 N_A_27_297#_c_342_n N_VGND_c_1135_n 0.00587047f $X=3.87 $Y=0.995 $X2=0
+ $Y2=0
cc_379 N_A_27_297#_c_343_n N_VGND_c_1135_n 0.006093f $X=4.34 $Y=0.995 $X2=0
+ $Y2=0
cc_380 N_A_27_297#_c_344_n N_VGND_c_1135_n 0.00608558f $X=4.81 $Y=0.995 $X2=0
+ $Y2=0
cc_381 N_A_27_297#_c_345_n N_VGND_c_1135_n 0.00745263f $X=5.33 $Y=0.995 $X2=0
+ $Y2=0
cc_382 N_A_27_297#_c_346_n N_VGND_c_1135_n 0.0137653f $X=0.28 $Y=0.39 $X2=0
+ $Y2=0
cc_383 N_A_27_297#_c_347_n N_VGND_c_1135_n 0.00567428f $X=0.665 $Y=0.81 $X2=0
+ $Y2=0
cc_384 N_B_c_494_n N_A_c_568_n 0.0243397f $X=7.73 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_385 N_B_c_500_n N_A_c_574_n 0.00971598f $X=7.705 $Y=1.41 $X2=0 $Y2=0
cc_386 N_B_c_495_n N_A_c_572_n 0.0121231f $X=7.59 $Y=1.16 $X2=0 $Y2=0
cc_387 N_B_c_496_n N_A_c_572_n 2.62535e-19 $X=7.705 $Y=1.202 $X2=0 $Y2=0
cc_388 N_B_c_495_n N_A_c_573_n 2.62535e-19 $X=7.59 $Y=1.16 $X2=0 $Y2=0
cc_389 N_B_c_496_n N_A_c_573_n 0.0243397f $X=7.705 $Y=1.202 $X2=0 $Y2=0
cc_390 N_B_c_497_n N_VPWR_c_641_n 0.00429453f $X=6.295 $Y=1.41 $X2=0 $Y2=0
cc_391 N_B_c_498_n N_VPWR_c_641_n 0.00429453f $X=6.765 $Y=1.41 $X2=0 $Y2=0
cc_392 N_B_c_499_n N_VPWR_c_641_n 0.00429453f $X=7.235 $Y=1.41 $X2=0 $Y2=0
cc_393 N_B_c_500_n N_VPWR_c_641_n 0.00429453f $X=7.705 $Y=1.41 $X2=0 $Y2=0
cc_394 N_B_c_497_n N_VPWR_c_637_n 0.00734734f $X=6.295 $Y=1.41 $X2=0 $Y2=0
cc_395 N_B_c_498_n N_VPWR_c_637_n 0.00606499f $X=6.765 $Y=1.41 $X2=0 $Y2=0
cc_396 N_B_c_499_n N_VPWR_c_637_n 0.00606499f $X=7.235 $Y=1.41 $X2=0 $Y2=0
cc_397 N_B_c_500_n N_VPWR_c_637_n 0.00609021f $X=7.705 $Y=1.41 $X2=0 $Y2=0
cc_398 N_B_c_491_n N_Y_c_796_n 0.0109318f $X=6.27 $Y=0.995 $X2=0 $Y2=0
cc_399 N_B_c_495_n N_Y_c_796_n 0.0501575f $X=7.59 $Y=1.16 $X2=0 $Y2=0
cc_400 N_B_c_491_n N_Y_c_874_n 0.0110728f $X=6.27 $Y=0.995 $X2=0 $Y2=0
cc_401 N_B_c_492_n N_Y_c_874_n 0.00686626f $X=6.74 $Y=0.995 $X2=0 $Y2=0
cc_402 N_B_c_493_n N_Y_c_874_n 5.45498e-19 $X=7.21 $Y=0.995 $X2=0 $Y2=0
cc_403 N_B_c_492_n N_Y_c_797_n 0.00901745f $X=6.74 $Y=0.995 $X2=0 $Y2=0
cc_404 N_B_c_493_n N_Y_c_797_n 0.00901745f $X=7.21 $Y=0.995 $X2=0 $Y2=0
cc_405 N_B_c_495_n N_Y_c_797_n 0.0398926f $X=7.59 $Y=1.16 $X2=0 $Y2=0
cc_406 N_B_c_496_n N_Y_c_797_n 0.00345541f $X=7.705 $Y=1.202 $X2=0 $Y2=0
cc_407 N_B_c_492_n N_Y_c_881_n 5.24597e-19 $X=6.74 $Y=0.995 $X2=0 $Y2=0
cc_408 N_B_c_493_n N_Y_c_881_n 0.00651696f $X=7.21 $Y=0.995 $X2=0 $Y2=0
cc_409 N_B_c_494_n N_Y_c_798_n 0.0106151f $X=7.73 $Y=0.995 $X2=0 $Y2=0
cc_410 N_B_c_495_n N_Y_c_798_n 0.0118017f $X=7.59 $Y=1.16 $X2=0 $Y2=0
cc_411 N_B_c_494_n N_Y_c_885_n 5.32212e-19 $X=7.73 $Y=0.995 $X2=0 $Y2=0
cc_412 N_B_c_491_n N_Y_c_803_n 0.00116636f $X=6.27 $Y=0.995 $X2=0 $Y2=0
cc_413 N_B_c_492_n N_Y_c_803_n 0.00116636f $X=6.74 $Y=0.995 $X2=0 $Y2=0
cc_414 N_B_c_495_n N_Y_c_803_n 0.0307014f $X=7.59 $Y=1.16 $X2=0 $Y2=0
cc_415 N_B_c_496_n N_Y_c_803_n 0.00358305f $X=7.705 $Y=1.202 $X2=0 $Y2=0
cc_416 N_B_c_493_n N_Y_c_804_n 0.00119564f $X=7.21 $Y=0.995 $X2=0 $Y2=0
cc_417 N_B_c_495_n N_Y_c_804_n 0.030835f $X=7.59 $Y=1.16 $X2=0 $Y2=0
cc_418 N_B_c_496_n N_Y_c_804_n 0.00486271f $X=7.705 $Y=1.202 $X2=0 $Y2=0
cc_419 N_B_c_497_n N_A_797_297#_c_984_n 0.0148794f $X=6.295 $Y=1.41 $X2=0 $Y2=0
cc_420 N_B_c_495_n N_A_797_297#_c_984_n 0.0562521f $X=7.59 $Y=1.16 $X2=0 $Y2=0
cc_421 N_B_c_496_n N_A_797_297#_c_984_n 8.84531e-19 $X=7.705 $Y=1.202 $X2=0
+ $Y2=0
cc_422 N_B_c_498_n N_A_797_297#_c_985_n 0.0128795f $X=6.765 $Y=1.41 $X2=0 $Y2=0
cc_423 N_B_c_499_n N_A_797_297#_c_985_n 0.0128188f $X=7.235 $Y=1.41 $X2=0 $Y2=0
cc_424 N_B_c_495_n N_A_797_297#_c_985_n 0.0486996f $X=7.59 $Y=1.16 $X2=0 $Y2=0
cc_425 N_B_c_496_n N_A_797_297#_c_985_n 0.00864922f $X=7.705 $Y=1.202 $X2=0
+ $Y2=0
cc_426 N_B_c_495_n N_A_797_297#_c_988_n 0.0204252f $X=7.59 $Y=1.16 $X2=0 $Y2=0
cc_427 N_B_c_496_n N_A_797_297#_c_988_n 0.00655199f $X=7.705 $Y=1.202 $X2=0
+ $Y2=0
cc_428 N_B_c_500_n N_A_797_297#_c_989_n 2.98195e-19 $X=7.705 $Y=1.41 $X2=0 $Y2=0
cc_429 N_B_c_495_n N_A_797_297#_c_989_n 0.0204252f $X=7.59 $Y=1.16 $X2=0 $Y2=0
cc_430 N_B_c_496_n N_A_797_297#_c_989_n 0.00634604f $X=7.705 $Y=1.202 $X2=0
+ $Y2=0
cc_431 N_B_c_497_n N_A_1187_297#_c_1052_n 0.01161f $X=6.295 $Y=1.41 $X2=0 $Y2=0
cc_432 N_B_c_498_n N_A_1187_297#_c_1052_n 0.01161f $X=6.765 $Y=1.41 $X2=0 $Y2=0
cc_433 N_B_c_499_n N_A_1187_297#_c_1054_n 0.01161f $X=7.235 $Y=1.41 $X2=0 $Y2=0
cc_434 N_B_c_500_n N_A_1187_297#_c_1054_n 0.0143578f $X=7.705 $Y=1.41 $X2=0
+ $Y2=0
cc_435 N_B_c_500_n N_A_1187_297#_c_1046_n 2.98195e-19 $X=7.705 $Y=1.41 $X2=0
+ $Y2=0
cc_436 N_B_c_492_n N_VGND_c_1112_n 0.00379224f $X=6.74 $Y=0.995 $X2=0 $Y2=0
cc_437 N_B_c_493_n N_VGND_c_1112_n 0.00276126f $X=7.21 $Y=0.995 $X2=0 $Y2=0
cc_438 N_B_c_494_n N_VGND_c_1113_n 0.00268723f $X=7.73 $Y=0.995 $X2=0 $Y2=0
cc_439 N_B_c_491_n N_VGND_c_1125_n 0.00423334f $X=6.27 $Y=0.995 $X2=0 $Y2=0
cc_440 N_B_c_492_n N_VGND_c_1125_n 0.00423334f $X=6.74 $Y=0.995 $X2=0 $Y2=0
cc_441 N_B_c_493_n N_VGND_c_1127_n 0.00423334f $X=7.21 $Y=0.995 $X2=0 $Y2=0
cc_442 N_B_c_494_n N_VGND_c_1127_n 0.00437852f $X=7.73 $Y=0.995 $X2=0 $Y2=0
cc_443 N_B_c_491_n N_VGND_c_1134_n 0.00481673f $X=6.27 $Y=0.995 $X2=0 $Y2=0
cc_444 N_B_c_491_n N_VGND_c_1135_n 0.00716687f $X=6.27 $Y=0.995 $X2=0 $Y2=0
cc_445 N_B_c_492_n N_VGND_c_1135_n 0.006093f $X=6.74 $Y=0.995 $X2=0 $Y2=0
cc_446 N_B_c_493_n N_VGND_c_1135_n 0.00608558f $X=7.21 $Y=0.995 $X2=0 $Y2=0
cc_447 N_B_c_494_n N_VGND_c_1135_n 0.00615622f $X=7.73 $Y=0.995 $X2=0 $Y2=0
cc_448 N_A_c_574_n N_VPWR_c_639_n 0.00300743f $X=8.175 $Y=1.41 $X2=0 $Y2=0
cc_449 N_A_c_575_n N_VPWR_c_639_n 0.00300743f $X=8.645 $Y=1.41 $X2=0 $Y2=0
cc_450 N_A_c_576_n N_VPWR_c_640_n 0.00300743f $X=9.115 $Y=1.41 $X2=0 $Y2=0
cc_451 N_A_c_577_n N_VPWR_c_640_n 0.00300743f $X=9.585 $Y=1.41 $X2=0 $Y2=0
cc_452 N_A_c_574_n N_VPWR_c_641_n 0.00702461f $X=8.175 $Y=1.41 $X2=0 $Y2=0
cc_453 N_A_c_575_n N_VPWR_c_643_n 0.00702461f $X=8.645 $Y=1.41 $X2=0 $Y2=0
cc_454 N_A_c_576_n N_VPWR_c_643_n 0.00702461f $X=9.115 $Y=1.41 $X2=0 $Y2=0
cc_455 N_A_c_577_n N_VPWR_c_646_n 0.00702461f $X=9.585 $Y=1.41 $X2=0 $Y2=0
cc_456 N_A_c_574_n N_VPWR_c_637_n 0.0124344f $X=8.175 $Y=1.41 $X2=0 $Y2=0
cc_457 N_A_c_575_n N_VPWR_c_637_n 0.0124092f $X=8.645 $Y=1.41 $X2=0 $Y2=0
cc_458 N_A_c_576_n N_VPWR_c_637_n 0.0124092f $X=9.115 $Y=1.41 $X2=0 $Y2=0
cc_459 N_A_c_577_n N_VPWR_c_637_n 0.0133558f $X=9.585 $Y=1.41 $X2=0 $Y2=0
cc_460 N_A_c_568_n N_Y_c_798_n 0.00865686f $X=8.15 $Y=0.995 $X2=0 $Y2=0
cc_461 N_A_c_572_n N_Y_c_798_n 0.00826974f $X=9.47 $Y=1.16 $X2=0 $Y2=0
cc_462 N_A_c_568_n N_Y_c_885_n 0.00644736f $X=8.15 $Y=0.995 $X2=0 $Y2=0
cc_463 N_A_c_569_n N_Y_c_885_n 0.00686626f $X=8.62 $Y=0.995 $X2=0 $Y2=0
cc_464 N_A_c_570_n N_Y_c_885_n 5.45498e-19 $X=9.09 $Y=0.995 $X2=0 $Y2=0
cc_465 N_A_c_569_n N_Y_c_799_n 0.00901745f $X=8.62 $Y=0.995 $X2=0 $Y2=0
cc_466 N_A_c_570_n N_Y_c_799_n 0.010179f $X=9.09 $Y=0.995 $X2=0 $Y2=0
cc_467 N_A_c_571_n N_Y_c_799_n 2.15189e-19 $X=9.61 $Y=0.995 $X2=0 $Y2=0
cc_468 N_A_c_572_n N_Y_c_799_n 0.0707276f $X=9.47 $Y=1.16 $X2=0 $Y2=0
cc_469 N_A_c_573_n N_Y_c_799_n 0.00831812f $X=9.585 $Y=1.202 $X2=0 $Y2=0
cc_470 N_A_c_569_n N_Y_c_903_n 5.24597e-19 $X=8.62 $Y=0.995 $X2=0 $Y2=0
cc_471 N_A_c_570_n N_Y_c_903_n 0.00651696f $X=9.09 $Y=0.995 $X2=0 $Y2=0
cc_472 N_A_c_568_n N_Y_c_805_n 0.00116636f $X=8.15 $Y=0.995 $X2=0 $Y2=0
cc_473 N_A_c_569_n N_Y_c_805_n 0.00116636f $X=8.62 $Y=0.995 $X2=0 $Y2=0
cc_474 N_A_c_572_n N_Y_c_805_n 0.0307014f $X=9.47 $Y=1.16 $X2=0 $Y2=0
cc_475 N_A_c_573_n N_Y_c_805_n 0.00358305f $X=9.585 $Y=1.202 $X2=0 $Y2=0
cc_476 N_A_c_574_n N_A_1187_297#_c_1047_n 0.0155666f $X=8.175 $Y=1.41 $X2=0
+ $Y2=0
cc_477 N_A_c_575_n N_A_1187_297#_c_1047_n 0.0156273f $X=8.645 $Y=1.41 $X2=0
+ $Y2=0
cc_478 N_A_c_572_n N_A_1187_297#_c_1047_n 0.0480109f $X=9.47 $Y=1.16 $X2=0 $Y2=0
cc_479 N_A_c_573_n N_A_1187_297#_c_1047_n 0.00837544f $X=9.585 $Y=1.202 $X2=0
+ $Y2=0
cc_480 N_A_c_576_n N_A_1187_297#_c_1048_n 0.0156273f $X=9.115 $Y=1.41 $X2=0
+ $Y2=0
cc_481 N_A_c_577_n N_A_1187_297#_c_1048_n 0.0158609f $X=9.585 $Y=1.41 $X2=0
+ $Y2=0
cc_482 N_A_c_572_n N_A_1187_297#_c_1048_n 0.0487385f $X=9.47 $Y=1.16 $X2=0 $Y2=0
cc_483 N_A_c_573_n N_A_1187_297#_c_1048_n 0.00816971f $X=9.585 $Y=1.202 $X2=0
+ $Y2=0
cc_484 N_A_c_572_n N_A_1187_297#_c_1049_n 0.0269937f $X=9.47 $Y=1.16 $X2=0 $Y2=0
cc_485 N_A_c_572_n N_A_1187_297#_c_1051_n 0.0204509f $X=9.47 $Y=1.16 $X2=0 $Y2=0
cc_486 N_A_c_573_n N_A_1187_297#_c_1051_n 0.00656533f $X=9.585 $Y=1.202 $X2=0
+ $Y2=0
cc_487 N_A_c_568_n N_VGND_c_1113_n 0.00268723f $X=8.15 $Y=0.995 $X2=0 $Y2=0
cc_488 N_A_c_569_n N_VGND_c_1114_n 0.00379224f $X=8.62 $Y=0.995 $X2=0 $Y2=0
cc_489 N_A_c_570_n N_VGND_c_1114_n 0.00276126f $X=9.09 $Y=0.995 $X2=0 $Y2=0
cc_490 N_A_c_571_n N_VGND_c_1116_n 0.00498331f $X=9.61 $Y=0.995 $X2=0 $Y2=0
cc_491 N_A_c_572_n N_VGND_c_1116_n 0.0233945f $X=9.47 $Y=1.16 $X2=0 $Y2=0
cc_492 N_A_c_568_n N_VGND_c_1129_n 0.00423334f $X=8.15 $Y=0.995 $X2=0 $Y2=0
cc_493 N_A_c_569_n N_VGND_c_1129_n 0.00423334f $X=8.62 $Y=0.995 $X2=0 $Y2=0
cc_494 N_A_c_570_n N_VGND_c_1131_n 0.00423334f $X=9.09 $Y=0.995 $X2=0 $Y2=0
cc_495 N_A_c_571_n N_VGND_c_1131_n 0.00585385f $X=9.61 $Y=0.995 $X2=0 $Y2=0
cc_496 N_A_c_568_n N_VGND_c_1135_n 0.00587047f $X=8.15 $Y=0.995 $X2=0 $Y2=0
cc_497 N_A_c_569_n N_VGND_c_1135_n 0.006093f $X=8.62 $Y=0.995 $X2=0 $Y2=0
cc_498 N_A_c_570_n N_VGND_c_1135_n 0.00608558f $X=9.09 $Y=0.995 $X2=0 $Y2=0
cc_499 N_A_c_571_n N_VGND_c_1135_n 0.0117699f $X=9.61 $Y=0.995 $X2=0 $Y2=0
cc_500 N_VPWR_c_637_n N_A_331_297#_M1000_s 0.00217543f $X=9.89 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_501 N_VPWR_c_637_n N_A_331_297#_M1010_s 0.00231289f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_502 N_VPWR_c_637_n N_A_331_297#_M1029_s 0.00231289f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_637_n N_A_331_297#_M1018_s 0.00231264f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_637_n N_A_331_297#_M1035_s 0.00217519f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_505 N_VPWR_c_641_n N_A_331_297#_c_743_n 0.163661f $X=8.285 $Y=2.72 $X2=0
+ $Y2=0
cc_506 N_VPWR_c_637_n N_A_331_297#_c_743_n 0.101859f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_507 N_VPWR_c_641_n N_A_331_297#_c_744_n 0.0571048f $X=8.285 $Y=2.72 $X2=0
+ $Y2=0
cc_508 N_VPWR_c_637_n N_A_331_297#_c_744_n 0.0346935f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_509 N_VPWR_c_641_n N_A_331_297#_c_773_n 0.0149886f $X=8.285 $Y=2.72 $X2=0
+ $Y2=0
cc_510 N_VPWR_c_637_n N_A_331_297#_c_773_n 0.00962421f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_511 N_VPWR_c_637_n N_Y_M1000_d 0.00232895f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_512 N_VPWR_c_637_n N_Y_M1016_d 0.00232895f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_513 N_VPWR_c_637_n N_A_797_297#_M1013_d 0.00232895f $X=9.89 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_514 N_VPWR_c_637_n N_A_797_297#_M1024_d 0.00232895f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_515 N_VPWR_c_637_n N_A_797_297#_M1001_s 0.00232895f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_516 N_VPWR_c_637_n N_A_797_297#_M1017_s 0.00232895f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_517 N_VPWR_c_637_n N_A_1187_297#_M1001_d 0.00217519f $X=9.89 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_518 N_VPWR_c_637_n N_A_1187_297#_M1011_d 0.00231264f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_519 N_VPWR_c_637_n N_A_1187_297#_M1022_d 0.00297222f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_520 N_VPWR_c_637_n N_A_1187_297#_M1025_s 0.00370124f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_521 N_VPWR_c_637_n N_A_1187_297#_M1032_s 0.00303344f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_522 N_VPWR_c_641_n N_A_1187_297#_c_1052_n 0.0386815f $X=8.285 $Y=2.72 $X2=0
+ $Y2=0
cc_523 N_VPWR_c_637_n N_A_1187_297#_c_1052_n 0.0239144f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_524 N_VPWR_c_641_n N_A_1187_297#_c_1045_n 0.0202137f $X=8.285 $Y=2.72 $X2=0
+ $Y2=0
cc_525 N_VPWR_c_637_n N_A_1187_297#_c_1045_n 0.0117415f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_526 N_VPWR_c_641_n N_A_1187_297#_c_1054_n 0.0386815f $X=8.285 $Y=2.72 $X2=0
+ $Y2=0
cc_527 N_VPWR_c_637_n N_A_1187_297#_c_1054_n 0.0239144f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_528 N_VPWR_c_641_n N_A_1187_297#_c_1079_n 0.015002f $X=8.285 $Y=2.72 $X2=0
+ $Y2=0
cc_529 N_VPWR_c_637_n N_A_1187_297#_c_1079_n 0.00962794f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_530 N_VPWR_M1020_d N_A_1187_297#_c_1047_n 0.00187091f $X=8.265 $Y=1.485 $X2=0
+ $Y2=0
cc_531 N_VPWR_c_639_n N_A_1187_297#_c_1047_n 0.0143191f $X=8.41 $Y=1.96 $X2=0
+ $Y2=0
cc_532 N_VPWR_c_643_n N_A_1187_297#_c_1083_n 0.0149311f $X=9.225 $Y=2.72 $X2=0
+ $Y2=0
cc_533 N_VPWR_c_637_n N_A_1187_297#_c_1083_n 0.00955092f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_534 N_VPWR_M1030_d N_A_1187_297#_c_1048_n 0.00187091f $X=9.205 $Y=1.485 $X2=0
+ $Y2=0
cc_535 N_VPWR_c_640_n N_A_1187_297#_c_1048_n 0.0143191f $X=9.35 $Y=1.96 $X2=0
+ $Y2=0
cc_536 N_VPWR_c_646_n N_A_1187_297#_c_1050_n 0.0208166f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_537 N_VPWR_c_637_n N_A_1187_297#_c_1050_n 0.0120542f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_641_n N_A_1187_297#_c_1089_n 0.0149886f $X=8.285 $Y=2.72 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_637_n N_A_1187_297#_c_1089_n 0.00962421f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_540 N_A_331_297#_c_743_n N_Y_M1000_d 0.00357068f $X=3.7 $Y=2.34 $X2=0 $Y2=0
cc_541 N_A_331_297#_c_743_n N_Y_M1016_d 0.00357068f $X=3.7 $Y=2.34 $X2=0 $Y2=0
cc_542 N_A_331_297#_M1010_s N_Y_c_807_n 0.00190658f $X=2.575 $Y=1.485 $X2=0
+ $Y2=0
cc_543 N_A_331_297#_c_758_n N_A_797_297#_M1013_d 0.00345323f $X=4.475 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_544 N_A_331_297#_c_744_n N_A_797_297#_M1024_d 0.00352392f $X=5.415 $Y=2.38
+ $X2=0 $Y2=0
cc_545 N_A_331_297#_M1018_s N_A_797_297#_c_983_n 0.00187091f $X=4.455 $Y=1.485
+ $X2=0 $Y2=0
cc_546 N_A_331_297#_c_758_n N_A_797_297#_c_983_n 0.00385532f $X=4.475 $Y=2.38
+ $X2=0 $Y2=0
cc_547 N_A_331_297#_c_782_p N_A_797_297#_c_983_n 0.0143018f $X=4.6 $Y=1.96 $X2=0
+ $Y2=0
cc_548 N_A_331_297#_c_744_n N_A_797_297#_c_983_n 0.00385532f $X=5.415 $Y=2.38
+ $X2=0 $Y2=0
cc_549 N_A_331_297#_M1035_s N_A_797_297#_c_984_n 0.00295666f $X=5.395 $Y=1.485
+ $X2=0 $Y2=0
cc_550 N_A_331_297#_c_744_n N_A_797_297#_c_984_n 0.00385532f $X=5.415 $Y=2.38
+ $X2=0 $Y2=0
cc_551 N_A_331_297#_c_745_n N_A_797_297#_c_984_n 0.0197547f $X=5.54 $Y=1.96
+ $X2=0 $Y2=0
cc_552 N_A_331_297#_c_758_n N_A_797_297#_c_986_n 0.0130906f $X=4.475 $Y=2.38
+ $X2=0 $Y2=0
cc_553 N_A_331_297#_c_744_n N_A_797_297#_c_987_n 0.013395f $X=5.415 $Y=2.38
+ $X2=0 $Y2=0
cc_554 N_A_331_297#_c_745_n N_A_1187_297#_c_1044_n 0.0384367f $X=5.54 $Y=1.96
+ $X2=0 $Y2=0
cc_555 N_A_331_297#_c_744_n N_A_1187_297#_c_1045_n 0.0149967f $X=5.415 $Y=2.38
+ $X2=0 $Y2=0
cc_556 N_Y_c_796_n N_A_797_297#_c_984_n 0.00820983f $X=6.315 $Y=0.815 $X2=0
+ $Y2=0
cc_557 N_Y_c_798_n N_A_1187_297#_c_1046_n 0.00936521f $X=8.195 $Y=0.815 $X2=0
+ $Y2=0
cc_558 N_Y_c_798_n N_A_1187_297#_c_1047_n 3.18413e-19 $X=8.195 $Y=0.815 $X2=0
+ $Y2=0
cc_559 N_Y_c_791_n N_VGND_M1019_d 0.00251047f $X=2.975 $Y=0.815 $X2=0 $Y2=0
cc_560 N_Y_c_794_n N_VGND_M1028_d 0.00162089f $X=3.915 $Y=0.815 $X2=0 $Y2=0
cc_561 N_Y_c_795_n N_VGND_M1005_s 0.00251047f $X=4.855 $Y=0.815 $X2=0 $Y2=0
cc_562 N_Y_c_796_n N_VGND_M1015_s 0.0108248f $X=6.315 $Y=0.815 $X2=0 $Y2=0
cc_563 N_Y_c_797_n N_VGND_M1014_s 0.00251047f $X=7.255 $Y=0.815 $X2=0 $Y2=0
cc_564 N_Y_c_798_n N_VGND_M1033_s 0.00162089f $X=8.195 $Y=0.815 $X2=0 $Y2=0
cc_565 N_Y_c_799_n N_VGND_M1021_s 0.00251047f $X=9.135 $Y=0.815 $X2=0 $Y2=0
cc_566 N_Y_c_808_n N_VGND_c_1109_n 0.0183628f $X=2.25 $Y=0.39 $X2=0 $Y2=0
cc_567 N_Y_c_791_n N_VGND_c_1109_n 0.0127273f $X=2.975 $Y=0.815 $X2=0 $Y2=0
cc_568 N_Y_c_794_n N_VGND_c_1110_n 0.0122559f $X=3.915 $Y=0.815 $X2=0 $Y2=0
cc_569 N_Y_c_829_n N_VGND_c_1111_n 0.0183628f $X=4.13 $Y=0.39 $X2=0 $Y2=0
cc_570 N_Y_c_795_n N_VGND_c_1111_n 0.0127273f $X=4.855 $Y=0.815 $X2=0 $Y2=0
cc_571 N_Y_c_874_n N_VGND_c_1112_n 0.0183628f $X=6.53 $Y=0.39 $X2=0 $Y2=0
cc_572 N_Y_c_797_n N_VGND_c_1112_n 0.0127273f $X=7.255 $Y=0.815 $X2=0 $Y2=0
cc_573 N_Y_c_798_n N_VGND_c_1113_n 0.0122559f $X=8.195 $Y=0.815 $X2=0 $Y2=0
cc_574 N_Y_c_885_n N_VGND_c_1114_n 0.0183628f $X=8.41 $Y=0.39 $X2=0 $Y2=0
cc_575 N_Y_c_799_n N_VGND_c_1114_n 0.0127273f $X=9.135 $Y=0.815 $X2=0 $Y2=0
cc_576 N_Y_c_799_n N_VGND_c_1116_n 0.00138214f $X=9.135 $Y=0.815 $X2=0 $Y2=0
cc_577 N_Y_c_808_n N_VGND_c_1119_n 0.0223596f $X=2.25 $Y=0.39 $X2=0 $Y2=0
cc_578 N_Y_c_791_n N_VGND_c_1119_n 0.00266636f $X=2.975 $Y=0.815 $X2=0 $Y2=0
cc_579 N_Y_c_791_n N_VGND_c_1121_n 0.00198695f $X=2.975 $Y=0.815 $X2=0 $Y2=0
cc_580 N_Y_c_822_n N_VGND_c_1121_n 0.0231929f $X=3.19 $Y=0.39 $X2=0 $Y2=0
cc_581 N_Y_c_794_n N_VGND_c_1121_n 0.00158379f $X=3.915 $Y=0.815 $X2=0 $Y2=0
cc_582 N_Y_c_800_n N_VGND_c_1121_n 0.00103384f $X=3.205 $Y=0.815 $X2=0 $Y2=0
cc_583 N_Y_c_794_n N_VGND_c_1123_n 0.00198695f $X=3.915 $Y=0.815 $X2=0 $Y2=0
cc_584 N_Y_c_829_n N_VGND_c_1123_n 0.0223596f $X=4.13 $Y=0.39 $X2=0 $Y2=0
cc_585 N_Y_c_795_n N_VGND_c_1123_n 0.00266636f $X=4.855 $Y=0.815 $X2=0 $Y2=0
cc_586 N_Y_c_796_n N_VGND_c_1125_n 0.00198695f $X=6.315 $Y=0.815 $X2=0 $Y2=0
cc_587 N_Y_c_874_n N_VGND_c_1125_n 0.0223596f $X=6.53 $Y=0.39 $X2=0 $Y2=0
cc_588 N_Y_c_797_n N_VGND_c_1125_n 0.00266636f $X=7.255 $Y=0.815 $X2=0 $Y2=0
cc_589 N_Y_c_797_n N_VGND_c_1127_n 0.00198695f $X=7.255 $Y=0.815 $X2=0 $Y2=0
cc_590 N_Y_c_881_n N_VGND_c_1127_n 0.0231806f $X=7.47 $Y=0.39 $X2=0 $Y2=0
cc_591 N_Y_c_798_n N_VGND_c_1127_n 0.00254521f $X=8.195 $Y=0.815 $X2=0 $Y2=0
cc_592 N_Y_c_798_n N_VGND_c_1129_n 0.00198695f $X=8.195 $Y=0.815 $X2=0 $Y2=0
cc_593 N_Y_c_885_n N_VGND_c_1129_n 0.0223596f $X=8.41 $Y=0.39 $X2=0 $Y2=0
cc_594 N_Y_c_799_n N_VGND_c_1129_n 0.00266636f $X=9.135 $Y=0.815 $X2=0 $Y2=0
cc_595 N_Y_c_799_n N_VGND_c_1131_n 0.00198695f $X=9.135 $Y=0.815 $X2=0 $Y2=0
cc_596 N_Y_c_903_n N_VGND_c_1131_n 0.0231806f $X=9.35 $Y=0.39 $X2=0 $Y2=0
cc_597 N_Y_c_795_n N_VGND_c_1133_n 0.00198695f $X=4.855 $Y=0.815 $X2=0 $Y2=0
cc_598 N_Y_c_858_n N_VGND_c_1133_n 0.0231806f $X=5.07 $Y=0.39 $X2=0 $Y2=0
cc_599 N_Y_c_796_n N_VGND_c_1133_n 0.00254521f $X=6.315 $Y=0.815 $X2=0 $Y2=0
cc_600 N_Y_c_796_n N_VGND_c_1134_n 0.0528344f $X=6.315 $Y=0.815 $X2=0 $Y2=0
cc_601 N_Y_M1007_s N_VGND_c_1135_n 0.0025535f $X=2.065 $Y=0.235 $X2=0 $Y2=0
cc_602 N_Y_M1027_s N_VGND_c_1135_n 0.00304114f $X=3.005 $Y=0.235 $X2=0 $Y2=0
cc_603 N_Y_M1004_d N_VGND_c_1135_n 0.0025535f $X=3.945 $Y=0.235 $X2=0 $Y2=0
cc_604 N_Y_M1012_d N_VGND_c_1135_n 0.00304143f $X=4.885 $Y=0.235 $X2=0 $Y2=0
cc_605 N_Y_M1009_d N_VGND_c_1135_n 0.0025535f $X=6.345 $Y=0.235 $X2=0 $Y2=0
cc_606 N_Y_M1031_d N_VGND_c_1135_n 0.00304143f $X=7.285 $Y=0.235 $X2=0 $Y2=0
cc_607 N_Y_M1008_d N_VGND_c_1135_n 0.0025535f $X=8.225 $Y=0.235 $X2=0 $Y2=0
cc_608 N_Y_M1023_d N_VGND_c_1135_n 0.00364931f $X=9.165 $Y=0.235 $X2=0 $Y2=0
cc_609 N_Y_c_808_n N_VGND_c_1135_n 0.0141302f $X=2.25 $Y=0.39 $X2=0 $Y2=0
cc_610 N_Y_c_791_n N_VGND_c_1135_n 0.00972452f $X=2.975 $Y=0.815 $X2=0 $Y2=0
cc_611 N_Y_c_822_n N_VGND_c_1135_n 0.0143393f $X=3.19 $Y=0.39 $X2=0 $Y2=0
cc_612 N_Y_c_794_n N_VGND_c_1135_n 0.00771335f $X=3.915 $Y=0.815 $X2=0 $Y2=0
cc_613 N_Y_c_829_n N_VGND_c_1135_n 0.0141302f $X=4.13 $Y=0.39 $X2=0 $Y2=0
cc_614 N_Y_c_795_n N_VGND_c_1135_n 0.00972452f $X=4.855 $Y=0.815 $X2=0 $Y2=0
cc_615 N_Y_c_858_n N_VGND_c_1135_n 0.0143352f $X=5.07 $Y=0.39 $X2=0 $Y2=0
cc_616 N_Y_c_796_n N_VGND_c_1135_n 0.0114512f $X=6.315 $Y=0.815 $X2=0 $Y2=0
cc_617 N_Y_c_874_n N_VGND_c_1135_n 0.0141302f $X=6.53 $Y=0.39 $X2=0 $Y2=0
cc_618 N_Y_c_797_n N_VGND_c_1135_n 0.00972452f $X=7.255 $Y=0.815 $X2=0 $Y2=0
cc_619 N_Y_c_881_n N_VGND_c_1135_n 0.0143352f $X=7.47 $Y=0.39 $X2=0 $Y2=0
cc_620 N_Y_c_798_n N_VGND_c_1135_n 0.0094839f $X=8.195 $Y=0.815 $X2=0 $Y2=0
cc_621 N_Y_c_885_n N_VGND_c_1135_n 0.0141302f $X=8.41 $Y=0.39 $X2=0 $Y2=0
cc_622 N_Y_c_799_n N_VGND_c_1135_n 0.00972452f $X=9.135 $Y=0.815 $X2=0 $Y2=0
cc_623 N_Y_c_903_n N_VGND_c_1135_n 0.0143352f $X=9.35 $Y=0.39 $X2=0 $Y2=0
cc_624 N_Y_c_800_n N_VGND_c_1135_n 0.00189268f $X=3.205 $Y=0.815 $X2=0 $Y2=0
cc_625 N_A_797_297#_c_984_n N_A_1187_297#_M1001_d 0.00295666f $X=6.405 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_626 N_A_797_297#_c_985_n N_A_1187_297#_M1011_d 0.00187091f $X=7.345 $Y=1.54
+ $X2=0 $Y2=0
cc_627 N_A_797_297#_c_984_n N_A_1187_297#_c_1044_n 0.0218636f $X=6.405 $Y=1.54
+ $X2=0 $Y2=0
cc_628 N_A_797_297#_M1001_s N_A_1187_297#_c_1052_n 0.00352392f $X=6.385 $Y=1.485
+ $X2=0 $Y2=0
cc_629 N_A_797_297#_c_984_n N_A_1187_297#_c_1052_n 0.00385532f $X=6.405 $Y=1.54
+ $X2=0 $Y2=0
cc_630 N_A_797_297#_c_985_n N_A_1187_297#_c_1052_n 0.00385532f $X=7.345 $Y=1.54
+ $X2=0 $Y2=0
cc_631 N_A_797_297#_c_988_n N_A_1187_297#_c_1052_n 0.013395f $X=6.53 $Y=1.62
+ $X2=0 $Y2=0
cc_632 N_A_797_297#_c_985_n N_A_1187_297#_c_1102_n 0.0143018f $X=7.345 $Y=1.54
+ $X2=0 $Y2=0
cc_633 N_A_797_297#_M1017_s N_A_1187_297#_c_1054_n 0.00352392f $X=7.325 $Y=1.485
+ $X2=0 $Y2=0
cc_634 N_A_797_297#_c_985_n N_A_1187_297#_c_1054_n 0.00385532f $X=7.345 $Y=1.54
+ $X2=0 $Y2=0
cc_635 N_A_797_297#_c_989_n N_A_1187_297#_c_1054_n 0.013395f $X=7.47 $Y=1.62
+ $X2=0 $Y2=0
cc_636 N_A_797_297#_c_989_n N_A_1187_297#_c_1046_n 0.00226124f $X=7.47 $Y=1.62
+ $X2=0 $Y2=0
