* File: sky130_fd_sc_hdll__nand4bb_2.pex.spice
* Created: Thu Aug 27 19:15:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_2%B_N 4 5 7 8 10 13 15 17 18 22 24
c43 17 0 1.71118e-19 $X=0.235 $Y=1.19
c44 15 0 1.28647e-19 $X=0.305 $Y=1.887
c45 5 0 7.16994e-20 $X=0.495 $Y=1.99
r46 22 25 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r47 22 24 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r48 17 18 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r49 17 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r50 15 16 50.8778 $w=1.8e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.887
+ $X2=0.495 $Y2=1.887
r51 11 13 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.52 $Y2=0.805
r52 8 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.805
r53 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.445
r54 5 16 2.83073 $w=1.8e-07 $l=1.03e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=1.887
r55 5 7 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r56 4 15 7.1379 $w=1.5e-07 $l=1.02e-07 $layer=POLY_cond $X=0.305 $Y=1.785
+ $X2=0.305 $Y2=1.887
r57 4 25 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.305 $Y=1.785
+ $X2=0.305 $Y2=1.4
r58 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r59 1 24 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_N 2 3 5 8 10 11 19
c41 8 0 1.47484e-20 $X=0.99 $Y=0.445
c42 2 0 1.56369e-19 $X=0.965 $Y=1.89
r43 18 19 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.255
+ $X2=0.99 $Y2=1.255
r44 15 18 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.775 $Y=1.255
+ $X2=0.965 $Y2=1.255
r45 10 11 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=0.75 $Y=1.19
+ $X2=0.75 $Y2=1.53
r46 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.775
+ $Y=1.255 $X2=0.775 $Y2=1.255
r47 6 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=1.09
+ $X2=0.99 $Y2=1.255
r48 6 8 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=0.99 $Y=1.09 $X2=0.99
+ $Y2=0.445
r49 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.965 $Y=1.99
+ $X2=0.965 $Y2=2.275
r50 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.89 $X2=0.965
+ $Y2=1.99
r51 1 18 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.42
+ $X2=0.965 $Y2=1.255
r52 1 2 155.841 $w=2e-07 $l=4.7e-07 $layer=POLY_cond $X=0.965 $Y=1.42 $X2=0.965
+ $Y2=1.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_211_413# 1 2 7 9 10 12 13 15 18 20 23
+ 25 29 36
c77 29 0 7.16994e-20 $X=1.5 $Y=2.307
r78 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.585
+ $Y=1.16 $X2=1.585 $Y2=1.16
r79 34 36 62.7429 $w=1.73e-07 $l=9.9e-07 $layer=LI1_cond $X=1.587 $Y=2.15
+ $X2=1.587 $Y2=1.16
r80 33 36 38.026 $w=1.73e-07 $l=6e-07 $layer=LI1_cond $X=1.587 $Y=0.56 $X2=1.587
+ $Y2=1.16
r81 29 34 7.5664 $w=3.15e-07 $l=1.95724e-07 $layer=LI1_cond $X=1.5 $Y=2.307
+ $X2=1.587 $Y2=2.15
r82 29 31 10.9756 $w=3.13e-07 $l=3e-07 $layer=LI1_cond $X=1.5 $Y=2.307 $X2=1.2
+ $Y2=2.307
r83 25 33 7.48781 $w=3.05e-07 $l=1.91625e-07 $layer=LI1_cond $X=1.5 $Y=0.407
+ $X2=1.587 $Y2=0.56
r84 25 27 11.3355 $w=3.03e-07 $l=3e-07 $layer=LI1_cond $X=1.5 $Y=0.407 $X2=1.2
+ $Y2=0.407
r85 23 24 3.47262 $w=3.47e-07 $l=2.5e-08 $layer=POLY_cond $X=2.635 $Y=1.202
+ $X2=2.66 $Y2=1.202
r86 22 23 61.8127 $w=3.47e-07 $l=4.45e-07 $layer=POLY_cond $X=2.19 $Y=1.202
+ $X2=2.635 $Y2=1.202
r87 21 22 3.47262 $w=3.47e-07 $l=2.5e-08 $layer=POLY_cond $X=2.165 $Y=1.202
+ $X2=2.19 $Y2=1.202
r88 20 37 83.9334 $w=3.3e-07 $l=4.8e-07 $layer=POLY_cond $X=2.065 $Y=1.16
+ $X2=1.585 $Y2=1.16
r89 20 21 14.0525 $w=3.47e-07 $l=1.19164e-07 $layer=POLY_cond $X=2.065 $Y=1.16
+ $X2=2.165 $Y2=1.202
r90 16 24 22.4223 $w=1.5e-07 $l=1.77e-07 $layer=POLY_cond $X=2.66 $Y=1.025
+ $X2=2.66 $Y2=1.202
r91 16 18 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.66 $Y=1.025
+ $X2=2.66 $Y2=0.56
r92 13 23 18.1053 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.635 $Y=1.41
+ $X2=2.635 $Y2=1.202
r93 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.635 $Y=1.41
+ $X2=2.635 $Y2=1.985
r94 10 22 22.4223 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.19 $Y=0.995
+ $X2=2.19 $Y2=1.202
r95 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.19 $Y=0.995
+ $X2=2.19 $Y2=0.56
r96 7 21 18.1053 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.165 $Y=1.41
+ $X2=2.165 $Y2=1.202
r97 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.165 $Y=1.41
+ $X2=2.165 $Y2=1.985
r98 2 31 600 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=2.065 $X2=1.2 $Y2=2.33
r99 1 27 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_27_47# 1 2 7 9 12 14 16 19 23 27 29 30
+ 31 32 37 40 46 48
c109 7 0 1.7445e-19 $X=3.105 $Y=1.41
r110 48 49 3.61862 $w=3.33e-07 $l=2.5e-08 $layer=POLY_cond $X=3.575 $Y=1.217
+ $X2=3.6 $Y2=1.217
r111 47 48 64.4114 $w=3.33e-07 $l=4.45e-07 $layer=POLY_cond $X=3.13 $Y=1.217
+ $X2=3.575 $Y2=1.217
r112 45 47 2.89489 $w=3.33e-07 $l=2e-08 $layer=POLY_cond $X=3.11 $Y=1.217
+ $X2=3.13 $Y2=1.217
r113 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.11
+ $Y=1.16 $X2=3.11 $Y2=1.16
r114 43 45 0.723724 $w=3.33e-07 $l=5e-09 $layer=POLY_cond $X=3.105 $Y=1.217
+ $X2=3.11 $Y2=1.217
r115 40 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.24 $Y=1.19
+ $X2=3.24 $Y2=1.19
r116 36 40 1.28 $w=2.3e-07 $l=1.995e-06 $layer=MET1_cond $X=1.245 $Y=1.19
+ $X2=3.24 $Y2=1.19
r117 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.245 $Y=1.19
+ $X2=1.245 $Y2=1.19
r118 34 37 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=1.245 $Y=1.785
+ $X2=1.245 $Y2=1.19
r119 33 37 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.245 $Y=0.9
+ $X2=1.245 $Y2=1.19
r120 31 34 6.85817 $w=1.95e-07 $l=1.32868e-07 $layer=LI1_cond $X=1.16 $Y=1.882
+ $X2=1.245 $Y2=1.785
r121 31 32 44.9324 $w=1.93e-07 $l=7.9e-07 $layer=LI1_cond $X=1.16 $Y=1.882
+ $X2=0.37 $Y2=1.882
r122 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.16 $Y=0.815
+ $X2=1.245 $Y2=0.9
r123 29 30 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=1.16 $Y=0.815
+ $X2=0.345 $Y2=0.815
r124 25 32 7.13288 $w=1.95e-07 $l=1.85642e-07 $layer=LI1_cond $X=0.227 $Y=1.98
+ $X2=0.37 $Y2=1.882
r125 25 27 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=0.227 $Y=1.98
+ $X2=0.227 $Y2=2.275
r126 21 30 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.73
+ $X2=0.345 $Y2=0.815
r127 21 23 11.9677 $w=2.58e-07 $l=2.7e-07 $layer=LI1_cond $X=0.215 $Y=0.73
+ $X2=0.215 $Y2=0.46
r128 17 49 21.4384 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.6 $Y=1.025
+ $X2=3.6 $Y2=1.217
r129 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.6 $Y=1.025
+ $X2=3.6 $Y2=0.56
r130 14 48 17.1428 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.575 $Y=1.41
+ $X2=3.575 $Y2=1.217
r131 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.575 $Y=1.41
+ $X2=3.575 $Y2=1.985
r132 10 47 21.4384 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.13 $Y=1.025
+ $X2=3.13 $Y2=1.217
r133 10 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.13 $Y=1.025
+ $X2=3.13 $Y2=0.56
r134 7 43 17.1428 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.105 $Y=1.41
+ $X2=3.105 $Y2=1.217
r135 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.105 $Y=1.41
+ $X2=3.105 $Y2=1.985
r136 2 27 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.275
r137 1 23 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_2%C 1 3 6 8 10 13 15 16 24 29 31
c45 16 0 1.97021e-19 $X=4.74 $Y=1.105
c46 13 0 1.91072e-19 $X=5.03 $Y=0.56
r47 29 31 21.0727 $w=1.98e-07 $l=3.8e-07 $layer=LI1_cond $X=4.39 $Y=1.175
+ $X2=4.77 $Y2=1.175
r48 24 25 3.53372 $w=3.41e-07 $l=2.5e-08 $layer=POLY_cond $X=5.005 $Y=1.212
+ $X2=5.03 $Y2=1.212
r49 22 24 33.217 $w=3.41e-07 $l=2.35e-07 $layer=POLY_cond $X=4.77 $Y=1.212
+ $X2=5.005 $Y2=1.212
r50 22 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.77
+ $Y=1.16 $X2=4.77 $Y2=1.16
r51 20 22 29.6833 $w=3.41e-07 $l=2.1e-07 $layer=POLY_cond $X=4.56 $Y=1.212
+ $X2=4.77 $Y2=1.212
r52 19 20 3.53372 $w=3.41e-07 $l=2.5e-08 $layer=POLY_cond $X=4.535 $Y=1.212
+ $X2=4.56 $Y2=1.212
r53 16 31 3.05 $w=1.98e-07 $l=5.5e-08 $layer=LI1_cond $X=4.825 $Y=1.175 $X2=4.77
+ $Y2=1.175
r54 15 29 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=4.375 $Y=1.175
+ $X2=4.39 $Y2=1.175
r55 11 25 22.0049 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=5.03 $Y=1.025
+ $X2=5.03 $Y2=1.212
r56 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.03 $Y=1.025
+ $X2=5.03 $Y2=0.56
r57 8 24 17.6972 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=5.005 $Y=1.41
+ $X2=5.005 $Y2=1.212
r58 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.005 $Y=1.41
+ $X2=5.005 $Y2=1.985
r59 4 20 22.0049 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=4.56 $Y=1.015
+ $X2=4.56 $Y2=1.212
r60 4 6 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.56 $Y=1.015
+ $X2=4.56 $Y2=0.56
r61 1 19 17.6972 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=4.535 $Y=1.41
+ $X2=4.535 $Y2=1.212
r62 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.535 $Y=1.41
+ $X2=4.535 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_2%D 1 3 6 8 10 13 15 16 22 29 31
c44 22 0 1.97021e-19 $X=5.97 $Y=1.212
r45 29 31 18.5773 $w=1.98e-07 $l=3.35e-07 $layer=LI1_cond $X=5.74 $Y=1.175
+ $X2=6.075 $Y2=1.175
r46 24 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.075
+ $Y=1.16 $X2=6.075 $Y2=1.16
r47 22 24 15.5723 $w=3.25e-07 $l=1.05e-07 $layer=POLY_cond $X=5.97 $Y=1.212
+ $X2=6.075 $Y2=1.212
r48 21 22 3.70769 $w=3.25e-07 $l=2.5e-08 $layer=POLY_cond $X=5.945 $Y=1.212
+ $X2=5.97 $Y2=1.212
r49 20 21 65.9969 $w=3.25e-07 $l=4.45e-07 $layer=POLY_cond $X=5.5 $Y=1.212
+ $X2=5.945 $Y2=1.212
r50 19 20 3.70769 $w=3.25e-07 $l=2.5e-08 $layer=POLY_cond $X=5.475 $Y=1.212
+ $X2=5.5 $Y2=1.212
r51 16 31 3.32727 $w=1.98e-07 $l=6e-08 $layer=LI1_cond $X=6.135 $Y=1.175
+ $X2=6.075 $Y2=1.175
r52 15 29 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=5.73 $Y=1.175
+ $X2=5.74 $Y2=1.175
r53 11 22 20.86 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=5.97 $Y=1.015
+ $X2=5.97 $Y2=1.212
r54 11 13 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=5.97 $Y=1.015
+ $X2=5.97 $Y2=0.56
r55 8 21 16.5763 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=5.945 $Y=1.41
+ $X2=5.945 $Y2=1.212
r56 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.945 $Y=1.41
+ $X2=5.945 $Y2=1.985
r57 4 20 20.86 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=5.5 $Y=1.025 $X2=5.5
+ $Y2=1.212
r58 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.5 $Y=1.025 $X2=5.5
+ $Y2=0.56
r59 1 19 16.5763 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=5.475 $Y=1.41
+ $X2=5.475 $Y2=1.212
r60 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.475 $Y=1.41
+ $X2=5.475 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_2%VPWR 1 2 3 4 5 6 21 25 31 35 39 41 43 48
+ 49 51 52 54 55 56 58 70 78 83 86 90
c100 58 0 1.28647e-19 $X=0.54 $Y=2.72
r101 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r102 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r103 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r104 81 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r105 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r106 78 89 4.04153 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=6.095 $Y=2.72
+ $X2=6.267 $Y2=2.72
r107 78 80 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.095 $Y=2.72
+ $X2=5.75 $Y2=2.72
r108 77 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r109 77 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=3.91 $Y2=2.72
r110 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r111 74 86 13.2376 $w=1.7e-07 $l=3.3e-07 $layer=LI1_cond $X=4.385 $Y=2.72
+ $X2=4.055 $Y2=2.72
r112 74 76 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=4.385 $Y=2.72
+ $X2=4.83 $Y2=2.72
r113 73 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r114 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r115 70 86 13.2376 $w=1.7e-07 $l=3.3e-07 $layer=LI1_cond $X=3.725 $Y=2.72
+ $X2=4.055 $Y2=2.72
r116 70 72 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.725 $Y=2.72
+ $X2=3.45 $Y2=2.72
r117 69 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r118 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r119 66 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r120 66 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r121 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r122 63 83 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.815 $Y=2.72
+ $X2=0.677 $Y2=2.72
r123 63 65 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=0.815 $Y=2.72
+ $X2=1.61 $Y2=2.72
r124 58 83 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=0.54 $Y=2.72
+ $X2=0.677 $Y2=2.72
r125 58 60 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.54 $Y=2.72
+ $X2=0.23 $Y2=2.72
r126 56 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r127 56 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r128 54 76 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.155 $Y=2.72
+ $X2=4.83 $Y2=2.72
r129 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=2.72
+ $X2=5.24 $Y2=2.72
r130 53 80 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=5.325 $Y=2.72
+ $X2=5.75 $Y2=2.72
r131 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.325 $Y=2.72
+ $X2=5.24 $Y2=2.72
r132 51 68 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.655 $Y=2.72
+ $X2=2.53 $Y2=2.72
r133 51 52 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.655 $Y=2.72
+ $X2=2.805 $Y2=2.72
r134 50 72 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.955 $Y=2.72
+ $X2=3.45 $Y2=2.72
r135 50 52 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.955 $Y=2.72
+ $X2=2.805 $Y2=2.72
r136 48 65 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r137 48 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.845 $Y=2.72
+ $X2=1.93 $Y2=2.72
r138 47 68 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.015 $Y=2.72
+ $X2=2.53 $Y2=2.72
r139 47 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=2.72
+ $X2=1.93 $Y2=2.72
r140 43 46 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=6.22 $Y=1.66
+ $X2=6.22 $Y2=2.34
r141 41 89 3.10164 $w=2.5e-07 $l=1.05924e-07 $layer=LI1_cond $X=6.22 $Y=2.635
+ $X2=6.267 $Y2=2.72
r142 41 46 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=6.22 $Y=2.635
+ $X2=6.22 $Y2=2.34
r143 37 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.24 $Y=2.635
+ $X2=5.24 $Y2=2.72
r144 37 39 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.24 $Y=2.635
+ $X2=5.24 $Y2=2
r145 33 86 2.7357 $w=6.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=2.635
+ $X2=4.055 $Y2=2.72
r146 33 35 11.5077 $w=6.58e-07 $l=6.35e-07 $layer=LI1_cond $X=4.055 $Y=2.635
+ $X2=4.055 $Y2=2
r147 29 52 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.805 $Y=2.635
+ $X2=2.805 $Y2=2.72
r148 29 31 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=2.805 $Y=2.635
+ $X2=2.805 $Y2=2
r149 25 28 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.93 $Y=1.66
+ $X2=1.93 $Y2=2.34
r150 23 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=2.635
+ $X2=1.93 $Y2=2.72
r151 23 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.93 $Y=2.635
+ $X2=1.93 $Y2=2.34
r152 19 83 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.677 $Y=2.635
+ $X2=0.677 $Y2=2.72
r153 19 21 11.5244 $w=2.73e-07 $l=2.75e-07 $layer=LI1_cond $X=0.677 $Y=2.635
+ $X2=0.677 $Y2=2.36
r154 6 46 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.035
+ $Y=1.485 $X2=6.18 $Y2=2.34
r155 6 43 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=6.035
+ $Y=1.485 $X2=6.18 $Y2=1.66
r156 5 39 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.095
+ $Y=1.485 $X2=5.24 $Y2=2
r157 4 35 150 $w=1.7e-07 $l=8.02185e-07 $layer=licon1_PDIFF $count=4 $X=3.665
+ $Y=1.485 $X2=4.25 $Y2=2
r158 3 31 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.725
+ $Y=1.485 $X2=2.87 $Y2=2
r159 2 28 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.93 $Y2=2.34
r160 2 25 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.93 $Y2=1.66
r161 1 21 600 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.065 $X2=0.73 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_2%Y 1 2 3 4 5 18 22 24 28 30 31 34 36 38
+ 40 42 44 47 48
c99 18 0 1.7445e-19 $X=2.4 $Y=0.74
r100 47 48 0.553288 $w=4.41e-07 $l=2e-08 $layer=LI1_cond $X=3.875 $Y=1.37
+ $X2=3.895 $Y2=1.37
r101 38 46 2.73777 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=5.685 $Y=1.665
+ $X2=5.685 $Y2=1.555
r102 38 40 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=5.685 $Y=1.665
+ $X2=5.685 $Y2=2.34
r103 37 44 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=4.935 $Y=1.555
+ $X2=4.745 $Y2=1.555
r104 36 46 4.72888 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=5.495 $Y=1.555
+ $X2=5.685 $Y2=1.555
r105 36 37 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=5.495 $Y=1.555
+ $X2=4.935 $Y2=1.555
r106 32 44 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=4.745 $Y=1.665
+ $X2=4.745 $Y2=1.555
r107 32 34 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=4.745 $Y=1.665
+ $X2=4.745 $Y2=2.34
r108 31 48 7.21215 $w=4.41e-07 $l=2.48948e-07 $layer=LI1_cond $X=4.045 $Y=1.555
+ $X2=3.895 $Y2=1.37
r109 30 44 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=4.555 $Y=1.555
+ $X2=4.745 $Y2=1.555
r110 30 31 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=4.555 $Y=1.555
+ $X2=4.045 $Y2=1.555
r111 26 47 15.4921 $w=4.41e-07 $l=6.91954e-07 $layer=LI1_cond $X=3.315 $Y=1.665
+ $X2=3.875 $Y2=1.37
r112 26 28 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=3.315 $Y=1.665
+ $X2=3.315 $Y2=2.34
r113 25 42 3.29167 $w=2.2e-07 $l=2.23e-07 $layer=LI1_cond $X=2.63 $Y=1.555
+ $X2=2.407 $Y2=1.555
r114 24 26 8.31873 $w=4.41e-07 $l=2.38747e-07 $layer=LI1_cond $X=3.125 $Y=1.555
+ $X2=3.315 $Y2=1.665
r115 24 25 25.93 $w=2.18e-07 $l=4.95e-07 $layer=LI1_cond $X=3.125 $Y=1.555
+ $X2=2.63 $Y2=1.555
r116 20 42 3.2688 $w=3.72e-07 $l=1.41492e-07 $layer=LI1_cond $X=2.335 $Y=1.665
+ $X2=2.407 $Y2=1.555
r117 20 22 4.60977 $w=2.98e-07 $l=1.2e-07 $layer=LI1_cond $X=2.335 $Y=1.665
+ $X2=2.335 $Y2=1.785
r118 16 42 3.2688 $w=3.72e-07 $l=1.1e-07 $layer=LI1_cond $X=2.407 $Y=1.445
+ $X2=2.407 $Y2=1.555
r119 16 18 18.2578 $w=4.43e-07 $l=7.05e-07 $layer=LI1_cond $X=2.407 $Y=1.445
+ $X2=2.407 $Y2=0.74
r120 5 46 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=1.485 $X2=5.71 $Y2=1.66
r121 5 40 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=1.485 $X2=5.71 $Y2=2.34
r122 4 44 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.625
+ $Y=1.485 $X2=4.77 $Y2=1.66
r123 4 34 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.625
+ $Y=1.485 $X2=4.77 $Y2=2.34
r124 3 26 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.195
+ $Y=1.485 $X2=3.34 $Y2=1.66
r125 3 28 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.195
+ $Y=1.485 $X2=3.34 $Y2=2.34
r126 2 22 300 $w=1.7e-07 $l=3.65377e-07 $layer=licon1_PDIFF $count=2 $X=2.255
+ $Y=1.485 $X2=2.4 $Y2=1.785
r127 1 18 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=2.265
+ $Y=0.235 $X2=2.4 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_2%VGND 1 2 9 13 16 17 18 20 33 34 37
r71 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r72 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r73 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r74 30 31 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r75 28 31 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=5.29
+ $Y2=0
r76 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r77 27 30 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=5.29
+ $Y2=0
r78 27 28 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r79 25 37 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.665
+ $Y2=0
r80 25 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=1.15
+ $Y2=0
r81 20 37 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.665
+ $Y2=0
r82 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r83 18 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r84 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r85 16 30 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.625 $Y=0 $X2=5.29
+ $Y2=0
r86 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.625 $Y=0 $X2=5.71
+ $Y2=0
r87 15 33 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=5.795 $Y=0 $X2=6.21
+ $Y2=0
r88 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.795 $Y=0 $X2=5.71
+ $Y2=0
r89 11 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.71 $Y=0.085
+ $X2=5.71 $Y2=0
r90 11 13 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.71 $Y=0.085
+ $X2=5.71 $Y2=0.4
r91 7 37 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=0.085
+ $X2=0.665 $Y2=0
r92 7 9 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.665 $Y=0.085
+ $X2=0.665 $Y2=0.38
r93 2 13 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.575
+ $Y=0.235 $X2=5.71 $Y2=0.4
r94 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_361_47# 1 2 3 14 19
r25 17 19 4.03881 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=0.42
+ $X2=2.015 $Y2=0.42
r26 12 14 47.0998 $w=2.28e-07 $l=9.4e-07 $layer=LI1_cond $X=2.87 $Y=0.37
+ $X2=3.81 $Y2=0.37
r27 12 19 42.8408 $w=2.28e-07 $l=8.55e-07 $layer=LI1_cond $X=2.87 $Y=0.37
+ $X2=2.015 $Y2=0.37
r28 3 14 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.675
+ $Y=0.235 $X2=3.81 $Y2=0.4
r29 2 12 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.735
+ $Y=0.235 $X2=2.87 $Y2=0.4
r30 1 17 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.93 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_641_47# 1 2 11
c24 11 0 1.91072e-19 $X=4.77 $Y=0.74
r25 8 11 65.9197 $w=2.48e-07 $l=1.43e-06 $layer=LI1_cond $X=3.34 $Y=0.78
+ $X2=4.77 $Y2=0.78
r26 2 11 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.635
+ $Y=0.235 $X2=4.77 $Y2=0.74
r27 1 8 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.205
+ $Y=0.235 $X2=3.34 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_841_47# 1 2 3 10 14 15 16 20
r37 18 20 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.155 $Y=0.735
+ $X2=6.155 $Y2=0.4
r38 17 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.405 $Y=0.82
+ $X2=5.28 $Y2=0.82
r39 16 18 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=5.965 $Y=0.82
+ $X2=6.155 $Y2=0.735
r40 16 17 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.965 $Y=0.82
+ $X2=5.405 $Y2=0.82
r41 15 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.28 $Y=0.735
+ $X2=5.28 $Y2=0.82
r42 14 23 3.27362 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=5.28 $Y=0.485
+ $X2=5.28 $Y2=0.37
r43 14 15 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=5.28 $Y=0.485
+ $X2=5.28 $Y2=0.735
r44 10 23 3.55828 $w=2.3e-07 $l=1.25e-07 $layer=LI1_cond $X=5.155 $Y=0.37
+ $X2=5.28 $Y2=0.37
r45 10 12 41.3376 $w=2.28e-07 $l=8.25e-07 $layer=LI1_cond $X=5.155 $Y=0.37
+ $X2=4.33 $Y2=0.37
r46 3 20 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=6.045
+ $Y=0.235 $X2=6.18 $Y2=0.4
r47 2 25 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=5.105
+ $Y=0.235 $X2=5.24 $Y2=0.74
r48 2 23 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.105
+ $Y=0.235 $X2=5.24 $Y2=0.4
r49 1 12 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=4.205
+ $Y=0.235 $X2=4.33 $Y2=0.4
.ends

