* NGSPICE file created from sky130_fd_sc_hdll__or2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__or2_1 A B VGND VNB VPB VPWR X
M1000 VPWR A a_128_297# VPB phighvt w=420000u l=180000u
+  ad=3.057e+11p pd=2.71e+06u as=9.66e+10p ps=1.3e+06u
M1001 a_128_297# B a_38_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1002 a_38_297# B VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=3.307e+11p ps=3.43e+06u
M1003 X a_38_297# VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=0p ps=0u
M1004 VGND A a_38_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_38_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.5e+11p pd=2.7e+06u as=0p ps=0u
.ends

