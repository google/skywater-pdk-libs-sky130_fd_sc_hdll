* File: sky130_fd_sc_hdll__nor4_2.pex.spice
* Created: Thu Aug 27 19:17:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR4_2%A 1 3 4 6 7 9 10 12 13 20 24
c37 13 0 1.93357e-19 $X=0.66 $Y=1.105
r38 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.01 $Y2=1.202
r39 18 20 43.1263 $w=3.8e-07 $l=3.4e-07 $layer=POLY_cond $X=0.645 $Y=1.202
+ $X2=0.985 $Y2=1.202
r40 18 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.645
+ $Y=1.16 $X2=0.645 $Y2=1.16
r41 16 18 16.4895 $w=3.8e-07 $l=1.3e-07 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.645 $Y2=1.202
r42 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.49 $Y=1.202
+ $X2=0.515 $Y2=1.202
r43 13 24 5.28139 $w=2.08e-07 $l=1e-07 $layer=LI1_cond $X=0.745 $Y=1.18
+ $X2=0.645 $Y2=1.18
r44 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=1.202
r45 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=0.56
r46 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r47 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r48 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r49 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r50 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.202
r51 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_2%B 1 3 4 6 7 9 10 12 13 20 23
c41 20 0 1.93357e-19 $X=1.925 $Y=1.202
r42 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.925 $Y=1.202
+ $X2=1.95 $Y2=1.202
r43 18 20 31.7105 $w=3.8e-07 $l=2.5e-07 $layer=POLY_cond $X=1.675 $Y=1.202
+ $X2=1.925 $Y2=1.202
r44 18 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.675
+ $Y=1.16 $X2=1.675 $Y2=1.16
r45 16 18 27.9053 $w=3.8e-07 $l=2.2e-07 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.675 $Y2=1.202
r46 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.43 $Y=1.202
+ $X2=1.455 $Y2=1.202
r47 13 23 7.92208 $w=2.08e-07 $l=1.5e-07 $layer=LI1_cond $X=1.765 $Y=1.18
+ $X2=1.615 $Y2=1.18
r48 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=1.202
r49 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=0.56
r50 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r51 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r52 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r53 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r54 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=1.202
r55 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995 $X2=1.43
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_2%C 1 3 4 6 7 9 10 12 13 19 20 23
c38 19 0 1.64881e-19 $X=3.19 $Y=1.16
r39 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.425 $Y=1.202
+ $X2=3.45 $Y2=1.202
r40 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=3.19 $Y=1.202
+ $X2=3.425 $Y2=1.202
r41 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.19
+ $Y=1.16 $X2=3.19 $Y2=1.16
r42 16 18 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=2.955 $Y=1.202
+ $X2=3.19 $Y2=1.202
r43 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=2.93 $Y=1.202
+ $X2=2.955 $Y2=1.202
r44 13 19 22.974 $w=2.08e-07 $l=4.35e-07 $layer=LI1_cond $X=2.755 $Y=1.18
+ $X2=3.19 $Y2=1.18
r45 13 23 0.528139 $w=2.08e-07 $l=1e-08 $layer=LI1_cond $X=2.755 $Y=1.18
+ $X2=2.745 $Y2=1.18
r46 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.45 $Y=0.995
+ $X2=3.45 $Y2=1.202
r47 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.45 $Y=0.995
+ $X2=3.45 $Y2=0.56
r48 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.425 $Y=1.41
+ $X2=3.425 $Y2=1.202
r49 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.425 $Y=1.41
+ $X2=3.425 $Y2=1.985
r50 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.955 $Y=1.41
+ $X2=2.955 $Y2=1.202
r51 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.955 $Y=1.41
+ $X2=2.955 $Y2=1.985
r52 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.93 $Y=0.995
+ $X2=2.93 $Y2=1.202
r53 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.93 $Y=0.995 $X2=2.93
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_2%D 1 3 4 6 7 9 10 12 13 19 20 23
c43 20 0 1.64881e-19 $X=4.365 $Y=1.202
r44 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.365 $Y=1.202
+ $X2=4.39 $Y2=1.202
r45 18 20 32.3447 $w=3.8e-07 $l=2.55e-07 $layer=POLY_cond $X=4.11 $Y=1.202
+ $X2=4.365 $Y2=1.202
r46 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.11
+ $Y=1.16 $X2=4.11 $Y2=1.16
r47 16 18 27.2711 $w=3.8e-07 $l=2.15e-07 $layer=POLY_cond $X=3.895 $Y=1.202
+ $X2=4.11 $Y2=1.202
r48 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.87 $Y=1.202
+ $X2=3.895 $Y2=1.202
r49 13 19 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=3.775 $Y=1.18
+ $X2=4.11 $Y2=1.18
r50 13 23 0.528139 $w=2.08e-07 $l=1e-08 $layer=LI1_cond $X=3.775 $Y=1.18
+ $X2=3.765 $Y2=1.18
r51 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.39 $Y=0.995
+ $X2=4.39 $Y2=1.202
r52 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.39 $Y=0.995
+ $X2=4.39 $Y2=0.56
r53 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.365 $Y=1.41
+ $X2=4.365 $Y2=1.202
r54 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.365 $Y=1.41
+ $X2=4.365 $Y2=1.985
r55 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.895 $Y=1.41
+ $X2=3.895 $Y2=1.202
r56 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.895 $Y=1.41
+ $X2=3.895 $Y2=1.985
r57 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.87 $Y=0.995
+ $X2=3.87 $Y2=1.202
r58 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.87 $Y=0.995 $X2=3.87
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_2%A_27_297# 1 2 3 10 12 14 18 20 27 29
r36 21 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=1.54
+ $X2=1.22 $Y2=1.54
r37 20 29 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=1.54
+ $X2=2.16 $Y2=1.54
r38 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.035 $Y=1.54
+ $X2=1.345 $Y2=1.54
r39 16 27 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=1.625
+ $X2=1.22 $Y2=1.54
r40 16 18 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.22 $Y=1.625
+ $X2=1.22 $Y2=2.3
r41 15 25 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.405 $Y=1.54
+ $X2=0.277 $Y2=1.54
r42 14 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=1.54
+ $X2=1.22 $Y2=1.54
r43 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=1.54
+ $X2=0.405 $Y2=1.54
r44 10 25 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.277 $Y=1.625
+ $X2=0.277 $Y2=1.54
r45 10 12 30.5058 $w=2.53e-07 $l=6.75e-07 $layer=LI1_cond $X=0.277 $Y=1.625
+ $X2=0.277 $Y2=2.3
r46 3 29 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=1.62
r47 2 27 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.62
r48 2 18 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.3
r49 1 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r50 1 12 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_2%VPWR 1 8 10 17 18 21 24
r46 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r47 17 18 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r48 15 18 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=4.83 $Y2=2.72
r49 15 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 14 17 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=4.83 $Y2=2.72
r51 14 15 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r52 12 21 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=0.75 $Y2=2.72
r53 12 14 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=1.15 $Y2=2.72
r54 10 22 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r55 10 24 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r56 6 21 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r57 6 8 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.75 $Y=2.635 $X2=0.75
+ $Y2=1.96
r58 1 8 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_2%A_309_297# 1 2 9 11 12 15
r19 13 15 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.19 $Y=2.295
+ $X2=3.19 $Y2=1.96
r20 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.065 $Y=2.38
+ $X2=3.19 $Y2=2.295
r21 11 12 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=3.065 $Y=2.38
+ $X2=1.815 $Y2=2.38
r22 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.69 $Y=2.295
+ $X2=1.815 $Y2=2.38
r23 7 9 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.69 $Y=2.295
+ $X2=1.69 $Y2=1.96
r24 2 15 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.045
+ $Y=1.485 $X2=3.19 $Y2=1.96
r25 1 9 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_2%A_515_297# 1 2 3 12 14 15 16 20 23
r36 18 20 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.6 $Y=2.295
+ $X2=4.6 $Y2=1.96
r37 17 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.785 $Y=2.38
+ $X2=3.66 $Y2=2.38
r38 16 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.475 $Y=2.38
+ $X2=4.6 $Y2=2.295
r39 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.475 $Y=2.38
+ $X2=3.785 $Y2=2.38
r40 15 27 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.66 $Y=2.295
+ $X2=3.66 $Y2=2.38
r41 14 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.66 $Y=1.625
+ $X2=3.66 $Y2=1.54
r42 14 15 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=3.66 $Y=1.625
+ $X2=3.66 $Y2=2.295
r43 13 23 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.845 $Y=1.54
+ $X2=2.72 $Y2=1.54
r44 12 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.535 $Y=1.54
+ $X2=3.66 $Y2=1.54
r45 12 13 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.535 $Y=1.54
+ $X2=2.845 $Y2=1.54
r46 3 20 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.455
+ $Y=1.485 $X2=4.6 $Y2=1.96
r47 2 27 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.485 $X2=3.66 $Y2=2.3
r48 2 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.485 $X2=3.66 $Y2=1.62
r49 1 23 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.575
+ $Y=1.485 $X2=2.72 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_2%Y 1 2 3 4 5 18 20 21 24 26 30 32 36 40 42
+ 44 45 46 48 50 53
r103 50 53 2.6797 $w=3.35e-07 $l=9e-08 $layer=LI1_cond $X=4.782 $Y=0.815
+ $X2=4.782 $Y2=0.905
r104 50 53 0.516019 $w=3.33e-07 $l=1.5e-08 $layer=LI1_cond $X=4.782 $Y=0.92
+ $X2=4.782 $Y2=0.905
r105 49 50 18.4047 $w=3.33e-07 $l=5.35e-07 $layer=LI1_cond $X=4.782 $Y=1.455
+ $X2=4.782 $Y2=0.92
r106 43 46 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.33 $Y=0.815
+ $X2=4.14 $Y2=0.815
r107 42 50 4.97233 $w=1.8e-07 $l=1.67e-07 $layer=LI1_cond $X=4.615 $Y=0.815
+ $X2=4.782 $Y2=0.815
r108 42 43 17.5606 $w=1.78e-07 $l=2.85e-07 $layer=LI1_cond $X=4.615 $Y=0.815
+ $X2=4.33 $Y2=0.815
r109 41 48 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.29 $Y=1.54
+ $X2=4.165 $Y2=1.54
r110 40 49 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=4.615 $Y=1.54
+ $X2=4.782 $Y2=1.455
r111 40 41 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.615 $Y=1.54
+ $X2=4.29 $Y2=1.54
r112 34 46 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=4.14 $Y=0.725 $X2=4.14
+ $Y2=0.815
r113 34 36 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.14 $Y=0.725
+ $X2=4.14 $Y2=0.39
r114 33 45 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.39 $Y=0.815
+ $X2=3.2 $Y2=0.815
r115 32 46 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.95 $Y=0.815
+ $X2=4.14 $Y2=0.815
r116 32 33 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.95 $Y=0.815
+ $X2=3.39 $Y2=0.815
r117 28 45 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=3.2 $Y=0.725 $X2=3.2
+ $Y2=0.815
r118 28 30 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.2 $Y=0.725
+ $X2=3.2 $Y2=0.39
r119 27 44 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.89 $Y=0.815
+ $X2=1.7 $Y2=0.815
r120 26 45 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.01 $Y=0.815
+ $X2=3.2 $Y2=0.815
r121 26 27 69.0101 $w=1.78e-07 $l=1.12e-06 $layer=LI1_cond $X=3.01 $Y=0.815
+ $X2=1.89 $Y2=0.815
r122 22 44 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=1.7 $Y=0.725 $X2=1.7
+ $Y2=0.815
r123 22 24 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.7 $Y=0.725
+ $X2=1.7 $Y2=0.39
r124 20 44 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.51 $Y=0.815
+ $X2=1.7 $Y2=0.815
r125 20 21 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.51 $Y=0.815
+ $X2=0.95 $Y2=0.815
r126 16 21 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=0.76 $Y=0.725
+ $X2=0.95 $Y2=0.815
r127 16 18 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.76 $Y=0.725
+ $X2=0.76 $Y2=0.39
r128 5 48 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.985
+ $Y=1.485 $X2=4.13 $Y2=1.62
r129 4 36 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.945
+ $Y=0.235 $X2=4.13 $Y2=0.39
r130 3 30 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.005
+ $Y=0.235 $X2=3.19 $Y2=0.39
r131 2 24 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.505
+ $Y=0.235 $X2=1.69 $Y2=0.39
r132 1 18 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_2%VGND 1 2 3 4 5 6 19 21 23 27 31 33 35 38 39
+ 40 51 59 63 69 72
r77 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r78 68 69 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.72 $Y=0.235
+ $X2=2.805 $Y2=0.235
r79 65 68 3.55086 $w=6.38e-07 $l=1.9e-07 $layer=LI1_cond $X=2.53 $Y=0.235
+ $X2=2.72 $Y2=0.235
r80 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r81 62 65 6.91483 $w=6.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=0.235
+ $X2=2.53 $Y2=0.235
r82 62 63 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.235
+ $X2=2.075 $Y2=0.235
r83 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r84 54 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r85 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r86 51 71 4.17994 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=4.515 $Y=0 $X2=4.787
+ $Y2=0
r87 51 53 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.515 $Y=0 $X2=4.37
+ $Y2=0
r88 50 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r89 50 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r90 49 69 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=2.805
+ $Y2=0
r91 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r92 46 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r93 46 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r94 45 63 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.075
+ $Y2=0
r95 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r96 43 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.22
+ $Y2=0
r97 43 45 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=2.07
+ $Y2=0
r98 40 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r99 40 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r100 38 49 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.575 $Y=0
+ $X2=3.45 $Y2=0
r101 38 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.575 $Y=0 $X2=3.66
+ $Y2=0
r102 37 53 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.745 $Y=0
+ $X2=4.37 $Y2=0
r103 37 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.745 $Y=0 $X2=3.66
+ $Y2=0
r104 33 71 3.2579 $w=2.9e-07 $l=1.64085e-07 $layer=LI1_cond $X=4.66 $Y=0.085
+ $X2=4.787 $Y2=0
r105 33 35 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=4.66 $Y=0.085
+ $X2=4.66 $Y2=0.39
r106 29 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.66 $Y=0.085
+ $X2=3.66 $Y2=0
r107 29 31 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.66 $Y=0.085
+ $X2=3.66 $Y2=0.39
r108 25 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r109 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.39
r110 24 56 4.28094 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r111 23 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.22
+ $Y2=0
r112 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=0
+ $X2=0.365 $Y2=0
r113 19 56 3.0411 $w=2.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.182 $Y2=0
r114 19 21 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.227 $Y2=0.39
r115 6 35 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.465
+ $Y=0.235 $X2=4.6 $Y2=0.39
r116 5 31 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.525
+ $Y=0.235 $X2=3.66 $Y2=0.39
r117 4 68 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=2.575
+ $Y=0.235 $X2=2.72 $Y2=0.39
r118 3 62 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.16 $Y2=0.39
r119 2 27 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.235 $X2=1.22 $Y2=0.39
r120 1 21 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

