* File: sky130_fd_sc_hdll__mux2_4.spice
* Created: Thu Aug 27 19:10:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__mux2_4.pex.spice"
.subckt sky130_fd_sc_hdll__mux2_4  VNB VPB S A0 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A0	A0
* S	S
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_S_M1010_g N_A_27_47#_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.125125 AS=0.2015 PD=1.035 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75005.2 A=0.0975 P=1.6 MULT=1
MM1015 A_226_47# N_A_27_47#_M1015_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.65
+ AD=0.27625 AS=0.125125 PD=1.5 PS=1.035 NRD=68.304 NRS=20.304 M=1 R=4.33333
+ SA=75000.8 SB=75004.6 A=0.0975 P=1.6 MULT=1
MM1011 N_A_424_297#_M1011_d N_A0_M1011_g A_226_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.27625 PD=1.02 PS=1.5 NRD=3.684 NRS=68.304 M=1 R=4.33333
+ SA=75001.8 SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1006 A_530_47# N_A1_M1006_g N_A_424_297#_M1011_d VNB NSHORT L=0.15 W=0.65
+ AD=0.290875 AS=0.12025 PD=1.545 PS=1.02 NRD=72.456 NRS=12.912 M=1 R=4.33333
+ SA=75002.3 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_S_M1008_g A_530_47# VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.290875 PD=0.97 PS=1.545 NRD=0 NRS=72.456 M=1 R=4.33333 SA=75003.3
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1003_d N_A_424_297#_M1003_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.8
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1005 N_X_M1003_d N_A_424_297#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75004.3
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1009_d N_A_424_297#_M1009_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.7
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1017 N_X_M1009_d N_A_424_297#_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.169 PD=0.97 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75005.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_S_M1004_g N_A_27_47#_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1725 AS=0.27 PD=1.345 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1016 N_A_222_297#_M1016_d N_A_27_47#_M1016_g N_VPWR_M1004_d VPB PHIGHVT L=0.18
+ W=1 AD=0.29 AS=0.1725 PD=2.58 PS=1.345 NRD=2.955 NRS=11.8003 M=1 R=5.55556
+ SA=90000.7 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1001 N_A_424_297#_M1001_d N_A0_M1001_g N_A_334_297#_M1001_s VPB PHIGHVT L=0.18
+ W=1 AD=0.17 AS=0.27 PD=1.34 PS=2.54 NRD=6.8753 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1014 N_A_222_297#_M1014_d N_A1_M1014_g N_A_424_297#_M1001_d VPB PHIGHVT L=0.18
+ W=1 AD=0.31 AS=0.17 PD=2.62 PS=1.34 NRD=4.9053 NRS=4.9053 M=1 R=5.55556
+ SA=90000.7 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_S_M1012_g N_A_334_297#_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1012_d N_A_424_297#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A_424_297#_M1002_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1002_d N_A_424_297#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1013_d N_A_424_297#_M1013_g N_X_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90000.2 A=0.18 P=2.36 MULT=1
DX18_noxref VNB VPB NWDIODE A=10.2078 P=15.93
*
.include "sky130_fd_sc_hdll__mux2_4.pxi.spice"
*
.ends
*
*
