* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nor4_6 A B C D VGND VNB VPB VPWR Y
X0 a_1263_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND D Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_1263_297# C a_685_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Y D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_685_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 a_685_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 a_1263_297# C a_685_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 VGND D Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_27_297# B a_685_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_685_297# C a_1263_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 Y D a_1263_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 Y D a_1263_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 VGND D Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_685_297# C a_1263_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_1263_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X31 a_27_297# B a_685_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X32 a_1263_297# C a_685_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 a_685_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X35 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 a_27_297# B a_685_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X37 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X38 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 Y D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X40 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X41 a_1263_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X42 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X43 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X44 a_685_297# C a_1263_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X45 Y D a_1263_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X46 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X47 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
