* File: sky130_fd_sc_hdll__nand4bb_4.pex.spice
* Created: Thu Aug 27 19:15:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_N 1 3 4 6 7 8 14
c28 1 0 7.16581e-20 $X=0.495 $Y=1.41
r29 14 15 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r30 12 14 33.1044 $w=3.64e-07 $l=2.5e-07 $layer=POLY_cond $X=0.245 $Y=1.202
+ $X2=0.495 $Y2=1.202
r31 7 8 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.215 $Y=1.16
+ $X2=0.215 $Y2=1.53
r32 7 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r33 4 15 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r34 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r35 1 14 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r36 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_4%B_N 1 3 4 6 7 8 13
r33 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r34 7 8 8.90524 $w=4.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.805 $Y=1.19
+ $X2=0.805 $Y2=1.53
r35 7 13 0.785757 $w=4.38e-07 $l=3e-08 $layer=LI1_cond $X=0.805 $Y=1.19
+ $X2=0.805 $Y2=1.16
r36 4 12 39.2931 $w=2.55e-07 $l=1.72337e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.94 $Y2=1.16
r37 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=0.56
r38 1 12 51.486 $w=2.55e-07 $l=2.62202e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.94 $Y2=1.16
r39 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_27_47# 1 2 7 9 10 12 13 15 18 20 22 25
+ 27 29 32 36 40 42 43 44 45 49 53 56 66
c142 66 0 4.77784e-20 $X=3.745 $Y=1.202
r143 66 67 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=3.745 $Y=1.202
+ $X2=3.77 $Y2=1.202
r144 65 66 64.997 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=3.3 $Y=1.202
+ $X2=3.745 $Y2=1.202
r145 64 65 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=3.275 $Y=1.202
+ $X2=3.3 $Y2=1.202
r146 61 62 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.805 $Y=1.202
+ $X2=2.83 $Y2=1.202
r147 60 61 64.997 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=2.36 $Y=1.202
+ $X2=2.805 $Y2=1.202
r148 59 60 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.335 $Y=1.202
+ $X2=2.36 $Y2=1.202
r149 56 59 14.6061 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=2.235 $Y=1.16
+ $X2=2.335 $Y2=1.202
r150 53 64 35.0545 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=3.035 $Y=1.202
+ $X2=3.275 $Y2=1.202
r151 53 62 29.9424 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.035 $Y=1.202
+ $X2=2.83 $Y2=1.202
r152 50 56 142.512 $w=3.3e-07 $l=8.15e-07 $layer=POLY_cond $X=1.42 $Y=1.16
+ $X2=2.235 $Y2=1.16
r153 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.42
+ $Y=1.16 $X2=1.42 $Y2=1.16
r154 47 49 23.2347 $w=3.08e-07 $l=6.25e-07 $layer=LI1_cond $X=1.35 $Y=1.785
+ $X2=1.35 $Y2=1.16
r155 46 49 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=1.35 $Y=0.805
+ $X2=1.35 $Y2=1.16
r156 44 47 7.28659 $w=1.95e-07 $l=1.97636e-07 $layer=LI1_cond $X=1.195 $Y=1.882
+ $X2=1.35 $Y2=1.785
r157 44 45 46.9231 $w=1.93e-07 $l=8.25e-07 $layer=LI1_cond $X=1.195 $Y=1.882
+ $X2=0.37 $Y2=1.882
r158 42 46 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=1.195 $Y=0.72
+ $X2=1.35 $Y2=0.805
r159 42 43 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.195 $Y=0.72
+ $X2=0.345 $Y2=0.72
r160 38 45 7.13288 $w=1.95e-07 $l=1.85642e-07 $layer=LI1_cond $X=0.227 $Y=1.98
+ $X2=0.37 $Y2=1.882
r161 38 40 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=0.227 $Y=1.98
+ $X2=0.227 $Y2=2.275
r162 34 43 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.345 $Y2=0.72
r163 34 36 7.75683 $w=2.58e-07 $l=1.75e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.215 $Y2=0.46
r164 30 67 21.2229 $w=1.5e-07 $l=1.77e-07 $layer=POLY_cond $X=3.77 $Y=1.025
+ $X2=3.77 $Y2=1.202
r165 30 32 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.77 $Y=1.025
+ $X2=3.77 $Y2=0.56
r166 27 66 16.9318 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.745 $Y=1.41
+ $X2=3.745 $Y2=1.202
r167 27 29 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.745 $Y=1.41
+ $X2=3.745 $Y2=1.985
r168 23 65 21.2229 $w=1.5e-07 $l=1.77e-07 $layer=POLY_cond $X=3.3 $Y=1.025
+ $X2=3.3 $Y2=1.202
r169 23 25 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.3 $Y=1.025
+ $X2=3.3 $Y2=0.56
r170 20 64 16.9318 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.275 $Y=1.41
+ $X2=3.275 $Y2=1.202
r171 20 22 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.275 $Y=1.41
+ $X2=3.275 $Y2=1.985
r172 16 62 21.2229 $w=1.5e-07 $l=1.77e-07 $layer=POLY_cond $X=2.83 $Y=1.025
+ $X2=2.83 $Y2=1.202
r173 16 18 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.83 $Y=1.025
+ $X2=2.83 $Y2=0.56
r174 13 61 16.9318 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.805 $Y=1.41
+ $X2=2.805 $Y2=1.202
r175 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.805 $Y=1.41
+ $X2=2.805 $Y2=1.985
r176 10 60 21.2229 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.36 $Y=0.995
+ $X2=2.36 $Y2=1.202
r177 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.36 $Y=0.995
+ $X2=2.36 $Y2=0.56
r178 7 59 16.9318 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.335 $Y=1.41
+ $X2=2.335 $Y2=1.202
r179 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.335 $Y=1.41
+ $X2=2.335 $Y2=1.985
r180 2 40 600 $w=1.7e-07 $l=8.50206e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.275
r181 1 36 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_206_47# 1 2 9 11 13 16 18 20 23 25 27
+ 28 30 33 35 39 44 46 47 48 51 54 68 69
c136 68 0 1.56636e-19 $X=5.39 $Y=1.16
c137 54 0 1.50024e-19 $X=4.415 $Y=1.19
c138 51 0 4.77784e-20 $X=1.88 $Y=1.19
c139 35 0 7.16581e-20 $X=1.675 $Y=2.307
r140 69 70 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=5.625 $Y=1.217
+ $X2=5.65 $Y2=1.217
r141 67 69 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=5.39 $Y=1.217
+ $X2=5.625 $Y2=1.217
r142 67 68 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.39
+ $Y=1.16 $X2=5.39 $Y2=1.16
r143 65 67 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=5.155 $Y=1.217
+ $X2=5.39 $Y2=1.217
r144 64 65 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=5.13 $Y=1.217
+ $X2=5.155 $Y2=1.217
r145 63 64 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=4.685 $Y=1.217
+ $X2=5.13 $Y2=1.217
r146 62 63 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=4.66 $Y=1.217
+ $X2=4.685 $Y2=1.217
r147 60 62 30.2171 $w=3.27e-07 $l=2.05e-07 $layer=POLY_cond $X=4.455 $Y=1.217
+ $X2=4.66 $Y2=1.217
r148 58 60 35.3761 $w=3.27e-07 $l=2.4e-07 $layer=POLY_cond $X=4.215 $Y=1.217
+ $X2=4.455 $Y2=1.217
r149 57 58 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=4.19 $Y=1.217
+ $X2=4.215 $Y2=1.217
r150 55 68 54.0682 $w=1.98e-07 $l=9.75e-07 $layer=LI1_cond $X=4.415 $Y=1.175
+ $X2=5.39 $Y2=1.175
r151 55 60 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.455
+ $Y=1.16 $X2=4.455 $Y2=1.16
r152 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.415 $Y=1.19
+ $X2=4.415 $Y2=1.19
r153 51 75 6.01275 $w=2.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.88 $Y=1.19
+ $X2=1.76 $Y2=1.19
r154 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.88 $Y=1.19
+ $X2=1.88 $Y2=1.19
r155 48 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.025 $Y=1.19
+ $X2=1.88 $Y2=1.19
r156 47 54 0.137923 $w=2.3e-07 $l=1.8e-07 $layer=MET1_cond $X=4.235 $Y=1.19
+ $X2=4.415 $Y2=1.19
r157 47 48 2.73514 $w=1.4e-07 $l=2.21e-06 $layer=MET1_cond $X=4.235 $Y=1.19
+ $X2=2.025 $Y2=1.19
r158 45 75 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.76 $Y=1.305
+ $X2=1.76 $Y2=1.19
r159 45 46 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.76 $Y=1.305
+ $X2=1.76 $Y2=2.15
r160 44 75 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.76 $Y=1.075
+ $X2=1.76 $Y2=1.19
r161 43 44 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.76 $Y=0.465
+ $X2=1.76 $Y2=1.075
r162 39 43 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.675 $Y=0.36
+ $X2=1.76 $Y2=0.465
r163 39 41 20.8615 $w=2.08e-07 $l=3.95e-07 $layer=LI1_cond $X=1.675 $Y=0.36
+ $X2=1.28 $Y2=0.36
r164 35 46 7.64049 $w=3.15e-07 $l=1.94921e-07 $layer=LI1_cond $X=1.675 $Y=2.307
+ $X2=1.76 $Y2=2.15
r165 35 37 17.3781 $w=3.13e-07 $l=4.75e-07 $layer=LI1_cond $X=1.675 $Y=2.307
+ $X2=1.2 $Y2=2.307
r166 31 70 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.65 $Y=1.025
+ $X2=5.65 $Y2=1.217
r167 31 33 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.65 $Y=1.025
+ $X2=5.65 $Y2=0.56
r168 28 69 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.625 $Y=1.41
+ $X2=5.625 $Y2=1.217
r169 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.625 $Y=1.41
+ $X2=5.625 $Y2=1.985
r170 25 65 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.155 $Y=1.41
+ $X2=5.155 $Y2=1.217
r171 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.155 $Y=1.41
+ $X2=5.155 $Y2=1.985
r172 21 64 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.13 $Y=1.025
+ $X2=5.13 $Y2=1.217
r173 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.13 $Y=1.025
+ $X2=5.13 $Y2=0.56
r174 18 63 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.685 $Y=1.41
+ $X2=4.685 $Y2=1.217
r175 18 20 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.685 $Y=1.41
+ $X2=4.685 $Y2=1.985
r176 14 62 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.66 $Y=1.025
+ $X2=4.66 $Y2=1.217
r177 14 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.66 $Y=1.025
+ $X2=4.66 $Y2=0.56
r178 11 58 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.215 $Y=1.41
+ $X2=4.215 $Y2=1.217
r179 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.215 $Y=1.41
+ $X2=4.215 $Y2=1.985
r180 7 57 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.19 $Y=1.025
+ $X2=4.19 $Y2=1.217
r181 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.19 $Y=1.025
+ $X2=4.19 $Y2=0.56
r182 2 37 600 $w=1.7e-07 $l=9.14631e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.33
r183 1 41 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.235 $X2=1.28 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_4%C 1 3 6 8 10 13 15 17 20 22 24 27 29 30
+ 31 32 37 50 51 56 60 63 65
c76 50 0 1.87801e-19 $X=7.82 $Y=1.16
c77 37 0 1.56636e-19 $X=6.545 $Y=1.16
r78 63 65 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=7.125 $Y=1.175
+ $X2=7.585 $Y2=1.175
r79 51 52 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=8.055 $Y=1.217
+ $X2=8.08 $Y2=1.217
r80 49 51 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=7.82 $Y=1.217
+ $X2=8.055 $Y2=1.217
r81 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.82
+ $Y=1.16 $X2=7.82 $Y2=1.16
r82 47 49 30.9541 $w=3.27e-07 $l=2.1e-07 $layer=POLY_cond $X=7.61 $Y=1.217
+ $X2=7.82 $Y2=1.217
r83 46 47 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=7.585 $Y=1.217
+ $X2=7.61 $Y2=1.217
r84 45 46 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=7.14 $Y=1.217
+ $X2=7.585 $Y2=1.217
r85 44 45 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=7.115 $Y=1.217
+ $X2=7.14 $Y2=1.217
r86 43 44 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=6.67 $Y=1.217
+ $X2=7.115 $Y2=1.217
r87 42 43 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=6.645 $Y=1.217
+ $X2=6.67 $Y2=1.217
r88 40 56 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=6.38 $Y=1.175
+ $X2=6.205 $Y2=1.175
r89 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.38
+ $Y=1.16 $X2=6.38 $Y2=1.16
r90 37 42 16.3472 $w=3.27e-07 $l=1.253e-07 $layer=POLY_cond $X=6.545 $Y=1.16
+ $X2=6.645 $Y2=1.217
r91 37 39 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.545 $Y=1.16
+ $X2=6.38 $Y2=1.16
r92 32 50 11.6455 $w=1.98e-07 $l=2.1e-07 $layer=LI1_cond $X=7.61 $Y=1.175
+ $X2=7.82 $Y2=1.175
r93 32 65 1.38636 $w=1.98e-07 $l=2.5e-08 $layer=LI1_cond $X=7.61 $Y=1.175
+ $X2=7.585 $Y2=1.175
r94 31 63 1.38636 $w=1.98e-07 $l=2.5e-08 $layer=LI1_cond $X=7.1 $Y=1.175
+ $X2=7.125 $Y2=1.175
r95 31 60 24.1227 $w=1.98e-07 $l=4.35e-07 $layer=LI1_cond $X=7.1 $Y=1.175
+ $X2=6.665 $Y2=1.175
r96 30 60 4.15909 $w=1.98e-07 $l=7.5e-08 $layer=LI1_cond $X=6.59 $Y=1.175
+ $X2=6.665 $Y2=1.175
r97 30 40 11.6455 $w=1.98e-07 $l=2.1e-07 $layer=LI1_cond $X=6.59 $Y=1.175
+ $X2=6.38 $Y2=1.175
r98 29 56 4.15909 $w=1.98e-07 $l=7.5e-08 $layer=LI1_cond $X=6.13 $Y=1.175
+ $X2=6.205 $Y2=1.175
r99 25 52 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=8.08 $Y=1.025
+ $X2=8.08 $Y2=1.217
r100 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.08 $Y=1.025
+ $X2=8.08 $Y2=0.56
r101 22 51 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=8.055 $Y=1.41
+ $X2=8.055 $Y2=1.217
r102 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.055 $Y=1.41
+ $X2=8.055 $Y2=1.985
r103 18 47 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.61 $Y=1.025
+ $X2=7.61 $Y2=1.217
r104 18 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.61 $Y=1.025
+ $X2=7.61 $Y2=0.56
r105 15 46 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.585 $Y=1.41
+ $X2=7.585 $Y2=1.217
r106 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.585 $Y=1.41
+ $X2=7.585 $Y2=1.985
r107 11 45 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.14 $Y=1.025
+ $X2=7.14 $Y2=1.217
r108 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.14 $Y=1.025
+ $X2=7.14 $Y2=0.56
r109 8 44 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.115 $Y=1.41
+ $X2=7.115 $Y2=1.217
r110 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.115 $Y=1.41
+ $X2=7.115 $Y2=1.985
r111 4 43 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.67 $Y=1.025
+ $X2=6.67 $Y2=1.217
r112 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.67 $Y=1.025
+ $X2=6.67 $Y2=0.56
r113 1 42 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.645 $Y=1.41
+ $X2=6.645 $Y2=1.217
r114 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.645 $Y=1.41
+ $X2=6.645 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_4%D 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 32 37 39 56 59 63
c74 37 0 1.87801e-19 $X=10.035 $Y=1.165
r75 51 52 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=9.91 $Y=1.217
+ $X2=9.935 $Y2=1.217
r76 50 51 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=9.465 $Y=1.217
+ $X2=9.91 $Y2=1.217
r77 49 50 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=9.44 $Y=1.217
+ $X2=9.465 $Y2=1.217
r78 48 49 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=8.995 $Y=1.217
+ $X2=9.44 $Y2=1.217
r79 47 48 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=8.97 $Y=1.217
+ $X2=8.995 $Y2=1.217
r80 45 47 30.9541 $w=3.27e-07 $l=2.1e-07 $layer=POLY_cond $X=8.76 $Y=1.217
+ $X2=8.97 $Y2=1.217
r81 45 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.76
+ $Y=1.16 $X2=8.76 $Y2=1.16
r82 43 45 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=8.525 $Y=1.217
+ $X2=8.76 $Y2=1.217
r83 42 43 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=8.5 $Y=1.217
+ $X2=8.525 $Y2=1.217
r84 39 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.17
+ $Y=1.16 $X2=10.17 $Y2=1.16
r85 37 52 15.8716 $w=3.27e-07 $l=1.23288e-07 $layer=POLY_cond $X=10.035 $Y=1.165
+ $X2=9.935 $Y2=1.217
r86 37 39 28.9223 $w=2.8e-07 $l=1.35e-07 $layer=POLY_cond $X=10.035 $Y=1.165
+ $X2=10.17 $Y2=1.165
r87 32 63 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=10.21 $Y=1.175
+ $X2=10.17 $Y2=1.175
r88 31 63 26.0636 $w=1.98e-07 $l=4.7e-07 $layer=LI1_cond $X=9.7 $Y=1.175
+ $X2=10.17 $Y2=1.175
r89 31 59 27.45 $w=1.98e-07 $l=4.95e-07 $layer=LI1_cond $X=9.7 $Y=1.175
+ $X2=9.205 $Y2=1.175
r90 30 59 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=9.19 $Y=1.175
+ $X2=9.205 $Y2=1.175
r91 30 56 27.7273 $w=1.98e-07 $l=5e-07 $layer=LI1_cond $X=9.19 $Y=1.175 $X2=8.69
+ $Y2=1.175
r92 29 56 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=8.68 $Y=1.175
+ $X2=8.69 $Y2=1.175
r93 26 52 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=9.935 $Y=1.41
+ $X2=9.935 $Y2=1.217
r94 26 28 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.935 $Y=1.41
+ $X2=9.935 $Y2=1.985
r95 22 51 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=9.91 $Y=1.025
+ $X2=9.91 $Y2=1.217
r96 22 24 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.91 $Y=1.025
+ $X2=9.91 $Y2=0.56
r97 19 50 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=9.465 $Y=1.41
+ $X2=9.465 $Y2=1.217
r98 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.465 $Y=1.41
+ $X2=9.465 $Y2=1.985
r99 15 49 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=9.44 $Y=1.025
+ $X2=9.44 $Y2=1.217
r100 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.44 $Y=1.025
+ $X2=9.44 $Y2=0.56
r101 12 48 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=8.995 $Y=1.41
+ $X2=8.995 $Y2=1.217
r102 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.995 $Y=1.41
+ $X2=8.995 $Y2=1.985
r103 8 47 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=8.97 $Y=1.025
+ $X2=8.97 $Y2=1.217
r104 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.97 $Y=1.025
+ $X2=8.97 $Y2=0.56
r105 5 43 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=8.525 $Y=1.41
+ $X2=8.525 $Y2=1.217
r106 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.525 $Y=1.41
+ $X2=8.525 $Y2=1.985
r107 1 42 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=8.5 $Y=1.025
+ $X2=8.5 $Y2=1.217
r108 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.5 $Y=1.025 $X2=8.5
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_4%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 43 45 49
+ 53 57 61 65 69 71 73 78 79 81 82 84 85 87 88 89 91 96 101 110 124 129 132 135
+ 138 141 145
r165 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r166 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r167 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r168 136 139 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r169 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r170 132 133 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r171 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r172 127 145 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.35 $Y2=2.72
r173 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r174 124 144 4.09173 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=10.085 $Y=2.72
+ $X2=10.332 $Y2=2.72
r175 124 126 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=10.085 $Y=2.72
+ $X2=9.89 $Y2=2.72
r176 123 127 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r177 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r178 120 123 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r179 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r180 117 120 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r181 117 142 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=6.21 $Y2=2.72
r182 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r183 114 141 13.0174 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=6.465 $Y=2.72
+ $X2=6.145 $Y2=2.72
r184 114 116 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=6.465 $Y=2.72
+ $X2=7.13 $Y2=2.72
r185 113 142 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r186 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r187 110 141 13.0174 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=5.825 $Y=2.72
+ $X2=6.145 $Y2=2.72
r188 110 112 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.825 $Y=2.72
+ $X2=5.75 $Y2=2.72
r189 109 113 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r190 109 139 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=3.91 $Y2=2.72
r191 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r192 106 138 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.065 $Y=2.72
+ $X2=3.98 $Y2=2.72
r193 106 108 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=4.065 $Y=2.72
+ $X2=4.83 $Y2=2.72
r194 105 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r195 105 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r196 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r197 102 132 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.185 $Y=2.72
+ $X2=2.1 $Y2=2.72
r198 102 104 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.185 $Y=2.72
+ $X2=2.53 $Y2=2.72
r199 101 135 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.825 $Y=2.72
+ $X2=2.975 $Y2=2.72
r200 101 104 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.825 $Y=2.72
+ $X2=2.53 $Y2=2.72
r201 100 133 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r202 100 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r203 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r204 97 129 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.815 $Y=2.72
+ $X2=0.677 $Y2=2.72
r205 97 99 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=2.72
+ $X2=1.15 $Y2=2.72
r206 96 132 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=2.72
+ $X2=2.1 $Y2=2.72
r207 96 99 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=2.015 $Y=2.72
+ $X2=1.15 $Y2=2.72
r208 91 129 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=0.54 $Y=2.72
+ $X2=0.677 $Y2=2.72
r209 91 93 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.54 $Y=2.72
+ $X2=0.23 $Y2=2.72
r210 89 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r211 89 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r212 87 122 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=9.145 $Y=2.72
+ $X2=8.97 $Y2=2.72
r213 87 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.145 $Y=2.72
+ $X2=9.23 $Y2=2.72
r214 86 126 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=9.315 $Y=2.72
+ $X2=9.89 $Y2=2.72
r215 86 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.315 $Y=2.72
+ $X2=9.23 $Y2=2.72
r216 84 119 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.205 $Y=2.72
+ $X2=8.05 $Y2=2.72
r217 84 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.205 $Y=2.72
+ $X2=8.29 $Y2=2.72
r218 83 122 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=8.375 $Y=2.72
+ $X2=8.97 $Y2=2.72
r219 83 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.375 $Y=2.72
+ $X2=8.29 $Y2=2.72
r220 81 116 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.265 $Y=2.72
+ $X2=7.13 $Y2=2.72
r221 81 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.265 $Y=2.72
+ $X2=7.35 $Y2=2.72
r222 80 119 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=7.435 $Y=2.72
+ $X2=8.05 $Y2=2.72
r223 80 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.435 $Y=2.72
+ $X2=7.35 $Y2=2.72
r224 78 108 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.835 $Y=2.72
+ $X2=4.83 $Y2=2.72
r225 78 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.835 $Y=2.72
+ $X2=4.92 $Y2=2.72
r226 77 112 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=5.005 $Y=2.72
+ $X2=5.75 $Y2=2.72
r227 77 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=2.72
+ $X2=4.92 $Y2=2.72
r228 73 76 28.4968 $w=2.73e-07 $l=6.8e-07 $layer=LI1_cond $X=10.222 $Y=1.66
+ $X2=10.222 $Y2=2.34
r229 71 144 3.23031 $w=2.75e-07 $l=1.46458e-07 $layer=LI1_cond $X=10.222
+ $Y=2.635 $X2=10.332 $Y2=2.72
r230 71 76 12.3626 $w=2.73e-07 $l=2.95e-07 $layer=LI1_cond $X=10.222 $Y=2.635
+ $X2=10.222 $Y2=2.34
r231 67 88 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.23 $Y=2.635
+ $X2=9.23 $Y2=2.72
r232 67 69 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=9.23 $Y=2.635
+ $X2=9.23 $Y2=2
r233 63 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.29 $Y=2.635
+ $X2=8.29 $Y2=2.72
r234 63 65 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.29 $Y=2.635
+ $X2=8.29 $Y2=2
r235 59 82 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.35 $Y=2.635
+ $X2=7.35 $Y2=2.72
r236 59 61 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.35 $Y=2.635
+ $X2=7.35 $Y2=2
r237 55 141 2.66764 $w=6.4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.145 $Y=2.635
+ $X2=6.145 $Y2=2.72
r238 55 57 11.8673 $w=6.38e-07 $l=6.35e-07 $layer=LI1_cond $X=6.145 $Y=2.635
+ $X2=6.145 $Y2=2
r239 51 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.92 $Y=2.635
+ $X2=4.92 $Y2=2.72
r240 51 53 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.92 $Y=2.635
+ $X2=4.92 $Y2=2
r241 47 138 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.98 $Y=2.635
+ $X2=3.98 $Y2=2.72
r242 47 49 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.98 $Y=2.635
+ $X2=3.98 $Y2=2
r243 46 135 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.125 $Y=2.72
+ $X2=2.975 $Y2=2.72
r244 45 138 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.895 $Y=2.72
+ $X2=3.98 $Y2=2.72
r245 45 46 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.895 $Y=2.72
+ $X2=3.125 $Y2=2.72
r246 41 135 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=2.635
+ $X2=2.975 $Y2=2.72
r247 41 43 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=2.975 $Y=2.635
+ $X2=2.975 $Y2=2
r248 37 40 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.1 $Y=1.66 $X2=2.1
+ $Y2=2.34
r249 35 132 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=2.635
+ $X2=2.1 $Y2=2.72
r250 35 40 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.1 $Y=2.635
+ $X2=2.1 $Y2=2.34
r251 31 129 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.677 $Y=2.635
+ $X2=0.677 $Y2=2.72
r252 31 33 11.5244 $w=2.73e-07 $l=2.75e-07 $layer=LI1_cond $X=0.677 $Y=2.635
+ $X2=0.677 $Y2=2.36
r253 10 76 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.025
+ $Y=1.485 $X2=10.17 $Y2=2.34
r254 10 73 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=10.025
+ $Y=1.485 $X2=10.17 $Y2=1.66
r255 9 69 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=9.085
+ $Y=1.485 $X2=9.23 $Y2=2
r256 8 65 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=8.145
+ $Y=1.485 $X2=8.29 $Y2=2
r257 7 61 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=7.205
+ $Y=1.485 $X2=7.35 $Y2=2
r258 6 57 150 $w=1.7e-07 $l=7.54785e-07 $layer=licon1_PDIFF $count=4 $X=5.715
+ $Y=1.485 $X2=6.255 $Y2=2
r259 5 53 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.775
+ $Y=1.485 $X2=4.92 $Y2=2
r260 4 49 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.835
+ $Y=1.485 $X2=3.98 $Y2=2
r261 3 43 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.895
+ $Y=1.485 $X2=3.04 $Y2=2
r262 2 40 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.975
+ $Y=1.485 $X2=2.1 $Y2=2.34
r263 2 37 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.975
+ $Y=1.485 $X2=2.1 $Y2=1.66
r264 1 33 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_4%Y 1 2 3 4 5 6 7 8 9 10 31 39 41 42 45 49
+ 51 52 55 57 61 63 67 69 73 75 77 79 82 84 86 88 91 92 97 108
c192 97 0 1.23116e-19 $X=3.84 $Y=0.905
r193 92 108 1.83343 $w=2.18e-07 $l=3.5e-08 $layer=LI1_cond $X=3.87 $Y=1.555
+ $X2=3.905 $Y2=1.555
r194 91 97 2.94404 $w=3.5e-07 $l=1.25e-07 $layer=LI1_cond $X=3.84 $Y=0.78
+ $X2=3.84 $Y2=0.905
r195 91 92 13.3593 $w=5.18e-07 $l=5.25e-07 $layer=LI1_cond $X=3.84 $Y=0.92
+ $X2=3.84 $Y2=1.445
r196 91 97 0.493904 $w=3.48e-07 $l=1.5e-08 $layer=LI1_cond $X=3.84 $Y=0.92
+ $X2=3.84 $Y2=0.905
r197 77 90 2.73777 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=9.675 $Y=1.665
+ $X2=9.675 $Y2=1.555
r198 77 79 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=9.675 $Y=1.665
+ $X2=9.675 $Y2=2.34
r199 76 88 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=8.925 $Y=1.555
+ $X2=8.735 $Y2=1.555
r200 75 90 4.72888 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=9.485 $Y=1.555
+ $X2=9.675 $Y2=1.555
r201 75 76 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=9.485 $Y=1.555
+ $X2=8.925 $Y2=1.555
r202 71 88 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=8.735 $Y=1.665
+ $X2=8.735 $Y2=1.555
r203 71 73 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=8.735 $Y=1.665
+ $X2=8.735 $Y2=2.34
r204 70 86 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=7.985 $Y=1.555
+ $X2=7.795 $Y2=1.555
r205 69 88 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=8.545 $Y=1.555
+ $X2=8.735 $Y2=1.555
r206 69 70 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=8.545 $Y=1.555
+ $X2=7.985 $Y2=1.555
r207 65 86 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=7.795 $Y=1.665
+ $X2=7.795 $Y2=1.555
r208 65 67 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=7.795 $Y=1.665
+ $X2=7.795 $Y2=2.34
r209 64 84 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=7.045 $Y=1.555
+ $X2=6.855 $Y2=1.555
r210 63 86 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=7.605 $Y=1.555
+ $X2=7.795 $Y2=1.555
r211 63 64 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=7.605 $Y=1.555
+ $X2=7.045 $Y2=1.555
r212 59 84 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=6.855 $Y=1.665
+ $X2=6.855 $Y2=1.555
r213 59 61 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=6.855 $Y=1.665
+ $X2=6.855 $Y2=2.34
r214 58 82 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=5.555 $Y=1.555
+ $X2=5.365 $Y2=1.555
r215 57 84 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=6.665 $Y=1.555
+ $X2=6.855 $Y2=1.555
r216 57 58 58.146 $w=2.18e-07 $l=1.11e-06 $layer=LI1_cond $X=6.665 $Y=1.555
+ $X2=5.555 $Y2=1.555
r217 53 82 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=5.365 $Y=1.665
+ $X2=5.365 $Y2=1.555
r218 53 55 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=5.365 $Y=1.665
+ $X2=5.365 $Y2=2.34
r219 51 82 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=5.175 $Y=1.555
+ $X2=5.365 $Y2=1.555
r220 51 52 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=5.175 $Y=1.555
+ $X2=4.615 $Y2=1.555
r221 47 52 9.95292 $w=2.18e-07 $l=1.9e-07 $layer=LI1_cond $X=4.425 $Y=1.555
+ $X2=4.615 $Y2=1.555
r222 47 108 27.2396 $w=2.18e-07 $l=5.2e-07 $layer=LI1_cond $X=4.425 $Y=1.555
+ $X2=3.905 $Y2=1.555
r223 47 49 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=4.425 $Y=1.665
+ $X2=4.425 $Y2=2.34
r224 43 92 18.5962 $w=2.18e-07 $l=3.55e-07 $layer=LI1_cond $X=3.485 $Y=1.555
+ $X2=3.84 $Y2=1.555
r225 43 45 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=3.485 $Y=1.665
+ $X2=3.485 $Y2=2.34
r226 41 43 9.95292 $w=2.18e-07 $l=1.9e-07 $layer=LI1_cond $X=3.295 $Y=1.555
+ $X2=3.485 $Y2=1.555
r227 41 42 33.5256 $w=2.18e-07 $l=6.4e-07 $layer=LI1_cond $X=3.295 $Y=1.555
+ $X2=2.655 $Y2=1.555
r228 37 42 7.02845 $w=2.2e-07 $l=1.97484e-07 $layer=LI1_cond $X=2.505 $Y=1.665
+ $X2=2.655 $Y2=1.555
r229 37 39 4.60977 $w=2.98e-07 $l=1.2e-07 $layer=LI1_cond $X=2.505 $Y=1.665
+ $X2=2.505 $Y2=1.785
r230 33 36 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=2.57 $Y=0.78
+ $X2=3.51 $Y2=0.78
r231 31 91 4.12165 $w=2.5e-07 $l=1.75e-07 $layer=LI1_cond $X=3.665 $Y=0.78
+ $X2=3.84 $Y2=0.78
r232 31 36 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=3.665 $Y=0.78
+ $X2=3.51 $Y2=0.78
r233 10 90 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=9.555
+ $Y=1.485 $X2=9.7 $Y2=1.66
r234 10 79 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=9.555
+ $Y=1.485 $X2=9.7 $Y2=2.34
r235 9 88 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=8.615
+ $Y=1.485 $X2=8.76 $Y2=1.66
r236 9 73 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=8.615
+ $Y=1.485 $X2=8.76 $Y2=2.34
r237 8 86 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=7.675
+ $Y=1.485 $X2=7.82 $Y2=1.66
r238 8 67 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.675
+ $Y=1.485 $X2=7.82 $Y2=2.34
r239 7 84 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=6.735
+ $Y=1.485 $X2=6.88 $Y2=1.66
r240 7 61 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.735
+ $Y=1.485 $X2=6.88 $Y2=2.34
r241 6 82 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.245
+ $Y=1.485 $X2=5.39 $Y2=1.66
r242 6 55 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.245
+ $Y=1.485 $X2=5.39 $Y2=2.34
r243 5 47 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.305
+ $Y=1.485 $X2=4.45 $Y2=1.66
r244 5 49 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.305
+ $Y=1.485 $X2=4.45 $Y2=2.34
r245 4 43 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.365
+ $Y=1.485 $X2=3.51 $Y2=1.66
r246 4 45 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.365
+ $Y=1.485 $X2=3.51 $Y2=2.34
r247 3 39 300 $w=1.7e-07 $l=3.65377e-07 $layer=licon1_PDIFF $count=2 $X=2.425
+ $Y=1.485 $X2=2.57 $Y2=1.785
r248 2 36 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.375
+ $Y=0.235 $X2=3.51 $Y2=0.74
r249 1 33 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=2.435
+ $Y=0.235 $X2=2.57 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_4%VGND 1 2 3 12 16 19 20 22 23 24 26 42 43
+ 47
r98 47 50 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0 $X2=0.705
+ $Y2=0.38
r99 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r100 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r101 40 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.35 $Y2=0
r102 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r103 37 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=9.43
+ $Y2=0
r104 36 37 1.09412 $w=1.7e-07 $l=1.445e-06 $layer=mcon $count=8 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r105 34 37 2.09423 $w=4.8e-07 $l=7.36e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=8.51
+ $Y2=0
r106 34 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r107 33 36 480.171 $w=1.68e-07 $l=7.36e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=8.51
+ $Y2=0
r108 33 34 1.09412 $w=1.7e-07 $l=1.445e-06 $layer=mcon $count=8 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r109 31 47 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r110 31 33 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r111 26 47 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r112 26 28 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r113 24 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r114 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r115 22 39 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=9.535 $Y=0
+ $X2=9.43 $Y2=0
r116 22 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.535 $Y=0 $X2=9.7
+ $Y2=0
r117 21 42 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=9.865 $Y=0
+ $X2=10.35 $Y2=0
r118 21 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.865 $Y=0 $X2=9.7
+ $Y2=0
r119 19 36 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=8.595 $Y=0 $X2=8.51
+ $Y2=0
r120 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.595 $Y=0 $X2=8.76
+ $Y2=0
r121 18 39 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=8.925 $Y=0
+ $X2=9.43 $Y2=0
r122 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.925 $Y=0 $X2=8.76
+ $Y2=0
r123 14 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.7 $Y=0.085 $X2=9.7
+ $Y2=0
r124 14 16 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=9.7 $Y=0.085
+ $X2=9.7 $Y2=0.4
r125 10 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.76 $Y=0.085
+ $X2=8.76 $Y2=0
r126 10 12 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=8.76 $Y=0.085
+ $X2=8.76 $Y2=0.4
r127 3 16 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=9.515
+ $Y=0.235 $X2=9.7 $Y2=0.4
r128 2 12 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=8.575
+ $Y=0.235 $X2=8.76 $Y2=0.4
r129 1 50 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_395_47# 1 2 3 4 5 18 20 28
r43 26 28 47.0998 $w=2.28e-07 $l=9.4e-07 $layer=LI1_cond $X=4.92 $Y=0.37
+ $X2=5.86 $Y2=0.37
r44 24 26 47.0998 $w=2.28e-07 $l=9.4e-07 $layer=LI1_cond $X=3.98 $Y=0.37
+ $X2=4.92 $Y2=0.37
r45 22 24 47.0998 $w=2.28e-07 $l=9.4e-07 $layer=LI1_cond $X=3.04 $Y=0.37
+ $X2=3.98 $Y2=0.37
r46 20 22 42.8408 $w=2.28e-07 $l=8.55e-07 $layer=LI1_cond $X=2.185 $Y=0.37
+ $X2=3.04 $Y2=0.37
r47 16 20 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.1 $Y=0.485
+ $X2=2.185 $Y2=0.37
r48 16 18 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.1 $Y=0.485
+ $X2=2.1 $Y2=0.74
r49 5 28 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.725
+ $Y=0.235 $X2=5.86 $Y2=0.4
r50 4 26 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=4.735
+ $Y=0.235 $X2=4.92 $Y2=0.4
r51 3 24 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.845
+ $Y=0.235 $X2=3.98 $Y2=0.4
r52 2 22 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.905
+ $Y=0.235 $X2=3.04 $Y2=0.4
r53 1 18 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.1 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_853_47# 1 2 3 4 21
r36 19 21 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=6.905 $Y=0.78
+ $X2=7.845 $Y2=0.78
r37 17 19 69.838 $w=2.48e-07 $l=1.515e-06 $layer=LI1_cond $X=5.39 $Y=0.78
+ $X2=6.905 $Y2=0.78
r38 14 17 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=4.45 $Y=0.78
+ $X2=5.39 $Y2=0.78
r39 4 21 182 $w=1.7e-07 $l=5.79504e-07 $layer=licon1_NDIFF $count=1 $X=7.685
+ $Y=0.235 $X2=7.845 $Y2=0.74
r40 3 19 182 $w=1.7e-07 $l=5.79504e-07 $layer=licon1_NDIFF $count=1 $X=6.745
+ $Y=0.235 $X2=6.905 $Y2=0.74
r41 2 17 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=5.205
+ $Y=0.235 $X2=5.39 $Y2=0.74
r42 1 14 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=4.265
+ $Y=0.235 $X2=4.45 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_1251_47# 1 2 3 4 5 16 26 30
r32 28 30 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=9.215 $Y=0.74
+ $X2=10.12 $Y2=0.74
r33 26 28 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=8.375 $Y=0.74
+ $X2=9.215 $Y2=0.74
r34 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.29 $Y=0.655
+ $X2=8.375 $Y2=0.74
r35 23 25 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=8.29 $Y=0.655
+ $X2=8.29 $Y2=0.535
r36 22 25 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=8.29 $Y=0.485 $X2=8.29
+ $Y2=0.535
r37 18 21 47.0998 $w=2.28e-07 $l=9.4e-07 $layer=LI1_cond $X=6.43 $Y=0.37
+ $X2=7.37 $Y2=0.37
r38 16 22 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=8.205 $Y=0.37
+ $X2=8.29 $Y2=0.485
r39 16 21 41.8387 $w=2.28e-07 $l=8.35e-07 $layer=LI1_cond $X=8.205 $Y=0.37
+ $X2=7.37 $Y2=0.37
r40 5 30 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=9.985
+ $Y=0.235 $X2=10.12 $Y2=0.74
r41 4 28 182 $w=1.7e-07 $l=5.83845e-07 $layer=licon1_NDIFF $count=1 $X=9.045
+ $Y=0.235 $X2=9.215 $Y2=0.74
r42 3 25 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=8.155
+ $Y=0.235 $X2=8.29 $Y2=0.535
r43 2 21 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=7.215
+ $Y=0.235 $X2=7.37 $Y2=0.4
r44 1 18 182 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_NDIFF $count=1 $X=6.255
+ $Y=0.235 $X2=6.43 $Y2=0.4
.ends

