# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__clkinv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkinv_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.42000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  5.328000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  1.615000 1.075000  2.415000 1.120000 ;
        RECT  1.615000 1.120000 11.135000 1.260000 ;
        RECT  1.615000 1.260000  2.415000 1.305000 ;
        RECT 10.285000 1.075000 11.135000 1.120000 ;
        RECT 10.285000 1.260000 11.135000 1.305000 ;
    END
  END A
  PIN VGND
    ANTENNADIFFAREA  1.228500 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.420000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  3.895000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.420000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  4.928900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.625000 1.455000 11.630000 1.665000 ;
        RECT  0.625000 1.665000  0.880000 2.465000 ;
        RECT  1.585000 1.665000  1.840000 2.450000 ;
        RECT  2.575000 0.280000  2.800000 1.415000 ;
        RECT  2.575000 1.415000  9.705000 1.455000 ;
        RECT  2.575000 1.665000  2.800000 2.465000 ;
        RECT  3.505000 0.280000  3.760000 1.415000 ;
        RECT  3.505000 1.665000  3.760000 2.450000 ;
        RECT  4.465000 0.280000  4.705000 1.415000 ;
        RECT  4.465000 1.665000  4.705000 2.450000 ;
        RECT  5.455000 0.280000  5.805000 1.415000 ;
        RECT  5.455000 1.665000  5.830000 2.450000 ;
        RECT  6.575000 0.280000  6.825000 1.415000 ;
        RECT  6.575000 1.665000  6.825000 2.450000 ;
        RECT  7.535000 0.280000  7.785000 1.415000 ;
        RECT  7.535000 1.665000  7.785000 2.450000 ;
        RECT  8.495000 0.280000  8.745000 1.415000 ;
        RECT  8.495000 1.665000  8.745000 2.450000 ;
        RECT  9.455000 0.280000  9.705000 1.415000 ;
        RECT  9.455000 1.665000  9.705000 2.450000 ;
        RECT 10.415000 1.665000 10.655000 2.450000 ;
        RECT 11.375000 1.665000 11.630000 2.450000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.420000 0.085000 ;
      RECT  0.000000  2.635000 12.420000 2.805000 ;
      RECT  0.140000  1.495000  0.405000 2.635000 ;
      RECT  0.345000  0.895000  2.355000 1.275000 ;
      RECT  1.100000  1.835000  1.360000 2.635000 ;
      RECT  2.055000  0.085000  2.325000 0.610000 ;
      RECT  2.065000  1.835000  2.320000 2.635000 ;
      RECT  3.020000  0.085000  3.285000 0.610000 ;
      RECT  3.020000  1.835000  3.280000 2.635000 ;
      RECT  3.980000  0.085000  4.245000 0.610000 ;
      RECT  3.985000  1.835000  4.240000 2.635000 ;
      RECT  4.965000  0.085000  5.230000 0.610000 ;
      RECT  4.965000  1.835000  5.220000 2.635000 ;
      RECT  6.090000  0.085000  6.355000 0.610000 ;
      RECT  6.090000  1.835000  6.345000 2.120000 ;
      RECT  6.090000  2.120000  6.350000 2.635000 ;
      RECT  7.050000  0.085000  7.275000 0.610000 ;
      RECT  7.055000  1.835000  7.310000 2.635000 ;
      RECT  8.010000  0.085000  8.275000 0.610000 ;
      RECT  8.015000  1.835000  8.270000 2.635000 ;
      RECT  8.970000  0.085000  9.235000 0.610000 ;
      RECT  8.975000  1.835000  9.230000 2.635000 ;
      RECT  9.930000  0.085000 10.195000 0.610000 ;
      RECT  9.930000  0.895000 11.910000 1.275000 ;
      RECT  9.935000  1.835000 10.190000 2.635000 ;
      RECT 10.895000  1.835000 11.150000 2.635000 ;
      RECT 11.850000  1.835000 12.110000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.675000  1.105000  1.845000 1.275000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.185000  1.105000  2.355000 1.275000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.395000  1.105000 10.565000 1.275000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 10.905000  1.105000 11.075000 1.275000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinv_16
