* NGSPICE file created from sky130_fd_sc_hdll__o32ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 VGND A2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=1.0595e+12p pd=7.16e+06u as=1.469e+12p ps=1.232e+07u
M1001 a_27_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=8.3e+11p pd=7.66e+06u as=5.8e+11p ps=5.16e+06u
M1002 Y A3 a_525_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.7e+11p ps=7.74e+06u
M1003 a_27_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.81e+11p ps=4.08e+06u
M1004 VGND A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_807_297# VPB phighvt w=1e+06u l=180000u
+  ad=8.5e+11p pd=7.7e+06u as=5.8e+11p ps=5.16e+06u
M1007 Y B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_525_297# A2 a_807_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_807_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_807_297# A2 a_525_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_525_297# A3 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A3 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

