* File: sky130_fd_sc_hdll__xnor2_4.pex.spice
* Created: Thu Aug 27 19:29:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__XNOR2_4%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 50 51 52 54 55 60 63 64 78
+ 88 93
c203 88 0 6.90269e-20 $X=8.14 $Y=1.202
c204 51 0 1.5003e-19 $X=6.1 $Y=1.53
c205 50 0 1.87257e-19 $X=1.92 $Y=1.445
c206 22 0 1.98558e-19 $X=2.005 $Y=0.995
r207 88 89 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.14 $Y=1.202
+ $X2=8.165 $Y2=1.202
r208 85 86 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.645 $Y=1.202
+ $X2=7.67 $Y2=1.202
r209 84 85 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=7.2 $Y=1.202
+ $X2=7.645 $Y2=1.202
r210 83 84 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.175 $Y=1.202
+ $X2=7.2 $Y2=1.202
r211 80 81 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.705 $Y=1.202
+ $X2=6.73 $Y2=1.202
r212 78 79 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.98 $Y=1.202
+ $X2=2.005 $Y2=1.202
r213 76 78 20.0833 $w=3.72e-07 $l=1.55e-07 $layer=POLY_cond $X=1.825 $Y=1.202
+ $X2=1.98 $Y2=1.202
r214 76 77 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.825
+ $Y=1.16 $X2=1.825 $Y2=1.16
r215 74 76 40.8145 $w=3.72e-07 $l=3.15e-07 $layer=POLY_cond $X=1.51 $Y=1.202
+ $X2=1.825 $Y2=1.202
r216 73 74 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.485 $Y=1.202
+ $X2=1.51 $Y2=1.202
r217 72 73 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=1.04 $Y=1.202
+ $X2=1.485 $Y2=1.202
r218 71 72 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.015 $Y=1.202
+ $X2=1.04 $Y2=1.202
r219 70 93 27.45 $w=1.98e-07 $l=4.95e-07 $layer=LI1_cond $X=0.655 $Y=1.175
+ $X2=1.15 $Y2=1.175
r220 69 71 46.6452 $w=3.72e-07 $l=3.6e-07 $layer=POLY_cond $X=0.655 $Y=1.202
+ $X2=1.015 $Y2=1.202
r221 69 70 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.655
+ $Y=1.16 $X2=0.655 $Y2=1.16
r222 67 69 11.0134 $w=3.72e-07 $l=8.5e-08 $layer=POLY_cond $X=0.57 $Y=1.202
+ $X2=0.655 $Y2=1.202
r223 66 67 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.545 $Y=1.202
+ $X2=0.57 $Y2=1.202
r224 64 77 37.1545 $w=1.98e-07 $l=6.7e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=1.825 $Y2=1.175
r225 64 93 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=1.15 $Y2=1.175
r226 63 77 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=1.835 $Y=1.175
+ $X2=1.825 $Y2=1.175
r227 61 88 18.1398 $w=3.72e-07 $l=1.4e-07 $layer=POLY_cond $X=8 $Y=1.202
+ $X2=8.14 $Y2=1.202
r228 61 86 42.7581 $w=3.72e-07 $l=3.3e-07 $layer=POLY_cond $X=8 $Y=1.202
+ $X2=7.67 $Y2=1.202
r229 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8 $Y=1.16
+ $X2=8 $Y2=1.16
r230 58 83 44.7016 $w=3.72e-07 $l=3.45e-07 $layer=POLY_cond $X=6.83 $Y=1.202
+ $X2=7.175 $Y2=1.202
r231 58 81 12.957 $w=3.72e-07 $l=1e-07 $layer=POLY_cond $X=6.83 $Y=1.202
+ $X2=6.73 $Y2=1.202
r232 57 60 64.8818 $w=1.98e-07 $l=1.17e-06 $layer=LI1_cond $X=6.83 $Y=1.175
+ $X2=8 $Y2=1.175
r233 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.83
+ $Y=1.16 $X2=6.83 $Y2=1.16
r234 55 57 31.0545 $w=1.98e-07 $l=5.6e-07 $layer=LI1_cond $X=6.27 $Y=1.175
+ $X2=6.83 $Y2=1.175
r235 53 55 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=6.185 $Y=1.275
+ $X2=6.27 $Y2=1.175
r236 53 54 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.185 $Y=1.275
+ $X2=6.185 $Y2=1.445
r237 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.1 $Y=1.53
+ $X2=6.185 $Y2=1.445
r238 51 52 267.16 $w=1.68e-07 $l=4.095e-06 $layer=LI1_cond $X=6.1 $Y=1.53
+ $X2=2.005 $Y2=1.53
r239 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.92 $Y=1.445
+ $X2=2.005 $Y2=1.53
r240 49 63 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.92 $Y=1.275
+ $X2=1.835 $Y2=1.175
r241 49 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.92 $Y=1.275
+ $X2=1.92 $Y2=1.445
r242 46 89 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.165 $Y=0.995
+ $X2=8.165 $Y2=1.202
r243 46 48 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.165 $Y=0.995
+ $X2=8.165 $Y2=0.56
r244 43 88 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.14 $Y=1.41
+ $X2=8.14 $Y2=1.202
r245 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.14 $Y=1.41
+ $X2=8.14 $Y2=1.985
r246 40 86 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.67 $Y=1.41
+ $X2=7.67 $Y2=1.202
r247 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.67 $Y=1.41
+ $X2=7.67 $Y2=1.985
r248 37 85 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.645 $Y=0.995
+ $X2=7.645 $Y2=1.202
r249 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.645 $Y=0.995
+ $X2=7.645 $Y2=0.56
r250 34 84 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.2 $Y=1.41
+ $X2=7.2 $Y2=1.202
r251 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.2 $Y=1.41
+ $X2=7.2 $Y2=1.985
r252 31 83 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.175 $Y=0.995
+ $X2=7.175 $Y2=1.202
r253 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.175 $Y=0.995
+ $X2=7.175 $Y2=0.56
r254 28 81 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.73 $Y=1.41
+ $X2=6.73 $Y2=1.202
r255 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.73 $Y=1.41
+ $X2=6.73 $Y2=1.985
r256 25 80 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.705 $Y=0.995
+ $X2=6.705 $Y2=1.202
r257 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.705 $Y=0.995
+ $X2=6.705 $Y2=0.56
r258 22 79 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.005 $Y=0.995
+ $X2=2.005 $Y2=1.202
r259 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.005 $Y=0.995
+ $X2=2.005 $Y2=0.56
r260 19 78 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.98 $Y=1.41
+ $X2=1.98 $Y2=1.202
r261 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.98 $Y=1.41
+ $X2=1.98 $Y2=1.985
r262 16 74 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.51 $Y=1.41
+ $X2=1.51 $Y2=1.202
r263 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.51 $Y=1.41
+ $X2=1.51 $Y2=1.985
r264 13 73 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.485 $Y=0.995
+ $X2=1.485 $Y2=1.202
r265 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.485 $Y=0.995
+ $X2=1.485 $Y2=0.56
r266 10 72 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.04 $Y=1.41
+ $X2=1.04 $Y2=1.202
r267 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.04 $Y=1.41
+ $X2=1.04 $Y2=1.985
r268 7 71 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.015 $Y=0.995
+ $X2=1.015 $Y2=1.202
r269 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.015 $Y=0.995
+ $X2=1.015 $Y2=0.56
r270 4 67 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.57 $Y=1.41
+ $X2=0.57 $Y2=1.202
r271 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.57 $Y=1.41
+ $X2=0.57 $Y2=1.985
r272 1 66 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.545 $Y=0.995
+ $X2=0.545 $Y2=1.202
r273 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.545 $Y=0.995
+ $X2=0.545 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 63 74 77 84
c152 74 0 6.90269e-20 $X=5.715 $Y=1.16
c153 4 0 1.87257e-19 $X=2.45 $Y=1.41
r154 77 78 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.26 $Y=1.202
+ $X2=6.285 $Y2=1.202
r155 76 77 60.8979 $w=3.72e-07 $l=4.7e-07 $layer=POLY_cond $X=5.79 $Y=1.202
+ $X2=6.26 $Y2=1.202
r156 75 76 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.765 $Y=1.202
+ $X2=5.79 $Y2=1.202
r157 73 75 6.47849 $w=3.72e-07 $l=5e-08 $layer=POLY_cond $X=5.715 $Y=1.202
+ $X2=5.765 $Y2=1.202
r158 73 74 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.715
+ $Y=1.16 $X2=5.715 $Y2=1.16
r159 71 73 51.1801 $w=3.72e-07 $l=3.95e-07 $layer=POLY_cond $X=5.32 $Y=1.202
+ $X2=5.715 $Y2=1.202
r160 70 71 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.295 $Y=1.202
+ $X2=5.32 $Y2=1.202
r161 69 74 43.2545 $w=1.98e-07 $l=7.8e-07 $layer=LI1_cond $X=4.935 $Y=1.175
+ $X2=5.715 $Y2=1.175
r162 69 84 30.5 $w=1.98e-07 $l=5.5e-07 $layer=LI1_cond $X=4.935 $Y=1.175
+ $X2=4.385 $Y2=1.175
r163 68 70 46.6452 $w=3.72e-07 $l=3.6e-07 $layer=POLY_cond $X=4.935 $Y=1.202
+ $X2=5.295 $Y2=1.202
r164 68 69 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.935
+ $Y=1.16 $X2=4.935 $Y2=1.16
r165 66 68 11.0134 $w=3.72e-07 $l=8.5e-08 $layer=POLY_cond $X=4.85 $Y=1.202
+ $X2=4.935 $Y2=1.202
r166 65 66 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.825 $Y=1.202
+ $X2=4.85 $Y2=1.202
r167 63 64 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.86 $Y=1.202
+ $X2=3.885 $Y2=1.202
r168 61 63 18.1398 $w=3.72e-07 $l=1.4e-07 $layer=POLY_cond $X=3.72 $Y=1.202
+ $X2=3.86 $Y2=1.202
r169 61 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.72
+ $Y=1.16 $X2=3.72 $Y2=1.16
r170 59 61 42.7581 $w=3.72e-07 $l=3.3e-07 $layer=POLY_cond $X=3.39 $Y=1.202
+ $X2=3.72 $Y2=1.202
r171 58 59 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.365 $Y=1.202
+ $X2=3.39 $Y2=1.202
r172 57 58 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=2.92 $Y=1.202
+ $X2=3.365 $Y2=1.202
r173 56 57 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.895 $Y=1.202
+ $X2=2.92 $Y2=1.202
r174 55 62 64.8818 $w=1.98e-07 $l=1.17e-06 $layer=LI1_cond $X=2.55 $Y=1.175
+ $X2=3.72 $Y2=1.175
r175 54 56 44.7016 $w=3.72e-07 $l=3.45e-07 $layer=POLY_cond $X=2.55 $Y=1.202
+ $X2=2.895 $Y2=1.202
r176 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.55
+ $Y=1.16 $X2=2.55 $Y2=1.16
r177 52 54 12.957 $w=3.72e-07 $l=1e-07 $layer=POLY_cond $X=2.45 $Y=1.202
+ $X2=2.55 $Y2=1.202
r178 51 52 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.425 $Y=1.202
+ $X2=2.45 $Y2=1.202
r179 49 84 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=4.37 $Y=1.175
+ $X2=4.385 $Y2=1.175
r180 49 62 36.0455 $w=1.98e-07 $l=6.5e-07 $layer=LI1_cond $X=4.37 $Y=1.175
+ $X2=3.72 $Y2=1.175
r181 46 78 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.285 $Y=0.995
+ $X2=6.285 $Y2=1.202
r182 46 48 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.285 $Y=0.995
+ $X2=6.285 $Y2=0.56
r183 43 77 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.26 $Y=1.41
+ $X2=6.26 $Y2=1.202
r184 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.26 $Y=1.41
+ $X2=6.26 $Y2=1.985
r185 40 76 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.79 $Y=1.41
+ $X2=5.79 $Y2=1.202
r186 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.79 $Y=1.41
+ $X2=5.79 $Y2=1.985
r187 37 75 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.765 $Y=0.995
+ $X2=5.765 $Y2=1.202
r188 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.765 $Y=0.995
+ $X2=5.765 $Y2=0.56
r189 34 71 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.32 $Y=1.41
+ $X2=5.32 $Y2=1.202
r190 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.32 $Y=1.41
+ $X2=5.32 $Y2=1.985
r191 31 70 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.295 $Y=0.995
+ $X2=5.295 $Y2=1.202
r192 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.295 $Y=0.995
+ $X2=5.295 $Y2=0.56
r193 28 66 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.85 $Y=1.41
+ $X2=4.85 $Y2=1.202
r194 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.85 $Y=1.41
+ $X2=4.85 $Y2=1.985
r195 25 65 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.825 $Y=0.995
+ $X2=4.825 $Y2=1.202
r196 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.825 $Y=0.995
+ $X2=4.825 $Y2=0.56
r197 22 64 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.885 $Y=0.995
+ $X2=3.885 $Y2=1.202
r198 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.885 $Y=0.995
+ $X2=3.885 $Y2=0.56
r199 19 63 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.86 $Y=1.41
+ $X2=3.86 $Y2=1.202
r200 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.86 $Y=1.41
+ $X2=3.86 $Y2=1.985
r201 16 59 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.39 $Y=1.41
+ $X2=3.39 $Y2=1.202
r202 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.39 $Y=1.41
+ $X2=3.39 $Y2=1.985
r203 13 58 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.365 $Y=0.995
+ $X2=3.365 $Y2=1.202
r204 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.365 $Y=0.995
+ $X2=3.365 $Y2=0.56
r205 10 57 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.92 $Y=1.41
+ $X2=2.92 $Y2=1.202
r206 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.92 $Y=1.41
+ $X2=2.92 $Y2=1.985
r207 7 56 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.895 $Y=0.995
+ $X2=2.895 $Y2=1.202
r208 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.895 $Y=0.995
+ $X2=2.895 $Y2=0.56
r209 4 52 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.45 $Y=1.41
+ $X2=2.45 $Y2=1.202
r210 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.45 $Y=1.41
+ $X2=2.45 $Y2=1.985
r211 1 51 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.425 $Y=0.995
+ $X2=2.425 $Y2=1.202
r212 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.425 $Y=0.995
+ $X2=2.425 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_4%A_38_297# 1 2 3 4 5 6 7 22 24 25 27 28 30
+ 31 33 34 36 37 39 40 42 43 45 47 50 54 58 60 62 68 72 76 81 82 87 90 92 94 96
+ 98 99 100 101 107 118
c223 107 0 1.5003e-19 $X=6.81 $Y=1.53
r224 118 119 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=10.54 $Y=1.202
+ $X2=10.565 $Y2=1.202
r225 115 116 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=10.045 $Y=1.202
+ $X2=10.07 $Y2=1.202
r226 114 115 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=9.6 $Y=1.202
+ $X2=10.045 $Y2=1.202
r227 113 114 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=9.575 $Y=1.202
+ $X2=9.6 $Y2=1.202
r228 110 111 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=9.105 $Y=1.202
+ $X2=9.13 $Y2=1.202
r229 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.81 $Y=1.53
+ $X2=6.81 $Y2=1.53
r230 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.25 $Y=1.53
+ $X2=1.25 $Y2=1.53
r231 101 103 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.395 $Y=1.53
+ $X2=1.25 $Y2=1.53
r232 100 107 0.121883 $w=2.3e-07 $l=1.55e-07 $layer=MET1_cond $X=6.655 $Y=1.53
+ $X2=6.81 $Y2=1.53
r233 100 101 6.50989 $w=1.4e-07 $l=5.26e-06 $layer=MET1_cond $X=6.655 $Y=1.53
+ $X2=1.395 $Y2=1.53
r234 99 108 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=8.39 $Y=1.53
+ $X2=6.81 $Y2=1.53
r235 88 118 22.0269 $w=3.72e-07 $l=1.7e-07 $layer=POLY_cond $X=10.37 $Y=1.202
+ $X2=10.54 $Y2=1.202
r236 88 116 38.871 $w=3.72e-07 $l=3e-07 $layer=POLY_cond $X=10.37 $Y=1.202
+ $X2=10.07 $Y2=1.202
r237 87 88 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.37
+ $Y=1.16 $X2=10.37 $Y2=1.16
r238 85 113 48.5887 $w=3.72e-07 $l=3.75e-07 $layer=POLY_cond $X=9.2 $Y=1.202
+ $X2=9.575 $Y2=1.202
r239 85 111 9.06989 $w=3.72e-07 $l=7e-08 $layer=POLY_cond $X=9.2 $Y=1.202
+ $X2=9.13 $Y2=1.202
r240 84 87 64.8818 $w=1.98e-07 $l=1.17e-06 $layer=LI1_cond $X=9.2 $Y=1.175
+ $X2=10.37 $Y2=1.175
r241 84 85 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.2
+ $Y=1.16 $X2=9.2 $Y2=1.16
r242 82 84 35.4909 $w=1.98e-07 $l=6.4e-07 $layer=LI1_cond $X=8.56 $Y=1.175
+ $X2=9.2 $Y2=1.175
r243 81 99 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.475 $Y=1.445
+ $X2=8.39 $Y2=1.53
r244 80 82 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=8.475 $Y=1.275
+ $X2=8.56 $Y2=1.175
r245 80 81 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.475 $Y=1.275
+ $X2=8.475 $Y2=1.445
r246 77 96 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=3.28 $Y=1.895
+ $X2=3.155 $Y2=1.895
r247 76 98 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=3.97 $Y=1.895
+ $X2=4.095 $Y2=1.895
r248 76 77 36.1448 $w=2.18e-07 $l=6.9e-07 $layer=LI1_cond $X=3.97 $Y=1.895
+ $X2=3.28 $Y2=1.895
r249 73 94 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=2.34 $Y=1.895
+ $X2=2.215 $Y2=1.895
r250 72 96 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=3.03 $Y=1.895
+ $X2=3.155 $Y2=1.895
r251 72 73 36.1448 $w=2.18e-07 $l=6.9e-07 $layer=LI1_cond $X=3.03 $Y=1.895
+ $X2=2.34 $Y2=1.895
r252 69 92 1.80668 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=1.4 $Y=1.895
+ $X2=1.275 $Y2=1.895
r253 68 94 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=2.09 $Y=1.895
+ $X2=2.215 $Y2=1.895
r254 68 69 36.1448 $w=2.18e-07 $l=6.9e-07 $layer=LI1_cond $X=2.09 $Y=1.895
+ $X2=1.4 $Y2=1.895
r255 63 92 4.63873 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=1.275 $Y=1.785
+ $X2=1.275 $Y2=1.895
r256 63 65 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.275 $Y=1.785
+ $X2=1.275 $Y2=1.62
r257 62 104 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.275 $Y=1.615
+ $X2=1.275 $Y2=1.53
r258 62 65 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.275 $Y=1.615
+ $X2=1.275 $Y2=1.62
r259 61 90 3.51065 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.46 $Y=1.53
+ $X2=0.272 $Y2=1.53
r260 60 104 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.15 $Y=1.53
+ $X2=1.275 $Y2=1.53
r261 60 61 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.15 $Y=1.53
+ $X2=0.46 $Y2=1.53
r262 56 58 41.6652 $w=2.58e-07 $l=9.4e-07 $layer=LI1_cond $X=0.805 $Y=0.775
+ $X2=1.745 $Y2=0.775
r263 54 56 21.4975 $w=2.58e-07 $l=4.85e-07 $layer=LI1_cond $X=0.32 $Y=0.775
+ $X2=0.805 $Y2=0.775
r264 50 52 20.8976 $w=3.73e-07 $l=6.8e-07 $layer=LI1_cond $X=0.272 $Y=1.62
+ $X2=0.272 $Y2=2.3
r265 48 90 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.272 $Y=1.615
+ $X2=0.272 $Y2=1.53
r266 48 50 0.153659 $w=3.73e-07 $l=5e-09 $layer=LI1_cond $X=0.272 $Y=1.615
+ $X2=0.272 $Y2=1.62
r267 47 90 3.10218 $w=3.05e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.202 $Y=1.445
+ $X2=0.272 $Y2=1.53
r268 46 54 6.83913 $w=2.6e-07 $l=1.79555e-07 $layer=LI1_cond $X=0.202 $Y=0.905
+ $X2=0.32 $Y2=0.775
r269 46 47 26.4817 $w=2.33e-07 $l=5.4e-07 $layer=LI1_cond $X=0.202 $Y=0.905
+ $X2=0.202 $Y2=1.445
r270 43 119 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.565 $Y=0.995
+ $X2=10.565 $Y2=1.202
r271 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.565 $Y=0.995
+ $X2=10.565 $Y2=0.56
r272 40 118 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.54 $Y=1.41
+ $X2=10.54 $Y2=1.202
r273 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.54 $Y=1.41
+ $X2=10.54 $Y2=1.985
r274 37 116 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.07 $Y=1.41
+ $X2=10.07 $Y2=1.202
r275 37 39 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.07 $Y=1.41
+ $X2=10.07 $Y2=1.985
r276 34 115 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.045 $Y=0.995
+ $X2=10.045 $Y2=1.202
r277 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.045 $Y=0.995
+ $X2=10.045 $Y2=0.56
r278 31 114 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.6 $Y=1.41
+ $X2=9.6 $Y2=1.202
r279 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.6 $Y=1.41
+ $X2=9.6 $Y2=1.985
r280 28 113 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.575 $Y=0.995
+ $X2=9.575 $Y2=1.202
r281 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.575 $Y=0.995
+ $X2=9.575 $Y2=0.56
r282 25 111 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.13 $Y=1.41
+ $X2=9.13 $Y2=1.202
r283 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.13 $Y=1.41
+ $X2=9.13 $Y2=1.985
r284 22 110 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.105 $Y=0.995
+ $X2=9.105 $Y2=1.202
r285 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.105 $Y=0.995
+ $X2=9.105 $Y2=0.56
r286 7 98 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.95
+ $Y=1.485 $X2=4.095 $Y2=1.96
r287 6 96 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.01
+ $Y=1.485 $X2=3.155 $Y2=1.96
r288 5 94 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.07
+ $Y=1.485 $X2=2.215 $Y2=1.96
r289 4 92 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.13
+ $Y=1.485 $X2=1.275 $Y2=1.96
r290 4 65 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=1.485 $X2=1.275 $Y2=1.62
r291 3 52 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.19
+ $Y=1.485 $X2=0.335 $Y2=2.3
r292 3 50 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.19
+ $Y=1.485 $X2=0.335 $Y2=1.62
r293 2 58 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.235 $X2=1.745 $Y2=0.73
r294 1 56 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=0.62
+ $Y=0.235 $X2=0.805 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_4%VPWR 1 2 3 4 5 6 7 8 29 33 37 41 45 49 53
+ 57 60 61 63 64 66 67 69 70 72 73 75 76 78 79 80 111 112 115
r159 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r160 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r161 109 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.81 $Y2=2.72
r162 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r163 106 109 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r164 105 106 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r165 103 106 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=8.97 $Y2=2.72
r166 102 105 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=6.21 $Y=2.72
+ $X2=8.97 $Y2=2.72
r167 102 103 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r168 100 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r169 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r170 97 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r171 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r172 94 97 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r173 93 96 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r174 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r175 91 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r176 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r177 88 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r178 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r179 85 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r180 85 116 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r181 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r182 82 115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.93 $Y=2.72
+ $X2=0.805 $Y2=2.72
r183 82 84 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.93 $Y=2.72
+ $X2=1.61 $Y2=2.72
r184 80 116 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r185 78 108 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=10.18 $Y=2.72
+ $X2=9.89 $Y2=2.72
r186 78 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.18 $Y=2.72
+ $X2=10.305 $Y2=2.72
r187 77 111 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=10.43 $Y=2.72
+ $X2=10.81 $Y2=2.72
r188 77 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.43 $Y=2.72
+ $X2=10.305 $Y2=2.72
r189 75 105 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.24 $Y=2.72
+ $X2=8.97 $Y2=2.72
r190 75 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.24 $Y=2.72
+ $X2=9.365 $Y2=2.72
r191 74 108 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=9.49 $Y=2.72
+ $X2=9.89 $Y2=2.72
r192 74 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.49 $Y=2.72
+ $X2=9.365 $Y2=2.72
r193 72 99 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.9 $Y=2.72 $X2=5.75
+ $Y2=2.72
r194 72 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.9 $Y=2.72
+ $X2=6.025 $Y2=2.72
r195 71 102 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=6.15 $Y=2.72
+ $X2=6.21 $Y2=2.72
r196 71 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.15 $Y=2.72
+ $X2=6.025 $Y2=2.72
r197 69 96 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.96 $Y=2.72
+ $X2=4.83 $Y2=2.72
r198 69 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.96 $Y=2.72
+ $X2=5.085 $Y2=2.72
r199 68 99 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=5.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r200 68 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.21 $Y=2.72
+ $X2=5.085 $Y2=2.72
r201 66 90 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=3.5 $Y=2.72 $X2=3.45
+ $Y2=2.72
r202 66 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.5 $Y=2.72
+ $X2=3.625 $Y2=2.72
r203 65 93 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.75 $Y=2.72
+ $X2=3.91 $Y2=2.72
r204 65 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.75 $Y=2.72
+ $X2=3.625 $Y2=2.72
r205 63 87 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.56 $Y=2.72 $X2=2.53
+ $Y2=2.72
r206 63 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.56 $Y=2.72
+ $X2=2.685 $Y2=2.72
r207 62 90 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.81 $Y=2.72
+ $X2=3.45 $Y2=2.72
r208 62 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.81 $Y=2.72
+ $X2=2.685 $Y2=2.72
r209 60 84 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.62 $Y=2.72
+ $X2=1.61 $Y2=2.72
r210 60 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.62 $Y=2.72
+ $X2=1.745 $Y2=2.72
r211 59 87 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.87 $Y=2.72
+ $X2=2.53 $Y2=2.72
r212 59 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.87 $Y=2.72
+ $X2=1.745 $Y2=2.72
r213 55 79 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.305 $Y=2.635
+ $X2=10.305 $Y2=2.72
r214 55 57 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=10.305 $Y=2.635
+ $X2=10.305 $Y2=2
r215 51 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.365 $Y=2.635
+ $X2=9.365 $Y2=2.72
r216 51 53 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=9.365 $Y=2.635
+ $X2=9.365 $Y2=2
r217 47 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.025 $Y=2.635
+ $X2=6.025 $Y2=2.72
r218 47 49 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=6.025 $Y=2.635
+ $X2=6.025 $Y2=2.34
r219 43 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.085 $Y=2.635
+ $X2=5.085 $Y2=2.72
r220 43 45 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=5.085 $Y=2.635
+ $X2=5.085 $Y2=2.34
r221 39 67 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=2.635
+ $X2=3.625 $Y2=2.72
r222 39 41 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.625 $Y=2.635
+ $X2=3.625 $Y2=2.34
r223 35 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.685 $Y=2.635
+ $X2=2.685 $Y2=2.72
r224 35 37 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.685 $Y=2.635
+ $X2=2.685 $Y2=2.34
r225 31 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.745 $Y=2.635
+ $X2=1.745 $Y2=2.72
r226 31 33 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.745 $Y=2.635
+ $X2=1.745 $Y2=2.34
r227 27 115 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=2.635
+ $X2=0.805 $Y2=2.72
r228 27 29 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.805 $Y=2.635
+ $X2=0.805 $Y2=2
r229 8 57 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=10.16
+ $Y=1.485 $X2=10.305 $Y2=2
r230 7 53 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=9.22
+ $Y=1.485 $X2=9.365 $Y2=2
r231 6 49 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.88
+ $Y=1.485 $X2=6.025 $Y2=2.34
r232 5 45 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.94
+ $Y=1.485 $X2=5.085 $Y2=2.34
r233 4 41 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.48
+ $Y=1.485 $X2=3.625 $Y2=2.34
r234 3 37 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.54
+ $Y=1.485 $X2=2.685 $Y2=2.34
r235 2 33 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.6
+ $Y=1.485 $X2=1.745 $Y2=2.34
r236 1 29 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.66
+ $Y=1.485 $X2=0.805 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_4%A_898_297# 1 2 3 4 5 18 22 24 25 30 33 35
r64 28 30 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=7.435 $Y=2.34
+ $X2=8.375 $Y2=2.34
r65 26 39 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=6.58 $Y=2.34
+ $X2=6.475 $Y2=2.34
r66 26 28 39.4136 $w=2.48e-07 $l=8.55e-07 $layer=LI1_cond $X=6.58 $Y=2.34
+ $X2=7.435 $Y2=2.34
r67 25 39 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=6.475 $Y=2.215
+ $X2=6.475 $Y2=2.34
r68 24 37 3.48996 $w=2.1e-07 $l=1.1e-07 $layer=LI1_cond $X=6.475 $Y=2.005
+ $X2=6.475 $Y2=1.895
r69 24 25 11.0909 $w=2.08e-07 $l=2.1e-07 $layer=LI1_cond $X=6.475 $Y=2.005
+ $X2=6.475 $Y2=2.215
r70 23 35 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=5.68 $Y=1.895
+ $X2=5.555 $Y2=1.895
r71 22 37 3.33133 $w=2.2e-07 $l=1.05e-07 $layer=LI1_cond $X=6.37 $Y=1.895
+ $X2=6.475 $Y2=1.895
r72 22 23 36.1448 $w=2.18e-07 $l=6.9e-07 $layer=LI1_cond $X=6.37 $Y=1.895
+ $X2=5.68 $Y2=1.895
r73 19 33 4.18571 $w=2.2e-07 $l=1.58e-07 $layer=LI1_cond $X=4.74 $Y=1.895
+ $X2=4.582 $Y2=1.895
r74 18 35 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=5.43 $Y=1.895
+ $X2=5.555 $Y2=1.895
r75 18 19 36.1448 $w=2.18e-07 $l=6.9e-07 $layer=LI1_cond $X=5.43 $Y=1.895
+ $X2=4.74 $Y2=1.895
r76 5 30 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=8.23
+ $Y=1.485 $X2=8.375 $Y2=2.3
r77 4 28 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=7.29
+ $Y=1.485 $X2=7.435 $Y2=2.3
r78 3 39 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=6.35
+ $Y=1.485 $X2=6.495 $Y2=2.3
r79 3 37 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=6.35
+ $Y=1.485 $X2=6.495 $Y2=1.96
r80 2 35 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.41
+ $Y=1.485 $X2=5.555 $Y2=1.96
r81 1 33 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=4.49
+ $Y=1.485 $X2=4.615 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_4%Y 1 2 3 4 5 6 7 22 30 32 34 42 44 48 50 56
+ 59 61 64
r84 61 64 0.735602 $w=2.33e-07 $l=1.5e-08 $layer=LI1_cond $X=10.822 $Y=1.19
+ $X2=10.822 $Y2=1.175
r85 60 64 13.2408 $w=2.33e-07 $l=2.7e-07 $layer=LI1_cond $X=10.822 $Y=0.905
+ $X2=10.822 $Y2=1.175
r86 57 61 12.5052 $w=2.33e-07 $l=2.55e-07 $layer=LI1_cond $X=10.822 $Y=1.445
+ $X2=10.822 $Y2=1.19
r87 57 59 4.1757 $w=2.82e-07 $l=1.31415e-07 $layer=LI1_cond $X=10.822 $Y=1.445
+ $X2=10.775 $Y2=1.555
r88 53 54 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=8.895 $Y=1.66
+ $X2=8.895 $Y2=1.915
r89 50 53 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=8.895 $Y=1.555
+ $X2=8.895 $Y2=1.66
r90 46 59 4.1757 $w=2.82e-07 $l=1.1e-07 $layer=LI1_cond $X=10.775 $Y=1.665
+ $X2=10.775 $Y2=1.555
r91 46 48 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=10.775 $Y=1.665
+ $X2=10.775 $Y2=2.34
r92 45 56 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=9.96 $Y=1.555
+ $X2=9.835 $Y2=1.555
r93 44 59 2.25663 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=10.61 $Y=1.555
+ $X2=10.775 $Y2=1.555
r94 44 45 34.0495 $w=2.18e-07 $l=6.5e-07 $layer=LI1_cond $X=10.61 $Y=1.555
+ $X2=9.96 $Y2=1.555
r95 40 56 0.886536 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=9.835 $Y=1.665
+ $X2=9.835 $Y2=1.555
r96 40 42 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=9.835 $Y=1.665
+ $X2=9.835 $Y2=2.3
r97 36 39 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=9.365 $Y=0.78
+ $X2=10.305 $Y2=0.78
r98 34 60 6.82498 $w=2.5e-07 $l=1.73925e-07 $layer=LI1_cond $X=10.705 $Y=0.78
+ $X2=10.822 $Y2=0.905
r99 34 39 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=10.705 $Y=0.78
+ $X2=10.305 $Y2=0.78
r100 33 50 3.11056 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=9.06 $Y=1.555
+ $X2=8.895 $Y2=1.555
r101 32 56 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=9.71 $Y=1.555
+ $X2=9.835 $Y2=1.555
r102 32 33 34.0495 $w=2.18e-07 $l=6.5e-07 $layer=LI1_cond $X=9.71 $Y=1.555
+ $X2=9.06 $Y2=1.555
r103 28 54 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=8.895 $Y=2.045
+ $X2=8.895 $Y2=1.915
r104 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.895 $Y=2.045
+ $X2=8.895 $Y2=2.34
r105 24 27 41.6652 $w=2.58e-07 $l=9.4e-07 $layer=LI1_cond $X=6.965 $Y=1.915
+ $X2=7.905 $Y2=1.915
r106 22 54 2.13598 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=8.73 $Y=1.915
+ $X2=8.895 $Y2=1.915
r107 22 27 36.5679 $w=2.58e-07 $l=8.25e-07 $layer=LI1_cond $X=8.73 $Y=1.915
+ $X2=7.905 $Y2=1.915
r108 7 59 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=10.63
+ $Y=1.485 $X2=10.775 $Y2=1.66
r109 7 48 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.63
+ $Y=1.485 $X2=10.775 $Y2=2.34
r110 6 56 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.69
+ $Y=1.485 $X2=9.835 $Y2=1.62
r111 6 42 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=9.69
+ $Y=1.485 $X2=9.835 $Y2=2.3
r112 5 53 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=8.77
+ $Y=1.485 $X2=8.895 $Y2=1.66
r113 5 30 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=8.77
+ $Y=1.485 $X2=8.895 $Y2=2.34
r114 4 27 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=1.485 $X2=7.905 $Y2=1.96
r115 3 24 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=6.82
+ $Y=1.485 $X2=6.965 $Y2=1.96
r116 2 39 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=10.12
+ $Y=0.235 $X2=10.305 $Y2=0.74
r117 1 36 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=9.18
+ $Y=0.235 $X2=9.365 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_4%A_38_47# 1 2 3 4 5 16 22 23 24 28 30 34 40
c72 23 0 1.98558e-19 $X=2.255 $Y=0.725
r73 32 34 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.07 $Y=0.725
+ $X2=4.07 $Y2=0.39
r74 31 40 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.32 $Y=0.815
+ $X2=3.13 $Y2=0.815
r75 30 32 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=3.88 $Y=0.815
+ $X2=4.07 $Y2=0.725
r76 30 31 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.88 $Y=0.815
+ $X2=3.32 $Y2=0.815
r77 26 40 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=3.13 $Y=0.725 $X2=3.13
+ $Y2=0.815
r78 26 28 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.13 $Y=0.725
+ $X2=3.13 $Y2=0.39
r79 25 39 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=2.38 $Y=0.815
+ $X2=2.255 $Y2=0.815
r80 24 40 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.94 $Y=0.815
+ $X2=3.13 $Y2=0.815
r81 24 25 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=2.94 $Y=0.815
+ $X2=2.38 $Y2=0.815
r82 23 39 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=2.255 $Y=0.725
+ $X2=2.255 $Y2=0.815
r83 22 37 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=2.255 $Y=0.475
+ $X2=2.255 $Y2=0.365
r84 22 23 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=2.255 $Y=0.475
+ $X2=2.255 $Y2=0.725
r85 18 21 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=0.335 $Y=0.365
+ $X2=1.275 $Y2=0.365
r86 16 37 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=2.13 $Y=0.365
+ $X2=2.255 $Y2=0.365
r87 16 21 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=2.13 $Y=0.365
+ $X2=1.275 $Y2=0.365
r88 5 34 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.96
+ $Y=0.235 $X2=4.095 $Y2=0.39
r89 4 28 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=2.97
+ $Y=0.235 $X2=3.155 $Y2=0.39
r90 3 39 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.08
+ $Y=0.235 $X2=2.215 $Y2=0.73
r91 3 37 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.08
+ $Y=0.235 $X2=2.215 $Y2=0.39
r92 2 21 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.235 $X2=1.275 $Y2=0.39
r93 1 18 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=0.19
+ $Y=0.235 $X2=0.335 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_4%VGND 1 2 3 4 5 6 7 24 28 32 36 40 44 48 51
+ 52 54 55 57 58 60 61 63 64 66 67 69 70 71 102 103
r159 102 103 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r160 100 103 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=10.81 $Y2=0
r161 99 102 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=8.51 $Y=0
+ $X2=10.81 $Y2=0
r162 99 100 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r163 97 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.51 $Y2=0
r164 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r165 94 97 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=8.05
+ $Y2=0
r166 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r167 91 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r168 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r169 88 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r170 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r171 85 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r172 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r173 82 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r174 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r175 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r176 78 79 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r177 74 78 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r178 71 79 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r179 71 74 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r180 69 96 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=8.29 $Y=0 $X2=8.05
+ $Y2=0
r181 69 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.29 $Y=0 $X2=8.375
+ $Y2=0
r182 68 99 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=8.46 $Y=0 $X2=8.51
+ $Y2=0
r183 68 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.46 $Y=0 $X2=8.375
+ $Y2=0
r184 66 93 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=7.35 $Y=0 $X2=7.13
+ $Y2=0
r185 66 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.35 $Y=0 $X2=7.435
+ $Y2=0
r186 65 96 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.52 $Y=0 $X2=8.05
+ $Y2=0
r187 65 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.52 $Y=0 $X2=7.435
+ $Y2=0
r188 63 90 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=6.41 $Y=0 $X2=6.21
+ $Y2=0
r189 63 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.41 $Y=0 $X2=6.495
+ $Y2=0
r190 62 93 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=6.58 $Y=0 $X2=7.13
+ $Y2=0
r191 62 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.58 $Y=0 $X2=6.495
+ $Y2=0
r192 60 87 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.47 $Y=0 $X2=5.29
+ $Y2=0
r193 60 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.47 $Y=0 $X2=5.555
+ $Y2=0
r194 59 90 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.64 $Y=0 $X2=6.21
+ $Y2=0
r195 59 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.64 $Y=0 $X2=5.555
+ $Y2=0
r196 57 84 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=4.43 $Y=0 $X2=4.37
+ $Y2=0
r197 57 58 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.43 $Y=0 $X2=4.565
+ $Y2=0
r198 56 87 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.7 $Y=0 $X2=5.29
+ $Y2=0
r199 56 58 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.7 $Y=0 $X2=4.565
+ $Y2=0
r200 54 81 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.54 $Y=0 $X2=3.45
+ $Y2=0
r201 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=0 $X2=3.625
+ $Y2=0
r202 53 84 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=3.71 $Y=0 $X2=4.37
+ $Y2=0
r203 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=0 $X2=3.625
+ $Y2=0
r204 51 78 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.6 $Y=0 $X2=2.53
+ $Y2=0
r205 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.6 $Y=0 $X2=2.685
+ $Y2=0
r206 50 81 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.77 $Y=0 $X2=3.45
+ $Y2=0
r207 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.77 $Y=0 $X2=2.685
+ $Y2=0
r208 46 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.375 $Y=0.085
+ $X2=8.375 $Y2=0
r209 46 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.375 $Y=0.085
+ $X2=8.375 $Y2=0.39
r210 42 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.435 $Y=0.085
+ $X2=7.435 $Y2=0
r211 42 44 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.435 $Y=0.085
+ $X2=7.435 $Y2=0.39
r212 38 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.495 $Y=0.085
+ $X2=6.495 $Y2=0
r213 38 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.495 $Y=0.085
+ $X2=6.495 $Y2=0.39
r214 34 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.555 $Y=0.085
+ $X2=5.555 $Y2=0
r215 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.555 $Y=0.085
+ $X2=5.555 $Y2=0.39
r216 30 58 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=0.085
+ $X2=4.565 $Y2=0
r217 30 32 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.565 $Y=0.085
+ $X2=4.565 $Y2=0.39
r218 26 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=0.085
+ $X2=3.625 $Y2=0
r219 26 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.625 $Y=0.085
+ $X2=3.625 $Y2=0.39
r220 22 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.685 $Y=0.085
+ $X2=2.685 $Y2=0
r221 22 24 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.685 $Y=0.085
+ $X2=2.685 $Y2=0.39
r222 7 48 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=8.24
+ $Y=0.235 $X2=8.375 $Y2=0.39
r223 6 44 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=7.25
+ $Y=0.235 $X2=7.435 $Y2=0.39
r224 5 40 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.36
+ $Y=0.235 $X2=6.495 $Y2=0.39
r225 4 36 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=5.37
+ $Y=0.235 $X2=5.555 $Y2=0.39
r226 3 32 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=4.49
+ $Y=0.235 $X2=4.615 $Y2=0.39
r227 2 28 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=3.44
+ $Y=0.235 $X2=3.625 $Y2=0.39
r228 1 24 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.5
+ $Y=0.235 $X2=2.685 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_4%A_980_47# 1 2 3 4 5 6 7 24 26 27 30 32 36
+ 38 42 44 46 49 54 56 57 58
r116 52 54 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=9.835 $Y=0.39
+ $X2=10.775 $Y2=0.39
r117 50 60 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.98 $Y=0.39
+ $X2=8.855 $Y2=0.39
r118 50 52 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=8.98 $Y=0.39
+ $X2=9.835 $Y2=0.39
r119 47 49 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=8.855 $Y=0.735
+ $X2=8.855 $Y2=0.73
r120 46 60 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.855 $Y=0.475
+ $X2=8.855 $Y2=0.39
r121 46 49 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=8.855 $Y=0.475
+ $X2=8.855 $Y2=0.73
r122 45 58 9.30075 $w=1.75e-07 $l=2.42487e-07 $layer=LI1_cond $X=8.17 $Y=0.82
+ $X2=7.93 $Y2=0.815
r123 44 47 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.73 $Y=0.82
+ $X2=8.855 $Y2=0.735
r124 44 45 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.73 $Y=0.82
+ $X2=8.17 $Y2=0.82
r125 40 58 1.23463 $w=3.8e-07 $l=1.1225e-07 $layer=LI1_cond $X=7.88 $Y=0.725
+ $X2=7.93 $Y2=0.815
r126 40 42 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.88 $Y=0.725
+ $X2=7.88 $Y2=0.39
r127 39 57 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=7.13 $Y=0.815
+ $X2=6.94 $Y2=0.815
r128 38 58 9.30075 $w=1.75e-07 $l=2.4e-07 $layer=LI1_cond $X=7.69 $Y=0.815
+ $X2=7.93 $Y2=0.815
r129 38 39 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=7.69 $Y=0.815
+ $X2=7.13 $Y2=0.815
r130 34 57 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=6.94 $Y=0.725 $X2=6.94
+ $Y2=0.815
r131 34 36 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.94 $Y=0.725
+ $X2=6.94 $Y2=0.39
r132 33 56 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.19 $Y=0.815 $X2=6
+ $Y2=0.815
r133 32 57 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.75 $Y=0.815
+ $X2=6.94 $Y2=0.815
r134 32 33 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=6.75 $Y=0.815
+ $X2=6.19 $Y2=0.815
r135 28 56 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=6 $Y=0.725 $X2=6
+ $Y2=0.815
r136 28 30 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6 $Y=0.725 $X2=6
+ $Y2=0.39
r137 26 56 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.81 $Y=0.815 $X2=6
+ $Y2=0.815
r138 26 27 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=5.81 $Y=0.815
+ $X2=5.25 $Y2=0.815
r139 22 27 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=5.06 $Y=0.725
+ $X2=5.25 $Y2=0.815
r140 22 24 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.06 $Y=0.725
+ $X2=5.06 $Y2=0.39
r141 7 54 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=10.64
+ $Y=0.235 $X2=10.775 $Y2=0.39
r142 6 52 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=9.65
+ $Y=0.235 $X2=9.835 $Y2=0.39
r143 5 60 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=8.77
+ $Y=0.235 $X2=8.895 $Y2=0.39
r144 5 49 182 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_NDIFF $count=1 $X=8.77
+ $Y=0.235 $X2=8.895 $Y2=0.73
r145 4 42 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=7.72
+ $Y=0.235 $X2=7.905 $Y2=0.39
r146 3 36 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=6.78
+ $Y=0.235 $X2=6.965 $Y2=0.39
r147 2 30 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=5.84
+ $Y=0.235 $X2=6.025 $Y2=0.39
r148 1 24 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.9
+ $Y=0.235 $X2=5.085 $Y2=0.39
.ends

