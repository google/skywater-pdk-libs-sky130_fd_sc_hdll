* File: sky130_fd_sc_hdll__a21o_6.pxi.spice
* Created: Wed Sep  2 08:17:26 2020
* 
x_PM_SKY130_FD_SC_HDLL__A21O_6%A2 N_A2_c_100_n N_A2_M1010_g N_A2_c_101_n
+ N_A2_M1000_g N_A2_c_102_n N_A2_M1012_g N_A2_c_103_n N_A2_M1015_g N_A2_c_109_n
+ N_A2_c_110_n N_A2_c_151_p N_A2_c_104_n N_A2_c_105_n N_A2_c_106_n A2
+ PM_SKY130_FD_SC_HDLL__A21O_6%A2
x_PM_SKY130_FD_SC_HDLL__A21O_6%A1 N_A1_c_192_n N_A1_M1002_g N_A1_c_188_n
+ N_A1_M1007_g N_A1_c_189_n N_A1_M1003_g N_A1_c_193_n N_A1_M1020_g A1
+ N_A1_c_190_n N_A1_c_191_n PM_SKY130_FD_SC_HDLL__A21O_6%A1
x_PM_SKY130_FD_SC_HDLL__A21O_6%B1 N_B1_c_244_n N_B1_M1008_g N_B1_c_240_n
+ N_B1_M1014_g N_B1_c_241_n N_B1_M1019_g N_B1_c_245_n N_B1_M1011_g B1
+ N_B1_c_243_n PM_SKY130_FD_SC_HDLL__A21O_6%B1
x_PM_SKY130_FD_SC_HDLL__A21O_6%A_213_47# N_A_213_47#_M1007_d N_A_213_47#_M1014_d
+ N_A_213_47#_M1008_s N_A_213_47#_c_305_n N_A_213_47#_M1004_g
+ N_A_213_47#_c_294_n N_A_213_47#_M1001_g N_A_213_47#_c_295_n
+ N_A_213_47#_M1005_g N_A_213_47#_c_306_n N_A_213_47#_M1006_g
+ N_A_213_47#_c_307_n N_A_213_47#_M1013_g N_A_213_47#_c_296_n
+ N_A_213_47#_M1009_g N_A_213_47#_c_297_n N_A_213_47#_M1016_g
+ N_A_213_47#_c_308_n N_A_213_47#_M1018_g N_A_213_47#_c_309_n
+ N_A_213_47#_M1021_g N_A_213_47#_c_298_n N_A_213_47#_M1017_g
+ N_A_213_47#_c_299_n N_A_213_47#_M1022_g N_A_213_47#_c_310_n
+ N_A_213_47#_M1023_g N_A_213_47#_c_313_n N_A_213_47#_c_315_n
+ N_A_213_47#_c_300_n N_A_213_47#_c_320_n N_A_213_47#_c_301_n
+ N_A_213_47#_c_342_n N_A_213_47#_c_302_n N_A_213_47#_c_303_n
+ N_A_213_47#_c_391_p N_A_213_47#_c_349_n N_A_213_47#_c_350_n
+ N_A_213_47#_c_304_n PM_SKY130_FD_SC_HDLL__A21O_6%A_213_47#
x_PM_SKY130_FD_SC_HDLL__A21O_6%A_27_297# N_A_27_297#_M1010_s N_A_27_297#_M1002_d
+ N_A_27_297#_M1015_s N_A_27_297#_M1011_d N_A_27_297#_c_474_n
+ N_A_27_297#_c_475_n N_A_27_297#_c_485_n N_A_27_297#_c_489_n
+ N_A_27_297#_c_492_n N_A_27_297#_c_476_n N_A_27_297#_c_477_n
+ N_A_27_297#_c_494_n N_A_27_297#_c_478_n N_A_27_297#_c_479_n
+ N_A_27_297#_c_497_n N_A_27_297#_c_500_n PM_SKY130_FD_SC_HDLL__A21O_6%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A21O_6%VPWR N_VPWR_M1010_d N_VPWR_M1020_s N_VPWR_M1004_s
+ N_VPWR_M1006_s N_VPWR_M1018_s N_VPWR_M1023_s N_VPWR_c_546_n N_VPWR_c_547_n
+ N_VPWR_c_548_n N_VPWR_c_549_n N_VPWR_c_550_n N_VPWR_c_551_n N_VPWR_c_552_n
+ N_VPWR_c_553_n N_VPWR_c_554_n N_VPWR_c_555_n N_VPWR_c_556_n N_VPWR_c_557_n
+ N_VPWR_c_558_n N_VPWR_c_559_n N_VPWR_c_560_n VPWR N_VPWR_c_561_n
+ N_VPWR_c_562_n N_VPWR_c_545_n N_VPWR_c_564_n N_VPWR_c_565_n
+ PM_SKY130_FD_SC_HDLL__A21O_6%VPWR
x_PM_SKY130_FD_SC_HDLL__A21O_6%X N_X_M1001_d N_X_M1009_d N_X_M1017_d N_X_M1004_d
+ N_X_M1013_d N_X_M1021_d N_X_c_660_n N_X_c_714_n N_X_c_654_n N_X_c_655_n
+ N_X_c_670_n N_X_c_674_n N_X_c_678_n N_X_c_718_n N_X_c_656_n N_X_c_685_n
+ N_X_c_688_n N_X_c_657_n N_X_c_723_n N_X_c_694_n N_X_c_658_n N_X_c_700_n X
+ PM_SKY130_FD_SC_HDLL__A21O_6%X
x_PM_SKY130_FD_SC_HDLL__A21O_6%VGND N_VGND_M1000_s N_VGND_M1012_s N_VGND_M1019_s
+ N_VGND_M1005_s N_VGND_M1016_s N_VGND_M1022_s N_VGND_c_746_n N_VGND_c_747_n
+ N_VGND_c_748_n N_VGND_c_749_n N_VGND_c_750_n N_VGND_c_751_n N_VGND_c_752_n
+ N_VGND_c_753_n N_VGND_c_754_n N_VGND_c_755_n N_VGND_c_756_n N_VGND_c_757_n
+ VGND N_VGND_c_758_n N_VGND_c_759_n N_VGND_c_760_n N_VGND_c_761_n
+ N_VGND_c_762_n N_VGND_c_763_n PM_SKY130_FD_SC_HDLL__A21O_6%VGND
cc_1 VNB N_A2_c_100_n 0.0293869f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_A2_c_101_n 0.0211848f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.995
cc_3 VNB N_A2_c_102_n 0.017665f $X=-0.19 $Y=-0.24 $X2=1.82 $Y2=0.995
cc_4 VNB N_A2_c_103_n 0.0197856f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_5 VNB N_A2_c_104_n 2.55318e-19 $X=-0.19 $Y=-0.24 $X2=1.79 $Y2=1.46
cc_6 VNB N_A2_c_105_n 0.0199748f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.172
cc_7 VNB N_A2_c_106_n 0.00458328f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_8 VNB N_A1_c_188_n 0.0161331f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.995
cc_9 VNB N_A1_c_189_n 0.0161021f $X=-0.19 $Y=-0.24 $X2=1.82 $Y2=0.995
cc_10 VNB N_A1_c_190_n 0.00291039f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.172
cc_11 VNB N_A1_c_191_n 0.035465f $X=-0.19 $Y=-0.24 $X2=1.79 $Y2=1.172
cc_12 VNB N_B1_c_240_n 0.0170767f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.995
cc_13 VNB N_B1_c_241_n 0.0201851f $X=-0.19 $Y=-0.24 $X2=1.82 $Y2=0.995
cc_14 VNB B1 0.00256212f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.29
cc_15 VNB N_B1_c_243_n 0.0540894f $X=-0.19 $Y=-0.24 $X2=1.79 $Y2=1.46
cc_16 VNB N_A_213_47#_c_294_n 0.0191654f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.29
cc_17 VNB N_A_213_47#_c_295_n 0.0169283f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.545
cc_18 VNB N_A_213_47#_c_296_n 0.0169331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_213_47#_c_297_n 0.0169084f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_20 VNB N_A_213_47#_c_298_n 0.0159577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_213_47#_c_299_n 0.0214437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_213_47#_c_300_n 0.00115748f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_213_47#_c_301_n 0.00103672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_213_47#_c_302_n 0.00339889f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_213_47#_c_303_n 0.00399351f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_213_47#_c_304_n 0.131914f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_545_n 0.288713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB X 0.00235332f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_746_n 0.0138449f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.172
cc_30 VNB N_VGND_c_747_n 0.0297009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_748_n 0.00501005f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_749_n 0.00413904f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_33 VNB N_VGND_c_750_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.172
cc_34 VNB N_VGND_c_751_n 0.0329125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_752_n 0.0172699f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_753_n 0.00515784f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_754_n 0.0165909f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_755_n 0.00515784f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_756_n 0.0172687f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_757_n 0.00480536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_758_n 0.0384028f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_759_n 0.0137583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_760_n 0.347996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_761_n 0.00631346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_762_n 0.0159607f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_763_n 0.0229593f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VPB N_A2_c_100_n 0.0332672f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_48 VPB N_A2_c_103_n 0.0243889f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_49 VPB N_A2_c_109_n 0.00148131f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.46
cc_50 VPB N_A2_c_110_n 0.0102624f $X=-0.19 $Y=1.305 $X2=1.705 $Y2=1.545
cc_51 VPB N_A2_c_104_n 0.00148131f $X=-0.19 $Y=1.305 $X2=1.79 $Y2=1.46
cc_52 VPB N_A1_c_192_n 0.016105f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_53 VPB N_A1_c_193_n 0.016105f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_54 VPB N_A1_c_191_n 0.0195118f $X=-0.19 $Y=1.305 $X2=1.79 $Y2=1.172
cc_55 VPB N_B1_c_244_n 0.0161061f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_56 VPB N_B1_c_245_n 0.0195953f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_57 VPB B1 0.00260515f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.29
cc_58 VPB N_B1_c_243_n 0.0295495f $X=-0.19 $Y=1.305 $X2=1.79 $Y2=1.46
cc_59 VPB N_A_213_47#_c_305_n 0.0197254f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_60 VPB N_A_213_47#_c_306_n 0.0157197f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.172
cc_61 VPB N_A_213_47#_c_307_n 0.0157197f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.172
cc_62 VPB N_A_213_47#_c_308_n 0.0156966f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_63 VPB N_A_213_47#_c_309_n 0.0155598f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_213_47#_c_310_n 0.0194579f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_213_47#_c_301_n 9.30672e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_213_47#_c_304_n 0.0772866f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_27_297#_c_474_n 0.0153465f $X=-0.19 $Y=1.305 $X2=1.705 $Y2=1.545
cc_68 VPB N_A_27_297#_c_475_n 0.0194072f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.172
cc_69 VPB N_A_27_297#_c_476_n 0.00407295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_27_297#_c_477_n 0.0019327f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.172
cc_71 VPB N_A_27_297#_c_478_n 0.00645964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_297#_c_479_n 0.00717518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_546_n 0.00466368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_547_n 0.0167297f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_75 VPB N_VPWR_c_548_n 0.0046582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_549_n 0.00462153f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_77 VPB N_VPWR_c_550_n 3.40287e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_551_n 3.37329e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_552_n 0.0495624f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_553_n 0.0404498f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_554_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_555_n 0.0167344f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_556_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_557_n 0.0147329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_558_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_559_n 0.0150512f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_560_n 0.00519718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_561_n 0.0172595f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_562_n 0.011849f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_545_n 0.0626784f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_564_n 0.00516022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_565_n 0.00515985f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_X_c_654_n 0.00180924f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_94 VPB N_X_c_655_n 0.00215492f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_95 VPB N_X_c_656_n 0.00213184f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_X_c_657_n 0.00211041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_X_c_658_n 0.00162501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB X 0.0014431f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 N_A2_c_100_n N_A1_c_192_n 0.0364735f $X=0.495 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_100 N_A2_c_109_n N_A1_c_192_n 0.00101315f $X=0.61 $Y=1.46 $X2=-0.19 $Y2=-0.24
cc_101 N_A2_c_110_n N_A1_c_192_n 0.0118662f $X=1.705 $Y=1.545 $X2=-0.19
+ $Y2=-0.24
cc_102 N_A2_c_101_n N_A1_c_188_n 0.0418602f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A2_c_102_n N_A1_c_189_n 0.0440841f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A2_c_103_n N_A1_c_193_n 0.0364735f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A2_c_110_n N_A1_c_193_n 0.0118662f $X=1.705 $Y=1.545 $X2=0 $Y2=0
cc_106 N_A2_c_104_n N_A1_c_193_n 0.00101315f $X=1.79 $Y=1.46 $X2=0 $Y2=0
cc_107 N_A2_c_100_n N_A1_c_190_n 2.66334e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A2_c_103_n N_A1_c_190_n 2.67076e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A2_c_110_n N_A1_c_190_n 0.0477309f $X=1.705 $Y=1.545 $X2=0 $Y2=0
cc_110 N_A2_c_105_n N_A1_c_190_n 0.0205474f $X=0.525 $Y=1.172 $X2=0 $Y2=0
cc_111 N_A2_c_106_n N_A1_c_190_n 0.0196709f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A2_c_100_n N_A1_c_191_n 0.0260406f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A2_c_103_n N_A1_c_191_n 0.0259586f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A2_c_109_n N_A1_c_191_n 0.0024835f $X=0.61 $Y=1.46 $X2=0 $Y2=0
cc_115 N_A2_c_110_n N_A1_c_191_n 0.0081936f $X=1.705 $Y=1.545 $X2=0 $Y2=0
cc_116 N_A2_c_104_n N_A1_c_191_n 0.00250084f $X=1.79 $Y=1.46 $X2=0 $Y2=0
cc_117 N_A2_c_105_n N_A1_c_191_n 8.47697e-19 $X=0.525 $Y=1.172 $X2=0 $Y2=0
cc_118 N_A2_c_106_n N_A1_c_191_n 7.65384e-19 $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A2_c_103_n N_B1_c_244_n 0.00914847f $X=1.905 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_120 N_A2_c_102_n N_B1_c_240_n 0.0223862f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A2_c_103_n N_B1_c_243_n 0.02115f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A2_c_104_n N_B1_c_243_n 3.96194e-19 $X=1.79 $Y=1.46 $X2=0 $Y2=0
cc_123 N_A2_c_106_n N_B1_c_243_n 0.00207728f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A2_c_101_n N_A_213_47#_c_313_n 0.00116223f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A2_c_102_n N_A_213_47#_c_313_n 0.00153389f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A2_c_102_n N_A_213_47#_c_315_n 0.0142266f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A2_c_103_n N_A_213_47#_c_315_n 0.00318656f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A2_c_110_n N_A_213_47#_c_315_n 0.00493675f $X=1.705 $Y=1.545 $X2=0
+ $Y2=0
cc_129 N_A2_c_106_n N_A_213_47#_c_315_n 0.0211231f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A2_c_101_n N_A_213_47#_c_300_n 6.08286e-19 $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A2_c_102_n N_A_213_47#_c_320_n 8.26073e-19 $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A2_c_102_n N_A_213_47#_c_301_n 4.98365e-19 $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A2_c_103_n N_A_213_47#_c_301_n 0.00110089f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A2_c_104_n N_A_213_47#_c_301_n 0.00434447f $X=1.79 $Y=1.46 $X2=0 $Y2=0
cc_135 N_A2_c_106_n N_A_213_47#_c_301_n 0.00960727f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A2_c_110_n N_A_27_297#_M1002_d 0.00187091f $X=1.705 $Y=1.545 $X2=0
+ $Y2=0
cc_137 N_A2_c_100_n N_A_27_297#_c_474_n 0.00128062f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A2_c_151_p N_A_27_297#_c_474_n 0.00812827f $X=0.695 $Y=1.545 $X2=0
+ $Y2=0
cc_139 N_A2_c_105_n N_A_27_297#_c_474_n 0.022168f $X=0.525 $Y=1.172 $X2=0 $Y2=0
cc_140 N_A2_c_100_n N_A_27_297#_c_475_n 0.00681523f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A2_c_100_n N_A_27_297#_c_485_n 0.0121086f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A2_c_110_n N_A_27_297#_c_485_n 0.0197085f $X=1.705 $Y=1.545 $X2=0 $Y2=0
cc_143 N_A2_c_151_p N_A_27_297#_c_485_n 0.00871932f $X=0.695 $Y=1.545 $X2=0
+ $Y2=0
cc_144 N_A2_c_105_n N_A_27_297#_c_485_n 0.00280628f $X=0.525 $Y=1.172 $X2=0
+ $Y2=0
cc_145 N_A2_c_103_n N_A_27_297#_c_489_n 0.0121086f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A2_c_110_n N_A_27_297#_c_489_n 0.0280721f $X=1.705 $Y=1.545 $X2=0 $Y2=0
cc_147 N_A2_c_106_n N_A_27_297#_c_489_n 0.00285382f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A2_c_103_n N_A_27_297#_c_492_n 0.00486243f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A2_c_110_n N_A_27_297#_c_476_n 0.00811046f $X=1.705 $Y=1.545 $X2=0
+ $Y2=0
cc_150 N_A2_c_103_n N_A_27_297#_c_494_n 0.00195885f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A2_c_100_n N_A_27_297#_c_479_n 7.83256e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A2_c_105_n N_A_27_297#_c_479_n 0.00134292f $X=0.525 $Y=1.172 $X2=0
+ $Y2=0
cc_153 N_A2_c_100_n N_A_27_297#_c_497_n 5.15302e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A2_c_103_n N_A_27_297#_c_497_n 5.15302e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A2_c_110_n N_A_27_297#_c_497_n 0.0172506f $X=1.705 $Y=1.545 $X2=0 $Y2=0
cc_156 N_A2_c_103_n N_A_27_297#_c_500_n 8.09873e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A2_c_106_n N_A_27_297#_c_500_n 0.00146178f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A2_c_110_n N_VPWR_M1010_d 0.00130005f $X=1.705 $Y=1.545 $X2=-0.19
+ $Y2=-0.24
cc_159 N_A2_c_151_p N_VPWR_M1010_d 5.84953e-19 $X=0.695 $Y=1.545 $X2=-0.19
+ $Y2=-0.24
cc_160 N_A2_c_110_n N_VPWR_M1020_s 0.00186483f $X=1.705 $Y=1.545 $X2=0 $Y2=0
cc_161 N_A2_c_100_n N_VPWR_c_546_n 0.00309049f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A2_c_103_n N_VPWR_c_548_n 0.00309049f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A2_c_103_n N_VPWR_c_553_n 0.00518316f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A2_c_100_n N_VPWR_c_561_n 0.00519834f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A2_c_100_n N_VPWR_c_545_n 0.00767899f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A2_c_103_n N_VPWR_c_545_n 0.00680185f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A2_c_100_n N_VGND_c_747_n 0.00474596f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A2_c_101_n N_VGND_c_747_n 0.0176088f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A2_c_105_n N_VGND_c_747_n 0.0243306f $X=0.525 $Y=1.172 $X2=0 $Y2=0
cc_170 N_A2_c_102_n N_VGND_c_748_n 0.00475459f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A2_c_101_n N_VGND_c_758_n 0.0046653f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A2_c_102_n N_VGND_c_758_n 0.00430895f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A2_c_101_n N_VGND_c_760_n 0.00796999f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A2_c_102_n N_VGND_c_760_n 0.00623871f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A1_c_188_n N_A_213_47#_c_313_n 0.00712196f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A1_c_189_n N_A_213_47#_c_313_n 0.00761603f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A1_c_189_n N_A_213_47#_c_315_n 0.00910922f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A1_c_190_n N_A_213_47#_c_315_n 0.0102215f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A1_c_188_n N_A_213_47#_c_300_n 0.0040234f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A1_c_189_n N_A_213_47#_c_300_n 9.7745e-19 $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A1_c_190_n N_A_213_47#_c_300_n 0.0211043f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A1_c_191_n N_A_213_47#_c_300_n 0.00224326f $X=1.41 $Y=1.202 $X2=0 $Y2=0
cc_183 N_A1_c_192_n N_A_27_297#_c_475_n 5.15302e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A1_c_192_n N_A_27_297#_c_485_n 0.0108454f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A1_c_193_n N_A_27_297#_c_489_n 0.0108454f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_186 N_A1_c_193_n N_A_27_297#_c_492_n 4.72751e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_187 N_A1_c_192_n N_A_27_297#_c_497_n 0.00769006f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A1_c_193_n N_A_27_297#_c_497_n 0.00769006f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A1_c_192_n N_VPWR_c_546_n 0.00173895f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_190 N_A1_c_192_n N_VPWR_c_547_n 0.00519834f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_191 N_A1_c_193_n N_VPWR_c_547_n 0.00519834f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_192 N_A1_c_193_n N_VPWR_c_548_n 0.00173895f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A1_c_192_n N_VPWR_c_545_n 0.00676756f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A1_c_193_n N_VPWR_c_545_n 0.00676756f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A1_c_188_n N_VGND_c_747_n 0.00302624f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A1_c_188_n N_VGND_c_758_n 0.00542163f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A1_c_189_n N_VGND_c_758_n 0.00418572f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A1_c_188_n N_VGND_c_760_n 0.00970348f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A1_c_189_n N_VGND_c_760_n 0.00578774f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_200 B1 N_A_213_47#_c_305_n 0.00228471f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_201 N_B1_c_240_n N_A_213_47#_c_315_n 0.0139202f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_202 N_B1_c_240_n N_A_213_47#_c_320_n 0.00640026f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_203 N_B1_c_244_n N_A_213_47#_c_301_n 0.00506273f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_204 N_B1_c_240_n N_A_213_47#_c_301_n 0.00314306f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_205 N_B1_c_241_n N_A_213_47#_c_301_n 0.00279934f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_206 N_B1_c_245_n N_A_213_47#_c_301_n 0.0046097f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_207 B1 N_A_213_47#_c_301_n 0.0421322f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_208 N_B1_c_243_n N_A_213_47#_c_301_n 0.0299017f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_209 N_B1_c_241_n N_A_213_47#_c_342_n 0.0172949f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_210 B1 N_A_213_47#_c_342_n 0.0235839f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_211 N_B1_c_243_n N_A_213_47#_c_342_n 0.00728832f $X=2.845 $Y=1.202 $X2=0
+ $Y2=0
cc_212 N_B1_c_241_n N_A_213_47#_c_302_n 0.00222925f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_213 N_B1_c_243_n N_A_213_47#_c_302_n 7.80627e-19 $X=2.845 $Y=1.202 $X2=0
+ $Y2=0
cc_214 B1 N_A_213_47#_c_303_n 0.0103841f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_215 N_B1_c_243_n N_A_213_47#_c_303_n 0.00164768f $X=2.845 $Y=1.202 $X2=0
+ $Y2=0
cc_216 N_B1_c_240_n N_A_213_47#_c_349_n 5.73461e-19 $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_217 N_B1_c_244_n N_A_213_47#_c_350_n 0.0037767f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_218 N_B1_c_243_n N_A_213_47#_c_350_n 9.13766e-19 $X=2.845 $Y=1.202 $X2=0
+ $Y2=0
cc_219 B1 N_A_213_47#_c_304_n 0.00275109f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_220 N_B1_c_243_n N_A_213_47#_c_304_n 0.00576975f $X=2.845 $Y=1.202 $X2=0
+ $Y2=0
cc_221 B1 N_A_27_297#_M1011_d 0.00431235f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_222 N_B1_c_244_n N_A_27_297#_c_476_n 2.03034e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_223 N_B1_c_244_n N_A_27_297#_c_477_n 0.0137768f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_224 N_B1_c_245_n N_A_27_297#_c_477_n 0.0134429f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_225 N_B1_c_244_n N_A_27_297#_c_478_n 4.38946e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_226 N_B1_c_245_n N_A_27_297#_c_478_n 0.00878804f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_227 B1 N_A_27_297#_c_478_n 0.0194936f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_228 N_B1_c_243_n N_A_27_297#_c_478_n 9.68667e-19 $X=2.845 $Y=1.202 $X2=0
+ $Y2=0
cc_229 N_B1_c_245_n N_VPWR_c_549_n 0.00677716f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_230 B1 N_VPWR_c_549_n 0.00633255f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_231 N_B1_c_244_n N_VPWR_c_553_n 0.00429453f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_232 N_B1_c_245_n N_VPWR_c_553_n 0.00429425f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_233 N_B1_c_244_n N_VPWR_c_545_n 0.00609021f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_234 N_B1_c_245_n N_VPWR_c_545_n 0.00734732f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_235 N_B1_c_240_n N_VGND_c_748_n 0.00338986f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_236 N_B1_c_240_n N_VGND_c_760_n 0.00604629f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_237 N_B1_c_241_n N_VGND_c_760_n 0.00701283f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_238 N_B1_c_240_n N_VGND_c_762_n 0.00417768f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_239 N_B1_c_241_n N_VGND_c_762_n 0.00430895f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_240 N_B1_c_241_n N_VGND_c_763_n 0.00353715f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A_213_47#_c_315_n N_A_27_297#_c_476_n 0.00791064f $X=2.445 $Y=0.78
+ $X2=0 $Y2=0
cc_242 N_A_213_47#_c_301_n N_A_27_297#_c_476_n 0.0131458f $X=2.61 $Y=1.62 $X2=0
+ $Y2=0
cc_243 N_A_213_47#_M1008_s N_A_27_297#_c_477_n 0.00344383f $X=2.465 $Y=1.485
+ $X2=0 $Y2=0
cc_244 N_A_213_47#_c_350_n N_A_27_297#_c_477_n 0.0147165f $X=2.61 $Y=1.96 $X2=0
+ $Y2=0
cc_245 N_A_213_47#_c_301_n N_A_27_297#_c_478_n 2.79839e-19 $X=2.61 $Y=1.62 $X2=0
+ $Y2=0
cc_246 N_A_213_47#_c_305_n N_VPWR_c_549_n 0.00349953f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_247 N_A_213_47#_c_342_n N_VPWR_c_549_n 0.00248426f $X=3.565 $Y=0.78 $X2=0
+ $Y2=0
cc_248 N_A_213_47#_c_303_n N_VPWR_c_549_n 0.0110476f $X=3.735 $Y=1.155 $X2=0
+ $Y2=0
cc_249 N_A_213_47#_c_305_n N_VPWR_c_550_n 6.17091e-19 $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_250 N_A_213_47#_c_306_n N_VPWR_c_550_n 0.0128989f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_251 N_A_213_47#_c_307_n N_VPWR_c_550_n 0.0128391f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_252 N_A_213_47#_c_308_n N_VPWR_c_550_n 6.06824e-19 $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_253 N_A_213_47#_c_307_n N_VPWR_c_551_n 6.06824e-19 $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_254 N_A_213_47#_c_308_n N_VPWR_c_551_n 0.0128391f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_255 N_A_213_47#_c_309_n N_VPWR_c_551_n 0.0128593f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_256 N_A_213_47#_c_310_n N_VPWR_c_551_n 6.10267e-19 $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_257 N_A_213_47#_c_309_n N_VPWR_c_552_n 7.09884e-19 $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_258 N_A_213_47#_c_310_n N_VPWR_c_552_n 0.0164203f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_259 N_A_213_47#_c_304_n N_VPWR_c_552_n 0.00222608f $X=6.16 $Y=1.202 $X2=0
+ $Y2=0
cc_260 N_A_213_47#_c_305_n N_VPWR_c_555_n 0.00702461f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_261 N_A_213_47#_c_306_n N_VPWR_c_555_n 0.00622633f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_262 N_A_213_47#_c_307_n N_VPWR_c_557_n 0.00622633f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_263 N_A_213_47#_c_308_n N_VPWR_c_557_n 0.00622633f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_264 N_A_213_47#_c_309_n N_VPWR_c_559_n 0.00622633f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_265 N_A_213_47#_c_310_n N_VPWR_c_559_n 0.00661659f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_266 N_A_213_47#_M1008_s N_VPWR_c_545_n 0.00232895f $X=2.465 $Y=1.485 $X2=0
+ $Y2=0
cc_267 N_A_213_47#_c_305_n N_VPWR_c_545_n 0.0136664f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_268 N_A_213_47#_c_306_n N_VPWR_c_545_n 0.0104011f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_269 N_A_213_47#_c_307_n N_VPWR_c_545_n 0.0104011f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_270 N_A_213_47#_c_308_n N_VPWR_c_545_n 0.0104011f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_271 N_A_213_47#_c_309_n N_VPWR_c_545_n 0.0104011f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_272 N_A_213_47#_c_310_n N_VPWR_c_545_n 0.0110154f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_273 N_A_213_47#_c_294_n N_X_c_660_n 0.0106602f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A_213_47#_c_295_n N_X_c_660_n 0.00639957f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A_213_47#_c_296_n N_X_c_660_n 5.17822e-19 $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_276 N_A_213_47#_c_306_n N_X_c_654_n 0.0150944f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_277 N_A_213_47#_c_307_n N_X_c_654_n 0.0151703f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_278 N_A_213_47#_c_391_p N_X_c_654_n 0.0477325f $X=5.29 $Y=1.16 $X2=0 $Y2=0
cc_279 N_A_213_47#_c_304_n N_X_c_654_n 0.00798413f $X=6.16 $Y=1.202 $X2=0 $Y2=0
cc_280 N_A_213_47#_c_305_n N_X_c_655_n 0.0013234f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_281 N_A_213_47#_c_391_p N_X_c_655_n 0.0222834f $X=5.29 $Y=1.16 $X2=0 $Y2=0
cc_282 N_A_213_47#_c_304_n N_X_c_655_n 0.00743165f $X=6.16 $Y=1.202 $X2=0 $Y2=0
cc_283 N_A_213_47#_c_295_n N_X_c_670_n 0.00893375f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_284 N_A_213_47#_c_296_n N_X_c_670_n 0.00893375f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_285 N_A_213_47#_c_391_p N_X_c_670_n 0.0391608f $X=5.29 $Y=1.16 $X2=0 $Y2=0
cc_286 N_A_213_47#_c_304_n N_X_c_670_n 0.00446519f $X=6.16 $Y=1.202 $X2=0 $Y2=0
cc_287 N_A_213_47#_c_294_n N_X_c_674_n 0.00227599f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_288 N_A_213_47#_c_295_n N_X_c_674_n 8.68219e-19 $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_289 N_A_213_47#_c_391_p N_X_c_674_n 0.0211425f $X=5.29 $Y=1.16 $X2=0 $Y2=0
cc_290 N_A_213_47#_c_304_n N_X_c_674_n 0.00218937f $X=6.16 $Y=1.202 $X2=0 $Y2=0
cc_291 N_A_213_47#_c_295_n N_X_c_678_n 5.17822e-19 $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_292 N_A_213_47#_c_296_n N_X_c_678_n 0.00639957f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_293 N_A_213_47#_c_297_n N_X_c_678_n 0.00639957f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_294 N_A_213_47#_c_298_n N_X_c_678_n 5.17822e-19 $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_295 N_A_213_47#_c_308_n N_X_c_656_n 0.0151703f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_296 N_A_213_47#_c_391_p N_X_c_656_n 0.0220321f $X=5.29 $Y=1.16 $X2=0 $Y2=0
cc_297 N_A_213_47#_c_304_n N_X_c_656_n 0.00845362f $X=6.16 $Y=1.202 $X2=0 $Y2=0
cc_298 N_A_213_47#_c_297_n N_X_c_685_n 0.00893375f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_299 N_A_213_47#_c_391_p N_X_c_685_n 0.0177792f $X=5.29 $Y=1.16 $X2=0 $Y2=0
cc_300 N_A_213_47#_c_304_n N_X_c_685_n 0.00500329f $X=6.16 $Y=1.202 $X2=0 $Y2=0
cc_301 N_A_213_47#_c_297_n N_X_c_688_n 5.17822e-19 $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_302 N_A_213_47#_c_298_n N_X_c_688_n 0.00639957f $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_303 N_A_213_47#_c_299_n N_X_c_688_n 0.00506666f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_304 N_A_213_47#_c_309_n N_X_c_657_n 0.0131812f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_305 N_A_213_47#_c_310_n N_X_c_657_n 3.64537e-19 $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_306 N_A_213_47#_c_304_n N_X_c_657_n 0.0069432f $X=6.16 $Y=1.202 $X2=0 $Y2=0
cc_307 N_A_213_47#_c_296_n N_X_c_694_n 8.68219e-19 $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_308 N_A_213_47#_c_297_n N_X_c_694_n 8.68219e-19 $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_309 N_A_213_47#_c_391_p N_X_c_694_n 0.0211425f $X=5.29 $Y=1.16 $X2=0 $Y2=0
cc_310 N_A_213_47#_c_304_n N_X_c_694_n 0.00218937f $X=6.16 $Y=1.202 $X2=0 $Y2=0
cc_311 N_A_213_47#_c_391_p N_X_c_658_n 0.0222834f $X=5.29 $Y=1.16 $X2=0 $Y2=0
cc_312 N_A_213_47#_c_304_n N_X_c_658_n 0.00743165f $X=6.16 $Y=1.202 $X2=0 $Y2=0
cc_313 N_A_213_47#_c_298_n N_X_c_700_n 0.00785862f $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_314 N_A_213_47#_c_299_n N_X_c_700_n 0.00328757f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_315 N_A_213_47#_c_304_n N_X_c_700_n 0.0027324f $X=6.16 $Y=1.202 $X2=0 $Y2=0
cc_316 N_A_213_47#_c_297_n X 0.00215078f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_317 N_A_213_47#_c_308_n X 2.16223e-19 $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_318 N_A_213_47#_c_309_n X 0.00177918f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_319 N_A_213_47#_c_298_n X 0.00309036f $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_320 N_A_213_47#_c_299_n X 0.00214937f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_321 N_A_213_47#_c_310_n X 7.39448e-19 $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_322 N_A_213_47#_c_391_p X 0.0186245f $X=5.29 $Y=1.16 $X2=0 $Y2=0
cc_323 N_A_213_47#_c_304_n X 0.036083f $X=6.16 $Y=1.202 $X2=0 $Y2=0
cc_324 N_A_213_47#_c_315_n N_VGND_M1012_s 0.00924222f $X=2.445 $Y=0.78 $X2=0
+ $Y2=0
cc_325 N_A_213_47#_c_342_n N_VGND_M1019_s 0.0301698f $X=3.565 $Y=0.78 $X2=0
+ $Y2=0
cc_326 N_A_213_47#_c_313_n N_VGND_c_747_n 0.0124356f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_327 N_A_213_47#_c_300_n N_VGND_c_747_n 0.00693247f $X=1.365 $Y=0.78 $X2=0
+ $Y2=0
cc_328 N_A_213_47#_c_315_n N_VGND_c_748_n 0.0247398f $X=2.445 $Y=0.78 $X2=0
+ $Y2=0
cc_329 N_A_213_47#_c_295_n N_VGND_c_749_n 0.00166738f $X=4.28 $Y=0.995 $X2=0
+ $Y2=0
cc_330 N_A_213_47#_c_296_n N_VGND_c_749_n 0.00166854f $X=4.8 $Y=0.995 $X2=0
+ $Y2=0
cc_331 N_A_213_47#_c_297_n N_VGND_c_750_n 0.00166854f $X=5.22 $Y=0.995 $X2=0
+ $Y2=0
cc_332 N_A_213_47#_c_298_n N_VGND_c_750_n 0.00166854f $X=5.74 $Y=0.995 $X2=0
+ $Y2=0
cc_333 N_A_213_47#_c_299_n N_VGND_c_751_n 0.00372401f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_334 N_A_213_47#_c_304_n N_VGND_c_751_n 0.00171941f $X=6.16 $Y=1.202 $X2=0
+ $Y2=0
cc_335 N_A_213_47#_c_294_n N_VGND_c_752_n 0.00541359f $X=3.86 $Y=0.995 $X2=0
+ $Y2=0
cc_336 N_A_213_47#_c_295_n N_VGND_c_752_n 0.00420025f $X=4.28 $Y=0.995 $X2=0
+ $Y2=0
cc_337 N_A_213_47#_c_296_n N_VGND_c_754_n 0.00420025f $X=4.8 $Y=0.995 $X2=0
+ $Y2=0
cc_338 N_A_213_47#_c_297_n N_VGND_c_754_n 0.00420025f $X=5.22 $Y=0.995 $X2=0
+ $Y2=0
cc_339 N_A_213_47#_c_298_n N_VGND_c_756_n 0.00419913f $X=5.74 $Y=0.995 $X2=0
+ $Y2=0
cc_340 N_A_213_47#_c_299_n N_VGND_c_756_n 0.00541359f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_341 N_A_213_47#_c_313_n N_VGND_c_758_n 0.0166744f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_342 N_A_213_47#_c_315_n N_VGND_c_758_n 0.00789631f $X=2.445 $Y=0.78 $X2=0
+ $Y2=0
cc_343 N_A_213_47#_M1007_d N_VGND_c_760_n 0.00216035f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_344 N_A_213_47#_M1014_d N_VGND_c_760_n 0.00215201f $X=2.475 $Y=0.235 $X2=0
+ $Y2=0
cc_345 N_A_213_47#_c_294_n N_VGND_c_760_n 0.0109518f $X=3.86 $Y=0.995 $X2=0
+ $Y2=0
cc_346 N_A_213_47#_c_295_n N_VGND_c_760_n 0.0058995f $X=4.28 $Y=0.995 $X2=0
+ $Y2=0
cc_347 N_A_213_47#_c_296_n N_VGND_c_760_n 0.0058995f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_348 N_A_213_47#_c_297_n N_VGND_c_760_n 0.0058995f $X=5.22 $Y=0.995 $X2=0
+ $Y2=0
cc_349 N_A_213_47#_c_298_n N_VGND_c_760_n 0.00589754f $X=5.74 $Y=0.995 $X2=0
+ $Y2=0
cc_350 N_A_213_47#_c_299_n N_VGND_c_760_n 0.0106331f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_351 N_A_213_47#_c_313_n N_VGND_c_760_n 0.0120611f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_352 N_A_213_47#_c_315_n N_VGND_c_760_n 0.0201864f $X=2.445 $Y=0.78 $X2=0
+ $Y2=0
cc_353 N_A_213_47#_c_320_n N_VGND_c_760_n 0.0112677f $X=2.61 $Y=0.42 $X2=0 $Y2=0
cc_354 N_A_213_47#_c_342_n N_VGND_c_760_n 0.00740747f $X=3.565 $Y=0.78 $X2=0
+ $Y2=0
cc_355 N_A_213_47#_c_315_n N_VGND_c_762_n 0.00224243f $X=2.445 $Y=0.78 $X2=0
+ $Y2=0
cc_356 N_A_213_47#_c_320_n N_VGND_c_762_n 0.0169239f $X=2.61 $Y=0.42 $X2=0 $Y2=0
cc_357 N_A_213_47#_c_342_n N_VGND_c_762_n 0.00243213f $X=3.565 $Y=0.78 $X2=0
+ $Y2=0
cc_358 N_A_213_47#_c_294_n N_VGND_c_763_n 0.00853918f $X=3.86 $Y=0.995 $X2=0
+ $Y2=0
cc_359 N_A_213_47#_c_342_n N_VGND_c_763_n 0.0614132f $X=3.565 $Y=0.78 $X2=0
+ $Y2=0
cc_360 N_A_213_47#_c_315_n A_131_47# 0.00554514f $X=2.445 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_361 N_A_27_297#_c_485_n N_VPWR_M1010_d 0.00368875f $X=1.035 $Y=1.885
+ $X2=-0.19 $Y2=1.305
cc_362 N_A_27_297#_c_489_n N_VPWR_M1020_s 0.00368875f $X=1.975 $Y=1.885 $X2=0
+ $Y2=0
cc_363 N_A_27_297#_c_485_n N_VPWR_c_546_n 0.0138616f $X=1.035 $Y=1.885 $X2=0
+ $Y2=0
cc_364 N_A_27_297#_c_485_n N_VPWR_c_547_n 0.00209157f $X=1.035 $Y=1.885 $X2=0
+ $Y2=0
cc_365 N_A_27_297#_c_489_n N_VPWR_c_547_n 0.00209157f $X=1.975 $Y=1.885 $X2=0
+ $Y2=0
cc_366 N_A_27_297#_c_497_n N_VPWR_c_547_n 0.0189225f $X=1.2 $Y=1.885 $X2=0 $Y2=0
cc_367 N_A_27_297#_c_489_n N_VPWR_c_548_n 0.0138616f $X=1.975 $Y=1.885 $X2=0
+ $Y2=0
cc_368 N_A_27_297#_c_477_n N_VPWR_c_549_n 0.0113145f $X=2.915 $Y=2.38 $X2=0
+ $Y2=0
cc_369 N_A_27_297#_c_478_n N_VPWR_c_549_n 0.0318764f $X=3.08 $Y=1.87 $X2=0 $Y2=0
cc_370 N_A_27_297#_c_489_n N_VPWR_c_553_n 0.00209157f $X=1.975 $Y=1.885 $X2=0
+ $Y2=0
cc_371 N_A_27_297#_c_477_n N_VPWR_c_553_n 0.0575925f $X=2.915 $Y=2.38 $X2=0
+ $Y2=0
cc_372 N_A_27_297#_c_494_n N_VPWR_c_553_n 0.0173953f $X=2.275 $Y=2.38 $X2=0
+ $Y2=0
cc_373 N_A_27_297#_c_475_n N_VPWR_c_561_n 0.0210576f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_374 N_A_27_297#_c_485_n N_VPWR_c_561_n 0.00209157f $X=1.035 $Y=1.885 $X2=0
+ $Y2=0
cc_375 N_A_27_297#_M1010_s N_VPWR_c_545_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_376 N_A_27_297#_M1002_d N_VPWR_c_545_n 0.00231261f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_377 N_A_27_297#_M1015_s N_VPWR_c_545_n 0.00231262f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_378 N_A_27_297#_M1011_d N_VPWR_c_545_n 0.00217517f $X=2.935 $Y=1.485 $X2=0
+ $Y2=0
cc_379 N_A_27_297#_c_475_n N_VPWR_c_545_n 0.0124606f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_380 N_A_27_297#_c_485_n N_VPWR_c_545_n 0.00811004f $X=1.035 $Y=1.885 $X2=0
+ $Y2=0
cc_381 N_A_27_297#_c_489_n N_VPWR_c_545_n 0.00811004f $X=1.975 $Y=1.885 $X2=0
+ $Y2=0
cc_382 N_A_27_297#_c_477_n N_VPWR_c_545_n 0.0347586f $X=2.915 $Y=2.38 $X2=0
+ $Y2=0
cc_383 N_A_27_297#_c_494_n N_VPWR_c_545_n 0.0113829f $X=2.275 $Y=2.38 $X2=0
+ $Y2=0
cc_384 N_A_27_297#_c_497_n N_VPWR_c_545_n 0.0123059f $X=1.2 $Y=1.885 $X2=0 $Y2=0
cc_385 N_VPWR_c_545_n N_X_M1004_d 0.00300692f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_386 N_VPWR_c_545_n N_X_M1013_d 0.00300692f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_387 N_VPWR_c_545_n N_X_M1021_d 0.00300692f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_388 N_VPWR_c_555_n N_X_c_714_n 0.0156407f $X=4.375 $Y=2.72 $X2=0 $Y2=0
cc_389 N_VPWR_c_545_n N_X_c_714_n 0.0103212f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_390 N_VPWR_M1006_s N_X_c_654_n 0.00187091f $X=4.395 $Y=1.485 $X2=0 $Y2=0
cc_391 N_VPWR_c_550_n N_X_c_654_n 0.0171295f $X=4.54 $Y=1.87 $X2=0 $Y2=0
cc_392 N_VPWR_c_557_n N_X_c_718_n 0.0156407f $X=5.315 $Y=2.72 $X2=0 $Y2=0
cc_393 N_VPWR_c_545_n N_X_c_718_n 0.0103212f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_394 N_VPWR_M1018_s N_X_c_656_n 0.00187091f $X=5.335 $Y=1.485 $X2=0 $Y2=0
cc_395 N_VPWR_c_551_n N_X_c_656_n 0.0170955f $X=5.48 $Y=1.87 $X2=0 $Y2=0
cc_396 N_VPWR_c_552_n N_X_c_657_n 0.00774923f $X=6.42 $Y=1.63 $X2=0 $Y2=0
cc_397 N_VPWR_c_559_n N_X_c_723_n 0.0156407f $X=6.265 $Y=2.72 $X2=0 $Y2=0
cc_398 N_VPWR_c_545_n N_X_c_723_n 0.0103212f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_399 N_VPWR_c_552_n N_VGND_c_751_n 0.0103464f $X=6.42 $Y=1.63 $X2=0 $Y2=0
cc_400 N_X_c_670_n N_VGND_M1005_s 0.00500678f $X=4.845 $Y=0.78 $X2=0 $Y2=0
cc_401 N_X_c_685_n N_VGND_M1016_s 0.00579152f $X=5.625 $Y=0.78 $X2=0 $Y2=0
cc_402 N_X_c_670_n N_VGND_c_749_n 0.0198794f $X=4.845 $Y=0.78 $X2=0 $Y2=0
cc_403 N_X_c_685_n N_VGND_c_750_n 0.0198794f $X=5.625 $Y=0.78 $X2=0 $Y2=0
cc_404 X N_VGND_c_751_n 0.00122525f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_405 N_X_c_660_n N_VGND_c_752_n 0.018787f $X=4.07 $Y=0.36 $X2=0 $Y2=0
cc_406 N_X_c_670_n N_VGND_c_752_n 0.00211912f $X=4.845 $Y=0.78 $X2=0 $Y2=0
cc_407 N_X_c_670_n N_VGND_c_754_n 0.00211912f $X=4.845 $Y=0.78 $X2=0 $Y2=0
cc_408 N_X_c_678_n N_VGND_c_754_n 0.018787f $X=5.01 $Y=0.36 $X2=0 $Y2=0
cc_409 N_X_c_685_n N_VGND_c_754_n 0.00211912f $X=5.625 $Y=0.78 $X2=0 $Y2=0
cc_410 N_X_c_688_n N_VGND_c_756_n 0.0188037f $X=5.95 $Y=0.36 $X2=0 $Y2=0
cc_411 N_X_c_700_n N_VGND_c_756_n 0.00222291f $X=5.87 $Y=0.78 $X2=0 $Y2=0
cc_412 N_X_M1001_d N_VGND_c_760_n 0.00215201f $X=3.935 $Y=0.235 $X2=0 $Y2=0
cc_413 N_X_M1009_d N_VGND_c_760_n 0.00215201f $X=4.875 $Y=0.235 $X2=0 $Y2=0
cc_414 N_X_M1017_d N_VGND_c_760_n 0.00215201f $X=5.815 $Y=0.235 $X2=0 $Y2=0
cc_415 N_X_c_660_n N_VGND_c_760_n 0.0121864f $X=4.07 $Y=0.36 $X2=0 $Y2=0
cc_416 N_X_c_670_n N_VGND_c_760_n 0.00897448f $X=4.845 $Y=0.78 $X2=0 $Y2=0
cc_417 N_X_c_678_n N_VGND_c_760_n 0.0121864f $X=5.01 $Y=0.36 $X2=0 $Y2=0
cc_418 N_X_c_685_n N_VGND_c_760_n 0.00528391f $X=5.625 $Y=0.78 $X2=0 $Y2=0
cc_419 N_X_c_688_n N_VGND_c_760_n 0.0121958f $X=5.95 $Y=0.36 $X2=0 $Y2=0
cc_420 N_X_c_700_n N_VGND_c_760_n 0.0039496f $X=5.87 $Y=0.78 $X2=0 $Y2=0
cc_421 N_VGND_c_760_n A_297_47# 0.0111139f $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24
cc_422 N_VGND_c_760_n A_131_47# 0.00318778f $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24
