* File: sky130_fd_sc_hdll__nor4b_2.pxi.spice
* Created: Thu Aug 27 19:17:35 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR4B_2%A N_A_c_91_n N_A_M1001_g N_A_c_95_n N_A_M1000_g
+ N_A_c_96_n N_A_M1008_g N_A_c_92_n N_A_M1015_g A A A N_A_c_94_n A
+ PM_SKY130_FD_SC_HDLL__NOR4B_2%A
x_PM_SKY130_FD_SC_HDLL__NOR4B_2%B N_B_c_134_n N_B_M1004_g N_B_c_138_n
+ N_B_M1010_g N_B_c_139_n N_B_M1014_g N_B_c_135_n N_B_M1011_g B B B N_B_c_137_n
+ B PM_SKY130_FD_SC_HDLL__NOR4B_2%B
x_PM_SKY130_FD_SC_HDLL__NOR4B_2%C N_C_c_174_n N_C_M1006_g N_C_c_178_n
+ N_C_M1007_g N_C_c_179_n N_C_M1009_g N_C_c_175_n N_C_M1012_g C C N_C_c_177_n C
+ PM_SKY130_FD_SC_HDLL__NOR4B_2%C
x_PM_SKY130_FD_SC_HDLL__NOR4B_2%A_754_21# N_A_754_21#_M1002_s
+ N_A_754_21#_M1005_s N_A_754_21#_c_220_n N_A_754_21#_M1013_g
+ N_A_754_21#_c_228_n N_A_754_21#_M1003_g N_A_754_21#_c_221_n
+ N_A_754_21#_M1016_g N_A_754_21#_c_229_n N_A_754_21#_M1017_g
+ N_A_754_21#_c_222_n N_A_754_21#_c_223_n N_A_754_21#_c_224_n
+ N_A_754_21#_c_225_n N_A_754_21#_c_226_n N_A_754_21#_c_232_n
+ N_A_754_21#_c_227_n PM_SKY130_FD_SC_HDLL__NOR4B_2%A_754_21#
x_PM_SKY130_FD_SC_HDLL__NOR4B_2%D_N N_D_N_M1002_g N_D_N_c_296_n N_D_N_c_297_n
+ N_D_N_M1005_g N_D_N_c_291_n N_D_N_c_292_n D_N D_N D_N N_D_N_c_294_n
+ N_D_N_c_295_n PM_SKY130_FD_SC_HDLL__NOR4B_2%D_N
x_PM_SKY130_FD_SC_HDLL__NOR4B_2%A_27_297# N_A_27_297#_M1000_d
+ N_A_27_297#_M1008_d N_A_27_297#_M1014_d N_A_27_297#_c_324_n
+ N_A_27_297#_c_325_n N_A_27_297#_c_326_n N_A_27_297#_c_351_p
+ N_A_27_297#_c_327_n N_A_27_297#_c_328_n N_A_27_297#_c_329_n
+ PM_SKY130_FD_SC_HDLL__NOR4B_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__NOR4B_2%VPWR N_VPWR_M1000_s N_VPWR_M1005_d
+ N_VPWR_c_370_n N_VPWR_c_371_n N_VPWR_c_372_n N_VPWR_c_373_n VPWR
+ N_VPWR_c_374_n N_VPWR_c_369_n N_VPWR_c_376_n
+ PM_SKY130_FD_SC_HDLL__NOR4B_2%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR4B_2%A_305_297# N_A_305_297#_M1010_s
+ N_A_305_297#_M1007_s N_A_305_297#_c_431_n N_A_305_297#_c_427_n
+ N_A_305_297#_c_440_n N_A_305_297#_c_444_p
+ PM_SKY130_FD_SC_HDLL__NOR4B_2%A_305_297#
x_PM_SKY130_FD_SC_HDLL__NOR4B_2%A_514_297# N_A_514_297#_M1007_d
+ N_A_514_297#_M1009_d N_A_514_297#_M1017_s N_A_514_297#_c_448_n
+ N_A_514_297#_c_449_n N_A_514_297#_c_450_n N_A_514_297#_c_451_n
+ N_A_514_297#_c_474_n N_A_514_297#_c_464_n N_A_514_297#_c_467_n
+ PM_SKY130_FD_SC_HDLL__NOR4B_2%A_514_297#
x_PM_SKY130_FD_SC_HDLL__NOR4B_2%Y N_Y_M1001_s N_Y_M1004_d N_Y_M1006_d
+ N_Y_M1013_s N_Y_M1003_d N_Y_c_500_n N_Y_c_491_n N_Y_c_492_n N_Y_c_506_n
+ N_Y_c_493_n N_Y_c_516_n N_Y_c_494_n N_Y_c_519_n N_Y_c_495_n N_Y_c_496_n
+ N_Y_c_497_n N_Y_c_498_n Y Y N_Y_c_499_n PM_SKY130_FD_SC_HDLL__NOR4B_2%Y
x_PM_SKY130_FD_SC_HDLL__NOR4B_2%VGND N_VGND_M1001_d N_VGND_M1015_d
+ N_VGND_M1011_s N_VGND_M1006_s N_VGND_M1012_s N_VGND_M1016_d N_VGND_M1002_d
+ N_VGND_c_584_n N_VGND_c_585_n N_VGND_c_586_n N_VGND_c_587_n N_VGND_c_588_n
+ N_VGND_c_589_n N_VGND_c_590_n N_VGND_c_591_n N_VGND_c_592_n N_VGND_c_593_n
+ N_VGND_c_594_n N_VGND_c_595_n N_VGND_c_596_n VGND N_VGND_c_597_n
+ N_VGND_c_598_n N_VGND_c_599_n N_VGND_c_600_n N_VGND_c_601_n
+ PM_SKY130_FD_SC_HDLL__NOR4B_2%VGND
cc_1 VNB N_A_c_91_n 0.0222857f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_c_92_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB A 0.0210886f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=1.105
cc_4 VNB N_A_c_94_n 0.0426802f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_5 VNB N_B_c_134_n 0.0169338f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_6 VNB N_B_c_135_n 0.0224149f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_7 VNB B 0.0212585f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=1.105
cc_8 VNB N_B_c_137_n 0.0426802f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_9 VNB N_C_c_174_n 0.0224106f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_10 VNB N_C_c_175_n 0.0169173f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_11 VNB C 0.00464355f $X=-0.19 $Y=-0.24 $X2=0.64 $Y2=1.105
cc_12 VNB N_C_c_177_n 0.0421532f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.16
cc_13 VNB N_A_754_21#_c_220_n 0.0164635f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_14 VNB N_A_754_21#_c_221_n 0.0198031f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_15 VNB N_A_754_21#_c_222_n 0.0344846f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.202
cc_16 VNB N_A_754_21#_c_223_n 0.00270102f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.202
cc_17 VNB N_A_754_21#_c_224_n 0.00110808f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=1.19
cc_18 VNB N_A_754_21#_c_225_n 0.0426408f $X=-0.19 $Y=-0.24 $X2=0.725 $Y2=1.18
cc_19 VNB N_A_754_21#_c_226_n 0.0169962f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_754_21#_c_227_n 4.66423e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_D_N_c_291_n 0.00538215f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_22 VNB N_D_N_c_292_n 0.0310875f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_23 VNB D_N 9.68566e-19 $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=1.105
cc_24 VNB N_D_N_c_294_n 0.0213759f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.202
cc_25 VNB N_D_N_c_295_n 0.0184197f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.16
cc_26 VNB N_VPWR_c_369_n 0.250759f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=1.18
cc_27 VNB N_Y_c_491_n 0.00265754f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_28 VNB N_Y_c_492_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.202
cc_29 VNB N_Y_c_493_n 0.0135598f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.18
cc_30 VNB N_Y_c_494_n 0.00351242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_Y_c_495_n 8.60263e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_496_n 0.00287455f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_Y_c_497_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_Y_c_498_n 0.0032614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_584_n 0.00991007f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.16
cc_36 VNB N_VGND_c_585_n 0.0332649f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_37 VNB N_VGND_c_586_n 0.0199314f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.18
cc_38 VNB N_VGND_c_587_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0.725 $Y2=1.18
cc_39 VNB N_VGND_c_588_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_589_n 0.00736823f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_590_n 0.0199258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_591_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_592_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_593_n 0.0200006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_594_n 0.00394313f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_595_n 0.0210437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_596_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_597_n 0.0113717f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_598_n 0.317185f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_599_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_600_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_601_n 0.0282059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VPB N_A_c_95_n 0.0203249f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_54 VPB N_A_c_96_n 0.0161064f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_55 VPB N_A_c_94_n 0.022695f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_56 VPB N_B_c_138_n 0.0161064f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_57 VPB N_B_c_139_n 0.0203249f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_58 VPB N_B_c_137_n 0.022695f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_59 VPB N_C_c_178_n 0.0203249f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_60 VPB N_C_c_179_n 0.0160856f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_61 VPB N_C_c_177_n 0.0226924f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.16
cc_62 VPB N_A_754_21#_c_228_n 0.0164093f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_63 VPB N_A_754_21#_c_229_n 0.0192858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_754_21#_c_222_n 0.021283f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.202
cc_65 VPB N_A_754_21#_c_225_n 0.0221207f $X=-0.19 $Y=1.305 $X2=0.725 $Y2=1.18
cc_66 VPB N_A_754_21#_c_232_n 0.0128965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_754_21#_c_227_n 0.0165709f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_D_N_c_296_n 0.038113f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_69 VPB N_D_N_c_297_n 0.0324146f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_70 VPB N_D_N_c_292_n 0.00786212f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_71 VPB D_N 0.0399569f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=1.105
cc_72 VPB N_A_27_297#_c_324_n 0.0332602f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_73 VPB N_A_27_297#_c_325_n 0.00185169f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_297#_c_326_n 0.0103829f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_297#_c_327_n 0.00634455f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.16
cc_76 VPB N_A_27_297#_c_328_n 0.0047306f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.18
cc_77 VPB N_A_27_297#_c_329_n 0.00234762f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.19
cc_78 VPB N_VPWR_c_370_n 0.00495424f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_79 VPB N_VPWR_c_371_n 0.00518f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=1.105
cc_80 VPB N_VPWR_c_372_n 0.112137f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_373_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.202
cc_82 VPB N_VPWR_c_374_n 0.0113717f $X=-0.19 $Y=1.305 $X2=0.725 $Y2=1.18
cc_83 VPB N_VPWR_c_369_n 0.0571001f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=1.18
cc_84 VPB N_VPWR_c_376_n 0.0233763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_305_297#_c_427_n 0.0111956f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_86 VPB N_A_514_297#_c_448_n 0.00610595f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_87 VPB N_A_514_297#_c_449_n 0.00185169f $X=-0.19 $Y=1.305 $X2=0.64 $Y2=1.105
cc_88 VPB N_A_514_297#_c_450_n 0.00646983f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=1.105
cc_89 VPB N_A_514_297#_c_451_n 0.00325504f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_Y_c_499_n 0.00424114f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 N_A_c_92_n N_B_c_134_n 0.0242921f $X=0.99 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_92 N_A_c_96_n N_B_c_138_n 0.00985632f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_93 A B 0.0164404f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_94 A N_B_c_137_n 0.00575962f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_95 N_A_c_94_n N_B_c_137_n 0.0242921f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_96 N_A_c_95_n N_A_27_297#_c_324_n 0.0113204f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A_c_96_n N_A_27_297#_c_324_n 6.54437e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A_c_95_n N_A_27_297#_c_325_n 0.0137916f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A_c_96_n N_A_27_297#_c_325_n 0.0156202f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_100 A N_A_27_297#_c_325_n 0.0459115f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_101 N_A_c_94_n N_A_27_297#_c_325_n 0.00759056f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_102 N_A_c_95_n N_A_27_297#_c_326_n 0.00118933f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_103 A N_A_27_297#_c_326_n 0.0276437f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_104 N_A_c_94_n N_A_27_297#_c_326_n 3.16729e-19 $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_105 A N_A_27_297#_c_327_n 0.00109081f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_106 A N_A_27_297#_c_329_n 0.0214236f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_107 N_A_c_95_n N_VPWR_c_370_n 0.00553644f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A_c_96_n N_VPWR_c_370_n 0.00295479f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A_c_96_n N_VPWR_c_372_n 0.00702461f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A_c_95_n N_VPWR_c_369_n 0.0127552f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A_c_96_n N_VPWR_c_369_n 0.0124344f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A_c_95_n N_VPWR_c_376_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_c_91_n N_Y_c_500_n 0.00539651f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A_c_92_n N_Y_c_491_n 0.0106151f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_115 A N_Y_c_491_n 0.0328995f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_116 N_A_c_91_n N_Y_c_492_n 0.00269085f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_117 A N_Y_c_492_n 0.030835f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_118 N_A_c_94_n N_Y_c_492_n 0.00486271f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_119 N_A_c_92_n N_Y_c_506_n 5.32212e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A_c_91_n N_VGND_c_585_n 0.00495051f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_121 A N_VGND_c_585_n 0.0209094f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_122 N_A_c_91_n N_VGND_c_586_n 0.00541359f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_c_92_n N_VGND_c_586_n 0.00437852f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A_c_92_n N_VGND_c_587_n 0.00268723f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_c_91_n N_VGND_c_598_n 0.0106981f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_c_92_n N_VGND_c_598_n 0.00615622f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_127 B C 0.0158042f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_128 B N_C_c_177_n 0.00564877f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_129 N_B_c_138_n N_A_27_297#_c_327_n 0.017847f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_130 N_B_c_139_n N_A_27_297#_c_327_n 0.0111266f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_131 B N_A_27_297#_c_327_n 0.0605092f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_132 N_B_c_137_n N_A_27_297#_c_327_n 0.00793122f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_133 N_B_c_138_n N_A_27_297#_c_328_n 5.70824e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_134 N_B_c_139_n N_A_27_297#_c_328_n 0.00937268f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_135 N_B_c_138_n N_VPWR_c_372_n 0.00702461f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_136 N_B_c_139_n N_VPWR_c_372_n 0.00429453f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_137 N_B_c_138_n N_VPWR_c_369_n 0.0126324f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_138 N_B_c_139_n N_VPWR_c_369_n 0.00739666f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_139 N_B_c_139_n N_A_305_297#_c_427_n 0.01253f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_140 N_B_c_139_n N_A_514_297#_c_450_n 3.61833e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_141 B N_A_514_297#_c_450_n 0.0149784f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_142 N_B_c_134_n N_Y_c_491_n 0.01006f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_143 N_B_c_134_n N_Y_c_506_n 0.00644736f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_144 N_B_c_135_n N_Y_c_493_n 0.01289f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_145 B N_Y_c_493_n 0.0613753f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_146 N_B_c_134_n N_Y_c_496_n 0.00157949f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_147 B N_Y_c_496_n 0.0252639f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_148 N_B_c_137_n N_Y_c_496_n 0.00486271f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_149 N_B_c_134_n N_VGND_c_587_n 0.00268723f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_150 N_B_c_134_n N_VGND_c_598_n 0.00598581f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_151 N_B_c_135_n N_VGND_c_598_n 0.00745263f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_152 N_B_c_134_n N_VGND_c_600_n 0.00423334f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_153 N_B_c_135_n N_VGND_c_600_n 0.00437852f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_154 N_B_c_135_n N_VGND_c_601_n 0.00483063f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_155 N_C_c_175_n N_A_754_21#_c_220_n 0.0236835f $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_156 N_C_c_179_n N_A_754_21#_c_228_n 0.00954312f $X=3.4 $Y=1.41 $X2=0 $Y2=0
cc_157 C N_A_754_21#_c_222_n 0.00262876f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_158 N_C_c_177_n N_A_754_21#_c_222_n 0.0236835f $X=3.4 $Y=1.202 $X2=0 $Y2=0
cc_159 N_C_c_178_n N_A_27_297#_c_327_n 3.29218e-19 $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_160 N_C_c_178_n N_VPWR_c_372_n 0.00429453f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_161 N_C_c_179_n N_VPWR_c_372_n 0.00702461f $X=3.4 $Y=1.41 $X2=0 $Y2=0
cc_162 N_C_c_178_n N_VPWR_c_369_n 0.00739666f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_163 N_C_c_179_n N_VPWR_c_369_n 0.0126324f $X=3.4 $Y=1.41 $X2=0 $Y2=0
cc_164 N_C_c_178_n N_A_305_297#_c_427_n 0.0132915f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_165 N_C_c_178_n N_A_514_297#_c_448_n 0.00745176f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_166 N_C_c_179_n N_A_514_297#_c_448_n 5.45151e-19 $X=3.4 $Y=1.41 $X2=0 $Y2=0
cc_167 N_C_c_178_n N_A_514_297#_c_449_n 0.0113508f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_168 N_C_c_179_n N_A_514_297#_c_449_n 0.0155666f $X=3.4 $Y=1.41 $X2=0 $Y2=0
cc_169 C N_A_514_297#_c_449_n 0.0459115f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_170 N_C_c_177_n N_A_514_297#_c_449_n 0.00759056f $X=3.4 $Y=1.202 $X2=0 $Y2=0
cc_171 N_C_c_178_n N_A_514_297#_c_450_n 0.00144466f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_172 N_C_c_177_n N_A_514_297#_c_450_n 3.83669e-19 $X=3.4 $Y=1.202 $X2=0 $Y2=0
cc_173 C N_A_514_297#_c_451_n 0.0128541f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_174 N_C_c_174_n N_Y_c_493_n 0.0112792f $X=2.905 $Y=0.995 $X2=0 $Y2=0
cc_175 C N_Y_c_493_n 0.00619376f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_176 N_C_c_174_n N_Y_c_516_n 0.0110728f $X=2.905 $Y=0.995 $X2=0 $Y2=0
cc_177 N_C_c_175_n N_Y_c_494_n 0.0106151f $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_178 C N_Y_c_494_n 0.024099f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_179 N_C_c_175_n N_Y_c_519_n 5.32212e-19 $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_180 N_C_c_177_n N_Y_c_495_n 3.42221e-19 $X=3.4 $Y=1.202 $X2=0 $Y2=0
cc_181 N_C_c_174_n N_Y_c_497_n 0.00119564f $X=2.905 $Y=0.995 $X2=0 $Y2=0
cc_182 C N_Y_c_497_n 0.030835f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_183 N_C_c_177_n N_Y_c_497_n 0.00486271f $X=3.4 $Y=1.202 $X2=0 $Y2=0
cc_184 C N_Y_c_499_n 0.00934461f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_185 N_C_c_177_n N_Y_c_499_n 3.21364e-19 $X=3.4 $Y=1.202 $X2=0 $Y2=0
cc_186 N_C_c_175_n N_VGND_c_588_n 0.00268723f $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_187 N_C_c_174_n N_VGND_c_591_n 0.00423334f $X=2.905 $Y=0.995 $X2=0 $Y2=0
cc_188 N_C_c_175_n N_VGND_c_591_n 0.00437852f $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_189 N_C_c_174_n N_VGND_c_598_n 0.00728222f $X=2.905 $Y=0.995 $X2=0 $Y2=0
cc_190 N_C_c_175_n N_VGND_c_598_n 0.00615622f $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_191 N_C_c_174_n N_VGND_c_601_n 0.00483063f $X=2.905 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_754_21#_c_232_n N_D_N_c_297_n 0.00184336f $X=5.095 $Y=2.285 $X2=0
+ $Y2=0
cc_193 N_A_754_21#_c_227_n N_D_N_c_297_n 0.00148108f $X=5.042 $Y=2.035 $X2=0
+ $Y2=0
cc_194 N_A_754_21#_c_224_n N_D_N_c_291_n 0.0148758f $X=4.885 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A_754_21#_c_225_n N_D_N_c_291_n 7.43407e-19 $X=4.885 $Y=1.16 $X2=0
+ $Y2=0
cc_196 N_A_754_21#_c_226_n N_D_N_c_291_n 0.0011748f $X=5.095 $Y=0.66 $X2=0 $Y2=0
cc_197 N_A_754_21#_c_227_n N_D_N_c_291_n 0.00329272f $X=5.042 $Y=2.035 $X2=0
+ $Y2=0
cc_198 N_A_754_21#_c_224_n N_D_N_c_292_n 5.13953e-19 $X=4.885 $Y=1.16 $X2=0
+ $Y2=0
cc_199 N_A_754_21#_c_225_n N_D_N_c_292_n 0.0212545f $X=4.885 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A_754_21#_c_227_n N_D_N_c_292_n 0.0165538f $X=5.042 $Y=2.035 $X2=0
+ $Y2=0
cc_201 N_A_754_21#_c_227_n D_N 0.0220439f $X=5.042 $Y=2.035 $X2=0 $Y2=0
cc_202 N_A_754_21#_c_223_n N_D_N_c_294_n 0.00455001f $X=4.95 $Y=1.075 $X2=0
+ $Y2=0
cc_203 N_A_754_21#_c_226_n N_D_N_c_294_n 0.00356691f $X=5.095 $Y=0.66 $X2=0
+ $Y2=0
cc_204 N_A_754_21#_c_228_n N_VPWR_c_372_n 0.00429453f $X=3.87 $Y=1.41 $X2=0
+ $Y2=0
cc_205 N_A_754_21#_c_229_n N_VPWR_c_372_n 0.00429453f $X=4.34 $Y=1.41 $X2=0
+ $Y2=0
cc_206 N_A_754_21#_c_232_n N_VPWR_c_372_n 0.0213169f $X=5.095 $Y=2.285 $X2=0
+ $Y2=0
cc_207 N_A_754_21#_M1005_s N_VPWR_c_369_n 0.00266577f $X=4.97 $Y=2.065 $X2=0
+ $Y2=0
cc_208 N_A_754_21#_c_228_n N_VPWR_c_369_n 0.00609021f $X=3.87 $Y=1.41 $X2=0
+ $Y2=0
cc_209 N_A_754_21#_c_229_n N_VPWR_c_369_n 0.00734734f $X=4.34 $Y=1.41 $X2=0
+ $Y2=0
cc_210 N_A_754_21#_c_232_n N_VPWR_c_369_n 0.0134053f $X=5.095 $Y=2.285 $X2=0
+ $Y2=0
cc_211 N_A_754_21#_c_228_n N_A_514_297#_c_451_n 2.98195e-19 $X=3.87 $Y=1.41
+ $X2=0 $Y2=0
cc_212 N_A_754_21#_c_228_n N_A_514_297#_c_464_n 0.0143578f $X=3.87 $Y=1.41 $X2=0
+ $Y2=0
cc_213 N_A_754_21#_c_229_n N_A_514_297#_c_464_n 0.0116061f $X=4.34 $Y=1.41 $X2=0
+ $Y2=0
cc_214 N_A_754_21#_c_232_n N_A_514_297#_c_464_n 0.0135088f $X=5.095 $Y=2.285
+ $X2=0 $Y2=0
cc_215 N_A_754_21#_c_225_n N_A_514_297#_c_467_n 0.00665307f $X=4.885 $Y=1.16
+ $X2=0 $Y2=0
cc_216 N_A_754_21#_c_227_n N_A_514_297#_c_467_n 0.0390848f $X=5.042 $Y=2.035
+ $X2=0 $Y2=0
cc_217 N_A_754_21#_c_220_n N_Y_c_494_n 0.0122977f $X=3.845 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A_754_21#_c_220_n N_Y_c_519_n 0.00644736f $X=3.845 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A_754_21#_c_221_n N_Y_c_519_n 0.00600712f $X=4.315 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_754_21#_c_220_n N_Y_c_495_n 0.00200685f $X=3.845 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A_754_21#_c_221_n N_Y_c_495_n 0.00265654f $X=4.315 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A_754_21#_c_222_n N_Y_c_495_n 0.00719288f $X=4.44 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A_754_21#_c_223_n N_Y_c_495_n 0.00443109f $X=4.95 $Y=1.075 $X2=0 $Y2=0
cc_224 N_A_754_21#_c_220_n N_Y_c_498_n 0.00224457f $X=3.845 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A_754_21#_c_221_n N_Y_c_498_n 0.00256543f $X=4.315 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A_754_21#_c_222_n N_Y_c_498_n 0.00174649f $X=4.44 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A_754_21#_c_226_n N_Y_c_498_n 3.25184e-19 $X=5.095 $Y=0.66 $X2=0 $Y2=0
cc_228 N_A_754_21#_c_228_n N_Y_c_499_n 0.00150282f $X=3.87 $Y=1.41 $X2=0 $Y2=0
cc_229 N_A_754_21#_c_229_n N_Y_c_499_n 0.013014f $X=4.34 $Y=1.41 $X2=0 $Y2=0
cc_230 N_A_754_21#_c_222_n N_Y_c_499_n 0.0345934f $X=4.44 $Y=1.16 $X2=0 $Y2=0
cc_231 N_A_754_21#_c_224_n N_Y_c_499_n 0.0101408f $X=4.885 $Y=1.16 $X2=0 $Y2=0
cc_232 N_A_754_21#_c_225_n N_Y_c_499_n 0.00880525f $X=4.885 $Y=1.16 $X2=0 $Y2=0
cc_233 N_A_754_21#_c_227_n N_Y_c_499_n 0.0170371f $X=5.042 $Y=2.035 $X2=0 $Y2=0
cc_234 N_A_754_21#_c_220_n N_VGND_c_588_n 0.00268723f $X=3.845 $Y=0.995 $X2=0
+ $Y2=0
cc_235 N_A_754_21#_c_221_n N_VGND_c_589_n 0.00672154f $X=4.315 $Y=0.995 $X2=0
+ $Y2=0
cc_236 N_A_754_21#_c_225_n N_VGND_c_589_n 0.00973477f $X=4.885 $Y=1.16 $X2=0
+ $Y2=0
cc_237 N_A_754_21#_c_226_n N_VGND_c_589_n 0.040929f $X=5.095 $Y=0.66 $X2=0 $Y2=0
cc_238 N_A_754_21#_c_226_n N_VGND_c_590_n 0.0172241f $X=5.095 $Y=0.66 $X2=0
+ $Y2=0
cc_239 N_A_754_21#_c_220_n N_VGND_c_593_n 0.00423334f $X=3.845 $Y=0.995 $X2=0
+ $Y2=0
cc_240 N_A_754_21#_c_221_n N_VGND_c_593_n 0.00541359f $X=4.315 $Y=0.995 $X2=0
+ $Y2=0
cc_241 N_A_754_21#_c_226_n N_VGND_c_595_n 0.0139512f $X=5.095 $Y=0.66 $X2=0
+ $Y2=0
cc_242 N_A_754_21#_c_220_n N_VGND_c_598_n 0.00587047f $X=3.845 $Y=0.995 $X2=0
+ $Y2=0
cc_243 N_A_754_21#_c_221_n N_VGND_c_598_n 0.0110773f $X=4.315 $Y=0.995 $X2=0
+ $Y2=0
cc_244 N_A_754_21#_c_226_n N_VGND_c_598_n 0.0126265f $X=5.095 $Y=0.66 $X2=0
+ $Y2=0
cc_245 N_D_N_c_297_n N_VPWR_c_371_n 0.00479105f $X=5.33 $Y=1.99 $X2=0 $Y2=0
cc_246 D_N N_VPWR_c_371_n 0.00618824f $X=5.67 $Y=1.445 $X2=0 $Y2=0
cc_247 N_D_N_c_297_n N_VPWR_c_372_n 0.00743866f $X=5.33 $Y=1.99 $X2=0 $Y2=0
cc_248 N_D_N_c_297_n N_VPWR_c_369_n 0.0153164f $X=5.33 $Y=1.99 $X2=0 $Y2=0
cc_249 D_N N_VPWR_c_369_n 0.00844898f $X=5.67 $Y=1.445 $X2=0 $Y2=0
cc_250 N_D_N_c_294_n N_VGND_c_589_n 0.00167989f $X=5.392 $Y=0.995 $X2=0 $Y2=0
cc_251 N_D_N_c_291_n N_VGND_c_590_n 0.0105684f $X=5.615 $Y=1.18 $X2=0 $Y2=0
cc_252 N_D_N_c_292_n N_VGND_c_590_n 0.00280284f $X=5.37 $Y=1.16 $X2=0 $Y2=0
cc_253 N_D_N_c_294_n N_VGND_c_590_n 0.00512723f $X=5.392 $Y=0.995 $X2=0 $Y2=0
cc_254 N_D_N_c_295_n N_VGND_c_590_n 0.00514577f $X=5.75 $Y=1.285 $X2=0 $Y2=0
cc_255 N_D_N_c_294_n N_VGND_c_595_n 0.00510437f $X=5.392 $Y=0.995 $X2=0 $Y2=0
cc_256 N_D_N_c_294_n N_VGND_c_598_n 0.00512902f $X=5.392 $Y=0.995 $X2=0 $Y2=0
cc_257 N_A_27_297#_c_325_n N_VPWR_M1000_s 0.00182839f $X=1.075 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_258 N_A_27_297#_c_324_n N_VPWR_c_370_n 0.0413039f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_259 N_A_27_297#_c_325_n N_VPWR_c_370_n 0.0139937f $X=1.075 $Y=1.54 $X2=0
+ $Y2=0
cc_260 N_A_27_297#_c_351_p N_VPWR_c_372_n 0.0149311f $X=1.2 $Y=2.3 $X2=0 $Y2=0
cc_261 N_A_27_297#_M1000_d N_VPWR_c_369_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_262 N_A_27_297#_M1008_d N_VPWR_c_369_n 0.00370124f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_263 N_A_27_297#_M1014_d N_VPWR_c_369_n 0.00218346f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_264 N_A_27_297#_c_324_n N_VPWR_c_369_n 0.0128576f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_265 N_A_27_297#_c_351_p N_VPWR_c_369_n 0.00955092f $X=1.2 $Y=2.3 $X2=0 $Y2=0
cc_266 N_A_27_297#_c_324_n N_VPWR_c_376_n 0.0217765f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_267 N_A_27_297#_c_327_n N_A_305_297#_M1010_s 0.00182839f $X=1.925 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_268 N_A_27_297#_c_327_n N_A_305_297#_c_431_n 0.0139767f $X=1.925 $Y=1.54
+ $X2=0 $Y2=0
cc_269 N_A_27_297#_c_328_n N_A_305_297#_c_431_n 0.0250219f $X=2.14 $Y=1.63 $X2=0
+ $Y2=0
cc_270 N_A_27_297#_M1014_d N_A_305_297#_c_427_n 0.00510164f $X=1.995 $Y=1.485
+ $X2=0 $Y2=0
cc_271 N_A_27_297#_c_327_n N_A_305_297#_c_427_n 0.00238643f $X=1.925 $Y=1.54
+ $X2=0 $Y2=0
cc_272 N_A_27_297#_c_328_n N_A_305_297#_c_427_n 0.0241709f $X=2.14 $Y=1.63 $X2=0
+ $Y2=0
cc_273 N_A_27_297#_c_328_n N_A_514_297#_c_448_n 0.042489f $X=2.14 $Y=1.63 $X2=0
+ $Y2=0
cc_274 N_A_27_297#_c_327_n N_A_514_297#_c_450_n 0.0159284f $X=1.925 $Y=1.54
+ $X2=0 $Y2=0
cc_275 N_A_27_297#_c_327_n N_Y_c_491_n 0.00299046f $X=1.925 $Y=1.54 $X2=0 $Y2=0
cc_276 N_A_27_297#_c_327_n N_Y_c_496_n 0.00220237f $X=1.925 $Y=1.54 $X2=0 $Y2=0
cc_277 N_A_27_297#_c_326_n N_VGND_c_585_n 5.77871e-19 $X=0.425 $Y=1.54 $X2=0
+ $Y2=0
cc_278 N_VPWR_c_369_n N_A_305_297#_M1010_s 0.00297226f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_279 N_VPWR_c_369_n N_A_305_297#_M1007_s 0.00297226f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_280 N_VPWR_c_372_n N_A_305_297#_c_427_n 0.0904664f $X=5.44 $Y=2.72 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_369_n N_A_305_297#_c_427_n 0.0556336f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_282 N_VPWR_c_372_n N_A_305_297#_c_440_n 0.0134651f $X=5.44 $Y=2.72 $X2=0
+ $Y2=0
cc_283 N_VPWR_c_369_n N_A_305_297#_c_440_n 0.00808434f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_369_n N_A_514_297#_M1007_d 0.00218346f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_285 N_VPWR_c_369_n N_A_514_297#_M1009_d 0.00297222f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_286 N_VPWR_c_369_n N_A_514_297#_M1017_s 0.00234877f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_287 N_VPWR_c_372_n N_A_514_297#_c_474_n 0.015002f $X=5.44 $Y=2.72 $X2=0 $Y2=0
cc_288 N_VPWR_c_369_n N_A_514_297#_c_474_n 0.00962794f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_289 N_VPWR_c_372_n N_A_514_297#_c_464_n 0.0546052f $X=5.44 $Y=2.72 $X2=0
+ $Y2=0
cc_290 N_VPWR_c_369_n N_A_514_297#_c_464_n 0.0333461f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_369_n N_Y_M1003_d 0.00232895f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_292 N_A_305_297#_c_427_n N_A_514_297#_M1007_d 0.00510164f $X=3.08 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_293 N_A_305_297#_c_427_n N_A_514_297#_c_448_n 0.0249537f $X=3.08 $Y=2.38
+ $X2=0 $Y2=0
cc_294 N_A_305_297#_c_444_p N_A_514_297#_c_448_n 0.0205381f $X=3.165 $Y=1.96
+ $X2=0 $Y2=0
cc_295 N_A_305_297#_M1007_s N_A_514_297#_c_449_n 0.00182839f $X=3.02 $Y=1.485
+ $X2=0 $Y2=0
cc_296 N_A_305_297#_c_427_n N_A_514_297#_c_449_n 0.00346334f $X=3.08 $Y=2.38
+ $X2=0 $Y2=0
cc_297 N_A_305_297#_c_444_p N_A_514_297#_c_449_n 0.0139767f $X=3.165 $Y=1.96
+ $X2=0 $Y2=0
cc_298 N_A_514_297#_c_464_n N_Y_M1003_d 0.00352392f $X=4.45 $Y=2.38 $X2=0 $Y2=0
cc_299 N_A_514_297#_c_450_n N_Y_c_493_n 0.00764905f $X=2.86 $Y=1.54 $X2=0 $Y2=0
cc_300 N_A_514_297#_c_451_n N_Y_c_494_n 0.00374609f $X=3.635 $Y=1.625 $X2=0
+ $Y2=0
cc_301 N_A_514_297#_M1017_s N_Y_c_499_n 0.00224845f $X=4.43 $Y=1.485 $X2=0 $Y2=0
cc_302 N_A_514_297#_c_451_n N_Y_c_499_n 0.00221338f $X=3.635 $Y=1.625 $X2=0
+ $Y2=0
cc_303 N_A_514_297#_c_464_n N_Y_c_499_n 0.0176569f $X=4.45 $Y=2.38 $X2=0 $Y2=0
cc_304 N_A_514_297#_c_467_n N_Y_c_499_n 2.65999e-19 $X=4.575 $Y=1.96 $X2=0 $Y2=0
cc_305 N_Y_c_491_n N_VGND_M1015_d 0.00162089f $X=1.455 $Y=0.815 $X2=0 $Y2=0
cc_306 N_Y_c_493_n N_VGND_M1011_s 0.00281828f $X=2.95 $Y=0.815 $X2=0 $Y2=0
cc_307 N_Y_c_493_n N_VGND_M1006_s 0.00281828f $X=2.95 $Y=0.815 $X2=0 $Y2=0
cc_308 N_Y_c_494_n N_VGND_M1012_s 0.00162089f $X=3.89 $Y=0.815 $X2=0 $Y2=0
cc_309 N_Y_c_492_n N_VGND_c_585_n 0.00834802f $X=0.895 $Y=0.815 $X2=0 $Y2=0
cc_310 N_Y_c_500_n N_VGND_c_586_n 0.0231806f $X=0.73 $Y=0.39 $X2=0 $Y2=0
cc_311 N_Y_c_491_n N_VGND_c_586_n 0.00254521f $X=1.455 $Y=0.815 $X2=0 $Y2=0
cc_312 N_Y_c_491_n N_VGND_c_587_n 0.0122559f $X=1.455 $Y=0.815 $X2=0 $Y2=0
cc_313 N_Y_c_494_n N_VGND_c_588_n 0.0122559f $X=3.89 $Y=0.815 $X2=0 $Y2=0
cc_314 N_Y_c_519_n N_VGND_c_589_n 0.0291386f $X=4.105 $Y=0.39 $X2=0 $Y2=0
cc_315 N_Y_c_498_n N_VGND_c_589_n 0.0110997f $X=4.08 $Y=0.815 $X2=0 $Y2=0
cc_316 N_Y_c_493_n N_VGND_c_591_n 0.00198695f $X=2.95 $Y=0.815 $X2=0 $Y2=0
cc_317 N_Y_c_516_n N_VGND_c_591_n 0.0231806f $X=3.165 $Y=0.39 $X2=0 $Y2=0
cc_318 N_Y_c_494_n N_VGND_c_591_n 0.00254521f $X=3.89 $Y=0.815 $X2=0 $Y2=0
cc_319 N_Y_c_494_n N_VGND_c_593_n 0.00198695f $X=3.89 $Y=0.815 $X2=0 $Y2=0
cc_320 N_Y_c_519_n N_VGND_c_593_n 0.0223932f $X=4.105 $Y=0.39 $X2=0 $Y2=0
cc_321 N_Y_M1001_s N_VGND_c_598_n 0.00304143f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_322 N_Y_M1004_d N_VGND_c_598_n 0.00304143f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_323 N_Y_M1006_d N_VGND_c_598_n 0.00304143f $X=2.98 $Y=0.235 $X2=0 $Y2=0
cc_324 N_Y_M1013_s N_VGND_c_598_n 0.0025535f $X=3.92 $Y=0.235 $X2=0 $Y2=0
cc_325 N_Y_c_500_n N_VGND_c_598_n 0.0143352f $X=0.73 $Y=0.39 $X2=0 $Y2=0
cc_326 N_Y_c_491_n N_VGND_c_598_n 0.0094839f $X=1.455 $Y=0.815 $X2=0 $Y2=0
cc_327 N_Y_c_506_n N_VGND_c_598_n 0.0143352f $X=1.67 $Y=0.39 $X2=0 $Y2=0
cc_328 N_Y_c_493_n N_VGND_c_598_n 0.0115853f $X=2.95 $Y=0.815 $X2=0 $Y2=0
cc_329 N_Y_c_516_n N_VGND_c_598_n 0.0143352f $X=3.165 $Y=0.39 $X2=0 $Y2=0
cc_330 N_Y_c_494_n N_VGND_c_598_n 0.0094839f $X=3.89 $Y=0.815 $X2=0 $Y2=0
cc_331 N_Y_c_519_n N_VGND_c_598_n 0.0141395f $X=4.105 $Y=0.39 $X2=0 $Y2=0
cc_332 N_Y_c_491_n N_VGND_c_600_n 0.00198695f $X=1.455 $Y=0.815 $X2=0 $Y2=0
cc_333 N_Y_c_506_n N_VGND_c_600_n 0.0231806f $X=1.67 $Y=0.39 $X2=0 $Y2=0
cc_334 N_Y_c_493_n N_VGND_c_600_n 0.00254521f $X=2.95 $Y=0.815 $X2=0 $Y2=0
cc_335 N_Y_c_493_n N_VGND_c_601_n 0.0564849f $X=2.95 $Y=0.815 $X2=0 $Y2=0
