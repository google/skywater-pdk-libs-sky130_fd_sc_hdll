* File: sky130_fd_sc_hdll__clkinv_8.spice
* Created: Thu Aug 27 19:03:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__clkinv_8.pex.spice"
.subckt sky130_fd_sc_hdll__clkinv_8  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_M1000_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0693 PD=1.37 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.2 SB=75003.8
+ A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.7 SB=75003.3
+ A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1004_d N_A_M1005_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0693 PD=0.75 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1 SB=75002.8
+ A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.6 SB=75002.4
+ A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1007_d N_A_M1010_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0798 PD=0.75 PS=0.8 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.1 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A_M1012_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.42 AD=0.0798
+ AS=0.0798 PD=0.8 PS=0.8 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75002.6 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1012_d N_A_M1015_g N_Y_M1015_s VNB NSHORT L=0.15 W=0.42 AD=0.0798
+ AS=0.0798 PD=0.8 PS=0.8 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75003.2 SB=75000.8
+ A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_M1019_g N_Y_M1015_s VNB NSHORT L=0.15 W=0.42 AD=0.1533
+ AS=0.0798 PD=1.57 PS=0.8 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75003.7 SB=75000.3
+ A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90005.5 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1 AD=0.1475
+ AS=0.145 PD=1.295 PS=1.29 NRD=1.9503 NRS=0.9653 M=1 R=5.55556 SA=90000.6
+ SB=90005 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1002_d N_A_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.1475
+ AS=0.145 PD=1.295 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.1
+ SB=90004.6 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.6
+ SB=90004.1 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1006_d N_A_M1008_g N_Y_M1008_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.1
+ SB=90003.6 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g N_Y_M1008_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.5
+ SB=90003.1 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1009_d N_A_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90002.7 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1013_d N_A_M1013_g N_Y_M1011_s VPB PHIGHVT L=0.18 W=1 AD=0.17
+ AS=0.145 PD=1.34 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003.5
+ SB=90002.2 A=0.18 P=2.36 MULT=1
MM1014 N_VPWR_M1013_d N_A_M1014_g N_Y_M1014_s VPB PHIGHVT L=0.18 W=1 AD=0.17
+ AS=0.17 PD=1.34 PS=1.34 NRD=10.8153 NRS=0.9653 M=1 R=5.55556 SA=90004
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1016 N_VPWR_M1016_d N_A_M1016_g N_Y_M1014_s VPB PHIGHVT L=0.18 W=1 AD=0.17
+ AS=0.17 PD=1.34 PS=1.34 NRD=0.9653 NRS=10.8153 M=1 R=5.55556 SA=90004.5
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1017 N_VPWR_M1016_d N_A_M1017_g N_Y_M1017_s VPB PHIGHVT L=0.18 W=1 AD=0.17
+ AS=0.145 PD=1.34 PS=1.29 NRD=10.8153 NRS=0.9653 M=1 R=5.55556 SA=90005
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1018_d N_A_M1018_g N_Y_M1017_s VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90005.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.9461 P=16.85
pX21_noxref noxref_7 A A PROBETYPE=1
pX22_noxref noxref_8 A A PROBETYPE=1
pX23_noxref noxref_9 A A PROBETYPE=1
pX24_noxref noxref_10 A A PROBETYPE=1
pX25_noxref noxref_11 A A PROBETYPE=1
*
.include "sky130_fd_sc_hdll__clkinv_8.pxi.spice"
*
.ends
*
*
