* File: sky130_fd_sc_hdll__and3_2.pxi.spice
* Created: Wed Sep  2 08:22:18 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND3_2%A N_A_c_54_n N_A_M1009_g N_A_M1008_g A
+ PM_SKY130_FD_SC_HDLL__AND3_2%A
x_PM_SKY130_FD_SC_HDLL__AND3_2%B N_B_c_80_n N_B_M1004_g N_B_c_83_n N_B_M1003_g B
+ B PM_SKY130_FD_SC_HDLL__AND3_2%B
x_PM_SKY130_FD_SC_HDLL__AND3_2%C N_C_M1001_g N_C_c_125_n N_C_M1002_g C C
+ PM_SKY130_FD_SC_HDLL__AND3_2%C
x_PM_SKY130_FD_SC_HDLL__AND3_2%A_29_311# N_A_29_311#_M1008_s N_A_29_311#_M1009_s
+ N_A_29_311#_M1003_d N_A_29_311#_c_175_n N_A_29_311#_M1005_g
+ N_A_29_311#_c_169_n N_A_29_311#_M1000_g N_A_29_311#_c_176_n
+ N_A_29_311#_M1007_g N_A_29_311#_c_170_n N_A_29_311#_M1006_g
+ N_A_29_311#_c_177_n N_A_29_311#_c_171_n N_A_29_311#_c_178_n
+ N_A_29_311#_c_179_n N_A_29_311#_c_172_n N_A_29_311#_c_181_n
+ N_A_29_311#_c_182_n N_A_29_311#_c_173_n N_A_29_311#_c_205_n
+ N_A_29_311#_c_184_n N_A_29_311#_c_174_n PM_SKY130_FD_SC_HDLL__AND3_2%A_29_311#
x_PM_SKY130_FD_SC_HDLL__AND3_2%VPWR N_VPWR_M1009_d N_VPWR_M1002_d N_VPWR_M1007_d
+ N_VPWR_c_275_n N_VPWR_c_276_n N_VPWR_c_277_n N_VPWR_c_278_n N_VPWR_c_285_n
+ N_VPWR_c_279_n N_VPWR_c_280_n VPWR N_VPWR_c_281_n N_VPWR_c_282_n
+ N_VPWR_c_274_n PM_SKY130_FD_SC_HDLL__AND3_2%VPWR
x_PM_SKY130_FD_SC_HDLL__AND3_2%X N_X_M1000_s N_X_M1005_s X X X N_X_c_345_n
+ N_X_c_332_n N_X_c_330_n PM_SKY130_FD_SC_HDLL__AND3_2%X
x_PM_SKY130_FD_SC_HDLL__AND3_2%VGND N_VGND_M1001_d N_VGND_M1006_d N_VGND_c_362_n
+ N_VGND_c_363_n N_VGND_c_364_n VGND N_VGND_c_365_n N_VGND_c_366_n
+ N_VGND_c_367_n N_VGND_c_368_n PM_SKY130_FD_SC_HDLL__AND3_2%VGND
cc_1 VNB N_A_c_54_n 0.0401015f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.48
cc_2 VNB N_A_M1008_g 0.0336848f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=0.475
cc_3 VNB A 0.0231074f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_4 VNB N_B_c_80_n 0.00733474f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.48
cc_5 VNB N_B_M1004_g 0.0370767f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.765
cc_6 VNB N_C_M1001_g 0.0285975f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.765
cc_7 VNB N_C_c_125_n 0.0244902f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=0.475
cc_8 VNB C 0.0119268f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_9 VNB C 4.23731e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_29_311#_c_169_n 0.0193135f $X=-0.19 $Y=-0.24 $X2=0.277 $Y2=0.85
cc_11 VNB N_A_29_311#_c_170_n 0.0210624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_29_311#_c_171_n 0.011913f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_29_311#_c_172_n 0.00434876f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_29_311#_c_173_n 0.00896058f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_29_311#_c_174_n 0.047328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_274_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB X 0.0246541f $X=-0.19 $Y=-0.24 $X2=0.277 $Y2=0.85
cc_18 VNB N_X_c_330_n 7.1556e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_362_n 0.00603992f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_363_n 0.0154652f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_21 VNB N_VGND_c_364_n 0.026561f $X=-0.19 $Y=-0.24 $X2=0.277 $Y2=0.85
cc_22 VNB N_VGND_c_365_n 0.039942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_366_n 0.0236077f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_367_n 0.0063175f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_368_n 0.196608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VPB N_A_c_54_n 0.0425098f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.48
cc_27 VPB N_B_c_80_n 0.0117634f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.48
cc_28 VPB N_B_c_83_n 0.0508101f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=0.475
cc_29 VPB N_B_M1003_g 0.011983f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_30 VPB B 0.0110007f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_C_c_125_n 0.0279489f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=0.475
cc_32 VPB N_A_29_311#_c_175_n 0.0186937f $X=-0.19 $Y=1.305 $X2=0.375 $Y2=1.16
cc_33 VPB N_A_29_311#_c_176_n 0.0192434f $X=-0.19 $Y=1.305 $X2=0.277 $Y2=1.16
cc_34 VPB N_A_29_311#_c_177_n 0.0141199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_29_311#_c_178_n 0.00305118f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_29_311#_c_179_n 0.00925693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_29_311#_c_172_n 0.0011162f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_29_311#_c_181_n 0.00118319f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_29_311#_c_182_n 0.0066042f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_29_311#_c_173_n 0.0012199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_29_311#_c_184_n 0.00181824f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_29_311#_c_174_n 0.0261263f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_275_n 0.00149543f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_44 VPB N_VPWR_c_276_n 0.00498307f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_277_n 0.0125989f $X=-0.19 $Y=1.305 $X2=0.277 $Y2=1.16
cc_46 VPB N_VPWR_c_278_n 0.0398159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_279_n 0.0242641f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_280_n 0.00410958f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_281_n 0.0232274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_282_n 0.053359f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_274_n 0.0539998f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB X 0.0151099f $X=-0.19 $Y=1.305 $X2=0.277 $Y2=0.85
cc_53 VPB N_X_c_332_n 0.00168378f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 N_A_c_54_n N_B_c_80_n 0.0463348f $X=0.505 $Y=1.48 $X2=-0.19 $Y2=-0.24
cc_55 N_A_M1008_g N_B_M1004_g 0.0370925f $X=0.535 $Y=0.475 $X2=0 $Y2=0
cc_56 A N_B_M1004_g 3.9475e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_57 N_A_c_54_n N_B_c_83_n 8.20678e-19 $X=0.505 $Y=1.48 $X2=0 $Y2=0
cc_58 N_A_c_54_n N_B_M1003_g 0.0125066f $X=0.505 $Y=1.48 $X2=0 $Y2=0
cc_59 N_A_c_54_n N_A_29_311#_c_177_n 0.00434893f $X=0.505 $Y=1.48 $X2=0 $Y2=0
cc_60 N_A_c_54_n N_A_29_311#_c_171_n 0.00128145f $X=0.505 $Y=1.48 $X2=0 $Y2=0
cc_61 N_A_M1008_g N_A_29_311#_c_171_n 0.0142536f $X=0.535 $Y=0.475 $X2=0 $Y2=0
cc_62 A N_A_29_311#_c_171_n 0.02408f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_63 N_A_c_54_n N_A_29_311#_c_178_n 0.0197968f $X=0.505 $Y=1.48 $X2=0 $Y2=0
cc_64 A N_A_29_311#_c_178_n 0.00820785f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_65 N_A_c_54_n N_A_29_311#_c_179_n 0.00543798f $X=0.505 $Y=1.48 $X2=0 $Y2=0
cc_66 A N_A_29_311#_c_179_n 0.0210059f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_67 N_A_c_54_n N_A_29_311#_c_172_n 0.00229932f $X=0.505 $Y=1.48 $X2=0 $Y2=0
cc_68 N_A_M1008_g N_A_29_311#_c_172_n 0.00977176f $X=0.535 $Y=0.475 $X2=0 $Y2=0
cc_69 A N_A_29_311#_c_172_n 0.030481f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_70 N_A_c_54_n N_VPWR_c_275_n 0.0107103f $X=0.505 $Y=1.48 $X2=0 $Y2=0
cc_71 N_A_c_54_n N_VPWR_c_285_n 0.00389701f $X=0.505 $Y=1.48 $X2=0 $Y2=0
cc_72 N_A_c_54_n N_VPWR_c_282_n 0.00448433f $X=0.505 $Y=1.48 $X2=0 $Y2=0
cc_73 N_A_M1008_g N_VGND_c_365_n 0.00347765f $X=0.535 $Y=0.475 $X2=0 $Y2=0
cc_74 N_A_M1008_g N_VGND_c_368_n 0.00567931f $X=0.535 $Y=0.475 $X2=0 $Y2=0
cc_75 A N_VGND_c_368_n 0.00156165f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_76 N_B_M1004_g N_C_M1001_g 0.0418265f $X=0.895 $Y=0.475 $X2=0 $Y2=0
cc_77 N_B_c_80_n N_C_c_125_n 0.0217479f $X=0.895 $Y=1.26 $X2=0 $Y2=0
cc_78 B N_C_c_125_n 0.00352515f $X=1.165 $Y=2.125 $X2=0 $Y2=0
cc_79 N_B_M1004_g C 0.00682912f $X=0.895 $Y=0.475 $X2=0 $Y2=0
cc_80 N_B_M1004_g N_A_29_311#_c_171_n 0.0067345f $X=0.895 $Y=0.475 $X2=0 $Y2=0
cc_81 N_B_c_80_n N_A_29_311#_c_172_n 0.00464789f $X=0.895 $Y=1.26 $X2=0 $Y2=0
cc_82 N_B_M1004_g N_A_29_311#_c_172_n 0.0129984f $X=0.895 $Y=0.475 $X2=0 $Y2=0
cc_83 N_B_c_80_n N_A_29_311#_c_181_n 0.008218f $X=0.895 $Y=1.26 $X2=0 $Y2=0
cc_84 N_B_c_83_n N_A_29_311#_c_181_n 4.03637e-19 $X=0.975 $Y=2.105 $X2=0 $Y2=0
cc_85 N_B_M1003_g N_A_29_311#_c_181_n 0.00765442f $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_86 B N_A_29_311#_c_181_n 0.00643772f $X=1.165 $Y=2.125 $X2=0 $Y2=0
cc_87 B N_A_29_311#_c_182_n 0.00128683f $X=1.165 $Y=2.125 $X2=0 $Y2=0
cc_88 N_B_c_80_n N_A_29_311#_c_205_n 0.00193228f $X=0.895 $Y=1.26 $X2=0 $Y2=0
cc_89 N_B_M1003_g N_A_29_311#_c_205_n 0.00162596f $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_90 N_B_c_80_n N_A_29_311#_c_184_n 2.58056e-19 $X=0.895 $Y=1.26 $X2=0 $Y2=0
cc_91 N_B_c_83_n N_A_29_311#_c_184_n 2.414e-19 $X=0.975 $Y=2.105 $X2=0 $Y2=0
cc_92 N_B_M1003_g N_A_29_311#_c_184_n 0.00552106f $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_93 B N_A_29_311#_c_184_n 0.0168986f $X=1.165 $Y=2.125 $X2=0 $Y2=0
cc_94 N_B_c_83_n N_VPWR_c_275_n 6.57524e-19 $X=0.975 $Y=2.105 $X2=0 $Y2=0
cc_95 N_B_M1003_g N_VPWR_c_275_n 0.0034845f $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_96 N_B_c_83_n N_VPWR_c_276_n 0.00248857f $X=0.975 $Y=2.105 $X2=0 $Y2=0
cc_97 N_B_M1003_g N_VPWR_c_276_n 0.0018025f $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_98 B N_VPWR_c_276_n 0.0264701f $X=1.165 $Y=2.125 $X2=0 $Y2=0
cc_99 N_B_c_80_n N_VPWR_c_285_n 2.16256e-19 $X=0.895 $Y=1.26 $X2=0 $Y2=0
cc_100 N_B_M1003_g N_VPWR_c_285_n 0.0035719f $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_101 N_B_c_83_n N_VPWR_c_279_n 0.00720942f $X=0.975 $Y=2.105 $X2=0 $Y2=0
cc_102 B N_VPWR_c_279_n 0.0380394f $X=1.165 $Y=2.125 $X2=0 $Y2=0
cc_103 N_B_c_83_n N_VPWR_c_282_n 0.00989316f $X=0.975 $Y=2.105 $X2=0 $Y2=0
cc_104 B N_VPWR_c_282_n 0.028168f $X=1.165 $Y=2.125 $X2=0 $Y2=0
cc_105 N_B_c_83_n N_VPWR_c_274_n 0.0101872f $X=0.975 $Y=2.105 $X2=0 $Y2=0
cc_106 B N_VPWR_c_274_n 0.020518f $X=1.165 $Y=2.125 $X2=0 $Y2=0
cc_107 N_B_M1004_g N_VGND_c_365_n 0.00451413f $X=0.895 $Y=0.475 $X2=0 $Y2=0
cc_108 N_B_M1004_g N_VGND_c_368_n 0.00771524f $X=0.895 $Y=0.475 $X2=0 $Y2=0
cc_109 N_C_c_125_n N_A_29_311#_c_175_n 0.0145349f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_110 N_C_M1001_g N_A_29_311#_c_169_n 0.0132891f $X=1.35 $Y=0.475 $X2=0 $Y2=0
cc_111 C N_A_29_311#_c_169_n 0.00263331f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_112 C N_A_29_311#_c_169_n 6.12055e-19 $X=1.08 $Y=0.425 $X2=0 $Y2=0
cc_113 N_C_M1001_g N_A_29_311#_c_171_n 2.18102e-19 $X=1.35 $Y=0.475 $X2=0 $Y2=0
cc_114 C N_A_29_311#_c_171_n 0.0214033f $X=1.08 $Y=0.425 $X2=0 $Y2=0
cc_115 N_C_M1001_g N_A_29_311#_c_172_n 5.60035e-19 $X=1.35 $Y=0.475 $X2=0 $Y2=0
cc_116 N_C_c_125_n N_A_29_311#_c_172_n 8.64293e-19 $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_117 C N_A_29_311#_c_172_n 0.0527966f $X=1.08 $Y=0.425 $X2=0 $Y2=0
cc_118 C N_A_29_311#_c_181_n 0.00924599f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_119 N_C_c_125_n N_A_29_311#_c_182_n 0.0105391f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_120 C N_A_29_311#_c_182_n 0.0103913f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_121 N_C_c_125_n N_A_29_311#_c_173_n 0.00458955f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_122 C N_A_29_311#_c_173_n 0.0198994f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_123 N_C_c_125_n N_A_29_311#_c_184_n 0.0145232f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_124 C N_A_29_311#_c_184_n 0.0245131f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_125 N_C_c_125_n N_A_29_311#_c_174_n 0.0240078f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_126 C N_A_29_311#_c_174_n 9.05841e-19 $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_127 N_C_c_125_n N_VPWR_c_276_n 0.00435022f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_128 N_C_c_125_n N_VPWR_c_285_n 2.56837e-19 $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_129 N_C_c_125_n N_VPWR_c_279_n 0.00159425f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_130 N_C_c_125_n N_VPWR_c_274_n 0.00194828f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_131 N_C_M1001_g X 5.61276e-19 $X=1.35 $Y=0.475 $X2=0 $Y2=0
cc_132 C X 0.00322662f $X=1.08 $Y=0.425 $X2=0 $Y2=0
cc_133 C N_X_c_330_n 0.00804073f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_134 C A_194_53# 0.0052042f $X=1.08 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_135 N_C_M1001_g N_VGND_c_362_n 0.00741778f $X=1.35 $Y=0.475 $X2=0 $Y2=0
cc_136 N_C_c_125_n N_VGND_c_362_n 5.58019e-19 $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_137 C N_VGND_c_362_n 0.0119552f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_138 C N_VGND_c_362_n 0.0209169f $X=1.08 $Y=0.425 $X2=0 $Y2=0
cc_139 N_C_M1001_g N_VGND_c_365_n 0.0039881f $X=1.35 $Y=0.475 $X2=0 $Y2=0
cc_140 C N_VGND_c_365_n 0.0024496f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_141 C N_VGND_c_365_n 0.0116437f $X=1.08 $Y=0.425 $X2=0 $Y2=0
cc_142 N_C_M1001_g N_VGND_c_368_n 0.0060562f $X=1.35 $Y=0.475 $X2=0 $Y2=0
cc_143 C N_VGND_c_368_n 0.00466102f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_144 C N_VGND_c_368_n 0.00912818f $X=1.08 $Y=0.425 $X2=0 $Y2=0
cc_145 N_A_29_311#_c_178_n N_VPWR_M1009_d 3.94276e-19 $X=0.69 $Y=1.51 $X2=-0.19
+ $Y2=-0.24
cc_146 N_A_29_311#_c_205_n N_VPWR_M1009_d 0.0015309f $X=0.792 $Y=1.51 $X2=-0.19
+ $Y2=-0.24
cc_147 N_A_29_311#_c_182_n N_VPWR_M1002_d 0.00442957f $X=1.81 $Y=1.51 $X2=0
+ $Y2=0
cc_148 N_A_29_311#_c_177_n N_VPWR_c_275_n 3.71611e-19 $X=0.27 $Y=1.76 $X2=0
+ $Y2=0
cc_149 N_A_29_311#_c_175_n N_VPWR_c_276_n 0.00462168f $X=2.045 $Y=1.41 $X2=0
+ $Y2=0
cc_150 N_A_29_311#_c_182_n N_VPWR_c_276_n 0.0146982f $X=1.81 $Y=1.51 $X2=0 $Y2=0
cc_151 N_A_29_311#_c_184_n N_VPWR_c_276_n 0.00601324f $X=1.33 $Y=1.51 $X2=0
+ $Y2=0
cc_152 N_A_29_311#_c_174_n N_VPWR_c_276_n 3.95938e-19 $X=2.515 $Y=1.202 $X2=0
+ $Y2=0
cc_153 N_A_29_311#_c_176_n N_VPWR_c_278_n 0.0101772f $X=2.515 $Y=1.41 $X2=0
+ $Y2=0
cc_154 N_A_29_311#_c_177_n N_VPWR_c_285_n 0.0145346f $X=0.27 $Y=1.76 $X2=0 $Y2=0
cc_155 N_A_29_311#_c_178_n N_VPWR_c_285_n 0.00749807f $X=0.69 $Y=1.51 $X2=0
+ $Y2=0
cc_156 N_A_29_311#_c_181_n N_VPWR_c_285_n 6.49764e-19 $X=1.18 $Y=1.51 $X2=0
+ $Y2=0
cc_157 N_A_29_311#_c_205_n N_VPWR_c_285_n 0.0120451f $X=0.792 $Y=1.51 $X2=0
+ $Y2=0
cc_158 N_A_29_311#_c_184_n N_VPWR_c_285_n 0.00669846f $X=1.33 $Y=1.51 $X2=0
+ $Y2=0
cc_159 N_A_29_311#_c_175_n N_VPWR_c_281_n 0.00702461f $X=2.045 $Y=1.41 $X2=0
+ $Y2=0
cc_160 N_A_29_311#_c_176_n N_VPWR_c_281_n 0.00429201f $X=2.515 $Y=1.41 $X2=0
+ $Y2=0
cc_161 N_A_29_311#_c_177_n N_VPWR_c_282_n 0.0222117f $X=0.27 $Y=1.76 $X2=0 $Y2=0
cc_162 N_A_29_311#_c_178_n N_VPWR_c_282_n 0.00498695f $X=0.69 $Y=1.51 $X2=0
+ $Y2=0
cc_163 N_A_29_311#_c_175_n N_VPWR_c_274_n 0.0137292f $X=2.045 $Y=1.41 $X2=0
+ $Y2=0
cc_164 N_A_29_311#_c_176_n N_VPWR_c_274_n 0.00716187f $X=2.515 $Y=1.41 $X2=0
+ $Y2=0
cc_165 N_A_29_311#_c_177_n N_VPWR_c_274_n 0.00100952f $X=0.27 $Y=1.76 $X2=0
+ $Y2=0
cc_166 N_A_29_311#_c_169_n X 0.0174424f $X=2.055 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_29_311#_c_173_n X 0.00288489f $X=1.955 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A_29_311#_c_174_n X 0.0014966f $X=2.515 $Y=1.202 $X2=0 $Y2=0
cc_169 N_A_29_311#_c_175_n X 0.0063111f $X=2.045 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_29_311#_c_176_n X 0.00154202f $X=2.515 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_29_311#_c_170_n X 0.01085f $X=2.545 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_29_311#_c_182_n X 0.0115101f $X=1.81 $Y=1.51 $X2=0 $Y2=0
cc_173 N_A_29_311#_c_173_n X 0.0274396f $X=1.955 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_29_311#_c_174_n X 0.0351377f $X=2.515 $Y=1.202 $X2=0 $Y2=0
cc_175 N_A_29_311#_c_176_n N_X_c_345_n 0.0222707f $X=2.515 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A_29_311#_c_174_n N_X_c_345_n 0.0026358f $X=2.515 $Y=1.202 $X2=0 $Y2=0
cc_177 N_A_29_311#_c_176_n N_X_c_332_n 0.0133498f $X=2.515 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A_29_311#_c_169_n N_X_c_330_n 0.00375326f $X=2.055 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_29_311#_c_170_n N_X_c_330_n 0.00420201f $X=2.545 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_29_311#_c_171_n A_122_53# 0.00191292f $X=0.69 $Y=0.437 $X2=-0.19
+ $Y2=-0.24
cc_181 N_A_29_311#_c_172_n A_122_53# 0.0012908f $X=0.792 $Y=1.425 $X2=-0.19
+ $Y2=-0.24
cc_182 N_A_29_311#_c_169_n N_VGND_c_362_n 0.00612553f $X=2.055 $Y=0.995 $X2=0
+ $Y2=0
cc_183 N_A_29_311#_c_170_n N_VGND_c_364_n 0.00911137f $X=2.545 $Y=0.995 $X2=0
+ $Y2=0
cc_184 N_A_29_311#_c_171_n N_VGND_c_365_n 0.0354833f $X=0.69 $Y=0.437 $X2=0
+ $Y2=0
cc_185 N_A_29_311#_c_169_n N_VGND_c_366_n 0.00366776f $X=2.055 $Y=0.995 $X2=0
+ $Y2=0
cc_186 N_A_29_311#_c_170_n N_VGND_c_366_n 0.00585385f $X=2.545 $Y=0.995 $X2=0
+ $Y2=0
cc_187 N_A_29_311#_c_169_n N_VGND_c_368_n 0.00643925f $X=2.055 $Y=0.995 $X2=0
+ $Y2=0
cc_188 N_A_29_311#_c_170_n N_VGND_c_368_n 0.012076f $X=2.545 $Y=0.995 $X2=0
+ $Y2=0
cc_189 N_A_29_311#_c_171_n N_VGND_c_368_n 0.027991f $X=0.69 $Y=0.437 $X2=0 $Y2=0
cc_190 N_VPWR_c_274_n N_X_M1005_s 0.00352766f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_191 N_VPWR_c_278_n X 0.0114887f $X=2.875 $Y=1.96 $X2=0 $Y2=0
cc_192 N_VPWR_c_281_n N_X_c_345_n 0.0278752f $X=2.79 $Y=2.72 $X2=0 $Y2=0
cc_193 N_VPWR_c_274_n N_X_c_345_n 0.0163563f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_194 X N_VGND_c_362_n 0.0257991f $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_195 X N_VGND_c_364_n 0.0197021f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_196 X N_VGND_c_366_n 0.0278854f $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_197 N_X_M1000_s N_VGND_c_368_n 0.00415351f $X=2.13 $Y=0.235 $X2=0 $Y2=0
cc_198 X N_VGND_c_368_n 0.016298f $X=2.01 $Y=0.425 $X2=0 $Y2=0
