* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 a_255_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.45e+11p pd=2.49e+06u as=9.7e+11p ps=7.94e+06u
M1001 a_245_47# B1 a_151_47# VNB nshort w=650000u l=150000u
+  ad=3.9325e+11p pd=3.81e+06u as=3.9975e+11p ps=3.83e+06u
M1002 a_151_47# C1 a_38_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.6975e+11p ps=2.13e+06u
M1003 a_151_47# B2 a_245_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A1 a_245_47# VNB nshort w=650000u l=150000u
+  ad=5.46e+11p pd=5.58e+06u as=0p ps=0u
M1005 VPWR A1 a_535_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.3e+11p ps=2.46e+06u
M1006 a_535_297# A2 a_38_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.13e+12p ps=6.26e+06u
M1007 VPWR C1 a_38_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_245_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_38_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1010 a_38_47# B2 a_255_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_38_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.405e+11p ps=2.04e+06u
M1012 X a_38_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_38_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
