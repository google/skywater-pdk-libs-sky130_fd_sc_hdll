* File: sky130_fd_sc_hdll__bufinv_16.pxi.spice
* Created: Thu Aug 27 19:01:07 2020
* 
x_PM_SKY130_FD_SC_HDLL__BUFINV_16%A N_A_M1014_g N_A_c_211_n N_A_M1001_g
+ N_A_M1042_g N_A_c_212_n N_A_M1019_g N_A_c_213_n N_A_M1041_g N_A_M1049_g A
+ N_A_c_209_n N_A_c_210_n PM_SKY130_FD_SC_HDLL__BUFINV_16%A
x_PM_SKY130_FD_SC_HDLL__BUFINV_16%A_27_47# N_A_27_47#_M1014_d N_A_27_47#_M1042_d
+ N_A_27_47#_M1001_d N_A_27_47#_M1019_d N_A_27_47#_M1021_g N_A_27_47#_c_291_n
+ N_A_27_47#_M1000_g N_A_27_47#_M1024_g N_A_27_47#_c_292_n N_A_27_47#_M1005_g
+ N_A_27_47#_M1036_g N_A_27_47#_c_293_n N_A_27_47#_M1013_g N_A_27_47#_M1040_g
+ N_A_27_47#_c_294_n N_A_27_47#_M1023_g N_A_27_47#_M1043_g N_A_27_47#_c_295_n
+ N_A_27_47#_M1030_g N_A_27_47#_c_296_n N_A_27_47#_M1035_g N_A_27_47#_M1048_g
+ N_A_27_47#_c_281_n N_A_27_47#_c_297_n N_A_27_47#_c_282_n N_A_27_47#_c_283_n
+ N_A_27_47#_c_298_n N_A_27_47#_c_299_n N_A_27_47#_c_323_n N_A_27_47#_c_325_n
+ N_A_27_47#_c_284_n N_A_27_47#_c_300_n N_A_27_47#_c_285_n N_A_27_47#_c_286_n
+ N_A_27_47#_c_287_n N_A_27_47#_c_288_n N_A_27_47#_c_302_n N_A_27_47#_c_289_n
+ N_A_27_47#_c_290_n PM_SKY130_FD_SC_HDLL__BUFINV_16%A_27_47#
x_PM_SKY130_FD_SC_HDLL__BUFINV_16%A_391_47# N_A_391_47#_M1021_d
+ N_A_391_47#_M1036_d N_A_391_47#_M1043_d N_A_391_47#_M1000_d
+ N_A_391_47#_M1013_d N_A_391_47#_M1030_d N_A_391_47#_M1004_g
+ N_A_391_47#_c_510_n N_A_391_47#_M1002_g N_A_391_47#_M1007_g
+ N_A_391_47#_c_511_n N_A_391_47#_M1003_g N_A_391_47#_M1008_g
+ N_A_391_47#_c_512_n N_A_391_47#_M1006_g N_A_391_47#_M1009_g
+ N_A_391_47#_c_513_n N_A_391_47#_M1010_g N_A_391_47#_M1012_g
+ N_A_391_47#_c_514_n N_A_391_47#_M1011_g N_A_391_47#_M1016_g
+ N_A_391_47#_c_515_n N_A_391_47#_M1015_g N_A_391_47#_M1018_g
+ N_A_391_47#_c_516_n N_A_391_47#_M1017_g N_A_391_47#_M1022_g
+ N_A_391_47#_c_517_n N_A_391_47#_M1020_g N_A_391_47#_M1025_g
+ N_A_391_47#_c_518_n N_A_391_47#_M1027_g N_A_391_47#_M1026_g
+ N_A_391_47#_c_519_n N_A_391_47#_M1028_g N_A_391_47#_M1029_g
+ N_A_391_47#_c_520_n N_A_391_47#_M1032_g N_A_391_47#_M1031_g
+ N_A_391_47#_c_521_n N_A_391_47#_M1033_g N_A_391_47#_M1034_g
+ N_A_391_47#_c_522_n N_A_391_47#_M1038_g N_A_391_47#_M1037_g
+ N_A_391_47#_c_523_n N_A_391_47#_M1039_g N_A_391_47#_M1044_g
+ N_A_391_47#_c_524_n N_A_391_47#_M1046_g N_A_391_47#_c_525_n
+ N_A_391_47#_M1047_g N_A_391_47#_M1045_g N_A_391_47#_c_534_n
+ N_A_391_47#_c_535_n N_A_391_47#_c_499_n N_A_391_47#_c_500_n
+ N_A_391_47#_c_526_n N_A_391_47#_c_527_n N_A_391_47#_c_563_n
+ N_A_391_47#_c_567_n N_A_391_47#_c_501_n N_A_391_47#_c_528_n
+ N_A_391_47#_c_579_n N_A_391_47#_c_581_n N_A_391_47#_c_502_n
+ N_A_391_47#_c_529_n N_A_391_47#_c_503_n N_A_391_47#_c_504_n
+ N_A_391_47#_c_505_n N_A_391_47#_c_506_n N_A_391_47#_c_531_n
+ N_A_391_47#_c_507_n N_A_391_47#_c_532_n N_A_391_47#_c_508_n
+ N_A_391_47#_c_509_n PM_SKY130_FD_SC_HDLL__BUFINV_16%A_391_47#
x_PM_SKY130_FD_SC_HDLL__BUFINV_16%VPWR N_VPWR_M1001_s N_VPWR_M1041_s
+ N_VPWR_M1005_s N_VPWR_M1023_s N_VPWR_M1035_s N_VPWR_M1003_s N_VPWR_M1010_s
+ N_VPWR_M1015_s N_VPWR_M1020_s N_VPWR_M1028_s N_VPWR_M1033_s N_VPWR_M1039_s
+ N_VPWR_M1047_s N_VPWR_c_946_n N_VPWR_c_947_n N_VPWR_c_948_n N_VPWR_c_949_n
+ N_VPWR_c_950_n N_VPWR_c_951_n N_VPWR_c_952_n N_VPWR_c_953_n N_VPWR_c_954_n
+ N_VPWR_c_955_n N_VPWR_c_956_n N_VPWR_c_957_n N_VPWR_c_958_n N_VPWR_c_959_n
+ N_VPWR_c_960_n N_VPWR_c_961_n N_VPWR_c_962_n N_VPWR_c_963_n N_VPWR_c_964_n
+ N_VPWR_c_965_n N_VPWR_c_966_n N_VPWR_c_967_n N_VPWR_c_968_n N_VPWR_c_969_n
+ N_VPWR_c_970_n N_VPWR_c_971_n N_VPWR_c_972_n N_VPWR_c_973_n N_VPWR_c_974_n
+ N_VPWR_c_975_n N_VPWR_c_976_n N_VPWR_c_977_n N_VPWR_c_978_n N_VPWR_c_979_n
+ N_VPWR_c_980_n VPWR N_VPWR_c_981_n N_VPWR_c_945_n N_VPWR_c_983_n
+ N_VPWR_c_984_n N_VPWR_c_985_n VPWR PM_SKY130_FD_SC_HDLL__BUFINV_16%VPWR
x_PM_SKY130_FD_SC_HDLL__BUFINV_16%Y N_Y_M1004_s N_Y_M1008_s N_Y_M1012_s
+ N_Y_M1018_s N_Y_M1025_s N_Y_M1029_s N_Y_M1034_s N_Y_M1044_s N_Y_M1002_d
+ N_Y_M1006_d N_Y_M1011_d N_Y_M1017_d N_Y_M1027_d N_Y_M1032_d N_Y_M1038_d
+ N_Y_M1046_d N_Y_c_1189_n N_Y_c_1187_n N_Y_c_1188_n N_Y_c_1152_n N_Y_c_1153_n
+ N_Y_c_1169_n N_Y_c_1170_n N_Y_c_1216_n N_Y_c_1218_n N_Y_c_1222_n N_Y_c_1154_n
+ N_Y_c_1171_n N_Y_c_1234_n N_Y_c_1236_n N_Y_c_1240_n N_Y_c_1155_n N_Y_c_1172_n
+ N_Y_c_1252_n N_Y_c_1256_n N_Y_c_1156_n N_Y_c_1173_n N_Y_c_1268_n N_Y_c_1272_n
+ N_Y_c_1157_n N_Y_c_1174_n N_Y_c_1284_n N_Y_c_1288_n N_Y_c_1158_n N_Y_c_1175_n
+ N_Y_c_1300_n N_Y_c_1304_n N_Y_c_1159_n N_Y_c_1176_n N_Y_c_1316_n N_Y_c_1318_n
+ N_Y_c_1160_n N_Y_c_1177_n N_Y_c_1161_n N_Y_c_1178_n N_Y_c_1162_n N_Y_c_1179_n
+ N_Y_c_1163_n N_Y_c_1180_n N_Y_c_1164_n N_Y_c_1181_n N_Y_c_1165_n N_Y_c_1182_n
+ N_Y_c_1166_n N_Y_c_1183_n N_Y_c_1167_n N_Y_c_1184_n Y Y
+ PM_SKY130_FD_SC_HDLL__BUFINV_16%Y
x_PM_SKY130_FD_SC_HDLL__BUFINV_16%VGND N_VGND_M1014_s N_VGND_M1049_s
+ N_VGND_M1024_s N_VGND_M1040_s N_VGND_M1048_s N_VGND_M1007_d N_VGND_M1009_d
+ N_VGND_M1016_d N_VGND_M1022_d N_VGND_M1026_d N_VGND_M1031_d N_VGND_M1037_d
+ N_VGND_M1045_d N_VGND_c_1515_n N_VGND_c_1516_n N_VGND_c_1517_n N_VGND_c_1518_n
+ N_VGND_c_1519_n N_VGND_c_1520_n N_VGND_c_1521_n N_VGND_c_1522_n
+ N_VGND_c_1523_n N_VGND_c_1524_n N_VGND_c_1525_n N_VGND_c_1526_n
+ N_VGND_c_1527_n N_VGND_c_1528_n N_VGND_c_1529_n N_VGND_c_1530_n
+ N_VGND_c_1531_n N_VGND_c_1532_n N_VGND_c_1533_n N_VGND_c_1534_n
+ N_VGND_c_1535_n N_VGND_c_1536_n N_VGND_c_1537_n N_VGND_c_1538_n
+ N_VGND_c_1539_n N_VGND_c_1540_n N_VGND_c_1541_n N_VGND_c_1542_n
+ N_VGND_c_1543_n N_VGND_c_1544_n N_VGND_c_1545_n N_VGND_c_1546_n
+ N_VGND_c_1547_n N_VGND_c_1548_n N_VGND_c_1549_n VGND N_VGND_c_1550_n
+ N_VGND_c_1551_n N_VGND_c_1552_n N_VGND_c_1553_n N_VGND_c_1554_n VGND
+ PM_SKY130_FD_SC_HDLL__BUFINV_16%VGND
cc_1 VNB N_A_M1014_g 0.0244194f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_A_M1042_g 0.0188756f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_3 VNB N_A_M1049_g 0.0185511f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_4 VNB N_A_c_209_n 0.0148466f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.16
cc_5 VNB N_A_c_210_n 0.070276f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.217
cc_6 VNB N_A_27_47#_M1021_g 0.0181991f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_7 VNB N_A_27_47#_M1024_g 0.0183796f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_8 VNB N_A_27_47#_M1036_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.16
cc_9 VNB N_A_27_47#_M1040_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.175
cc_10 VNB N_A_27_47#_M1043_g 0.0188753f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_M1048_g 0.0185509f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_281_n 0.0186353f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_282_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_283_n 0.0100396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_284_n 0.00102469f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_285_n 0.00304777f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_286_n 5.26104e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_287_n 0.00343466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_288_n 0.00263423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_289_n 0.00153756f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_290_n 0.13593f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_391_47#_M1004_g 0.0181991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_391_47#_M1007_g 0.0183796f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.217
cc_24 VNB N_A_391_47#_M1008_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_391_47#_M1009_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_391_47#_M1012_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_391_47#_M1016_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_391_47#_M1018_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_391_47#_M1022_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_391_47#_M1025_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_391_47#_M1026_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_391_47#_M1029_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_391_47#_M1031_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_391_47#_M1034_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_391_47#_M1037_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_391_47#_M1044_g 0.0188758f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_391_47#_M1045_g 0.0218157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_391_47#_c_499_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_391_47#_c_500_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_391_47#_c_501_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_391_47#_c_502_n 9.58484e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_391_47#_c_503_n 0.00305698f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_391_47#_c_504_n 5.27693e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_391_47#_c_505_n 0.00343466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_391_47#_c_506_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_391_47#_c_507_n 0.00278347f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_391_47#_c_508_n 0.00163661f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_391_47#_c_509_n 0.376438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VPWR_c_945_n 0.516438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_Y_c_1152_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_Y_c_1153_n 0.00253087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_Y_c_1154_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_Y_c_1155_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_Y_c_1156_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_Y_c_1157_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_Y_c_1158_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_Y_c_1159_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_Y_c_1160_n 0.00938092f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_Y_c_1161_n 0.00253075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_Y_c_1162_n 0.00253075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_Y_c_1163_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_Y_c_1164_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_Y_c_1165_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_Y_c_1166_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_Y_c_1167_n 0.00263423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB Y 0.0207773f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1515_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1516_n 0.0194241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1517_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1518_n 0.0200002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1519_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1520_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1521_n 0.00466605f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1522_n 0.00467908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1523_n 0.00467908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1524_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1525_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1526_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1527_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1528_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1529_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1530_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1531_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1532_n 0.0193874f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1533_n 0.00323954f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1534_n 0.0198969f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1535_n 0.00324139f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1536_n 0.0193636f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1537_n 0.00324139f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1538_n 0.0193636f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1539_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1540_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1541_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1542_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1543_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1544_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1545_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1546_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1547_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1548_n 0.0194241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1549_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1550_n 0.0120879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1551_n 0.567295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1552_n 0.0219871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1553_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1554_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VPB N_A_c_211_n 0.0200897f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_108 VPB N_A_c_212_n 0.0158858f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_109 VPB N_A_c_213_n 0.0159693f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_110 VPB N_A_c_210_n 0.0223834f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.217
cc_111 VPB N_A_27_47#_c_291_n 0.0162292f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_112 VPB N_A_27_47#_c_292_n 0.0158858f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.217
cc_113 VPB N_A_27_47#_c_293_n 0.0158869f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.217
cc_114 VPB N_A_27_47#_c_294_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_27_47#_c_295_n 0.0158857f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_27_47#_c_296_n 0.0159692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_27_47#_c_297_n 0.0331497f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_27_47#_c_298_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_27_47#_c_299_n 0.0101812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_27_47#_c_300_n 0.00100785f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_27_47#_c_286_n 0.00252324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_27_47#_c_302_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_27_47#_c_290_n 0.0384682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_391_47#_c_510_n 0.0162292f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_391_47#_c_511_n 0.0158858f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.16
cc_126 VPB N_A_391_47#_c_512_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_391_47#_c_513_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_391_47#_c_514_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_391_47#_c_515_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_391_47#_c_516_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_391_47#_c_517_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_391_47#_c_518_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_391_47#_c_519_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_391_47#_c_520_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_391_47#_c_521_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_391_47#_c_522_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_391_47#_c_523_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_391_47#_c_524_n 0.0158858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_391_47#_c_525_n 0.0191645f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_391_47#_c_526_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_391_47#_c_527_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_391_47#_c_528_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_391_47#_c_529_n 9.4165e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_391_47#_c_504_n 0.0025308f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_391_47#_c_531_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_391_47#_c_532_n 0.00179747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_391_47#_c_509_n 0.101888f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_946_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_947_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_948_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_949_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_950_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_951_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_952_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_953_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_954_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_955_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_956_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_957_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_958_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_959_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_960_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_961_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_962_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_963_n 0.020564f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_964_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_965_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_966_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_967_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_968_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_969_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_970_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_971_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_972_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_973_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_974_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_975_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_976_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_977_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_978_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_979_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_980_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_981_n 0.0124854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_945_n 0.0528234f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_983_n 0.0226976f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_984_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_985_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_Y_c_1169_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_Y_c_1170_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_Y_c_1171_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_Y_c_1172_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_Y_c_1173_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_Y_c_1174_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_Y_c_1175_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_Y_c_1176_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_Y_c_1177_n 7.91715e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_Y_c_1178_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_Y_c_1179_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_Y_c_1180_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_Y_c_1181_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_Y_c_1182_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_Y_c_1183_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_Y_c_1184_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB Y 0.00722345f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB Y 0.0103072f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 N_A_M1049_g N_A_27_47#_M1021_g 0.0207193f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_207 N_A_c_213_n N_A_27_47#_c_291_n 0.0215651f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A_M1014_g N_A_27_47#_c_281_n 0.00693104f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_209 N_A_M1042_g N_A_27_47#_c_281_n 5.47935e-19 $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_210 N_A_c_211_n N_A_27_47#_c_297_n 0.0112091f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A_c_212_n N_A_27_47#_c_297_n 7.06303e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A_M1014_g N_A_27_47#_c_282_n 0.00879805f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_213 N_A_M1042_g N_A_27_47#_c_282_n 0.00879805f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_214 N_A_c_209_n N_A_27_47#_c_282_n 0.03957f $X=1.07 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A_c_210_n N_A_27_47#_c_282_n 0.0031956f $X=1.435 $Y=1.217 $X2=0 $Y2=0
cc_216 N_A_M1014_g N_A_27_47#_c_283_n 0.00126794f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_217 N_A_c_209_n N_A_27_47#_c_283_n 0.0278128f $X=1.07 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A_c_211_n N_A_27_47#_c_298_n 0.0137916f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_219 N_A_c_212_n N_A_27_47#_c_298_n 0.0101048f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_220 N_A_c_209_n N_A_27_47#_c_298_n 0.0394547f $X=1.07 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A_c_210_n N_A_27_47#_c_298_n 0.00720931f $X=1.435 $Y=1.217 $X2=0 $Y2=0
cc_222 N_A_c_211_n N_A_27_47#_c_299_n 0.00138874f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A_c_209_n N_A_27_47#_c_299_n 0.0279779f $X=1.07 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A_c_210_n N_A_27_47#_c_299_n 3.20658e-19 $X=1.435 $Y=1.217 $X2=0 $Y2=0
cc_225 N_A_M1014_g N_A_27_47#_c_323_n 5.25882e-19 $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_226 N_A_M1042_g N_A_27_47#_c_323_n 0.00657592f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_227 N_A_c_211_n N_A_27_47#_c_325_n 7.33057e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_228 N_A_c_212_n N_A_27_47#_c_325_n 0.0137692f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_229 N_A_c_213_n N_A_27_47#_c_325_n 0.0112091f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_230 N_A_M1049_g N_A_27_47#_c_284_n 0.0116573f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_231 N_A_c_213_n N_A_27_47#_c_300_n 0.0151183f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_232 N_A_c_210_n N_A_27_47#_c_300_n 3.58038e-19 $X=1.435 $Y=1.217 $X2=0 $Y2=0
cc_233 N_A_M1049_g N_A_27_47#_c_285_n 0.00410511f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_234 N_A_c_213_n N_A_27_47#_c_286_n 8.16926e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A_c_210_n N_A_27_47#_c_286_n 0.00327205f $X=1.435 $Y=1.217 $X2=0 $Y2=0
cc_236 N_A_M1042_g N_A_27_47#_c_288_n 0.0011682f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_237 N_A_c_209_n N_A_27_47#_c_288_n 0.0307156f $X=1.07 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A_c_210_n N_A_27_47#_c_288_n 0.00450461f $X=1.435 $Y=1.217 $X2=0 $Y2=0
cc_239 N_A_c_212_n N_A_27_47#_c_302_n 0.00259297f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_240 N_A_c_213_n N_A_27_47#_c_302_n 0.00107777f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_241 N_A_c_209_n N_A_27_47#_c_302_n 0.0305808f $X=1.07 $Y=1.16 $X2=0 $Y2=0
cc_242 N_A_c_210_n N_A_27_47#_c_302_n 0.00723098f $X=1.435 $Y=1.217 $X2=0 $Y2=0
cc_243 N_A_c_209_n N_A_27_47#_c_289_n 0.014524f $X=1.07 $Y=1.16 $X2=0 $Y2=0
cc_244 N_A_c_210_n N_A_27_47#_c_289_n 0.00220849f $X=1.435 $Y=1.217 $X2=0 $Y2=0
cc_245 N_A_c_210_n N_A_27_47#_c_290_n 0.0207193f $X=1.435 $Y=1.217 $X2=0 $Y2=0
cc_246 N_A_M1049_g N_A_391_47#_c_534_n 5.33681e-19 $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_247 N_A_c_213_n N_A_391_47#_c_535_n 7.33057e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_248 N_A_c_211_n N_VPWR_c_946_n 0.00547044f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_249 N_A_c_212_n N_VPWR_c_946_n 0.00497803f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_250 N_A_c_212_n N_VPWR_c_947_n 0.00597712f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_251 N_A_c_213_n N_VPWR_c_947_n 0.00673617f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_252 N_A_c_213_n N_VPWR_c_948_n 0.00547044f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_253 N_A_c_211_n N_VPWR_c_945_n 0.0127552f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_254 N_A_c_212_n N_VPWR_c_945_n 0.00999457f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_255 N_A_c_213_n N_VPWR_c_945_n 0.011869f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_256 N_A_c_211_n N_VPWR_c_983_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_257 N_A_M1014_g N_VGND_c_1515_n 0.00390178f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_258 N_A_M1042_g N_VGND_c_1515_n 0.00276126f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_259 N_A_M1042_g N_VGND_c_1516_n 0.00424619f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_260 N_A_M1049_g N_VGND_c_1516_n 0.00439206f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_261 N_A_M1049_g N_VGND_c_1517_n 0.00268723f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_262 N_A_M1014_g N_VGND_c_1551_n 0.00694018f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_263 N_A_M1042_g N_VGND_c_1551_n 0.00610552f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_264 N_A_M1049_g N_VGND_c_1551_n 0.00618081f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_265 N_A_M1014_g N_VGND_c_1552_n 0.00424619f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_266 N_A_27_47#_M1048_g N_A_391_47#_M1004_g 0.0207158f $X=4.28 $Y=0.56 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_296_n N_A_391_47#_c_510_n 0.0216821f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_M1021_g N_A_391_47#_c_534_n 0.0065059f $X=1.88 $Y=0.56 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_M1024_g N_A_391_47#_c_534_n 0.00693104f $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_M1036_g N_A_391_47#_c_534_n 5.47131e-19 $X=2.82 $Y=0.56 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_291_n N_A_391_47#_c_535_n 0.0137692f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_292_n N_A_391_47#_c_535_n 0.0115459f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_293_n N_A_391_47#_c_535_n 7.68612e-19 $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_325_n N_A_391_47#_c_535_n 0.00486061f $X=1.2 $Y=1.63 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_M1024_g N_A_391_47#_c_499_n 0.00879805f $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_M1036_g N_A_391_47#_c_499_n 0.00879805f $X=2.82 $Y=0.56 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_287_n N_A_391_47#_c_499_n 0.03957f $X=3.91 $Y=1.16 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_290_n N_A_391_47#_c_499_n 0.0031956f $X=4.255 $Y=1.217 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_M1021_g N_A_391_47#_c_500_n 0.00243606f $X=1.88 $Y=0.56 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_M1024_g N_A_391_47#_c_500_n 0.00113891f $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_284_n N_A_391_47#_c_500_n 0.00808484f $X=1.585 $Y=0.82 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_287_n N_A_391_47#_c_500_n 0.030582f $X=3.91 $Y=1.16 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_290_n N_A_391_47#_c_500_n 0.00331919f $X=4.255 $Y=1.217
+ $X2=0 $Y2=0
cc_284 N_A_27_47#_c_292_n N_A_391_47#_c_526_n 0.0137916f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_293_n N_A_391_47#_c_526_n 0.0101048f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_287_n N_A_391_47#_c_526_n 0.0394547f $X=3.91 $Y=1.16 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_290_n N_A_391_47#_c_526_n 0.00720931f $X=4.255 $Y=1.217
+ $X2=0 $Y2=0
cc_288 N_A_27_47#_c_291_n N_A_391_47#_c_527_n 0.00386185f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_292_n N_A_391_47#_c_527_n 0.00107777f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_300_n N_A_391_47#_c_527_n 0.0149281f $X=1.585 $Y=1.53 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_287_n N_A_391_47#_c_527_n 0.0305808f $X=3.91 $Y=1.16 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_290_n N_A_391_47#_c_527_n 0.0074788f $X=4.255 $Y=1.217 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_M1024_g N_A_391_47#_c_563_n 5.25882e-19 $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_M1036_g N_A_391_47#_c_563_n 0.00657592f $X=2.82 $Y=0.56 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_M1040_g N_A_391_47#_c_563_n 0.00693104f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_M1043_g N_A_391_47#_c_563_n 5.47131e-19 $X=3.76 $Y=0.56 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_292_n N_A_391_47#_c_567_n 8.07084e-19 $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_293_n N_A_391_47#_c_567_n 0.0141618f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_294_n N_A_391_47#_c_567_n 0.0115459f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_295_n N_A_391_47#_c_567_n 7.68612e-19 $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_M1040_g N_A_391_47#_c_501_n 0.00879805f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_M1043_g N_A_391_47#_c_501_n 0.00879805f $X=3.76 $Y=0.56 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_287_n N_A_391_47#_c_501_n 0.03957f $X=3.91 $Y=1.16 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_290_n N_A_391_47#_c_501_n 0.0031956f $X=4.255 $Y=1.217 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_294_n N_A_391_47#_c_528_n 0.0137916f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_295_n N_A_391_47#_c_528_n 0.0101048f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_287_n N_A_391_47#_c_528_n 0.0394547f $X=3.91 $Y=1.16 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_290_n N_A_391_47#_c_528_n 0.00720931f $X=4.255 $Y=1.217
+ $X2=0 $Y2=0
cc_309 N_A_27_47#_M1040_g N_A_391_47#_c_579_n 5.25882e-19 $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_M1043_g N_A_391_47#_c_579_n 0.00657592f $X=3.76 $Y=0.56 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_294_n N_A_391_47#_c_581_n 8.07084e-19 $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_295_n N_A_391_47#_c_581_n 0.0141618f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_296_n N_A_391_47#_c_581_n 0.0115459f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_M1048_g N_A_391_47#_c_502_n 0.0116573f $X=4.28 $Y=0.56 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_296_n N_A_391_47#_c_529_n 0.0151183f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_290_n N_A_391_47#_c_529_n 3.58038e-19 $X=4.255 $Y=1.217
+ $X2=0 $Y2=0
cc_317 N_A_27_47#_M1048_g N_A_391_47#_c_503_n 0.00415408f $X=4.28 $Y=0.56 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_296_n N_A_391_47#_c_504_n 8.26658e-19 $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_290_n N_A_391_47#_c_504_n 0.00331109f $X=4.255 $Y=1.217
+ $X2=0 $Y2=0
cc_320 N_A_27_47#_M1036_g N_A_391_47#_c_506_n 0.00113891f $X=2.82 $Y=0.56 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_M1040_g N_A_391_47#_c_506_n 0.00113891f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_287_n N_A_391_47#_c_506_n 0.030582f $X=3.91 $Y=1.16 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_290_n N_A_391_47#_c_506_n 0.00331919f $X=4.255 $Y=1.217
+ $X2=0 $Y2=0
cc_324 N_A_27_47#_c_293_n N_A_391_47#_c_531_n 0.00260297f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_294_n N_A_391_47#_c_531_n 0.00107777f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_287_n N_A_391_47#_c_531_n 0.0305808f $X=3.91 $Y=1.16 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_290_n N_A_391_47#_c_531_n 0.0074788f $X=4.255 $Y=1.217 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_M1043_g N_A_391_47#_c_507_n 0.0011682f $X=3.76 $Y=0.56 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_287_n N_A_391_47#_c_507_n 0.0274674f $X=3.91 $Y=1.16 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_290_n N_A_391_47#_c_507_n 0.00450461f $X=4.255 $Y=1.217
+ $X2=0 $Y2=0
cc_331 N_A_27_47#_c_295_n N_A_391_47#_c_532_n 0.00259297f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_296_n N_A_391_47#_c_532_n 0.00128868f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_c_287_n N_A_391_47#_c_532_n 0.0274092f $X=3.91 $Y=1.16 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_290_n N_A_391_47#_c_532_n 0.00735453f $X=4.255 $Y=1.217
+ $X2=0 $Y2=0
cc_335 N_A_27_47#_c_287_n N_A_391_47#_c_508_n 0.0130035f $X=3.91 $Y=1.16 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_290_n N_A_391_47#_c_508_n 0.00237077f $X=4.255 $Y=1.217
+ $X2=0 $Y2=0
cc_337 N_A_27_47#_c_290_n N_A_391_47#_c_509_n 0.0207158f $X=4.255 $Y=1.217 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_c_298_n N_VPWR_M1001_s 0.00178587f $X=0.985 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_339 N_A_27_47#_c_300_n N_VPWR_M1041_s 0.00324655f $X=1.585 $Y=1.53 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_c_297_n N_VPWR_c_946_n 0.0411685f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_341 N_A_27_47#_c_298_n N_VPWR_c_946_n 0.0136682f $X=0.985 $Y=1.53 $X2=0 $Y2=0
cc_342 N_A_27_47#_c_325_n N_VPWR_c_946_n 0.0507655f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_343 N_A_27_47#_c_325_n N_VPWR_c_947_n 0.0223557f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_344 N_A_27_47#_c_291_n N_VPWR_c_948_n 0.00497803f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_325_n N_VPWR_c_948_n 0.0416217f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_346 N_A_27_47#_c_300_n N_VPWR_c_948_n 0.0151472f $X=1.585 $Y=1.53 $X2=0 $Y2=0
cc_347 N_A_27_47#_c_291_n N_VPWR_c_949_n 0.00597712f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_292_n N_VPWR_c_949_n 0.00673617f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_292_n N_VPWR_c_950_n 0.0052072f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_350 N_A_27_47#_c_293_n N_VPWR_c_950_n 0.004751f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_351 N_A_27_47#_c_294_n N_VPWR_c_951_n 0.0052072f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_352 N_A_27_47#_c_295_n N_VPWR_c_951_n 0.004751f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_353 N_A_27_47#_c_296_n N_VPWR_c_952_n 0.0052072f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_354 N_A_27_47#_c_293_n N_VPWR_c_961_n 0.00597712f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_294_n N_VPWR_c_961_n 0.00673617f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_295_n N_VPWR_c_963_n 0.00597712f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_296_n N_VPWR_c_963_n 0.00673617f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_M1001_d N_VPWR_c_945_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_M1019_d N_VPWR_c_945_n 0.00231261f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_291_n N_VPWR_c_945_n 0.0100198f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_361 N_A_27_47#_c_292_n N_VPWR_c_945_n 0.0118438f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_362 N_A_27_47#_c_293_n N_VPWR_c_945_n 0.00999457f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_294_n N_VPWR_c_945_n 0.0118438f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_364 N_A_27_47#_c_295_n N_VPWR_c_945_n 0.00999457f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_296_n N_VPWR_c_945_n 0.011869f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_366 N_A_27_47#_c_297_n N_VPWR_c_945_n 0.0124725f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_367 N_A_27_47#_c_325_n N_VPWR_c_945_n 0.0140101f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_368 N_A_27_47#_c_297_n N_VPWR_c_983_n 0.0210596f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_369 N_A_27_47#_M1048_g N_Y_c_1187_n 4.77587e-19 $X=4.28 $Y=0.56 $X2=0 $Y2=0
cc_370 N_A_27_47#_c_296_n N_Y_c_1188_n 8.07084e-19 $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_371 N_A_27_47#_c_282_n N_VGND_M1014_s 0.00251598f $X=0.985 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_372 N_A_27_47#_c_284_n N_VGND_M1049_s 0.00193551f $X=1.585 $Y=0.82 $X2=0
+ $Y2=0
cc_373 N_A_27_47#_c_281_n N_VGND_c_1515_n 0.0184656f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_374 N_A_27_47#_c_282_n N_VGND_c_1515_n 0.0127122f $X=0.985 $Y=0.82 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_c_282_n N_VGND_c_1516_n 0.00193763f $X=0.985 $Y=0.82 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_c_323_n N_VGND_c_1516_n 0.022456f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_377 N_A_27_47#_c_284_n N_VGND_c_1516_n 0.00248202f $X=1.585 $Y=0.82 $X2=0
+ $Y2=0
cc_378 N_A_27_47#_M1021_g N_VGND_c_1517_n 0.00268723f $X=1.88 $Y=0.56 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_c_284_n N_VGND_c_1517_n 0.0135251f $X=1.585 $Y=0.82 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_M1021_g N_VGND_c_1518_n 0.00541562f $X=1.88 $Y=0.56 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_M1024_g N_VGND_c_1518_n 0.00424619f $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_M1024_g N_VGND_c_1519_n 0.00390178f $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_M1036_g N_VGND_c_1519_n 0.00276126f $X=2.82 $Y=0.56 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_M1040_g N_VGND_c_1520_n 0.00390178f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_M1043_g N_VGND_c_1520_n 0.00276126f $X=3.76 $Y=0.56 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_M1048_g N_VGND_c_1521_n 0.00268723f $X=4.28 $Y=0.56 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_M1036_g N_VGND_c_1530_n 0.00424619f $X=2.82 $Y=0.56 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_M1040_g N_VGND_c_1530_n 0.00424619f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_M1043_g N_VGND_c_1532_n 0.00424619f $X=3.76 $Y=0.56 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_M1048_g N_VGND_c_1532_n 0.00439206f $X=4.28 $Y=0.56 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_M1014_d N_VGND_c_1551_n 0.0020946f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_M1042_d N_VGND_c_1551_n 0.00304616f $X=1.015 $Y=0.235 $X2=0
+ $Y2=0
cc_393 N_A_27_47#_M1021_g N_VGND_c_1551_n 0.00965588f $X=1.88 $Y=0.56 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_M1024_g N_VGND_c_1551_n 0.00611295f $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_395 N_A_27_47#_M1036_g N_VGND_c_1551_n 0.00599018f $X=2.82 $Y=0.56 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_M1040_g N_VGND_c_1551_n 0.00611295f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_M1043_g N_VGND_c_1551_n 0.00610552f $X=3.76 $Y=0.56 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_M1048_g N_VGND_c_1551_n 0.00618081f $X=4.28 $Y=0.56 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_c_281_n N_VGND_c_1551_n 0.0123792f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_400 N_A_27_47#_c_282_n N_VGND_c_1551_n 0.00961016f $X=0.985 $Y=0.82 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_c_323_n N_VGND_c_1551_n 0.0142976f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_402 N_A_27_47#_c_284_n N_VGND_c_1551_n 0.00561929f $X=1.585 $Y=0.82 $X2=0
+ $Y2=0
cc_403 N_A_27_47#_c_281_n N_VGND_c_1552_n 0.020318f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_404 N_A_27_47#_c_282_n N_VGND_c_1552_n 0.00260082f $X=0.985 $Y=0.82 $X2=0
+ $Y2=0
cc_405 N_A_391_47#_c_526_n N_VPWR_M1005_s 0.00199888f $X=2.865 $Y=1.53 $X2=0
+ $Y2=0
cc_406 N_A_391_47#_c_528_n N_VPWR_M1023_s 0.00199888f $X=3.805 $Y=1.53 $X2=0
+ $Y2=0
cc_407 N_A_391_47#_c_529_n N_VPWR_M1035_s 0.00347056f $X=4.4 $Y=1.53 $X2=0 $Y2=0
cc_408 N_A_391_47#_c_535_n N_VPWR_c_948_n 0.0507655f $X=2.14 $Y=1.63 $X2=0 $Y2=0
cc_409 N_A_391_47#_c_535_n N_VPWR_c_949_n 0.0223557f $X=2.14 $Y=1.63 $X2=0 $Y2=0
cc_410 N_A_391_47#_c_535_n N_VPWR_c_950_n 0.0385613f $X=2.14 $Y=1.63 $X2=0 $Y2=0
cc_411 N_A_391_47#_c_526_n N_VPWR_c_950_n 0.0112848f $X=2.865 $Y=1.53 $X2=0
+ $Y2=0
cc_412 N_A_391_47#_c_567_n N_VPWR_c_950_n 0.0470327f $X=3.08 $Y=1.63 $X2=0 $Y2=0
cc_413 N_A_391_47#_c_567_n N_VPWR_c_951_n 0.0385613f $X=3.08 $Y=1.63 $X2=0 $Y2=0
cc_414 N_A_391_47#_c_528_n N_VPWR_c_951_n 0.0112848f $X=3.805 $Y=1.53 $X2=0
+ $Y2=0
cc_415 N_A_391_47#_c_581_n N_VPWR_c_951_n 0.0470327f $X=4.02 $Y=1.63 $X2=0 $Y2=0
cc_416 N_A_391_47#_c_510_n N_VPWR_c_952_n 0.004751f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_417 N_A_391_47#_c_581_n N_VPWR_c_952_n 0.0385613f $X=4.02 $Y=1.63 $X2=0 $Y2=0
cc_418 N_A_391_47#_c_529_n N_VPWR_c_952_n 0.0124926f $X=4.4 $Y=1.53 $X2=0 $Y2=0
cc_419 N_A_391_47#_c_511_n N_VPWR_c_953_n 0.0052072f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_420 N_A_391_47#_c_512_n N_VPWR_c_953_n 0.004751f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_421 N_A_391_47#_c_513_n N_VPWR_c_954_n 0.0052072f $X=6.135 $Y=1.41 $X2=0
+ $Y2=0
cc_422 N_A_391_47#_c_514_n N_VPWR_c_954_n 0.004751f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_423 N_A_391_47#_c_515_n N_VPWR_c_955_n 0.0052072f $X=7.075 $Y=1.41 $X2=0
+ $Y2=0
cc_424 N_A_391_47#_c_516_n N_VPWR_c_955_n 0.004751f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_425 N_A_391_47#_c_517_n N_VPWR_c_956_n 0.0052072f $X=8.015 $Y=1.41 $X2=0
+ $Y2=0
cc_426 N_A_391_47#_c_518_n N_VPWR_c_956_n 0.004751f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_427 N_A_391_47#_c_519_n N_VPWR_c_957_n 0.0052072f $X=8.955 $Y=1.41 $X2=0
+ $Y2=0
cc_428 N_A_391_47#_c_520_n N_VPWR_c_957_n 0.004751f $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_429 N_A_391_47#_c_521_n N_VPWR_c_958_n 0.0052072f $X=9.895 $Y=1.41 $X2=0
+ $Y2=0
cc_430 N_A_391_47#_c_522_n N_VPWR_c_958_n 0.004751f $X=10.365 $Y=1.41 $X2=0
+ $Y2=0
cc_431 N_A_391_47#_c_523_n N_VPWR_c_959_n 0.0052072f $X=10.835 $Y=1.41 $X2=0
+ $Y2=0
cc_432 N_A_391_47#_c_524_n N_VPWR_c_959_n 0.004751f $X=11.305 $Y=1.41 $X2=0
+ $Y2=0
cc_433 N_A_391_47#_c_525_n N_VPWR_c_960_n 0.00688901f $X=11.775 $Y=1.41 $X2=0
+ $Y2=0
cc_434 N_A_391_47#_c_567_n N_VPWR_c_961_n 0.0223557f $X=3.08 $Y=1.63 $X2=0 $Y2=0
cc_435 N_A_391_47#_c_581_n N_VPWR_c_963_n 0.0223557f $X=4.02 $Y=1.63 $X2=0 $Y2=0
cc_436 N_A_391_47#_c_510_n N_VPWR_c_965_n 0.00597712f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_437 N_A_391_47#_c_511_n N_VPWR_c_965_n 0.00673617f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_438 N_A_391_47#_c_512_n N_VPWR_c_967_n 0.00597712f $X=5.665 $Y=1.41 $X2=0
+ $Y2=0
cc_439 N_A_391_47#_c_513_n N_VPWR_c_967_n 0.00673617f $X=6.135 $Y=1.41 $X2=0
+ $Y2=0
cc_440 N_A_391_47#_c_514_n N_VPWR_c_969_n 0.00597712f $X=6.605 $Y=1.41 $X2=0
+ $Y2=0
cc_441 N_A_391_47#_c_515_n N_VPWR_c_969_n 0.00673617f $X=7.075 $Y=1.41 $X2=0
+ $Y2=0
cc_442 N_A_391_47#_c_516_n N_VPWR_c_971_n 0.00597712f $X=7.545 $Y=1.41 $X2=0
+ $Y2=0
cc_443 N_A_391_47#_c_517_n N_VPWR_c_971_n 0.00673617f $X=8.015 $Y=1.41 $X2=0
+ $Y2=0
cc_444 N_A_391_47#_c_518_n N_VPWR_c_973_n 0.00597712f $X=8.485 $Y=1.41 $X2=0
+ $Y2=0
cc_445 N_A_391_47#_c_519_n N_VPWR_c_973_n 0.00673617f $X=8.955 $Y=1.41 $X2=0
+ $Y2=0
cc_446 N_A_391_47#_c_520_n N_VPWR_c_975_n 0.00597712f $X=9.425 $Y=1.41 $X2=0
+ $Y2=0
cc_447 N_A_391_47#_c_521_n N_VPWR_c_975_n 0.00673617f $X=9.895 $Y=1.41 $X2=0
+ $Y2=0
cc_448 N_A_391_47#_c_522_n N_VPWR_c_977_n 0.00597712f $X=10.365 $Y=1.41 $X2=0
+ $Y2=0
cc_449 N_A_391_47#_c_523_n N_VPWR_c_977_n 0.00673617f $X=10.835 $Y=1.41 $X2=0
+ $Y2=0
cc_450 N_A_391_47#_c_524_n N_VPWR_c_979_n 0.00597712f $X=11.305 $Y=1.41 $X2=0
+ $Y2=0
cc_451 N_A_391_47#_c_525_n N_VPWR_c_979_n 0.00673617f $X=11.775 $Y=1.41 $X2=0
+ $Y2=0
cc_452 N_A_391_47#_M1000_d N_VPWR_c_945_n 0.00231261f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_453 N_A_391_47#_M1013_d N_VPWR_c_945_n 0.00231261f $X=2.935 $Y=1.485 $X2=0
+ $Y2=0
cc_454 N_A_391_47#_M1030_d N_VPWR_c_945_n 0.00231261f $X=3.875 $Y=1.485 $X2=0
+ $Y2=0
cc_455 N_A_391_47#_c_510_n N_VPWR_c_945_n 0.0100198f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_456 N_A_391_47#_c_511_n N_VPWR_c_945_n 0.0118438f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_457 N_A_391_47#_c_512_n N_VPWR_c_945_n 0.00999457f $X=5.665 $Y=1.41 $X2=0
+ $Y2=0
cc_458 N_A_391_47#_c_513_n N_VPWR_c_945_n 0.0118438f $X=6.135 $Y=1.41 $X2=0
+ $Y2=0
cc_459 N_A_391_47#_c_514_n N_VPWR_c_945_n 0.00999457f $X=6.605 $Y=1.41 $X2=0
+ $Y2=0
cc_460 N_A_391_47#_c_515_n N_VPWR_c_945_n 0.0118438f $X=7.075 $Y=1.41 $X2=0
+ $Y2=0
cc_461 N_A_391_47#_c_516_n N_VPWR_c_945_n 0.00999457f $X=7.545 $Y=1.41 $X2=0
+ $Y2=0
cc_462 N_A_391_47#_c_517_n N_VPWR_c_945_n 0.0118438f $X=8.015 $Y=1.41 $X2=0
+ $Y2=0
cc_463 N_A_391_47#_c_518_n N_VPWR_c_945_n 0.00999457f $X=8.485 $Y=1.41 $X2=0
+ $Y2=0
cc_464 N_A_391_47#_c_519_n N_VPWR_c_945_n 0.0118438f $X=8.955 $Y=1.41 $X2=0
+ $Y2=0
cc_465 N_A_391_47#_c_520_n N_VPWR_c_945_n 0.00999457f $X=9.425 $Y=1.41 $X2=0
+ $Y2=0
cc_466 N_A_391_47#_c_521_n N_VPWR_c_945_n 0.0118438f $X=9.895 $Y=1.41 $X2=0
+ $Y2=0
cc_467 N_A_391_47#_c_522_n N_VPWR_c_945_n 0.00999457f $X=10.365 $Y=1.41 $X2=0
+ $Y2=0
cc_468 N_A_391_47#_c_523_n N_VPWR_c_945_n 0.0118438f $X=10.835 $Y=1.41 $X2=0
+ $Y2=0
cc_469 N_A_391_47#_c_524_n N_VPWR_c_945_n 0.00999457f $X=11.305 $Y=1.41 $X2=0
+ $Y2=0
cc_470 N_A_391_47#_c_525_n N_VPWR_c_945_n 0.0128678f $X=11.775 $Y=1.41 $X2=0
+ $Y2=0
cc_471 N_A_391_47#_c_535_n N_VPWR_c_945_n 0.0140101f $X=2.14 $Y=1.63 $X2=0 $Y2=0
cc_472 N_A_391_47#_c_567_n N_VPWR_c_945_n 0.0140101f $X=3.08 $Y=1.63 $X2=0 $Y2=0
cc_473 N_A_391_47#_c_581_n N_VPWR_c_945_n 0.0140101f $X=4.02 $Y=1.63 $X2=0 $Y2=0
cc_474 N_A_391_47#_M1004_g N_Y_c_1189_n 0.00229101f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_475 N_A_391_47#_M1007_g N_Y_c_1189_n 0.00248233f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_476 N_A_391_47#_M1004_g N_Y_c_1187_n 0.00426764f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_477 N_A_391_47#_M1007_g N_Y_c_1187_n 0.00445433f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_478 N_A_391_47#_M1008_g N_Y_c_1187_n 4.84753e-19 $X=5.64 $Y=0.56 $X2=0 $Y2=0
cc_479 N_A_391_47#_c_510_n N_Y_c_1188_n 0.0141618f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_480 N_A_391_47#_c_511_n N_Y_c_1188_n 0.0115459f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_481 N_A_391_47#_c_512_n N_Y_c_1188_n 7.68612e-19 $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_482 N_A_391_47#_c_581_n N_Y_c_1188_n 0.00629866f $X=4.02 $Y=1.63 $X2=0 $Y2=0
cc_483 N_A_391_47#_M1007_g N_Y_c_1152_n 0.00879805f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_484 N_A_391_47#_M1008_g N_Y_c_1152_n 0.00879805f $X=5.64 $Y=0.56 $X2=0 $Y2=0
cc_485 N_A_391_47#_c_505_n N_Y_c_1152_n 0.03957f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_486 N_A_391_47#_c_509_n N_Y_c_1152_n 0.0031956f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_487 N_A_391_47#_M1004_g N_Y_c_1153_n 0.00245067f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_488 N_A_391_47#_M1007_g N_Y_c_1153_n 0.00115337f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_489 N_A_391_47#_c_502_n N_Y_c_1153_n 0.00808484f $X=4.4 $Y=0.82 $X2=0 $Y2=0
cc_490 N_A_391_47#_c_505_n N_Y_c_1153_n 0.0305973f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_491 N_A_391_47#_c_509_n N_Y_c_1153_n 0.00332f $X=11.775 $Y=1.217 $X2=0 $Y2=0
cc_492 N_A_391_47#_c_511_n N_Y_c_1169_n 0.0137916f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_493 N_A_391_47#_c_512_n N_Y_c_1169_n 0.0101048f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_494 N_A_391_47#_c_505_n N_Y_c_1169_n 0.0394547f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_495 N_A_391_47#_c_509_n N_Y_c_1169_n 0.00720931f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_496 N_A_391_47#_c_510_n N_Y_c_1170_n 0.00386185f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_497 N_A_391_47#_c_511_n N_Y_c_1170_n 0.00107777f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_498 N_A_391_47#_c_529_n N_Y_c_1170_n 0.0149281f $X=4.4 $Y=1.53 $X2=0 $Y2=0
cc_499 N_A_391_47#_c_505_n N_Y_c_1170_n 0.0305808f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_500 N_A_391_47#_c_509_n N_Y_c_1170_n 0.0074788f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_501 N_A_391_47#_M1008_g N_Y_c_1216_n 0.00226116f $X=5.64 $Y=0.56 $X2=0 $Y2=0
cc_502 N_A_391_47#_M1009_g N_Y_c_1216_n 0.00248233f $X=6.11 $Y=0.56 $X2=0 $Y2=0
cc_503 N_A_391_47#_M1007_g N_Y_c_1218_n 4.7681e-19 $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_504 N_A_391_47#_M1008_g N_Y_c_1218_n 0.0043216f $X=5.64 $Y=0.56 $X2=0 $Y2=0
cc_505 N_A_391_47#_M1009_g N_Y_c_1218_n 0.00445433f $X=6.11 $Y=0.56 $X2=0 $Y2=0
cc_506 N_A_391_47#_M1012_g N_Y_c_1218_n 4.84753e-19 $X=6.58 $Y=0.56 $X2=0 $Y2=0
cc_507 N_A_391_47#_c_511_n N_Y_c_1222_n 8.07084e-19 $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_508 N_A_391_47#_c_512_n N_Y_c_1222_n 0.0141618f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_509 N_A_391_47#_c_513_n N_Y_c_1222_n 0.0115459f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_510 N_A_391_47#_c_514_n N_Y_c_1222_n 7.68612e-19 $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_511 N_A_391_47#_M1009_g N_Y_c_1154_n 0.00879805f $X=6.11 $Y=0.56 $X2=0 $Y2=0
cc_512 N_A_391_47#_M1012_g N_Y_c_1154_n 0.00879805f $X=6.58 $Y=0.56 $X2=0 $Y2=0
cc_513 N_A_391_47#_c_505_n N_Y_c_1154_n 0.03957f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_514 N_A_391_47#_c_509_n N_Y_c_1154_n 0.0031956f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_515 N_A_391_47#_c_513_n N_Y_c_1171_n 0.0137916f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_516 N_A_391_47#_c_514_n N_Y_c_1171_n 0.0101048f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_517 N_A_391_47#_c_505_n N_Y_c_1171_n 0.0394547f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_518 N_A_391_47#_c_509_n N_Y_c_1171_n 0.00720931f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_519 N_A_391_47#_M1012_g N_Y_c_1234_n 0.00226116f $X=6.58 $Y=0.56 $X2=0 $Y2=0
cc_520 N_A_391_47#_M1016_g N_Y_c_1234_n 0.00248233f $X=7.05 $Y=0.56 $X2=0 $Y2=0
cc_521 N_A_391_47#_M1009_g N_Y_c_1236_n 4.7681e-19 $X=6.11 $Y=0.56 $X2=0 $Y2=0
cc_522 N_A_391_47#_M1012_g N_Y_c_1236_n 0.0043216f $X=6.58 $Y=0.56 $X2=0 $Y2=0
cc_523 N_A_391_47#_M1016_g N_Y_c_1236_n 0.00445433f $X=7.05 $Y=0.56 $X2=0 $Y2=0
cc_524 N_A_391_47#_M1018_g N_Y_c_1236_n 4.84753e-19 $X=7.52 $Y=0.56 $X2=0 $Y2=0
cc_525 N_A_391_47#_c_513_n N_Y_c_1240_n 8.07084e-19 $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_526 N_A_391_47#_c_514_n N_Y_c_1240_n 0.0141618f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_527 N_A_391_47#_c_515_n N_Y_c_1240_n 0.0115459f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_528 N_A_391_47#_c_516_n N_Y_c_1240_n 7.68612e-19 $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_529 N_A_391_47#_M1016_g N_Y_c_1155_n 0.00879805f $X=7.05 $Y=0.56 $X2=0 $Y2=0
cc_530 N_A_391_47#_M1018_g N_Y_c_1155_n 0.00879805f $X=7.52 $Y=0.56 $X2=0 $Y2=0
cc_531 N_A_391_47#_c_505_n N_Y_c_1155_n 0.03957f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_532 N_A_391_47#_c_509_n N_Y_c_1155_n 0.0031956f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_533 N_A_391_47#_c_515_n N_Y_c_1172_n 0.0137916f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_534 N_A_391_47#_c_516_n N_Y_c_1172_n 0.0101048f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_535 N_A_391_47#_c_505_n N_Y_c_1172_n 0.0394547f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_536 N_A_391_47#_c_509_n N_Y_c_1172_n 0.00720931f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_537 N_A_391_47#_M1016_g N_Y_c_1252_n 5.25882e-19 $X=7.05 $Y=0.56 $X2=0 $Y2=0
cc_538 N_A_391_47#_M1018_g N_Y_c_1252_n 0.00657592f $X=7.52 $Y=0.56 $X2=0 $Y2=0
cc_539 N_A_391_47#_M1022_g N_Y_c_1252_n 0.00693104f $X=7.99 $Y=0.56 $X2=0 $Y2=0
cc_540 N_A_391_47#_M1025_g N_Y_c_1252_n 5.47131e-19 $X=8.46 $Y=0.56 $X2=0 $Y2=0
cc_541 N_A_391_47#_c_515_n N_Y_c_1256_n 8.07084e-19 $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_542 N_A_391_47#_c_516_n N_Y_c_1256_n 0.0141618f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_543 N_A_391_47#_c_517_n N_Y_c_1256_n 0.0115459f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_544 N_A_391_47#_c_518_n N_Y_c_1256_n 7.68612e-19 $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_545 N_A_391_47#_M1022_g N_Y_c_1156_n 0.00879805f $X=7.99 $Y=0.56 $X2=0 $Y2=0
cc_546 N_A_391_47#_M1025_g N_Y_c_1156_n 0.00879805f $X=8.46 $Y=0.56 $X2=0 $Y2=0
cc_547 N_A_391_47#_c_505_n N_Y_c_1156_n 0.03957f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_548 N_A_391_47#_c_509_n N_Y_c_1156_n 0.0031956f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_549 N_A_391_47#_c_517_n N_Y_c_1173_n 0.0137916f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_550 N_A_391_47#_c_518_n N_Y_c_1173_n 0.0101048f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_551 N_A_391_47#_c_505_n N_Y_c_1173_n 0.0394547f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_552 N_A_391_47#_c_509_n N_Y_c_1173_n 0.00720931f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_553 N_A_391_47#_M1022_g N_Y_c_1268_n 5.25882e-19 $X=7.99 $Y=0.56 $X2=0 $Y2=0
cc_554 N_A_391_47#_M1025_g N_Y_c_1268_n 0.00657592f $X=8.46 $Y=0.56 $X2=0 $Y2=0
cc_555 N_A_391_47#_M1026_g N_Y_c_1268_n 0.00693104f $X=8.93 $Y=0.56 $X2=0 $Y2=0
cc_556 N_A_391_47#_M1029_g N_Y_c_1268_n 5.47131e-19 $X=9.4 $Y=0.56 $X2=0 $Y2=0
cc_557 N_A_391_47#_c_517_n N_Y_c_1272_n 8.07084e-19 $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_558 N_A_391_47#_c_518_n N_Y_c_1272_n 0.0141618f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_559 N_A_391_47#_c_519_n N_Y_c_1272_n 0.0115459f $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_560 N_A_391_47#_c_520_n N_Y_c_1272_n 7.68612e-19 $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_561 N_A_391_47#_M1026_g N_Y_c_1157_n 0.00879805f $X=8.93 $Y=0.56 $X2=0 $Y2=0
cc_562 N_A_391_47#_M1029_g N_Y_c_1157_n 0.00879805f $X=9.4 $Y=0.56 $X2=0 $Y2=0
cc_563 N_A_391_47#_c_505_n N_Y_c_1157_n 0.03957f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_564 N_A_391_47#_c_509_n N_Y_c_1157_n 0.0031956f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_565 N_A_391_47#_c_519_n N_Y_c_1174_n 0.0137916f $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_566 N_A_391_47#_c_520_n N_Y_c_1174_n 0.0101048f $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_567 N_A_391_47#_c_505_n N_Y_c_1174_n 0.0394547f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_568 N_A_391_47#_c_509_n N_Y_c_1174_n 0.00720931f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_569 N_A_391_47#_M1026_g N_Y_c_1284_n 5.25882e-19 $X=8.93 $Y=0.56 $X2=0 $Y2=0
cc_570 N_A_391_47#_M1029_g N_Y_c_1284_n 0.00657592f $X=9.4 $Y=0.56 $X2=0 $Y2=0
cc_571 N_A_391_47#_M1031_g N_Y_c_1284_n 0.00693104f $X=9.87 $Y=0.56 $X2=0 $Y2=0
cc_572 N_A_391_47#_M1034_g N_Y_c_1284_n 5.47131e-19 $X=10.34 $Y=0.56 $X2=0 $Y2=0
cc_573 N_A_391_47#_c_519_n N_Y_c_1288_n 8.07084e-19 $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_574 N_A_391_47#_c_520_n N_Y_c_1288_n 0.0141618f $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_575 N_A_391_47#_c_521_n N_Y_c_1288_n 0.0115459f $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_576 N_A_391_47#_c_522_n N_Y_c_1288_n 7.68612e-19 $X=10.365 $Y=1.41 $X2=0
+ $Y2=0
cc_577 N_A_391_47#_M1031_g N_Y_c_1158_n 0.00879805f $X=9.87 $Y=0.56 $X2=0 $Y2=0
cc_578 N_A_391_47#_M1034_g N_Y_c_1158_n 0.00879805f $X=10.34 $Y=0.56 $X2=0 $Y2=0
cc_579 N_A_391_47#_c_505_n N_Y_c_1158_n 0.03957f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_580 N_A_391_47#_c_509_n N_Y_c_1158_n 0.0031956f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_581 N_A_391_47#_c_521_n N_Y_c_1175_n 0.0137916f $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_582 N_A_391_47#_c_522_n N_Y_c_1175_n 0.0101048f $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_583 N_A_391_47#_c_505_n N_Y_c_1175_n 0.0394547f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_584 N_A_391_47#_c_509_n N_Y_c_1175_n 0.00720931f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_585 N_A_391_47#_M1031_g N_Y_c_1300_n 5.25882e-19 $X=9.87 $Y=0.56 $X2=0 $Y2=0
cc_586 N_A_391_47#_M1034_g N_Y_c_1300_n 0.00657592f $X=10.34 $Y=0.56 $X2=0 $Y2=0
cc_587 N_A_391_47#_M1037_g N_Y_c_1300_n 0.00693104f $X=10.81 $Y=0.56 $X2=0 $Y2=0
cc_588 N_A_391_47#_M1044_g N_Y_c_1300_n 5.47131e-19 $X=11.28 $Y=0.56 $X2=0 $Y2=0
cc_589 N_A_391_47#_c_521_n N_Y_c_1304_n 8.07084e-19 $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_590 N_A_391_47#_c_522_n N_Y_c_1304_n 0.0141618f $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_591 N_A_391_47#_c_523_n N_Y_c_1304_n 0.0115459f $X=10.835 $Y=1.41 $X2=0 $Y2=0
cc_592 N_A_391_47#_c_524_n N_Y_c_1304_n 7.68612e-19 $X=11.305 $Y=1.41 $X2=0
+ $Y2=0
cc_593 N_A_391_47#_M1037_g N_Y_c_1159_n 0.00879805f $X=10.81 $Y=0.56 $X2=0 $Y2=0
cc_594 N_A_391_47#_M1044_g N_Y_c_1159_n 0.00879805f $X=11.28 $Y=0.56 $X2=0 $Y2=0
cc_595 N_A_391_47#_c_505_n N_Y_c_1159_n 0.03957f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_596 N_A_391_47#_c_509_n N_Y_c_1159_n 0.0031956f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_597 N_A_391_47#_c_523_n N_Y_c_1176_n 0.0137916f $X=10.835 $Y=1.41 $X2=0 $Y2=0
cc_598 N_A_391_47#_c_524_n N_Y_c_1176_n 0.0101048f $X=11.305 $Y=1.41 $X2=0 $Y2=0
cc_599 N_A_391_47#_c_505_n N_Y_c_1176_n 0.0394547f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_600 N_A_391_47#_c_509_n N_Y_c_1176_n 0.00720931f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_601 N_A_391_47#_M1037_g N_Y_c_1316_n 5.25882e-19 $X=10.81 $Y=0.56 $X2=0 $Y2=0
cc_602 N_A_391_47#_M1044_g N_Y_c_1316_n 0.00657592f $X=11.28 $Y=0.56 $X2=0 $Y2=0
cc_603 N_A_391_47#_c_523_n N_Y_c_1318_n 8.07084e-19 $X=10.835 $Y=1.41 $X2=0
+ $Y2=0
cc_604 N_A_391_47#_c_524_n N_Y_c_1318_n 0.0141618f $X=11.305 $Y=1.41 $X2=0 $Y2=0
cc_605 N_A_391_47#_c_525_n N_Y_c_1318_n 0.017566f $X=11.775 $Y=1.41 $X2=0 $Y2=0
cc_606 N_A_391_47#_M1045_g N_Y_c_1160_n 0.013646f $X=11.8 $Y=0.56 $X2=0 $Y2=0
cc_607 N_A_391_47#_c_505_n N_Y_c_1160_n 3.24343e-19 $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_608 N_A_391_47#_c_525_n N_Y_c_1177_n 0.0169182f $X=11.775 $Y=1.41 $X2=0 $Y2=0
cc_609 N_A_391_47#_c_505_n N_Y_c_1177_n 3.09302e-19 $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_610 N_A_391_47#_c_509_n N_Y_c_1177_n 3.58038e-19 $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_611 N_A_391_47#_M1008_g N_Y_c_1161_n 0.00115337f $X=5.64 $Y=0.56 $X2=0 $Y2=0
cc_612 N_A_391_47#_M1009_g N_Y_c_1161_n 0.00115337f $X=6.11 $Y=0.56 $X2=0 $Y2=0
cc_613 N_A_391_47#_c_505_n N_Y_c_1161_n 0.0305905f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_614 N_A_391_47#_c_509_n N_Y_c_1161_n 0.00331994f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_615 N_A_391_47#_c_512_n N_Y_c_1178_n 0.00260297f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_616 N_A_391_47#_c_513_n N_Y_c_1178_n 0.00107777f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_617 N_A_391_47#_c_505_n N_Y_c_1178_n 0.0305808f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_618 N_A_391_47#_c_509_n N_Y_c_1178_n 0.0074788f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_619 N_A_391_47#_M1012_g N_Y_c_1162_n 0.00115337f $X=6.58 $Y=0.56 $X2=0 $Y2=0
cc_620 N_A_391_47#_M1016_g N_Y_c_1162_n 0.00115337f $X=7.05 $Y=0.56 $X2=0 $Y2=0
cc_621 N_A_391_47#_c_505_n N_Y_c_1162_n 0.0305905f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_622 N_A_391_47#_c_509_n N_Y_c_1162_n 0.00331994f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_623 N_A_391_47#_c_514_n N_Y_c_1179_n 0.00260297f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_624 N_A_391_47#_c_515_n N_Y_c_1179_n 0.00107777f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_625 N_A_391_47#_c_505_n N_Y_c_1179_n 0.0305808f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_626 N_A_391_47#_c_509_n N_Y_c_1179_n 0.0074788f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_627 N_A_391_47#_M1018_g N_Y_c_1163_n 0.00113891f $X=7.52 $Y=0.56 $X2=0 $Y2=0
cc_628 N_A_391_47#_M1022_g N_Y_c_1163_n 0.00113891f $X=7.99 $Y=0.56 $X2=0 $Y2=0
cc_629 N_A_391_47#_c_505_n N_Y_c_1163_n 0.030582f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_630 N_A_391_47#_c_509_n N_Y_c_1163_n 0.00331919f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_631 N_A_391_47#_c_516_n N_Y_c_1180_n 0.00260297f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_632 N_A_391_47#_c_517_n N_Y_c_1180_n 0.00107777f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_633 N_A_391_47#_c_505_n N_Y_c_1180_n 0.0305808f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_634 N_A_391_47#_c_509_n N_Y_c_1180_n 0.0074788f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_635 N_A_391_47#_M1025_g N_Y_c_1164_n 0.00113891f $X=8.46 $Y=0.56 $X2=0 $Y2=0
cc_636 N_A_391_47#_M1026_g N_Y_c_1164_n 0.00113891f $X=8.93 $Y=0.56 $X2=0 $Y2=0
cc_637 N_A_391_47#_c_505_n N_Y_c_1164_n 0.030582f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_638 N_A_391_47#_c_509_n N_Y_c_1164_n 0.00331919f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_639 N_A_391_47#_c_518_n N_Y_c_1181_n 0.00260297f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_640 N_A_391_47#_c_519_n N_Y_c_1181_n 0.00107777f $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_641 N_A_391_47#_c_505_n N_Y_c_1181_n 0.0305808f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_642 N_A_391_47#_c_509_n N_Y_c_1181_n 0.0074788f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_643 N_A_391_47#_M1029_g N_Y_c_1165_n 0.00113891f $X=9.4 $Y=0.56 $X2=0 $Y2=0
cc_644 N_A_391_47#_M1031_g N_Y_c_1165_n 0.00113891f $X=9.87 $Y=0.56 $X2=0 $Y2=0
cc_645 N_A_391_47#_c_505_n N_Y_c_1165_n 0.030582f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_646 N_A_391_47#_c_509_n N_Y_c_1165_n 0.00331919f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_647 N_A_391_47#_c_520_n N_Y_c_1182_n 0.00260297f $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_648 N_A_391_47#_c_521_n N_Y_c_1182_n 0.00107777f $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_649 N_A_391_47#_c_505_n N_Y_c_1182_n 0.0305808f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_650 N_A_391_47#_c_509_n N_Y_c_1182_n 0.0074788f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_651 N_A_391_47#_M1034_g N_Y_c_1166_n 0.00113891f $X=10.34 $Y=0.56 $X2=0 $Y2=0
cc_652 N_A_391_47#_M1037_g N_Y_c_1166_n 0.00113891f $X=10.81 $Y=0.56 $X2=0 $Y2=0
cc_653 N_A_391_47#_c_505_n N_Y_c_1166_n 0.030582f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_654 N_A_391_47#_c_509_n N_Y_c_1166_n 0.00331919f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_655 N_A_391_47#_c_522_n N_Y_c_1183_n 0.00260297f $X=10.365 $Y=1.41 $X2=0
+ $Y2=0
cc_656 N_A_391_47#_c_523_n N_Y_c_1183_n 0.00107777f $X=10.835 $Y=1.41 $X2=0
+ $Y2=0
cc_657 N_A_391_47#_c_505_n N_Y_c_1183_n 0.0305808f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_658 N_A_391_47#_c_509_n N_Y_c_1183_n 0.0074788f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_659 N_A_391_47#_M1044_g N_Y_c_1167_n 0.0011682f $X=11.28 $Y=0.56 $X2=0 $Y2=0
cc_660 N_A_391_47#_c_505_n N_Y_c_1167_n 0.0307156f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_661 N_A_391_47#_c_509_n N_Y_c_1167_n 0.00450461f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_662 N_A_391_47#_c_524_n N_Y_c_1184_n 0.00260297f $X=11.305 $Y=1.41 $X2=0
+ $Y2=0
cc_663 N_A_391_47#_c_525_n N_Y_c_1184_n 0.00107777f $X=11.775 $Y=1.41 $X2=0
+ $Y2=0
cc_664 N_A_391_47#_c_505_n N_Y_c_1184_n 0.0305808f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_665 N_A_391_47#_c_509_n N_Y_c_1184_n 0.00723098f $X=11.775 $Y=1.217 $X2=0
+ $Y2=0
cc_666 N_A_391_47#_c_525_n Y 0.00140994f $X=11.775 $Y=1.41 $X2=0 $Y2=0
cc_667 N_A_391_47#_M1045_g Y 0.0195212f $X=11.8 $Y=0.56 $X2=0 $Y2=0
cc_668 N_A_391_47#_c_505_n Y 0.0134881f $X=11.29 $Y=1.16 $X2=0 $Y2=0
cc_669 N_A_391_47#_c_499_n N_VGND_M1024_s 0.00251598f $X=2.865 $Y=0.82 $X2=0
+ $Y2=0
cc_670 N_A_391_47#_c_501_n N_VGND_M1040_s 0.00251598f $X=3.805 $Y=0.82 $X2=0
+ $Y2=0
cc_671 N_A_391_47#_c_502_n N_VGND_M1048_s 0.00193551f $X=4.4 $Y=0.82 $X2=0 $Y2=0
cc_672 N_A_391_47#_c_534_n N_VGND_c_1518_n 0.0216617f $X=2.14 $Y=0.4 $X2=0 $Y2=0
cc_673 N_A_391_47#_c_499_n N_VGND_c_1518_n 0.00260082f $X=2.865 $Y=0.82 $X2=0
+ $Y2=0
cc_674 N_A_391_47#_c_534_n N_VGND_c_1519_n 0.0186688f $X=2.14 $Y=0.4 $X2=0 $Y2=0
cc_675 N_A_391_47#_c_499_n N_VGND_c_1519_n 0.0127122f $X=2.865 $Y=0.82 $X2=0
+ $Y2=0
cc_676 N_A_391_47#_c_563_n N_VGND_c_1520_n 0.0186688f $X=3.08 $Y=0.4 $X2=0 $Y2=0
cc_677 N_A_391_47#_c_501_n N_VGND_c_1520_n 0.0127122f $X=3.805 $Y=0.82 $X2=0
+ $Y2=0
cc_678 N_A_391_47#_M1004_g N_VGND_c_1521_n 0.00268723f $X=4.7 $Y=0.56 $X2=0
+ $Y2=0
cc_679 N_A_391_47#_c_502_n N_VGND_c_1521_n 0.0135251f $X=4.4 $Y=0.82 $X2=0 $Y2=0
cc_680 N_A_391_47#_M1007_g N_VGND_c_1522_n 0.00382673f $X=5.17 $Y=0.56 $X2=0
+ $Y2=0
cc_681 N_A_391_47#_M1008_g N_VGND_c_1522_n 0.00276126f $X=5.64 $Y=0.56 $X2=0
+ $Y2=0
cc_682 N_A_391_47#_M1009_g N_VGND_c_1523_n 0.00382673f $X=6.11 $Y=0.56 $X2=0
+ $Y2=0
cc_683 N_A_391_47#_M1012_g N_VGND_c_1523_n 0.00276126f $X=6.58 $Y=0.56 $X2=0
+ $Y2=0
cc_684 N_A_391_47#_M1016_g N_VGND_c_1524_n 0.00382673f $X=7.05 $Y=0.56 $X2=0
+ $Y2=0
cc_685 N_A_391_47#_M1018_g N_VGND_c_1524_n 0.00276126f $X=7.52 $Y=0.56 $X2=0
+ $Y2=0
cc_686 N_A_391_47#_M1022_g N_VGND_c_1525_n 0.00390178f $X=7.99 $Y=0.56 $X2=0
+ $Y2=0
cc_687 N_A_391_47#_M1025_g N_VGND_c_1525_n 0.00276126f $X=8.46 $Y=0.56 $X2=0
+ $Y2=0
cc_688 N_A_391_47#_M1026_g N_VGND_c_1526_n 0.00390178f $X=8.93 $Y=0.56 $X2=0
+ $Y2=0
cc_689 N_A_391_47#_M1029_g N_VGND_c_1526_n 0.00276126f $X=9.4 $Y=0.56 $X2=0
+ $Y2=0
cc_690 N_A_391_47#_M1031_g N_VGND_c_1527_n 0.00390178f $X=9.87 $Y=0.56 $X2=0
+ $Y2=0
cc_691 N_A_391_47#_M1034_g N_VGND_c_1527_n 0.00276126f $X=10.34 $Y=0.56 $X2=0
+ $Y2=0
cc_692 N_A_391_47#_M1037_g N_VGND_c_1528_n 0.00390178f $X=10.81 $Y=0.56 $X2=0
+ $Y2=0
cc_693 N_A_391_47#_M1044_g N_VGND_c_1528_n 0.00276126f $X=11.28 $Y=0.56 $X2=0
+ $Y2=0
cc_694 N_A_391_47#_M1045_g N_VGND_c_1529_n 0.00438629f $X=11.8 $Y=0.56 $X2=0
+ $Y2=0
cc_695 N_A_391_47#_c_499_n N_VGND_c_1530_n 0.00193763f $X=2.865 $Y=0.82 $X2=0
+ $Y2=0
cc_696 N_A_391_47#_c_563_n N_VGND_c_1530_n 0.0216617f $X=3.08 $Y=0.4 $X2=0 $Y2=0
cc_697 N_A_391_47#_c_501_n N_VGND_c_1530_n 0.00260082f $X=3.805 $Y=0.82 $X2=0
+ $Y2=0
cc_698 N_A_391_47#_c_501_n N_VGND_c_1532_n 0.00193763f $X=3.805 $Y=0.82 $X2=0
+ $Y2=0
cc_699 N_A_391_47#_c_579_n N_VGND_c_1532_n 0.022456f $X=4.02 $Y=0.4 $X2=0 $Y2=0
cc_700 N_A_391_47#_c_502_n N_VGND_c_1532_n 0.00245178f $X=4.4 $Y=0.82 $X2=0
+ $Y2=0
cc_701 N_A_391_47#_M1004_g N_VGND_c_1534_n 0.00539841f $X=4.7 $Y=0.56 $X2=0
+ $Y2=0
cc_702 N_A_391_47#_M1007_g N_VGND_c_1534_n 0.00423108f $X=5.17 $Y=0.56 $X2=0
+ $Y2=0
cc_703 N_A_391_47#_M1008_g N_VGND_c_1536_n 0.00423108f $X=5.64 $Y=0.56 $X2=0
+ $Y2=0
cc_704 N_A_391_47#_M1009_g N_VGND_c_1536_n 0.00423108f $X=6.11 $Y=0.56 $X2=0
+ $Y2=0
cc_705 N_A_391_47#_M1012_g N_VGND_c_1538_n 0.00423108f $X=6.58 $Y=0.56 $X2=0
+ $Y2=0
cc_706 N_A_391_47#_M1016_g N_VGND_c_1538_n 0.00423108f $X=7.05 $Y=0.56 $X2=0
+ $Y2=0
cc_707 N_A_391_47#_M1018_g N_VGND_c_1540_n 0.00424619f $X=7.52 $Y=0.56 $X2=0
+ $Y2=0
cc_708 N_A_391_47#_M1022_g N_VGND_c_1540_n 0.00424619f $X=7.99 $Y=0.56 $X2=0
+ $Y2=0
cc_709 N_A_391_47#_M1025_g N_VGND_c_1542_n 0.00424619f $X=8.46 $Y=0.56 $X2=0
+ $Y2=0
cc_710 N_A_391_47#_M1026_g N_VGND_c_1542_n 0.00424619f $X=8.93 $Y=0.56 $X2=0
+ $Y2=0
cc_711 N_A_391_47#_M1029_g N_VGND_c_1544_n 0.00424619f $X=9.4 $Y=0.56 $X2=0
+ $Y2=0
cc_712 N_A_391_47#_M1031_g N_VGND_c_1544_n 0.00424619f $X=9.87 $Y=0.56 $X2=0
+ $Y2=0
cc_713 N_A_391_47#_M1034_g N_VGND_c_1546_n 0.00424619f $X=10.34 $Y=0.56 $X2=0
+ $Y2=0
cc_714 N_A_391_47#_M1037_g N_VGND_c_1546_n 0.00424619f $X=10.81 $Y=0.56 $X2=0
+ $Y2=0
cc_715 N_A_391_47#_M1044_g N_VGND_c_1548_n 0.00424619f $X=11.28 $Y=0.56 $X2=0
+ $Y2=0
cc_716 N_A_391_47#_M1045_g N_VGND_c_1548_n 0.00439206f $X=11.8 $Y=0.56 $X2=0
+ $Y2=0
cc_717 N_A_391_47#_M1021_d N_VGND_c_1551_n 0.00255524f $X=1.955 $Y=0.235 $X2=0
+ $Y2=0
cc_718 N_A_391_47#_M1036_d N_VGND_c_1551_n 0.00255524f $X=2.895 $Y=0.235 $X2=0
+ $Y2=0
cc_719 N_A_391_47#_M1043_d N_VGND_c_1551_n 0.00304616f $X=3.835 $Y=0.235 $X2=0
+ $Y2=0
cc_720 N_A_391_47#_M1004_g N_VGND_c_1551_n 0.00961873f $X=4.7 $Y=0.56 $X2=0
+ $Y2=0
cc_721 N_A_391_47#_M1007_g N_VGND_c_1551_n 0.00612203f $X=5.17 $Y=0.56 $X2=0
+ $Y2=0
cc_722 N_A_391_47#_M1008_g N_VGND_c_1551_n 0.00599926f $X=5.64 $Y=0.56 $X2=0
+ $Y2=0
cc_723 N_A_391_47#_M1009_g N_VGND_c_1551_n 0.00612203f $X=6.11 $Y=0.56 $X2=0
+ $Y2=0
cc_724 N_A_391_47#_M1012_g N_VGND_c_1551_n 0.00599926f $X=6.58 $Y=0.56 $X2=0
+ $Y2=0
cc_725 N_A_391_47#_M1016_g N_VGND_c_1551_n 0.00612203f $X=7.05 $Y=0.56 $X2=0
+ $Y2=0
cc_726 N_A_391_47#_M1018_g N_VGND_c_1551_n 0.00599018f $X=7.52 $Y=0.56 $X2=0
+ $Y2=0
cc_727 N_A_391_47#_M1022_g N_VGND_c_1551_n 0.00611295f $X=7.99 $Y=0.56 $X2=0
+ $Y2=0
cc_728 N_A_391_47#_M1025_g N_VGND_c_1551_n 0.00599018f $X=8.46 $Y=0.56 $X2=0
+ $Y2=0
cc_729 N_A_391_47#_M1026_g N_VGND_c_1551_n 0.00611295f $X=8.93 $Y=0.56 $X2=0
+ $Y2=0
cc_730 N_A_391_47#_M1029_g N_VGND_c_1551_n 0.00599018f $X=9.4 $Y=0.56 $X2=0
+ $Y2=0
cc_731 N_A_391_47#_M1031_g N_VGND_c_1551_n 0.00611295f $X=9.87 $Y=0.56 $X2=0
+ $Y2=0
cc_732 N_A_391_47#_M1034_g N_VGND_c_1551_n 0.00599018f $X=10.34 $Y=0.56 $X2=0
+ $Y2=0
cc_733 N_A_391_47#_M1037_g N_VGND_c_1551_n 0.00611295f $X=10.81 $Y=0.56 $X2=0
+ $Y2=0
cc_734 N_A_391_47#_M1044_g N_VGND_c_1551_n 0.00610552f $X=11.28 $Y=0.56 $X2=0
+ $Y2=0
cc_735 N_A_391_47#_M1045_g N_VGND_c_1551_n 0.00722383f $X=11.8 $Y=0.56 $X2=0
+ $Y2=0
cc_736 N_A_391_47#_c_534_n N_VGND_c_1551_n 0.0140924f $X=2.14 $Y=0.4 $X2=0 $Y2=0
cc_737 N_A_391_47#_c_499_n N_VGND_c_1551_n 0.00961016f $X=2.865 $Y=0.82 $X2=0
+ $Y2=0
cc_738 N_A_391_47#_c_563_n N_VGND_c_1551_n 0.0140924f $X=3.08 $Y=0.4 $X2=0 $Y2=0
cc_739 N_A_391_47#_c_501_n N_VGND_c_1551_n 0.00961016f $X=3.805 $Y=0.82 $X2=0
+ $Y2=0
cc_740 N_A_391_47#_c_579_n N_VGND_c_1551_n 0.0142976f $X=4.02 $Y=0.4 $X2=0 $Y2=0
cc_741 N_A_391_47#_c_502_n N_VGND_c_1551_n 0.00565014f $X=4.4 $Y=0.82 $X2=0
+ $Y2=0
cc_742 N_VPWR_c_945_n N_Y_M1002_d 0.00231261f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_743 N_VPWR_c_945_n N_Y_M1006_d 0.00231261f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_744 N_VPWR_c_945_n N_Y_M1011_d 0.00231261f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_745 N_VPWR_c_945_n N_Y_M1017_d 0.00231261f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_746 N_VPWR_c_945_n N_Y_M1027_d 0.00231261f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_747 N_VPWR_c_945_n N_Y_M1032_d 0.00231261f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_748 N_VPWR_c_945_n N_Y_M1038_d 0.00231261f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_749 N_VPWR_c_945_n N_Y_M1046_d 0.00231261f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_750 N_VPWR_c_952_n N_Y_c_1188_n 0.0470327f $X=4.49 $Y=2 $X2=0 $Y2=0
cc_751 N_VPWR_c_953_n N_Y_c_1188_n 0.0385613f $X=5.43 $Y=2 $X2=0 $Y2=0
cc_752 N_VPWR_c_965_n N_Y_c_1188_n 0.0223557f $X=5.345 $Y=2.72 $X2=0 $Y2=0
cc_753 N_VPWR_c_945_n N_Y_c_1188_n 0.0140101f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_754 N_VPWR_M1003_s N_Y_c_1169_n 0.00199888f $X=5.285 $Y=1.485 $X2=0 $Y2=0
cc_755 N_VPWR_c_953_n N_Y_c_1169_n 0.0112848f $X=5.43 $Y=2 $X2=0 $Y2=0
cc_756 N_VPWR_c_953_n N_Y_c_1222_n 0.0470327f $X=5.43 $Y=2 $X2=0 $Y2=0
cc_757 N_VPWR_c_954_n N_Y_c_1222_n 0.0385613f $X=6.37 $Y=2 $X2=0 $Y2=0
cc_758 N_VPWR_c_967_n N_Y_c_1222_n 0.0223557f $X=6.285 $Y=2.72 $X2=0 $Y2=0
cc_759 N_VPWR_c_945_n N_Y_c_1222_n 0.0140101f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_760 N_VPWR_M1010_s N_Y_c_1171_n 0.00199888f $X=6.225 $Y=1.485 $X2=0 $Y2=0
cc_761 N_VPWR_c_954_n N_Y_c_1171_n 0.0112848f $X=6.37 $Y=2 $X2=0 $Y2=0
cc_762 N_VPWR_c_954_n N_Y_c_1240_n 0.0470327f $X=6.37 $Y=2 $X2=0 $Y2=0
cc_763 N_VPWR_c_955_n N_Y_c_1240_n 0.0385613f $X=7.31 $Y=2 $X2=0 $Y2=0
cc_764 N_VPWR_c_969_n N_Y_c_1240_n 0.0223557f $X=7.225 $Y=2.72 $X2=0 $Y2=0
cc_765 N_VPWR_c_945_n N_Y_c_1240_n 0.0140101f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_766 N_VPWR_M1015_s N_Y_c_1172_n 0.00199888f $X=7.165 $Y=1.485 $X2=0 $Y2=0
cc_767 N_VPWR_c_955_n N_Y_c_1172_n 0.0112848f $X=7.31 $Y=2 $X2=0 $Y2=0
cc_768 N_VPWR_c_955_n N_Y_c_1256_n 0.0470327f $X=7.31 $Y=2 $X2=0 $Y2=0
cc_769 N_VPWR_c_956_n N_Y_c_1256_n 0.0385613f $X=8.25 $Y=2 $X2=0 $Y2=0
cc_770 N_VPWR_c_971_n N_Y_c_1256_n 0.0223557f $X=8.165 $Y=2.72 $X2=0 $Y2=0
cc_771 N_VPWR_c_945_n N_Y_c_1256_n 0.0140101f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_772 N_VPWR_M1020_s N_Y_c_1173_n 0.00199888f $X=8.105 $Y=1.485 $X2=0 $Y2=0
cc_773 N_VPWR_c_956_n N_Y_c_1173_n 0.0112848f $X=8.25 $Y=2 $X2=0 $Y2=0
cc_774 N_VPWR_c_956_n N_Y_c_1272_n 0.0470327f $X=8.25 $Y=2 $X2=0 $Y2=0
cc_775 N_VPWR_c_957_n N_Y_c_1272_n 0.0385613f $X=9.19 $Y=2 $X2=0 $Y2=0
cc_776 N_VPWR_c_973_n N_Y_c_1272_n 0.0223557f $X=9.105 $Y=2.72 $X2=0 $Y2=0
cc_777 N_VPWR_c_945_n N_Y_c_1272_n 0.0140101f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_778 N_VPWR_M1028_s N_Y_c_1174_n 0.00199888f $X=9.045 $Y=1.485 $X2=0 $Y2=0
cc_779 N_VPWR_c_957_n N_Y_c_1174_n 0.0112848f $X=9.19 $Y=2 $X2=0 $Y2=0
cc_780 N_VPWR_c_957_n N_Y_c_1288_n 0.0470327f $X=9.19 $Y=2 $X2=0 $Y2=0
cc_781 N_VPWR_c_958_n N_Y_c_1288_n 0.0385613f $X=10.13 $Y=2 $X2=0 $Y2=0
cc_782 N_VPWR_c_975_n N_Y_c_1288_n 0.0223557f $X=10.045 $Y=2.72 $X2=0 $Y2=0
cc_783 N_VPWR_c_945_n N_Y_c_1288_n 0.0140101f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_784 N_VPWR_M1033_s N_Y_c_1175_n 0.00199888f $X=9.985 $Y=1.485 $X2=0 $Y2=0
cc_785 N_VPWR_c_958_n N_Y_c_1175_n 0.0112848f $X=10.13 $Y=2 $X2=0 $Y2=0
cc_786 N_VPWR_c_958_n N_Y_c_1304_n 0.0470327f $X=10.13 $Y=2 $X2=0 $Y2=0
cc_787 N_VPWR_c_959_n N_Y_c_1304_n 0.0385613f $X=11.07 $Y=2 $X2=0 $Y2=0
cc_788 N_VPWR_c_977_n N_Y_c_1304_n 0.0223557f $X=10.985 $Y=2.72 $X2=0 $Y2=0
cc_789 N_VPWR_c_945_n N_Y_c_1304_n 0.0140101f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_790 N_VPWR_M1039_s N_Y_c_1176_n 0.00199888f $X=10.925 $Y=1.485 $X2=0 $Y2=0
cc_791 N_VPWR_c_959_n N_Y_c_1176_n 0.0112848f $X=11.07 $Y=2 $X2=0 $Y2=0
cc_792 N_VPWR_c_959_n N_Y_c_1318_n 0.0470327f $X=11.07 $Y=2 $X2=0 $Y2=0
cc_793 N_VPWR_c_960_n N_Y_c_1318_n 0.0385613f $X=12.01 $Y=2 $X2=0 $Y2=0
cc_794 N_VPWR_c_979_n N_Y_c_1318_n 0.0223557f $X=11.925 $Y=2.72 $X2=0 $Y2=0
cc_795 N_VPWR_c_945_n N_Y_c_1318_n 0.0140101f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_796 N_VPWR_M1047_s N_Y_c_1177_n 2.67089e-19 $X=11.865 $Y=1.485 $X2=0 $Y2=0
cc_797 N_VPWR_M1047_s Y 0.00453067f $X=11.865 $Y=1.485 $X2=0 $Y2=0
cc_798 N_VPWR_c_960_n Y 0.0121952f $X=12.01 $Y=2 $X2=0 $Y2=0
cc_799 N_Y_c_1152_n N_VGND_M1007_d 0.00251598f $X=5.685 $Y=0.82 $X2=0 $Y2=0
cc_800 N_Y_c_1154_n N_VGND_M1009_d 0.00251598f $X=6.625 $Y=0.82 $X2=0 $Y2=0
cc_801 N_Y_c_1155_n N_VGND_M1016_d 0.00251598f $X=7.565 $Y=0.82 $X2=0 $Y2=0
cc_802 N_Y_c_1156_n N_VGND_M1022_d 0.00251598f $X=8.505 $Y=0.82 $X2=0 $Y2=0
cc_803 N_Y_c_1157_n N_VGND_M1026_d 0.00251598f $X=9.445 $Y=0.82 $X2=0 $Y2=0
cc_804 N_Y_c_1158_n N_VGND_M1031_d 0.00251598f $X=10.385 $Y=0.82 $X2=0 $Y2=0
cc_805 N_Y_c_1159_n N_VGND_M1037_d 0.00251598f $X=11.325 $Y=0.82 $X2=0 $Y2=0
cc_806 N_Y_c_1160_n N_VGND_M1045_d 0.00322964f $X=11.93 $Y=0.82 $X2=0 $Y2=0
cc_807 N_Y_c_1189_n N_VGND_c_1522_n 0.0116752f $X=4.935 $Y=0.45 $X2=0 $Y2=0
cc_808 N_Y_c_1187_n N_VGND_c_1522_n 0.00700786f $X=4.935 $Y=0.735 $X2=0 $Y2=0
cc_809 N_Y_c_1152_n N_VGND_c_1522_n 0.0127122f $X=5.685 $Y=0.82 $X2=0 $Y2=0
cc_810 N_Y_c_1216_n N_VGND_c_1523_n 0.0116752f $X=5.875 $Y=0.45 $X2=0 $Y2=0
cc_811 N_Y_c_1218_n N_VGND_c_1523_n 0.00700786f $X=5.875 $Y=0.735 $X2=0 $Y2=0
cc_812 N_Y_c_1154_n N_VGND_c_1523_n 0.0127122f $X=6.625 $Y=0.82 $X2=0 $Y2=0
cc_813 N_Y_c_1234_n N_VGND_c_1524_n 0.0116752f $X=6.815 $Y=0.45 $X2=0 $Y2=0
cc_814 N_Y_c_1236_n N_VGND_c_1524_n 0.00700786f $X=6.815 $Y=0.735 $X2=0 $Y2=0
cc_815 N_Y_c_1155_n N_VGND_c_1524_n 0.0127122f $X=7.565 $Y=0.82 $X2=0 $Y2=0
cc_816 N_Y_c_1252_n N_VGND_c_1525_n 0.0186688f $X=7.78 $Y=0.4 $X2=0 $Y2=0
cc_817 N_Y_c_1156_n N_VGND_c_1525_n 0.0127122f $X=8.505 $Y=0.82 $X2=0 $Y2=0
cc_818 N_Y_c_1268_n N_VGND_c_1526_n 0.0186688f $X=8.72 $Y=0.4 $X2=0 $Y2=0
cc_819 N_Y_c_1157_n N_VGND_c_1526_n 0.0127122f $X=9.445 $Y=0.82 $X2=0 $Y2=0
cc_820 N_Y_c_1284_n N_VGND_c_1527_n 0.0186688f $X=9.66 $Y=0.4 $X2=0 $Y2=0
cc_821 N_Y_c_1158_n N_VGND_c_1527_n 0.0127122f $X=10.385 $Y=0.82 $X2=0 $Y2=0
cc_822 N_Y_c_1300_n N_VGND_c_1528_n 0.0186688f $X=10.6 $Y=0.4 $X2=0 $Y2=0
cc_823 N_Y_c_1159_n N_VGND_c_1528_n 0.0127122f $X=11.325 $Y=0.82 $X2=0 $Y2=0
cc_824 N_Y_c_1160_n N_VGND_c_1529_n 0.0140453f $X=11.93 $Y=0.82 $X2=0 $Y2=0
cc_825 N_Y_c_1189_n N_VGND_c_1534_n 0.0223797f $X=4.935 $Y=0.45 $X2=0 $Y2=0
cc_826 N_Y_c_1152_n N_VGND_c_1534_n 0.00260082f $X=5.685 $Y=0.82 $X2=0 $Y2=0
cc_827 N_Y_c_1152_n N_VGND_c_1536_n 0.00193763f $X=5.685 $Y=0.82 $X2=0 $Y2=0
cc_828 N_Y_c_1216_n N_VGND_c_1536_n 0.0221615f $X=5.875 $Y=0.45 $X2=0 $Y2=0
cc_829 N_Y_c_1154_n N_VGND_c_1536_n 0.00260082f $X=6.625 $Y=0.82 $X2=0 $Y2=0
cc_830 N_Y_c_1154_n N_VGND_c_1538_n 0.00193763f $X=6.625 $Y=0.82 $X2=0 $Y2=0
cc_831 N_Y_c_1234_n N_VGND_c_1538_n 0.0221615f $X=6.815 $Y=0.45 $X2=0 $Y2=0
cc_832 N_Y_c_1155_n N_VGND_c_1538_n 0.00260082f $X=7.565 $Y=0.82 $X2=0 $Y2=0
cc_833 N_Y_c_1155_n N_VGND_c_1540_n 0.00193763f $X=7.565 $Y=0.82 $X2=0 $Y2=0
cc_834 N_Y_c_1252_n N_VGND_c_1540_n 0.0216617f $X=7.78 $Y=0.4 $X2=0 $Y2=0
cc_835 N_Y_c_1156_n N_VGND_c_1540_n 0.00260082f $X=8.505 $Y=0.82 $X2=0 $Y2=0
cc_836 N_Y_c_1156_n N_VGND_c_1542_n 0.00193763f $X=8.505 $Y=0.82 $X2=0 $Y2=0
cc_837 N_Y_c_1268_n N_VGND_c_1542_n 0.0216617f $X=8.72 $Y=0.4 $X2=0 $Y2=0
cc_838 N_Y_c_1157_n N_VGND_c_1542_n 0.00260082f $X=9.445 $Y=0.82 $X2=0 $Y2=0
cc_839 N_Y_c_1157_n N_VGND_c_1544_n 0.00193763f $X=9.445 $Y=0.82 $X2=0 $Y2=0
cc_840 N_Y_c_1284_n N_VGND_c_1544_n 0.0216617f $X=9.66 $Y=0.4 $X2=0 $Y2=0
cc_841 N_Y_c_1158_n N_VGND_c_1544_n 0.00260082f $X=10.385 $Y=0.82 $X2=0 $Y2=0
cc_842 N_Y_c_1158_n N_VGND_c_1546_n 0.00193763f $X=10.385 $Y=0.82 $X2=0 $Y2=0
cc_843 N_Y_c_1300_n N_VGND_c_1546_n 0.0216617f $X=10.6 $Y=0.4 $X2=0 $Y2=0
cc_844 N_Y_c_1159_n N_VGND_c_1546_n 0.00260082f $X=11.325 $Y=0.82 $X2=0 $Y2=0
cc_845 N_Y_c_1159_n N_VGND_c_1548_n 0.00193763f $X=11.325 $Y=0.82 $X2=0 $Y2=0
cc_846 N_Y_c_1316_n N_VGND_c_1548_n 0.022456f $X=11.54 $Y=0.4 $X2=0 $Y2=0
cc_847 N_Y_c_1160_n N_VGND_c_1548_n 0.00248202f $X=11.93 $Y=0.82 $X2=0 $Y2=0
cc_848 N_Y_c_1160_n N_VGND_c_1550_n 0.00179231f $X=11.93 $Y=0.82 $X2=0 $Y2=0
cc_849 N_Y_M1004_s N_VGND_c_1551_n 0.00255377f $X=4.775 $Y=0.235 $X2=0 $Y2=0
cc_850 N_Y_M1008_s N_VGND_c_1551_n 0.00255431f $X=5.715 $Y=0.235 $X2=0 $Y2=0
cc_851 N_Y_M1012_s N_VGND_c_1551_n 0.00255431f $X=6.655 $Y=0.235 $X2=0 $Y2=0
cc_852 N_Y_M1018_s N_VGND_c_1551_n 0.00255524f $X=7.595 $Y=0.235 $X2=0 $Y2=0
cc_853 N_Y_M1025_s N_VGND_c_1551_n 0.00255524f $X=8.535 $Y=0.235 $X2=0 $Y2=0
cc_854 N_Y_M1029_s N_VGND_c_1551_n 0.00255524f $X=9.475 $Y=0.235 $X2=0 $Y2=0
cc_855 N_Y_M1034_s N_VGND_c_1551_n 0.00255524f $X=10.415 $Y=0.235 $X2=0 $Y2=0
cc_856 N_Y_M1044_s N_VGND_c_1551_n 0.00304616f $X=11.355 $Y=0.235 $X2=0 $Y2=0
cc_857 N_Y_c_1189_n N_VGND_c_1551_n 0.0141899f $X=4.935 $Y=0.45 $X2=0 $Y2=0
cc_858 N_Y_c_1152_n N_VGND_c_1551_n 0.00961016f $X=5.685 $Y=0.82 $X2=0 $Y2=0
cc_859 N_Y_c_1216_n N_VGND_c_1551_n 0.0141768f $X=5.875 $Y=0.45 $X2=0 $Y2=0
cc_860 N_Y_c_1154_n N_VGND_c_1551_n 0.00961016f $X=6.625 $Y=0.82 $X2=0 $Y2=0
cc_861 N_Y_c_1234_n N_VGND_c_1551_n 0.0141768f $X=6.815 $Y=0.45 $X2=0 $Y2=0
cc_862 N_Y_c_1155_n N_VGND_c_1551_n 0.00961016f $X=7.565 $Y=0.82 $X2=0 $Y2=0
cc_863 N_Y_c_1252_n N_VGND_c_1551_n 0.0140924f $X=7.78 $Y=0.4 $X2=0 $Y2=0
cc_864 N_Y_c_1156_n N_VGND_c_1551_n 0.00961016f $X=8.505 $Y=0.82 $X2=0 $Y2=0
cc_865 N_Y_c_1268_n N_VGND_c_1551_n 0.0140924f $X=8.72 $Y=0.4 $X2=0 $Y2=0
cc_866 N_Y_c_1157_n N_VGND_c_1551_n 0.00961016f $X=9.445 $Y=0.82 $X2=0 $Y2=0
cc_867 N_Y_c_1284_n N_VGND_c_1551_n 0.0140924f $X=9.66 $Y=0.4 $X2=0 $Y2=0
cc_868 N_Y_c_1158_n N_VGND_c_1551_n 0.00961016f $X=10.385 $Y=0.82 $X2=0 $Y2=0
cc_869 N_Y_c_1300_n N_VGND_c_1551_n 0.0140924f $X=10.6 $Y=0.4 $X2=0 $Y2=0
cc_870 N_Y_c_1159_n N_VGND_c_1551_n 0.00961016f $X=11.325 $Y=0.82 $X2=0 $Y2=0
cc_871 N_Y_c_1316_n N_VGND_c_1551_n 0.0142976f $X=11.54 $Y=0.4 $X2=0 $Y2=0
cc_872 N_Y_c_1160_n N_VGND_c_1551_n 0.00873756f $X=11.93 $Y=0.82 $X2=0 $Y2=0
