* File: sky130_fd_sc_hdll__muxb16to1_2.pxi.spice
* Created: Thu Aug 27 19:11:31 2020
* 
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[0] N_D[0]_M1010_g N_D[0]_M1042_g
+ N_D[0]_M1108_g N_D[0]_M1075_g D[0] N_D[0]_c_852_n N_D[0]_c_853_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[0]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[8] N_D[8]_M1014_g N_D[8]_M1047_g
+ N_D[8]_M1118_g N_D[8]_M1078_g D[8] N_D[8]_c_903_n N_D[8]_c_904_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[8]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_278_265# N_A_278_265#_M1081_s
+ N_A_278_265#_M1023_s N_A_278_265#_M1013_g N_A_278_265#_c_956_n
+ N_A_278_265#_c_957_n N_A_278_265#_M1031_g N_A_278_265#_c_951_n
+ N_A_278_265#_c_952_n N_A_278_265#_c_959_n N_A_278_265#_c_953_n
+ N_A_278_265#_c_954_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_278_265#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_278_793# N_A_278_793#_M1115_s
+ N_A_278_793#_M1027_s N_A_278_793#_M1099_g N_A_278_793#_c_1039_n
+ N_A_278_793#_c_1040_n N_A_278_793#_M1111_g N_A_278_793#_c_1035_n
+ N_A_278_793#_c_1036_n N_A_278_793#_c_1043_n N_A_278_793#_c_1037_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_278_793#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[0] N_S[0]_c_1114_n N_S[0]_M1032_g
+ N_S[0]_c_1115_n N_S[0]_c_1116_n N_S[0]_c_1117_n N_S[0]_M1041_g N_S[0]_c_1118_n
+ N_S[0]_c_1119_n N_S[0]_c_1120_n N_S[0]_c_1121_n N_S[0]_c_1122_n N_S[0]_M1023_g
+ N_S[0]_c_1123_n N_S[0]_M1081_g N_S[0]_c_1124_n S[0]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[0]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[8] N_S[8]_c_1180_n N_S[8]_M1020_g
+ N_S[8]_c_1181_n N_S[8]_c_1182_n N_S[8]_c_1183_n N_S[8]_M1104_g N_S[8]_c_1184_n
+ N_S[8]_c_1185_n N_S[8]_c_1186_n N_S[8]_c_1187_n N_S[8]_c_1191_n N_S[8]_M1027_g
+ N_S[8]_c_1188_n N_S[8]_M1115_g N_S[8]_c_1189_n S[8]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[8]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[1] N_S[1]_c_1246_n N_S[1]_M1072_g
+ N_S[1]_c_1247_n N_S[1]_M1089_g N_S[1]_c_1248_n N_S[1]_c_1249_n N_S[1]_c_1250_n
+ N_S[1]_c_1251_n N_S[1]_c_1252_n N_S[1]_M1028_g N_S[1]_c_1253_n N_S[1]_c_1254_n
+ N_S[1]_M1037_g N_S[1]_c_1255_n S[1] PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[1]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[9] N_S[9]_c_1309_n N_S[9]_M1039_g
+ N_S[9]_c_1320_n N_S[9]_M1092_g N_S[9]_c_1310_n N_S[9]_c_1311_n N_S[9]_c_1312_n
+ N_S[9]_c_1313_n N_S[9]_c_1314_n N_S[9]_M1048_g N_S[9]_c_1315_n N_S[9]_c_1316_n
+ N_S[9]_M1130_g N_S[9]_c_1317_n S[9] PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[9]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_701_47# N_A_701_47#_M1072_d
+ N_A_701_47#_M1089_d N_A_701_47#_M1084_g N_A_701_47#_c_1380_n
+ N_A_701_47#_c_1375_n N_A_701_47#_M1113_g N_A_701_47#_c_1383_n
+ N_A_701_47#_c_1376_n N_A_701_47#_c_1377_n N_A_701_47#_c_1378_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_701_47#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_701_937# N_A_701_937#_M1039_d
+ N_A_701_937#_M1092_d N_A_701_937#_M1036_g N_A_701_937#_c_1461_n
+ N_A_701_937#_c_1456_n N_A_701_937#_M1157_g N_A_701_937#_c_1464_n
+ N_A_701_937#_c_1457_n N_A_701_937#_c_1458_n N_A_701_937#_c_1459_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_701_937#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[1] N_D[1]_M1052_g N_D[1]_M1074_g
+ N_D[1]_M1105_g N_D[1]_M1097_g D[1] N_D[1]_c_1542_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[1]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[9] N_D[9]_M1056_g N_D[9]_M1026_g
+ N_D[9]_M1059_g N_D[9]_M1101_g D[9] N_D[9]_c_1599_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[9]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[2] N_D[2]_M1003_g N_D[2]_M1117_g
+ N_D[2]_M1127_g N_D[2]_M1120_g D[2] N_D[2]_c_1655_n N_D[2]_c_1656_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[2]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[10] N_D[10]_M1009_g N_D[10]_M1035_g
+ N_D[10]_M1109_g N_D[10]_M1126_g D[10] N_D[10]_c_1713_n N_D[10]_c_1714_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[10]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1566_265# N_A_1566_265#_M1150_s
+ N_A_1566_265#_M1133_s N_A_1566_265#_M1005_g N_A_1566_265#_c_1773_n
+ N_A_1566_265#_c_1774_n N_A_1566_265#_M1124_g N_A_1566_265#_c_1768_n
+ N_A_1566_265#_c_1769_n N_A_1566_265#_c_1776_n N_A_1566_265#_c_1770_n
+ N_A_1566_265#_c_1771_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1566_265#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1566_793# N_A_1566_793#_M1033_s
+ N_A_1566_793#_M1137_s N_A_1566_793#_M1044_g N_A_1566_793#_c_1857_n
+ N_A_1566_793#_c_1858_n N_A_1566_793#_M1095_g N_A_1566_793#_c_1853_n
+ N_A_1566_793#_c_1854_n N_A_1566_793#_c_1861_n N_A_1566_793#_c_1855_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1566_793#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[2] N_S[2]_c_1933_n N_S[2]_M1116_g
+ N_S[2]_c_1934_n N_S[2]_c_1935_n N_S[2]_c_1936_n N_S[2]_M1151_g N_S[2]_c_1937_n
+ N_S[2]_c_1938_n N_S[2]_c_1939_n N_S[2]_c_1940_n N_S[2]_c_1941_n N_S[2]_M1133_g
+ N_S[2]_c_1942_n N_S[2]_M1150_g N_S[2]_c_1943_n S[2]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[2]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[10] N_S[10]_c_1999_n N_S[10]_M1015_g
+ N_S[10]_c_2000_n N_S[10]_c_2001_n N_S[10]_c_2002_n N_S[10]_M1043_g
+ N_S[10]_c_2003_n N_S[10]_c_2004_n N_S[10]_c_2005_n N_S[10]_c_2006_n
+ N_S[10]_c_2010_n N_S[10]_M1137_g N_S[10]_c_2007_n N_S[10]_M1033_g
+ N_S[10]_c_2008_n S[10] PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[10]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[3] N_S[3]_c_2065_n N_S[3]_M1019_g
+ N_S[3]_c_2066_n N_S[3]_M1053_g N_S[3]_c_2067_n N_S[3]_c_2068_n N_S[3]_c_2069_n
+ N_S[3]_c_2070_n N_S[3]_c_2071_n N_S[3]_M1102_g N_S[3]_c_2072_n N_S[3]_c_2073_n
+ N_S[3]_M1125_g N_S[3]_c_2074_n S[3] PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[3]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[11] N_S[11]_c_2128_n N_S[11]_M1071_g
+ N_S[11]_c_2139_n N_S[11]_M1060_g N_S[11]_c_2129_n N_S[11]_c_2130_n
+ N_S[11]_c_2131_n N_S[11]_c_2132_n N_S[11]_c_2133_n N_S[11]_M1029_g
+ N_S[11]_c_2134_n N_S[11]_c_2135_n N_S[11]_M1067_g N_S[11]_c_2136_n S[11]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[11]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1989_47# N_A_1989_47#_M1019_d
+ N_A_1989_47#_M1053_d N_A_1989_47#_M1004_g N_A_1989_47#_c_2199_n
+ N_A_1989_47#_c_2194_n N_A_1989_47#_M1123_g N_A_1989_47#_c_2202_n
+ N_A_1989_47#_c_2195_n N_A_1989_47#_c_2196_n N_A_1989_47#_c_2197_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1989_47#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1989_937# N_A_1989_937#_M1071_d
+ N_A_1989_937#_M1060_d N_A_1989_937#_M1045_g N_A_1989_937#_c_2280_n
+ N_A_1989_937#_c_2275_n N_A_1989_937#_M1093_g N_A_1989_937#_c_2283_n
+ N_A_1989_937#_c_2276_n N_A_1989_937#_c_2277_n N_A_1989_937#_c_2278_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1989_937#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[3] N_D[3]_M1002_g N_D[3]_M1025_g
+ N_D[3]_M1156_g N_D[3]_M1135_g D[3] N_D[3]_c_2361_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[3]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[11] N_D[11]_M1008_g N_D[11]_M1011_g
+ N_D[11]_M1136_g N_D[11]_M1141_g D[11] N_D[11]_c_2418_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[11]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[4] N_D[4]_M1030_g N_D[4]_M1057_g
+ N_D[4]_M1094_g N_D[4]_M1080_g D[4] N_D[4]_c_2474_n N_D[4]_c_2475_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[4]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[12] N_D[12]_M1038_g N_D[12]_M1073_g
+ N_D[12]_M1103_g N_D[12]_M1088_g D[12] N_D[12]_c_2532_n N_D[12]_c_2533_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[12]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2854_265# N_A_2854_265#_M1064_s
+ N_A_2854_265#_M1001_s N_A_2854_265#_M1034_g N_A_2854_265#_c_2592_n
+ N_A_2854_265#_c_2593_n N_A_2854_265#_M1083_g N_A_2854_265#_c_2587_n
+ N_A_2854_265#_c_2588_n N_A_2854_265#_c_2595_n N_A_2854_265#_c_2589_n
+ N_A_2854_265#_c_2590_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2854_265#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2854_793# N_A_2854_793#_M1063_s
+ N_A_2854_793#_M1007_s N_A_2854_793#_M1114_g N_A_2854_793#_c_2676_n
+ N_A_2854_793#_c_2677_n N_A_2854_793#_M1159_g N_A_2854_793#_c_2672_n
+ N_A_2854_793#_c_2673_n N_A_2854_793#_c_2680_n N_A_2854_793#_c_2674_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2854_793#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[4] N_S[4]_c_2752_n N_S[4]_M1046_g
+ N_S[4]_c_2753_n N_S[4]_c_2754_n N_S[4]_c_2755_n N_S[4]_M1086_g N_S[4]_c_2756_n
+ N_S[4]_c_2757_n N_S[4]_c_2758_n N_S[4]_c_2759_n N_S[4]_c_2760_n N_S[4]_M1001_g
+ N_S[4]_c_2761_n N_S[4]_M1064_g N_S[4]_c_2762_n S[4]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[4]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[12] N_S[12]_c_2818_n N_S[12]_M1000_g
+ N_S[12]_c_2819_n N_S[12]_c_2820_n N_S[12]_c_2821_n N_S[12]_M1128_g
+ N_S[12]_c_2822_n N_S[12]_c_2823_n N_S[12]_c_2824_n N_S[12]_c_2825_n
+ N_S[12]_c_2829_n N_S[12]_M1007_g N_S[12]_c_2826_n N_S[12]_M1063_g
+ N_S[12]_c_2827_n S[12] PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[12]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[5] N_S[5]_c_2884_n N_S[5]_M1098_g
+ N_S[5]_c_2885_n N_S[5]_M1065_g N_S[5]_c_2886_n N_S[5]_c_2887_n N_S[5]_c_2888_n
+ N_S[5]_c_2889_n N_S[5]_c_2890_n N_S[5]_M1022_g N_S[5]_c_2891_n N_S[5]_c_2892_n
+ N_S[5]_M1054_g N_S[5]_c_2893_n S[5] PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[5]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[13] N_S[13]_c_2947_n N_S[13]_M1096_g
+ N_S[13]_c_2958_n N_S[13]_M1070_g N_S[13]_c_2948_n N_S[13]_c_2949_n
+ N_S[13]_c_2950_n N_S[13]_c_2951_n N_S[13]_c_2952_n N_S[13]_M1016_g
+ N_S[13]_c_2953_n N_S[13]_c_2954_n N_S[13]_M1146_g N_S[13]_c_2955_n S[13]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[13]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3277_47# N_A_3277_47#_M1098_d
+ N_A_3277_47#_M1065_d N_A_3277_47#_M1055_g N_A_3277_47#_c_3018_n
+ N_A_3277_47#_c_3013_n N_A_3277_47#_M1082_g N_A_3277_47#_c_3021_n
+ N_A_3277_47#_c_3014_n N_A_3277_47#_c_3015_n N_A_3277_47#_c_3016_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3277_47#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3277_937# N_A_3277_937#_M1096_d
+ N_A_3277_937#_M1070_d N_A_3277_937#_M1134_g N_A_3277_937#_c_3099_n
+ N_A_3277_937#_c_3094_n N_A_3277_937#_M1158_g N_A_3277_937#_c_3102_n
+ N_A_3277_937#_c_3095_n N_A_3277_937#_c_3096_n N_A_3277_937#_c_3097_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3277_937#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[5] N_D[5]_M1051_g N_D[5]_M1090_g
+ N_D[5]_M1110_g N_D[5]_M1079_g D[5] N_D[5]_c_3180_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[5]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[13] N_D[13]_M1058_g N_D[13]_M1100_g
+ N_D[13]_M1121_g N_D[13]_M1087_g D[13] N_D[13]_c_3237_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[13]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[6] N_D[6]_M1062_g N_D[6]_M1139_g
+ N_D[6]_M1155_g N_D[6]_M1143_g D[6] N_D[6]_c_3293_n N_D[6]_c_3294_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[6]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[14] N_D[14]_M1069_g N_D[14]_M1018_g
+ N_D[14]_M1119_g N_D[14]_M1152_g D[14] N_D[14]_c_3351_n N_D[14]_c_3352_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[14]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4142_265# N_A_4142_265#_M1144_s
+ N_A_4142_265#_M1077_s N_A_4142_265#_M1066_g N_A_4142_265#_c_3411_n
+ N_A_4142_265#_c_3412_n N_A_4142_265#_M1091_g N_A_4142_265#_c_3406_n
+ N_A_4142_265#_c_3407_n N_A_4142_265#_c_3414_n N_A_4142_265#_c_3408_n
+ N_A_4142_265#_c_3409_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4142_265#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4142_793# N_A_4142_793#_M1012_s
+ N_A_4142_793#_M1085_s N_A_4142_793#_M1006_g N_A_4142_793#_c_3495_n
+ N_A_4142_793#_c_3496_n N_A_4142_793#_M1140_g N_A_4142_793#_c_3491_n
+ N_A_4142_793#_c_3492_n N_A_4142_793#_c_3499_n N_A_4142_793#_c_3493_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4142_793#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[6] N_S[6]_c_3571_n N_S[6]_M1112_g
+ N_S[6]_c_3572_n N_S[6]_c_3573_n N_S[6]_c_3574_n N_S[6]_M1145_g N_S[6]_c_3575_n
+ N_S[6]_c_3576_n N_S[6]_c_3577_n N_S[6]_c_3578_n N_S[6]_c_3579_n N_S[6]_M1077_g
+ N_S[6]_c_3580_n N_S[6]_M1144_g N_S[6]_c_3581_n S[6]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[6]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[14] N_S[14]_c_3637_n N_S[14]_M1021_g
+ N_S[14]_c_3638_n N_S[14]_c_3639_n N_S[14]_c_3640_n N_S[14]_M1153_g
+ N_S[14]_c_3641_n N_S[14]_c_3642_n N_S[14]_c_3643_n N_S[14]_c_3644_n
+ N_S[14]_c_3648_n N_S[14]_M1085_g N_S[14]_c_3645_n N_S[14]_M1012_g
+ N_S[14]_c_3646_n S[14] PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[14]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[7] N_S[7]_c_3703_n N_S[7]_M1017_g
+ N_S[7]_c_3704_n N_S[7]_M1129_g N_S[7]_c_3705_n N_S[7]_c_3706_n N_S[7]_c_3707_n
+ N_S[7]_c_3708_n N_S[7]_c_3709_n N_S[7]_M1107_g N_S[7]_c_3710_n N_S[7]_c_3711_n
+ N_S[7]_M1138_g N_S[7]_c_3712_n S[7] PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[7]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[15] N_S[15]_c_3766_n N_S[15]_M1040_g
+ N_S[15]_c_3777_n N_S[15]_M1132_g N_S[15]_c_3767_n N_S[15]_c_3768_n
+ N_S[15]_c_3769_n N_S[15]_c_3770_n N_S[15]_c_3771_n N_S[15]_M1106_g
+ N_S[15]_c_3772_n N_S[15]_c_3773_n N_S[15]_M1131_g N_S[15]_c_3774_n S[15]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%S[15]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4565_47# N_A_4565_47#_M1017_d
+ N_A_4565_47#_M1129_d N_A_4565_47#_M1122_g N_A_4565_47#_c_3837_n
+ N_A_4565_47#_c_3832_n N_A_4565_47#_M1148_g N_A_4565_47#_c_3840_n
+ N_A_4565_47#_c_3833_n N_A_4565_47#_c_3834_n N_A_4565_47#_c_3835_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4565_47#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4565_937# N_A_4565_937#_M1040_d
+ N_A_4565_937#_M1132_d N_A_4565_937#_M1049_g N_A_4565_937#_c_3917_n
+ N_A_4565_937#_c_3912_n N_A_4565_937#_M1076_g N_A_4565_937#_c_3920_n
+ N_A_4565_937#_c_3913_n N_A_4565_937#_c_3914_n N_A_4565_937#_c_3915_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4565_937#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[7] N_D[7]_M1061_g N_D[7]_M1024_g
+ N_D[7]_M1050_g N_D[7]_M1142_g D[7] N_D[7]_c_3997_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[7]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[15] N_D[15]_M1068_g N_D[15]_M1147_g
+ N_D[15]_M1154_g N_D[15]_M1149_g D[15] N_D[15]_c_4047_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%D[15]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_27_297# N_A_27_297#_M1010_d
+ N_A_27_297#_M1075_d N_A_27_297#_M1031_d N_A_27_297#_c_4092_n
+ N_A_27_297#_c_4099_n N_A_27_297#_c_4103_n N_A_27_297#_c_4121_p
+ N_A_27_297#_c_4108_n N_A_27_297#_c_4110_n N_A_27_297#_c_4093_n
+ N_A_27_297#_c_4111_n N_A_27_297#_c_4094_n N_A_27_297#_c_4113_n
+ N_A_27_297#_c_4106_n N_A_27_297#_c_4095_n N_A_27_297#_c_4096_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_27_591# N_A_27_591#_M1014_d
+ N_A_27_591#_M1078_d N_A_27_591#_M1111_d N_A_27_591#_c_4170_n
+ N_A_27_591#_c_4175_n N_A_27_591#_c_4171_n N_A_27_591#_c_4186_n
+ N_A_27_591#_c_4172_n N_A_27_591#_c_4181_n N_A_27_591#_c_4200_p
+ N_A_27_591#_c_4191_n N_A_27_591#_c_4193_n N_A_27_591#_c_4183_n
+ N_A_27_591#_c_4173_n N_A_27_591#_c_4174_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_27_591#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%VPWR N_VPWR_M1010_s N_VPWR_M1014_s
+ N_VPWR_M1023_d N_VPWR_M1027_d N_VPWR_M1052_s N_VPWR_M1056_s N_VPWR_M1003_d
+ N_VPWR_M1009_d N_VPWR_M1133_d N_VPWR_M1137_d N_VPWR_M1002_d N_VPWR_M1008_d
+ N_VPWR_M1030_s N_VPWR_M1038_s N_VPWR_M1001_d N_VPWR_M1007_d N_VPWR_M1051_s
+ N_VPWR_M1058_s N_VPWR_M1062_s N_VPWR_M1069_s N_VPWR_M1077_d N_VPWR_M1085_d
+ N_VPWR_M1061_s N_VPWR_M1068_s N_VPWR_c_4246_n N_VPWR_c_4247_n N_VPWR_c_4248_n
+ N_VPWR_c_4249_n N_VPWR_c_4250_n N_VPWR_c_4251_n N_VPWR_c_4252_n
+ N_VPWR_c_4253_n N_VPWR_c_4254_n N_VPWR_c_4255_n N_VPWR_c_4256_n
+ N_VPWR_c_4257_n N_VPWR_c_4258_n N_VPWR_c_4259_n N_VPWR_c_4260_n
+ N_VPWR_c_4261_n N_VPWR_c_4262_n N_VPWR_c_4263_n N_VPWR_c_4264_n
+ N_VPWR_c_4265_n N_VPWR_c_4266_n N_VPWR_c_4267_n N_VPWR_c_4268_n
+ N_VPWR_c_4269_n N_VPWR_c_4306_n N_VPWR_c_4314_n N_VPWR_c_4270_n
+ N_VPWR_c_4271_n N_VPWR_c_4376_n N_VPWR_c_4384_n N_VPWR_c_4392_n
+ N_VPWR_c_4400_n N_VPWR_c_4272_n N_VPWR_c_4273_n N_VPWR_c_4462_n
+ N_VPWR_c_4470_n N_VPWR_c_4478_n N_VPWR_c_4486_n N_VPWR_c_4274_n
+ N_VPWR_c_4275_n N_VPWR_c_4548_n N_VPWR_c_4556_n N_VPWR_c_4564_n
+ N_VPWR_c_4572_n N_VPWR_c_4276_n N_VPWR_c_4277_n N_VPWR_c_4634_n
+ N_VPWR_c_4642_n VPWR VPWR VPWR VPWR VPWR VPWR VPWR VPWR N_VPWR_c_4279_n
+ N_VPWR_c_4280_n N_VPWR_c_4281_n N_VPWR_c_4282_n N_VPWR_c_4283_n
+ N_VPWR_c_4284_n N_VPWR_c_4285_n N_VPWR_c_4286_n N_VPWR_c_4287_n
+ N_VPWR_c_4288_n N_VPWR_c_4289_n N_VPWR_c_4290_n N_VPWR_c_4291_n
+ N_VPWR_c_4292_n N_VPWR_c_4293_n N_VPWR_c_4294_n N_VPWR_c_4295_n
+ N_VPWR_c_4296_n N_VPWR_c_4297_n N_VPWR_c_4298_n N_VPWR_c_4299_n
+ N_VPWR_c_4300_n N_VPWR_c_4301_n N_VPWR_c_4302_n N_VPWR_c_4303_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%VPWR
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%Z N_Z_M1032_s N_Z_M1020_s N_Z_M1028_s
+ N_Z_M1048_d N_Z_M1116_d N_Z_M1015_d N_Z_M1102_d N_Z_M1029_d N_Z_M1046_d
+ N_Z_M1000_s N_Z_M1022_d N_Z_M1016_s N_Z_M1112_d N_Z_M1021_s N_Z_M1107_d
+ N_Z_M1106_d N_Z_M1013_s N_Z_M1099_s N_Z_M1084_s N_Z_M1036_d N_Z_M1005_d
+ N_Z_M1044_s N_Z_M1004_d N_Z_M1045_s N_Z_M1034_s N_Z_M1114_s N_Z_M1055_s
+ N_Z_M1134_s N_Z_M1066_s N_Z_M1006_d N_Z_M1122_s N_Z_M1049_s N_Z_c_5202_n
+ N_Z_c_5203_n N_Z_c_5204_n N_Z_c_5205_n N_Z_c_5206_n N_Z_c_5207_n N_Z_c_5208_n
+ N_Z_c_5209_n N_Z_c_5210_n N_Z_c_5211_n N_Z_c_5212_n N_Z_c_5213_n N_Z_c_5214_n
+ N_Z_c_5215_n N_Z_c_5216_n N_Z_c_5217_n N_Z_c_5218_n N_Z_c_5219_n N_Z_c_5220_n
+ N_Z_c_5221_n N_Z_c_5222_n N_Z_c_5223_n N_Z_c_5224_n N_Z_c_5225_n N_Z_c_5242_n
+ N_Z_c_5287_n N_Z_c_5243_n N_Z_c_5313_n N_Z_c_5244_n N_Z_c_5357_n N_Z_c_5245_n
+ N_Z_c_5383_n N_Z_c_5246_n N_Z_c_5426_n N_Z_c_5247_n N_Z_c_5453_n N_Z_c_5248_n
+ N_Z_c_5497_n N_Z_c_5249_n N_Z_c_5523_n N_Z_c_5250_n N_Z_c_5566_n N_Z_c_5251_n
+ N_Z_c_5593_n N_Z_c_5252_n N_Z_c_5637_n N_Z_c_5253_n N_Z_c_5663_n N_Z_c_5254_n
+ N_Z_c_5706_n N_Z_c_5255_n N_Z_c_5733_n Z Z Z Z Z Z Z Z Z Z Z Z Z Z Z Z
+ N_Z_c_5288_n N_Z_c_5226_n N_Z_c_5297_n N_Z_c_5257_n N_Z_c_5358_n N_Z_c_5227_n
+ N_Z_c_5367_n N_Z_c_5259_n N_Z_c_5427_n N_Z_c_5228_n N_Z_c_5436_n N_Z_c_5261_n
+ N_Z_c_5498_n N_Z_c_5229_n N_Z_c_5507_n N_Z_c_5263_n N_Z_c_5567_n N_Z_c_5230_n
+ N_Z_c_5576_n N_Z_c_5265_n N_Z_c_5638_n N_Z_c_5231_n N_Z_c_5647_n N_Z_c_5267_n
+ N_Z_c_5707_n N_Z_c_5232_n N_Z_c_5716_n N_Z_c_5269_n N_Z_c_5777_n N_Z_c_5233_n
+ N_Z_c_5786_n N_Z_c_5271_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%Z
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_824_333# N_A_824_333#_M1084_d
+ N_A_824_333#_M1113_d N_A_824_333#_M1097_d N_A_824_333#_c_6435_n
+ N_A_824_333#_c_6423_n N_A_824_333#_c_6418_n N_A_824_333#_c_6424_n
+ N_A_824_333#_c_6419_n N_A_824_333#_c_6441_n N_A_824_333#_c_6427_n
+ N_A_824_333#_c_6428_n N_A_824_333#_c_6429_n N_A_824_333#_c_6466_n
+ N_A_824_333#_c_6420_n N_A_824_333#_c_6421_n N_A_824_333#_c_6434_n
+ N_A_824_333#_c_6422_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_824_333#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_824_591# N_A_824_591#_M1036_s
+ N_A_824_591#_M1157_s N_A_824_591#_M1101_d N_A_824_591#_c_6514_n
+ N_A_824_591#_c_6519_n N_A_824_591#_c_6515_n N_A_824_591#_c_6516_n
+ N_A_824_591#_c_6524_n N_A_824_591#_c_6525_n N_A_824_591#_c_6517_n
+ N_A_824_591#_c_6534_n N_A_824_591#_c_6528_n N_A_824_591#_c_6529_n
+ N_A_824_591#_c_6562_n N_A_824_591#_c_6518_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_824_591#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1315_297# N_A_1315_297#_M1003_s
+ N_A_1315_297#_M1120_s N_A_1315_297#_M1124_s N_A_1315_297#_c_6605_n
+ N_A_1315_297#_c_6612_n N_A_1315_297#_c_6616_n N_A_1315_297#_c_6642_n
+ N_A_1315_297#_c_6621_n N_A_1315_297#_c_6623_n N_A_1315_297#_c_6606_n
+ N_A_1315_297#_c_6624_n N_A_1315_297#_c_6607_n N_A_1315_297#_c_6626_n
+ N_A_1315_297#_c_6619_n N_A_1315_297#_c_6608_n N_A_1315_297#_c_6609_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1315_297#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1315_591# N_A_1315_591#_M1009_s
+ N_A_1315_591#_M1126_s N_A_1315_591#_M1095_d N_A_1315_591#_c_6699_n
+ N_A_1315_591#_c_6704_n N_A_1315_591#_c_6700_n N_A_1315_591#_c_6715_n
+ N_A_1315_591#_c_6701_n N_A_1315_591#_c_6710_n N_A_1315_591#_c_6742_n
+ N_A_1315_591#_c_6720_n N_A_1315_591#_c_6722_n N_A_1315_591#_c_6712_n
+ N_A_1315_591#_c_6702_n N_A_1315_591#_c_6703_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1315_591#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2112_333# N_A_2112_333#_M1004_s
+ N_A_2112_333#_M1123_s N_A_2112_333#_M1135_s N_A_2112_333#_c_6808_n
+ N_A_2112_333#_c_6796_n N_A_2112_333#_c_6791_n N_A_2112_333#_c_6797_n
+ N_A_2112_333#_c_6792_n N_A_2112_333#_c_6814_n N_A_2112_333#_c_6800_n
+ N_A_2112_333#_c_6801_n N_A_2112_333#_c_6802_n N_A_2112_333#_c_6839_n
+ N_A_2112_333#_c_6793_n N_A_2112_333#_c_6794_n N_A_2112_333#_c_6807_n
+ N_A_2112_333#_c_6795_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2112_333#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2112_591# N_A_2112_591#_M1045_d
+ N_A_2112_591#_M1093_d N_A_2112_591#_M1141_s N_A_2112_591#_c_6887_n
+ N_A_2112_591#_c_6892_n N_A_2112_591#_c_6888_n N_A_2112_591#_c_6889_n
+ N_A_2112_591#_c_6897_n N_A_2112_591#_c_6898_n N_A_2112_591#_c_6890_n
+ N_A_2112_591#_c_6907_n N_A_2112_591#_c_6901_n N_A_2112_591#_c_6902_n
+ N_A_2112_591#_c_6935_n N_A_2112_591#_c_6891_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2112_591#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2603_297# N_A_2603_297#_M1030_d
+ N_A_2603_297#_M1080_d N_A_2603_297#_M1083_d N_A_2603_297#_c_6978_n
+ N_A_2603_297#_c_6985_n N_A_2603_297#_c_6989_n N_A_2603_297#_c_7015_n
+ N_A_2603_297#_c_6994_n N_A_2603_297#_c_6996_n N_A_2603_297#_c_6979_n
+ N_A_2603_297#_c_6997_n N_A_2603_297#_c_6980_n N_A_2603_297#_c_6999_n
+ N_A_2603_297#_c_6992_n N_A_2603_297#_c_6981_n N_A_2603_297#_c_6982_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2603_297#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2603_591# N_A_2603_591#_M1038_d
+ N_A_2603_591#_M1088_d N_A_2603_591#_M1159_d N_A_2603_591#_c_7072_n
+ N_A_2603_591#_c_7077_n N_A_2603_591#_c_7073_n N_A_2603_591#_c_7088_n
+ N_A_2603_591#_c_7074_n N_A_2603_591#_c_7083_n N_A_2603_591#_c_7115_n
+ N_A_2603_591#_c_7093_n N_A_2603_591#_c_7095_n N_A_2603_591#_c_7085_n
+ N_A_2603_591#_c_7075_n N_A_2603_591#_c_7076_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2603_591#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3400_333# N_A_3400_333#_M1055_d
+ N_A_3400_333#_M1082_d N_A_3400_333#_M1079_d N_A_3400_333#_c_7181_n
+ N_A_3400_333#_c_7169_n N_A_3400_333#_c_7164_n N_A_3400_333#_c_7170_n
+ N_A_3400_333#_c_7165_n N_A_3400_333#_c_7187_n N_A_3400_333#_c_7173_n
+ N_A_3400_333#_c_7174_n N_A_3400_333#_c_7175_n N_A_3400_333#_c_7212_n
+ N_A_3400_333#_c_7166_n N_A_3400_333#_c_7167_n N_A_3400_333#_c_7180_n
+ N_A_3400_333#_c_7168_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3400_333#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3400_591# N_A_3400_591#_M1134_d
+ N_A_3400_591#_M1158_d N_A_3400_591#_M1087_d N_A_3400_591#_c_7260_n
+ N_A_3400_591#_c_7265_n N_A_3400_591#_c_7261_n N_A_3400_591#_c_7262_n
+ N_A_3400_591#_c_7270_n N_A_3400_591#_c_7271_n N_A_3400_591#_c_7263_n
+ N_A_3400_591#_c_7280_n N_A_3400_591#_c_7274_n N_A_3400_591#_c_7275_n
+ N_A_3400_591#_c_7308_n N_A_3400_591#_c_7264_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3400_591#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3891_297# N_A_3891_297#_M1062_d
+ N_A_3891_297#_M1143_d N_A_3891_297#_M1091_d N_A_3891_297#_c_7351_n
+ N_A_3891_297#_c_7358_n N_A_3891_297#_c_7362_n N_A_3891_297#_c_7388_n
+ N_A_3891_297#_c_7367_n N_A_3891_297#_c_7369_n N_A_3891_297#_c_7352_n
+ N_A_3891_297#_c_7370_n N_A_3891_297#_c_7353_n N_A_3891_297#_c_7372_n
+ N_A_3891_297#_c_7365_n N_A_3891_297#_c_7354_n N_A_3891_297#_c_7355_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3891_297#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3891_591# N_A_3891_591#_M1069_d
+ N_A_3891_591#_M1152_d N_A_3891_591#_M1140_s N_A_3891_591#_c_7445_n
+ N_A_3891_591#_c_7450_n N_A_3891_591#_c_7446_n N_A_3891_591#_c_7461_n
+ N_A_3891_591#_c_7447_n N_A_3891_591#_c_7456_n N_A_3891_591#_c_7488_n
+ N_A_3891_591#_c_7466_n N_A_3891_591#_c_7468_n N_A_3891_591#_c_7458_n
+ N_A_3891_591#_c_7448_n N_A_3891_591#_c_7449_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3891_591#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4688_333# N_A_4688_333#_M1122_d
+ N_A_4688_333#_M1148_d N_A_4688_333#_M1142_d N_A_4688_333#_c_7554_n
+ N_A_4688_333#_c_7542_n N_A_4688_333#_c_7537_n N_A_4688_333#_c_7543_n
+ N_A_4688_333#_c_7538_n N_A_4688_333#_c_7560_n N_A_4688_333#_c_7546_n
+ N_A_4688_333#_c_7547_n N_A_4688_333#_c_7548_n N_A_4688_333#_c_7585_n
+ N_A_4688_333#_c_7539_n N_A_4688_333#_c_7540_n N_A_4688_333#_c_7553_n
+ N_A_4688_333#_c_7541_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4688_333#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4688_591# N_A_4688_591#_M1049_d
+ N_A_4688_591#_M1076_d N_A_4688_591#_M1149_d N_A_4688_591#_c_7617_n
+ N_A_4688_591#_c_7622_n N_A_4688_591#_c_7618_n N_A_4688_591#_c_7619_n
+ N_A_4688_591#_c_7627_n N_A_4688_591#_c_7628_n N_A_4688_591#_c_7620_n
+ N_A_4688_591#_c_7637_n N_A_4688_591#_c_7631_n N_A_4688_591#_c_7632_n
+ N_A_4688_591#_c_7664_n N_A_4688_591#_c_7621_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4688_591#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_27_47# N_A_27_47#_M1042_d
+ N_A_27_47#_M1108_d N_A_27_47#_M1041_d N_A_27_47#_c_7695_n N_A_27_47#_c_7692_n
+ N_A_27_47#_c_7693_n N_A_27_47#_c_7724_p N_A_27_47#_c_7694_n
+ N_A_27_47#_c_7705_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_27_911# N_A_27_911#_M1047_s
+ N_A_27_911#_M1118_s N_A_27_911#_M1104_d N_A_27_911#_c_7737_n
+ N_A_27_911#_c_7734_n N_A_27_911#_c_7735_n N_A_27_911#_c_7768_p
+ N_A_27_911#_c_7748_n N_A_27_911#_c_7736_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_27_911#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%VGND N_VGND_M1042_s N_VGND_M1047_d
+ N_VGND_M1081_d N_VGND_M1115_d N_VGND_M1074_d N_VGND_M1026_d N_VGND_M1117_s
+ N_VGND_M1035_s N_VGND_M1150_d N_VGND_M1033_d N_VGND_M1025_s N_VGND_M1011_s
+ N_VGND_M1057_d N_VGND_M1073_d N_VGND_M1064_d N_VGND_M1063_d N_VGND_M1090_d
+ N_VGND_M1100_d N_VGND_M1139_d N_VGND_M1018_d N_VGND_M1144_d N_VGND_M1012_d
+ N_VGND_M1024_s N_VGND_M1147_s N_VGND_c_7777_n N_VGND_c_7778_n N_VGND_c_7779_n
+ N_VGND_c_7780_n N_VGND_c_7781_n N_VGND_c_7782_n N_VGND_c_7783_n
+ N_VGND_c_7784_n N_VGND_c_7785_n N_VGND_c_7786_n N_VGND_c_7787_n
+ N_VGND_c_7788_n N_VGND_c_7789_n N_VGND_c_7790_n N_VGND_c_7791_n
+ N_VGND_c_7792_n N_VGND_c_7793_n N_VGND_c_7794_n N_VGND_c_7795_n
+ N_VGND_c_7796_n N_VGND_c_7797_n N_VGND_c_7798_n N_VGND_c_7799_n
+ N_VGND_c_7800_n N_VGND_c_7801_n N_VGND_c_7802_n N_VGND_c_7803_n
+ N_VGND_c_7804_n N_VGND_c_7805_n N_VGND_c_7806_n N_VGND_c_7807_n
+ N_VGND_c_7808_n N_VGND_c_7809_n N_VGND_c_7810_n N_VGND_c_7811_n
+ N_VGND_c_7812_n N_VGND_c_7813_n N_VGND_c_7814_n N_VGND_c_7815_n
+ N_VGND_c_7816_n N_VGND_c_7817_n N_VGND_c_7818_n N_VGND_c_7819_n
+ N_VGND_c_7820_n N_VGND_c_7821_n N_VGND_c_7822_n N_VGND_c_7823_n
+ N_VGND_c_7824_n N_VGND_c_7825_n N_VGND_c_7826_n VGND VGND VGND VGND VGND VGND
+ VGND VGND VGND VGND VGND VGND VGND VGND VGND VGND N_VGND_c_7829_n
+ N_VGND_c_7830_n N_VGND_c_7831_n N_VGND_c_7832_n N_VGND_c_7833_n
+ N_VGND_c_7834_n N_VGND_c_7835_n N_VGND_c_7836_n N_VGND_c_7837_n
+ N_VGND_c_7838_n N_VGND_c_7839_n N_VGND_c_7840_n N_VGND_c_7841_n
+ N_VGND_c_7842_n N_VGND_c_7843_n N_VGND_c_7844_n N_VGND_c_7845_n
+ N_VGND_c_7846_n N_VGND_c_7847_n N_VGND_c_7848_n N_VGND_c_7849_n
+ N_VGND_c_7850_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%VGND
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_845_69# N_A_845_69#_M1028_d
+ N_A_845_69#_M1037_d N_A_845_69#_M1105_s N_A_845_69#_c_8343_n
+ N_A_845_69#_c_8339_n N_A_845_69#_c_8340_n N_A_845_69#_c_8376_n
+ N_A_845_69#_c_8341_n N_A_845_69#_c_8342_n N_A_845_69#_c_8361_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_845_69#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_845_915# N_A_845_915#_M1048_s
+ N_A_845_915#_M1130_s N_A_845_915#_M1059_s N_A_845_915#_c_8391_n
+ N_A_845_915#_c_8387_n N_A_845_915#_c_8388_n N_A_845_915#_c_8389_n
+ N_A_845_915#_c_8405_n N_A_845_915#_c_8390_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_845_915#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1315_47# N_A_1315_47#_M1117_d
+ N_A_1315_47#_M1127_d N_A_1315_47#_M1151_s N_A_1315_47#_c_8437_n
+ N_A_1315_47#_c_8434_n N_A_1315_47#_c_8435_n N_A_1315_47#_c_8472_n
+ N_A_1315_47#_c_8436_n N_A_1315_47#_c_8447_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1315_47#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1315_911# N_A_1315_911#_M1035_d
+ N_A_1315_911#_M1109_d N_A_1315_911#_M1043_s N_A_1315_911#_c_8481_n
+ N_A_1315_911#_c_8478_n N_A_1315_911#_c_8479_n N_A_1315_911#_c_8517_n
+ N_A_1315_911#_c_8492_n N_A_1315_911#_c_8480_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_1315_911#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2133_69# N_A_2133_69#_M1102_s
+ N_A_2133_69#_M1125_s N_A_2133_69#_M1156_d N_A_2133_69#_c_8526_n
+ N_A_2133_69#_c_8522_n N_A_2133_69#_c_8523_n N_A_2133_69#_c_8559_n
+ N_A_2133_69#_c_8524_n N_A_2133_69#_c_8525_n N_A_2133_69#_c_8544_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2133_69#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2133_915# N_A_2133_915#_M1029_s
+ N_A_2133_915#_M1067_s N_A_2133_915#_M1136_d N_A_2133_915#_c_8574_n
+ N_A_2133_915#_c_8570_n N_A_2133_915#_c_8571_n N_A_2133_915#_c_8572_n
+ N_A_2133_915#_c_8588_n N_A_2133_915#_c_8573_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2133_915#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2603_47# N_A_2603_47#_M1057_s
+ N_A_2603_47#_M1094_s N_A_2603_47#_M1086_s N_A_2603_47#_c_8620_n
+ N_A_2603_47#_c_8617_n N_A_2603_47#_c_8618_n N_A_2603_47#_c_8655_n
+ N_A_2603_47#_c_8619_n N_A_2603_47#_c_8630_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2603_47#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2603_911# N_A_2603_911#_M1073_s
+ N_A_2603_911#_M1103_s N_A_2603_911#_M1128_d N_A_2603_911#_c_8664_n
+ N_A_2603_911#_c_8661_n N_A_2603_911#_c_8662_n N_A_2603_911#_c_8700_n
+ N_A_2603_911#_c_8675_n N_A_2603_911#_c_8663_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_2603_911#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3421_69# N_A_3421_69#_M1022_s
+ N_A_3421_69#_M1054_s N_A_3421_69#_M1110_s N_A_3421_69#_c_8709_n
+ N_A_3421_69#_c_8705_n N_A_3421_69#_c_8706_n N_A_3421_69#_c_8742_n
+ N_A_3421_69#_c_8707_n N_A_3421_69#_c_8708_n N_A_3421_69#_c_8727_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3421_69#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3421_915# N_A_3421_915#_M1016_d
+ N_A_3421_915#_M1146_d N_A_3421_915#_M1121_s N_A_3421_915#_c_8757_n
+ N_A_3421_915#_c_8753_n N_A_3421_915#_c_8754_n N_A_3421_915#_c_8755_n
+ N_A_3421_915#_c_8771_n N_A_3421_915#_c_8756_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3421_915#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3891_47# N_A_3891_47#_M1139_s
+ N_A_3891_47#_M1155_s N_A_3891_47#_M1145_s N_A_3891_47#_c_8803_n
+ N_A_3891_47#_c_8800_n N_A_3891_47#_c_8801_n N_A_3891_47#_c_8838_n
+ N_A_3891_47#_c_8802_n N_A_3891_47#_c_8813_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3891_47#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3891_911# N_A_3891_911#_M1018_s
+ N_A_3891_911#_M1119_s N_A_3891_911#_M1153_d N_A_3891_911#_c_8847_n
+ N_A_3891_911#_c_8844_n N_A_3891_911#_c_8845_n N_A_3891_911#_c_8883_n
+ N_A_3891_911#_c_8858_n N_A_3891_911#_c_8846_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_3891_911#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4709_69# N_A_4709_69#_M1107_s
+ N_A_4709_69#_M1138_s N_A_4709_69#_M1050_d N_A_4709_69#_c_8892_n
+ N_A_4709_69#_c_8888_n N_A_4709_69#_c_8889_n N_A_4709_69#_c_8925_n
+ N_A_4709_69#_c_8890_n N_A_4709_69#_c_8891_n N_A_4709_69#_c_8910_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4709_69#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4709_915# N_A_4709_915#_M1106_s
+ N_A_4709_915#_M1131_s N_A_4709_915#_M1154_d N_A_4709_915#_c_8938_n
+ N_A_4709_915#_c_8934_n N_A_4709_915#_c_8935_n N_A_4709_915#_c_8936_n
+ N_A_4709_915#_c_8952_n N_A_4709_915#_c_8937_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_2%A_4709_915#
cc_1 VNB N_D[0]_M1010_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_2 VNB N_D[0]_M1042_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_3 VNB N_D[0]_M1108_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_4 VNB N_D[0]_M1075_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_5 VNB N_D[0]_c_852_n 0.0128835f $X=-0.19 $Y=-0.24 $X2=0.75 $Y2=1.16
cc_6 VNB N_D[0]_c_853_n 0.0571683f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_7 VNB N_D[8]_M1014_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_8 VNB N_D[8]_M1047_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_9 VNB N_D[8]_M1118_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_10 VNB N_D[8]_M1078_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_11 VNB N_D[8]_c_903_n 0.0128835f $X=-0.19 $Y=-0.24 $X2=0.75 $Y2=1.16
cc_12 VNB N_D[8]_c_904_n 0.0571683f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_13 VNB N_A_278_265#_c_951_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_14 VNB N_A_278_265#_c_952_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_278_265#_c_953_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_16 VNB N_A_278_265#_c_954_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_278_793#_c_1035_n 0.0147415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_278_793#_c_1036_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_19 VNB N_A_278_793#_c_1037_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_S[0]_c_1114_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_21 VNB N_S[0]_c_1115_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_S[0]_c_1116_n 0.0101495f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.025
cc_23 VNB N_S[0]_c_1117_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_24 VNB N_S[0]_c_1118_n 0.032124f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_25 VNB N_S[0]_c_1119_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_S[0]_c_1120_n 0.0222544f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_27 VNB N_S[0]_c_1121_n 0.0073997f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_28 VNB N_S[0]_c_1122_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_29 VNB N_S[0]_c_1123_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_S[0]_c_1124_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_31 VNB S[0] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_S[8]_c_1180_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_33 VNB N_S[8]_c_1181_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_S[8]_c_1182_n 0.0101495f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.025
cc_35 VNB N_S[8]_c_1183_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_36 VNB N_S[8]_c_1184_n 0.032124f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_37 VNB N_S[8]_c_1185_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_S[8]_c_1186_n 0.0222544f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_39 VNB N_S[8]_c_1187_n 0.0073997f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_40 VNB N_S[8]_c_1188_n 0.0456684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_S[8]_c_1189_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_42 VNB S[8] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_S[1]_c_1246_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_44 VNB N_S[1]_c_1247_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_S[1]_c_1248_n 0.0296541f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_46 VNB N_S[1]_c_1249_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_47 VNB N_S[1]_c_1250_n 0.0214653f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_48 VNB N_S[1]_c_1251_n 0.0106587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_S[1]_c_1252_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_50 VNB N_S[1]_c_1253_n 0.0254151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_S[1]_c_1254_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_S[1]_c_1255_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_53 VNB S[1] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_S[9]_c_1309_n 0.0456684f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_55 VNB N_S[9]_c_1310_n 0.0296541f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_56 VNB N_S[9]_c_1311_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_57 VNB N_S[9]_c_1312_n 0.0214653f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_58 VNB N_S[9]_c_1313_n 0.0106587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_S[9]_c_1314_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_60 VNB N_S[9]_c_1315_n 0.0254151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_S[9]_c_1316_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_S[9]_c_1317_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_63 VNB S[9] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_701_47#_c_1375_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_701_47#_c_1376_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_701_47#_c_1377_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_67 VNB N_A_701_47#_c_1378_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_68 VNB N_A_701_937#_c_1456_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_701_937#_c_1457_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_701_937#_c_1458_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_71 VNB N_A_701_937#_c_1459_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_72 VNB N_D[1]_M1052_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_73 VNB N_D[1]_M1074_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_74 VNB N_D[1]_M1105_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_75 VNB N_D[1]_M1097_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_76 VNB D[1] 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_77 VNB N_D[1]_c_1542_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_78 VNB N_D[9]_M1056_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_79 VNB N_D[9]_M1026_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_80 VNB N_D[9]_M1059_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_81 VNB N_D[9]_M1101_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_82 VNB D[9] 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_83 VNB N_D[9]_c_1599_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_84 VNB N_D[2]_M1003_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_85 VNB N_D[2]_M1117_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_86 VNB N_D[2]_M1127_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_87 VNB N_D[2]_M1120_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_88 VNB N_D[2]_c_1655_n 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.75 $Y2=1.16
cc_89 VNB N_D[2]_c_1656_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_90 VNB N_D[10]_M1009_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_91 VNB N_D[10]_M1035_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_92 VNB N_D[10]_M1109_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_93 VNB N_D[10]_M1126_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_94 VNB N_D[10]_c_1713_n 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.75 $Y2=1.16
cc_95 VNB N_D[10]_c_1714_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_96 VNB N_A_1566_265#_c_1768_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.105
cc_97 VNB N_A_1566_265#_c_1769_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_A_1566_265#_c_1770_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_99 VNB N_A_1566_265#_c_1771_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_A_1566_793#_c_1853_n 0.0147415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_A_1566_793#_c_1854_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.41
+ $Y2=1.16
cc_102 VNB N_A_1566_793#_c_1855_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_S[2]_c_1933_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_104 VNB N_S[2]_c_1934_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_S[2]_c_1935_n 0.0101495f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.025
cc_106 VNB N_S[2]_c_1936_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_107 VNB N_S[2]_c_1937_n 0.032124f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_108 VNB N_S[2]_c_1938_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_S[2]_c_1939_n 0.0222544f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_110 VNB N_S[2]_c_1940_n 0.0073997f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_111 VNB N_S[2]_c_1941_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_112 VNB N_S[2]_c_1942_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_S[2]_c_1943_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_114 VNB S[2] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_S[10]_c_1999_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_116 VNB N_S[10]_c_2000_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_S[10]_c_2001_n 0.0101495f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.025
cc_118 VNB N_S[10]_c_2002_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_119 VNB N_S[10]_c_2003_n 0.032124f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_120 VNB N_S[10]_c_2004_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_S[10]_c_2005_n 0.0222544f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_122 VNB N_S[10]_c_2006_n 0.0073997f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_123 VNB N_S[10]_c_2007_n 0.0456684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_S[10]_c_2008_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_125 VNB S[10] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_S[3]_c_2065_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_127 VNB N_S[3]_c_2066_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_S[3]_c_2067_n 0.0296541f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_129 VNB N_S[3]_c_2068_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_130 VNB N_S[3]_c_2069_n 0.0214653f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_131 VNB N_S[3]_c_2070_n 0.0106587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_132 VNB N_S[3]_c_2071_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_133 VNB N_S[3]_c_2072_n 0.0254151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_134 VNB N_S[3]_c_2073_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_135 VNB N_S[3]_c_2074_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_136 VNB S[3] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_137 VNB N_S[11]_c_2128_n 0.0456684f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_138 VNB N_S[11]_c_2129_n 0.0296541f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_139 VNB N_S[11]_c_2130_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_140 VNB N_S[11]_c_2131_n 0.0214653f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_141 VNB N_S[11]_c_2132_n 0.0106587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_142 VNB N_S[11]_c_2133_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_143 VNB N_S[11]_c_2134_n 0.0254151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_144 VNB N_S[11]_c_2135_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_145 VNB N_S[11]_c_2136_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_146 VNB S[11] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_147 VNB N_A_1989_47#_c_2194_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_148 VNB N_A_1989_47#_c_2195_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_149 VNB N_A_1989_47#_c_2196_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_150 VNB N_A_1989_47#_c_2197_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_151 VNB N_A_1989_937#_c_2275_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_152 VNB N_A_1989_937#_c_2276_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_153 VNB N_A_1989_937#_c_2277_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.52
+ $Y2=1.16
cc_154 VNB N_A_1989_937#_c_2278_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94
+ $Y2=1.16
cc_155 VNB N_D[3]_M1002_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_156 VNB N_D[3]_M1025_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_157 VNB N_D[3]_M1156_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_158 VNB N_D[3]_M1135_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_159 VNB D[3] 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_160 VNB N_D[3]_c_2361_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_161 VNB N_D[11]_M1008_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_162 VNB N_D[11]_M1011_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_163 VNB N_D[11]_M1136_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_164 VNB N_D[11]_M1141_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_165 VNB D[11] 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_166 VNB N_D[11]_c_2418_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_167 VNB N_D[4]_M1030_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_168 VNB N_D[4]_M1057_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_169 VNB N_D[4]_M1094_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_170 VNB N_D[4]_M1080_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_171 VNB N_D[4]_c_2474_n 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.75 $Y2=1.16
cc_172 VNB N_D[4]_c_2475_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_173 VNB N_D[12]_M1038_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_174 VNB N_D[12]_M1073_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_175 VNB N_D[12]_M1103_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_176 VNB N_D[12]_M1088_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_177 VNB N_D[12]_c_2532_n 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.75 $Y2=1.16
cc_178 VNB N_D[12]_c_2533_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_179 VNB N_A_2854_265#_c_2587_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.105
cc_180 VNB N_A_2854_265#_c_2588_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_181 VNB N_A_2854_265#_c_2589_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94
+ $Y2=1.16
cc_182 VNB N_A_2854_265#_c_2590_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_183 VNB N_A_2854_793#_c_2672_n 0.0147415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_184 VNB N_A_2854_793#_c_2673_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.41
+ $Y2=1.16
cc_185 VNB N_A_2854_793#_c_2674_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_186 VNB N_S[4]_c_2752_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_187 VNB N_S[4]_c_2753_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_188 VNB N_S[4]_c_2754_n 0.0101495f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.025
cc_189 VNB N_S[4]_c_2755_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_190 VNB N_S[4]_c_2756_n 0.032124f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_191 VNB N_S[4]_c_2757_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_192 VNB N_S[4]_c_2758_n 0.0222544f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_193 VNB N_S[4]_c_2759_n 0.0073997f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_194 VNB N_S[4]_c_2760_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_195 VNB N_S[4]_c_2761_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_196 VNB N_S[4]_c_2762_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_197 VNB S[4] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_198 VNB N_S[12]_c_2818_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_199 VNB N_S[12]_c_2819_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_200 VNB N_S[12]_c_2820_n 0.0101495f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.025
cc_201 VNB N_S[12]_c_2821_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_202 VNB N_S[12]_c_2822_n 0.032124f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_203 VNB N_S[12]_c_2823_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_204 VNB N_S[12]_c_2824_n 0.0222544f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_205 VNB N_S[12]_c_2825_n 0.0073997f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_206 VNB N_S[12]_c_2826_n 0.0456684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_207 VNB N_S[12]_c_2827_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_208 VNB S[12] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_209 VNB N_S[5]_c_2884_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_210 VNB N_S[5]_c_2885_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_211 VNB N_S[5]_c_2886_n 0.0296541f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_212 VNB N_S[5]_c_2887_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_213 VNB N_S[5]_c_2888_n 0.0214653f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_214 VNB N_S[5]_c_2889_n 0.0106587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_215 VNB N_S[5]_c_2890_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_216 VNB N_S[5]_c_2891_n 0.0254151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_217 VNB N_S[5]_c_2892_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_218 VNB N_S[5]_c_2893_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_219 VNB S[5] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_220 VNB N_S[13]_c_2947_n 0.0456684f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_221 VNB N_S[13]_c_2948_n 0.0296541f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_222 VNB N_S[13]_c_2949_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_223 VNB N_S[13]_c_2950_n 0.0214653f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_224 VNB N_S[13]_c_2951_n 0.0106587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_225 VNB N_S[13]_c_2952_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_226 VNB N_S[13]_c_2953_n 0.0254151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_227 VNB N_S[13]_c_2954_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_228 VNB N_S[13]_c_2955_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_229 VNB S[13] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_230 VNB N_A_3277_47#_c_3013_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_231 VNB N_A_3277_47#_c_3014_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_232 VNB N_A_3277_47#_c_3015_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_233 VNB N_A_3277_47#_c_3016_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_234 VNB N_A_3277_937#_c_3094_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_235 VNB N_A_3277_937#_c_3095_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_236 VNB N_A_3277_937#_c_3096_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.52
+ $Y2=1.16
cc_237 VNB N_A_3277_937#_c_3097_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94
+ $Y2=1.16
cc_238 VNB N_D[5]_M1051_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_239 VNB N_D[5]_M1090_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_240 VNB N_D[5]_M1110_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_241 VNB N_D[5]_M1079_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_242 VNB D[5] 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_243 VNB N_D[5]_c_3180_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_244 VNB N_D[13]_M1058_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_245 VNB N_D[13]_M1100_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_246 VNB N_D[13]_M1121_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_247 VNB N_D[13]_M1087_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_248 VNB D[13] 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_249 VNB N_D[13]_c_3237_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_250 VNB N_D[6]_M1062_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_251 VNB N_D[6]_M1139_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_252 VNB N_D[6]_M1155_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_253 VNB N_D[6]_M1143_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_254 VNB N_D[6]_c_3293_n 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.75 $Y2=1.16
cc_255 VNB N_D[6]_c_3294_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_256 VNB N_D[14]_M1069_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_257 VNB N_D[14]_M1018_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_258 VNB N_D[14]_M1119_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_259 VNB N_D[14]_M1152_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_260 VNB N_D[14]_c_3351_n 0.00447828f $X=-0.19 $Y=-0.24 $X2=0.75 $Y2=1.16
cc_261 VNB N_D[14]_c_3352_n 0.0542469f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_262 VNB N_A_4142_265#_c_3406_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.105
cc_263 VNB N_A_4142_265#_c_3407_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_264 VNB N_A_4142_265#_c_3408_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94
+ $Y2=1.16
cc_265 VNB N_A_4142_265#_c_3409_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_266 VNB N_A_4142_793#_c_3491_n 0.0147415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_267 VNB N_A_4142_793#_c_3492_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.41
+ $Y2=1.16
cc_268 VNB N_A_4142_793#_c_3493_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_269 VNB N_S[6]_c_3571_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_270 VNB N_S[6]_c_3572_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_271 VNB N_S[6]_c_3573_n 0.0101495f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.025
cc_272 VNB N_S[6]_c_3574_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_273 VNB N_S[6]_c_3575_n 0.032124f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_274 VNB N_S[6]_c_3576_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_275 VNB N_S[6]_c_3577_n 0.0222544f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_276 VNB N_S[6]_c_3578_n 0.0073997f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_277 VNB N_S[6]_c_3579_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_278 VNB N_S[6]_c_3580_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_279 VNB N_S[6]_c_3581_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_280 VNB S[6] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_281 VNB N_S[14]_c_3637_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_282 VNB N_S[14]_c_3638_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_283 VNB N_S[14]_c_3639_n 0.0101495f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.025
cc_284 VNB N_S[14]_c_3640_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_285 VNB N_S[14]_c_3641_n 0.032124f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_286 VNB N_S[14]_c_3642_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_287 VNB N_S[14]_c_3643_n 0.0222544f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_288 VNB N_S[14]_c_3644_n 0.0073997f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_289 VNB N_S[14]_c_3645_n 0.0456684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_290 VNB N_S[14]_c_3646_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_291 VNB S[14] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_292 VNB N_S[7]_c_3703_n 0.0169105f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_293 VNB N_S[7]_c_3704_n 0.0287579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_294 VNB N_S[7]_c_3705_n 0.0296541f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_295 VNB N_S[7]_c_3706_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_296 VNB N_S[7]_c_3707_n 0.0214653f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_297 VNB N_S[7]_c_3708_n 0.0106587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_298 VNB N_S[7]_c_3709_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_299 VNB N_S[7]_c_3710_n 0.0254151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_300 VNB N_S[7]_c_3711_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_301 VNB N_S[7]_c_3712_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_302 VNB S[7] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_303 VNB N_S[15]_c_3766_n 0.0456684f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_304 VNB N_S[15]_c_3767_n 0.0296541f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_305 VNB N_S[15]_c_3768_n 0.0340051f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_306 VNB N_S[15]_c_3769_n 0.0214653f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_307 VNB N_S[15]_c_3770_n 0.0106587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_308 VNB N_S[15]_c_3771_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.295
cc_309 VNB N_S[15]_c_3772_n 0.0254151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_310 VNB N_S[15]_c_3773_n 0.014497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_311 VNB N_S[15]_c_3774_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_312 VNB S[15] 0.00576383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_313 VNB N_A_4565_47#_c_3832_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_314 VNB N_A_4565_47#_c_3833_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_315 VNB N_A_4565_47#_c_3834_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_316 VNB N_A_4565_47#_c_3835_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_317 VNB N_A_4565_937#_c_3912_n 0.014946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_318 VNB N_A_4565_937#_c_3913_n 0.00602901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_319 VNB N_A_4565_937#_c_3914_n 0.00871246f $X=-0.19 $Y=-0.24 $X2=0.52
+ $Y2=1.16
cc_320 VNB N_A_4565_937#_c_3915_n 0.00877362f $X=-0.19 $Y=-0.24 $X2=0.94
+ $Y2=1.16
cc_321 VNB N_D[7]_M1061_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_322 VNB N_D[7]_M1024_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_323 VNB N_D[7]_M1050_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_324 VNB N_D[7]_M1142_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_325 VNB D[7] 0.0128835f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_326 VNB N_D[7]_c_3997_n 0.0571683f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_327 VNB N_D[15]_M1068_g 5.5957e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_328 VNB N_D[15]_M1147_g 0.0189129f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_329 VNB N_D[15]_M1154_g 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_330 VNB N_D[15]_M1149_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_331 VNB D[15] 0.0128835f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_332 VNB N_D[15]_c_4047_n 0.0571683f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_333 VNB N_Z_c_5202_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_334 VNB N_Z_c_5203_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_335 VNB N_Z_c_5204_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_336 VNB N_Z_c_5205_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_337 VNB N_Z_c_5206_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_338 VNB N_Z_c_5207_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_339 VNB N_Z_c_5208_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_340 VNB N_Z_c_5209_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_341 VNB N_Z_c_5210_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_342 VNB N_Z_c_5211_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_343 VNB N_Z_c_5212_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_344 VNB N_Z_c_5213_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_345 VNB N_Z_c_5214_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_346 VNB N_Z_c_5215_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_347 VNB N_Z_c_5216_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_348 VNB N_Z_c_5217_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_349 VNB N_Z_c_5218_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_350 VNB N_Z_c_5219_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_351 VNB N_Z_c_5220_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_352 VNB N_Z_c_5221_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_353 VNB N_Z_c_5222_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_354 VNB N_Z_c_5223_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_355 VNB N_Z_c_5224_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_356 VNB N_Z_c_5225_n 0.00129655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_357 VNB N_Z_c_5226_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_358 VNB N_Z_c_5227_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_359 VNB N_Z_c_5228_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_360 VNB N_Z_c_5229_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_361 VNB N_Z_c_5230_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_362 VNB N_Z_c_5231_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_363 VNB N_Z_c_5232_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_364 VNB N_Z_c_5233_n 0.0103781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_365 VNB N_A_27_47#_c_7692_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_366 VNB N_A_27_47#_c_7693_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_367 VNB N_A_27_47#_c_7694_n 0.0034739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_368 VNB N_A_27_911#_c_7734_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_369 VNB N_A_27_911#_c_7735_n 0.0034739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_370 VNB N_A_27_911#_c_7736_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_371 VNB N_VGND_c_7777_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_372 VNB N_VGND_c_7778_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_373 VNB N_VGND_c_7779_n 0.00516508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_374 VNB N_VGND_c_7780_n 0.00516508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_375 VNB N_VGND_c_7781_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_376 VNB N_VGND_c_7782_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_377 VNB N_VGND_c_7783_n 0.0332577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_378 VNB N_VGND_c_7784_n 0.0332577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_379 VNB N_VGND_c_7785_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_380 VNB N_VGND_c_7786_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_381 VNB N_VGND_c_7787_n 0.00516508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_382 VNB N_VGND_c_7788_n 0.00516508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_383 VNB N_VGND_c_7789_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_384 VNB N_VGND_c_7790_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_385 VNB N_VGND_c_7791_n 0.0332577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_386 VNB N_VGND_c_7792_n 0.0332577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_387 VNB N_VGND_c_7793_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_388 VNB N_VGND_c_7794_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_389 VNB N_VGND_c_7795_n 0.00516508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_390 VNB N_VGND_c_7796_n 0.00516508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_391 VNB N_VGND_c_7797_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_392 VNB N_VGND_c_7798_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_393 VNB N_VGND_c_7799_n 0.0332577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_394 VNB N_VGND_c_7800_n 0.0332577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_395 VNB N_VGND_c_7801_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_396 VNB N_VGND_c_7802_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_397 VNB N_VGND_c_7803_n 0.00516508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_398 VNB N_VGND_c_7804_n 0.00516508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_399 VNB N_VGND_c_7805_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_400 VNB N_VGND_c_7806_n 0.00492504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_401 VNB N_VGND_c_7807_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_402 VNB N_VGND_c_7808_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_403 VNB N_VGND_c_7809_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_404 VNB N_VGND_c_7810_n 0.0047828f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_405 VNB N_VGND_c_7811_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_406 VNB N_VGND_c_7812_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_407 VNB N_VGND_c_7813_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_408 VNB N_VGND_c_7814_n 0.0047828f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_409 VNB N_VGND_c_7815_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_410 VNB N_VGND_c_7816_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_411 VNB N_VGND_c_7817_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_412 VNB N_VGND_c_7818_n 0.0047828f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_413 VNB N_VGND_c_7819_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_414 VNB N_VGND_c_7820_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_415 VNB N_VGND_c_7821_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_416 VNB N_VGND_c_7822_n 0.0047828f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_417 VNB N_VGND_c_7823_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_418 VNB N_VGND_c_7824_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_419 VNB N_VGND_c_7825_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_420 VNB N_VGND_c_7826_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_421 VNB VGND 1.17536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_422 VNB VGND 1.17536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_423 VNB N_VGND_c_7829_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_424 VNB N_VGND_c_7830_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_425 VNB N_VGND_c_7831_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_426 VNB N_VGND_c_7832_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_427 VNB N_VGND_c_7833_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_428 VNB N_VGND_c_7834_n 0.0556942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_429 VNB N_VGND_c_7835_n 0.0188039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_430 VNB N_VGND_c_7836_n 0.0188039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_431 VNB N_VGND_c_7837_n 0.0229085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_432 VNB N_VGND_c_7838_n 0.0229085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_433 VNB N_VGND_c_7839_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_434 VNB N_VGND_c_7840_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_435 VNB N_VGND_c_7841_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_436 VNB N_VGND_c_7842_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_437 VNB N_VGND_c_7843_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_438 VNB N_VGND_c_7844_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_439 VNB N_VGND_c_7845_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_440 VNB N_VGND_c_7846_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_441 VNB N_VGND_c_7847_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_442 VNB N_VGND_c_7848_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_443 VNB N_VGND_c_7849_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_444 VNB N_VGND_c_7850_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_445 VNB N_A_845_69#_c_8339_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_446 VNB N_A_845_69#_c_8340_n 0.00109213f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_447 VNB N_A_845_69#_c_8341_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_448 VNB N_A_845_69#_c_8342_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_449 VNB N_A_845_915#_c_8387_n 0.00256375f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_450 VNB N_A_845_915#_c_8388_n 0.00109213f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_451 VNB N_A_845_915#_c_8389_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_452 VNB N_A_845_915#_c_8390_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.75 $Y2=1.16
cc_453 VNB N_A_1315_47#_c_8434_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_454 VNB N_A_1315_47#_c_8435_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_455 VNB N_A_1315_47#_c_8436_n 0.0034739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_456 VNB N_A_1315_911#_c_8478_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_457 VNB N_A_1315_911#_c_8479_n 0.0034739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_458 VNB N_A_1315_911#_c_8480_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.495
+ $Y2=1.16
cc_459 VNB N_A_2133_69#_c_8522_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_460 VNB N_A_2133_69#_c_8523_n 0.00109213f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_461 VNB N_A_2133_69#_c_8524_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_462 VNB N_A_2133_69#_c_8525_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_463 VNB N_A_2133_915#_c_8570_n 0.00256375f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_464 VNB N_A_2133_915#_c_8571_n 0.00109213f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_465 VNB N_A_2133_915#_c_8572_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_466 VNB N_A_2133_915#_c_8573_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.75
+ $Y2=1.16
cc_467 VNB N_A_2603_47#_c_8617_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_468 VNB N_A_2603_47#_c_8618_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_469 VNB N_A_2603_47#_c_8619_n 0.0034739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_470 VNB N_A_2603_911#_c_8661_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_471 VNB N_A_2603_911#_c_8662_n 0.0034739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_472 VNB N_A_2603_911#_c_8663_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.495
+ $Y2=1.16
cc_473 VNB N_A_3421_69#_c_8705_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_474 VNB N_A_3421_69#_c_8706_n 0.00109213f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_475 VNB N_A_3421_69#_c_8707_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_476 VNB N_A_3421_69#_c_8708_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_477 VNB N_A_3421_915#_c_8753_n 0.00256375f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_478 VNB N_A_3421_915#_c_8754_n 0.00109213f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_479 VNB N_A_3421_915#_c_8755_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_480 VNB N_A_3421_915#_c_8756_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.75
+ $Y2=1.16
cc_481 VNB N_A_3891_47#_c_8800_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_482 VNB N_A_3891_47#_c_8801_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_483 VNB N_A_3891_47#_c_8802_n 0.0034739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_484 VNB N_A_3891_911#_c_8844_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_485 VNB N_A_3891_911#_c_8845_n 0.0034739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_486 VNB N_A_3891_911#_c_8846_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.495
+ $Y2=1.16
cc_487 VNB N_A_4709_69#_c_8888_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_488 VNB N_A_4709_69#_c_8889_n 0.00109213f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_489 VNB N_A_4709_69#_c_8890_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_490 VNB N_A_4709_69#_c_8891_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_491 VNB N_A_4709_915#_c_8934_n 0.00256375f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_492 VNB N_A_4709_915#_c_8935_n 0.00109213f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.985
cc_493 VNB N_A_4709_915#_c_8936_n 0.00682663f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_494 VNB N_A_4709_915#_c_8937_n 0.00179433f $X=-0.19 $Y=-0.24 $X2=0.75
+ $Y2=1.16
cc_495 VPB N_D[0]_M1010_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_496 VPB N_D[0]_M1075_g 0.0188543f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_497 VPB N_D[0]_c_852_n 0.00632455f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_498 VPB N_D[8]_M1014_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_499 VPB N_D[8]_M1078_g 0.0188543f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_500 VPB N_D[8]_c_903_n 0.00632455f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_501 VPB N_A_278_265#_M1013_g 0.0192795f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_502 VPB N_A_278_265#_c_956_n 0.0152663f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_503 VPB N_A_278_265#_c_957_n 0.0114291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_504 VPB N_A_278_265#_M1031_g 0.0225258f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_505 VPB N_A_278_265#_c_959_n 0.0076904f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_506 VPB N_A_278_265#_c_953_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_507 VPB N_A_278_265#_c_954_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_508 VPB N_A_278_793#_M1099_g 0.0192687f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_509 VPB N_A_278_793#_c_1039_n 0.0152663f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_510 VPB N_A_278_793#_c_1040_n 0.0114291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_511 VPB N_A_278_793#_M1111_g 0.022515f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_512 VPB N_A_278_793#_c_1036_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_513 VPB N_A_278_793#_c_1043_n 0.00768858f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_514 VPB N_A_278_793#_c_1037_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_515 VPB N_S[0]_c_1122_n 0.0253646f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_516 VPB N_S[8]_c_1191_n 0.0157866f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_517 VPB N_S[8]_c_1188_n 0.00957797f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_518 VPB N_S[1]_c_1247_n 0.0253646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_519 VPB N_S[9]_c_1309_n 0.00957797f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.295
cc_520 VPB N_S[9]_c_1320_n 0.0157866f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_521 VPB N_A_701_47#_M1084_g 0.0225258f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_522 VPB N_A_701_47#_c_1380_n 0.0265655f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_523 VPB N_A_701_47#_c_1375_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_524 VPB N_A_701_47#_M1113_g 0.0192795f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_525 VPB N_A_701_47#_c_1383_n 0.0076904f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_526 VPB N_A_701_47#_c_1378_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_527 VPB N_A_701_937#_M1036_g 0.022515f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_528 VPB N_A_701_937#_c_1461_n 0.0265655f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_529 VPB N_A_701_937#_c_1456_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_530 VPB N_A_701_937#_M1157_g 0.0192687f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_531 VPB N_A_701_937#_c_1464_n 0.00768858f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_532 VPB N_A_701_937#_c_1459_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_533 VPB N_D[1]_M1052_g 0.0188543f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_534 VPB N_D[1]_M1097_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_535 VPB D[1] 0.00525107f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_536 VPB N_D[9]_M1056_g 0.0188543f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_537 VPB N_D[9]_M1101_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_538 VPB D[9] 0.00525107f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_539 VPB N_D[2]_M1003_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_540 VPB N_D[2]_M1120_g 0.0188543f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_541 VPB N_D[2]_c_1655_n 0.00525107f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_542 VPB N_D[10]_M1009_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_543 VPB N_D[10]_M1126_g 0.0188543f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_544 VPB N_D[10]_c_1713_n 0.00525107f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_545 VPB N_A_1566_265#_M1005_g 0.0192795f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_546 VPB N_A_1566_265#_c_1773_n 0.0152663f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_547 VPB N_A_1566_265#_c_1774_n 0.0112992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_548 VPB N_A_1566_265#_M1124_g 0.0225258f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_549 VPB N_A_1566_265#_c_1776_n 0.0076904f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_550 VPB N_A_1566_265#_c_1770_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_551 VPB N_A_1566_265#_c_1771_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_552 VPB N_A_1566_793#_M1044_g 0.0192687f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_553 VPB N_A_1566_793#_c_1857_n 0.0152663f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_554 VPB N_A_1566_793#_c_1858_n 0.0112992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_555 VPB N_A_1566_793#_M1095_g 0.022515f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_556 VPB N_A_1566_793#_c_1854_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_557 VPB N_A_1566_793#_c_1861_n 0.00768858f $X=-0.19 $Y=1.305 $X2=0.41
+ $Y2=1.16
cc_558 VPB N_A_1566_793#_c_1855_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_559 VPB N_S[2]_c_1941_n 0.0253646f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_560 VPB N_S[10]_c_2010_n 0.0157866f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_561 VPB N_S[10]_c_2007_n 0.00957797f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_562 VPB N_S[3]_c_2066_n 0.0253646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_563 VPB N_S[11]_c_2128_n 0.00957797f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.295
cc_564 VPB N_S[11]_c_2139_n 0.0157866f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_565 VPB N_A_1989_47#_M1004_g 0.0225258f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_566 VPB N_A_1989_47#_c_2199_n 0.0265655f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_567 VPB N_A_1989_47#_c_2194_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_568 VPB N_A_1989_47#_M1123_g 0.0192795f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_569 VPB N_A_1989_47#_c_2202_n 0.0076904f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_570 VPB N_A_1989_47#_c_2197_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_571 VPB N_A_1989_937#_M1045_g 0.022515f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_572 VPB N_A_1989_937#_c_2280_n 0.0265655f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_573 VPB N_A_1989_937#_c_2275_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_574 VPB N_A_1989_937#_M1093_g 0.0192687f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_575 VPB N_A_1989_937#_c_2283_n 0.00768858f $X=-0.19 $Y=1.305 $X2=0.41
+ $Y2=1.16
cc_576 VPB N_A_1989_937#_c_2278_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_577 VPB N_D[3]_M1002_g 0.0188543f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_578 VPB N_D[3]_M1135_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_579 VPB D[3] 0.00525107f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_580 VPB N_D[11]_M1008_g 0.0188543f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_581 VPB N_D[11]_M1141_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_582 VPB D[11] 0.00525107f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_583 VPB N_D[4]_M1030_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_584 VPB N_D[4]_M1080_g 0.0188543f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_585 VPB N_D[4]_c_2474_n 0.00525107f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_586 VPB N_D[12]_M1038_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_587 VPB N_D[12]_M1088_g 0.0188543f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_588 VPB N_D[12]_c_2532_n 0.00525107f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_589 VPB N_A_2854_265#_M1034_g 0.0192795f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_590 VPB N_A_2854_265#_c_2592_n 0.0152663f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_591 VPB N_A_2854_265#_c_2593_n 0.0112992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_592 VPB N_A_2854_265#_M1083_g 0.0225258f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_593 VPB N_A_2854_265#_c_2595_n 0.0076904f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_594 VPB N_A_2854_265#_c_2589_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_595 VPB N_A_2854_265#_c_2590_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_596 VPB N_A_2854_793#_M1114_g 0.0192687f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_597 VPB N_A_2854_793#_c_2676_n 0.0152663f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_598 VPB N_A_2854_793#_c_2677_n 0.0112992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_599 VPB N_A_2854_793#_M1159_g 0.022515f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_600 VPB N_A_2854_793#_c_2673_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_601 VPB N_A_2854_793#_c_2680_n 0.00768858f $X=-0.19 $Y=1.305 $X2=0.41
+ $Y2=1.16
cc_602 VPB N_A_2854_793#_c_2674_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_603 VPB N_S[4]_c_2760_n 0.0253646f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_604 VPB N_S[12]_c_2829_n 0.0157866f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_605 VPB N_S[12]_c_2826_n 0.00957797f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_606 VPB N_S[5]_c_2885_n 0.0253646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_607 VPB N_S[13]_c_2947_n 0.00957797f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.295
cc_608 VPB N_S[13]_c_2958_n 0.0157866f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_609 VPB N_A_3277_47#_M1055_g 0.0225258f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_610 VPB N_A_3277_47#_c_3018_n 0.0265655f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_611 VPB N_A_3277_47#_c_3013_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_612 VPB N_A_3277_47#_M1082_g 0.0192795f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_613 VPB N_A_3277_47#_c_3021_n 0.0076904f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_614 VPB N_A_3277_47#_c_3016_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_615 VPB N_A_3277_937#_M1134_g 0.022515f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_616 VPB N_A_3277_937#_c_3099_n 0.0265655f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_617 VPB N_A_3277_937#_c_3094_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_618 VPB N_A_3277_937#_M1158_g 0.0192687f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_619 VPB N_A_3277_937#_c_3102_n 0.00768858f $X=-0.19 $Y=1.305 $X2=0.41
+ $Y2=1.16
cc_620 VPB N_A_3277_937#_c_3097_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_621 VPB N_D[5]_M1051_g 0.0188543f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_622 VPB N_D[5]_M1079_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_623 VPB D[5] 0.00525107f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_624 VPB N_D[13]_M1058_g 0.0188543f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_625 VPB N_D[13]_M1087_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_626 VPB D[13] 0.00525107f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_627 VPB N_D[6]_M1062_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_628 VPB N_D[6]_M1143_g 0.0188543f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_629 VPB N_D[6]_c_3293_n 0.00525107f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_630 VPB N_D[14]_M1069_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_631 VPB N_D[14]_M1152_g 0.0188543f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_632 VPB N_D[14]_c_3351_n 0.00525107f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_633 VPB N_A_4142_265#_M1066_g 0.0192795f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_634 VPB N_A_4142_265#_c_3411_n 0.0152663f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_635 VPB N_A_4142_265#_c_3412_n 0.0112992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_636 VPB N_A_4142_265#_M1091_g 0.0225258f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_637 VPB N_A_4142_265#_c_3414_n 0.0076904f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_638 VPB N_A_4142_265#_c_3408_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_639 VPB N_A_4142_265#_c_3409_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_640 VPB N_A_4142_793#_M1006_g 0.0192687f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_641 VPB N_A_4142_793#_c_3495_n 0.0152663f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_642 VPB N_A_4142_793#_c_3496_n 0.0112992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_643 VPB N_A_4142_793#_M1140_g 0.022515f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_644 VPB N_A_4142_793#_c_3492_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_645 VPB N_A_4142_793#_c_3499_n 0.00768858f $X=-0.19 $Y=1.305 $X2=0.41
+ $Y2=1.16
cc_646 VPB N_A_4142_793#_c_3493_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_647 VPB N_S[6]_c_3579_n 0.0253646f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_648 VPB N_S[14]_c_3648_n 0.0157866f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_649 VPB N_S[14]_c_3645_n 0.00957797f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_650 VPB N_S[7]_c_3704_n 0.0253646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_651 VPB N_S[15]_c_3766_n 0.00957797f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.295
cc_652 VPB N_S[15]_c_3777_n 0.0157866f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_653 VPB N_A_4565_47#_M1122_g 0.0225258f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_654 VPB N_A_4565_47#_c_3837_n 0.0266954f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_655 VPB N_A_4565_47#_c_3832_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_656 VPB N_A_4565_47#_M1148_g 0.0192795f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_657 VPB N_A_4565_47#_c_3840_n 0.0076904f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_658 VPB N_A_4565_47#_c_3835_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_659 VPB N_A_4565_937#_M1049_g 0.022515f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.025
cc_660 VPB N_A_4565_937#_c_3917_n 0.0266954f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_661 VPB N_A_4565_937#_c_3912_n 0.0320766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_662 VPB N_A_4565_937#_M1076_g 0.0192687f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_663 VPB N_A_4565_937#_c_3920_n 0.00768858f $X=-0.19 $Y=1.305 $X2=0.41
+ $Y2=1.16
cc_664 VPB N_A_4565_937#_c_3915_n 0.0134732f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_665 VPB N_D[7]_M1061_g 0.0188543f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_666 VPB N_D[7]_M1142_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_667 VPB D[7] 0.00632455f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_668 VPB N_D[15]_M1068_g 0.0188543f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_669 VPB N_D[15]_M1149_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_670 VPB D[15] 0.00632455f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_671 VPB N_A_27_297#_c_4092_n 0.0075508f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_672 VPB N_A_27_297#_c_4093_n 0.0101553f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.16
cc_673 VPB N_A_27_297#_c_4094_n 0.00205034f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.19
cc_674 VPB N_A_27_297#_c_4095_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_675 VPB N_A_27_297#_c_4096_n 0.0207852f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_676 VPB N_A_27_591#_c_4170_n 0.0207852f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.295
cc_677 VPB N_A_27_591#_c_4171_n 0.0075508f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_678 VPB N_A_27_591#_c_4172_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.16
cc_679 VPB N_A_27_591#_c_4173_n 0.00205034f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_680 VPB N_A_27_591#_c_4174_n 0.0101553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_681 VPB N_VPWR_c_4246_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_682 VPB N_VPWR_c_4247_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_683 VPB N_VPWR_c_4248_n 0.0147403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_684 VPB N_VPWR_c_4249_n 0.0147403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_685 VPB N_VPWR_c_4250_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_686 VPB N_VPWR_c_4251_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_687 VPB N_VPWR_c_4252_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_688 VPB N_VPWR_c_4253_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_689 VPB N_VPWR_c_4254_n 0.0147403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_690 VPB N_VPWR_c_4255_n 0.0147403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_691 VPB N_VPWR_c_4256_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_692 VPB N_VPWR_c_4257_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_693 VPB N_VPWR_c_4258_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_694 VPB N_VPWR_c_4259_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_695 VPB N_VPWR_c_4260_n 0.0147403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_696 VPB N_VPWR_c_4261_n 0.0147403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_697 VPB N_VPWR_c_4262_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_698 VPB N_VPWR_c_4263_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_699 VPB N_VPWR_c_4264_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_700 VPB N_VPWR_c_4265_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_701 VPB N_VPWR_c_4266_n 0.0147403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_702 VPB N_VPWR_c_4267_n 0.0147403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_703 VPB N_VPWR_c_4268_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_704 VPB N_VPWR_c_4269_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_705 VPB N_VPWR_c_4270_n 0.0232055f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_706 VPB N_VPWR_c_4271_n 0.00206903f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_707 VPB N_VPWR_c_4272_n 0.0232055f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_708 VPB N_VPWR_c_4273_n 0.00206903f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_709 VPB N_VPWR_c_4274_n 0.0232055f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_710 VPB N_VPWR_c_4275_n 0.00206903f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_711 VPB N_VPWR_c_4276_n 0.0232055f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_712 VPB N_VPWR_c_4277_n 0.00206903f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_713 VPB VPWR 0.134327f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_714 VPB N_VPWR_c_4279_n 0.0143733f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_715 VPB N_VPWR_c_4280_n 0.0102245f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_716 VPB N_VPWR_c_4281_n 0.0232055f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_717 VPB N_VPWR_c_4282_n 0.0102245f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_718 VPB N_VPWR_c_4283_n 0.0243964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_719 VPB N_VPWR_c_4284_n 0.0102245f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_720 VPB N_VPWR_c_4285_n 0.0232055f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_721 VPB N_VPWR_c_4286_n 0.0102245f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_722 VPB N_VPWR_c_4287_n 0.0243964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_723 VPB N_VPWR_c_4288_n 0.0102245f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_724 VPB N_VPWR_c_4289_n 0.0232055f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_725 VPB N_VPWR_c_4290_n 0.0102245f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_726 VPB N_VPWR_c_4291_n 0.0243964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_727 VPB N_VPWR_c_4292_n 0.0102245f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_728 VPB N_VPWR_c_4293_n 0.0232055f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_729 VPB N_VPWR_c_4294_n 0.0102245f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_730 VPB N_VPWR_c_4295_n 0.0143733f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_731 VPB N_VPWR_c_4296_n 6.22115e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_732 VPB N_VPWR_c_4297_n 6.22115e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_733 VPB N_VPWR_c_4298_n 6.22115e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_734 VPB N_VPWR_c_4299_n 6.22115e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_735 VPB N_VPWR_c_4300_n 6.22115e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_736 VPB N_VPWR_c_4301_n 6.22115e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_737 VPB N_VPWR_c_4302_n 6.22115e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_738 VPB N_VPWR_c_4303_n 6.22115e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_739 VPB N_Z_c_5202_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_740 VPB N_Z_c_5203_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_741 VPB N_Z_c_5204_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_742 VPB N_Z_c_5205_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_743 VPB N_Z_c_5206_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_744 VPB N_Z_c_5207_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_745 VPB N_Z_c_5208_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_746 VPB N_Z_c_5209_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_747 VPB N_Z_c_5242_n 0.0096248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_748 VPB N_Z_c_5243_n 0.0096248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_749 VPB N_Z_c_5244_n 0.00920862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_750 VPB N_Z_c_5245_n 0.00920862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_751 VPB N_Z_c_5246_n 0.0096248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_752 VPB N_Z_c_5247_n 0.0096248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_753 VPB N_Z_c_5248_n 0.00920862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_754 VPB N_Z_c_5249_n 0.00920862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_755 VPB N_Z_c_5250_n 0.0096248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_756 VPB N_Z_c_5251_n 0.0096248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_757 VPB N_Z_c_5252_n 0.00920862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_758 VPB N_Z_c_5253_n 0.00920862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_759 VPB N_Z_c_5254_n 0.0096248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_760 VPB N_Z_c_5255_n 0.0096248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_761 VPB N_Z_c_5226_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_762 VPB N_Z_c_5257_n 0.0115657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_763 VPB N_Z_c_5227_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_764 VPB N_Z_c_5259_n 0.0115657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_765 VPB N_Z_c_5228_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_766 VPB N_Z_c_5261_n 0.0115657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_767 VPB N_Z_c_5229_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_768 VPB N_Z_c_5263_n 0.0115657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_769 VPB N_Z_c_5230_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_770 VPB N_Z_c_5265_n 0.0115657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_771 VPB N_Z_c_5231_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_772 VPB N_Z_c_5267_n 0.0115657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_773 VPB N_Z_c_5232_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_774 VPB N_Z_c_5269_n 0.0115657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_775 VPB N_Z_c_5233_n 0.00348015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_776 VPB N_Z_c_5271_n 0.0115657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_777 VPB N_A_824_333#_c_6418_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_778 VPB N_A_824_333#_c_6419_n 0.00205034f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_779 VPB N_A_824_333#_c_6420_n 0.00239382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_780 VPB N_A_824_333#_c_6421_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_781 VPB N_A_824_333#_c_6422_n 0.0042022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_782 VPB N_A_824_591#_c_6514_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_783 VPB N_A_824_591#_c_6515_n 0.0042022f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_784 VPB N_A_824_591#_c_6516_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_785 VPB N_A_824_591#_c_6517_n 0.00205034f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_786 VPB N_A_824_591#_c_6518_n 0.00239382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_787 VPB N_A_1315_297#_c_6605_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=0.56
cc_788 VPB N_A_1315_297#_c_6606_n 0.00239382f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.16
cc_789 VPB N_A_1315_297#_c_6607_n 0.00205034f $X=-0.19 $Y=1.305 $X2=0.75
+ $Y2=1.19
cc_790 VPB N_A_1315_297#_c_6608_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_791 VPB N_A_1315_297#_c_6609_n 0.0042022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_792 VPB N_A_1315_591#_c_6699_n 0.0042022f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.295
cc_793 VPB N_A_1315_591#_c_6700_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_794 VPB N_A_1315_591#_c_6701_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.16
cc_795 VPB N_A_1315_591#_c_6702_n 0.00205034f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_796 VPB N_A_1315_591#_c_6703_n 0.00239382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_797 VPB N_A_2112_333#_c_6791_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_798 VPB N_A_2112_333#_c_6792_n 0.00205034f $X=-0.19 $Y=1.305 $X2=0.52
+ $Y2=1.16
cc_799 VPB N_A_2112_333#_c_6793_n 0.00239382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_800 VPB N_A_2112_333#_c_6794_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_801 VPB N_A_2112_333#_c_6795_n 0.0042022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_802 VPB N_A_2112_591#_c_6887_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=0.56
cc_803 VPB N_A_2112_591#_c_6888_n 0.0042022f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_804 VPB N_A_2112_591#_c_6889_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_805 VPB N_A_2112_591#_c_6890_n 0.00205034f $X=-0.19 $Y=1.305 $X2=0.75
+ $Y2=1.16
cc_806 VPB N_A_2112_591#_c_6891_n 0.00239382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_807 VPB N_A_2603_297#_c_6978_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=0.56
cc_808 VPB N_A_2603_297#_c_6979_n 0.00239382f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.16
cc_809 VPB N_A_2603_297#_c_6980_n 0.00205034f $X=-0.19 $Y=1.305 $X2=0.75
+ $Y2=1.19
cc_810 VPB N_A_2603_297#_c_6981_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_811 VPB N_A_2603_297#_c_6982_n 0.0042022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_812 VPB N_A_2603_591#_c_7072_n 0.0042022f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.295
cc_813 VPB N_A_2603_591#_c_7073_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_814 VPB N_A_2603_591#_c_7074_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.16
cc_815 VPB N_A_2603_591#_c_7075_n 0.00205034f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_816 VPB N_A_2603_591#_c_7076_n 0.00239382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_817 VPB N_A_3400_333#_c_7164_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_818 VPB N_A_3400_333#_c_7165_n 0.00205034f $X=-0.19 $Y=1.305 $X2=0.52
+ $Y2=1.16
cc_819 VPB N_A_3400_333#_c_7166_n 0.00239382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_820 VPB N_A_3400_333#_c_7167_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_821 VPB N_A_3400_333#_c_7168_n 0.0042022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_822 VPB N_A_3400_591#_c_7260_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=0.56
cc_823 VPB N_A_3400_591#_c_7261_n 0.0042022f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_824 VPB N_A_3400_591#_c_7262_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_825 VPB N_A_3400_591#_c_7263_n 0.00205034f $X=-0.19 $Y=1.305 $X2=0.75
+ $Y2=1.16
cc_826 VPB N_A_3400_591#_c_7264_n 0.00239382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_827 VPB N_A_3891_297#_c_7351_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=0.56
cc_828 VPB N_A_3891_297#_c_7352_n 0.00239382f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.16
cc_829 VPB N_A_3891_297#_c_7353_n 0.00205034f $X=-0.19 $Y=1.305 $X2=0.75
+ $Y2=1.19
cc_830 VPB N_A_3891_297#_c_7354_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_831 VPB N_A_3891_297#_c_7355_n 0.0042022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_832 VPB N_A_3891_591#_c_7445_n 0.0042022f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.295
cc_833 VPB N_A_3891_591#_c_7446_n 0.00189928f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_834 VPB N_A_3891_591#_c_7447_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.16
cc_835 VPB N_A_3891_591#_c_7448_n 0.00205034f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_836 VPB N_A_3891_591#_c_7449_n 0.00239382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_837 VPB N_A_4688_333#_c_7537_n 0.0075508f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_838 VPB N_A_4688_333#_c_7538_n 0.00205034f $X=-0.19 $Y=1.305 $X2=0.52
+ $Y2=1.16
cc_839 VPB N_A_4688_333#_c_7539_n 0.0101553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_840 VPB N_A_4688_333#_c_7540_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_841 VPB N_A_4688_333#_c_7541_n 0.0207852f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_842 VPB N_A_4688_591#_c_7617_n 0.0075508f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_843 VPB N_A_4688_591#_c_7618_n 0.0207852f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_844 VPB N_A_4688_591#_c_7619_n 0.00141501f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_845 VPB N_A_4688_591#_c_7620_n 0.00205034f $X=-0.19 $Y=1.305 $X2=0.75
+ $Y2=1.16
cc_846 VPB N_A_4688_591#_c_7621_n 0.0101553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_847 N_D[0]_M1010_g N_D[8]_M1014_g 0.0130744f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_848 N_D[0]_M1075_g N_D[8]_M1078_g 0.0129371f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_849 N_D[0]_M1075_g N_A_278_265#_M1013_g 0.0241487f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_850 N_D[0]_M1075_g N_A_278_265#_c_957_n 0.00671996f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_851 N_D[0]_M1108_g N_S[0]_c_1116_n 0.0165585f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_852 N_D[0]_c_852_n N_A_27_297#_c_4092_n 0.0235932f $X=0.75 $Y=1.16 $X2=0
+ $Y2=0
cc_853 N_D[0]_c_853_n N_A_27_297#_c_4092_n 9.6385e-19 $X=0.965 $Y=1.16 $X2=0
+ $Y2=0
cc_854 N_D[0]_M1010_g N_A_27_297#_c_4099_n 0.0111151f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_855 N_D[0]_M1075_g N_A_27_297#_c_4099_n 0.0138742f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_856 N_D[0]_c_852_n N_A_27_297#_c_4099_n 0.0339353f $X=0.75 $Y=1.16 $X2=0
+ $Y2=0
cc_857 N_D[0]_c_853_n N_A_27_297#_c_4099_n 7.13708e-19 $X=0.965 $Y=1.16 $X2=0
+ $Y2=0
cc_858 N_D[0]_M1010_g N_A_27_297#_c_4103_n 0.00332247f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_859 N_D[0]_M1075_g N_A_27_297#_c_4103_n 0.00330676f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_860 N_D[0]_M1010_g N_A_27_297#_c_4093_n 0.00290175f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_861 N_D[0]_M1075_g N_A_27_297#_c_4106_n 0.00611417f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_862 N_D[0]_M1010_g N_VPWR_c_4246_n 0.00338721f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_863 N_D[0]_M1075_g N_VPWR_c_4246_n 0.00848021f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_864 N_D[0]_M1010_g N_VPWR_c_4306_n 0.00359955f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_865 N_D[0]_M1075_g N_VPWR_c_4306_n 0.00343746f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_866 N_D[0]_M1010_g VPWR 0.00531592f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_867 N_D[0]_M1075_g VPWR 0.00350923f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_868 N_D[0]_M1010_g N_VPWR_c_4279_n 0.0033767f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_869 N_D[0]_M1075_g N_VPWR_c_4280_n 0.00342413f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_870 N_D[0]_M1108_g N_Z_c_5226_n 8.13311e-19 $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_871 N_D[0]_M1075_g N_Z_c_5226_n 0.00112534f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_872 N_D[0]_c_852_n N_Z_c_5226_n 0.00742792f $X=0.75 $Y=1.16 $X2=0 $Y2=0
cc_873 N_D[0]_c_853_n N_Z_c_5226_n 0.00583073f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_874 N_D[0]_M1042_g N_A_27_47#_c_7695_n 0.00633603f $X=0.52 $Y=0.56 $X2=0
+ $Y2=0
cc_875 N_D[0]_M1108_g N_A_27_47#_c_7695_n 5.29024e-19 $X=0.94 $Y=0.56 $X2=0
+ $Y2=0
cc_876 N_D[0]_M1042_g N_A_27_47#_c_7692_n 0.0084485f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_877 N_D[0]_M1108_g N_A_27_47#_c_7692_n 0.0125955f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_878 N_D[0]_c_852_n N_A_27_47#_c_7692_n 0.0274027f $X=0.75 $Y=1.16 $X2=0 $Y2=0
cc_879 N_D[0]_c_853_n N_A_27_47#_c_7692_n 0.00321151f $X=0.965 $Y=1.16 $X2=0
+ $Y2=0
cc_880 N_D[0]_M1042_g N_A_27_47#_c_7693_n 8.68782e-19 $X=0.52 $Y=0.56 $X2=0
+ $Y2=0
cc_881 N_D[0]_c_852_n N_A_27_47#_c_7693_n 0.024456f $X=0.75 $Y=1.16 $X2=0 $Y2=0
cc_882 N_D[0]_c_853_n N_A_27_47#_c_7693_n 0.00464565f $X=0.965 $Y=1.16 $X2=0
+ $Y2=0
cc_883 N_D[0]_M1042_g N_VGND_c_7777_n 0.0030929f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_884 N_D[0]_M1108_g N_VGND_c_7777_n 0.00300333f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_885 N_D[0]_M1108_g N_VGND_c_7807_n 0.00436487f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_886 N_D[0]_M1042_g VGND 0.00697949f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_887 N_D[0]_M1108_g VGND 0.00600262f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_888 N_D[0]_M1042_g N_VGND_c_7837_n 0.00430643f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_889 N_D[8]_M1078_g N_A_278_793#_M1099_g 0.0241475f $X=0.965 $Y=3.455 $X2=0
+ $Y2=0
cc_890 N_D[8]_M1078_g N_A_278_793#_c_1040_n 0.00671996f $X=0.965 $Y=3.455 $X2=0
+ $Y2=0
cc_891 N_D[8]_M1118_g N_S[8]_c_1180_n 0.0165585f $X=0.94 $Y=4.88 $X2=-0.19
+ $Y2=-0.24
cc_892 N_D[8]_M1014_g N_A_27_591#_c_4175_n 0.0111151f $X=0.495 $Y=3.455 $X2=0
+ $Y2=0
cc_893 N_D[8]_M1078_g N_A_27_591#_c_4175_n 0.0138742f $X=0.965 $Y=3.455 $X2=0
+ $Y2=0
cc_894 N_D[8]_c_903_n N_A_27_591#_c_4175_n 0.0339353f $X=0.75 $Y=4.28 $X2=0
+ $Y2=0
cc_895 N_D[8]_c_904_n N_A_27_591#_c_4175_n 7.13708e-19 $X=0.965 $Y=4.28 $X2=0
+ $Y2=0
cc_896 N_D[8]_c_903_n N_A_27_591#_c_4171_n 0.0235932f $X=0.75 $Y=4.28 $X2=0
+ $Y2=0
cc_897 N_D[8]_c_904_n N_A_27_591#_c_4171_n 9.6385e-19 $X=0.965 $Y=4.28 $X2=0
+ $Y2=0
cc_898 N_D[8]_M1014_g N_A_27_591#_c_4181_n 0.00332247f $X=0.495 $Y=3.455 $X2=0
+ $Y2=0
cc_899 N_D[8]_M1078_g N_A_27_591#_c_4181_n 0.00330232f $X=0.965 $Y=3.455 $X2=0
+ $Y2=0
cc_900 N_D[8]_M1078_g N_A_27_591#_c_4183_n 0.00548019f $X=0.965 $Y=3.455 $X2=0
+ $Y2=0
cc_901 N_D[8]_M1014_g N_A_27_591#_c_4174_n 0.00290175f $X=0.495 $Y=3.455 $X2=0
+ $Y2=0
cc_902 N_D[8]_M1014_g N_VPWR_c_4247_n 0.00338721f $X=0.495 $Y=3.455 $X2=0 $Y2=0
cc_903 N_D[8]_M1078_g N_VPWR_c_4247_n 0.00847423f $X=0.965 $Y=3.455 $X2=0 $Y2=0
cc_904 N_D[8]_M1014_g N_VPWR_c_4314_n 0.00359955f $X=0.495 $Y=3.455 $X2=0 $Y2=0
cc_905 N_D[8]_M1078_g N_VPWR_c_4314_n 0.00343746f $X=0.965 $Y=3.455 $X2=0 $Y2=0
cc_906 N_D[8]_M1014_g VPWR 0.00531592f $X=0.495 $Y=3.455 $X2=0 $Y2=0
cc_907 N_D[8]_M1078_g VPWR 0.00350923f $X=0.965 $Y=3.455 $X2=0 $Y2=0
cc_908 N_D[8]_M1014_g N_VPWR_c_4279_n 0.0033767f $X=0.495 $Y=3.455 $X2=0 $Y2=0
cc_909 N_D[8]_M1078_g N_VPWR_c_4280_n 0.00342413f $X=0.965 $Y=3.455 $X2=0 $Y2=0
cc_910 N_D[8]_M1118_g N_Z_c_5202_n 8.13311e-19 $X=0.94 $Y=4.88 $X2=0 $Y2=0
cc_911 N_D[8]_M1078_g N_Z_c_5202_n 0.00112534f $X=0.965 $Y=3.455 $X2=0 $Y2=0
cc_912 N_D[8]_c_903_n N_Z_c_5202_n 0.00742792f $X=0.75 $Y=4.28 $X2=0 $Y2=0
cc_913 N_D[8]_c_904_n N_Z_c_5202_n 0.00583073f $X=0.965 $Y=4.28 $X2=0 $Y2=0
cc_914 N_D[8]_M1047_g N_A_27_911#_c_7737_n 0.0084485f $X=0.52 $Y=4.88 $X2=0
+ $Y2=0
cc_915 N_D[8]_M1118_g N_A_27_911#_c_7737_n 0.0114493f $X=0.94 $Y=4.88 $X2=0
+ $Y2=0
cc_916 N_D[8]_c_903_n N_A_27_911#_c_7737_n 0.0274027f $X=0.75 $Y=4.28 $X2=0
+ $Y2=0
cc_917 N_D[8]_c_904_n N_A_27_911#_c_7737_n 0.0020061f $X=0.965 $Y=4.28 $X2=0
+ $Y2=0
cc_918 N_D[8]_M1118_g N_A_27_911#_c_7734_n 0.00114614f $X=0.94 $Y=4.88 $X2=0
+ $Y2=0
cc_919 N_D[8]_c_904_n N_A_27_911#_c_7734_n 0.00120541f $X=0.965 $Y=4.28 $X2=0
+ $Y2=0
cc_920 N_D[8]_M1047_g N_A_27_911#_c_7736_n 0.00720482f $X=0.52 $Y=4.88 $X2=0
+ $Y2=0
cc_921 N_D[8]_M1118_g N_A_27_911#_c_7736_n 5.29024e-19 $X=0.94 $Y=4.88 $X2=0
+ $Y2=0
cc_922 N_D[8]_c_903_n N_A_27_911#_c_7736_n 0.024456f $X=0.75 $Y=4.28 $X2=0 $Y2=0
cc_923 N_D[8]_c_904_n N_A_27_911#_c_7736_n 0.00464565f $X=0.965 $Y=4.28 $X2=0
+ $Y2=0
cc_924 N_D[8]_M1047_g N_VGND_c_7778_n 0.0030929f $X=0.52 $Y=4.88 $X2=0 $Y2=0
cc_925 N_D[8]_M1118_g N_VGND_c_7778_n 0.00300333f $X=0.94 $Y=4.88 $X2=0 $Y2=0
cc_926 N_D[8]_M1118_g N_VGND_c_7809_n 0.00436487f $X=0.94 $Y=4.88 $X2=0 $Y2=0
cc_927 N_D[8]_M1047_g VGND 0.00697949f $X=0.52 $Y=4.88 $X2=0 $Y2=0
cc_928 N_D[8]_M1118_g VGND 0.00600262f $X=0.94 $Y=4.88 $X2=0 $Y2=0
cc_929 N_D[8]_M1047_g N_VGND_c_7838_n 0.00430643f $X=0.52 $Y=4.88 $X2=0 $Y2=0
cc_930 N_A_278_265#_M1013_g N_A_278_793#_M1099_g 0.0130744f $X=1.49 $Y=2.075
+ $X2=0 $Y2=0
cc_931 N_A_278_265#_M1031_g N_A_278_793#_M1111_g 0.0130744f $X=1.96 $Y=2.075
+ $X2=0 $Y2=0
cc_932 N_A_278_265#_c_957_n N_S[0]_c_1114_n 0.00779314f $X=1.58 $Y=1.4 $X2=-0.19
+ $Y2=-0.24
cc_933 N_A_278_265#_c_956_n N_S[0]_c_1117_n 0.00810157f $X=1.87 $Y=1.4 $X2=0
+ $Y2=0
cc_934 N_A_278_265#_c_952_n N_S[0]_c_1117_n 7.04048e-19 $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_935 N_A_278_265#_c_951_n N_S[0]_c_1119_n 0.0100587f $X=2.43 $Y=0.755 $X2=0
+ $Y2=0
cc_936 N_A_278_265#_c_952_n N_S[0]_c_1119_n 0.00267287f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_937 N_A_278_265#_c_951_n N_S[0]_c_1120_n 0.0105766f $X=2.43 $Y=0.755 $X2=0
+ $Y2=0
cc_938 N_A_278_265#_c_952_n N_S[0]_c_1120_n 0.0090765f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_939 N_A_278_265#_c_953_n N_S[0]_c_1120_n 0.00742826f $X=2.715 $Y=1.63 $X2=0
+ $Y2=0
cc_940 N_A_278_265#_c_952_n N_S[0]_c_1121_n 0.00445422f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_941 N_A_278_265#_c_953_n N_S[0]_c_1121_n 4.25171e-19 $X=2.715 $Y=1.63 $X2=0
+ $Y2=0
cc_942 N_A_278_265#_c_954_n N_S[0]_c_1121_n 0.00920672f $X=1.96 $Y=1.34 $X2=0
+ $Y2=0
cc_943 N_A_278_265#_c_952_n N_S[0]_c_1122_n 0.00205356f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_944 N_A_278_265#_c_959_n N_S[0]_c_1122_n 0.00861299f $X=2.715 $Y=2.31 $X2=0
+ $Y2=0
cc_945 N_A_278_265#_c_953_n N_S[0]_c_1122_n 0.00828481f $X=2.715 $Y=1.63 $X2=0
+ $Y2=0
cc_946 N_A_278_265#_c_954_n N_S[0]_c_1122_n 0.00692516f $X=1.96 $Y=1.34 $X2=0
+ $Y2=0
cc_947 N_A_278_265#_c_952_n N_S[0]_c_1123_n 0.00149517f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_948 N_A_278_265#_c_951_n S[0] 0.0061421f $X=2.43 $Y=0.755 $X2=0 $Y2=0
cc_949 N_A_278_265#_c_952_n S[0] 0.0101733f $X=2.43 $Y=1.205 $X2=0 $Y2=0
cc_950 N_A_278_265#_c_953_n S[0] 0.0127184f $X=2.715 $Y=1.63 $X2=0 $Y2=0
cc_951 N_A_278_265#_c_954_n S[0] 3.07062e-19 $X=1.96 $Y=1.34 $X2=0 $Y2=0
cc_952 N_A_278_265#_M1013_g N_A_27_297#_c_4099_n 0.00176121f $X=1.49 $Y=2.075
+ $X2=0 $Y2=0
cc_953 N_A_278_265#_M1013_g N_A_27_297#_c_4108_n 0.00663284f $X=1.49 $Y=2.075
+ $X2=0 $Y2=0
cc_954 N_A_278_265#_M1031_g N_A_27_297#_c_4108_n 0.00334959f $X=1.96 $Y=2.075
+ $X2=0 $Y2=0
cc_955 N_A_278_265#_M1013_g N_A_27_297#_c_4110_n 7.75952e-19 $X=1.49 $Y=2.075
+ $X2=0 $Y2=0
cc_956 N_A_278_265#_M1013_g N_A_27_297#_c_4111_n 0.00415998f $X=1.49 $Y=2.075
+ $X2=0 $Y2=0
cc_957 N_A_278_265#_c_959_n N_A_27_297#_c_4094_n 0.00738363f $X=2.715 $Y=2.31
+ $X2=0 $Y2=0
cc_958 N_A_278_265#_M1031_g N_A_27_297#_c_4113_n 0.00692695f $X=1.96 $Y=2.075
+ $X2=0 $Y2=0
cc_959 N_A_278_265#_M1013_g N_A_27_297#_c_4106_n 0.00527462f $X=1.49 $Y=2.075
+ $X2=0 $Y2=0
cc_960 N_A_278_265#_M1031_g N_A_27_297#_c_4095_n 0.00550198f $X=1.96 $Y=2.075
+ $X2=0 $Y2=0
cc_961 N_A_278_265#_c_959_n N_A_27_297#_c_4095_n 0.0413447f $X=2.715 $Y=2.31
+ $X2=0 $Y2=0
cc_962 N_A_278_265#_c_953_n N_A_27_297#_c_4095_n 0.0132748f $X=2.715 $Y=1.63
+ $X2=0 $Y2=0
cc_963 N_A_278_265#_c_954_n N_A_27_297#_c_4095_n 0.00133381f $X=1.96 $Y=1.34
+ $X2=0 $Y2=0
cc_964 N_A_278_265#_M1013_g N_VPWR_c_4246_n 0.00107878f $X=1.49 $Y=2.075 $X2=0
+ $Y2=0
cc_965 N_A_278_265#_c_959_n N_VPWR_c_4248_n 0.0321301f $X=2.715 $Y=2.31 $X2=0
+ $Y2=0
cc_966 N_A_278_265#_c_953_n N_VPWR_c_4248_n 0.00732952f $X=2.715 $Y=1.63 $X2=0
+ $Y2=0
cc_967 N_A_278_265#_M1031_g N_VPWR_c_4270_n 8.06528e-19 $X=1.96 $Y=2.075 $X2=0
+ $Y2=0
cc_968 N_A_278_265#_c_959_n N_VPWR_c_4270_n 0.0210596f $X=2.715 $Y=2.31 $X2=0
+ $Y2=0
cc_969 N_A_278_265#_M1023_s VPWR 0.00179197f $X=2.59 $Y=1.485 $X2=0 $Y2=0
cc_970 N_A_278_265#_M1013_g VPWR 0.00435072f $X=1.49 $Y=2.075 $X2=0 $Y2=0
cc_971 N_A_278_265#_M1031_g VPWR 0.0054792f $X=1.96 $Y=2.075 $X2=0 $Y2=0
cc_972 N_A_278_265#_c_959_n VPWR 0.00594162f $X=2.715 $Y=2.31 $X2=0 $Y2=0
cc_973 N_A_278_265#_c_956_n N_Z_c_5210_n 0.00168443f $X=1.87 $Y=1.4 $X2=0 $Y2=0
cc_974 N_A_278_265#_c_957_n N_Z_c_5210_n 0.00180308f $X=1.58 $Y=1.4 $X2=0 $Y2=0
cc_975 N_A_278_265#_c_952_n N_Z_c_5210_n 0.0033343f $X=2.43 $Y=1.205 $X2=0 $Y2=0
cc_976 N_A_278_265#_M1031_g N_Z_c_5242_n 0.00708998f $X=1.96 $Y=2.075 $X2=0
+ $Y2=0
cc_977 N_A_278_265#_c_959_n N_Z_c_5242_n 0.0308332f $X=2.715 $Y=2.31 $X2=0 $Y2=0
cc_978 N_A_278_265#_c_953_n N_Z_c_5242_n 0.0132841f $X=2.715 $Y=1.63 $X2=0 $Y2=0
cc_979 N_A_278_265#_c_954_n N_Z_c_5242_n 9.57301e-19 $X=1.96 $Y=1.34 $X2=0 $Y2=0
cc_980 N_A_278_265#_M1013_g N_Z_c_5287_n 0.00635853f $X=1.49 $Y=2.075 $X2=0
+ $Y2=0
cc_981 N_A_278_265#_M1013_g N_Z_c_5288_n 0.00978858f $X=1.49 $Y=2.075 $X2=0
+ $Y2=0
cc_982 N_A_278_265#_c_956_n N_Z_c_5288_n 8.37785e-19 $X=1.87 $Y=1.4 $X2=0 $Y2=0
cc_983 N_A_278_265#_M1031_g N_Z_c_5288_n 0.00619657f $X=1.96 $Y=2.075 $X2=0
+ $Y2=0
cc_984 N_A_278_265#_M1013_g N_Z_c_5226_n 0.00268051f $X=1.49 $Y=2.075 $X2=0
+ $Y2=0
cc_985 N_A_278_265#_c_956_n N_Z_c_5226_n 0.0140957f $X=1.87 $Y=1.4 $X2=0 $Y2=0
cc_986 N_A_278_265#_M1031_g N_Z_c_5226_n 0.00476154f $X=1.96 $Y=2.075 $X2=0
+ $Y2=0
cc_987 N_A_278_265#_c_952_n N_Z_c_5226_n 0.00967956f $X=2.43 $Y=1.205 $X2=0
+ $Y2=0
cc_988 N_A_278_265#_c_953_n N_Z_c_5226_n 0.0117695f $X=2.715 $Y=1.63 $X2=0 $Y2=0
cc_989 N_A_278_265#_c_954_n N_Z_c_5226_n 7.26438e-19 $X=1.96 $Y=1.34 $X2=0 $Y2=0
cc_990 N_A_278_265#_M1013_g N_Z_c_5297_n 2.61869e-19 $X=1.49 $Y=2.075 $X2=0
+ $Y2=0
cc_991 N_A_278_265#_M1013_g N_Z_c_5257_n 0.00455034f $X=1.49 $Y=2.075 $X2=0
+ $Y2=0
cc_992 N_A_278_265#_M1031_g N_Z_c_5257_n 0.00462462f $X=1.96 $Y=2.075 $X2=0
+ $Y2=0
cc_993 N_A_278_265#_c_951_n N_A_27_47#_c_7694_n 0.00358194f $X=2.43 $Y=0.755
+ $X2=0 $Y2=0
cc_994 N_A_278_265#_c_951_n N_A_27_47#_c_7705_n 0.0185512f $X=2.43 $Y=0.755
+ $X2=0 $Y2=0
cc_995 N_A_278_265#_c_952_n N_A_27_47#_c_7705_n 0.00101918f $X=2.43 $Y=1.205
+ $X2=0 $Y2=0
cc_996 N_A_278_265#_c_953_n N_A_27_47#_c_7705_n 0.00285813f $X=2.715 $Y=1.63
+ $X2=0 $Y2=0
cc_997 N_A_278_265#_c_954_n N_A_27_47#_c_7705_n 0.00308807f $X=1.96 $Y=1.34
+ $X2=0 $Y2=0
cc_998 N_A_278_265#_c_951_n N_VGND_c_7807_n 0.0173492f $X=2.43 $Y=0.755 $X2=0
+ $Y2=0
cc_999 N_A_278_265#_M1081_s VGND 0.00250855f $X=2.675 $Y=0.235 $X2=0 $Y2=0
cc_1000 N_A_278_265#_c_951_n VGND 0.0186564f $X=2.43 $Y=0.755 $X2=0 $Y2=0
cc_1001 N_A_278_793#_c_1040_n N_S[8]_c_1180_n 0.00779314f $X=1.58 $Y=4.04
+ $X2=-0.19 $Y2=-0.24
cc_1002 N_A_278_793#_c_1039_n N_S[8]_c_1183_n 0.00810157f $X=1.87 $Y=4.04 $X2=0
+ $Y2=0
cc_1003 N_A_278_793#_c_1035_n N_S[8]_c_1183_n 7.04048e-19 $X=2.43 $Y=4.685 $X2=0
+ $Y2=0
cc_1004 N_A_278_793#_c_1035_n N_S[8]_c_1185_n 0.0127103f $X=2.43 $Y=4.685 $X2=0
+ $Y2=0
cc_1005 N_A_278_793#_c_1035_n N_S[8]_c_1186_n 0.0196531f $X=2.43 $Y=4.685 $X2=0
+ $Y2=0
cc_1006 N_A_278_793#_c_1036_n N_S[8]_c_1186_n 0.00742826f $X=2.715 $Y=3.805
+ $X2=0 $Y2=0
cc_1007 N_A_278_793#_c_1035_n N_S[8]_c_1187_n 0.00445422f $X=2.43 $Y=4.685 $X2=0
+ $Y2=0
cc_1008 N_A_278_793#_c_1036_n N_S[8]_c_1187_n 4.25171e-19 $X=2.715 $Y=3.805
+ $X2=0 $Y2=0
cc_1009 N_A_278_793#_c_1037_n N_S[8]_c_1187_n 0.00920672f $X=1.96 $Y=4.1 $X2=0
+ $Y2=0
cc_1010 N_A_278_793#_c_1036_n N_S[8]_c_1191_n 0.00386817f $X=2.715 $Y=3.805
+ $X2=0 $Y2=0
cc_1011 N_A_278_793#_c_1043_n N_S[8]_c_1191_n 0.00861299f $X=2.715 $Y=3.13 $X2=0
+ $Y2=0
cc_1012 N_A_278_793#_c_1037_n N_S[8]_c_1191_n 0.00149275f $X=1.96 $Y=4.1 $X2=0
+ $Y2=0
cc_1013 N_A_278_793#_c_1035_n N_S[8]_c_1188_n 0.00354873f $X=2.43 $Y=4.685 $X2=0
+ $Y2=0
cc_1014 N_A_278_793#_c_1036_n N_S[8]_c_1188_n 0.00441664f $X=2.715 $Y=3.805
+ $X2=0 $Y2=0
cc_1015 N_A_278_793#_c_1037_n N_S[8]_c_1188_n 0.00543241f $X=1.96 $Y=4.1 $X2=0
+ $Y2=0
cc_1016 N_A_278_793#_c_1035_n S[8] 0.0163154f $X=2.43 $Y=4.685 $X2=0 $Y2=0
cc_1017 N_A_278_793#_c_1036_n S[8] 0.0127184f $X=2.715 $Y=3.805 $X2=0 $Y2=0
cc_1018 N_A_278_793#_c_1037_n S[8] 3.07062e-19 $X=1.96 $Y=4.1 $X2=0 $Y2=0
cc_1019 N_A_278_793#_M1099_g N_A_27_591#_c_4175_n 0.00176121f $X=1.49 $Y=3.365
+ $X2=0 $Y2=0
cc_1020 N_A_278_793#_M1099_g N_A_27_591#_c_4186_n 0.00400484f $X=1.49 $Y=3.365
+ $X2=0 $Y2=0
cc_1021 N_A_278_793#_M1111_g N_A_27_591#_c_4172_n 0.0124482f $X=1.96 $Y=3.365
+ $X2=0 $Y2=0
cc_1022 N_A_278_793#_c_1036_n N_A_27_591#_c_4172_n 0.0132748f $X=2.715 $Y=3.805
+ $X2=0 $Y2=0
cc_1023 N_A_278_793#_c_1043_n N_A_27_591#_c_4172_n 0.0413753f $X=2.715 $Y=3.13
+ $X2=0 $Y2=0
cc_1024 N_A_278_793#_c_1037_n N_A_27_591#_c_4172_n 0.00133381f $X=1.96 $Y=4.1
+ $X2=0 $Y2=0
cc_1025 N_A_278_793#_M1099_g N_A_27_591#_c_4191_n 0.00670811f $X=1.49 $Y=3.365
+ $X2=0 $Y2=0
cc_1026 N_A_278_793#_M1111_g N_A_27_591#_c_4191_n 0.00334069f $X=1.96 $Y=3.365
+ $X2=0 $Y2=0
cc_1027 N_A_278_793#_M1099_g N_A_27_591#_c_4193_n 7.75952e-19 $X=1.49 $Y=3.365
+ $X2=0 $Y2=0
cc_1028 N_A_278_793#_M1099_g N_A_27_591#_c_4183_n 0.00527796f $X=1.49 $Y=3.365
+ $X2=0 $Y2=0
cc_1029 N_A_278_793#_c_1043_n N_A_27_591#_c_4173_n 0.00738293f $X=2.715 $Y=3.13
+ $X2=0 $Y2=0
cc_1030 N_A_278_793#_M1099_g N_VPWR_c_4247_n 0.0012647f $X=1.49 $Y=3.365 $X2=0
+ $Y2=0
cc_1031 N_A_278_793#_c_1036_n N_VPWR_c_4249_n 0.00732952f $X=2.715 $Y=3.805
+ $X2=0 $Y2=0
cc_1032 N_A_278_793#_c_1043_n N_VPWR_c_4249_n 0.0321301f $X=2.715 $Y=3.13 $X2=0
+ $Y2=0
cc_1033 N_A_278_793#_M1111_g N_VPWR_c_4270_n 7.91347e-19 $X=1.96 $Y=3.365 $X2=0
+ $Y2=0
cc_1034 N_A_278_793#_c_1043_n N_VPWR_c_4270_n 0.0210596f $X=2.715 $Y=3.13 $X2=0
+ $Y2=0
cc_1035 N_A_278_793#_M1027_s VPWR 0.00179197f $X=2.59 $Y=2.955 $X2=0 $Y2=0
cc_1036 N_A_278_793#_M1099_g VPWR 0.00434142f $X=1.49 $Y=3.365 $X2=0 $Y2=0
cc_1037 N_A_278_793#_M1111_g VPWR 0.00546988f $X=1.96 $Y=3.365 $X2=0 $Y2=0
cc_1038 N_A_278_793#_c_1043_n VPWR 0.00594162f $X=2.715 $Y=3.13 $X2=0 $Y2=0
cc_1039 N_A_278_793#_M1099_g N_Z_c_5202_n 0.00268051f $X=1.49 $Y=3.365 $X2=0
+ $Y2=0
cc_1040 N_A_278_793#_c_1039_n N_Z_c_5202_n 0.0140957f $X=1.87 $Y=4.04 $X2=0
+ $Y2=0
cc_1041 N_A_278_793#_M1111_g N_Z_c_5202_n 0.00476154f $X=1.96 $Y=3.365 $X2=0
+ $Y2=0
cc_1042 N_A_278_793#_c_1035_n N_Z_c_5202_n 0.00967956f $X=2.43 $Y=4.685 $X2=0
+ $Y2=0
cc_1043 N_A_278_793#_c_1036_n N_Z_c_5202_n 0.0117695f $X=2.715 $Y=3.805 $X2=0
+ $Y2=0
cc_1044 N_A_278_793#_c_1037_n N_Z_c_5202_n 7.26438e-19 $X=1.96 $Y=4.1 $X2=0
+ $Y2=0
cc_1045 N_A_278_793#_c_1039_n N_Z_c_5211_n 0.00168443f $X=1.87 $Y=4.04 $X2=0
+ $Y2=0
cc_1046 N_A_278_793#_c_1040_n N_Z_c_5211_n 0.00180308f $X=1.58 $Y=4.04 $X2=0
+ $Y2=0
cc_1047 N_A_278_793#_c_1035_n N_Z_c_5211_n 0.0033343f $X=2.43 $Y=4.685 $X2=0
+ $Y2=0
cc_1048 N_A_278_793#_M1111_g N_Z_c_5243_n 0.00708682f $X=1.96 $Y=3.365 $X2=0
+ $Y2=0
cc_1049 N_A_278_793#_c_1036_n N_Z_c_5243_n 0.0132841f $X=2.715 $Y=3.805 $X2=0
+ $Y2=0
cc_1050 N_A_278_793#_c_1043_n N_Z_c_5243_n 0.0308332f $X=2.715 $Y=3.13 $X2=0
+ $Y2=0
cc_1051 N_A_278_793#_c_1037_n N_Z_c_5243_n 9.57301e-19 $X=1.96 $Y=4.1 $X2=0
+ $Y2=0
cc_1052 N_A_278_793#_M1099_g N_Z_c_5313_n 0.00635853f $X=1.49 $Y=3.365 $X2=0
+ $Y2=0
cc_1053 N_A_278_793#_M1099_g N_Z_c_5288_n 2.61869e-19 $X=1.49 $Y=3.365 $X2=0
+ $Y2=0
cc_1054 N_A_278_793#_M1099_g N_Z_c_5297_n 0.00978858f $X=1.49 $Y=3.365 $X2=0
+ $Y2=0
cc_1055 N_A_278_793#_c_1039_n N_Z_c_5297_n 8.37785e-19 $X=1.87 $Y=4.04 $X2=0
+ $Y2=0
cc_1056 N_A_278_793#_M1111_g N_Z_c_5297_n 0.00619657f $X=1.96 $Y=3.365 $X2=0
+ $Y2=0
cc_1057 N_A_278_793#_M1099_g N_Z_c_5257_n 0.00455034f $X=1.49 $Y=3.365 $X2=0
+ $Y2=0
cc_1058 N_A_278_793#_M1111_g N_Z_c_5257_n 0.00462236f $X=1.96 $Y=3.365 $X2=0
+ $Y2=0
cc_1059 N_A_278_793#_c_1035_n N_A_27_911#_c_7735_n 0.00358194f $X=2.43 $Y=4.685
+ $X2=0 $Y2=0
cc_1060 N_A_278_793#_c_1035_n N_A_27_911#_c_7748_n 0.0195704f $X=2.43 $Y=4.685
+ $X2=0 $Y2=0
cc_1061 N_A_278_793#_c_1036_n N_A_27_911#_c_7748_n 0.00285813f $X=2.715 $Y=3.805
+ $X2=0 $Y2=0
cc_1062 N_A_278_793#_c_1037_n N_A_27_911#_c_7748_n 0.00308807f $X=1.96 $Y=4.1
+ $X2=0 $Y2=0
cc_1063 N_A_278_793#_c_1035_n N_VGND_c_7809_n 0.0173402f $X=2.43 $Y=4.685 $X2=0
+ $Y2=0
cc_1064 N_A_278_793#_M1115_s VGND 0.00250855f $X=2.675 $Y=4.685 $X2=0 $Y2=0
cc_1065 N_A_278_793#_c_1035_n VGND 0.0186503f $X=2.43 $Y=4.685 $X2=0 $Y2=0
cc_1066 N_S[0]_c_1122_n N_S[8]_c_1191_n 0.0130744f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_1067 N_S[0]_c_1123_n N_S[1]_c_1246_n 0.0133556f $X=3.01 $Y=0.845 $X2=-0.19
+ $Y2=-0.24
cc_1068 N_S[0]_c_1122_n N_S[1]_c_1247_n 0.0418422f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_1069 S[0] N_S[1]_c_1247_n 8.74983e-19 $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_1070 N_S[0]_c_1122_n S[1] 8.74983e-19 $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_1071 S[0] S[1] 0.0208489f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_1072 N_S[0]_c_1122_n N_VPWR_c_4248_n 0.00456891f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_1073 S[0] N_VPWR_c_4248_n 0.00569857f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_1074 N_S[0]_c_1122_n N_VPWR_c_4270_n 0.0035837f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_1075 N_S[0]_c_1122_n VPWR 0.00710985f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_1076 N_S[0]_c_1114_n N_Z_c_5210_n 0.00413022f $X=1.46 $Y=0.255 $X2=0 $Y2=0
cc_1077 N_S[0]_c_1117_n N_Z_c_5210_n 0.00495983f $X=1.88 $Y=0.255 $X2=0 $Y2=0
cc_1078 N_S[0]_c_1119_n N_Z_c_5210_n 4.25992e-19 $X=2.365 $Y=0.845 $X2=0 $Y2=0
cc_1079 N_S[0]_c_1122_n N_Z_c_5242_n 0.00513674f $X=2.95 $Y=1.41 $X2=0 $Y2=0
cc_1080 S[0] N_Z_c_5242_n 0.00545567f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_1081 N_S[0]_c_1114_n N_Z_c_5226_n 0.00199103f $X=1.46 $Y=0.255 $X2=0 $Y2=0
cc_1082 N_S[0]_c_1117_n N_Z_c_5226_n 0.00133607f $X=1.88 $Y=0.255 $X2=0 $Y2=0
cc_1083 N_S[0]_c_1114_n N_A_27_47#_c_7692_n 0.00139422f $X=1.46 $Y=0.255 $X2=0
+ $Y2=0
cc_1084 N_S[0]_c_1114_n N_A_27_47#_c_7694_n 0.0132844f $X=1.46 $Y=0.255 $X2=0
+ $Y2=0
cc_1085 N_S[0]_c_1115_n N_A_27_47#_c_7694_n 0.00211351f $X=1.805 $Y=0.18 $X2=0
+ $Y2=0
cc_1086 N_S[0]_c_1117_n N_A_27_47#_c_7694_n 0.0126455f $X=1.88 $Y=0.255 $X2=0
+ $Y2=0
cc_1087 N_S[0]_c_1118_n N_A_27_47#_c_7694_n 0.00436105f $X=2.29 $Y=0.18 $X2=0
+ $Y2=0
cc_1088 N_S[0]_c_1119_n N_A_27_47#_c_7694_n 0.00349455f $X=2.365 $Y=0.845 $X2=0
+ $Y2=0
cc_1089 N_S[0]_c_1119_n N_A_27_47#_c_7705_n 0.00295202f $X=2.365 $Y=0.845 $X2=0
+ $Y2=0
cc_1090 N_S[0]_c_1123_n N_VGND_c_7779_n 0.00330937f $X=3.01 $Y=0.845 $X2=0 $Y2=0
cc_1091 N_S[0]_c_1116_n N_VGND_c_7807_n 0.0271255f $X=1.535 $Y=0.18 $X2=0 $Y2=0
cc_1092 N_S[0]_c_1123_n N_VGND_c_7807_n 0.00585385f $X=3.01 $Y=0.845 $X2=0 $Y2=0
cc_1093 N_S[0]_c_1115_n VGND 0.00642387f $X=1.805 $Y=0.18 $X2=0 $Y2=0
cc_1094 N_S[0]_c_1116_n VGND 0.00474746f $X=1.535 $Y=0.18 $X2=0 $Y2=0
cc_1095 N_S[0]_c_1118_n VGND 0.0193094f $X=2.29 $Y=0.18 $X2=0 $Y2=0
cc_1096 N_S[0]_c_1123_n VGND 0.0111218f $X=3.01 $Y=0.845 $X2=0 $Y2=0
cc_1097 N_S[0]_c_1124_n VGND 0.00366655f $X=1.88 $Y=0.18 $X2=0 $Y2=0
cc_1098 N_S[8]_c_1188_n N_S[9]_c_1309_n 0.0474978f $X=3.01 $Y=4.595 $X2=-0.19
+ $Y2=-0.24
cc_1099 S[8] N_S[9]_c_1309_n 8.74983e-19 $X=2.905 $Y=4.165 $X2=-0.19 $Y2=-0.24
cc_1100 N_S[8]_c_1191_n N_S[9]_c_1320_n 0.00770012f $X=2.95 $Y=4.03 $X2=0 $Y2=0
cc_1101 N_S[8]_c_1188_n S[9] 8.74983e-19 $X=3.01 $Y=4.595 $X2=0 $Y2=0
cc_1102 S[8] S[9] 0.0208489f $X=2.905 $Y=4.165 $X2=0 $Y2=0
cc_1103 N_S[8]_c_1191_n N_VPWR_c_4249_n 0.00362951f $X=2.95 $Y=4.03 $X2=0 $Y2=0
cc_1104 N_S[8]_c_1188_n N_VPWR_c_4249_n 9.39395e-19 $X=3.01 $Y=4.595 $X2=0 $Y2=0
cc_1105 S[8] N_VPWR_c_4249_n 0.00569857f $X=2.905 $Y=4.165 $X2=0 $Y2=0
cc_1106 N_S[8]_c_1191_n N_VPWR_c_4270_n 0.0035837f $X=2.95 $Y=4.03 $X2=0 $Y2=0
cc_1107 N_S[8]_c_1191_n VPWR 0.00710985f $X=2.95 $Y=4.03 $X2=0 $Y2=0
cc_1108 N_S[8]_c_1180_n N_Z_c_5202_n 0.00199103f $X=1.46 $Y=5.185 $X2=0 $Y2=0
cc_1109 N_S[8]_c_1183_n N_Z_c_5202_n 0.00133607f $X=1.88 $Y=5.185 $X2=0 $Y2=0
cc_1110 N_S[8]_c_1180_n N_Z_c_5211_n 0.00413022f $X=1.46 $Y=5.185 $X2=0 $Y2=0
cc_1111 N_S[8]_c_1183_n N_Z_c_5211_n 0.00495983f $X=1.88 $Y=5.185 $X2=0 $Y2=0
cc_1112 N_S[8]_c_1187_n N_Z_c_5211_n 4.25992e-19 $X=2.44 $Y=4.52 $X2=0 $Y2=0
cc_1113 N_S[8]_c_1191_n N_Z_c_5243_n 0.00477894f $X=2.95 $Y=4.03 $X2=0 $Y2=0
cc_1114 N_S[8]_c_1188_n N_Z_c_5243_n 3.57797e-19 $X=3.01 $Y=4.595 $X2=0 $Y2=0
cc_1115 S[8] N_Z_c_5243_n 0.00545567f $X=2.905 $Y=4.165 $X2=0 $Y2=0
cc_1116 N_S[8]_c_1180_n N_A_27_911#_c_7734_n 0.00139422f $X=1.46 $Y=5.185 $X2=0
+ $Y2=0
cc_1117 N_S[8]_c_1180_n N_A_27_911#_c_7735_n 0.0132844f $X=1.46 $Y=5.185 $X2=0
+ $Y2=0
cc_1118 N_S[8]_c_1181_n N_A_27_911#_c_7735_n 0.00211351f $X=1.805 $Y=5.26 $X2=0
+ $Y2=0
cc_1119 N_S[8]_c_1183_n N_A_27_911#_c_7735_n 0.0126455f $X=1.88 $Y=5.185 $X2=0
+ $Y2=0
cc_1120 N_S[8]_c_1184_n N_A_27_911#_c_7735_n 0.00436105f $X=2.29 $Y=5.26 $X2=0
+ $Y2=0
cc_1121 N_S[8]_c_1185_n N_A_27_911#_c_7735_n 0.00349455f $X=2.365 $Y=5.185 $X2=0
+ $Y2=0
cc_1122 N_S[8]_c_1185_n N_A_27_911#_c_7748_n 0.00295202f $X=2.365 $Y=5.185 $X2=0
+ $Y2=0
cc_1123 N_S[8]_c_1188_n N_VGND_c_7780_n 0.00330937f $X=3.01 $Y=4.595 $X2=0 $Y2=0
cc_1124 N_S[8]_c_1182_n N_VGND_c_7809_n 0.0271255f $X=1.535 $Y=5.26 $X2=0 $Y2=0
cc_1125 N_S[8]_c_1188_n N_VGND_c_7809_n 0.00585385f $X=3.01 $Y=4.595 $X2=0 $Y2=0
cc_1126 N_S[8]_c_1181_n VGND 0.00642387f $X=1.805 $Y=5.26 $X2=0 $Y2=0
cc_1127 N_S[8]_c_1182_n VGND 0.00474746f $X=1.535 $Y=5.26 $X2=0 $Y2=0
cc_1128 N_S[8]_c_1184_n VGND 0.0193094f $X=2.29 $Y=5.26 $X2=0 $Y2=0
cc_1129 N_S[8]_c_1188_n VGND 0.0111218f $X=3.01 $Y=4.595 $X2=0 $Y2=0
cc_1130 N_S[8]_c_1189_n VGND 0.00366655f $X=1.88 $Y=5.26 $X2=0 $Y2=0
cc_1131 N_S[1]_c_1247_n N_S[9]_c_1320_n 0.0130744f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_1132 N_S[1]_c_1254_n N_A_701_47#_c_1380_n 0.00779314f $X=4.98 $Y=0.255 $X2=0
+ $Y2=0
cc_1133 N_S[1]_c_1247_n N_A_701_47#_c_1375_n 0.00692516f $X=3.49 $Y=1.41 $X2=0
+ $Y2=0
cc_1134 N_S[1]_c_1248_n N_A_701_47#_c_1375_n 0.00920672f $X=4 $Y=0.92 $X2=0
+ $Y2=0
cc_1135 N_S[1]_c_1252_n N_A_701_47#_c_1375_n 0.00810157f $X=4.56 $Y=0.255 $X2=0
+ $Y2=0
cc_1136 S[1] N_A_701_47#_c_1375_n 3.07062e-19 $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_1137 N_S[1]_c_1247_n N_A_701_47#_c_1383_n 0.00861299f $X=3.49 $Y=1.41 $X2=0
+ $Y2=0
cc_1138 N_S[1]_c_1246_n N_A_701_47#_c_1376_n 0.00149517f $X=3.43 $Y=0.845 $X2=0
+ $Y2=0
cc_1139 N_S[1]_c_1247_n N_A_701_47#_c_1376_n 0.00205356f $X=3.49 $Y=1.41 $X2=0
+ $Y2=0
cc_1140 N_S[1]_c_1248_n N_A_701_47#_c_1376_n 0.0135307f $X=4 $Y=0.92 $X2=0 $Y2=0
cc_1141 N_S[1]_c_1249_n N_A_701_47#_c_1376_n 0.00267287f $X=4.075 $Y=0.845 $X2=0
+ $Y2=0
cc_1142 N_S[1]_c_1252_n N_A_701_47#_c_1376_n 7.04048e-19 $X=4.56 $Y=0.255 $X2=0
+ $Y2=0
cc_1143 S[1] N_A_701_47#_c_1376_n 0.0101733f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_1144 N_S[1]_c_1247_n N_A_701_47#_c_1377_n 0.0105766f $X=3.49 $Y=1.41 $X2=0
+ $Y2=0
cc_1145 N_S[1]_c_1249_n N_A_701_47#_c_1377_n 0.0100587f $X=4.075 $Y=0.845 $X2=0
+ $Y2=0
cc_1146 S[1] N_A_701_47#_c_1377_n 0.0061421f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_1147 N_S[1]_c_1247_n N_A_701_47#_c_1378_n 0.00828481f $X=3.49 $Y=1.41 $X2=0
+ $Y2=0
cc_1148 N_S[1]_c_1248_n N_A_701_47#_c_1378_n 0.00785343f $X=4 $Y=0.92 $X2=0
+ $Y2=0
cc_1149 S[1] N_A_701_47#_c_1378_n 0.0127184f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_1150 N_S[1]_c_1253_n N_D[1]_M1074_g 0.0165585f $X=4.905 $Y=0.18 $X2=0 $Y2=0
cc_1151 N_S[1]_c_1247_n N_VPWR_c_4248_n 0.00456891f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_1152 S[1] N_VPWR_c_4248_n 0.00569857f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_1153 N_S[1]_c_1247_n VPWR 0.00710985f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_1154 N_S[1]_c_1247_n N_VPWR_c_4281_n 0.0035837f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_1155 N_S[1]_c_1249_n N_Z_c_5212_n 4.25992e-19 $X=4.075 $Y=0.845 $X2=0 $Y2=0
cc_1156 N_S[1]_c_1252_n N_Z_c_5212_n 0.00495983f $X=4.56 $Y=0.255 $X2=0 $Y2=0
cc_1157 N_S[1]_c_1254_n N_Z_c_5212_n 0.00413022f $X=4.98 $Y=0.255 $X2=0 $Y2=0
cc_1158 N_S[1]_c_1247_n N_Z_c_5242_n 0.00513674f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_1159 S[1] N_Z_c_5242_n 0.00545567f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_1160 N_S[1]_c_1252_n N_Z_c_5227_n 0.00133607f $X=4.56 $Y=0.255 $X2=0 $Y2=0
cc_1161 N_S[1]_c_1254_n N_Z_c_5227_n 0.00199103f $X=4.98 $Y=0.255 $X2=0 $Y2=0
cc_1162 N_S[1]_c_1246_n N_VGND_c_7779_n 0.00330937f $X=3.43 $Y=0.845 $X2=0 $Y2=0
cc_1163 N_S[1]_c_1246_n VGND 0.0111218f $X=3.43 $Y=0.845 $X2=0 $Y2=0
cc_1164 N_S[1]_c_1250_n VGND 0.0119932f $X=4.485 $Y=0.18 $X2=0 $Y2=0
cc_1165 N_S[1]_c_1251_n VGND 0.00731624f $X=4.15 $Y=0.18 $X2=0 $Y2=0
cc_1166 N_S[1]_c_1253_n VGND 0.0111713f $X=4.905 $Y=0.18 $X2=0 $Y2=0
cc_1167 N_S[1]_c_1255_n VGND 0.00366655f $X=4.56 $Y=0.18 $X2=0 $Y2=0
cc_1168 N_S[1]_c_1246_n N_VGND_c_7829_n 0.00585385f $X=3.43 $Y=0.845 $X2=0 $Y2=0
cc_1169 N_S[1]_c_1251_n N_VGND_c_7829_n 0.0271255f $X=4.15 $Y=0.18 $X2=0 $Y2=0
cc_1170 N_S[1]_c_1249_n N_A_845_69#_c_8343_n 0.00295202f $X=4.075 $Y=0.845 $X2=0
+ $Y2=0
cc_1171 N_S[1]_c_1252_n N_A_845_69#_c_8339_n 0.0126455f $X=4.56 $Y=0.255 $X2=0
+ $Y2=0
cc_1172 N_S[1]_c_1253_n N_A_845_69#_c_8339_n 0.00211351f $X=4.905 $Y=0.18 $X2=0
+ $Y2=0
cc_1173 N_S[1]_c_1254_n N_A_845_69#_c_8339_n 0.0132844f $X=4.98 $Y=0.255 $X2=0
+ $Y2=0
cc_1174 N_S[1]_c_1249_n N_A_845_69#_c_8340_n 0.00349455f $X=4.075 $Y=0.845 $X2=0
+ $Y2=0
cc_1175 N_S[1]_c_1250_n N_A_845_69#_c_8340_n 0.00436105f $X=4.485 $Y=0.18 $X2=0
+ $Y2=0
cc_1176 N_S[1]_c_1254_n N_A_845_69#_c_8342_n 0.00139422f $X=4.98 $Y=0.255 $X2=0
+ $Y2=0
cc_1177 N_S[9]_c_1316_n N_A_701_937#_c_1461_n 0.00779314f $X=4.98 $Y=5.185 $X2=0
+ $Y2=0
cc_1178 N_S[9]_c_1309_n N_A_701_937#_c_1456_n 0.00543241f $X=3.43 $Y=4.595 $X2=0
+ $Y2=0
cc_1179 N_S[9]_c_1320_n N_A_701_937#_c_1456_n 0.00149275f $X=3.49 $Y=4.03 $X2=0
+ $Y2=0
cc_1180 N_S[9]_c_1310_n N_A_701_937#_c_1456_n 0.00920672f $X=4 $Y=4.52 $X2=0
+ $Y2=0
cc_1181 N_S[9]_c_1314_n N_A_701_937#_c_1456_n 0.00810157f $X=4.56 $Y=5.185 $X2=0
+ $Y2=0
cc_1182 S[9] N_A_701_937#_c_1456_n 3.07062e-19 $X=3.365 $Y=4.165 $X2=0 $Y2=0
cc_1183 N_S[9]_c_1320_n N_A_701_937#_c_1464_n 0.00861299f $X=3.49 $Y=4.03 $X2=0
+ $Y2=0
cc_1184 N_S[9]_c_1309_n N_A_701_937#_c_1457_n 0.00354873f $X=3.43 $Y=4.595 $X2=0
+ $Y2=0
cc_1185 N_S[9]_c_1310_n N_A_701_937#_c_1457_n 0.0135307f $X=4 $Y=4.52 $X2=0
+ $Y2=0
cc_1186 N_S[9]_c_1311_n N_A_701_937#_c_1457_n 0.00267287f $X=4.075 $Y=5.185
+ $X2=0 $Y2=0
cc_1187 N_S[9]_c_1314_n N_A_701_937#_c_1457_n 7.04048e-19 $X=4.56 $Y=5.185 $X2=0
+ $Y2=0
cc_1188 S[9] N_A_701_937#_c_1457_n 0.0101733f $X=3.365 $Y=4.165 $X2=0 $Y2=0
cc_1189 N_S[9]_c_1309_n N_A_701_937#_c_1458_n 0.0105766f $X=3.43 $Y=4.595 $X2=0
+ $Y2=0
cc_1190 N_S[9]_c_1311_n N_A_701_937#_c_1458_n 0.0100374f $X=4.075 $Y=5.185 $X2=0
+ $Y2=0
cc_1191 S[9] N_A_701_937#_c_1458_n 0.0061421f $X=3.365 $Y=4.165 $X2=0 $Y2=0
cc_1192 N_S[9]_c_1309_n N_A_701_937#_c_1459_n 0.00441664f $X=3.43 $Y=4.595 $X2=0
+ $Y2=0
cc_1193 N_S[9]_c_1320_n N_A_701_937#_c_1459_n 0.00386817f $X=3.49 $Y=4.03 $X2=0
+ $Y2=0
cc_1194 N_S[9]_c_1310_n N_A_701_937#_c_1459_n 0.00785343f $X=4 $Y=4.52 $X2=0
+ $Y2=0
cc_1195 S[9] N_A_701_937#_c_1459_n 0.0127184f $X=3.365 $Y=4.165 $X2=0 $Y2=0
cc_1196 N_S[9]_c_1316_n N_D[9]_M1026_g 0.0165585f $X=4.98 $Y=5.185 $X2=0 $Y2=0
cc_1197 N_S[9]_c_1309_n N_VPWR_c_4249_n 9.39395e-19 $X=3.43 $Y=4.595 $X2=0 $Y2=0
cc_1198 N_S[9]_c_1320_n N_VPWR_c_4249_n 0.00362951f $X=3.49 $Y=4.03 $X2=0 $Y2=0
cc_1199 S[9] N_VPWR_c_4249_n 0.00569857f $X=3.365 $Y=4.165 $X2=0 $Y2=0
cc_1200 N_S[9]_c_1320_n VPWR 0.00710985f $X=3.49 $Y=4.03 $X2=0 $Y2=0
cc_1201 N_S[9]_c_1320_n N_VPWR_c_4281_n 0.0035837f $X=3.49 $Y=4.03 $X2=0 $Y2=0
cc_1202 N_S[9]_c_1314_n N_Z_c_5203_n 0.00133607f $X=4.56 $Y=5.185 $X2=0 $Y2=0
cc_1203 N_S[9]_c_1316_n N_Z_c_5203_n 0.00199103f $X=4.98 $Y=5.185 $X2=0 $Y2=0
cc_1204 N_S[9]_c_1310_n N_Z_c_5213_n 4.25992e-19 $X=4 $Y=4.52 $X2=0 $Y2=0
cc_1205 N_S[9]_c_1314_n N_Z_c_5213_n 0.00495983f $X=4.56 $Y=5.185 $X2=0 $Y2=0
cc_1206 N_S[9]_c_1316_n N_Z_c_5213_n 0.00413022f $X=4.98 $Y=5.185 $X2=0 $Y2=0
cc_1207 N_S[9]_c_1309_n N_Z_c_5243_n 3.57797e-19 $X=3.43 $Y=4.595 $X2=0 $Y2=0
cc_1208 N_S[9]_c_1320_n N_Z_c_5243_n 0.00477894f $X=3.49 $Y=4.03 $X2=0 $Y2=0
cc_1209 S[9] N_Z_c_5243_n 0.00545567f $X=3.365 $Y=4.165 $X2=0 $Y2=0
cc_1210 N_S[9]_c_1309_n N_VGND_c_7780_n 0.00330937f $X=3.43 $Y=4.595 $X2=0 $Y2=0
cc_1211 N_S[9]_c_1309_n VGND 0.0111218f $X=3.43 $Y=4.595 $X2=0 $Y2=0
cc_1212 N_S[9]_c_1312_n VGND 0.0119932f $X=4.485 $Y=5.26 $X2=0 $Y2=0
cc_1213 N_S[9]_c_1313_n VGND 0.00731624f $X=4.15 $Y=5.26 $X2=0 $Y2=0
cc_1214 N_S[9]_c_1315_n VGND 0.0111713f $X=4.905 $Y=5.26 $X2=0 $Y2=0
cc_1215 N_S[9]_c_1317_n VGND 0.00366655f $X=4.56 $Y=5.26 $X2=0 $Y2=0
cc_1216 N_S[9]_c_1309_n N_VGND_c_7830_n 0.00585385f $X=3.43 $Y=4.595 $X2=0 $Y2=0
cc_1217 N_S[9]_c_1313_n N_VGND_c_7830_n 0.0271255f $X=4.15 $Y=5.26 $X2=0 $Y2=0
cc_1218 N_S[9]_c_1311_n N_A_845_915#_c_8391_n 0.00295202f $X=4.075 $Y=5.185
+ $X2=0 $Y2=0
cc_1219 N_S[9]_c_1314_n N_A_845_915#_c_8387_n 0.0126455f $X=4.56 $Y=5.185 $X2=0
+ $Y2=0
cc_1220 N_S[9]_c_1315_n N_A_845_915#_c_8387_n 0.00211351f $X=4.905 $Y=5.26 $X2=0
+ $Y2=0
cc_1221 N_S[9]_c_1316_n N_A_845_915#_c_8387_n 0.0132844f $X=4.98 $Y=5.185 $X2=0
+ $Y2=0
cc_1222 N_S[9]_c_1311_n N_A_845_915#_c_8388_n 0.00349455f $X=4.075 $Y=5.185
+ $X2=0 $Y2=0
cc_1223 N_S[9]_c_1312_n N_A_845_915#_c_8388_n 0.00436105f $X=4.485 $Y=5.26 $X2=0
+ $Y2=0
cc_1224 N_S[9]_c_1316_n N_A_845_915#_c_8389_n 0.00139422f $X=4.98 $Y=5.185 $X2=0
+ $Y2=0
cc_1225 N_A_701_47#_M1084_g N_A_701_937#_M1036_g 0.0130744f $X=4.48 $Y=2.075
+ $X2=0 $Y2=0
cc_1226 N_A_701_47#_M1113_g N_A_701_937#_M1157_g 0.0130744f $X=4.95 $Y=2.075
+ $X2=0 $Y2=0
cc_1227 N_A_701_47#_c_1380_n N_D[1]_M1052_g 0.00671996f $X=4.86 $Y=1.4 $X2=0
+ $Y2=0
cc_1228 N_A_701_47#_M1113_g N_D[1]_M1052_g 0.025073f $X=4.95 $Y=2.075 $X2=0
+ $Y2=0
cc_1229 N_A_701_47#_c_1383_n N_VPWR_c_4248_n 0.0321301f $X=3.725 $Y=2.31 $X2=0
+ $Y2=0
cc_1230 N_A_701_47#_c_1378_n N_VPWR_c_4248_n 0.00732952f $X=4.01 $Y=1.42 $X2=0
+ $Y2=0
cc_1231 N_A_701_47#_M1113_g N_VPWR_c_4250_n 0.00107878f $X=4.95 $Y=2.075 $X2=0
+ $Y2=0
cc_1232 N_A_701_47#_M1089_d VPWR 0.00179197f $X=3.58 $Y=1.485 $X2=0 $Y2=0
cc_1233 N_A_701_47#_M1084_g VPWR 0.0054792f $X=4.48 $Y=2.075 $X2=0 $Y2=0
cc_1234 N_A_701_47#_M1113_g VPWR 0.00435072f $X=4.95 $Y=2.075 $X2=0 $Y2=0
cc_1235 N_A_701_47#_c_1383_n VPWR 0.00594162f $X=3.725 $Y=2.31 $X2=0 $Y2=0
cc_1236 N_A_701_47#_M1084_g N_VPWR_c_4281_n 8.06528e-19 $X=4.48 $Y=2.075 $X2=0
+ $Y2=0
cc_1237 N_A_701_47#_c_1383_n N_VPWR_c_4281_n 0.0210596f $X=3.725 $Y=2.31 $X2=0
+ $Y2=0
cc_1238 N_A_701_47#_c_1380_n N_Z_c_5212_n 0.00348752f $X=4.86 $Y=1.4 $X2=0 $Y2=0
cc_1239 N_A_701_47#_c_1376_n N_Z_c_5212_n 0.0033343f $X=4.01 $Y=1.205 $X2=0
+ $Y2=0
cc_1240 N_A_701_47#_M1084_g N_Z_c_5242_n 0.00708998f $X=4.48 $Y=2.075 $X2=0
+ $Y2=0
cc_1241 N_A_701_47#_c_1375_n N_Z_c_5242_n 9.57301e-19 $X=4.57 $Y=1.4 $X2=0 $Y2=0
cc_1242 N_A_701_47#_c_1383_n N_Z_c_5242_n 0.0308332f $X=3.725 $Y=2.31 $X2=0
+ $Y2=0
cc_1243 N_A_701_47#_c_1378_n N_Z_c_5242_n 0.0132841f $X=4.01 $Y=1.42 $X2=0 $Y2=0
cc_1244 N_A_701_47#_M1113_g N_Z_c_5244_n 0.00404618f $X=4.95 $Y=2.075 $X2=0
+ $Y2=0
cc_1245 N_A_701_47#_M1113_g N_Z_c_5357_n 0.00513826f $X=4.95 $Y=2.075 $X2=0
+ $Y2=0
cc_1246 N_A_701_47#_M1084_g N_Z_c_5358_n 0.00619657f $X=4.48 $Y=2.075 $X2=0
+ $Y2=0
cc_1247 N_A_701_47#_c_1380_n N_Z_c_5358_n 8.37785e-19 $X=4.86 $Y=1.4 $X2=0 $Y2=0
cc_1248 N_A_701_47#_M1113_g N_Z_c_5358_n 0.00978858f $X=4.95 $Y=2.075 $X2=0
+ $Y2=0
cc_1249 N_A_701_47#_M1084_g N_Z_c_5227_n 0.00476154f $X=4.48 $Y=2.075 $X2=0
+ $Y2=0
cc_1250 N_A_701_47#_c_1380_n N_Z_c_5227_n 0.0140957f $X=4.86 $Y=1.4 $X2=0 $Y2=0
cc_1251 N_A_701_47#_c_1375_n N_Z_c_5227_n 7.26438e-19 $X=4.57 $Y=1.4 $X2=0 $Y2=0
cc_1252 N_A_701_47#_M1113_g N_Z_c_5227_n 0.00268051f $X=4.95 $Y=2.075 $X2=0
+ $Y2=0
cc_1253 N_A_701_47#_c_1376_n N_Z_c_5227_n 0.00967956f $X=4.01 $Y=1.205 $X2=0
+ $Y2=0
cc_1254 N_A_701_47#_c_1378_n N_Z_c_5227_n 0.0117695f $X=4.01 $Y=1.42 $X2=0 $Y2=0
cc_1255 N_A_701_47#_M1113_g N_Z_c_5367_n 2.61869e-19 $X=4.95 $Y=2.075 $X2=0
+ $Y2=0
cc_1256 N_A_701_47#_M1084_g N_Z_c_5259_n 0.00462462f $X=4.48 $Y=2.075 $X2=0
+ $Y2=0
cc_1257 N_A_701_47#_M1113_g N_Z_c_5259_n 0.00455034f $X=4.95 $Y=2.075 $X2=0
+ $Y2=0
cc_1258 N_A_701_47#_M1113_g N_A_824_333#_c_6423_n 0.00176121f $X=4.95 $Y=2.075
+ $X2=0 $Y2=0
cc_1259 N_A_701_47#_M1084_g N_A_824_333#_c_6424_n 0.00334959f $X=4.48 $Y=2.075
+ $X2=0 $Y2=0
cc_1260 N_A_701_47#_M1113_g N_A_824_333#_c_6424_n 0.00463461f $X=4.95 $Y=2.075
+ $X2=0 $Y2=0
cc_1261 N_A_701_47#_c_1383_n N_A_824_333#_c_6419_n 0.00738363f $X=3.725 $Y=2.31
+ $X2=0 $Y2=0
cc_1262 N_A_701_47#_M1113_g N_A_824_333#_c_6427_n 7.75952e-19 $X=4.95 $Y=2.075
+ $X2=0 $Y2=0
cc_1263 N_A_701_47#_M1084_g N_A_824_333#_c_6428_n 0.00692695f $X=4.48 $Y=2.075
+ $X2=0 $Y2=0
cc_1264 N_A_701_47#_M1113_g N_A_824_333#_c_6429_n 0.00415998f $X=4.95 $Y=2.075
+ $X2=0 $Y2=0
cc_1265 N_A_701_47#_M1084_g N_A_824_333#_c_6421_n 0.00550198f $X=4.48 $Y=2.075
+ $X2=0 $Y2=0
cc_1266 N_A_701_47#_c_1375_n N_A_824_333#_c_6421_n 0.00133381f $X=4.57 $Y=1.4
+ $X2=0 $Y2=0
cc_1267 N_A_701_47#_c_1383_n N_A_824_333#_c_6421_n 0.0413447f $X=3.725 $Y=2.31
+ $X2=0 $Y2=0
cc_1268 N_A_701_47#_c_1378_n N_A_824_333#_c_6421_n 0.0132748f $X=4.01 $Y=1.42
+ $X2=0 $Y2=0
cc_1269 N_A_701_47#_M1113_g N_A_824_333#_c_6434_n 0.00508488f $X=4.95 $Y=2.075
+ $X2=0 $Y2=0
cc_1270 N_A_701_47#_M1072_d VGND 0.00250855f $X=3.505 $Y=0.235 $X2=0 $Y2=0
cc_1271 N_A_701_47#_c_1377_n VGND 0.0186564f $X=3.64 $Y=0.495 $X2=0 $Y2=0
cc_1272 N_A_701_47#_c_1377_n N_VGND_c_7829_n 0.0173492f $X=3.64 $Y=0.495 $X2=0
+ $Y2=0
cc_1273 N_A_701_47#_c_1375_n N_A_845_69#_c_8343_n 0.00308807f $X=4.57 $Y=1.4
+ $X2=0 $Y2=0
cc_1274 N_A_701_47#_c_1376_n N_A_845_69#_c_8343_n 0.00101918f $X=4.01 $Y=1.205
+ $X2=0 $Y2=0
cc_1275 N_A_701_47#_c_1377_n N_A_845_69#_c_8343_n 0.0185512f $X=3.64 $Y=0.495
+ $X2=0 $Y2=0
cc_1276 N_A_701_47#_c_1378_n N_A_845_69#_c_8343_n 0.00285813f $X=4.01 $Y=1.42
+ $X2=0 $Y2=0
cc_1277 N_A_701_47#_c_1377_n N_A_845_69#_c_8340_n 0.00358194f $X=3.64 $Y=0.495
+ $X2=0 $Y2=0
cc_1278 N_A_701_937#_c_1461_n N_D[9]_M1056_g 0.00671996f $X=4.86 $Y=4.04 $X2=0
+ $Y2=0
cc_1279 N_A_701_937#_M1157_g N_D[9]_M1056_g 0.0250718f $X=4.95 $Y=3.365 $X2=0
+ $Y2=0
cc_1280 N_A_701_937#_c_1464_n N_VPWR_c_4249_n 0.0321301f $X=3.725 $Y=3.13 $X2=0
+ $Y2=0
cc_1281 N_A_701_937#_c_1459_n N_VPWR_c_4249_n 0.00732952f $X=4.01 $Y=4.02 $X2=0
+ $Y2=0
cc_1282 N_A_701_937#_M1157_g N_VPWR_c_4251_n 0.0013032f $X=4.95 $Y=3.365 $X2=0
+ $Y2=0
cc_1283 N_A_701_937#_M1092_d VPWR 0.00179197f $X=3.58 $Y=2.955 $X2=0 $Y2=0
cc_1284 N_A_701_937#_M1036_g VPWR 0.00546988f $X=4.48 $Y=3.365 $X2=0 $Y2=0
cc_1285 N_A_701_937#_M1157_g VPWR 0.00434142f $X=4.95 $Y=3.365 $X2=0 $Y2=0
cc_1286 N_A_701_937#_c_1464_n VPWR 0.00594162f $X=3.725 $Y=3.13 $X2=0 $Y2=0
cc_1287 N_A_701_937#_M1036_g N_VPWR_c_4281_n 7.91347e-19 $X=4.48 $Y=3.365 $X2=0
+ $Y2=0
cc_1288 N_A_701_937#_c_1464_n N_VPWR_c_4281_n 0.0210596f $X=3.725 $Y=3.13 $X2=0
+ $Y2=0
cc_1289 N_A_701_937#_M1036_g N_Z_c_5203_n 0.00476154f $X=4.48 $Y=3.365 $X2=0
+ $Y2=0
cc_1290 N_A_701_937#_c_1461_n N_Z_c_5203_n 0.0140957f $X=4.86 $Y=4.04 $X2=0
+ $Y2=0
cc_1291 N_A_701_937#_c_1456_n N_Z_c_5203_n 7.26438e-19 $X=4.57 $Y=4.04 $X2=0
+ $Y2=0
cc_1292 N_A_701_937#_M1157_g N_Z_c_5203_n 0.00268051f $X=4.95 $Y=3.365 $X2=0
+ $Y2=0
cc_1293 N_A_701_937#_c_1457_n N_Z_c_5203_n 0.00967956f $X=4.01 $Y=4.685 $X2=0
+ $Y2=0
cc_1294 N_A_701_937#_c_1459_n N_Z_c_5203_n 0.0117695f $X=4.01 $Y=4.02 $X2=0
+ $Y2=0
cc_1295 N_A_701_937#_c_1461_n N_Z_c_5213_n 0.00348752f $X=4.86 $Y=4.04 $X2=0
+ $Y2=0
cc_1296 N_A_701_937#_c_1457_n N_Z_c_5213_n 0.0033343f $X=4.01 $Y=4.685 $X2=0
+ $Y2=0
cc_1297 N_A_701_937#_M1036_g N_Z_c_5243_n 0.00708682f $X=4.48 $Y=3.365 $X2=0
+ $Y2=0
cc_1298 N_A_701_937#_c_1456_n N_Z_c_5243_n 9.57301e-19 $X=4.57 $Y=4.04 $X2=0
+ $Y2=0
cc_1299 N_A_701_937#_c_1464_n N_Z_c_5243_n 0.0308332f $X=3.725 $Y=3.13 $X2=0
+ $Y2=0
cc_1300 N_A_701_937#_c_1459_n N_Z_c_5243_n 0.0132841f $X=4.01 $Y=4.02 $X2=0
+ $Y2=0
cc_1301 N_A_701_937#_M1157_g N_Z_c_5245_n 0.0040431f $X=4.95 $Y=3.365 $X2=0
+ $Y2=0
cc_1302 N_A_701_937#_M1157_g N_Z_c_5383_n 0.00513826f $X=4.95 $Y=3.365 $X2=0
+ $Y2=0
cc_1303 N_A_701_937#_M1157_g N_Z_c_5358_n 2.61869e-19 $X=4.95 $Y=3.365 $X2=0
+ $Y2=0
cc_1304 N_A_701_937#_M1036_g N_Z_c_5367_n 0.00619657f $X=4.48 $Y=3.365 $X2=0
+ $Y2=0
cc_1305 N_A_701_937#_c_1461_n N_Z_c_5367_n 8.37785e-19 $X=4.86 $Y=4.04 $X2=0
+ $Y2=0
cc_1306 N_A_701_937#_M1157_g N_Z_c_5367_n 0.00978858f $X=4.95 $Y=3.365 $X2=0
+ $Y2=0
cc_1307 N_A_701_937#_M1036_g N_Z_c_5259_n 0.00462236f $X=4.48 $Y=3.365 $X2=0
+ $Y2=0
cc_1308 N_A_701_937#_M1157_g N_Z_c_5259_n 0.00455034f $X=4.95 $Y=3.365 $X2=0
+ $Y2=0
cc_1309 N_A_701_937#_M1157_g N_A_824_591#_c_6519_n 0.00176121f $X=4.95 $Y=3.365
+ $X2=0 $Y2=0
cc_1310 N_A_701_937#_M1036_g N_A_824_591#_c_6516_n 0.0124482f $X=4.48 $Y=3.365
+ $X2=0 $Y2=0
cc_1311 N_A_701_937#_c_1456_n N_A_824_591#_c_6516_n 0.00133381f $X=4.57 $Y=4.04
+ $X2=0 $Y2=0
cc_1312 N_A_701_937#_c_1464_n N_A_824_591#_c_6516_n 0.0413753f $X=3.725 $Y=3.13
+ $X2=0 $Y2=0
cc_1313 N_A_701_937#_c_1459_n N_A_824_591#_c_6516_n 0.0132748f $X=4.01 $Y=4.02
+ $X2=0 $Y2=0
cc_1314 N_A_701_937#_M1157_g N_A_824_591#_c_6524_n 0.00400484f $X=4.95 $Y=3.365
+ $X2=0 $Y2=0
cc_1315 N_A_701_937#_M1036_g N_A_824_591#_c_6525_n 0.00334069f $X=4.48 $Y=3.365
+ $X2=0 $Y2=0
cc_1316 N_A_701_937#_M1157_g N_A_824_591#_c_6525_n 0.00470988f $X=4.95 $Y=3.365
+ $X2=0 $Y2=0
cc_1317 N_A_701_937#_c_1464_n N_A_824_591#_c_6517_n 0.00738293f $X=3.725 $Y=3.13
+ $X2=0 $Y2=0
cc_1318 N_A_701_937#_M1157_g N_A_824_591#_c_6528_n 7.75952e-19 $X=4.95 $Y=3.365
+ $X2=0 $Y2=0
cc_1319 N_A_701_937#_M1157_g N_A_824_591#_c_6529_n 0.00508821f $X=4.95 $Y=3.365
+ $X2=0 $Y2=0
cc_1320 N_A_701_937#_M1039_d VGND 0.00250855f $X=3.505 $Y=4.685 $X2=0 $Y2=0
cc_1321 N_A_701_937#_c_1458_n VGND 0.0186503f $X=3.64 $Y=4.945 $X2=0 $Y2=0
cc_1322 N_A_701_937#_c_1458_n N_VGND_c_7830_n 0.0173402f $X=3.64 $Y=4.945 $X2=0
+ $Y2=0
cc_1323 N_A_701_937#_c_1456_n N_A_845_915#_c_8391_n 0.00308807f $X=4.57 $Y=4.04
+ $X2=0 $Y2=0
cc_1324 N_A_701_937#_c_1457_n N_A_845_915#_c_8391_n 0.00101918f $X=4.01 $Y=4.685
+ $X2=0 $Y2=0
cc_1325 N_A_701_937#_c_1458_n N_A_845_915#_c_8391_n 0.0185512f $X=3.64 $Y=4.945
+ $X2=0 $Y2=0
cc_1326 N_A_701_937#_c_1459_n N_A_845_915#_c_8391_n 0.00285813f $X=4.01 $Y=4.02
+ $X2=0 $Y2=0
cc_1327 N_A_701_937#_c_1458_n N_A_845_915#_c_8388_n 0.00358194f $X=3.64 $Y=4.945
+ $X2=0 $Y2=0
cc_1328 N_D[1]_M1052_g N_D[9]_M1056_g 0.0129371f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_1329 N_D[1]_M1097_g N_D[9]_M1101_g 0.0130744f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_1330 D[1] N_D[2]_c_1655_n 0.0231965f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_1331 N_D[1]_c_1542_n N_D[2]_c_1655_n 7.85936e-19 $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_1332 D[1] N_D[2]_c_1656_n 7.85936e-19 $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_1333 N_D[1]_c_1542_n N_D[2]_c_1656_n 0.00603597f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_1334 N_D[1]_M1052_g N_VPWR_c_4250_n 0.00848021f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_1335 N_D[1]_M1097_g N_VPWR_c_4250_n 0.00338721f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_1336 N_D[1]_M1052_g N_VPWR_c_4376_n 0.00295119f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_1337 N_D[1]_M1097_g N_VPWR_c_4376_n 0.00311479f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_1338 N_D[1]_M1052_g VPWR 0.00350923f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_1339 N_D[1]_M1097_g VPWR 0.00568683f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_1340 N_D[1]_M1052_g N_VPWR_c_4282_n 0.00342413f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_1341 N_D[1]_M1097_g N_VPWR_c_4283_n 0.0033767f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_1342 N_D[1]_M1052_g N_Z_c_5244_n 0.0033316f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_1343 N_D[1]_M1097_g N_Z_c_5244_n 0.00312829f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_1344 D[1] N_Z_c_5244_n 0.00125914f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_1345 N_D[1]_M1052_g N_Z_c_5227_n 0.00112534f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_1346 N_D[1]_M1074_g N_Z_c_5227_n 8.13311e-19 $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_1347 D[1] N_Z_c_5227_n 0.00742792f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_1348 N_D[1]_c_1542_n N_Z_c_5227_n 0.00583073f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_1349 N_D[1]_M1052_g N_A_824_333#_c_6435_n 0.0127833f $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_1350 N_D[1]_M1097_g N_A_824_333#_c_6435_n 0.0101085f $X=5.945 $Y=1.985 $X2=0
+ $Y2=0
cc_1351 D[1] N_A_824_333#_c_6435_n 0.0323774f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_1352 N_D[1]_c_1542_n N_A_824_333#_c_6435_n 7.13708e-19 $X=6.03 $Y=1.16 $X2=0
+ $Y2=0
cc_1353 D[1] N_A_824_333#_c_6418_n 0.0226682f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_1354 N_D[1]_c_1542_n N_A_824_333#_c_6418_n 9.6385e-19 $X=6.03 $Y=1.16 $X2=0
+ $Y2=0
cc_1355 N_D[1]_M1052_g N_A_824_333#_c_6441_n 0.00246916f $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_1356 N_D[1]_M1097_g N_A_824_333#_c_6441_n 0.00244285f $X=5.945 $Y=1.985 $X2=0
+ $Y2=0
cc_1357 N_D[1]_M1097_g N_A_824_333#_c_6420_n 0.00290175f $X=5.945 $Y=1.985 $X2=0
+ $Y2=0
cc_1358 N_D[1]_M1052_g N_A_824_333#_c_6434_n 0.00595395f $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_1359 N_D[1]_M1074_g N_VGND_c_7781_n 0.00300333f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_1360 N_D[1]_M1105_g N_VGND_c_7781_n 0.0030929f $X=5.92 $Y=0.56 $X2=0 $Y2=0
cc_1361 N_D[1]_M1105_g N_VGND_c_7783_n 0.00430643f $X=5.92 $Y=0.56 $X2=0 $Y2=0
cc_1362 N_D[1]_M1074_g VGND 0.00600262f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_1363 N_D[1]_M1105_g VGND 0.00733187f $X=5.92 $Y=0.56 $X2=0 $Y2=0
cc_1364 N_D[1]_M1074_g N_VGND_c_7829_n 0.00436487f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_1365 N_D[1]_M1074_g N_A_845_69#_c_8341_n 0.0114493f $X=5.5 $Y=0.56 $X2=0
+ $Y2=0
cc_1366 N_D[1]_M1105_g N_A_845_69#_c_8341_n 0.00931728f $X=5.92 $Y=0.56 $X2=0
+ $Y2=0
cc_1367 D[1] N_A_845_69#_c_8341_n 0.0518587f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_1368 N_D[1]_c_1542_n N_A_845_69#_c_8341_n 0.00665175f $X=6.03 $Y=1.16 $X2=0
+ $Y2=0
cc_1369 N_D[1]_M1074_g N_A_845_69#_c_8342_n 0.00114614f $X=5.5 $Y=0.56 $X2=0
+ $Y2=0
cc_1370 N_D[1]_c_1542_n N_A_845_69#_c_8342_n 0.00120541f $X=6.03 $Y=1.16 $X2=0
+ $Y2=0
cc_1371 N_D[1]_M1074_g N_A_845_69#_c_8361_n 5.29024e-19 $X=5.5 $Y=0.56 $X2=0
+ $Y2=0
cc_1372 N_D[1]_M1105_g N_A_845_69#_c_8361_n 0.00633603f $X=5.92 $Y=0.56 $X2=0
+ $Y2=0
cc_1373 D[9] N_D[10]_c_1713_n 0.0231965f $X=6.125 $Y=4.165 $X2=0 $Y2=0
cc_1374 N_D[9]_c_1599_n N_D[10]_c_1713_n 7.85936e-19 $X=6.03 $Y=4.28 $X2=0 $Y2=0
cc_1375 D[9] N_D[10]_c_1714_n 7.85936e-19 $X=6.125 $Y=4.165 $X2=0 $Y2=0
cc_1376 N_D[9]_c_1599_n N_D[10]_c_1714_n 0.00603597f $X=6.03 $Y=4.28 $X2=0 $Y2=0
cc_1377 N_D[9]_M1056_g N_VPWR_c_4251_n 0.00847423f $X=5.475 $Y=3.455 $X2=0 $Y2=0
cc_1378 N_D[9]_M1101_g N_VPWR_c_4251_n 0.00338721f $X=5.945 $Y=3.455 $X2=0 $Y2=0
cc_1379 N_D[9]_M1056_g N_VPWR_c_4384_n 0.00295119f $X=5.475 $Y=3.455 $X2=0 $Y2=0
cc_1380 N_D[9]_M1101_g N_VPWR_c_4384_n 0.00311479f $X=5.945 $Y=3.455 $X2=0 $Y2=0
cc_1381 N_D[9]_M1056_g VPWR 0.00350923f $X=5.475 $Y=3.455 $X2=0 $Y2=0
cc_1382 N_D[9]_M1101_g VPWR 0.00568683f $X=5.945 $Y=3.455 $X2=0 $Y2=0
cc_1383 N_D[9]_M1056_g N_VPWR_c_4282_n 0.00342413f $X=5.475 $Y=3.455 $X2=0 $Y2=0
cc_1384 N_D[9]_M1101_g N_VPWR_c_4283_n 0.0033767f $X=5.945 $Y=3.455 $X2=0 $Y2=0
cc_1385 N_D[9]_M1056_g N_Z_c_5203_n 0.00112534f $X=5.475 $Y=3.455 $X2=0 $Y2=0
cc_1386 N_D[9]_M1026_g N_Z_c_5203_n 8.13311e-19 $X=5.5 $Y=4.88 $X2=0 $Y2=0
cc_1387 D[9] N_Z_c_5203_n 0.00742792f $X=6.125 $Y=4.165 $X2=0 $Y2=0
cc_1388 N_D[9]_c_1599_n N_Z_c_5203_n 0.00583073f $X=6.03 $Y=4.28 $X2=0 $Y2=0
cc_1389 N_D[9]_M1056_g N_Z_c_5245_n 0.0033316f $X=5.475 $Y=3.455 $X2=0 $Y2=0
cc_1390 N_D[9]_M1101_g N_Z_c_5245_n 0.00312829f $X=5.945 $Y=3.455 $X2=0 $Y2=0
cc_1391 D[9] N_Z_c_5245_n 0.00125914f $X=6.125 $Y=4.165 $X2=0 $Y2=0
cc_1392 N_D[9]_M1056_g N_A_824_591#_c_6514_n 0.0127833f $X=5.475 $Y=3.455 $X2=0
+ $Y2=0
cc_1393 N_D[9]_M1101_g N_A_824_591#_c_6514_n 0.0101085f $X=5.945 $Y=3.455 $X2=0
+ $Y2=0
cc_1394 D[9] N_A_824_591#_c_6514_n 0.0550456f $X=6.125 $Y=4.165 $X2=0 $Y2=0
cc_1395 N_D[9]_c_1599_n N_A_824_591#_c_6514_n 0.00167756f $X=6.03 $Y=4.28 $X2=0
+ $Y2=0
cc_1396 N_D[9]_M1056_g N_A_824_591#_c_6534_n 0.00246473f $X=5.475 $Y=3.455 $X2=0
+ $Y2=0
cc_1397 N_D[9]_M1101_g N_A_824_591#_c_6534_n 0.00244285f $X=5.945 $Y=3.455 $X2=0
+ $Y2=0
cc_1398 N_D[9]_M1056_g N_A_824_591#_c_6529_n 0.00531997f $X=5.475 $Y=3.455 $X2=0
+ $Y2=0
cc_1399 N_D[9]_M1101_g N_A_824_591#_c_6518_n 0.00290175f $X=5.945 $Y=3.455 $X2=0
+ $Y2=0
cc_1400 N_D[9]_M1026_g N_VGND_c_7782_n 0.00300333f $X=5.5 $Y=4.88 $X2=0 $Y2=0
cc_1401 N_D[9]_M1059_g N_VGND_c_7782_n 0.0030929f $X=5.92 $Y=4.88 $X2=0 $Y2=0
cc_1402 N_D[9]_M1059_g N_VGND_c_7784_n 0.00430643f $X=5.92 $Y=4.88 $X2=0 $Y2=0
cc_1403 N_D[9]_M1026_g VGND 0.00600262f $X=5.5 $Y=4.88 $X2=0 $Y2=0
cc_1404 N_D[9]_M1059_g VGND 0.00733187f $X=5.92 $Y=4.88 $X2=0 $Y2=0
cc_1405 N_D[9]_M1026_g N_VGND_c_7830_n 0.00436487f $X=5.5 $Y=4.88 $X2=0 $Y2=0
cc_1406 N_D[9]_M1026_g N_A_845_915#_c_8389_n 0.00114614f $X=5.5 $Y=4.88 $X2=0
+ $Y2=0
cc_1407 N_D[9]_c_1599_n N_A_845_915#_c_8389_n 0.00120541f $X=6.03 $Y=4.28 $X2=0
+ $Y2=0
cc_1408 N_D[9]_M1026_g N_A_845_915#_c_8405_n 0.0114493f $X=5.5 $Y=4.88 $X2=0
+ $Y2=0
cc_1409 N_D[9]_M1059_g N_A_845_915#_c_8405_n 0.0084485f $X=5.92 $Y=4.88 $X2=0
+ $Y2=0
cc_1410 D[9] N_A_845_915#_c_8405_n 0.0274027f $X=6.125 $Y=4.165 $X2=0 $Y2=0
cc_1411 N_D[9]_c_1599_n N_A_845_915#_c_8405_n 0.0020061f $X=6.03 $Y=4.28 $X2=0
+ $Y2=0
cc_1412 N_D[9]_M1026_g N_A_845_915#_c_8390_n 5.29024e-19 $X=5.5 $Y=4.88 $X2=0
+ $Y2=0
cc_1413 N_D[9]_M1059_g N_A_845_915#_c_8390_n 0.00720482f $X=5.92 $Y=4.88 $X2=0
+ $Y2=0
cc_1414 D[9] N_A_845_915#_c_8390_n 0.024456f $X=6.125 $Y=4.165 $X2=0 $Y2=0
cc_1415 N_D[9]_c_1599_n N_A_845_915#_c_8390_n 0.00464565f $X=6.03 $Y=4.28 $X2=0
+ $Y2=0
cc_1416 N_D[2]_M1003_g N_D[10]_M1009_g 0.0130744f $X=6.935 $Y=1.985 $X2=0 $Y2=0
cc_1417 N_D[2]_M1120_g N_D[10]_M1126_g 0.0129371f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_1418 N_D[2]_M1120_g N_A_1566_265#_M1005_g 0.025073f $X=7.405 $Y=1.985 $X2=0
+ $Y2=0
cc_1419 N_D[2]_M1120_g N_A_1566_265#_c_1774_n 0.00671996f $X=7.405 $Y=1.985
+ $X2=0 $Y2=0
cc_1420 N_D[2]_M1127_g N_S[2]_c_1935_n 0.0165585f $X=7.38 $Y=0.56 $X2=0 $Y2=0
cc_1421 N_D[2]_M1003_g N_VPWR_c_4252_n 0.00338721f $X=6.935 $Y=1.985 $X2=0 $Y2=0
cc_1422 N_D[2]_M1120_g N_VPWR_c_4252_n 0.00848021f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_1423 N_D[2]_M1003_g N_VPWR_c_4392_n 0.00311479f $X=6.935 $Y=1.985 $X2=0 $Y2=0
cc_1424 N_D[2]_M1120_g N_VPWR_c_4392_n 0.00295119f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_1425 N_D[2]_M1003_g VPWR 0.00568683f $X=6.935 $Y=1.985 $X2=0 $Y2=0
cc_1426 N_D[2]_M1120_g VPWR 0.00350923f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_1427 N_D[2]_M1003_g N_VPWR_c_4283_n 0.0033767f $X=6.935 $Y=1.985 $X2=0 $Y2=0
cc_1428 N_D[2]_M1120_g N_VPWR_c_4284_n 0.00342413f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_1429 N_D[2]_M1003_g N_Z_c_5244_n 0.00312829f $X=6.935 $Y=1.985 $X2=0 $Y2=0
cc_1430 N_D[2]_M1120_g N_Z_c_5244_n 0.0033316f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_1431 N_D[2]_c_1655_n N_Z_c_5244_n 0.00125914f $X=7.19 $Y=1.16 $X2=0 $Y2=0
cc_1432 N_D[2]_M1127_g N_Z_c_5228_n 8.13311e-19 $X=7.38 $Y=0.56 $X2=0 $Y2=0
cc_1433 N_D[2]_M1120_g N_Z_c_5228_n 0.00112534f $X=7.405 $Y=1.985 $X2=0 $Y2=0
cc_1434 N_D[2]_c_1655_n N_Z_c_5228_n 0.00742792f $X=7.19 $Y=1.16 $X2=0 $Y2=0
cc_1435 N_D[2]_c_1656_n N_Z_c_5228_n 0.00583073f $X=7.405 $Y=1.16 $X2=0 $Y2=0
cc_1436 N_D[2]_c_1655_n N_A_1315_297#_c_6605_n 0.0226682f $X=7.19 $Y=1.16 $X2=0
+ $Y2=0
cc_1437 N_D[2]_c_1656_n N_A_1315_297#_c_6605_n 9.6385e-19 $X=7.405 $Y=1.16 $X2=0
+ $Y2=0
cc_1438 N_D[2]_M1003_g N_A_1315_297#_c_6612_n 0.0101085f $X=6.935 $Y=1.985 $X2=0
+ $Y2=0
cc_1439 N_D[2]_M1120_g N_A_1315_297#_c_6612_n 0.0127833f $X=7.405 $Y=1.985 $X2=0
+ $Y2=0
cc_1440 N_D[2]_c_1655_n N_A_1315_297#_c_6612_n 0.0323774f $X=7.19 $Y=1.16 $X2=0
+ $Y2=0
cc_1441 N_D[2]_c_1656_n N_A_1315_297#_c_6612_n 7.13708e-19 $X=7.405 $Y=1.16
+ $X2=0 $Y2=0
cc_1442 N_D[2]_M1003_g N_A_1315_297#_c_6616_n 0.00244285f $X=6.935 $Y=1.985
+ $X2=0 $Y2=0
cc_1443 N_D[2]_M1120_g N_A_1315_297#_c_6616_n 0.00246916f $X=7.405 $Y=1.985
+ $X2=0 $Y2=0
cc_1444 N_D[2]_M1003_g N_A_1315_297#_c_6606_n 0.00290175f $X=6.935 $Y=1.985
+ $X2=0 $Y2=0
cc_1445 N_D[2]_M1120_g N_A_1315_297#_c_6619_n 0.00595395f $X=7.405 $Y=1.985
+ $X2=0 $Y2=0
cc_1446 N_D[2]_M1117_g N_VGND_c_7783_n 0.00430643f $X=6.96 $Y=0.56 $X2=0 $Y2=0
cc_1447 N_D[2]_M1117_g N_VGND_c_7785_n 0.0030929f $X=6.96 $Y=0.56 $X2=0 $Y2=0
cc_1448 N_D[2]_M1127_g N_VGND_c_7785_n 0.00300333f $X=7.38 $Y=0.56 $X2=0 $Y2=0
cc_1449 N_D[2]_M1127_g N_VGND_c_7811_n 0.00436487f $X=7.38 $Y=0.56 $X2=0 $Y2=0
cc_1450 N_D[2]_M1117_g VGND 0.00733187f $X=6.96 $Y=0.56 $X2=0 $Y2=0
cc_1451 N_D[2]_M1127_g VGND 0.00600262f $X=7.38 $Y=0.56 $X2=0 $Y2=0
cc_1452 N_D[2]_M1117_g N_A_1315_47#_c_8437_n 0.00633603f $X=6.96 $Y=0.56 $X2=0
+ $Y2=0
cc_1453 N_D[2]_M1127_g N_A_1315_47#_c_8437_n 5.29024e-19 $X=7.38 $Y=0.56 $X2=0
+ $Y2=0
cc_1454 N_D[2]_M1117_g N_A_1315_47#_c_8434_n 0.0084485f $X=6.96 $Y=0.56 $X2=0
+ $Y2=0
cc_1455 N_D[2]_M1127_g N_A_1315_47#_c_8434_n 0.0125955f $X=7.38 $Y=0.56 $X2=0
+ $Y2=0
cc_1456 N_D[2]_c_1655_n N_A_1315_47#_c_8434_n 0.0274027f $X=7.19 $Y=1.16 $X2=0
+ $Y2=0
cc_1457 N_D[2]_c_1656_n N_A_1315_47#_c_8434_n 0.00321151f $X=7.405 $Y=1.16 $X2=0
+ $Y2=0
cc_1458 N_D[2]_M1117_g N_A_1315_47#_c_8435_n 8.68782e-19 $X=6.96 $Y=0.56 $X2=0
+ $Y2=0
cc_1459 N_D[2]_c_1655_n N_A_1315_47#_c_8435_n 0.024456f $X=7.19 $Y=1.16 $X2=0
+ $Y2=0
cc_1460 N_D[2]_c_1656_n N_A_1315_47#_c_8435_n 0.00464565f $X=7.405 $Y=1.16 $X2=0
+ $Y2=0
cc_1461 N_D[10]_M1126_g N_A_1566_793#_M1044_g 0.0250718f $X=7.405 $Y=3.455 $X2=0
+ $Y2=0
cc_1462 N_D[10]_M1126_g N_A_1566_793#_c_1858_n 0.00671996f $X=7.405 $Y=3.455
+ $X2=0 $Y2=0
cc_1463 N_D[10]_M1109_g N_S[10]_c_1999_n 0.0165585f $X=7.38 $Y=4.88 $X2=-0.19
+ $Y2=-0.24
cc_1464 N_D[10]_M1009_g N_VPWR_c_4253_n 0.00338721f $X=6.935 $Y=3.455 $X2=0
+ $Y2=0
cc_1465 N_D[10]_M1126_g N_VPWR_c_4253_n 0.00847423f $X=7.405 $Y=3.455 $X2=0
+ $Y2=0
cc_1466 N_D[10]_M1009_g N_VPWR_c_4400_n 0.00311479f $X=6.935 $Y=3.455 $X2=0
+ $Y2=0
cc_1467 N_D[10]_M1126_g N_VPWR_c_4400_n 0.00295119f $X=7.405 $Y=3.455 $X2=0
+ $Y2=0
cc_1468 N_D[10]_M1009_g VPWR 0.00568683f $X=6.935 $Y=3.455 $X2=0 $Y2=0
cc_1469 N_D[10]_M1126_g VPWR 0.00350923f $X=7.405 $Y=3.455 $X2=0 $Y2=0
cc_1470 N_D[10]_M1009_g N_VPWR_c_4283_n 0.0033767f $X=6.935 $Y=3.455 $X2=0 $Y2=0
cc_1471 N_D[10]_M1126_g N_VPWR_c_4284_n 0.00342413f $X=7.405 $Y=3.455 $X2=0
+ $Y2=0
cc_1472 N_D[10]_M1109_g N_Z_c_5204_n 8.13311e-19 $X=7.38 $Y=4.88 $X2=0 $Y2=0
cc_1473 N_D[10]_M1126_g N_Z_c_5204_n 0.00112534f $X=7.405 $Y=3.455 $X2=0 $Y2=0
cc_1474 N_D[10]_c_1713_n N_Z_c_5204_n 0.00742792f $X=7.19 $Y=4.28 $X2=0 $Y2=0
cc_1475 N_D[10]_c_1714_n N_Z_c_5204_n 0.00583073f $X=7.405 $Y=4.28 $X2=0 $Y2=0
cc_1476 N_D[10]_M1009_g N_Z_c_5245_n 0.00312829f $X=6.935 $Y=3.455 $X2=0 $Y2=0
cc_1477 N_D[10]_M1126_g N_Z_c_5245_n 0.0033316f $X=7.405 $Y=3.455 $X2=0 $Y2=0
cc_1478 N_D[10]_c_1713_n N_Z_c_5245_n 0.00125914f $X=7.19 $Y=4.28 $X2=0 $Y2=0
cc_1479 N_D[10]_M1009_g N_A_1315_591#_c_6704_n 0.0101085f $X=6.935 $Y=3.455
+ $X2=0 $Y2=0
cc_1480 N_D[10]_M1126_g N_A_1315_591#_c_6704_n 0.0127833f $X=7.405 $Y=3.455
+ $X2=0 $Y2=0
cc_1481 N_D[10]_c_1713_n N_A_1315_591#_c_6704_n 0.0323774f $X=7.19 $Y=4.28 $X2=0
+ $Y2=0
cc_1482 N_D[10]_c_1714_n N_A_1315_591#_c_6704_n 7.13708e-19 $X=7.405 $Y=4.28
+ $X2=0 $Y2=0
cc_1483 N_D[10]_c_1713_n N_A_1315_591#_c_6700_n 0.0226682f $X=7.19 $Y=4.28 $X2=0
+ $Y2=0
cc_1484 N_D[10]_c_1714_n N_A_1315_591#_c_6700_n 9.6385e-19 $X=7.405 $Y=4.28
+ $X2=0 $Y2=0
cc_1485 N_D[10]_M1009_g N_A_1315_591#_c_6710_n 0.00244285f $X=6.935 $Y=3.455
+ $X2=0 $Y2=0
cc_1486 N_D[10]_M1126_g N_A_1315_591#_c_6710_n 0.00246473f $X=7.405 $Y=3.455
+ $X2=0 $Y2=0
cc_1487 N_D[10]_M1126_g N_A_1315_591#_c_6712_n 0.00531997f $X=7.405 $Y=3.455
+ $X2=0 $Y2=0
cc_1488 N_D[10]_M1009_g N_A_1315_591#_c_6703_n 0.00290175f $X=6.935 $Y=3.455
+ $X2=0 $Y2=0
cc_1489 N_D[10]_M1035_g N_VGND_c_7784_n 0.00430643f $X=6.96 $Y=4.88 $X2=0 $Y2=0
cc_1490 N_D[10]_M1035_g N_VGND_c_7786_n 0.0030929f $X=6.96 $Y=4.88 $X2=0 $Y2=0
cc_1491 N_D[10]_M1109_g N_VGND_c_7786_n 0.00300333f $X=7.38 $Y=4.88 $X2=0 $Y2=0
cc_1492 N_D[10]_M1109_g N_VGND_c_7813_n 0.00436487f $X=7.38 $Y=4.88 $X2=0 $Y2=0
cc_1493 N_D[10]_M1035_g VGND 0.00733187f $X=6.96 $Y=4.88 $X2=0 $Y2=0
cc_1494 N_D[10]_M1109_g VGND 0.00600262f $X=7.38 $Y=4.88 $X2=0 $Y2=0
cc_1495 N_D[10]_M1035_g N_A_1315_911#_c_8481_n 0.0084485f $X=6.96 $Y=4.88 $X2=0
+ $Y2=0
cc_1496 N_D[10]_M1109_g N_A_1315_911#_c_8481_n 0.0114493f $X=7.38 $Y=4.88 $X2=0
+ $Y2=0
cc_1497 N_D[10]_c_1713_n N_A_1315_911#_c_8481_n 0.0274027f $X=7.19 $Y=4.28 $X2=0
+ $Y2=0
cc_1498 N_D[10]_c_1714_n N_A_1315_911#_c_8481_n 0.0020061f $X=7.405 $Y=4.28
+ $X2=0 $Y2=0
cc_1499 N_D[10]_M1109_g N_A_1315_911#_c_8478_n 0.00114614f $X=7.38 $Y=4.88 $X2=0
+ $Y2=0
cc_1500 N_D[10]_c_1714_n N_A_1315_911#_c_8478_n 0.00120541f $X=7.405 $Y=4.28
+ $X2=0 $Y2=0
cc_1501 N_D[10]_M1035_g N_A_1315_911#_c_8480_n 0.00720482f $X=6.96 $Y=4.88 $X2=0
+ $Y2=0
cc_1502 N_D[10]_M1109_g N_A_1315_911#_c_8480_n 5.29024e-19 $X=7.38 $Y=4.88 $X2=0
+ $Y2=0
cc_1503 N_D[10]_c_1713_n N_A_1315_911#_c_8480_n 0.024456f $X=7.19 $Y=4.28 $X2=0
+ $Y2=0
cc_1504 N_D[10]_c_1714_n N_A_1315_911#_c_8480_n 0.00464565f $X=7.405 $Y=4.28
+ $X2=0 $Y2=0
cc_1505 N_A_1566_265#_M1005_g N_A_1566_793#_M1044_g 0.0130744f $X=7.93 $Y=2.075
+ $X2=0 $Y2=0
cc_1506 N_A_1566_265#_M1124_g N_A_1566_793#_M1095_g 0.0130744f $X=8.4 $Y=2.075
+ $X2=0 $Y2=0
cc_1507 N_A_1566_265#_c_1774_n N_S[2]_c_1933_n 0.00779314f $X=8.02 $Y=1.4
+ $X2=-0.19 $Y2=-0.24
cc_1508 N_A_1566_265#_c_1773_n N_S[2]_c_1936_n 0.00810157f $X=8.31 $Y=1.4 $X2=0
+ $Y2=0
cc_1509 N_A_1566_265#_c_1769_n N_S[2]_c_1936_n 7.04048e-19 $X=8.87 $Y=1.205
+ $X2=0 $Y2=0
cc_1510 N_A_1566_265#_c_1768_n N_S[2]_c_1938_n 0.0100587f $X=8.87 $Y=0.755 $X2=0
+ $Y2=0
cc_1511 N_A_1566_265#_c_1769_n N_S[2]_c_1938_n 0.00267287f $X=8.87 $Y=1.205
+ $X2=0 $Y2=0
cc_1512 N_A_1566_265#_c_1768_n N_S[2]_c_1939_n 0.0105766f $X=8.87 $Y=0.755 $X2=0
+ $Y2=0
cc_1513 N_A_1566_265#_c_1769_n N_S[2]_c_1939_n 0.0090765f $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_1514 N_A_1566_265#_c_1770_n N_S[2]_c_1939_n 0.00742826f $X=9.155 $Y=1.63
+ $X2=0 $Y2=0
cc_1515 N_A_1566_265#_c_1769_n N_S[2]_c_1940_n 0.00445422f $X=8.87 $Y=1.205
+ $X2=0 $Y2=0
cc_1516 N_A_1566_265#_c_1770_n N_S[2]_c_1940_n 4.25171e-19 $X=9.155 $Y=1.63
+ $X2=0 $Y2=0
cc_1517 N_A_1566_265#_c_1771_n N_S[2]_c_1940_n 0.00920672f $X=8.4 $Y=1.34 $X2=0
+ $Y2=0
cc_1518 N_A_1566_265#_c_1769_n N_S[2]_c_1941_n 0.00205356f $X=8.87 $Y=1.205
+ $X2=0 $Y2=0
cc_1519 N_A_1566_265#_c_1776_n N_S[2]_c_1941_n 0.00861299f $X=9.155 $Y=2.31
+ $X2=0 $Y2=0
cc_1520 N_A_1566_265#_c_1770_n N_S[2]_c_1941_n 0.00828481f $X=9.155 $Y=1.63
+ $X2=0 $Y2=0
cc_1521 N_A_1566_265#_c_1771_n N_S[2]_c_1941_n 0.00692516f $X=8.4 $Y=1.34 $X2=0
+ $Y2=0
cc_1522 N_A_1566_265#_c_1769_n N_S[2]_c_1942_n 0.00149517f $X=8.87 $Y=1.205
+ $X2=0 $Y2=0
cc_1523 N_A_1566_265#_c_1768_n S[2] 0.0061421f $X=8.87 $Y=0.755 $X2=0 $Y2=0
cc_1524 N_A_1566_265#_c_1769_n S[2] 0.0101733f $X=8.87 $Y=1.205 $X2=0 $Y2=0
cc_1525 N_A_1566_265#_c_1770_n S[2] 0.0127184f $X=9.155 $Y=1.63 $X2=0 $Y2=0
cc_1526 N_A_1566_265#_c_1771_n S[2] 3.07062e-19 $X=8.4 $Y=1.34 $X2=0 $Y2=0
cc_1527 N_A_1566_265#_M1005_g N_VPWR_c_4252_n 0.00107878f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_1528 N_A_1566_265#_c_1776_n N_VPWR_c_4254_n 0.0321301f $X=9.155 $Y=2.31 $X2=0
+ $Y2=0
cc_1529 N_A_1566_265#_c_1770_n N_VPWR_c_4254_n 0.00732952f $X=9.155 $Y=1.63
+ $X2=0 $Y2=0
cc_1530 N_A_1566_265#_M1124_g N_VPWR_c_4272_n 8.06528e-19 $X=8.4 $Y=2.075 $X2=0
+ $Y2=0
cc_1531 N_A_1566_265#_c_1776_n N_VPWR_c_4272_n 0.0210596f $X=9.155 $Y=2.31 $X2=0
+ $Y2=0
cc_1532 N_A_1566_265#_M1133_s VPWR 0.00179197f $X=9.03 $Y=1.485 $X2=0 $Y2=0
cc_1533 N_A_1566_265#_M1005_g VPWR 0.00435072f $X=7.93 $Y=2.075 $X2=0 $Y2=0
cc_1534 N_A_1566_265#_M1124_g VPWR 0.0054792f $X=8.4 $Y=2.075 $X2=0 $Y2=0
cc_1535 N_A_1566_265#_c_1776_n VPWR 0.00594162f $X=9.155 $Y=2.31 $X2=0 $Y2=0
cc_1536 N_A_1566_265#_c_1773_n N_Z_c_5214_n 0.00168443f $X=8.31 $Y=1.4 $X2=0
+ $Y2=0
cc_1537 N_A_1566_265#_c_1774_n N_Z_c_5214_n 0.00180308f $X=8.02 $Y=1.4 $X2=0
+ $Y2=0
cc_1538 N_A_1566_265#_c_1769_n N_Z_c_5214_n 0.0033343f $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_1539 N_A_1566_265#_M1005_g N_Z_c_5244_n 0.00404618f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_1540 N_A_1566_265#_M1124_g N_Z_c_5246_n 0.00708998f $X=8.4 $Y=2.075 $X2=0
+ $Y2=0
cc_1541 N_A_1566_265#_c_1776_n N_Z_c_5246_n 0.0308332f $X=9.155 $Y=2.31 $X2=0
+ $Y2=0
cc_1542 N_A_1566_265#_c_1770_n N_Z_c_5246_n 0.0132841f $X=9.155 $Y=1.63 $X2=0
+ $Y2=0
cc_1543 N_A_1566_265#_c_1771_n N_Z_c_5246_n 9.57301e-19 $X=8.4 $Y=1.34 $X2=0
+ $Y2=0
cc_1544 N_A_1566_265#_M1005_g N_Z_c_5426_n 0.00513826f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_1545 N_A_1566_265#_M1005_g N_Z_c_5427_n 0.00978858f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_1546 N_A_1566_265#_c_1773_n N_Z_c_5427_n 8.37785e-19 $X=8.31 $Y=1.4 $X2=0
+ $Y2=0
cc_1547 N_A_1566_265#_M1124_g N_Z_c_5427_n 0.00619657f $X=8.4 $Y=2.075 $X2=0
+ $Y2=0
cc_1548 N_A_1566_265#_M1005_g N_Z_c_5228_n 0.00268051f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_1549 N_A_1566_265#_c_1773_n N_Z_c_5228_n 0.0140957f $X=8.31 $Y=1.4 $X2=0
+ $Y2=0
cc_1550 N_A_1566_265#_M1124_g N_Z_c_5228_n 0.00476154f $X=8.4 $Y=2.075 $X2=0
+ $Y2=0
cc_1551 N_A_1566_265#_c_1769_n N_Z_c_5228_n 0.00967956f $X=8.87 $Y=1.205 $X2=0
+ $Y2=0
cc_1552 N_A_1566_265#_c_1770_n N_Z_c_5228_n 0.0117695f $X=9.155 $Y=1.63 $X2=0
+ $Y2=0
cc_1553 N_A_1566_265#_c_1771_n N_Z_c_5228_n 7.26438e-19 $X=8.4 $Y=1.34 $X2=0
+ $Y2=0
cc_1554 N_A_1566_265#_M1005_g N_Z_c_5436_n 2.61869e-19 $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_1555 N_A_1566_265#_M1005_g N_Z_c_5261_n 0.00455034f $X=7.93 $Y=2.075 $X2=0
+ $Y2=0
cc_1556 N_A_1566_265#_M1124_g N_Z_c_5261_n 0.00462462f $X=8.4 $Y=2.075 $X2=0
+ $Y2=0
cc_1557 N_A_1566_265#_M1005_g N_A_1315_297#_c_6612_n 0.00176121f $X=7.93
+ $Y=2.075 $X2=0 $Y2=0
cc_1558 N_A_1566_265#_M1005_g N_A_1315_297#_c_6621_n 0.00463461f $X=7.93
+ $Y=2.075 $X2=0 $Y2=0
cc_1559 N_A_1566_265#_M1124_g N_A_1315_297#_c_6621_n 0.00334959f $X=8.4 $Y=2.075
+ $X2=0 $Y2=0
cc_1560 N_A_1566_265#_M1005_g N_A_1315_297#_c_6623_n 7.75952e-19 $X=7.93
+ $Y=2.075 $X2=0 $Y2=0
cc_1561 N_A_1566_265#_M1005_g N_A_1315_297#_c_6624_n 0.00415998f $X=7.93
+ $Y=2.075 $X2=0 $Y2=0
cc_1562 N_A_1566_265#_c_1776_n N_A_1315_297#_c_6607_n 0.00738363f $X=9.155
+ $Y=2.31 $X2=0 $Y2=0
cc_1563 N_A_1566_265#_M1124_g N_A_1315_297#_c_6626_n 0.00692695f $X=8.4 $Y=2.075
+ $X2=0 $Y2=0
cc_1564 N_A_1566_265#_M1005_g N_A_1315_297#_c_6619_n 0.00508488f $X=7.93
+ $Y=2.075 $X2=0 $Y2=0
cc_1565 N_A_1566_265#_M1124_g N_A_1315_297#_c_6608_n 0.00550198f $X=8.4 $Y=2.075
+ $X2=0 $Y2=0
cc_1566 N_A_1566_265#_c_1776_n N_A_1315_297#_c_6608_n 0.0413447f $X=9.155
+ $Y=2.31 $X2=0 $Y2=0
cc_1567 N_A_1566_265#_c_1770_n N_A_1315_297#_c_6608_n 0.0132748f $X=9.155
+ $Y=1.63 $X2=0 $Y2=0
cc_1568 N_A_1566_265#_c_1771_n N_A_1315_297#_c_6608_n 0.00133381f $X=8.4 $Y=1.34
+ $X2=0 $Y2=0
cc_1569 N_A_1566_265#_c_1768_n N_VGND_c_7811_n 0.0173492f $X=8.87 $Y=0.755 $X2=0
+ $Y2=0
cc_1570 N_A_1566_265#_M1150_s VGND 0.00250855f $X=9.115 $Y=0.235 $X2=0 $Y2=0
cc_1571 N_A_1566_265#_c_1768_n VGND 0.0186564f $X=8.87 $Y=0.755 $X2=0 $Y2=0
cc_1572 N_A_1566_265#_c_1768_n N_A_1315_47#_c_8436_n 0.00358194f $X=8.87
+ $Y=0.755 $X2=0 $Y2=0
cc_1573 N_A_1566_265#_c_1768_n N_A_1315_47#_c_8447_n 0.0185512f $X=8.87 $Y=0.755
+ $X2=0 $Y2=0
cc_1574 N_A_1566_265#_c_1769_n N_A_1315_47#_c_8447_n 0.00101918f $X=8.87
+ $Y=1.205 $X2=0 $Y2=0
cc_1575 N_A_1566_265#_c_1770_n N_A_1315_47#_c_8447_n 0.00285813f $X=9.155
+ $Y=1.63 $X2=0 $Y2=0
cc_1576 N_A_1566_265#_c_1771_n N_A_1315_47#_c_8447_n 0.00308807f $X=8.4 $Y=1.34
+ $X2=0 $Y2=0
cc_1577 N_A_1566_793#_c_1858_n N_S[10]_c_1999_n 0.00779314f $X=8.02 $Y=4.04
+ $X2=-0.19 $Y2=-0.24
cc_1578 N_A_1566_793#_c_1857_n N_S[10]_c_2002_n 0.00810157f $X=8.31 $Y=4.04
+ $X2=0 $Y2=0
cc_1579 N_A_1566_793#_c_1853_n N_S[10]_c_2002_n 7.04048e-19 $X=8.87 $Y=4.685
+ $X2=0 $Y2=0
cc_1580 N_A_1566_793#_c_1853_n N_S[10]_c_2004_n 0.0127103f $X=8.87 $Y=4.685
+ $X2=0 $Y2=0
cc_1581 N_A_1566_793#_c_1853_n N_S[10]_c_2005_n 0.0196531f $X=8.87 $Y=4.685
+ $X2=0 $Y2=0
cc_1582 N_A_1566_793#_c_1854_n N_S[10]_c_2005_n 0.00742826f $X=9.155 $Y=3.805
+ $X2=0 $Y2=0
cc_1583 N_A_1566_793#_c_1853_n N_S[10]_c_2006_n 0.00445422f $X=8.87 $Y=4.685
+ $X2=0 $Y2=0
cc_1584 N_A_1566_793#_c_1854_n N_S[10]_c_2006_n 4.25171e-19 $X=9.155 $Y=3.805
+ $X2=0 $Y2=0
cc_1585 N_A_1566_793#_c_1855_n N_S[10]_c_2006_n 0.00920672f $X=8.4 $Y=4.1 $X2=0
+ $Y2=0
cc_1586 N_A_1566_793#_c_1854_n N_S[10]_c_2010_n 0.00386817f $X=9.155 $Y=3.805
+ $X2=0 $Y2=0
cc_1587 N_A_1566_793#_c_1861_n N_S[10]_c_2010_n 0.00861299f $X=9.155 $Y=3.13
+ $X2=0 $Y2=0
cc_1588 N_A_1566_793#_c_1855_n N_S[10]_c_2010_n 0.00149275f $X=8.4 $Y=4.1 $X2=0
+ $Y2=0
cc_1589 N_A_1566_793#_c_1853_n N_S[10]_c_2007_n 0.00354873f $X=8.87 $Y=4.685
+ $X2=0 $Y2=0
cc_1590 N_A_1566_793#_c_1854_n N_S[10]_c_2007_n 0.00441664f $X=9.155 $Y=3.805
+ $X2=0 $Y2=0
cc_1591 N_A_1566_793#_c_1855_n N_S[10]_c_2007_n 0.00543241f $X=8.4 $Y=4.1 $X2=0
+ $Y2=0
cc_1592 N_A_1566_793#_c_1853_n S[10] 0.0163154f $X=8.87 $Y=4.685 $X2=0 $Y2=0
cc_1593 N_A_1566_793#_c_1854_n S[10] 0.0127184f $X=9.155 $Y=3.805 $X2=0 $Y2=0
cc_1594 N_A_1566_793#_c_1855_n S[10] 3.07062e-19 $X=8.4 $Y=4.1 $X2=0 $Y2=0
cc_1595 N_A_1566_793#_M1044_g N_VPWR_c_4253_n 0.0013032f $X=7.93 $Y=3.365 $X2=0
+ $Y2=0
cc_1596 N_A_1566_793#_c_1854_n N_VPWR_c_4255_n 0.00732952f $X=9.155 $Y=3.805
+ $X2=0 $Y2=0
cc_1597 N_A_1566_793#_c_1861_n N_VPWR_c_4255_n 0.0321301f $X=9.155 $Y=3.13 $X2=0
+ $Y2=0
cc_1598 N_A_1566_793#_M1095_g N_VPWR_c_4272_n 7.91347e-19 $X=8.4 $Y=3.365 $X2=0
+ $Y2=0
cc_1599 N_A_1566_793#_c_1861_n N_VPWR_c_4272_n 0.0210596f $X=9.155 $Y=3.13 $X2=0
+ $Y2=0
cc_1600 N_A_1566_793#_M1137_s VPWR 0.00179197f $X=9.03 $Y=2.955 $X2=0 $Y2=0
cc_1601 N_A_1566_793#_M1044_g VPWR 0.00434142f $X=7.93 $Y=3.365 $X2=0 $Y2=0
cc_1602 N_A_1566_793#_M1095_g VPWR 0.00546988f $X=8.4 $Y=3.365 $X2=0 $Y2=0
cc_1603 N_A_1566_793#_c_1861_n VPWR 0.00594162f $X=9.155 $Y=3.13 $X2=0 $Y2=0
cc_1604 N_A_1566_793#_M1044_g N_Z_c_5204_n 0.00268051f $X=7.93 $Y=3.365 $X2=0
+ $Y2=0
cc_1605 N_A_1566_793#_c_1857_n N_Z_c_5204_n 0.0140957f $X=8.31 $Y=4.04 $X2=0
+ $Y2=0
cc_1606 N_A_1566_793#_M1095_g N_Z_c_5204_n 0.00476154f $X=8.4 $Y=3.365 $X2=0
+ $Y2=0
cc_1607 N_A_1566_793#_c_1853_n N_Z_c_5204_n 0.00967956f $X=8.87 $Y=4.685 $X2=0
+ $Y2=0
cc_1608 N_A_1566_793#_c_1854_n N_Z_c_5204_n 0.0117695f $X=9.155 $Y=3.805 $X2=0
+ $Y2=0
cc_1609 N_A_1566_793#_c_1855_n N_Z_c_5204_n 7.26438e-19 $X=8.4 $Y=4.1 $X2=0
+ $Y2=0
cc_1610 N_A_1566_793#_c_1857_n N_Z_c_5215_n 0.00168443f $X=8.31 $Y=4.04 $X2=0
+ $Y2=0
cc_1611 N_A_1566_793#_c_1858_n N_Z_c_5215_n 0.00180308f $X=8.02 $Y=4.04 $X2=0
+ $Y2=0
cc_1612 N_A_1566_793#_c_1853_n N_Z_c_5215_n 0.0033343f $X=8.87 $Y=4.685 $X2=0
+ $Y2=0
cc_1613 N_A_1566_793#_M1044_g N_Z_c_5245_n 0.0040431f $X=7.93 $Y=3.365 $X2=0
+ $Y2=0
cc_1614 N_A_1566_793#_M1095_g N_Z_c_5247_n 0.00708682f $X=8.4 $Y=3.365 $X2=0
+ $Y2=0
cc_1615 N_A_1566_793#_c_1854_n N_Z_c_5247_n 0.0132841f $X=9.155 $Y=3.805 $X2=0
+ $Y2=0
cc_1616 N_A_1566_793#_c_1861_n N_Z_c_5247_n 0.0308332f $X=9.155 $Y=3.13 $X2=0
+ $Y2=0
cc_1617 N_A_1566_793#_c_1855_n N_Z_c_5247_n 9.57301e-19 $X=8.4 $Y=4.1 $X2=0
+ $Y2=0
cc_1618 N_A_1566_793#_M1044_g N_Z_c_5453_n 0.00513826f $X=7.93 $Y=3.365 $X2=0
+ $Y2=0
cc_1619 N_A_1566_793#_M1044_g N_Z_c_5427_n 2.61869e-19 $X=7.93 $Y=3.365 $X2=0
+ $Y2=0
cc_1620 N_A_1566_793#_M1044_g N_Z_c_5436_n 0.00978858f $X=7.93 $Y=3.365 $X2=0
+ $Y2=0
cc_1621 N_A_1566_793#_c_1857_n N_Z_c_5436_n 8.37785e-19 $X=8.31 $Y=4.04 $X2=0
+ $Y2=0
cc_1622 N_A_1566_793#_M1095_g N_Z_c_5436_n 0.00619657f $X=8.4 $Y=3.365 $X2=0
+ $Y2=0
cc_1623 N_A_1566_793#_M1044_g N_Z_c_5261_n 0.00455034f $X=7.93 $Y=3.365 $X2=0
+ $Y2=0
cc_1624 N_A_1566_793#_M1095_g N_Z_c_5261_n 0.00462236f $X=8.4 $Y=3.365 $X2=0
+ $Y2=0
cc_1625 N_A_1566_793#_M1044_g N_A_1315_591#_c_6704_n 0.00176121f $X=7.93
+ $Y=3.365 $X2=0 $Y2=0
cc_1626 N_A_1566_793#_M1044_g N_A_1315_591#_c_6715_n 0.00400484f $X=7.93
+ $Y=3.365 $X2=0 $Y2=0
cc_1627 N_A_1566_793#_M1095_g N_A_1315_591#_c_6701_n 0.0124482f $X=8.4 $Y=3.365
+ $X2=0 $Y2=0
cc_1628 N_A_1566_793#_c_1854_n N_A_1315_591#_c_6701_n 0.0132748f $X=9.155
+ $Y=3.805 $X2=0 $Y2=0
cc_1629 N_A_1566_793#_c_1861_n N_A_1315_591#_c_6701_n 0.0413753f $X=9.155
+ $Y=3.13 $X2=0 $Y2=0
cc_1630 N_A_1566_793#_c_1855_n N_A_1315_591#_c_6701_n 0.00133381f $X=8.4 $Y=4.1
+ $X2=0 $Y2=0
cc_1631 N_A_1566_793#_M1044_g N_A_1315_591#_c_6720_n 0.00470988f $X=7.93
+ $Y=3.365 $X2=0 $Y2=0
cc_1632 N_A_1566_793#_M1095_g N_A_1315_591#_c_6720_n 0.00334069f $X=8.4 $Y=3.365
+ $X2=0 $Y2=0
cc_1633 N_A_1566_793#_M1044_g N_A_1315_591#_c_6722_n 7.75952e-19 $X=7.93
+ $Y=3.365 $X2=0 $Y2=0
cc_1634 N_A_1566_793#_M1044_g N_A_1315_591#_c_6712_n 0.00508821f $X=7.93
+ $Y=3.365 $X2=0 $Y2=0
cc_1635 N_A_1566_793#_c_1861_n N_A_1315_591#_c_6702_n 0.00738293f $X=9.155
+ $Y=3.13 $X2=0 $Y2=0
cc_1636 N_A_1566_793#_c_1853_n N_VGND_c_7813_n 0.0173402f $X=8.87 $Y=4.685 $X2=0
+ $Y2=0
cc_1637 N_A_1566_793#_M1033_s VGND 0.00250855f $X=9.115 $Y=4.685 $X2=0 $Y2=0
cc_1638 N_A_1566_793#_c_1853_n VGND 0.0186503f $X=8.87 $Y=4.685 $X2=0 $Y2=0
cc_1639 N_A_1566_793#_c_1853_n N_A_1315_911#_c_8479_n 0.00358194f $X=8.87
+ $Y=4.685 $X2=0 $Y2=0
cc_1640 N_A_1566_793#_c_1853_n N_A_1315_911#_c_8492_n 0.0195704f $X=8.87
+ $Y=4.685 $X2=0 $Y2=0
cc_1641 N_A_1566_793#_c_1854_n N_A_1315_911#_c_8492_n 0.00285813f $X=9.155
+ $Y=3.805 $X2=0 $Y2=0
cc_1642 N_A_1566_793#_c_1855_n N_A_1315_911#_c_8492_n 0.00308807f $X=8.4 $Y=4.1
+ $X2=0 $Y2=0
cc_1643 N_S[2]_c_1941_n N_S[10]_c_2010_n 0.0130744f $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_1644 N_S[2]_c_1942_n N_S[3]_c_2065_n 0.0133556f $X=9.45 $Y=0.845 $X2=-0.19
+ $Y2=-0.24
cc_1645 N_S[2]_c_1941_n N_S[3]_c_2066_n 0.0418422f $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_1646 S[2] N_S[3]_c_2066_n 8.74983e-19 $X=9.345 $Y=1.105 $X2=0 $Y2=0
cc_1647 N_S[2]_c_1941_n S[3] 8.74983e-19 $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_1648 S[2] S[3] 0.0208489f $X=9.345 $Y=1.105 $X2=0 $Y2=0
cc_1649 N_S[2]_c_1941_n N_VPWR_c_4254_n 0.00456891f $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_1650 S[2] N_VPWR_c_4254_n 0.00569857f $X=9.345 $Y=1.105 $X2=0 $Y2=0
cc_1651 N_S[2]_c_1941_n N_VPWR_c_4272_n 0.0035837f $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_1652 N_S[2]_c_1941_n VPWR 0.00710985f $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_1653 N_S[2]_c_1933_n N_Z_c_5214_n 0.00413022f $X=7.9 $Y=0.255 $X2=0 $Y2=0
cc_1654 N_S[2]_c_1936_n N_Z_c_5214_n 0.00495983f $X=8.32 $Y=0.255 $X2=0 $Y2=0
cc_1655 N_S[2]_c_1938_n N_Z_c_5214_n 4.25992e-19 $X=8.805 $Y=0.845 $X2=0 $Y2=0
cc_1656 N_S[2]_c_1941_n N_Z_c_5246_n 0.00513674f $X=9.39 $Y=1.41 $X2=0 $Y2=0
cc_1657 S[2] N_Z_c_5246_n 0.00545567f $X=9.345 $Y=1.105 $X2=0 $Y2=0
cc_1658 N_S[2]_c_1933_n N_Z_c_5228_n 0.00199103f $X=7.9 $Y=0.255 $X2=0 $Y2=0
cc_1659 N_S[2]_c_1936_n N_Z_c_5228_n 0.00133607f $X=8.32 $Y=0.255 $X2=0 $Y2=0
cc_1660 N_S[2]_c_1942_n N_VGND_c_7787_n 0.00330937f $X=9.45 $Y=0.845 $X2=0 $Y2=0
cc_1661 N_S[2]_c_1935_n N_VGND_c_7811_n 0.0271255f $X=7.975 $Y=0.18 $X2=0 $Y2=0
cc_1662 N_S[2]_c_1942_n N_VGND_c_7811_n 0.00585385f $X=9.45 $Y=0.845 $X2=0 $Y2=0
cc_1663 N_S[2]_c_1934_n VGND 0.00642387f $X=8.245 $Y=0.18 $X2=0 $Y2=0
cc_1664 N_S[2]_c_1935_n VGND 0.00474746f $X=7.975 $Y=0.18 $X2=0 $Y2=0
cc_1665 N_S[2]_c_1937_n VGND 0.0193094f $X=8.73 $Y=0.18 $X2=0 $Y2=0
cc_1666 N_S[2]_c_1942_n VGND 0.0111218f $X=9.45 $Y=0.845 $X2=0 $Y2=0
cc_1667 N_S[2]_c_1943_n VGND 0.00366655f $X=8.32 $Y=0.18 $X2=0 $Y2=0
cc_1668 N_S[2]_c_1933_n N_A_1315_47#_c_8434_n 0.00139422f $X=7.9 $Y=0.255 $X2=0
+ $Y2=0
cc_1669 N_S[2]_c_1933_n N_A_1315_47#_c_8436_n 0.0132844f $X=7.9 $Y=0.255 $X2=0
+ $Y2=0
cc_1670 N_S[2]_c_1934_n N_A_1315_47#_c_8436_n 0.00211351f $X=8.245 $Y=0.18 $X2=0
+ $Y2=0
cc_1671 N_S[2]_c_1936_n N_A_1315_47#_c_8436_n 0.0126455f $X=8.32 $Y=0.255 $X2=0
+ $Y2=0
cc_1672 N_S[2]_c_1937_n N_A_1315_47#_c_8436_n 0.00436105f $X=8.73 $Y=0.18 $X2=0
+ $Y2=0
cc_1673 N_S[2]_c_1938_n N_A_1315_47#_c_8436_n 0.00349455f $X=8.805 $Y=0.845
+ $X2=0 $Y2=0
cc_1674 N_S[2]_c_1938_n N_A_1315_47#_c_8447_n 0.00295202f $X=8.805 $Y=0.845
+ $X2=0 $Y2=0
cc_1675 N_S[10]_c_2007_n N_S[11]_c_2128_n 0.0474978f $X=9.45 $Y=4.595 $X2=-0.19
+ $Y2=-0.24
cc_1676 S[10] N_S[11]_c_2128_n 8.74983e-19 $X=9.345 $Y=4.165 $X2=-0.19 $Y2=-0.24
cc_1677 N_S[10]_c_2010_n N_S[11]_c_2139_n 0.00770012f $X=9.39 $Y=4.03 $X2=0
+ $Y2=0
cc_1678 N_S[10]_c_2007_n S[11] 8.74983e-19 $X=9.45 $Y=4.595 $X2=0 $Y2=0
cc_1679 S[10] S[11] 0.0208489f $X=9.345 $Y=4.165 $X2=0 $Y2=0
cc_1680 N_S[10]_c_2010_n N_VPWR_c_4255_n 0.00362951f $X=9.39 $Y=4.03 $X2=0 $Y2=0
cc_1681 N_S[10]_c_2007_n N_VPWR_c_4255_n 9.39395e-19 $X=9.45 $Y=4.595 $X2=0
+ $Y2=0
cc_1682 S[10] N_VPWR_c_4255_n 0.00569857f $X=9.345 $Y=4.165 $X2=0 $Y2=0
cc_1683 N_S[10]_c_2010_n N_VPWR_c_4272_n 0.0035837f $X=9.39 $Y=4.03 $X2=0 $Y2=0
cc_1684 N_S[10]_c_2010_n VPWR 0.00710985f $X=9.39 $Y=4.03 $X2=0 $Y2=0
cc_1685 N_S[10]_c_1999_n N_Z_c_5204_n 0.00199103f $X=7.9 $Y=5.185 $X2=0 $Y2=0
cc_1686 N_S[10]_c_2002_n N_Z_c_5204_n 0.00133607f $X=8.32 $Y=5.185 $X2=0 $Y2=0
cc_1687 N_S[10]_c_1999_n N_Z_c_5215_n 0.00413022f $X=7.9 $Y=5.185 $X2=0 $Y2=0
cc_1688 N_S[10]_c_2002_n N_Z_c_5215_n 0.00495983f $X=8.32 $Y=5.185 $X2=0 $Y2=0
cc_1689 N_S[10]_c_2006_n N_Z_c_5215_n 4.25992e-19 $X=8.88 $Y=4.52 $X2=0 $Y2=0
cc_1690 N_S[10]_c_2010_n N_Z_c_5247_n 0.00477894f $X=9.39 $Y=4.03 $X2=0 $Y2=0
cc_1691 N_S[10]_c_2007_n N_Z_c_5247_n 3.57797e-19 $X=9.45 $Y=4.595 $X2=0 $Y2=0
cc_1692 S[10] N_Z_c_5247_n 0.00545567f $X=9.345 $Y=4.165 $X2=0 $Y2=0
cc_1693 N_S[10]_c_2007_n N_VGND_c_7788_n 0.00330937f $X=9.45 $Y=4.595 $X2=0
+ $Y2=0
cc_1694 N_S[10]_c_2001_n N_VGND_c_7813_n 0.0271255f $X=7.975 $Y=5.26 $X2=0 $Y2=0
cc_1695 N_S[10]_c_2007_n N_VGND_c_7813_n 0.00585385f $X=9.45 $Y=4.595 $X2=0
+ $Y2=0
cc_1696 N_S[10]_c_2000_n VGND 0.00642387f $X=8.245 $Y=5.26 $X2=0 $Y2=0
cc_1697 N_S[10]_c_2001_n VGND 0.00474746f $X=7.975 $Y=5.26 $X2=0 $Y2=0
cc_1698 N_S[10]_c_2003_n VGND 0.0193094f $X=8.73 $Y=5.26 $X2=0 $Y2=0
cc_1699 N_S[10]_c_2007_n VGND 0.0111218f $X=9.45 $Y=4.595 $X2=0 $Y2=0
cc_1700 N_S[10]_c_2008_n VGND 0.00366655f $X=8.32 $Y=5.26 $X2=0 $Y2=0
cc_1701 N_S[10]_c_1999_n N_A_1315_911#_c_8478_n 0.00139422f $X=7.9 $Y=5.185
+ $X2=0 $Y2=0
cc_1702 N_S[10]_c_1999_n N_A_1315_911#_c_8479_n 0.0132844f $X=7.9 $Y=5.185 $X2=0
+ $Y2=0
cc_1703 N_S[10]_c_2000_n N_A_1315_911#_c_8479_n 0.00211351f $X=8.245 $Y=5.26
+ $X2=0 $Y2=0
cc_1704 N_S[10]_c_2002_n N_A_1315_911#_c_8479_n 0.0126455f $X=8.32 $Y=5.185
+ $X2=0 $Y2=0
cc_1705 N_S[10]_c_2003_n N_A_1315_911#_c_8479_n 0.00436105f $X=8.73 $Y=5.26
+ $X2=0 $Y2=0
cc_1706 N_S[10]_c_2004_n N_A_1315_911#_c_8479_n 0.00349455f $X=8.805 $Y=5.185
+ $X2=0 $Y2=0
cc_1707 N_S[10]_c_2004_n N_A_1315_911#_c_8492_n 0.00295202f $X=8.805 $Y=5.185
+ $X2=0 $Y2=0
cc_1708 N_S[3]_c_2066_n N_S[11]_c_2139_n 0.0130744f $X=9.93 $Y=1.41 $X2=0 $Y2=0
cc_1709 N_S[3]_c_2073_n N_A_1989_47#_c_2199_n 0.00779314f $X=11.42 $Y=0.255
+ $X2=0 $Y2=0
cc_1710 N_S[3]_c_2066_n N_A_1989_47#_c_2194_n 0.00692516f $X=9.93 $Y=1.41 $X2=0
+ $Y2=0
cc_1711 N_S[3]_c_2067_n N_A_1989_47#_c_2194_n 0.00920672f $X=10.44 $Y=0.92 $X2=0
+ $Y2=0
cc_1712 N_S[3]_c_2071_n N_A_1989_47#_c_2194_n 0.00810157f $X=11 $Y=0.255 $X2=0
+ $Y2=0
cc_1713 S[3] N_A_1989_47#_c_2194_n 3.07062e-19 $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_1714 N_S[3]_c_2066_n N_A_1989_47#_c_2202_n 0.00861299f $X=9.93 $Y=1.41 $X2=0
+ $Y2=0
cc_1715 N_S[3]_c_2065_n N_A_1989_47#_c_2195_n 0.00149517f $X=9.87 $Y=0.845 $X2=0
+ $Y2=0
cc_1716 N_S[3]_c_2066_n N_A_1989_47#_c_2195_n 0.00205356f $X=9.93 $Y=1.41 $X2=0
+ $Y2=0
cc_1717 N_S[3]_c_2067_n N_A_1989_47#_c_2195_n 0.0135307f $X=10.44 $Y=0.92 $X2=0
+ $Y2=0
cc_1718 N_S[3]_c_2068_n N_A_1989_47#_c_2195_n 0.00267287f $X=10.515 $Y=0.845
+ $X2=0 $Y2=0
cc_1719 N_S[3]_c_2071_n N_A_1989_47#_c_2195_n 7.04048e-19 $X=11 $Y=0.255 $X2=0
+ $Y2=0
cc_1720 S[3] N_A_1989_47#_c_2195_n 0.0101733f $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_1721 N_S[3]_c_2066_n N_A_1989_47#_c_2196_n 0.0105766f $X=9.93 $Y=1.41 $X2=0
+ $Y2=0
cc_1722 N_S[3]_c_2068_n N_A_1989_47#_c_2196_n 0.0100587f $X=10.515 $Y=0.845
+ $X2=0 $Y2=0
cc_1723 S[3] N_A_1989_47#_c_2196_n 0.0061421f $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_1724 N_S[3]_c_2066_n N_A_1989_47#_c_2197_n 0.00828481f $X=9.93 $Y=1.41 $X2=0
+ $Y2=0
cc_1725 N_S[3]_c_2067_n N_A_1989_47#_c_2197_n 0.00785343f $X=10.44 $Y=0.92 $X2=0
+ $Y2=0
cc_1726 S[3] N_A_1989_47#_c_2197_n 0.0127184f $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_1727 N_S[3]_c_2072_n N_D[3]_M1025_g 0.0165585f $X=11.345 $Y=0.18 $X2=0 $Y2=0
cc_1728 N_S[3]_c_2066_n N_VPWR_c_4254_n 0.00456891f $X=9.93 $Y=1.41 $X2=0 $Y2=0
cc_1729 S[3] N_VPWR_c_4254_n 0.00569857f $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_1730 N_S[3]_c_2066_n VPWR 0.00710985f $X=9.93 $Y=1.41 $X2=0 $Y2=0
cc_1731 N_S[3]_c_2066_n N_VPWR_c_4285_n 0.0035837f $X=9.93 $Y=1.41 $X2=0 $Y2=0
cc_1732 N_S[3]_c_2068_n N_Z_c_5216_n 4.25992e-19 $X=10.515 $Y=0.845 $X2=0 $Y2=0
cc_1733 N_S[3]_c_2071_n N_Z_c_5216_n 0.00495983f $X=11 $Y=0.255 $X2=0 $Y2=0
cc_1734 N_S[3]_c_2073_n N_Z_c_5216_n 0.00413022f $X=11.42 $Y=0.255 $X2=0 $Y2=0
cc_1735 N_S[3]_c_2066_n N_Z_c_5246_n 0.00513674f $X=9.93 $Y=1.41 $X2=0 $Y2=0
cc_1736 S[3] N_Z_c_5246_n 0.00545567f $X=9.805 $Y=1.105 $X2=0 $Y2=0
cc_1737 N_S[3]_c_2071_n N_Z_c_5229_n 0.00133607f $X=11 $Y=0.255 $X2=0 $Y2=0
cc_1738 N_S[3]_c_2073_n N_Z_c_5229_n 0.00199103f $X=11.42 $Y=0.255 $X2=0 $Y2=0
cc_1739 N_S[3]_c_2065_n N_VGND_c_7787_n 0.00330937f $X=9.87 $Y=0.845 $X2=0 $Y2=0
cc_1740 N_S[3]_c_2065_n VGND 0.0111218f $X=9.87 $Y=0.845 $X2=0 $Y2=0
cc_1741 N_S[3]_c_2069_n VGND 0.0119932f $X=10.925 $Y=0.18 $X2=0 $Y2=0
cc_1742 N_S[3]_c_2070_n VGND 0.00731624f $X=10.59 $Y=0.18 $X2=0 $Y2=0
cc_1743 N_S[3]_c_2072_n VGND 0.0111713f $X=11.345 $Y=0.18 $X2=0 $Y2=0
cc_1744 N_S[3]_c_2074_n VGND 0.00366655f $X=11 $Y=0.18 $X2=0 $Y2=0
cc_1745 N_S[3]_c_2065_n N_VGND_c_7831_n 0.00585385f $X=9.87 $Y=0.845 $X2=0 $Y2=0
cc_1746 N_S[3]_c_2070_n N_VGND_c_7831_n 0.0271255f $X=10.59 $Y=0.18 $X2=0 $Y2=0
cc_1747 N_S[3]_c_2068_n N_A_2133_69#_c_8526_n 0.00295202f $X=10.515 $Y=0.845
+ $X2=0 $Y2=0
cc_1748 N_S[3]_c_2071_n N_A_2133_69#_c_8522_n 0.0126455f $X=11 $Y=0.255 $X2=0
+ $Y2=0
cc_1749 N_S[3]_c_2072_n N_A_2133_69#_c_8522_n 0.00211351f $X=11.345 $Y=0.18
+ $X2=0 $Y2=0
cc_1750 N_S[3]_c_2073_n N_A_2133_69#_c_8522_n 0.0132844f $X=11.42 $Y=0.255 $X2=0
+ $Y2=0
cc_1751 N_S[3]_c_2068_n N_A_2133_69#_c_8523_n 0.00349455f $X=10.515 $Y=0.845
+ $X2=0 $Y2=0
cc_1752 N_S[3]_c_2069_n N_A_2133_69#_c_8523_n 0.00436105f $X=10.925 $Y=0.18
+ $X2=0 $Y2=0
cc_1753 N_S[3]_c_2073_n N_A_2133_69#_c_8525_n 0.00139422f $X=11.42 $Y=0.255
+ $X2=0 $Y2=0
cc_1754 N_S[11]_c_2135_n N_A_1989_937#_c_2280_n 0.00779314f $X=11.42 $Y=5.185
+ $X2=0 $Y2=0
cc_1755 N_S[11]_c_2128_n N_A_1989_937#_c_2275_n 0.00543241f $X=9.87 $Y=4.595
+ $X2=0 $Y2=0
cc_1756 N_S[11]_c_2139_n N_A_1989_937#_c_2275_n 0.00149275f $X=9.93 $Y=4.03
+ $X2=0 $Y2=0
cc_1757 N_S[11]_c_2129_n N_A_1989_937#_c_2275_n 0.00920672f $X=10.44 $Y=4.52
+ $X2=0 $Y2=0
cc_1758 N_S[11]_c_2133_n N_A_1989_937#_c_2275_n 0.00810157f $X=11 $Y=5.185 $X2=0
+ $Y2=0
cc_1759 S[11] N_A_1989_937#_c_2275_n 3.07062e-19 $X=9.805 $Y=4.165 $X2=0 $Y2=0
cc_1760 N_S[11]_c_2139_n N_A_1989_937#_c_2283_n 0.00861299f $X=9.93 $Y=4.03
+ $X2=0 $Y2=0
cc_1761 N_S[11]_c_2128_n N_A_1989_937#_c_2276_n 0.00354873f $X=9.87 $Y=4.595
+ $X2=0 $Y2=0
cc_1762 N_S[11]_c_2129_n N_A_1989_937#_c_2276_n 0.0135307f $X=10.44 $Y=4.52
+ $X2=0 $Y2=0
cc_1763 N_S[11]_c_2130_n N_A_1989_937#_c_2276_n 0.00267287f $X=10.515 $Y=5.185
+ $X2=0 $Y2=0
cc_1764 N_S[11]_c_2133_n N_A_1989_937#_c_2276_n 7.04048e-19 $X=11 $Y=5.185 $X2=0
+ $Y2=0
cc_1765 S[11] N_A_1989_937#_c_2276_n 0.0101733f $X=9.805 $Y=4.165 $X2=0 $Y2=0
cc_1766 N_S[11]_c_2128_n N_A_1989_937#_c_2277_n 0.0105766f $X=9.87 $Y=4.595
+ $X2=0 $Y2=0
cc_1767 N_S[11]_c_2130_n N_A_1989_937#_c_2277_n 0.0100374f $X=10.515 $Y=5.185
+ $X2=0 $Y2=0
cc_1768 S[11] N_A_1989_937#_c_2277_n 0.0061421f $X=9.805 $Y=4.165 $X2=0 $Y2=0
cc_1769 N_S[11]_c_2128_n N_A_1989_937#_c_2278_n 0.00441664f $X=9.87 $Y=4.595
+ $X2=0 $Y2=0
cc_1770 N_S[11]_c_2139_n N_A_1989_937#_c_2278_n 0.00386817f $X=9.93 $Y=4.03
+ $X2=0 $Y2=0
cc_1771 N_S[11]_c_2129_n N_A_1989_937#_c_2278_n 0.00785343f $X=10.44 $Y=4.52
+ $X2=0 $Y2=0
cc_1772 S[11] N_A_1989_937#_c_2278_n 0.0127184f $X=9.805 $Y=4.165 $X2=0 $Y2=0
cc_1773 N_S[11]_c_2135_n N_D[11]_M1011_g 0.0165585f $X=11.42 $Y=5.185 $X2=0
+ $Y2=0
cc_1774 N_S[11]_c_2128_n N_VPWR_c_4255_n 9.39395e-19 $X=9.87 $Y=4.595 $X2=0
+ $Y2=0
cc_1775 N_S[11]_c_2139_n N_VPWR_c_4255_n 0.00362951f $X=9.93 $Y=4.03 $X2=0 $Y2=0
cc_1776 S[11] N_VPWR_c_4255_n 0.00569857f $X=9.805 $Y=4.165 $X2=0 $Y2=0
cc_1777 N_S[11]_c_2139_n VPWR 0.00710985f $X=9.93 $Y=4.03 $X2=0 $Y2=0
cc_1778 N_S[11]_c_2139_n N_VPWR_c_4285_n 0.0035837f $X=9.93 $Y=4.03 $X2=0 $Y2=0
cc_1779 N_S[11]_c_2133_n N_Z_c_5205_n 0.00133607f $X=11 $Y=5.185 $X2=0 $Y2=0
cc_1780 N_S[11]_c_2135_n N_Z_c_5205_n 0.00199103f $X=11.42 $Y=5.185 $X2=0 $Y2=0
cc_1781 N_S[11]_c_2129_n N_Z_c_5217_n 4.25992e-19 $X=10.44 $Y=4.52 $X2=0 $Y2=0
cc_1782 N_S[11]_c_2133_n N_Z_c_5217_n 0.00495983f $X=11 $Y=5.185 $X2=0 $Y2=0
cc_1783 N_S[11]_c_2135_n N_Z_c_5217_n 0.00413022f $X=11.42 $Y=5.185 $X2=0 $Y2=0
cc_1784 N_S[11]_c_2128_n N_Z_c_5247_n 3.57797e-19 $X=9.87 $Y=4.595 $X2=0 $Y2=0
cc_1785 N_S[11]_c_2139_n N_Z_c_5247_n 0.00477894f $X=9.93 $Y=4.03 $X2=0 $Y2=0
cc_1786 S[11] N_Z_c_5247_n 0.00545567f $X=9.805 $Y=4.165 $X2=0 $Y2=0
cc_1787 N_S[11]_c_2128_n N_VGND_c_7788_n 0.00330937f $X=9.87 $Y=4.595 $X2=0
+ $Y2=0
cc_1788 N_S[11]_c_2128_n VGND 0.0111218f $X=9.87 $Y=4.595 $X2=0 $Y2=0
cc_1789 N_S[11]_c_2131_n VGND 0.0119932f $X=10.925 $Y=5.26 $X2=0 $Y2=0
cc_1790 N_S[11]_c_2132_n VGND 0.00731624f $X=10.59 $Y=5.26 $X2=0 $Y2=0
cc_1791 N_S[11]_c_2134_n VGND 0.0111713f $X=11.345 $Y=5.26 $X2=0 $Y2=0
cc_1792 N_S[11]_c_2136_n VGND 0.00366655f $X=11 $Y=5.26 $X2=0 $Y2=0
cc_1793 N_S[11]_c_2128_n N_VGND_c_7832_n 0.00585385f $X=9.87 $Y=4.595 $X2=0
+ $Y2=0
cc_1794 N_S[11]_c_2132_n N_VGND_c_7832_n 0.0271255f $X=10.59 $Y=5.26 $X2=0 $Y2=0
cc_1795 N_S[11]_c_2130_n N_A_2133_915#_c_8574_n 0.00295202f $X=10.515 $Y=5.185
+ $X2=0 $Y2=0
cc_1796 N_S[11]_c_2133_n N_A_2133_915#_c_8570_n 0.0126455f $X=11 $Y=5.185 $X2=0
+ $Y2=0
cc_1797 N_S[11]_c_2134_n N_A_2133_915#_c_8570_n 0.00211351f $X=11.345 $Y=5.26
+ $X2=0 $Y2=0
cc_1798 N_S[11]_c_2135_n N_A_2133_915#_c_8570_n 0.0132844f $X=11.42 $Y=5.185
+ $X2=0 $Y2=0
cc_1799 N_S[11]_c_2130_n N_A_2133_915#_c_8571_n 0.00349455f $X=10.515 $Y=5.185
+ $X2=0 $Y2=0
cc_1800 N_S[11]_c_2131_n N_A_2133_915#_c_8571_n 0.00436105f $X=10.925 $Y=5.26
+ $X2=0 $Y2=0
cc_1801 N_S[11]_c_2135_n N_A_2133_915#_c_8572_n 0.00139422f $X=11.42 $Y=5.185
+ $X2=0 $Y2=0
cc_1802 N_A_1989_47#_M1004_g N_A_1989_937#_M1045_g 0.0130744f $X=10.92 $Y=2.075
+ $X2=0 $Y2=0
cc_1803 N_A_1989_47#_M1123_g N_A_1989_937#_M1093_g 0.0130744f $X=11.39 $Y=2.075
+ $X2=0 $Y2=0
cc_1804 N_A_1989_47#_c_2199_n N_D[3]_M1002_g 0.00671996f $X=11.3 $Y=1.4 $X2=0
+ $Y2=0
cc_1805 N_A_1989_47#_M1123_g N_D[3]_M1002_g 0.025073f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_1806 N_A_1989_47#_c_2202_n N_VPWR_c_4254_n 0.0321301f $X=10.165 $Y=2.31 $X2=0
+ $Y2=0
cc_1807 N_A_1989_47#_c_2197_n N_VPWR_c_4254_n 0.00732952f $X=10.45 $Y=1.42 $X2=0
+ $Y2=0
cc_1808 N_A_1989_47#_M1123_g N_VPWR_c_4256_n 0.00107878f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_1809 N_A_1989_47#_M1053_d VPWR 0.00179197f $X=10.02 $Y=1.485 $X2=0 $Y2=0
cc_1810 N_A_1989_47#_M1004_g VPWR 0.0054792f $X=10.92 $Y=2.075 $X2=0 $Y2=0
cc_1811 N_A_1989_47#_M1123_g VPWR 0.00435072f $X=11.39 $Y=2.075 $X2=0 $Y2=0
cc_1812 N_A_1989_47#_c_2202_n VPWR 0.00594162f $X=10.165 $Y=2.31 $X2=0 $Y2=0
cc_1813 N_A_1989_47#_M1004_g N_VPWR_c_4285_n 8.06528e-19 $X=10.92 $Y=2.075 $X2=0
+ $Y2=0
cc_1814 N_A_1989_47#_c_2202_n N_VPWR_c_4285_n 0.0210596f $X=10.165 $Y=2.31 $X2=0
+ $Y2=0
cc_1815 N_A_1989_47#_c_2199_n N_Z_c_5216_n 0.00348752f $X=11.3 $Y=1.4 $X2=0
+ $Y2=0
cc_1816 N_A_1989_47#_c_2195_n N_Z_c_5216_n 0.0033343f $X=10.45 $Y=1.205 $X2=0
+ $Y2=0
cc_1817 N_A_1989_47#_M1004_g N_Z_c_5246_n 0.00708998f $X=10.92 $Y=2.075 $X2=0
+ $Y2=0
cc_1818 N_A_1989_47#_c_2194_n N_Z_c_5246_n 9.57301e-19 $X=11.01 $Y=1.4 $X2=0
+ $Y2=0
cc_1819 N_A_1989_47#_c_2202_n N_Z_c_5246_n 0.0308332f $X=10.165 $Y=2.31 $X2=0
+ $Y2=0
cc_1820 N_A_1989_47#_c_2197_n N_Z_c_5246_n 0.0132841f $X=10.45 $Y=1.42 $X2=0
+ $Y2=0
cc_1821 N_A_1989_47#_M1123_g N_Z_c_5248_n 0.00404618f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_1822 N_A_1989_47#_M1123_g N_Z_c_5497_n 0.00513826f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_1823 N_A_1989_47#_M1004_g N_Z_c_5498_n 0.00619657f $X=10.92 $Y=2.075 $X2=0
+ $Y2=0
cc_1824 N_A_1989_47#_c_2199_n N_Z_c_5498_n 8.37785e-19 $X=11.3 $Y=1.4 $X2=0
+ $Y2=0
cc_1825 N_A_1989_47#_M1123_g N_Z_c_5498_n 0.00978858f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_1826 N_A_1989_47#_M1004_g N_Z_c_5229_n 0.00476154f $X=10.92 $Y=2.075 $X2=0
+ $Y2=0
cc_1827 N_A_1989_47#_c_2199_n N_Z_c_5229_n 0.0140957f $X=11.3 $Y=1.4 $X2=0 $Y2=0
cc_1828 N_A_1989_47#_c_2194_n N_Z_c_5229_n 7.26438e-19 $X=11.01 $Y=1.4 $X2=0
+ $Y2=0
cc_1829 N_A_1989_47#_M1123_g N_Z_c_5229_n 0.00268051f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_1830 N_A_1989_47#_c_2195_n N_Z_c_5229_n 0.00967956f $X=10.45 $Y=1.205 $X2=0
+ $Y2=0
cc_1831 N_A_1989_47#_c_2197_n N_Z_c_5229_n 0.0117695f $X=10.45 $Y=1.42 $X2=0
+ $Y2=0
cc_1832 N_A_1989_47#_M1123_g N_Z_c_5507_n 2.61869e-19 $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_1833 N_A_1989_47#_M1004_g N_Z_c_5263_n 0.00462462f $X=10.92 $Y=2.075 $X2=0
+ $Y2=0
cc_1834 N_A_1989_47#_M1123_g N_Z_c_5263_n 0.00455034f $X=11.39 $Y=2.075 $X2=0
+ $Y2=0
cc_1835 N_A_1989_47#_M1123_g N_A_2112_333#_c_6796_n 0.00176121f $X=11.39
+ $Y=2.075 $X2=0 $Y2=0
cc_1836 N_A_1989_47#_M1004_g N_A_2112_333#_c_6797_n 0.00334959f $X=10.92
+ $Y=2.075 $X2=0 $Y2=0
cc_1837 N_A_1989_47#_M1123_g N_A_2112_333#_c_6797_n 0.00463461f $X=11.39
+ $Y=2.075 $X2=0 $Y2=0
cc_1838 N_A_1989_47#_c_2202_n N_A_2112_333#_c_6792_n 0.00738363f $X=10.165
+ $Y=2.31 $X2=0 $Y2=0
cc_1839 N_A_1989_47#_M1123_g N_A_2112_333#_c_6800_n 7.75952e-19 $X=11.39
+ $Y=2.075 $X2=0 $Y2=0
cc_1840 N_A_1989_47#_M1004_g N_A_2112_333#_c_6801_n 0.00692695f $X=10.92
+ $Y=2.075 $X2=0 $Y2=0
cc_1841 N_A_1989_47#_M1123_g N_A_2112_333#_c_6802_n 0.00415998f $X=11.39
+ $Y=2.075 $X2=0 $Y2=0
cc_1842 N_A_1989_47#_M1004_g N_A_2112_333#_c_6794_n 0.00550198f $X=10.92
+ $Y=2.075 $X2=0 $Y2=0
cc_1843 N_A_1989_47#_c_2194_n N_A_2112_333#_c_6794_n 0.00133381f $X=11.01 $Y=1.4
+ $X2=0 $Y2=0
cc_1844 N_A_1989_47#_c_2202_n N_A_2112_333#_c_6794_n 0.0413447f $X=10.165
+ $Y=2.31 $X2=0 $Y2=0
cc_1845 N_A_1989_47#_c_2197_n N_A_2112_333#_c_6794_n 0.0132748f $X=10.45 $Y=1.42
+ $X2=0 $Y2=0
cc_1846 N_A_1989_47#_M1123_g N_A_2112_333#_c_6807_n 0.00508488f $X=11.39
+ $Y=2.075 $X2=0 $Y2=0
cc_1847 N_A_1989_47#_M1019_d VGND 0.00250855f $X=9.945 $Y=0.235 $X2=0 $Y2=0
cc_1848 N_A_1989_47#_c_2196_n VGND 0.0186564f $X=10.08 $Y=0.495 $X2=0 $Y2=0
cc_1849 N_A_1989_47#_c_2196_n N_VGND_c_7831_n 0.0173492f $X=10.08 $Y=0.495 $X2=0
+ $Y2=0
cc_1850 N_A_1989_47#_c_2194_n N_A_2133_69#_c_8526_n 0.00308807f $X=11.01 $Y=1.4
+ $X2=0 $Y2=0
cc_1851 N_A_1989_47#_c_2195_n N_A_2133_69#_c_8526_n 0.00101918f $X=10.45
+ $Y=1.205 $X2=0 $Y2=0
cc_1852 N_A_1989_47#_c_2196_n N_A_2133_69#_c_8526_n 0.0185512f $X=10.08 $Y=0.495
+ $X2=0 $Y2=0
cc_1853 N_A_1989_47#_c_2197_n N_A_2133_69#_c_8526_n 0.00285813f $X=10.45 $Y=1.42
+ $X2=0 $Y2=0
cc_1854 N_A_1989_47#_c_2196_n N_A_2133_69#_c_8523_n 0.00358194f $X=10.08
+ $Y=0.495 $X2=0 $Y2=0
cc_1855 N_A_1989_937#_c_2280_n N_D[11]_M1008_g 0.00671996f $X=11.3 $Y=4.04 $X2=0
+ $Y2=0
cc_1856 N_A_1989_937#_M1093_g N_D[11]_M1008_g 0.0250718f $X=11.39 $Y=3.365 $X2=0
+ $Y2=0
cc_1857 N_A_1989_937#_c_2283_n N_VPWR_c_4255_n 0.0321301f $X=10.165 $Y=3.13
+ $X2=0 $Y2=0
cc_1858 N_A_1989_937#_c_2278_n N_VPWR_c_4255_n 0.00732952f $X=10.45 $Y=4.02
+ $X2=0 $Y2=0
cc_1859 N_A_1989_937#_M1093_g N_VPWR_c_4257_n 0.0013032f $X=11.39 $Y=3.365 $X2=0
+ $Y2=0
cc_1860 N_A_1989_937#_M1060_d VPWR 0.00179197f $X=10.02 $Y=2.955 $X2=0 $Y2=0
cc_1861 N_A_1989_937#_M1045_g VPWR 0.00546988f $X=10.92 $Y=3.365 $X2=0 $Y2=0
cc_1862 N_A_1989_937#_M1093_g VPWR 0.00434142f $X=11.39 $Y=3.365 $X2=0 $Y2=0
cc_1863 N_A_1989_937#_c_2283_n VPWR 0.00594162f $X=10.165 $Y=3.13 $X2=0 $Y2=0
cc_1864 N_A_1989_937#_M1045_g N_VPWR_c_4285_n 7.91347e-19 $X=10.92 $Y=3.365
+ $X2=0 $Y2=0
cc_1865 N_A_1989_937#_c_2283_n N_VPWR_c_4285_n 0.0210596f $X=10.165 $Y=3.13
+ $X2=0 $Y2=0
cc_1866 N_A_1989_937#_M1045_g N_Z_c_5205_n 0.00476154f $X=10.92 $Y=3.365 $X2=0
+ $Y2=0
cc_1867 N_A_1989_937#_c_2280_n N_Z_c_5205_n 0.0140957f $X=11.3 $Y=4.04 $X2=0
+ $Y2=0
cc_1868 N_A_1989_937#_c_2275_n N_Z_c_5205_n 7.26438e-19 $X=11.01 $Y=4.04 $X2=0
+ $Y2=0
cc_1869 N_A_1989_937#_M1093_g N_Z_c_5205_n 0.00268051f $X=11.39 $Y=3.365 $X2=0
+ $Y2=0
cc_1870 N_A_1989_937#_c_2276_n N_Z_c_5205_n 0.00967956f $X=10.45 $Y=4.685 $X2=0
+ $Y2=0
cc_1871 N_A_1989_937#_c_2278_n N_Z_c_5205_n 0.0117695f $X=10.45 $Y=4.02 $X2=0
+ $Y2=0
cc_1872 N_A_1989_937#_c_2280_n N_Z_c_5217_n 0.00348752f $X=11.3 $Y=4.04 $X2=0
+ $Y2=0
cc_1873 N_A_1989_937#_c_2276_n N_Z_c_5217_n 0.0033343f $X=10.45 $Y=4.685 $X2=0
+ $Y2=0
cc_1874 N_A_1989_937#_M1045_g N_Z_c_5247_n 0.00708682f $X=10.92 $Y=3.365 $X2=0
+ $Y2=0
cc_1875 N_A_1989_937#_c_2275_n N_Z_c_5247_n 9.57301e-19 $X=11.01 $Y=4.04 $X2=0
+ $Y2=0
cc_1876 N_A_1989_937#_c_2283_n N_Z_c_5247_n 0.0308332f $X=10.165 $Y=3.13 $X2=0
+ $Y2=0
cc_1877 N_A_1989_937#_c_2278_n N_Z_c_5247_n 0.0132841f $X=10.45 $Y=4.02 $X2=0
+ $Y2=0
cc_1878 N_A_1989_937#_M1093_g N_Z_c_5249_n 0.0040431f $X=11.39 $Y=3.365 $X2=0
+ $Y2=0
cc_1879 N_A_1989_937#_M1093_g N_Z_c_5523_n 0.00513826f $X=11.39 $Y=3.365 $X2=0
+ $Y2=0
cc_1880 N_A_1989_937#_M1093_g N_Z_c_5498_n 2.61869e-19 $X=11.39 $Y=3.365 $X2=0
+ $Y2=0
cc_1881 N_A_1989_937#_M1045_g N_Z_c_5507_n 0.00619657f $X=10.92 $Y=3.365 $X2=0
+ $Y2=0
cc_1882 N_A_1989_937#_c_2280_n N_Z_c_5507_n 8.37785e-19 $X=11.3 $Y=4.04 $X2=0
+ $Y2=0
cc_1883 N_A_1989_937#_M1093_g N_Z_c_5507_n 0.00978858f $X=11.39 $Y=3.365 $X2=0
+ $Y2=0
cc_1884 N_A_1989_937#_M1045_g N_Z_c_5263_n 0.00462236f $X=10.92 $Y=3.365 $X2=0
+ $Y2=0
cc_1885 N_A_1989_937#_M1093_g N_Z_c_5263_n 0.00455034f $X=11.39 $Y=3.365 $X2=0
+ $Y2=0
cc_1886 N_A_1989_937#_M1093_g N_A_2112_591#_c_6892_n 0.00176121f $X=11.39
+ $Y=3.365 $X2=0 $Y2=0
cc_1887 N_A_1989_937#_M1045_g N_A_2112_591#_c_6889_n 0.0124482f $X=10.92
+ $Y=3.365 $X2=0 $Y2=0
cc_1888 N_A_1989_937#_c_2275_n N_A_2112_591#_c_6889_n 0.00133381f $X=11.01
+ $Y=4.04 $X2=0 $Y2=0
cc_1889 N_A_1989_937#_c_2283_n N_A_2112_591#_c_6889_n 0.0413753f $X=10.165
+ $Y=3.13 $X2=0 $Y2=0
cc_1890 N_A_1989_937#_c_2278_n N_A_2112_591#_c_6889_n 0.0132748f $X=10.45
+ $Y=4.02 $X2=0 $Y2=0
cc_1891 N_A_1989_937#_M1093_g N_A_2112_591#_c_6897_n 0.00400484f $X=11.39
+ $Y=3.365 $X2=0 $Y2=0
cc_1892 N_A_1989_937#_M1045_g N_A_2112_591#_c_6898_n 0.00334069f $X=10.92
+ $Y=3.365 $X2=0 $Y2=0
cc_1893 N_A_1989_937#_M1093_g N_A_2112_591#_c_6898_n 0.00470988f $X=11.39
+ $Y=3.365 $X2=0 $Y2=0
cc_1894 N_A_1989_937#_c_2283_n N_A_2112_591#_c_6890_n 0.00738293f $X=10.165
+ $Y=3.13 $X2=0 $Y2=0
cc_1895 N_A_1989_937#_M1093_g N_A_2112_591#_c_6901_n 7.75952e-19 $X=11.39
+ $Y=3.365 $X2=0 $Y2=0
cc_1896 N_A_1989_937#_M1093_g N_A_2112_591#_c_6902_n 0.00508821f $X=11.39
+ $Y=3.365 $X2=0 $Y2=0
cc_1897 N_A_1989_937#_M1071_d VGND 0.00250855f $X=9.945 $Y=4.685 $X2=0 $Y2=0
cc_1898 N_A_1989_937#_c_2277_n VGND 0.0186503f $X=10.08 $Y=4.945 $X2=0 $Y2=0
cc_1899 N_A_1989_937#_c_2277_n N_VGND_c_7832_n 0.0173402f $X=10.08 $Y=4.945
+ $X2=0 $Y2=0
cc_1900 N_A_1989_937#_c_2275_n N_A_2133_915#_c_8574_n 0.00308807f $X=11.01
+ $Y=4.04 $X2=0 $Y2=0
cc_1901 N_A_1989_937#_c_2276_n N_A_2133_915#_c_8574_n 0.00101918f $X=10.45
+ $Y=4.685 $X2=0 $Y2=0
cc_1902 N_A_1989_937#_c_2277_n N_A_2133_915#_c_8574_n 0.0185512f $X=10.08
+ $Y=4.945 $X2=0 $Y2=0
cc_1903 N_A_1989_937#_c_2278_n N_A_2133_915#_c_8574_n 0.00285813f $X=10.45
+ $Y=4.02 $X2=0 $Y2=0
cc_1904 N_A_1989_937#_c_2277_n N_A_2133_915#_c_8571_n 0.00358194f $X=10.08
+ $Y=4.945 $X2=0 $Y2=0
cc_1905 N_D[3]_M1002_g N_D[11]_M1008_g 0.0129371f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_1906 N_D[3]_M1135_g N_D[11]_M1141_g 0.0130744f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_1907 D[3] N_D[4]_c_2474_n 0.0231965f $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_1908 N_D[3]_c_2361_n N_D[4]_c_2474_n 7.85936e-19 $X=12.47 $Y=1.16 $X2=0 $Y2=0
cc_1909 D[3] N_D[4]_c_2475_n 7.85936e-19 $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_1910 N_D[3]_c_2361_n N_D[4]_c_2475_n 0.00603597f $X=12.47 $Y=1.16 $X2=0 $Y2=0
cc_1911 N_D[3]_M1002_g N_VPWR_c_4256_n 0.00848021f $X=11.915 $Y=1.985 $X2=0
+ $Y2=0
cc_1912 N_D[3]_M1135_g N_VPWR_c_4256_n 0.00338721f $X=12.385 $Y=1.985 $X2=0
+ $Y2=0
cc_1913 N_D[3]_M1002_g N_VPWR_c_4462_n 0.00295119f $X=11.915 $Y=1.985 $X2=0
+ $Y2=0
cc_1914 N_D[3]_M1135_g N_VPWR_c_4462_n 0.00311479f $X=12.385 $Y=1.985 $X2=0
+ $Y2=0
cc_1915 N_D[3]_M1002_g VPWR 0.00350923f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_1916 N_D[3]_M1135_g VPWR 0.00568683f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_1917 N_D[3]_M1002_g N_VPWR_c_4286_n 0.00342413f $X=11.915 $Y=1.985 $X2=0
+ $Y2=0
cc_1918 N_D[3]_M1135_g N_VPWR_c_4287_n 0.0033767f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_1919 N_D[3]_M1002_g N_Z_c_5248_n 0.0033316f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_1920 N_D[3]_M1135_g N_Z_c_5248_n 0.00312829f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_1921 D[3] N_Z_c_5248_n 0.00125914f $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_1922 N_D[3]_M1002_g N_Z_c_5229_n 0.00112534f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_1923 N_D[3]_M1025_g N_Z_c_5229_n 8.13311e-19 $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_1924 D[3] N_Z_c_5229_n 0.00742792f $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_1925 N_D[3]_c_2361_n N_Z_c_5229_n 0.00583073f $X=12.47 $Y=1.16 $X2=0 $Y2=0
cc_1926 N_D[3]_M1002_g N_A_2112_333#_c_6808_n 0.0127833f $X=11.915 $Y=1.985
+ $X2=0 $Y2=0
cc_1927 N_D[3]_M1135_g N_A_2112_333#_c_6808_n 0.0101085f $X=12.385 $Y=1.985
+ $X2=0 $Y2=0
cc_1928 D[3] N_A_2112_333#_c_6808_n 0.0323774f $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_1929 N_D[3]_c_2361_n N_A_2112_333#_c_6808_n 7.13708e-19 $X=12.47 $Y=1.16
+ $X2=0 $Y2=0
cc_1930 D[3] N_A_2112_333#_c_6791_n 0.0226682f $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_1931 N_D[3]_c_2361_n N_A_2112_333#_c_6791_n 9.6385e-19 $X=12.47 $Y=1.16 $X2=0
+ $Y2=0
cc_1932 N_D[3]_M1002_g N_A_2112_333#_c_6814_n 0.00246916f $X=11.915 $Y=1.985
+ $X2=0 $Y2=0
cc_1933 N_D[3]_M1135_g N_A_2112_333#_c_6814_n 0.00244285f $X=12.385 $Y=1.985
+ $X2=0 $Y2=0
cc_1934 N_D[3]_M1135_g N_A_2112_333#_c_6793_n 0.00290175f $X=12.385 $Y=1.985
+ $X2=0 $Y2=0
cc_1935 N_D[3]_M1002_g N_A_2112_333#_c_6807_n 0.00595395f $X=11.915 $Y=1.985
+ $X2=0 $Y2=0
cc_1936 N_D[3]_M1025_g N_VGND_c_7789_n 0.00300333f $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_1937 N_D[3]_M1156_g N_VGND_c_7789_n 0.0030929f $X=12.36 $Y=0.56 $X2=0 $Y2=0
cc_1938 N_D[3]_M1156_g N_VGND_c_7791_n 0.00430643f $X=12.36 $Y=0.56 $X2=0 $Y2=0
cc_1939 N_D[3]_M1025_g VGND 0.00600262f $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_1940 N_D[3]_M1156_g VGND 0.00733187f $X=12.36 $Y=0.56 $X2=0 $Y2=0
cc_1941 N_D[3]_M1025_g N_VGND_c_7831_n 0.00436487f $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_1942 N_D[3]_M1025_g N_A_2133_69#_c_8524_n 0.0114493f $X=11.94 $Y=0.56 $X2=0
+ $Y2=0
cc_1943 N_D[3]_M1156_g N_A_2133_69#_c_8524_n 0.00931728f $X=12.36 $Y=0.56 $X2=0
+ $Y2=0
cc_1944 D[3] N_A_2133_69#_c_8524_n 0.0518587f $X=12.565 $Y=1.105 $X2=0 $Y2=0
cc_1945 N_D[3]_c_2361_n N_A_2133_69#_c_8524_n 0.00665175f $X=12.47 $Y=1.16 $X2=0
+ $Y2=0
cc_1946 N_D[3]_M1025_g N_A_2133_69#_c_8525_n 0.00114614f $X=11.94 $Y=0.56 $X2=0
+ $Y2=0
cc_1947 N_D[3]_c_2361_n N_A_2133_69#_c_8525_n 0.00120541f $X=12.47 $Y=1.16 $X2=0
+ $Y2=0
cc_1948 N_D[3]_M1025_g N_A_2133_69#_c_8544_n 5.29024e-19 $X=11.94 $Y=0.56 $X2=0
+ $Y2=0
cc_1949 N_D[3]_M1156_g N_A_2133_69#_c_8544_n 0.00633603f $X=12.36 $Y=0.56 $X2=0
+ $Y2=0
cc_1950 D[11] N_D[12]_c_2532_n 0.0231965f $X=12.565 $Y=4.165 $X2=0 $Y2=0
cc_1951 N_D[11]_c_2418_n N_D[12]_c_2532_n 7.85936e-19 $X=12.47 $Y=4.28 $X2=0
+ $Y2=0
cc_1952 D[11] N_D[12]_c_2533_n 7.85936e-19 $X=12.565 $Y=4.165 $X2=0 $Y2=0
cc_1953 N_D[11]_c_2418_n N_D[12]_c_2533_n 0.00603597f $X=12.47 $Y=4.28 $X2=0
+ $Y2=0
cc_1954 N_D[11]_M1008_g N_VPWR_c_4257_n 0.00847423f $X=11.915 $Y=3.455 $X2=0
+ $Y2=0
cc_1955 N_D[11]_M1141_g N_VPWR_c_4257_n 0.00338721f $X=12.385 $Y=3.455 $X2=0
+ $Y2=0
cc_1956 N_D[11]_M1008_g N_VPWR_c_4470_n 0.00295119f $X=11.915 $Y=3.455 $X2=0
+ $Y2=0
cc_1957 N_D[11]_M1141_g N_VPWR_c_4470_n 0.00311479f $X=12.385 $Y=3.455 $X2=0
+ $Y2=0
cc_1958 N_D[11]_M1008_g VPWR 0.00350923f $X=11.915 $Y=3.455 $X2=0 $Y2=0
cc_1959 N_D[11]_M1141_g VPWR 0.00568683f $X=12.385 $Y=3.455 $X2=0 $Y2=0
cc_1960 N_D[11]_M1008_g N_VPWR_c_4286_n 0.00342413f $X=11.915 $Y=3.455 $X2=0
+ $Y2=0
cc_1961 N_D[11]_M1141_g N_VPWR_c_4287_n 0.0033767f $X=12.385 $Y=3.455 $X2=0
+ $Y2=0
cc_1962 N_D[11]_M1008_g N_Z_c_5205_n 0.00112534f $X=11.915 $Y=3.455 $X2=0 $Y2=0
cc_1963 N_D[11]_M1011_g N_Z_c_5205_n 8.13311e-19 $X=11.94 $Y=4.88 $X2=0 $Y2=0
cc_1964 D[11] N_Z_c_5205_n 0.00742792f $X=12.565 $Y=4.165 $X2=0 $Y2=0
cc_1965 N_D[11]_c_2418_n N_Z_c_5205_n 0.00583073f $X=12.47 $Y=4.28 $X2=0 $Y2=0
cc_1966 N_D[11]_M1008_g N_Z_c_5249_n 0.0033316f $X=11.915 $Y=3.455 $X2=0 $Y2=0
cc_1967 N_D[11]_M1141_g N_Z_c_5249_n 0.00312829f $X=12.385 $Y=3.455 $X2=0 $Y2=0
cc_1968 D[11] N_Z_c_5249_n 0.00125914f $X=12.565 $Y=4.165 $X2=0 $Y2=0
cc_1969 N_D[11]_M1008_g N_A_2112_591#_c_6887_n 0.0127833f $X=11.915 $Y=3.455
+ $X2=0 $Y2=0
cc_1970 N_D[11]_M1141_g N_A_2112_591#_c_6887_n 0.0101085f $X=12.385 $Y=3.455
+ $X2=0 $Y2=0
cc_1971 D[11] N_A_2112_591#_c_6887_n 0.0550456f $X=12.565 $Y=4.165 $X2=0 $Y2=0
cc_1972 N_D[11]_c_2418_n N_A_2112_591#_c_6887_n 0.00167756f $X=12.47 $Y=4.28
+ $X2=0 $Y2=0
cc_1973 N_D[11]_M1008_g N_A_2112_591#_c_6907_n 0.00246473f $X=11.915 $Y=3.455
+ $X2=0 $Y2=0
cc_1974 N_D[11]_M1141_g N_A_2112_591#_c_6907_n 0.00244285f $X=12.385 $Y=3.455
+ $X2=0 $Y2=0
cc_1975 N_D[11]_M1008_g N_A_2112_591#_c_6902_n 0.00531997f $X=11.915 $Y=3.455
+ $X2=0 $Y2=0
cc_1976 N_D[11]_M1141_g N_A_2112_591#_c_6891_n 0.00290175f $X=12.385 $Y=3.455
+ $X2=0 $Y2=0
cc_1977 N_D[11]_M1011_g N_VGND_c_7790_n 0.00300333f $X=11.94 $Y=4.88 $X2=0 $Y2=0
cc_1978 N_D[11]_M1136_g N_VGND_c_7790_n 0.0030929f $X=12.36 $Y=4.88 $X2=0 $Y2=0
cc_1979 N_D[11]_M1136_g N_VGND_c_7792_n 0.00430643f $X=12.36 $Y=4.88 $X2=0 $Y2=0
cc_1980 N_D[11]_M1011_g VGND 0.00600262f $X=11.94 $Y=4.88 $X2=0 $Y2=0
cc_1981 N_D[11]_M1136_g VGND 0.00733187f $X=12.36 $Y=4.88 $X2=0 $Y2=0
cc_1982 N_D[11]_M1011_g N_VGND_c_7832_n 0.00436487f $X=11.94 $Y=4.88 $X2=0 $Y2=0
cc_1983 N_D[11]_M1011_g N_A_2133_915#_c_8572_n 0.00114614f $X=11.94 $Y=4.88
+ $X2=0 $Y2=0
cc_1984 N_D[11]_c_2418_n N_A_2133_915#_c_8572_n 0.00120541f $X=12.47 $Y=4.28
+ $X2=0 $Y2=0
cc_1985 N_D[11]_M1011_g N_A_2133_915#_c_8588_n 0.0114493f $X=11.94 $Y=4.88 $X2=0
+ $Y2=0
cc_1986 N_D[11]_M1136_g N_A_2133_915#_c_8588_n 0.0084485f $X=12.36 $Y=4.88 $X2=0
+ $Y2=0
cc_1987 D[11] N_A_2133_915#_c_8588_n 0.0274027f $X=12.565 $Y=4.165 $X2=0 $Y2=0
cc_1988 N_D[11]_c_2418_n N_A_2133_915#_c_8588_n 0.0020061f $X=12.47 $Y=4.28
+ $X2=0 $Y2=0
cc_1989 N_D[11]_M1011_g N_A_2133_915#_c_8573_n 5.29024e-19 $X=11.94 $Y=4.88
+ $X2=0 $Y2=0
cc_1990 N_D[11]_M1136_g N_A_2133_915#_c_8573_n 0.00720482f $X=12.36 $Y=4.88
+ $X2=0 $Y2=0
cc_1991 D[11] N_A_2133_915#_c_8573_n 0.024456f $X=12.565 $Y=4.165 $X2=0 $Y2=0
cc_1992 N_D[11]_c_2418_n N_A_2133_915#_c_8573_n 0.00464565f $X=12.47 $Y=4.28
+ $X2=0 $Y2=0
cc_1993 N_D[4]_M1030_g N_D[12]_M1038_g 0.0130744f $X=13.375 $Y=1.985 $X2=0 $Y2=0
cc_1994 N_D[4]_M1080_g N_D[12]_M1088_g 0.0129371f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_1995 N_D[4]_M1080_g N_A_2854_265#_M1034_g 0.025073f $X=13.845 $Y=1.985 $X2=0
+ $Y2=0
cc_1996 N_D[4]_M1080_g N_A_2854_265#_c_2593_n 0.00671996f $X=13.845 $Y=1.985
+ $X2=0 $Y2=0
cc_1997 N_D[4]_M1094_g N_S[4]_c_2754_n 0.0165585f $X=13.82 $Y=0.56 $X2=0 $Y2=0
cc_1998 N_D[4]_M1030_g N_VPWR_c_4258_n 0.00338721f $X=13.375 $Y=1.985 $X2=0
+ $Y2=0
cc_1999 N_D[4]_M1080_g N_VPWR_c_4258_n 0.00848021f $X=13.845 $Y=1.985 $X2=0
+ $Y2=0
cc_2000 N_D[4]_M1030_g N_VPWR_c_4478_n 0.00311479f $X=13.375 $Y=1.985 $X2=0
+ $Y2=0
cc_2001 N_D[4]_M1080_g N_VPWR_c_4478_n 0.00295119f $X=13.845 $Y=1.985 $X2=0
+ $Y2=0
cc_2002 N_D[4]_M1030_g VPWR 0.00568683f $X=13.375 $Y=1.985 $X2=0 $Y2=0
cc_2003 N_D[4]_M1080_g VPWR 0.00350923f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_2004 N_D[4]_M1030_g N_VPWR_c_4287_n 0.0033767f $X=13.375 $Y=1.985 $X2=0 $Y2=0
cc_2005 N_D[4]_M1080_g N_VPWR_c_4288_n 0.00342413f $X=13.845 $Y=1.985 $X2=0
+ $Y2=0
cc_2006 N_D[4]_M1030_g N_Z_c_5248_n 0.00312829f $X=13.375 $Y=1.985 $X2=0 $Y2=0
cc_2007 N_D[4]_M1080_g N_Z_c_5248_n 0.0033316f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_2008 N_D[4]_c_2474_n N_Z_c_5248_n 0.00125914f $X=13.63 $Y=1.16 $X2=0 $Y2=0
cc_2009 N_D[4]_M1094_g N_Z_c_5230_n 8.13311e-19 $X=13.82 $Y=0.56 $X2=0 $Y2=0
cc_2010 N_D[4]_M1080_g N_Z_c_5230_n 0.00112534f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_2011 N_D[4]_c_2474_n N_Z_c_5230_n 0.00742792f $X=13.63 $Y=1.16 $X2=0 $Y2=0
cc_2012 N_D[4]_c_2475_n N_Z_c_5230_n 0.00583073f $X=13.845 $Y=1.16 $X2=0 $Y2=0
cc_2013 N_D[4]_c_2474_n N_A_2603_297#_c_6978_n 0.0226682f $X=13.63 $Y=1.16 $X2=0
+ $Y2=0
cc_2014 N_D[4]_c_2475_n N_A_2603_297#_c_6978_n 9.6385e-19 $X=13.845 $Y=1.16
+ $X2=0 $Y2=0
cc_2015 N_D[4]_M1030_g N_A_2603_297#_c_6985_n 0.0101085f $X=13.375 $Y=1.985
+ $X2=0 $Y2=0
cc_2016 N_D[4]_M1080_g N_A_2603_297#_c_6985_n 0.0127833f $X=13.845 $Y=1.985
+ $X2=0 $Y2=0
cc_2017 N_D[4]_c_2474_n N_A_2603_297#_c_6985_n 0.0323774f $X=13.63 $Y=1.16 $X2=0
+ $Y2=0
cc_2018 N_D[4]_c_2475_n N_A_2603_297#_c_6985_n 7.13708e-19 $X=13.845 $Y=1.16
+ $X2=0 $Y2=0
cc_2019 N_D[4]_M1030_g N_A_2603_297#_c_6989_n 0.00244285f $X=13.375 $Y=1.985
+ $X2=0 $Y2=0
cc_2020 N_D[4]_M1080_g N_A_2603_297#_c_6989_n 0.00246916f $X=13.845 $Y=1.985
+ $X2=0 $Y2=0
cc_2021 N_D[4]_M1030_g N_A_2603_297#_c_6979_n 0.00290175f $X=13.375 $Y=1.985
+ $X2=0 $Y2=0
cc_2022 N_D[4]_M1080_g N_A_2603_297#_c_6992_n 0.00595395f $X=13.845 $Y=1.985
+ $X2=0 $Y2=0
cc_2023 N_D[4]_M1057_g N_VGND_c_7791_n 0.00430643f $X=13.4 $Y=0.56 $X2=0 $Y2=0
cc_2024 N_D[4]_M1057_g N_VGND_c_7793_n 0.0030929f $X=13.4 $Y=0.56 $X2=0 $Y2=0
cc_2025 N_D[4]_M1094_g N_VGND_c_7793_n 0.00300333f $X=13.82 $Y=0.56 $X2=0 $Y2=0
cc_2026 N_D[4]_M1094_g N_VGND_c_7815_n 0.00436487f $X=13.82 $Y=0.56 $X2=0 $Y2=0
cc_2027 N_D[4]_M1057_g VGND 0.00733187f $X=13.4 $Y=0.56 $X2=0 $Y2=0
cc_2028 N_D[4]_M1094_g VGND 0.00600262f $X=13.82 $Y=0.56 $X2=0 $Y2=0
cc_2029 N_D[4]_M1057_g N_A_2603_47#_c_8620_n 0.00633603f $X=13.4 $Y=0.56 $X2=0
+ $Y2=0
cc_2030 N_D[4]_M1094_g N_A_2603_47#_c_8620_n 5.29024e-19 $X=13.82 $Y=0.56 $X2=0
+ $Y2=0
cc_2031 N_D[4]_M1057_g N_A_2603_47#_c_8617_n 0.0084485f $X=13.4 $Y=0.56 $X2=0
+ $Y2=0
cc_2032 N_D[4]_M1094_g N_A_2603_47#_c_8617_n 0.0125955f $X=13.82 $Y=0.56 $X2=0
+ $Y2=0
cc_2033 N_D[4]_c_2474_n N_A_2603_47#_c_8617_n 0.0274027f $X=13.63 $Y=1.16 $X2=0
+ $Y2=0
cc_2034 N_D[4]_c_2475_n N_A_2603_47#_c_8617_n 0.00321151f $X=13.845 $Y=1.16
+ $X2=0 $Y2=0
cc_2035 N_D[4]_M1057_g N_A_2603_47#_c_8618_n 8.68782e-19 $X=13.4 $Y=0.56 $X2=0
+ $Y2=0
cc_2036 N_D[4]_c_2474_n N_A_2603_47#_c_8618_n 0.024456f $X=13.63 $Y=1.16 $X2=0
+ $Y2=0
cc_2037 N_D[4]_c_2475_n N_A_2603_47#_c_8618_n 0.00464565f $X=13.845 $Y=1.16
+ $X2=0 $Y2=0
cc_2038 N_D[12]_M1088_g N_A_2854_793#_M1114_g 0.0250718f $X=13.845 $Y=3.455
+ $X2=0 $Y2=0
cc_2039 N_D[12]_M1088_g N_A_2854_793#_c_2677_n 0.00671996f $X=13.845 $Y=3.455
+ $X2=0 $Y2=0
cc_2040 N_D[12]_M1103_g N_S[12]_c_2818_n 0.0165585f $X=13.82 $Y=4.88 $X2=-0.19
+ $Y2=-0.24
cc_2041 N_D[12]_M1038_g N_VPWR_c_4259_n 0.00338721f $X=13.375 $Y=3.455 $X2=0
+ $Y2=0
cc_2042 N_D[12]_M1088_g N_VPWR_c_4259_n 0.00847423f $X=13.845 $Y=3.455 $X2=0
+ $Y2=0
cc_2043 N_D[12]_M1038_g N_VPWR_c_4486_n 0.00311479f $X=13.375 $Y=3.455 $X2=0
+ $Y2=0
cc_2044 N_D[12]_M1088_g N_VPWR_c_4486_n 0.00295119f $X=13.845 $Y=3.455 $X2=0
+ $Y2=0
cc_2045 N_D[12]_M1038_g VPWR 0.00568683f $X=13.375 $Y=3.455 $X2=0 $Y2=0
cc_2046 N_D[12]_M1088_g VPWR 0.00350923f $X=13.845 $Y=3.455 $X2=0 $Y2=0
cc_2047 N_D[12]_M1038_g N_VPWR_c_4287_n 0.0033767f $X=13.375 $Y=3.455 $X2=0
+ $Y2=0
cc_2048 N_D[12]_M1088_g N_VPWR_c_4288_n 0.00342413f $X=13.845 $Y=3.455 $X2=0
+ $Y2=0
cc_2049 N_D[12]_M1103_g N_Z_c_5206_n 8.13311e-19 $X=13.82 $Y=4.88 $X2=0 $Y2=0
cc_2050 N_D[12]_M1088_g N_Z_c_5206_n 0.00112534f $X=13.845 $Y=3.455 $X2=0 $Y2=0
cc_2051 N_D[12]_c_2532_n N_Z_c_5206_n 0.00742792f $X=13.63 $Y=4.28 $X2=0 $Y2=0
cc_2052 N_D[12]_c_2533_n N_Z_c_5206_n 0.00583073f $X=13.845 $Y=4.28 $X2=0 $Y2=0
cc_2053 N_D[12]_M1038_g N_Z_c_5249_n 0.00312829f $X=13.375 $Y=3.455 $X2=0 $Y2=0
cc_2054 N_D[12]_M1088_g N_Z_c_5249_n 0.0033316f $X=13.845 $Y=3.455 $X2=0 $Y2=0
cc_2055 N_D[12]_c_2532_n N_Z_c_5249_n 0.00125914f $X=13.63 $Y=4.28 $X2=0 $Y2=0
cc_2056 N_D[12]_M1038_g N_A_2603_591#_c_7077_n 0.0101085f $X=13.375 $Y=3.455
+ $X2=0 $Y2=0
cc_2057 N_D[12]_M1088_g N_A_2603_591#_c_7077_n 0.0127833f $X=13.845 $Y=3.455
+ $X2=0 $Y2=0
cc_2058 N_D[12]_c_2532_n N_A_2603_591#_c_7077_n 0.0323774f $X=13.63 $Y=4.28
+ $X2=0 $Y2=0
cc_2059 N_D[12]_c_2533_n N_A_2603_591#_c_7077_n 7.13708e-19 $X=13.845 $Y=4.28
+ $X2=0 $Y2=0
cc_2060 N_D[12]_c_2532_n N_A_2603_591#_c_7073_n 0.0226682f $X=13.63 $Y=4.28
+ $X2=0 $Y2=0
cc_2061 N_D[12]_c_2533_n N_A_2603_591#_c_7073_n 9.6385e-19 $X=13.845 $Y=4.28
+ $X2=0 $Y2=0
cc_2062 N_D[12]_M1038_g N_A_2603_591#_c_7083_n 0.00244285f $X=13.375 $Y=3.455
+ $X2=0 $Y2=0
cc_2063 N_D[12]_M1088_g N_A_2603_591#_c_7083_n 0.00246473f $X=13.845 $Y=3.455
+ $X2=0 $Y2=0
cc_2064 N_D[12]_M1088_g N_A_2603_591#_c_7085_n 0.00531997f $X=13.845 $Y=3.455
+ $X2=0 $Y2=0
cc_2065 N_D[12]_M1038_g N_A_2603_591#_c_7076_n 0.00290175f $X=13.375 $Y=3.455
+ $X2=0 $Y2=0
cc_2066 N_D[12]_M1073_g N_VGND_c_7792_n 0.00430643f $X=13.4 $Y=4.88 $X2=0 $Y2=0
cc_2067 N_D[12]_M1073_g N_VGND_c_7794_n 0.0030929f $X=13.4 $Y=4.88 $X2=0 $Y2=0
cc_2068 N_D[12]_M1103_g N_VGND_c_7794_n 0.00300333f $X=13.82 $Y=4.88 $X2=0 $Y2=0
cc_2069 N_D[12]_M1103_g N_VGND_c_7817_n 0.00436487f $X=13.82 $Y=4.88 $X2=0 $Y2=0
cc_2070 N_D[12]_M1073_g VGND 0.00733187f $X=13.4 $Y=4.88 $X2=0 $Y2=0
cc_2071 N_D[12]_M1103_g VGND 0.00600262f $X=13.82 $Y=4.88 $X2=0 $Y2=0
cc_2072 N_D[12]_M1073_g N_A_2603_911#_c_8664_n 0.0084485f $X=13.4 $Y=4.88 $X2=0
+ $Y2=0
cc_2073 N_D[12]_M1103_g N_A_2603_911#_c_8664_n 0.0114493f $X=13.82 $Y=4.88 $X2=0
+ $Y2=0
cc_2074 N_D[12]_c_2532_n N_A_2603_911#_c_8664_n 0.0274027f $X=13.63 $Y=4.28
+ $X2=0 $Y2=0
cc_2075 N_D[12]_c_2533_n N_A_2603_911#_c_8664_n 0.0020061f $X=13.845 $Y=4.28
+ $X2=0 $Y2=0
cc_2076 N_D[12]_M1103_g N_A_2603_911#_c_8661_n 0.00114614f $X=13.82 $Y=4.88
+ $X2=0 $Y2=0
cc_2077 N_D[12]_c_2533_n N_A_2603_911#_c_8661_n 0.00120541f $X=13.845 $Y=4.28
+ $X2=0 $Y2=0
cc_2078 N_D[12]_M1073_g N_A_2603_911#_c_8663_n 0.00720482f $X=13.4 $Y=4.88 $X2=0
+ $Y2=0
cc_2079 N_D[12]_M1103_g N_A_2603_911#_c_8663_n 5.29024e-19 $X=13.82 $Y=4.88
+ $X2=0 $Y2=0
cc_2080 N_D[12]_c_2532_n N_A_2603_911#_c_8663_n 0.024456f $X=13.63 $Y=4.28 $X2=0
+ $Y2=0
cc_2081 N_D[12]_c_2533_n N_A_2603_911#_c_8663_n 0.00464565f $X=13.845 $Y=4.28
+ $X2=0 $Y2=0
cc_2082 N_A_2854_265#_M1034_g N_A_2854_793#_M1114_g 0.0130744f $X=14.37 $Y=2.075
+ $X2=0 $Y2=0
cc_2083 N_A_2854_265#_M1083_g N_A_2854_793#_M1159_g 0.0130744f $X=14.84 $Y=2.075
+ $X2=0 $Y2=0
cc_2084 N_A_2854_265#_c_2593_n N_S[4]_c_2752_n 0.00779314f $X=14.46 $Y=1.4
+ $X2=-0.19 $Y2=-0.24
cc_2085 N_A_2854_265#_c_2592_n N_S[4]_c_2755_n 0.00810157f $X=14.75 $Y=1.4 $X2=0
+ $Y2=0
cc_2086 N_A_2854_265#_c_2588_n N_S[4]_c_2755_n 7.04048e-19 $X=15.31 $Y=1.205
+ $X2=0 $Y2=0
cc_2087 N_A_2854_265#_c_2587_n N_S[4]_c_2757_n 0.0100587f $X=15.31 $Y=0.755
+ $X2=0 $Y2=0
cc_2088 N_A_2854_265#_c_2588_n N_S[4]_c_2757_n 0.00267287f $X=15.31 $Y=1.205
+ $X2=0 $Y2=0
cc_2089 N_A_2854_265#_c_2587_n N_S[4]_c_2758_n 0.0105766f $X=15.31 $Y=0.755
+ $X2=0 $Y2=0
cc_2090 N_A_2854_265#_c_2588_n N_S[4]_c_2758_n 0.0090765f $X=15.31 $Y=1.205
+ $X2=0 $Y2=0
cc_2091 N_A_2854_265#_c_2589_n N_S[4]_c_2758_n 0.00742826f $X=15.595 $Y=1.63
+ $X2=0 $Y2=0
cc_2092 N_A_2854_265#_c_2588_n N_S[4]_c_2759_n 0.00445422f $X=15.31 $Y=1.205
+ $X2=0 $Y2=0
cc_2093 N_A_2854_265#_c_2589_n N_S[4]_c_2759_n 4.25171e-19 $X=15.595 $Y=1.63
+ $X2=0 $Y2=0
cc_2094 N_A_2854_265#_c_2590_n N_S[4]_c_2759_n 0.00920672f $X=14.84 $Y=1.34
+ $X2=0 $Y2=0
cc_2095 N_A_2854_265#_c_2588_n N_S[4]_c_2760_n 0.00205356f $X=15.31 $Y=1.205
+ $X2=0 $Y2=0
cc_2096 N_A_2854_265#_c_2595_n N_S[4]_c_2760_n 0.00861299f $X=15.595 $Y=2.31
+ $X2=0 $Y2=0
cc_2097 N_A_2854_265#_c_2589_n N_S[4]_c_2760_n 0.00828481f $X=15.595 $Y=1.63
+ $X2=0 $Y2=0
cc_2098 N_A_2854_265#_c_2590_n N_S[4]_c_2760_n 0.00692516f $X=14.84 $Y=1.34
+ $X2=0 $Y2=0
cc_2099 N_A_2854_265#_c_2588_n N_S[4]_c_2761_n 0.00149517f $X=15.31 $Y=1.205
+ $X2=0 $Y2=0
cc_2100 N_A_2854_265#_c_2587_n S[4] 0.0061421f $X=15.31 $Y=0.755 $X2=0 $Y2=0
cc_2101 N_A_2854_265#_c_2588_n S[4] 0.0101733f $X=15.31 $Y=1.205 $X2=0 $Y2=0
cc_2102 N_A_2854_265#_c_2589_n S[4] 0.0127184f $X=15.595 $Y=1.63 $X2=0 $Y2=0
cc_2103 N_A_2854_265#_c_2590_n S[4] 3.07062e-19 $X=14.84 $Y=1.34 $X2=0 $Y2=0
cc_2104 N_A_2854_265#_M1034_g N_VPWR_c_4258_n 0.00107878f $X=14.37 $Y=2.075
+ $X2=0 $Y2=0
cc_2105 N_A_2854_265#_c_2595_n N_VPWR_c_4260_n 0.0321301f $X=15.595 $Y=2.31
+ $X2=0 $Y2=0
cc_2106 N_A_2854_265#_c_2589_n N_VPWR_c_4260_n 0.00732952f $X=15.595 $Y=1.63
+ $X2=0 $Y2=0
cc_2107 N_A_2854_265#_M1083_g N_VPWR_c_4274_n 8.06528e-19 $X=14.84 $Y=2.075
+ $X2=0 $Y2=0
cc_2108 N_A_2854_265#_c_2595_n N_VPWR_c_4274_n 0.0210596f $X=15.595 $Y=2.31
+ $X2=0 $Y2=0
cc_2109 N_A_2854_265#_M1001_s VPWR 0.00179197f $X=15.47 $Y=1.485 $X2=0 $Y2=0
cc_2110 N_A_2854_265#_M1034_g VPWR 0.00435072f $X=14.37 $Y=2.075 $X2=0 $Y2=0
cc_2111 N_A_2854_265#_M1083_g VPWR 0.0054792f $X=14.84 $Y=2.075 $X2=0 $Y2=0
cc_2112 N_A_2854_265#_c_2595_n VPWR 0.00594162f $X=15.595 $Y=2.31 $X2=0 $Y2=0
cc_2113 N_A_2854_265#_c_2592_n N_Z_c_5218_n 0.00168443f $X=14.75 $Y=1.4 $X2=0
+ $Y2=0
cc_2114 N_A_2854_265#_c_2593_n N_Z_c_5218_n 0.00180308f $X=14.46 $Y=1.4 $X2=0
+ $Y2=0
cc_2115 N_A_2854_265#_c_2588_n N_Z_c_5218_n 0.0033343f $X=15.31 $Y=1.205 $X2=0
+ $Y2=0
cc_2116 N_A_2854_265#_M1034_g N_Z_c_5248_n 0.00404618f $X=14.37 $Y=2.075 $X2=0
+ $Y2=0
cc_2117 N_A_2854_265#_M1083_g N_Z_c_5250_n 0.00708998f $X=14.84 $Y=2.075 $X2=0
+ $Y2=0
cc_2118 N_A_2854_265#_c_2595_n N_Z_c_5250_n 0.0308332f $X=15.595 $Y=2.31 $X2=0
+ $Y2=0
cc_2119 N_A_2854_265#_c_2589_n N_Z_c_5250_n 0.0132841f $X=15.595 $Y=1.63 $X2=0
+ $Y2=0
cc_2120 N_A_2854_265#_c_2590_n N_Z_c_5250_n 9.57301e-19 $X=14.84 $Y=1.34 $X2=0
+ $Y2=0
cc_2121 N_A_2854_265#_M1034_g N_Z_c_5566_n 0.00513826f $X=14.37 $Y=2.075 $X2=0
+ $Y2=0
cc_2122 N_A_2854_265#_M1034_g N_Z_c_5567_n 0.00978858f $X=14.37 $Y=2.075 $X2=0
+ $Y2=0
cc_2123 N_A_2854_265#_c_2592_n N_Z_c_5567_n 8.37785e-19 $X=14.75 $Y=1.4 $X2=0
+ $Y2=0
cc_2124 N_A_2854_265#_M1083_g N_Z_c_5567_n 0.00619657f $X=14.84 $Y=2.075 $X2=0
+ $Y2=0
cc_2125 N_A_2854_265#_M1034_g N_Z_c_5230_n 0.00268051f $X=14.37 $Y=2.075 $X2=0
+ $Y2=0
cc_2126 N_A_2854_265#_c_2592_n N_Z_c_5230_n 0.0140957f $X=14.75 $Y=1.4 $X2=0
+ $Y2=0
cc_2127 N_A_2854_265#_M1083_g N_Z_c_5230_n 0.00476154f $X=14.84 $Y=2.075 $X2=0
+ $Y2=0
cc_2128 N_A_2854_265#_c_2588_n N_Z_c_5230_n 0.00967956f $X=15.31 $Y=1.205 $X2=0
+ $Y2=0
cc_2129 N_A_2854_265#_c_2589_n N_Z_c_5230_n 0.0117695f $X=15.595 $Y=1.63 $X2=0
+ $Y2=0
cc_2130 N_A_2854_265#_c_2590_n N_Z_c_5230_n 7.26438e-19 $X=14.84 $Y=1.34 $X2=0
+ $Y2=0
cc_2131 N_A_2854_265#_M1034_g N_Z_c_5576_n 2.61869e-19 $X=14.37 $Y=2.075 $X2=0
+ $Y2=0
cc_2132 N_A_2854_265#_M1034_g N_Z_c_5265_n 0.00455034f $X=14.37 $Y=2.075 $X2=0
+ $Y2=0
cc_2133 N_A_2854_265#_M1083_g N_Z_c_5265_n 0.00462462f $X=14.84 $Y=2.075 $X2=0
+ $Y2=0
cc_2134 N_A_2854_265#_M1034_g N_A_2603_297#_c_6985_n 0.00176121f $X=14.37
+ $Y=2.075 $X2=0 $Y2=0
cc_2135 N_A_2854_265#_M1034_g N_A_2603_297#_c_6994_n 0.00463461f $X=14.37
+ $Y=2.075 $X2=0 $Y2=0
cc_2136 N_A_2854_265#_M1083_g N_A_2603_297#_c_6994_n 0.00334959f $X=14.84
+ $Y=2.075 $X2=0 $Y2=0
cc_2137 N_A_2854_265#_M1034_g N_A_2603_297#_c_6996_n 7.75952e-19 $X=14.37
+ $Y=2.075 $X2=0 $Y2=0
cc_2138 N_A_2854_265#_M1034_g N_A_2603_297#_c_6997_n 0.00415998f $X=14.37
+ $Y=2.075 $X2=0 $Y2=0
cc_2139 N_A_2854_265#_c_2595_n N_A_2603_297#_c_6980_n 0.00738363f $X=15.595
+ $Y=2.31 $X2=0 $Y2=0
cc_2140 N_A_2854_265#_M1083_g N_A_2603_297#_c_6999_n 0.00692695f $X=14.84
+ $Y=2.075 $X2=0 $Y2=0
cc_2141 N_A_2854_265#_M1034_g N_A_2603_297#_c_6992_n 0.00508488f $X=14.37
+ $Y=2.075 $X2=0 $Y2=0
cc_2142 N_A_2854_265#_M1083_g N_A_2603_297#_c_6981_n 0.00550198f $X=14.84
+ $Y=2.075 $X2=0 $Y2=0
cc_2143 N_A_2854_265#_c_2595_n N_A_2603_297#_c_6981_n 0.0413447f $X=15.595
+ $Y=2.31 $X2=0 $Y2=0
cc_2144 N_A_2854_265#_c_2589_n N_A_2603_297#_c_6981_n 0.0132748f $X=15.595
+ $Y=1.63 $X2=0 $Y2=0
cc_2145 N_A_2854_265#_c_2590_n N_A_2603_297#_c_6981_n 0.00133381f $X=14.84
+ $Y=1.34 $X2=0 $Y2=0
cc_2146 N_A_2854_265#_c_2587_n N_VGND_c_7815_n 0.0173492f $X=15.31 $Y=0.755
+ $X2=0 $Y2=0
cc_2147 N_A_2854_265#_M1064_s VGND 0.00250855f $X=15.555 $Y=0.235 $X2=0 $Y2=0
cc_2148 N_A_2854_265#_c_2587_n VGND 0.0186564f $X=15.31 $Y=0.755 $X2=0 $Y2=0
cc_2149 N_A_2854_265#_c_2587_n N_A_2603_47#_c_8619_n 0.00358194f $X=15.31
+ $Y=0.755 $X2=0 $Y2=0
cc_2150 N_A_2854_265#_c_2587_n N_A_2603_47#_c_8630_n 0.0185512f $X=15.31
+ $Y=0.755 $X2=0 $Y2=0
cc_2151 N_A_2854_265#_c_2588_n N_A_2603_47#_c_8630_n 0.00101918f $X=15.31
+ $Y=1.205 $X2=0 $Y2=0
cc_2152 N_A_2854_265#_c_2589_n N_A_2603_47#_c_8630_n 0.00285813f $X=15.595
+ $Y=1.63 $X2=0 $Y2=0
cc_2153 N_A_2854_265#_c_2590_n N_A_2603_47#_c_8630_n 0.00308807f $X=14.84
+ $Y=1.34 $X2=0 $Y2=0
cc_2154 N_A_2854_793#_c_2677_n N_S[12]_c_2818_n 0.00779314f $X=14.46 $Y=4.04
+ $X2=-0.19 $Y2=-0.24
cc_2155 N_A_2854_793#_c_2676_n N_S[12]_c_2821_n 0.00810157f $X=14.75 $Y=4.04
+ $X2=0 $Y2=0
cc_2156 N_A_2854_793#_c_2672_n N_S[12]_c_2821_n 7.04048e-19 $X=15.31 $Y=4.685
+ $X2=0 $Y2=0
cc_2157 N_A_2854_793#_c_2672_n N_S[12]_c_2823_n 0.0127103f $X=15.31 $Y=4.685
+ $X2=0 $Y2=0
cc_2158 N_A_2854_793#_c_2672_n N_S[12]_c_2824_n 0.0196531f $X=15.31 $Y=4.685
+ $X2=0 $Y2=0
cc_2159 N_A_2854_793#_c_2673_n N_S[12]_c_2824_n 0.00742826f $X=15.595 $Y=3.805
+ $X2=0 $Y2=0
cc_2160 N_A_2854_793#_c_2672_n N_S[12]_c_2825_n 0.00445422f $X=15.31 $Y=4.685
+ $X2=0 $Y2=0
cc_2161 N_A_2854_793#_c_2673_n N_S[12]_c_2825_n 4.25171e-19 $X=15.595 $Y=3.805
+ $X2=0 $Y2=0
cc_2162 N_A_2854_793#_c_2674_n N_S[12]_c_2825_n 0.00920672f $X=14.84 $Y=4.1
+ $X2=0 $Y2=0
cc_2163 N_A_2854_793#_c_2673_n N_S[12]_c_2829_n 0.00386817f $X=15.595 $Y=3.805
+ $X2=0 $Y2=0
cc_2164 N_A_2854_793#_c_2680_n N_S[12]_c_2829_n 0.00861299f $X=15.595 $Y=3.13
+ $X2=0 $Y2=0
cc_2165 N_A_2854_793#_c_2674_n N_S[12]_c_2829_n 0.00149275f $X=14.84 $Y=4.1
+ $X2=0 $Y2=0
cc_2166 N_A_2854_793#_c_2672_n N_S[12]_c_2826_n 0.00354873f $X=15.31 $Y=4.685
+ $X2=0 $Y2=0
cc_2167 N_A_2854_793#_c_2673_n N_S[12]_c_2826_n 0.00441664f $X=15.595 $Y=3.805
+ $X2=0 $Y2=0
cc_2168 N_A_2854_793#_c_2674_n N_S[12]_c_2826_n 0.00543241f $X=14.84 $Y=4.1
+ $X2=0 $Y2=0
cc_2169 N_A_2854_793#_c_2672_n S[12] 0.0163154f $X=15.31 $Y=4.685 $X2=0 $Y2=0
cc_2170 N_A_2854_793#_c_2673_n S[12] 0.0127184f $X=15.595 $Y=3.805 $X2=0 $Y2=0
cc_2171 N_A_2854_793#_c_2674_n S[12] 3.07062e-19 $X=14.84 $Y=4.1 $X2=0 $Y2=0
cc_2172 N_A_2854_793#_M1114_g N_VPWR_c_4259_n 0.0013032f $X=14.37 $Y=3.365 $X2=0
+ $Y2=0
cc_2173 N_A_2854_793#_c_2673_n N_VPWR_c_4261_n 0.00732952f $X=15.595 $Y=3.805
+ $X2=0 $Y2=0
cc_2174 N_A_2854_793#_c_2680_n N_VPWR_c_4261_n 0.0321301f $X=15.595 $Y=3.13
+ $X2=0 $Y2=0
cc_2175 N_A_2854_793#_M1159_g N_VPWR_c_4274_n 7.91347e-19 $X=14.84 $Y=3.365
+ $X2=0 $Y2=0
cc_2176 N_A_2854_793#_c_2680_n N_VPWR_c_4274_n 0.0210596f $X=15.595 $Y=3.13
+ $X2=0 $Y2=0
cc_2177 N_A_2854_793#_M1007_s VPWR 0.00179197f $X=15.47 $Y=2.955 $X2=0 $Y2=0
cc_2178 N_A_2854_793#_M1114_g VPWR 0.00434142f $X=14.37 $Y=3.365 $X2=0 $Y2=0
cc_2179 N_A_2854_793#_M1159_g VPWR 0.00546988f $X=14.84 $Y=3.365 $X2=0 $Y2=0
cc_2180 N_A_2854_793#_c_2680_n VPWR 0.00594162f $X=15.595 $Y=3.13 $X2=0 $Y2=0
cc_2181 N_A_2854_793#_M1114_g N_Z_c_5206_n 0.00268051f $X=14.37 $Y=3.365 $X2=0
+ $Y2=0
cc_2182 N_A_2854_793#_c_2676_n N_Z_c_5206_n 0.0140957f $X=14.75 $Y=4.04 $X2=0
+ $Y2=0
cc_2183 N_A_2854_793#_M1159_g N_Z_c_5206_n 0.00476154f $X=14.84 $Y=3.365 $X2=0
+ $Y2=0
cc_2184 N_A_2854_793#_c_2672_n N_Z_c_5206_n 0.00967956f $X=15.31 $Y=4.685 $X2=0
+ $Y2=0
cc_2185 N_A_2854_793#_c_2673_n N_Z_c_5206_n 0.0117695f $X=15.595 $Y=3.805 $X2=0
+ $Y2=0
cc_2186 N_A_2854_793#_c_2674_n N_Z_c_5206_n 7.26438e-19 $X=14.84 $Y=4.1 $X2=0
+ $Y2=0
cc_2187 N_A_2854_793#_c_2676_n N_Z_c_5219_n 0.00168443f $X=14.75 $Y=4.04 $X2=0
+ $Y2=0
cc_2188 N_A_2854_793#_c_2677_n N_Z_c_5219_n 0.00180308f $X=14.46 $Y=4.04 $X2=0
+ $Y2=0
cc_2189 N_A_2854_793#_c_2672_n N_Z_c_5219_n 0.0033343f $X=15.31 $Y=4.685 $X2=0
+ $Y2=0
cc_2190 N_A_2854_793#_M1114_g N_Z_c_5249_n 0.0040431f $X=14.37 $Y=3.365 $X2=0
+ $Y2=0
cc_2191 N_A_2854_793#_M1159_g N_Z_c_5251_n 0.00708682f $X=14.84 $Y=3.365 $X2=0
+ $Y2=0
cc_2192 N_A_2854_793#_c_2673_n N_Z_c_5251_n 0.0132841f $X=15.595 $Y=3.805 $X2=0
+ $Y2=0
cc_2193 N_A_2854_793#_c_2680_n N_Z_c_5251_n 0.0308332f $X=15.595 $Y=3.13 $X2=0
+ $Y2=0
cc_2194 N_A_2854_793#_c_2674_n N_Z_c_5251_n 9.57301e-19 $X=14.84 $Y=4.1 $X2=0
+ $Y2=0
cc_2195 N_A_2854_793#_M1114_g N_Z_c_5593_n 0.00513826f $X=14.37 $Y=3.365 $X2=0
+ $Y2=0
cc_2196 N_A_2854_793#_M1114_g N_Z_c_5567_n 2.61869e-19 $X=14.37 $Y=3.365 $X2=0
+ $Y2=0
cc_2197 N_A_2854_793#_M1114_g N_Z_c_5576_n 0.00978858f $X=14.37 $Y=3.365 $X2=0
+ $Y2=0
cc_2198 N_A_2854_793#_c_2676_n N_Z_c_5576_n 8.37785e-19 $X=14.75 $Y=4.04 $X2=0
+ $Y2=0
cc_2199 N_A_2854_793#_M1159_g N_Z_c_5576_n 0.00619657f $X=14.84 $Y=3.365 $X2=0
+ $Y2=0
cc_2200 N_A_2854_793#_M1114_g N_Z_c_5265_n 0.00455034f $X=14.37 $Y=3.365 $X2=0
+ $Y2=0
cc_2201 N_A_2854_793#_M1159_g N_Z_c_5265_n 0.00462236f $X=14.84 $Y=3.365 $X2=0
+ $Y2=0
cc_2202 N_A_2854_793#_M1114_g N_A_2603_591#_c_7077_n 0.00176121f $X=14.37
+ $Y=3.365 $X2=0 $Y2=0
cc_2203 N_A_2854_793#_M1114_g N_A_2603_591#_c_7088_n 0.00400484f $X=14.37
+ $Y=3.365 $X2=0 $Y2=0
cc_2204 N_A_2854_793#_M1159_g N_A_2603_591#_c_7074_n 0.0124482f $X=14.84
+ $Y=3.365 $X2=0 $Y2=0
cc_2205 N_A_2854_793#_c_2673_n N_A_2603_591#_c_7074_n 0.0132748f $X=15.595
+ $Y=3.805 $X2=0 $Y2=0
cc_2206 N_A_2854_793#_c_2680_n N_A_2603_591#_c_7074_n 0.0413753f $X=15.595
+ $Y=3.13 $X2=0 $Y2=0
cc_2207 N_A_2854_793#_c_2674_n N_A_2603_591#_c_7074_n 0.00133381f $X=14.84
+ $Y=4.1 $X2=0 $Y2=0
cc_2208 N_A_2854_793#_M1114_g N_A_2603_591#_c_7093_n 0.00470988f $X=14.37
+ $Y=3.365 $X2=0 $Y2=0
cc_2209 N_A_2854_793#_M1159_g N_A_2603_591#_c_7093_n 0.00334069f $X=14.84
+ $Y=3.365 $X2=0 $Y2=0
cc_2210 N_A_2854_793#_M1114_g N_A_2603_591#_c_7095_n 7.75952e-19 $X=14.37
+ $Y=3.365 $X2=0 $Y2=0
cc_2211 N_A_2854_793#_M1114_g N_A_2603_591#_c_7085_n 0.00508821f $X=14.37
+ $Y=3.365 $X2=0 $Y2=0
cc_2212 N_A_2854_793#_c_2680_n N_A_2603_591#_c_7075_n 0.00738293f $X=15.595
+ $Y=3.13 $X2=0 $Y2=0
cc_2213 N_A_2854_793#_c_2672_n N_VGND_c_7817_n 0.0173402f $X=15.31 $Y=4.685
+ $X2=0 $Y2=0
cc_2214 N_A_2854_793#_M1063_s VGND 0.00250855f $X=15.555 $Y=4.685 $X2=0 $Y2=0
cc_2215 N_A_2854_793#_c_2672_n VGND 0.0186503f $X=15.31 $Y=4.685 $X2=0 $Y2=0
cc_2216 N_A_2854_793#_c_2672_n N_A_2603_911#_c_8662_n 0.00358194f $X=15.31
+ $Y=4.685 $X2=0 $Y2=0
cc_2217 N_A_2854_793#_c_2672_n N_A_2603_911#_c_8675_n 0.0195704f $X=15.31
+ $Y=4.685 $X2=0 $Y2=0
cc_2218 N_A_2854_793#_c_2673_n N_A_2603_911#_c_8675_n 0.00285813f $X=15.595
+ $Y=3.805 $X2=0 $Y2=0
cc_2219 N_A_2854_793#_c_2674_n N_A_2603_911#_c_8675_n 0.00308807f $X=14.84
+ $Y=4.1 $X2=0 $Y2=0
cc_2220 N_S[4]_c_2760_n N_S[12]_c_2829_n 0.0130744f $X=15.83 $Y=1.41 $X2=0 $Y2=0
cc_2221 N_S[4]_c_2761_n N_S[5]_c_2884_n 0.0133556f $X=15.89 $Y=0.845 $X2=-0.19
+ $Y2=-0.24
cc_2222 N_S[4]_c_2760_n N_S[5]_c_2885_n 0.0418422f $X=15.83 $Y=1.41 $X2=0 $Y2=0
cc_2223 S[4] N_S[5]_c_2885_n 8.74983e-19 $X=15.785 $Y=1.105 $X2=0 $Y2=0
cc_2224 N_S[4]_c_2760_n S[5] 8.74983e-19 $X=15.83 $Y=1.41 $X2=0 $Y2=0
cc_2225 S[4] S[5] 0.0208489f $X=15.785 $Y=1.105 $X2=0 $Y2=0
cc_2226 N_S[4]_c_2760_n N_VPWR_c_4260_n 0.00456891f $X=15.83 $Y=1.41 $X2=0 $Y2=0
cc_2227 S[4] N_VPWR_c_4260_n 0.00569857f $X=15.785 $Y=1.105 $X2=0 $Y2=0
cc_2228 N_S[4]_c_2760_n N_VPWR_c_4274_n 0.0035837f $X=15.83 $Y=1.41 $X2=0 $Y2=0
cc_2229 N_S[4]_c_2760_n VPWR 0.00710985f $X=15.83 $Y=1.41 $X2=0 $Y2=0
cc_2230 N_S[4]_c_2752_n N_Z_c_5218_n 0.00413022f $X=14.34 $Y=0.255 $X2=0 $Y2=0
cc_2231 N_S[4]_c_2755_n N_Z_c_5218_n 0.00495983f $X=14.76 $Y=0.255 $X2=0 $Y2=0
cc_2232 N_S[4]_c_2757_n N_Z_c_5218_n 4.25992e-19 $X=15.245 $Y=0.845 $X2=0 $Y2=0
cc_2233 N_S[4]_c_2760_n N_Z_c_5250_n 0.00513674f $X=15.83 $Y=1.41 $X2=0 $Y2=0
cc_2234 S[4] N_Z_c_5250_n 0.00545567f $X=15.785 $Y=1.105 $X2=0 $Y2=0
cc_2235 N_S[4]_c_2752_n N_Z_c_5230_n 0.00199103f $X=14.34 $Y=0.255 $X2=0 $Y2=0
cc_2236 N_S[4]_c_2755_n N_Z_c_5230_n 0.00133607f $X=14.76 $Y=0.255 $X2=0 $Y2=0
cc_2237 N_S[4]_c_2761_n N_VGND_c_7795_n 0.00330937f $X=15.89 $Y=0.845 $X2=0
+ $Y2=0
cc_2238 N_S[4]_c_2754_n N_VGND_c_7815_n 0.0271255f $X=14.415 $Y=0.18 $X2=0 $Y2=0
cc_2239 N_S[4]_c_2761_n N_VGND_c_7815_n 0.00585385f $X=15.89 $Y=0.845 $X2=0
+ $Y2=0
cc_2240 N_S[4]_c_2753_n VGND 0.00642387f $X=14.685 $Y=0.18 $X2=0 $Y2=0
cc_2241 N_S[4]_c_2754_n VGND 0.00474746f $X=14.415 $Y=0.18 $X2=0 $Y2=0
cc_2242 N_S[4]_c_2756_n VGND 0.0193094f $X=15.17 $Y=0.18 $X2=0 $Y2=0
cc_2243 N_S[4]_c_2761_n VGND 0.0111218f $X=15.89 $Y=0.845 $X2=0 $Y2=0
cc_2244 N_S[4]_c_2762_n VGND 0.00366655f $X=14.76 $Y=0.18 $X2=0 $Y2=0
cc_2245 N_S[4]_c_2752_n N_A_2603_47#_c_8617_n 0.00139422f $X=14.34 $Y=0.255
+ $X2=0 $Y2=0
cc_2246 N_S[4]_c_2752_n N_A_2603_47#_c_8619_n 0.0132844f $X=14.34 $Y=0.255 $X2=0
+ $Y2=0
cc_2247 N_S[4]_c_2753_n N_A_2603_47#_c_8619_n 0.00211351f $X=14.685 $Y=0.18
+ $X2=0 $Y2=0
cc_2248 N_S[4]_c_2755_n N_A_2603_47#_c_8619_n 0.0126455f $X=14.76 $Y=0.255 $X2=0
+ $Y2=0
cc_2249 N_S[4]_c_2756_n N_A_2603_47#_c_8619_n 0.00436105f $X=15.17 $Y=0.18 $X2=0
+ $Y2=0
cc_2250 N_S[4]_c_2757_n N_A_2603_47#_c_8619_n 0.00349455f $X=15.245 $Y=0.845
+ $X2=0 $Y2=0
cc_2251 N_S[4]_c_2757_n N_A_2603_47#_c_8630_n 0.00295202f $X=15.245 $Y=0.845
+ $X2=0 $Y2=0
cc_2252 N_S[12]_c_2826_n N_S[13]_c_2947_n 0.0474978f $X=15.89 $Y=4.595 $X2=-0.19
+ $Y2=-0.24
cc_2253 S[12] N_S[13]_c_2947_n 8.74983e-19 $X=15.785 $Y=4.165 $X2=-0.19
+ $Y2=-0.24
cc_2254 N_S[12]_c_2829_n N_S[13]_c_2958_n 0.00770012f $X=15.83 $Y=4.03 $X2=0
+ $Y2=0
cc_2255 N_S[12]_c_2826_n S[13] 8.74983e-19 $X=15.89 $Y=4.595 $X2=0 $Y2=0
cc_2256 S[12] S[13] 0.0208489f $X=15.785 $Y=4.165 $X2=0 $Y2=0
cc_2257 N_S[12]_c_2829_n N_VPWR_c_4261_n 0.00362951f $X=15.83 $Y=4.03 $X2=0
+ $Y2=0
cc_2258 N_S[12]_c_2826_n N_VPWR_c_4261_n 9.39395e-19 $X=15.89 $Y=4.595 $X2=0
+ $Y2=0
cc_2259 S[12] N_VPWR_c_4261_n 0.00569857f $X=15.785 $Y=4.165 $X2=0 $Y2=0
cc_2260 N_S[12]_c_2829_n N_VPWR_c_4274_n 0.0035837f $X=15.83 $Y=4.03 $X2=0 $Y2=0
cc_2261 N_S[12]_c_2829_n VPWR 0.00710985f $X=15.83 $Y=4.03 $X2=0 $Y2=0
cc_2262 N_S[12]_c_2818_n N_Z_c_5206_n 0.00199103f $X=14.34 $Y=5.185 $X2=0 $Y2=0
cc_2263 N_S[12]_c_2821_n N_Z_c_5206_n 0.00133607f $X=14.76 $Y=5.185 $X2=0 $Y2=0
cc_2264 N_S[12]_c_2818_n N_Z_c_5219_n 0.00413022f $X=14.34 $Y=5.185 $X2=0 $Y2=0
cc_2265 N_S[12]_c_2821_n N_Z_c_5219_n 0.00495983f $X=14.76 $Y=5.185 $X2=0 $Y2=0
cc_2266 N_S[12]_c_2825_n N_Z_c_5219_n 4.25992e-19 $X=15.32 $Y=4.52 $X2=0 $Y2=0
cc_2267 N_S[12]_c_2829_n N_Z_c_5251_n 0.00477894f $X=15.83 $Y=4.03 $X2=0 $Y2=0
cc_2268 N_S[12]_c_2826_n N_Z_c_5251_n 3.57797e-19 $X=15.89 $Y=4.595 $X2=0 $Y2=0
cc_2269 S[12] N_Z_c_5251_n 0.00545567f $X=15.785 $Y=4.165 $X2=0 $Y2=0
cc_2270 N_S[12]_c_2826_n N_VGND_c_7796_n 0.00330937f $X=15.89 $Y=4.595 $X2=0
+ $Y2=0
cc_2271 N_S[12]_c_2820_n N_VGND_c_7817_n 0.0271255f $X=14.415 $Y=5.26 $X2=0
+ $Y2=0
cc_2272 N_S[12]_c_2826_n N_VGND_c_7817_n 0.00585385f $X=15.89 $Y=4.595 $X2=0
+ $Y2=0
cc_2273 N_S[12]_c_2819_n VGND 0.00642387f $X=14.685 $Y=5.26 $X2=0 $Y2=0
cc_2274 N_S[12]_c_2820_n VGND 0.00474746f $X=14.415 $Y=5.26 $X2=0 $Y2=0
cc_2275 N_S[12]_c_2822_n VGND 0.0193094f $X=15.17 $Y=5.26 $X2=0 $Y2=0
cc_2276 N_S[12]_c_2826_n VGND 0.0111218f $X=15.89 $Y=4.595 $X2=0 $Y2=0
cc_2277 N_S[12]_c_2827_n VGND 0.00366655f $X=14.76 $Y=5.26 $X2=0 $Y2=0
cc_2278 N_S[12]_c_2818_n N_A_2603_911#_c_8661_n 0.00139422f $X=14.34 $Y=5.185
+ $X2=0 $Y2=0
cc_2279 N_S[12]_c_2818_n N_A_2603_911#_c_8662_n 0.0132844f $X=14.34 $Y=5.185
+ $X2=0 $Y2=0
cc_2280 N_S[12]_c_2819_n N_A_2603_911#_c_8662_n 0.00211351f $X=14.685 $Y=5.26
+ $X2=0 $Y2=0
cc_2281 N_S[12]_c_2821_n N_A_2603_911#_c_8662_n 0.0126455f $X=14.76 $Y=5.185
+ $X2=0 $Y2=0
cc_2282 N_S[12]_c_2822_n N_A_2603_911#_c_8662_n 0.00436105f $X=15.17 $Y=5.26
+ $X2=0 $Y2=0
cc_2283 N_S[12]_c_2823_n N_A_2603_911#_c_8662_n 0.00349455f $X=15.245 $Y=5.185
+ $X2=0 $Y2=0
cc_2284 N_S[12]_c_2823_n N_A_2603_911#_c_8675_n 0.00295202f $X=15.245 $Y=5.185
+ $X2=0 $Y2=0
cc_2285 N_S[5]_c_2885_n N_S[13]_c_2958_n 0.0130744f $X=16.37 $Y=1.41 $X2=0 $Y2=0
cc_2286 N_S[5]_c_2892_n N_A_3277_47#_c_3018_n 0.00779314f $X=17.86 $Y=0.255
+ $X2=0 $Y2=0
cc_2287 N_S[5]_c_2885_n N_A_3277_47#_c_3013_n 0.00692516f $X=16.37 $Y=1.41 $X2=0
+ $Y2=0
cc_2288 N_S[5]_c_2886_n N_A_3277_47#_c_3013_n 0.00920672f $X=16.88 $Y=0.92 $X2=0
+ $Y2=0
cc_2289 N_S[5]_c_2890_n N_A_3277_47#_c_3013_n 0.00810157f $X=17.44 $Y=0.255
+ $X2=0 $Y2=0
cc_2290 S[5] N_A_3277_47#_c_3013_n 3.07062e-19 $X=16.245 $Y=1.105 $X2=0 $Y2=0
cc_2291 N_S[5]_c_2885_n N_A_3277_47#_c_3021_n 0.00861299f $X=16.37 $Y=1.41 $X2=0
+ $Y2=0
cc_2292 N_S[5]_c_2884_n N_A_3277_47#_c_3014_n 0.00149517f $X=16.31 $Y=0.845
+ $X2=0 $Y2=0
cc_2293 N_S[5]_c_2885_n N_A_3277_47#_c_3014_n 0.00205356f $X=16.37 $Y=1.41 $X2=0
+ $Y2=0
cc_2294 N_S[5]_c_2886_n N_A_3277_47#_c_3014_n 0.0135307f $X=16.88 $Y=0.92 $X2=0
+ $Y2=0
cc_2295 N_S[5]_c_2887_n N_A_3277_47#_c_3014_n 0.00267287f $X=16.955 $Y=0.845
+ $X2=0 $Y2=0
cc_2296 N_S[5]_c_2890_n N_A_3277_47#_c_3014_n 7.04048e-19 $X=17.44 $Y=0.255
+ $X2=0 $Y2=0
cc_2297 S[5] N_A_3277_47#_c_3014_n 0.0101733f $X=16.245 $Y=1.105 $X2=0 $Y2=0
cc_2298 N_S[5]_c_2885_n N_A_3277_47#_c_3015_n 0.0105766f $X=16.37 $Y=1.41 $X2=0
+ $Y2=0
cc_2299 N_S[5]_c_2887_n N_A_3277_47#_c_3015_n 0.0100587f $X=16.955 $Y=0.845
+ $X2=0 $Y2=0
cc_2300 S[5] N_A_3277_47#_c_3015_n 0.0061421f $X=16.245 $Y=1.105 $X2=0 $Y2=0
cc_2301 N_S[5]_c_2885_n N_A_3277_47#_c_3016_n 0.00828481f $X=16.37 $Y=1.41 $X2=0
+ $Y2=0
cc_2302 N_S[5]_c_2886_n N_A_3277_47#_c_3016_n 0.00785343f $X=16.88 $Y=0.92 $X2=0
+ $Y2=0
cc_2303 S[5] N_A_3277_47#_c_3016_n 0.0127184f $X=16.245 $Y=1.105 $X2=0 $Y2=0
cc_2304 N_S[5]_c_2891_n N_D[5]_M1090_g 0.0165585f $X=17.785 $Y=0.18 $X2=0 $Y2=0
cc_2305 N_S[5]_c_2885_n N_VPWR_c_4260_n 0.00456891f $X=16.37 $Y=1.41 $X2=0 $Y2=0
cc_2306 S[5] N_VPWR_c_4260_n 0.00569857f $X=16.245 $Y=1.105 $X2=0 $Y2=0
cc_2307 N_S[5]_c_2885_n VPWR 0.00710985f $X=16.37 $Y=1.41 $X2=0 $Y2=0
cc_2308 N_S[5]_c_2885_n N_VPWR_c_4289_n 0.0035837f $X=16.37 $Y=1.41 $X2=0 $Y2=0
cc_2309 N_S[5]_c_2887_n N_Z_c_5220_n 4.25992e-19 $X=16.955 $Y=0.845 $X2=0 $Y2=0
cc_2310 N_S[5]_c_2890_n N_Z_c_5220_n 0.00495983f $X=17.44 $Y=0.255 $X2=0 $Y2=0
cc_2311 N_S[5]_c_2892_n N_Z_c_5220_n 0.00413022f $X=17.86 $Y=0.255 $X2=0 $Y2=0
cc_2312 N_S[5]_c_2885_n N_Z_c_5250_n 0.00513674f $X=16.37 $Y=1.41 $X2=0 $Y2=0
cc_2313 S[5] N_Z_c_5250_n 0.00545567f $X=16.245 $Y=1.105 $X2=0 $Y2=0
cc_2314 N_S[5]_c_2890_n N_Z_c_5231_n 0.00133607f $X=17.44 $Y=0.255 $X2=0 $Y2=0
cc_2315 N_S[5]_c_2892_n N_Z_c_5231_n 0.00199103f $X=17.86 $Y=0.255 $X2=0 $Y2=0
cc_2316 N_S[5]_c_2884_n N_VGND_c_7795_n 0.00330937f $X=16.31 $Y=0.845 $X2=0
+ $Y2=0
cc_2317 N_S[5]_c_2884_n VGND 0.0111218f $X=16.31 $Y=0.845 $X2=0 $Y2=0
cc_2318 N_S[5]_c_2888_n VGND 0.0119932f $X=17.365 $Y=0.18 $X2=0 $Y2=0
cc_2319 N_S[5]_c_2889_n VGND 0.00731624f $X=17.03 $Y=0.18 $X2=0 $Y2=0
cc_2320 N_S[5]_c_2891_n VGND 0.0111713f $X=17.785 $Y=0.18 $X2=0 $Y2=0
cc_2321 N_S[5]_c_2893_n VGND 0.00366655f $X=17.44 $Y=0.18 $X2=0 $Y2=0
cc_2322 N_S[5]_c_2884_n N_VGND_c_7833_n 0.00585385f $X=16.31 $Y=0.845 $X2=0
+ $Y2=0
cc_2323 N_S[5]_c_2889_n N_VGND_c_7833_n 0.0271255f $X=17.03 $Y=0.18 $X2=0 $Y2=0
cc_2324 N_S[5]_c_2887_n N_A_3421_69#_c_8709_n 0.00295202f $X=16.955 $Y=0.845
+ $X2=0 $Y2=0
cc_2325 N_S[5]_c_2890_n N_A_3421_69#_c_8705_n 0.0126455f $X=17.44 $Y=0.255 $X2=0
+ $Y2=0
cc_2326 N_S[5]_c_2891_n N_A_3421_69#_c_8705_n 0.00211351f $X=17.785 $Y=0.18
+ $X2=0 $Y2=0
cc_2327 N_S[5]_c_2892_n N_A_3421_69#_c_8705_n 0.0132844f $X=17.86 $Y=0.255 $X2=0
+ $Y2=0
cc_2328 N_S[5]_c_2887_n N_A_3421_69#_c_8706_n 0.00349455f $X=16.955 $Y=0.845
+ $X2=0 $Y2=0
cc_2329 N_S[5]_c_2888_n N_A_3421_69#_c_8706_n 0.00436105f $X=17.365 $Y=0.18
+ $X2=0 $Y2=0
cc_2330 N_S[5]_c_2892_n N_A_3421_69#_c_8708_n 0.00139422f $X=17.86 $Y=0.255
+ $X2=0 $Y2=0
cc_2331 N_S[13]_c_2954_n N_A_3277_937#_c_3099_n 0.00779314f $X=17.86 $Y=5.185
+ $X2=0 $Y2=0
cc_2332 N_S[13]_c_2947_n N_A_3277_937#_c_3094_n 0.00543241f $X=16.31 $Y=4.595
+ $X2=0 $Y2=0
cc_2333 N_S[13]_c_2958_n N_A_3277_937#_c_3094_n 0.00149275f $X=16.37 $Y=4.03
+ $X2=0 $Y2=0
cc_2334 N_S[13]_c_2948_n N_A_3277_937#_c_3094_n 0.00920672f $X=16.88 $Y=4.52
+ $X2=0 $Y2=0
cc_2335 N_S[13]_c_2952_n N_A_3277_937#_c_3094_n 0.00810157f $X=17.44 $Y=5.185
+ $X2=0 $Y2=0
cc_2336 S[13] N_A_3277_937#_c_3094_n 3.07062e-19 $X=16.245 $Y=4.165 $X2=0 $Y2=0
cc_2337 N_S[13]_c_2958_n N_A_3277_937#_c_3102_n 0.00861299f $X=16.37 $Y=4.03
+ $X2=0 $Y2=0
cc_2338 N_S[13]_c_2947_n N_A_3277_937#_c_3095_n 0.00354873f $X=16.31 $Y=4.595
+ $X2=0 $Y2=0
cc_2339 N_S[13]_c_2948_n N_A_3277_937#_c_3095_n 0.0135307f $X=16.88 $Y=4.52
+ $X2=0 $Y2=0
cc_2340 N_S[13]_c_2949_n N_A_3277_937#_c_3095_n 0.00267287f $X=16.955 $Y=5.185
+ $X2=0 $Y2=0
cc_2341 N_S[13]_c_2952_n N_A_3277_937#_c_3095_n 7.04048e-19 $X=17.44 $Y=5.185
+ $X2=0 $Y2=0
cc_2342 S[13] N_A_3277_937#_c_3095_n 0.0101733f $X=16.245 $Y=4.165 $X2=0 $Y2=0
cc_2343 N_S[13]_c_2947_n N_A_3277_937#_c_3096_n 0.0105766f $X=16.31 $Y=4.595
+ $X2=0 $Y2=0
cc_2344 N_S[13]_c_2949_n N_A_3277_937#_c_3096_n 0.0100374f $X=16.955 $Y=5.185
+ $X2=0 $Y2=0
cc_2345 S[13] N_A_3277_937#_c_3096_n 0.0061421f $X=16.245 $Y=4.165 $X2=0 $Y2=0
cc_2346 N_S[13]_c_2947_n N_A_3277_937#_c_3097_n 0.00441664f $X=16.31 $Y=4.595
+ $X2=0 $Y2=0
cc_2347 N_S[13]_c_2958_n N_A_3277_937#_c_3097_n 0.00386817f $X=16.37 $Y=4.03
+ $X2=0 $Y2=0
cc_2348 N_S[13]_c_2948_n N_A_3277_937#_c_3097_n 0.00785343f $X=16.88 $Y=4.52
+ $X2=0 $Y2=0
cc_2349 S[13] N_A_3277_937#_c_3097_n 0.0127184f $X=16.245 $Y=4.165 $X2=0 $Y2=0
cc_2350 N_S[13]_c_2954_n N_D[13]_M1100_g 0.0165585f $X=17.86 $Y=5.185 $X2=0
+ $Y2=0
cc_2351 N_S[13]_c_2947_n N_VPWR_c_4261_n 9.39395e-19 $X=16.31 $Y=4.595 $X2=0
+ $Y2=0
cc_2352 N_S[13]_c_2958_n N_VPWR_c_4261_n 0.00362951f $X=16.37 $Y=4.03 $X2=0
+ $Y2=0
cc_2353 S[13] N_VPWR_c_4261_n 0.00569857f $X=16.245 $Y=4.165 $X2=0 $Y2=0
cc_2354 N_S[13]_c_2958_n VPWR 0.00710985f $X=16.37 $Y=4.03 $X2=0 $Y2=0
cc_2355 N_S[13]_c_2958_n N_VPWR_c_4289_n 0.0035837f $X=16.37 $Y=4.03 $X2=0 $Y2=0
cc_2356 N_S[13]_c_2952_n N_Z_c_5207_n 0.00133607f $X=17.44 $Y=5.185 $X2=0 $Y2=0
cc_2357 N_S[13]_c_2954_n N_Z_c_5207_n 0.00199103f $X=17.86 $Y=5.185 $X2=0 $Y2=0
cc_2358 N_S[13]_c_2948_n N_Z_c_5221_n 4.25992e-19 $X=16.88 $Y=4.52 $X2=0 $Y2=0
cc_2359 N_S[13]_c_2952_n N_Z_c_5221_n 0.00495983f $X=17.44 $Y=5.185 $X2=0 $Y2=0
cc_2360 N_S[13]_c_2954_n N_Z_c_5221_n 0.00413022f $X=17.86 $Y=5.185 $X2=0 $Y2=0
cc_2361 N_S[13]_c_2947_n N_Z_c_5251_n 3.57797e-19 $X=16.31 $Y=4.595 $X2=0 $Y2=0
cc_2362 N_S[13]_c_2958_n N_Z_c_5251_n 0.00477894f $X=16.37 $Y=4.03 $X2=0 $Y2=0
cc_2363 S[13] N_Z_c_5251_n 0.00545567f $X=16.245 $Y=4.165 $X2=0 $Y2=0
cc_2364 N_S[13]_c_2947_n N_VGND_c_7796_n 0.00330937f $X=16.31 $Y=4.595 $X2=0
+ $Y2=0
cc_2365 N_S[13]_c_2947_n VGND 0.0111218f $X=16.31 $Y=4.595 $X2=0 $Y2=0
cc_2366 N_S[13]_c_2950_n VGND 0.0119932f $X=17.365 $Y=5.26 $X2=0 $Y2=0
cc_2367 N_S[13]_c_2951_n VGND 0.00731624f $X=17.03 $Y=5.26 $X2=0 $Y2=0
cc_2368 N_S[13]_c_2953_n VGND 0.0111713f $X=17.785 $Y=5.26 $X2=0 $Y2=0
cc_2369 N_S[13]_c_2955_n VGND 0.00366655f $X=17.44 $Y=5.26 $X2=0 $Y2=0
cc_2370 N_S[13]_c_2947_n N_VGND_c_7834_n 0.00585385f $X=16.31 $Y=4.595 $X2=0
+ $Y2=0
cc_2371 N_S[13]_c_2951_n N_VGND_c_7834_n 0.0271255f $X=17.03 $Y=5.26 $X2=0 $Y2=0
cc_2372 N_S[13]_c_2949_n N_A_3421_915#_c_8757_n 0.00295202f $X=16.955 $Y=5.185
+ $X2=0 $Y2=0
cc_2373 N_S[13]_c_2952_n N_A_3421_915#_c_8753_n 0.0126455f $X=17.44 $Y=5.185
+ $X2=0 $Y2=0
cc_2374 N_S[13]_c_2953_n N_A_3421_915#_c_8753_n 0.00211351f $X=17.785 $Y=5.26
+ $X2=0 $Y2=0
cc_2375 N_S[13]_c_2954_n N_A_3421_915#_c_8753_n 0.0132844f $X=17.86 $Y=5.185
+ $X2=0 $Y2=0
cc_2376 N_S[13]_c_2949_n N_A_3421_915#_c_8754_n 0.00349455f $X=16.955 $Y=5.185
+ $X2=0 $Y2=0
cc_2377 N_S[13]_c_2950_n N_A_3421_915#_c_8754_n 0.00436105f $X=17.365 $Y=5.26
+ $X2=0 $Y2=0
cc_2378 N_S[13]_c_2954_n N_A_3421_915#_c_8755_n 0.00139422f $X=17.86 $Y=5.185
+ $X2=0 $Y2=0
cc_2379 N_A_3277_47#_M1055_g N_A_3277_937#_M1134_g 0.0130744f $X=17.36 $Y=2.075
+ $X2=0 $Y2=0
cc_2380 N_A_3277_47#_M1082_g N_A_3277_937#_M1158_g 0.0130744f $X=17.83 $Y=2.075
+ $X2=0 $Y2=0
cc_2381 N_A_3277_47#_c_3018_n N_D[5]_M1051_g 0.00671996f $X=17.74 $Y=1.4 $X2=0
+ $Y2=0
cc_2382 N_A_3277_47#_M1082_g N_D[5]_M1051_g 0.025073f $X=17.83 $Y=2.075 $X2=0
+ $Y2=0
cc_2383 N_A_3277_47#_c_3021_n N_VPWR_c_4260_n 0.0321301f $X=16.605 $Y=2.31 $X2=0
+ $Y2=0
cc_2384 N_A_3277_47#_c_3016_n N_VPWR_c_4260_n 0.00732952f $X=16.89 $Y=1.42 $X2=0
+ $Y2=0
cc_2385 N_A_3277_47#_M1082_g N_VPWR_c_4262_n 0.00107878f $X=17.83 $Y=2.075 $X2=0
+ $Y2=0
cc_2386 N_A_3277_47#_M1065_d VPWR 0.00179197f $X=16.46 $Y=1.485 $X2=0 $Y2=0
cc_2387 N_A_3277_47#_M1055_g VPWR 0.0054792f $X=17.36 $Y=2.075 $X2=0 $Y2=0
cc_2388 N_A_3277_47#_M1082_g VPWR 0.00435072f $X=17.83 $Y=2.075 $X2=0 $Y2=0
cc_2389 N_A_3277_47#_c_3021_n VPWR 0.00594162f $X=16.605 $Y=2.31 $X2=0 $Y2=0
cc_2390 N_A_3277_47#_M1055_g N_VPWR_c_4289_n 8.06528e-19 $X=17.36 $Y=2.075 $X2=0
+ $Y2=0
cc_2391 N_A_3277_47#_c_3021_n N_VPWR_c_4289_n 0.0210596f $X=16.605 $Y=2.31 $X2=0
+ $Y2=0
cc_2392 N_A_3277_47#_c_3018_n N_Z_c_5220_n 0.00348752f $X=17.74 $Y=1.4 $X2=0
+ $Y2=0
cc_2393 N_A_3277_47#_c_3014_n N_Z_c_5220_n 0.0033343f $X=16.89 $Y=1.205 $X2=0
+ $Y2=0
cc_2394 N_A_3277_47#_M1055_g N_Z_c_5250_n 0.00708998f $X=17.36 $Y=2.075 $X2=0
+ $Y2=0
cc_2395 N_A_3277_47#_c_3013_n N_Z_c_5250_n 9.57301e-19 $X=17.45 $Y=1.4 $X2=0
+ $Y2=0
cc_2396 N_A_3277_47#_c_3021_n N_Z_c_5250_n 0.0308332f $X=16.605 $Y=2.31 $X2=0
+ $Y2=0
cc_2397 N_A_3277_47#_c_3016_n N_Z_c_5250_n 0.0132841f $X=16.89 $Y=1.42 $X2=0
+ $Y2=0
cc_2398 N_A_3277_47#_M1082_g N_Z_c_5252_n 0.00404618f $X=17.83 $Y=2.075 $X2=0
+ $Y2=0
cc_2399 N_A_3277_47#_M1082_g N_Z_c_5637_n 0.00513826f $X=17.83 $Y=2.075 $X2=0
+ $Y2=0
cc_2400 N_A_3277_47#_M1055_g N_Z_c_5638_n 0.00619657f $X=17.36 $Y=2.075 $X2=0
+ $Y2=0
cc_2401 N_A_3277_47#_c_3018_n N_Z_c_5638_n 8.37785e-19 $X=17.74 $Y=1.4 $X2=0
+ $Y2=0
cc_2402 N_A_3277_47#_M1082_g N_Z_c_5638_n 0.00978858f $X=17.83 $Y=2.075 $X2=0
+ $Y2=0
cc_2403 N_A_3277_47#_M1055_g N_Z_c_5231_n 0.00476154f $X=17.36 $Y=2.075 $X2=0
+ $Y2=0
cc_2404 N_A_3277_47#_c_3018_n N_Z_c_5231_n 0.0140957f $X=17.74 $Y=1.4 $X2=0
+ $Y2=0
cc_2405 N_A_3277_47#_c_3013_n N_Z_c_5231_n 7.26438e-19 $X=17.45 $Y=1.4 $X2=0
+ $Y2=0
cc_2406 N_A_3277_47#_M1082_g N_Z_c_5231_n 0.00268051f $X=17.83 $Y=2.075 $X2=0
+ $Y2=0
cc_2407 N_A_3277_47#_c_3014_n N_Z_c_5231_n 0.00967956f $X=16.89 $Y=1.205 $X2=0
+ $Y2=0
cc_2408 N_A_3277_47#_c_3016_n N_Z_c_5231_n 0.0117695f $X=16.89 $Y=1.42 $X2=0
+ $Y2=0
cc_2409 N_A_3277_47#_M1082_g N_Z_c_5647_n 2.61869e-19 $X=17.83 $Y=2.075 $X2=0
+ $Y2=0
cc_2410 N_A_3277_47#_M1055_g N_Z_c_5267_n 0.00462462f $X=17.36 $Y=2.075 $X2=0
+ $Y2=0
cc_2411 N_A_3277_47#_M1082_g N_Z_c_5267_n 0.00455034f $X=17.83 $Y=2.075 $X2=0
+ $Y2=0
cc_2412 N_A_3277_47#_M1082_g N_A_3400_333#_c_7169_n 0.00176121f $X=17.83
+ $Y=2.075 $X2=0 $Y2=0
cc_2413 N_A_3277_47#_M1055_g N_A_3400_333#_c_7170_n 0.00334959f $X=17.36
+ $Y=2.075 $X2=0 $Y2=0
cc_2414 N_A_3277_47#_M1082_g N_A_3400_333#_c_7170_n 0.00463461f $X=17.83
+ $Y=2.075 $X2=0 $Y2=0
cc_2415 N_A_3277_47#_c_3021_n N_A_3400_333#_c_7165_n 0.00738363f $X=16.605
+ $Y=2.31 $X2=0 $Y2=0
cc_2416 N_A_3277_47#_M1082_g N_A_3400_333#_c_7173_n 7.75952e-19 $X=17.83
+ $Y=2.075 $X2=0 $Y2=0
cc_2417 N_A_3277_47#_M1055_g N_A_3400_333#_c_7174_n 0.00692695f $X=17.36
+ $Y=2.075 $X2=0 $Y2=0
cc_2418 N_A_3277_47#_M1082_g N_A_3400_333#_c_7175_n 0.00415998f $X=17.83
+ $Y=2.075 $X2=0 $Y2=0
cc_2419 N_A_3277_47#_M1055_g N_A_3400_333#_c_7167_n 0.00550198f $X=17.36
+ $Y=2.075 $X2=0 $Y2=0
cc_2420 N_A_3277_47#_c_3013_n N_A_3400_333#_c_7167_n 0.00133381f $X=17.45 $Y=1.4
+ $X2=0 $Y2=0
cc_2421 N_A_3277_47#_c_3021_n N_A_3400_333#_c_7167_n 0.0413447f $X=16.605
+ $Y=2.31 $X2=0 $Y2=0
cc_2422 N_A_3277_47#_c_3016_n N_A_3400_333#_c_7167_n 0.0132748f $X=16.89 $Y=1.42
+ $X2=0 $Y2=0
cc_2423 N_A_3277_47#_M1082_g N_A_3400_333#_c_7180_n 0.00508488f $X=17.83
+ $Y=2.075 $X2=0 $Y2=0
cc_2424 N_A_3277_47#_M1098_d VGND 0.00250855f $X=16.385 $Y=0.235 $X2=0 $Y2=0
cc_2425 N_A_3277_47#_c_3015_n VGND 0.0186564f $X=16.52 $Y=0.495 $X2=0 $Y2=0
cc_2426 N_A_3277_47#_c_3015_n N_VGND_c_7833_n 0.0173492f $X=16.52 $Y=0.495 $X2=0
+ $Y2=0
cc_2427 N_A_3277_47#_c_3013_n N_A_3421_69#_c_8709_n 0.00308807f $X=17.45 $Y=1.4
+ $X2=0 $Y2=0
cc_2428 N_A_3277_47#_c_3014_n N_A_3421_69#_c_8709_n 0.00101918f $X=16.89
+ $Y=1.205 $X2=0 $Y2=0
cc_2429 N_A_3277_47#_c_3015_n N_A_3421_69#_c_8709_n 0.0185512f $X=16.52 $Y=0.495
+ $X2=0 $Y2=0
cc_2430 N_A_3277_47#_c_3016_n N_A_3421_69#_c_8709_n 0.00285813f $X=16.89 $Y=1.42
+ $X2=0 $Y2=0
cc_2431 N_A_3277_47#_c_3015_n N_A_3421_69#_c_8706_n 0.00358194f $X=16.52
+ $Y=0.495 $X2=0 $Y2=0
cc_2432 N_A_3277_937#_c_3099_n N_D[13]_M1058_g 0.00671996f $X=17.74 $Y=4.04
+ $X2=0 $Y2=0
cc_2433 N_A_3277_937#_M1158_g N_D[13]_M1058_g 0.0250718f $X=17.83 $Y=3.365 $X2=0
+ $Y2=0
cc_2434 N_A_3277_937#_c_3102_n N_VPWR_c_4261_n 0.0321301f $X=16.605 $Y=3.13
+ $X2=0 $Y2=0
cc_2435 N_A_3277_937#_c_3097_n N_VPWR_c_4261_n 0.00732952f $X=16.89 $Y=4.02
+ $X2=0 $Y2=0
cc_2436 N_A_3277_937#_M1158_g N_VPWR_c_4263_n 0.0013032f $X=17.83 $Y=3.365 $X2=0
+ $Y2=0
cc_2437 N_A_3277_937#_M1070_d VPWR 0.00179197f $X=16.46 $Y=2.955 $X2=0 $Y2=0
cc_2438 N_A_3277_937#_M1134_g VPWR 0.00546988f $X=17.36 $Y=3.365 $X2=0 $Y2=0
cc_2439 N_A_3277_937#_M1158_g VPWR 0.00434142f $X=17.83 $Y=3.365 $X2=0 $Y2=0
cc_2440 N_A_3277_937#_c_3102_n VPWR 0.00594162f $X=16.605 $Y=3.13 $X2=0 $Y2=0
cc_2441 N_A_3277_937#_M1134_g N_VPWR_c_4289_n 7.91347e-19 $X=17.36 $Y=3.365
+ $X2=0 $Y2=0
cc_2442 N_A_3277_937#_c_3102_n N_VPWR_c_4289_n 0.0210596f $X=16.605 $Y=3.13
+ $X2=0 $Y2=0
cc_2443 N_A_3277_937#_M1134_g N_Z_c_5207_n 0.00476154f $X=17.36 $Y=3.365 $X2=0
+ $Y2=0
cc_2444 N_A_3277_937#_c_3099_n N_Z_c_5207_n 0.0140957f $X=17.74 $Y=4.04 $X2=0
+ $Y2=0
cc_2445 N_A_3277_937#_c_3094_n N_Z_c_5207_n 7.26438e-19 $X=17.45 $Y=4.04 $X2=0
+ $Y2=0
cc_2446 N_A_3277_937#_M1158_g N_Z_c_5207_n 0.00268051f $X=17.83 $Y=3.365 $X2=0
+ $Y2=0
cc_2447 N_A_3277_937#_c_3095_n N_Z_c_5207_n 0.00967956f $X=16.89 $Y=4.685 $X2=0
+ $Y2=0
cc_2448 N_A_3277_937#_c_3097_n N_Z_c_5207_n 0.0117695f $X=16.89 $Y=4.02 $X2=0
+ $Y2=0
cc_2449 N_A_3277_937#_c_3099_n N_Z_c_5221_n 0.00348752f $X=17.74 $Y=4.04 $X2=0
+ $Y2=0
cc_2450 N_A_3277_937#_c_3095_n N_Z_c_5221_n 0.0033343f $X=16.89 $Y=4.685 $X2=0
+ $Y2=0
cc_2451 N_A_3277_937#_M1134_g N_Z_c_5251_n 0.00708682f $X=17.36 $Y=3.365 $X2=0
+ $Y2=0
cc_2452 N_A_3277_937#_c_3094_n N_Z_c_5251_n 9.57301e-19 $X=17.45 $Y=4.04 $X2=0
+ $Y2=0
cc_2453 N_A_3277_937#_c_3102_n N_Z_c_5251_n 0.0308332f $X=16.605 $Y=3.13 $X2=0
+ $Y2=0
cc_2454 N_A_3277_937#_c_3097_n N_Z_c_5251_n 0.0132841f $X=16.89 $Y=4.02 $X2=0
+ $Y2=0
cc_2455 N_A_3277_937#_M1158_g N_Z_c_5253_n 0.0040431f $X=17.83 $Y=3.365 $X2=0
+ $Y2=0
cc_2456 N_A_3277_937#_M1158_g N_Z_c_5663_n 0.00513826f $X=17.83 $Y=3.365 $X2=0
+ $Y2=0
cc_2457 N_A_3277_937#_M1158_g N_Z_c_5638_n 2.61869e-19 $X=17.83 $Y=3.365 $X2=0
+ $Y2=0
cc_2458 N_A_3277_937#_M1134_g N_Z_c_5647_n 0.00619657f $X=17.36 $Y=3.365 $X2=0
+ $Y2=0
cc_2459 N_A_3277_937#_c_3099_n N_Z_c_5647_n 8.37785e-19 $X=17.74 $Y=4.04 $X2=0
+ $Y2=0
cc_2460 N_A_3277_937#_M1158_g N_Z_c_5647_n 0.00978858f $X=17.83 $Y=3.365 $X2=0
+ $Y2=0
cc_2461 N_A_3277_937#_M1134_g N_Z_c_5267_n 0.00462236f $X=17.36 $Y=3.365 $X2=0
+ $Y2=0
cc_2462 N_A_3277_937#_M1158_g N_Z_c_5267_n 0.00455034f $X=17.83 $Y=3.365 $X2=0
+ $Y2=0
cc_2463 N_A_3277_937#_M1158_g N_A_3400_591#_c_7265_n 0.00176121f $X=17.83
+ $Y=3.365 $X2=0 $Y2=0
cc_2464 N_A_3277_937#_M1134_g N_A_3400_591#_c_7262_n 0.0124482f $X=17.36
+ $Y=3.365 $X2=0 $Y2=0
cc_2465 N_A_3277_937#_c_3094_n N_A_3400_591#_c_7262_n 0.00133381f $X=17.45
+ $Y=4.04 $X2=0 $Y2=0
cc_2466 N_A_3277_937#_c_3102_n N_A_3400_591#_c_7262_n 0.0413753f $X=16.605
+ $Y=3.13 $X2=0 $Y2=0
cc_2467 N_A_3277_937#_c_3097_n N_A_3400_591#_c_7262_n 0.0132748f $X=16.89
+ $Y=4.02 $X2=0 $Y2=0
cc_2468 N_A_3277_937#_M1158_g N_A_3400_591#_c_7270_n 0.00400484f $X=17.83
+ $Y=3.365 $X2=0 $Y2=0
cc_2469 N_A_3277_937#_M1134_g N_A_3400_591#_c_7271_n 0.00334069f $X=17.36
+ $Y=3.365 $X2=0 $Y2=0
cc_2470 N_A_3277_937#_M1158_g N_A_3400_591#_c_7271_n 0.00470988f $X=17.83
+ $Y=3.365 $X2=0 $Y2=0
cc_2471 N_A_3277_937#_c_3102_n N_A_3400_591#_c_7263_n 0.00738293f $X=16.605
+ $Y=3.13 $X2=0 $Y2=0
cc_2472 N_A_3277_937#_M1158_g N_A_3400_591#_c_7274_n 7.75952e-19 $X=17.83
+ $Y=3.365 $X2=0 $Y2=0
cc_2473 N_A_3277_937#_M1158_g N_A_3400_591#_c_7275_n 0.00508821f $X=17.83
+ $Y=3.365 $X2=0 $Y2=0
cc_2474 N_A_3277_937#_M1096_d VGND 0.00250855f $X=16.385 $Y=4.685 $X2=0 $Y2=0
cc_2475 N_A_3277_937#_c_3096_n VGND 0.0186503f $X=16.52 $Y=4.945 $X2=0 $Y2=0
cc_2476 N_A_3277_937#_c_3096_n N_VGND_c_7834_n 0.0173402f $X=16.52 $Y=4.945
+ $X2=0 $Y2=0
cc_2477 N_A_3277_937#_c_3094_n N_A_3421_915#_c_8757_n 0.00308807f $X=17.45
+ $Y=4.04 $X2=0 $Y2=0
cc_2478 N_A_3277_937#_c_3095_n N_A_3421_915#_c_8757_n 0.00101918f $X=16.89
+ $Y=4.685 $X2=0 $Y2=0
cc_2479 N_A_3277_937#_c_3096_n N_A_3421_915#_c_8757_n 0.0185512f $X=16.52
+ $Y=4.945 $X2=0 $Y2=0
cc_2480 N_A_3277_937#_c_3097_n N_A_3421_915#_c_8757_n 0.00285813f $X=16.89
+ $Y=4.02 $X2=0 $Y2=0
cc_2481 N_A_3277_937#_c_3096_n N_A_3421_915#_c_8754_n 0.00358194f $X=16.52
+ $Y=4.945 $X2=0 $Y2=0
cc_2482 N_D[5]_M1051_g N_D[13]_M1058_g 0.0129371f $X=18.355 $Y=1.985 $X2=0 $Y2=0
cc_2483 N_D[5]_M1079_g N_D[13]_M1087_g 0.0130744f $X=18.825 $Y=1.985 $X2=0 $Y2=0
cc_2484 D[5] N_D[6]_c_3293_n 0.0231965f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_2485 N_D[5]_c_3180_n N_D[6]_c_3293_n 7.85936e-19 $X=18.91 $Y=1.16 $X2=0 $Y2=0
cc_2486 D[5] N_D[6]_c_3294_n 7.85936e-19 $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_2487 N_D[5]_c_3180_n N_D[6]_c_3294_n 0.00603597f $X=18.91 $Y=1.16 $X2=0 $Y2=0
cc_2488 N_D[5]_M1051_g N_VPWR_c_4262_n 0.00848021f $X=18.355 $Y=1.985 $X2=0
+ $Y2=0
cc_2489 N_D[5]_M1079_g N_VPWR_c_4262_n 0.00338721f $X=18.825 $Y=1.985 $X2=0
+ $Y2=0
cc_2490 N_D[5]_M1051_g N_VPWR_c_4548_n 0.00295119f $X=18.355 $Y=1.985 $X2=0
+ $Y2=0
cc_2491 N_D[5]_M1079_g N_VPWR_c_4548_n 0.00311479f $X=18.825 $Y=1.985 $X2=0
+ $Y2=0
cc_2492 N_D[5]_M1051_g VPWR 0.00350923f $X=18.355 $Y=1.985 $X2=0 $Y2=0
cc_2493 N_D[5]_M1079_g VPWR 0.00568683f $X=18.825 $Y=1.985 $X2=0 $Y2=0
cc_2494 N_D[5]_M1051_g N_VPWR_c_4290_n 0.00342413f $X=18.355 $Y=1.985 $X2=0
+ $Y2=0
cc_2495 N_D[5]_M1079_g N_VPWR_c_4291_n 0.0033767f $X=18.825 $Y=1.985 $X2=0 $Y2=0
cc_2496 N_D[5]_M1051_g N_Z_c_5252_n 0.0033316f $X=18.355 $Y=1.985 $X2=0 $Y2=0
cc_2497 N_D[5]_M1079_g N_Z_c_5252_n 0.00312829f $X=18.825 $Y=1.985 $X2=0 $Y2=0
cc_2498 D[5] N_Z_c_5252_n 0.00125914f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_2499 N_D[5]_M1051_g N_Z_c_5231_n 0.00112534f $X=18.355 $Y=1.985 $X2=0 $Y2=0
cc_2500 N_D[5]_M1090_g N_Z_c_5231_n 8.13311e-19 $X=18.38 $Y=0.56 $X2=0 $Y2=0
cc_2501 D[5] N_Z_c_5231_n 0.00742792f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_2502 N_D[5]_c_3180_n N_Z_c_5231_n 0.00583073f $X=18.91 $Y=1.16 $X2=0 $Y2=0
cc_2503 N_D[5]_M1051_g N_A_3400_333#_c_7181_n 0.0127833f $X=18.355 $Y=1.985
+ $X2=0 $Y2=0
cc_2504 N_D[5]_M1079_g N_A_3400_333#_c_7181_n 0.0101085f $X=18.825 $Y=1.985
+ $X2=0 $Y2=0
cc_2505 D[5] N_A_3400_333#_c_7181_n 0.0323774f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_2506 N_D[5]_c_3180_n N_A_3400_333#_c_7181_n 7.13708e-19 $X=18.91 $Y=1.16
+ $X2=0 $Y2=0
cc_2507 D[5] N_A_3400_333#_c_7164_n 0.0226682f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_2508 N_D[5]_c_3180_n N_A_3400_333#_c_7164_n 9.6385e-19 $X=18.91 $Y=1.16 $X2=0
+ $Y2=0
cc_2509 N_D[5]_M1051_g N_A_3400_333#_c_7187_n 0.00246916f $X=18.355 $Y=1.985
+ $X2=0 $Y2=0
cc_2510 N_D[5]_M1079_g N_A_3400_333#_c_7187_n 0.00244285f $X=18.825 $Y=1.985
+ $X2=0 $Y2=0
cc_2511 N_D[5]_M1079_g N_A_3400_333#_c_7166_n 0.00290175f $X=18.825 $Y=1.985
+ $X2=0 $Y2=0
cc_2512 N_D[5]_M1051_g N_A_3400_333#_c_7180_n 0.00595395f $X=18.355 $Y=1.985
+ $X2=0 $Y2=0
cc_2513 N_D[5]_M1090_g N_VGND_c_7797_n 0.00300333f $X=18.38 $Y=0.56 $X2=0 $Y2=0
cc_2514 N_D[5]_M1110_g N_VGND_c_7797_n 0.0030929f $X=18.8 $Y=0.56 $X2=0 $Y2=0
cc_2515 N_D[5]_M1110_g N_VGND_c_7799_n 0.00430643f $X=18.8 $Y=0.56 $X2=0 $Y2=0
cc_2516 N_D[5]_M1090_g VGND 0.00600262f $X=18.38 $Y=0.56 $X2=0 $Y2=0
cc_2517 N_D[5]_M1110_g VGND 0.00733187f $X=18.8 $Y=0.56 $X2=0 $Y2=0
cc_2518 N_D[5]_M1090_g N_VGND_c_7833_n 0.00436487f $X=18.38 $Y=0.56 $X2=0 $Y2=0
cc_2519 N_D[5]_M1090_g N_A_3421_69#_c_8707_n 0.0114493f $X=18.38 $Y=0.56 $X2=0
+ $Y2=0
cc_2520 N_D[5]_M1110_g N_A_3421_69#_c_8707_n 0.00931728f $X=18.8 $Y=0.56 $X2=0
+ $Y2=0
cc_2521 D[5] N_A_3421_69#_c_8707_n 0.0518587f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_2522 N_D[5]_c_3180_n N_A_3421_69#_c_8707_n 0.00665175f $X=18.91 $Y=1.16 $X2=0
+ $Y2=0
cc_2523 N_D[5]_M1090_g N_A_3421_69#_c_8708_n 0.00114614f $X=18.38 $Y=0.56 $X2=0
+ $Y2=0
cc_2524 N_D[5]_c_3180_n N_A_3421_69#_c_8708_n 0.00120541f $X=18.91 $Y=1.16 $X2=0
+ $Y2=0
cc_2525 N_D[5]_M1090_g N_A_3421_69#_c_8727_n 5.29024e-19 $X=18.38 $Y=0.56 $X2=0
+ $Y2=0
cc_2526 N_D[5]_M1110_g N_A_3421_69#_c_8727_n 0.00633603f $X=18.8 $Y=0.56 $X2=0
+ $Y2=0
cc_2527 D[13] N_D[14]_c_3351_n 0.0231965f $X=19.005 $Y=4.165 $X2=0 $Y2=0
cc_2528 N_D[13]_c_3237_n N_D[14]_c_3351_n 7.85936e-19 $X=18.91 $Y=4.28 $X2=0
+ $Y2=0
cc_2529 D[13] N_D[14]_c_3352_n 7.85936e-19 $X=19.005 $Y=4.165 $X2=0 $Y2=0
cc_2530 N_D[13]_c_3237_n N_D[14]_c_3352_n 0.00603597f $X=18.91 $Y=4.28 $X2=0
+ $Y2=0
cc_2531 N_D[13]_M1058_g N_VPWR_c_4263_n 0.00847423f $X=18.355 $Y=3.455 $X2=0
+ $Y2=0
cc_2532 N_D[13]_M1087_g N_VPWR_c_4263_n 0.00338721f $X=18.825 $Y=3.455 $X2=0
+ $Y2=0
cc_2533 N_D[13]_M1058_g N_VPWR_c_4556_n 0.00295119f $X=18.355 $Y=3.455 $X2=0
+ $Y2=0
cc_2534 N_D[13]_M1087_g N_VPWR_c_4556_n 0.00311479f $X=18.825 $Y=3.455 $X2=0
+ $Y2=0
cc_2535 N_D[13]_M1058_g VPWR 0.00350923f $X=18.355 $Y=3.455 $X2=0 $Y2=0
cc_2536 N_D[13]_M1087_g VPWR 0.00568683f $X=18.825 $Y=3.455 $X2=0 $Y2=0
cc_2537 N_D[13]_M1058_g N_VPWR_c_4290_n 0.00342413f $X=18.355 $Y=3.455 $X2=0
+ $Y2=0
cc_2538 N_D[13]_M1087_g N_VPWR_c_4291_n 0.0033767f $X=18.825 $Y=3.455 $X2=0
+ $Y2=0
cc_2539 N_D[13]_M1058_g N_Z_c_5207_n 0.00112534f $X=18.355 $Y=3.455 $X2=0 $Y2=0
cc_2540 N_D[13]_M1100_g N_Z_c_5207_n 8.13311e-19 $X=18.38 $Y=4.88 $X2=0 $Y2=0
cc_2541 D[13] N_Z_c_5207_n 0.00742792f $X=19.005 $Y=4.165 $X2=0 $Y2=0
cc_2542 N_D[13]_c_3237_n N_Z_c_5207_n 0.00583073f $X=18.91 $Y=4.28 $X2=0 $Y2=0
cc_2543 N_D[13]_M1058_g N_Z_c_5253_n 0.0033316f $X=18.355 $Y=3.455 $X2=0 $Y2=0
cc_2544 N_D[13]_M1087_g N_Z_c_5253_n 0.00312829f $X=18.825 $Y=3.455 $X2=0 $Y2=0
cc_2545 D[13] N_Z_c_5253_n 0.00125914f $X=19.005 $Y=4.165 $X2=0 $Y2=0
cc_2546 N_D[13]_M1058_g N_A_3400_591#_c_7260_n 0.0127833f $X=18.355 $Y=3.455
+ $X2=0 $Y2=0
cc_2547 N_D[13]_M1087_g N_A_3400_591#_c_7260_n 0.0101085f $X=18.825 $Y=3.455
+ $X2=0 $Y2=0
cc_2548 D[13] N_A_3400_591#_c_7260_n 0.0550456f $X=19.005 $Y=4.165 $X2=0 $Y2=0
cc_2549 N_D[13]_c_3237_n N_A_3400_591#_c_7260_n 0.00167756f $X=18.91 $Y=4.28
+ $X2=0 $Y2=0
cc_2550 N_D[13]_M1058_g N_A_3400_591#_c_7280_n 0.00246473f $X=18.355 $Y=3.455
+ $X2=0 $Y2=0
cc_2551 N_D[13]_M1087_g N_A_3400_591#_c_7280_n 0.00244285f $X=18.825 $Y=3.455
+ $X2=0 $Y2=0
cc_2552 N_D[13]_M1058_g N_A_3400_591#_c_7275_n 0.00531997f $X=18.355 $Y=3.455
+ $X2=0 $Y2=0
cc_2553 N_D[13]_M1087_g N_A_3400_591#_c_7264_n 0.00290175f $X=18.825 $Y=3.455
+ $X2=0 $Y2=0
cc_2554 N_D[13]_M1100_g N_VGND_c_7798_n 0.00300333f $X=18.38 $Y=4.88 $X2=0 $Y2=0
cc_2555 N_D[13]_M1121_g N_VGND_c_7798_n 0.0030929f $X=18.8 $Y=4.88 $X2=0 $Y2=0
cc_2556 N_D[13]_M1121_g N_VGND_c_7800_n 0.00430643f $X=18.8 $Y=4.88 $X2=0 $Y2=0
cc_2557 N_D[13]_M1100_g VGND 0.00600262f $X=18.38 $Y=4.88 $X2=0 $Y2=0
cc_2558 N_D[13]_M1121_g VGND 0.00733187f $X=18.8 $Y=4.88 $X2=0 $Y2=0
cc_2559 N_D[13]_M1100_g N_VGND_c_7834_n 0.00436487f $X=18.38 $Y=4.88 $X2=0 $Y2=0
cc_2560 N_D[13]_M1100_g N_A_3421_915#_c_8755_n 0.00114614f $X=18.38 $Y=4.88
+ $X2=0 $Y2=0
cc_2561 N_D[13]_c_3237_n N_A_3421_915#_c_8755_n 0.00120541f $X=18.91 $Y=4.28
+ $X2=0 $Y2=0
cc_2562 N_D[13]_M1100_g N_A_3421_915#_c_8771_n 0.0114493f $X=18.38 $Y=4.88 $X2=0
+ $Y2=0
cc_2563 N_D[13]_M1121_g N_A_3421_915#_c_8771_n 0.0084485f $X=18.8 $Y=4.88 $X2=0
+ $Y2=0
cc_2564 D[13] N_A_3421_915#_c_8771_n 0.0274027f $X=19.005 $Y=4.165 $X2=0 $Y2=0
cc_2565 N_D[13]_c_3237_n N_A_3421_915#_c_8771_n 0.0020061f $X=18.91 $Y=4.28
+ $X2=0 $Y2=0
cc_2566 N_D[13]_M1100_g N_A_3421_915#_c_8756_n 5.29024e-19 $X=18.38 $Y=4.88
+ $X2=0 $Y2=0
cc_2567 N_D[13]_M1121_g N_A_3421_915#_c_8756_n 0.00720482f $X=18.8 $Y=4.88 $X2=0
+ $Y2=0
cc_2568 D[13] N_A_3421_915#_c_8756_n 0.024456f $X=19.005 $Y=4.165 $X2=0 $Y2=0
cc_2569 N_D[13]_c_3237_n N_A_3421_915#_c_8756_n 0.00464565f $X=18.91 $Y=4.28
+ $X2=0 $Y2=0
cc_2570 N_D[6]_M1062_g N_D[14]_M1069_g 0.0130744f $X=19.815 $Y=1.985 $X2=0 $Y2=0
cc_2571 N_D[6]_M1143_g N_D[14]_M1152_g 0.0129371f $X=20.285 $Y=1.985 $X2=0 $Y2=0
cc_2572 N_D[6]_M1143_g N_A_4142_265#_M1066_g 0.025073f $X=20.285 $Y=1.985 $X2=0
+ $Y2=0
cc_2573 N_D[6]_M1143_g N_A_4142_265#_c_3412_n 0.00671996f $X=20.285 $Y=1.985
+ $X2=0 $Y2=0
cc_2574 N_D[6]_M1155_g N_S[6]_c_3573_n 0.0165585f $X=20.26 $Y=0.56 $X2=0 $Y2=0
cc_2575 N_D[6]_M1062_g N_VPWR_c_4264_n 0.00338721f $X=19.815 $Y=1.985 $X2=0
+ $Y2=0
cc_2576 N_D[6]_M1143_g N_VPWR_c_4264_n 0.00848021f $X=20.285 $Y=1.985 $X2=0
+ $Y2=0
cc_2577 N_D[6]_M1062_g N_VPWR_c_4564_n 0.00311479f $X=19.815 $Y=1.985 $X2=0
+ $Y2=0
cc_2578 N_D[6]_M1143_g N_VPWR_c_4564_n 0.00295119f $X=20.285 $Y=1.985 $X2=0
+ $Y2=0
cc_2579 N_D[6]_M1062_g VPWR 0.00568683f $X=19.815 $Y=1.985 $X2=0 $Y2=0
cc_2580 N_D[6]_M1143_g VPWR 0.00350923f $X=20.285 $Y=1.985 $X2=0 $Y2=0
cc_2581 N_D[6]_M1062_g N_VPWR_c_4291_n 0.0033767f $X=19.815 $Y=1.985 $X2=0 $Y2=0
cc_2582 N_D[6]_M1143_g N_VPWR_c_4292_n 0.00342413f $X=20.285 $Y=1.985 $X2=0
+ $Y2=0
cc_2583 N_D[6]_M1062_g N_Z_c_5252_n 0.00312829f $X=19.815 $Y=1.985 $X2=0 $Y2=0
cc_2584 N_D[6]_M1143_g N_Z_c_5252_n 0.0033316f $X=20.285 $Y=1.985 $X2=0 $Y2=0
cc_2585 N_D[6]_c_3293_n N_Z_c_5252_n 0.00125914f $X=20.07 $Y=1.16 $X2=0 $Y2=0
cc_2586 N_D[6]_M1155_g N_Z_c_5232_n 8.13311e-19 $X=20.26 $Y=0.56 $X2=0 $Y2=0
cc_2587 N_D[6]_M1143_g N_Z_c_5232_n 0.00112534f $X=20.285 $Y=1.985 $X2=0 $Y2=0
cc_2588 N_D[6]_c_3293_n N_Z_c_5232_n 0.00742792f $X=20.07 $Y=1.16 $X2=0 $Y2=0
cc_2589 N_D[6]_c_3294_n N_Z_c_5232_n 0.00583073f $X=20.285 $Y=1.16 $X2=0 $Y2=0
cc_2590 N_D[6]_c_3293_n N_A_3891_297#_c_7351_n 0.0226682f $X=20.07 $Y=1.16 $X2=0
+ $Y2=0
cc_2591 N_D[6]_c_3294_n N_A_3891_297#_c_7351_n 9.6385e-19 $X=20.285 $Y=1.16
+ $X2=0 $Y2=0
cc_2592 N_D[6]_M1062_g N_A_3891_297#_c_7358_n 0.0101085f $X=19.815 $Y=1.985
+ $X2=0 $Y2=0
cc_2593 N_D[6]_M1143_g N_A_3891_297#_c_7358_n 0.0127833f $X=20.285 $Y=1.985
+ $X2=0 $Y2=0
cc_2594 N_D[6]_c_3293_n N_A_3891_297#_c_7358_n 0.0323774f $X=20.07 $Y=1.16 $X2=0
+ $Y2=0
cc_2595 N_D[6]_c_3294_n N_A_3891_297#_c_7358_n 7.13708e-19 $X=20.285 $Y=1.16
+ $X2=0 $Y2=0
cc_2596 N_D[6]_M1062_g N_A_3891_297#_c_7362_n 0.00244285f $X=19.815 $Y=1.985
+ $X2=0 $Y2=0
cc_2597 N_D[6]_M1143_g N_A_3891_297#_c_7362_n 0.00246916f $X=20.285 $Y=1.985
+ $X2=0 $Y2=0
cc_2598 N_D[6]_M1062_g N_A_3891_297#_c_7352_n 0.00290175f $X=19.815 $Y=1.985
+ $X2=0 $Y2=0
cc_2599 N_D[6]_M1143_g N_A_3891_297#_c_7365_n 0.00595395f $X=20.285 $Y=1.985
+ $X2=0 $Y2=0
cc_2600 N_D[6]_M1139_g N_VGND_c_7799_n 0.00430643f $X=19.84 $Y=0.56 $X2=0 $Y2=0
cc_2601 N_D[6]_M1139_g N_VGND_c_7801_n 0.0030929f $X=19.84 $Y=0.56 $X2=0 $Y2=0
cc_2602 N_D[6]_M1155_g N_VGND_c_7801_n 0.00300333f $X=20.26 $Y=0.56 $X2=0 $Y2=0
cc_2603 N_D[6]_M1155_g N_VGND_c_7819_n 0.00436487f $X=20.26 $Y=0.56 $X2=0 $Y2=0
cc_2604 N_D[6]_M1139_g VGND 0.00733187f $X=19.84 $Y=0.56 $X2=0 $Y2=0
cc_2605 N_D[6]_M1155_g VGND 0.00600262f $X=20.26 $Y=0.56 $X2=0 $Y2=0
cc_2606 N_D[6]_M1139_g N_A_3891_47#_c_8803_n 0.00633603f $X=19.84 $Y=0.56 $X2=0
+ $Y2=0
cc_2607 N_D[6]_M1155_g N_A_3891_47#_c_8803_n 5.29024e-19 $X=20.26 $Y=0.56 $X2=0
+ $Y2=0
cc_2608 N_D[6]_M1139_g N_A_3891_47#_c_8800_n 0.0084485f $X=19.84 $Y=0.56 $X2=0
+ $Y2=0
cc_2609 N_D[6]_M1155_g N_A_3891_47#_c_8800_n 0.0125955f $X=20.26 $Y=0.56 $X2=0
+ $Y2=0
cc_2610 N_D[6]_c_3293_n N_A_3891_47#_c_8800_n 0.0274027f $X=20.07 $Y=1.16 $X2=0
+ $Y2=0
cc_2611 N_D[6]_c_3294_n N_A_3891_47#_c_8800_n 0.00321151f $X=20.285 $Y=1.16
+ $X2=0 $Y2=0
cc_2612 N_D[6]_M1139_g N_A_3891_47#_c_8801_n 8.68782e-19 $X=19.84 $Y=0.56 $X2=0
+ $Y2=0
cc_2613 N_D[6]_c_3293_n N_A_3891_47#_c_8801_n 0.024456f $X=20.07 $Y=1.16 $X2=0
+ $Y2=0
cc_2614 N_D[6]_c_3294_n N_A_3891_47#_c_8801_n 0.00464565f $X=20.285 $Y=1.16
+ $X2=0 $Y2=0
cc_2615 N_D[14]_M1152_g N_A_4142_793#_M1006_g 0.0250718f $X=20.285 $Y=3.455
+ $X2=0 $Y2=0
cc_2616 N_D[14]_M1152_g N_A_4142_793#_c_3496_n 0.00671996f $X=20.285 $Y=3.455
+ $X2=0 $Y2=0
cc_2617 N_D[14]_M1119_g N_S[14]_c_3637_n 0.0165585f $X=20.26 $Y=4.88 $X2=-0.19
+ $Y2=-0.24
cc_2618 N_D[14]_M1069_g N_VPWR_c_4265_n 0.00338721f $X=19.815 $Y=3.455 $X2=0
+ $Y2=0
cc_2619 N_D[14]_M1152_g N_VPWR_c_4265_n 0.00847423f $X=20.285 $Y=3.455 $X2=0
+ $Y2=0
cc_2620 N_D[14]_M1069_g N_VPWR_c_4572_n 0.00311479f $X=19.815 $Y=3.455 $X2=0
+ $Y2=0
cc_2621 N_D[14]_M1152_g N_VPWR_c_4572_n 0.00295119f $X=20.285 $Y=3.455 $X2=0
+ $Y2=0
cc_2622 N_D[14]_M1069_g VPWR 0.00568683f $X=19.815 $Y=3.455 $X2=0 $Y2=0
cc_2623 N_D[14]_M1152_g VPWR 0.00350923f $X=20.285 $Y=3.455 $X2=0 $Y2=0
cc_2624 N_D[14]_M1069_g N_VPWR_c_4291_n 0.0033767f $X=19.815 $Y=3.455 $X2=0
+ $Y2=0
cc_2625 N_D[14]_M1152_g N_VPWR_c_4292_n 0.00342413f $X=20.285 $Y=3.455 $X2=0
+ $Y2=0
cc_2626 N_D[14]_M1119_g N_Z_c_5208_n 8.13311e-19 $X=20.26 $Y=4.88 $X2=0 $Y2=0
cc_2627 N_D[14]_M1152_g N_Z_c_5208_n 0.00112534f $X=20.285 $Y=3.455 $X2=0 $Y2=0
cc_2628 N_D[14]_c_3351_n N_Z_c_5208_n 0.00742792f $X=20.07 $Y=4.28 $X2=0 $Y2=0
cc_2629 N_D[14]_c_3352_n N_Z_c_5208_n 0.00583073f $X=20.285 $Y=4.28 $X2=0 $Y2=0
cc_2630 N_D[14]_M1069_g N_Z_c_5253_n 0.00312829f $X=19.815 $Y=3.455 $X2=0 $Y2=0
cc_2631 N_D[14]_M1152_g N_Z_c_5253_n 0.0033316f $X=20.285 $Y=3.455 $X2=0 $Y2=0
cc_2632 N_D[14]_c_3351_n N_Z_c_5253_n 0.00125914f $X=20.07 $Y=4.28 $X2=0 $Y2=0
cc_2633 N_D[14]_M1069_g N_A_3891_591#_c_7450_n 0.0101085f $X=19.815 $Y=3.455
+ $X2=0 $Y2=0
cc_2634 N_D[14]_M1152_g N_A_3891_591#_c_7450_n 0.0127833f $X=20.285 $Y=3.455
+ $X2=0 $Y2=0
cc_2635 N_D[14]_c_3351_n N_A_3891_591#_c_7450_n 0.0323774f $X=20.07 $Y=4.28
+ $X2=0 $Y2=0
cc_2636 N_D[14]_c_3352_n N_A_3891_591#_c_7450_n 7.13708e-19 $X=20.285 $Y=4.28
+ $X2=0 $Y2=0
cc_2637 N_D[14]_c_3351_n N_A_3891_591#_c_7446_n 0.0226682f $X=20.07 $Y=4.28
+ $X2=0 $Y2=0
cc_2638 N_D[14]_c_3352_n N_A_3891_591#_c_7446_n 9.6385e-19 $X=20.285 $Y=4.28
+ $X2=0 $Y2=0
cc_2639 N_D[14]_M1069_g N_A_3891_591#_c_7456_n 0.00244285f $X=19.815 $Y=3.455
+ $X2=0 $Y2=0
cc_2640 N_D[14]_M1152_g N_A_3891_591#_c_7456_n 0.00246473f $X=20.285 $Y=3.455
+ $X2=0 $Y2=0
cc_2641 N_D[14]_M1152_g N_A_3891_591#_c_7458_n 0.00531997f $X=20.285 $Y=3.455
+ $X2=0 $Y2=0
cc_2642 N_D[14]_M1069_g N_A_3891_591#_c_7449_n 0.00290175f $X=19.815 $Y=3.455
+ $X2=0 $Y2=0
cc_2643 N_D[14]_M1018_g N_VGND_c_7800_n 0.00430643f $X=19.84 $Y=4.88 $X2=0 $Y2=0
cc_2644 N_D[14]_M1018_g N_VGND_c_7802_n 0.0030929f $X=19.84 $Y=4.88 $X2=0 $Y2=0
cc_2645 N_D[14]_M1119_g N_VGND_c_7802_n 0.00300333f $X=20.26 $Y=4.88 $X2=0 $Y2=0
cc_2646 N_D[14]_M1119_g N_VGND_c_7821_n 0.00436487f $X=20.26 $Y=4.88 $X2=0 $Y2=0
cc_2647 N_D[14]_M1018_g VGND 0.00733187f $X=19.84 $Y=4.88 $X2=0 $Y2=0
cc_2648 N_D[14]_M1119_g VGND 0.00600262f $X=20.26 $Y=4.88 $X2=0 $Y2=0
cc_2649 N_D[14]_M1018_g N_A_3891_911#_c_8847_n 0.0084485f $X=19.84 $Y=4.88 $X2=0
+ $Y2=0
cc_2650 N_D[14]_M1119_g N_A_3891_911#_c_8847_n 0.0114493f $X=20.26 $Y=4.88 $X2=0
+ $Y2=0
cc_2651 N_D[14]_c_3351_n N_A_3891_911#_c_8847_n 0.0274027f $X=20.07 $Y=4.28
+ $X2=0 $Y2=0
cc_2652 N_D[14]_c_3352_n N_A_3891_911#_c_8847_n 0.0020061f $X=20.285 $Y=4.28
+ $X2=0 $Y2=0
cc_2653 N_D[14]_M1119_g N_A_3891_911#_c_8844_n 0.00114614f $X=20.26 $Y=4.88
+ $X2=0 $Y2=0
cc_2654 N_D[14]_c_3352_n N_A_3891_911#_c_8844_n 0.00120541f $X=20.285 $Y=4.28
+ $X2=0 $Y2=0
cc_2655 N_D[14]_M1018_g N_A_3891_911#_c_8846_n 0.00720482f $X=19.84 $Y=4.88
+ $X2=0 $Y2=0
cc_2656 N_D[14]_M1119_g N_A_3891_911#_c_8846_n 5.29024e-19 $X=20.26 $Y=4.88
+ $X2=0 $Y2=0
cc_2657 N_D[14]_c_3351_n N_A_3891_911#_c_8846_n 0.024456f $X=20.07 $Y=4.28 $X2=0
+ $Y2=0
cc_2658 N_D[14]_c_3352_n N_A_3891_911#_c_8846_n 0.00464565f $X=20.285 $Y=4.28
+ $X2=0 $Y2=0
cc_2659 N_A_4142_265#_M1066_g N_A_4142_793#_M1006_g 0.0130744f $X=20.81 $Y=2.075
+ $X2=0 $Y2=0
cc_2660 N_A_4142_265#_M1091_g N_A_4142_793#_M1140_g 0.0130744f $X=21.28 $Y=2.075
+ $X2=0 $Y2=0
cc_2661 N_A_4142_265#_c_3412_n N_S[6]_c_3571_n 0.00779314f $X=20.9 $Y=1.4
+ $X2=-0.19 $Y2=-0.24
cc_2662 N_A_4142_265#_c_3411_n N_S[6]_c_3574_n 0.00810157f $X=21.19 $Y=1.4 $X2=0
+ $Y2=0
cc_2663 N_A_4142_265#_c_3407_n N_S[6]_c_3574_n 7.04048e-19 $X=21.75 $Y=1.205
+ $X2=0 $Y2=0
cc_2664 N_A_4142_265#_c_3406_n N_S[6]_c_3576_n 0.0100587f $X=21.75 $Y=0.755
+ $X2=0 $Y2=0
cc_2665 N_A_4142_265#_c_3407_n N_S[6]_c_3576_n 0.00267287f $X=21.75 $Y=1.205
+ $X2=0 $Y2=0
cc_2666 N_A_4142_265#_c_3406_n N_S[6]_c_3577_n 0.0105766f $X=21.75 $Y=0.755
+ $X2=0 $Y2=0
cc_2667 N_A_4142_265#_c_3407_n N_S[6]_c_3577_n 0.0090765f $X=21.75 $Y=1.205
+ $X2=0 $Y2=0
cc_2668 N_A_4142_265#_c_3408_n N_S[6]_c_3577_n 0.00742826f $X=22.035 $Y=1.63
+ $X2=0 $Y2=0
cc_2669 N_A_4142_265#_c_3407_n N_S[6]_c_3578_n 0.00445422f $X=21.75 $Y=1.205
+ $X2=0 $Y2=0
cc_2670 N_A_4142_265#_c_3408_n N_S[6]_c_3578_n 4.25171e-19 $X=22.035 $Y=1.63
+ $X2=0 $Y2=0
cc_2671 N_A_4142_265#_c_3409_n N_S[6]_c_3578_n 0.00920672f $X=21.28 $Y=1.34
+ $X2=0 $Y2=0
cc_2672 N_A_4142_265#_c_3407_n N_S[6]_c_3579_n 0.00205356f $X=21.75 $Y=1.205
+ $X2=0 $Y2=0
cc_2673 N_A_4142_265#_c_3414_n N_S[6]_c_3579_n 0.00861299f $X=22.035 $Y=2.31
+ $X2=0 $Y2=0
cc_2674 N_A_4142_265#_c_3408_n N_S[6]_c_3579_n 0.00828481f $X=22.035 $Y=1.63
+ $X2=0 $Y2=0
cc_2675 N_A_4142_265#_c_3409_n N_S[6]_c_3579_n 0.00692516f $X=21.28 $Y=1.34
+ $X2=0 $Y2=0
cc_2676 N_A_4142_265#_c_3407_n N_S[6]_c_3580_n 0.00149517f $X=21.75 $Y=1.205
+ $X2=0 $Y2=0
cc_2677 N_A_4142_265#_c_3406_n S[6] 0.0061421f $X=21.75 $Y=0.755 $X2=0 $Y2=0
cc_2678 N_A_4142_265#_c_3407_n S[6] 0.0101733f $X=21.75 $Y=1.205 $X2=0 $Y2=0
cc_2679 N_A_4142_265#_c_3408_n S[6] 0.0127184f $X=22.035 $Y=1.63 $X2=0 $Y2=0
cc_2680 N_A_4142_265#_c_3409_n S[6] 3.07062e-19 $X=21.28 $Y=1.34 $X2=0 $Y2=0
cc_2681 N_A_4142_265#_M1066_g N_VPWR_c_4264_n 0.00107878f $X=20.81 $Y=2.075
+ $X2=0 $Y2=0
cc_2682 N_A_4142_265#_c_3414_n N_VPWR_c_4266_n 0.0321301f $X=22.035 $Y=2.31
+ $X2=0 $Y2=0
cc_2683 N_A_4142_265#_c_3408_n N_VPWR_c_4266_n 0.00732952f $X=22.035 $Y=1.63
+ $X2=0 $Y2=0
cc_2684 N_A_4142_265#_M1091_g N_VPWR_c_4276_n 8.06528e-19 $X=21.28 $Y=2.075
+ $X2=0 $Y2=0
cc_2685 N_A_4142_265#_c_3414_n N_VPWR_c_4276_n 0.0210596f $X=22.035 $Y=2.31
+ $X2=0 $Y2=0
cc_2686 N_A_4142_265#_M1077_s VPWR 0.00179197f $X=21.91 $Y=1.485 $X2=0 $Y2=0
cc_2687 N_A_4142_265#_M1066_g VPWR 0.00435072f $X=20.81 $Y=2.075 $X2=0 $Y2=0
cc_2688 N_A_4142_265#_M1091_g VPWR 0.0054792f $X=21.28 $Y=2.075 $X2=0 $Y2=0
cc_2689 N_A_4142_265#_c_3414_n VPWR 0.00594162f $X=22.035 $Y=2.31 $X2=0 $Y2=0
cc_2690 N_A_4142_265#_c_3411_n N_Z_c_5222_n 0.00168443f $X=21.19 $Y=1.4 $X2=0
+ $Y2=0
cc_2691 N_A_4142_265#_c_3412_n N_Z_c_5222_n 0.00180308f $X=20.9 $Y=1.4 $X2=0
+ $Y2=0
cc_2692 N_A_4142_265#_c_3407_n N_Z_c_5222_n 0.0033343f $X=21.75 $Y=1.205 $X2=0
+ $Y2=0
cc_2693 N_A_4142_265#_M1066_g N_Z_c_5252_n 0.00404618f $X=20.81 $Y=2.075 $X2=0
+ $Y2=0
cc_2694 N_A_4142_265#_M1091_g N_Z_c_5254_n 0.00708998f $X=21.28 $Y=2.075 $X2=0
+ $Y2=0
cc_2695 N_A_4142_265#_c_3414_n N_Z_c_5254_n 0.0308332f $X=22.035 $Y=2.31 $X2=0
+ $Y2=0
cc_2696 N_A_4142_265#_c_3408_n N_Z_c_5254_n 0.0132841f $X=22.035 $Y=1.63 $X2=0
+ $Y2=0
cc_2697 N_A_4142_265#_c_3409_n N_Z_c_5254_n 9.57301e-19 $X=21.28 $Y=1.34 $X2=0
+ $Y2=0
cc_2698 N_A_4142_265#_M1066_g N_Z_c_5706_n 0.00513826f $X=20.81 $Y=2.075 $X2=0
+ $Y2=0
cc_2699 N_A_4142_265#_M1066_g N_Z_c_5707_n 0.00978858f $X=20.81 $Y=2.075 $X2=0
+ $Y2=0
cc_2700 N_A_4142_265#_c_3411_n N_Z_c_5707_n 8.37785e-19 $X=21.19 $Y=1.4 $X2=0
+ $Y2=0
cc_2701 N_A_4142_265#_M1091_g N_Z_c_5707_n 0.00619657f $X=21.28 $Y=2.075 $X2=0
+ $Y2=0
cc_2702 N_A_4142_265#_M1066_g N_Z_c_5232_n 0.00268051f $X=20.81 $Y=2.075 $X2=0
+ $Y2=0
cc_2703 N_A_4142_265#_c_3411_n N_Z_c_5232_n 0.0140957f $X=21.19 $Y=1.4 $X2=0
+ $Y2=0
cc_2704 N_A_4142_265#_M1091_g N_Z_c_5232_n 0.00476154f $X=21.28 $Y=2.075 $X2=0
+ $Y2=0
cc_2705 N_A_4142_265#_c_3407_n N_Z_c_5232_n 0.00967956f $X=21.75 $Y=1.205 $X2=0
+ $Y2=0
cc_2706 N_A_4142_265#_c_3408_n N_Z_c_5232_n 0.0117695f $X=22.035 $Y=1.63 $X2=0
+ $Y2=0
cc_2707 N_A_4142_265#_c_3409_n N_Z_c_5232_n 7.26438e-19 $X=21.28 $Y=1.34 $X2=0
+ $Y2=0
cc_2708 N_A_4142_265#_M1066_g N_Z_c_5716_n 2.61869e-19 $X=20.81 $Y=2.075 $X2=0
+ $Y2=0
cc_2709 N_A_4142_265#_M1066_g N_Z_c_5269_n 0.00455034f $X=20.81 $Y=2.075 $X2=0
+ $Y2=0
cc_2710 N_A_4142_265#_M1091_g N_Z_c_5269_n 0.00462462f $X=21.28 $Y=2.075 $X2=0
+ $Y2=0
cc_2711 N_A_4142_265#_M1066_g N_A_3891_297#_c_7358_n 0.00176121f $X=20.81
+ $Y=2.075 $X2=0 $Y2=0
cc_2712 N_A_4142_265#_M1066_g N_A_3891_297#_c_7367_n 0.00463461f $X=20.81
+ $Y=2.075 $X2=0 $Y2=0
cc_2713 N_A_4142_265#_M1091_g N_A_3891_297#_c_7367_n 0.00334959f $X=21.28
+ $Y=2.075 $X2=0 $Y2=0
cc_2714 N_A_4142_265#_M1066_g N_A_3891_297#_c_7369_n 7.75952e-19 $X=20.81
+ $Y=2.075 $X2=0 $Y2=0
cc_2715 N_A_4142_265#_M1066_g N_A_3891_297#_c_7370_n 0.00415998f $X=20.81
+ $Y=2.075 $X2=0 $Y2=0
cc_2716 N_A_4142_265#_c_3414_n N_A_3891_297#_c_7353_n 0.00738363f $X=22.035
+ $Y=2.31 $X2=0 $Y2=0
cc_2717 N_A_4142_265#_M1091_g N_A_3891_297#_c_7372_n 0.00692695f $X=21.28
+ $Y=2.075 $X2=0 $Y2=0
cc_2718 N_A_4142_265#_M1066_g N_A_3891_297#_c_7365_n 0.00508488f $X=20.81
+ $Y=2.075 $X2=0 $Y2=0
cc_2719 N_A_4142_265#_M1091_g N_A_3891_297#_c_7354_n 0.00550198f $X=21.28
+ $Y=2.075 $X2=0 $Y2=0
cc_2720 N_A_4142_265#_c_3414_n N_A_3891_297#_c_7354_n 0.0413447f $X=22.035
+ $Y=2.31 $X2=0 $Y2=0
cc_2721 N_A_4142_265#_c_3408_n N_A_3891_297#_c_7354_n 0.0132748f $X=22.035
+ $Y=1.63 $X2=0 $Y2=0
cc_2722 N_A_4142_265#_c_3409_n N_A_3891_297#_c_7354_n 0.00133381f $X=21.28
+ $Y=1.34 $X2=0 $Y2=0
cc_2723 N_A_4142_265#_c_3406_n N_VGND_c_7819_n 0.0173492f $X=21.75 $Y=0.755
+ $X2=0 $Y2=0
cc_2724 N_A_4142_265#_M1144_s VGND 0.00250855f $X=21.995 $Y=0.235 $X2=0 $Y2=0
cc_2725 N_A_4142_265#_c_3406_n VGND 0.0186564f $X=21.75 $Y=0.755 $X2=0 $Y2=0
cc_2726 N_A_4142_265#_c_3406_n N_A_3891_47#_c_8802_n 0.00358194f $X=21.75
+ $Y=0.755 $X2=0 $Y2=0
cc_2727 N_A_4142_265#_c_3406_n N_A_3891_47#_c_8813_n 0.0185512f $X=21.75
+ $Y=0.755 $X2=0 $Y2=0
cc_2728 N_A_4142_265#_c_3407_n N_A_3891_47#_c_8813_n 0.00101918f $X=21.75
+ $Y=1.205 $X2=0 $Y2=0
cc_2729 N_A_4142_265#_c_3408_n N_A_3891_47#_c_8813_n 0.00285813f $X=22.035
+ $Y=1.63 $X2=0 $Y2=0
cc_2730 N_A_4142_265#_c_3409_n N_A_3891_47#_c_8813_n 0.00308807f $X=21.28
+ $Y=1.34 $X2=0 $Y2=0
cc_2731 N_A_4142_793#_c_3496_n N_S[14]_c_3637_n 0.00779314f $X=20.9 $Y=4.04
+ $X2=-0.19 $Y2=-0.24
cc_2732 N_A_4142_793#_c_3495_n N_S[14]_c_3640_n 0.00810157f $X=21.19 $Y=4.04
+ $X2=0 $Y2=0
cc_2733 N_A_4142_793#_c_3491_n N_S[14]_c_3640_n 7.04048e-19 $X=21.75 $Y=4.685
+ $X2=0 $Y2=0
cc_2734 N_A_4142_793#_c_3491_n N_S[14]_c_3642_n 0.0127103f $X=21.75 $Y=4.685
+ $X2=0 $Y2=0
cc_2735 N_A_4142_793#_c_3491_n N_S[14]_c_3643_n 0.0196531f $X=21.75 $Y=4.685
+ $X2=0 $Y2=0
cc_2736 N_A_4142_793#_c_3492_n N_S[14]_c_3643_n 0.00742826f $X=22.035 $Y=3.805
+ $X2=0 $Y2=0
cc_2737 N_A_4142_793#_c_3491_n N_S[14]_c_3644_n 0.00445422f $X=21.75 $Y=4.685
+ $X2=0 $Y2=0
cc_2738 N_A_4142_793#_c_3492_n N_S[14]_c_3644_n 4.25171e-19 $X=22.035 $Y=3.805
+ $X2=0 $Y2=0
cc_2739 N_A_4142_793#_c_3493_n N_S[14]_c_3644_n 0.00920672f $X=21.28 $Y=4.1
+ $X2=0 $Y2=0
cc_2740 N_A_4142_793#_c_3492_n N_S[14]_c_3648_n 0.00386817f $X=22.035 $Y=3.805
+ $X2=0 $Y2=0
cc_2741 N_A_4142_793#_c_3499_n N_S[14]_c_3648_n 0.00861299f $X=22.035 $Y=3.13
+ $X2=0 $Y2=0
cc_2742 N_A_4142_793#_c_3493_n N_S[14]_c_3648_n 0.00149275f $X=21.28 $Y=4.1
+ $X2=0 $Y2=0
cc_2743 N_A_4142_793#_c_3491_n N_S[14]_c_3645_n 0.00354873f $X=21.75 $Y=4.685
+ $X2=0 $Y2=0
cc_2744 N_A_4142_793#_c_3492_n N_S[14]_c_3645_n 0.00441664f $X=22.035 $Y=3.805
+ $X2=0 $Y2=0
cc_2745 N_A_4142_793#_c_3493_n N_S[14]_c_3645_n 0.00543241f $X=21.28 $Y=4.1
+ $X2=0 $Y2=0
cc_2746 N_A_4142_793#_c_3491_n S[14] 0.0163154f $X=21.75 $Y=4.685 $X2=0 $Y2=0
cc_2747 N_A_4142_793#_c_3492_n S[14] 0.0127184f $X=22.035 $Y=3.805 $X2=0 $Y2=0
cc_2748 N_A_4142_793#_c_3493_n S[14] 3.07062e-19 $X=21.28 $Y=4.1 $X2=0 $Y2=0
cc_2749 N_A_4142_793#_M1006_g N_VPWR_c_4265_n 0.0013032f $X=20.81 $Y=3.365 $X2=0
+ $Y2=0
cc_2750 N_A_4142_793#_c_3492_n N_VPWR_c_4267_n 0.00732952f $X=22.035 $Y=3.805
+ $X2=0 $Y2=0
cc_2751 N_A_4142_793#_c_3499_n N_VPWR_c_4267_n 0.0321301f $X=22.035 $Y=3.13
+ $X2=0 $Y2=0
cc_2752 N_A_4142_793#_M1140_g N_VPWR_c_4276_n 7.91347e-19 $X=21.28 $Y=3.365
+ $X2=0 $Y2=0
cc_2753 N_A_4142_793#_c_3499_n N_VPWR_c_4276_n 0.0210596f $X=22.035 $Y=3.13
+ $X2=0 $Y2=0
cc_2754 N_A_4142_793#_M1085_s VPWR 0.00179197f $X=21.91 $Y=2.955 $X2=0 $Y2=0
cc_2755 N_A_4142_793#_M1006_g VPWR 0.00434142f $X=20.81 $Y=3.365 $X2=0 $Y2=0
cc_2756 N_A_4142_793#_M1140_g VPWR 0.00546988f $X=21.28 $Y=3.365 $X2=0 $Y2=0
cc_2757 N_A_4142_793#_c_3499_n VPWR 0.00594162f $X=22.035 $Y=3.13 $X2=0 $Y2=0
cc_2758 N_A_4142_793#_M1006_g N_Z_c_5208_n 0.00268051f $X=20.81 $Y=3.365 $X2=0
+ $Y2=0
cc_2759 N_A_4142_793#_c_3495_n N_Z_c_5208_n 0.0140957f $X=21.19 $Y=4.04 $X2=0
+ $Y2=0
cc_2760 N_A_4142_793#_M1140_g N_Z_c_5208_n 0.00476154f $X=21.28 $Y=3.365 $X2=0
+ $Y2=0
cc_2761 N_A_4142_793#_c_3491_n N_Z_c_5208_n 0.00967956f $X=21.75 $Y=4.685 $X2=0
+ $Y2=0
cc_2762 N_A_4142_793#_c_3492_n N_Z_c_5208_n 0.0117695f $X=22.035 $Y=3.805 $X2=0
+ $Y2=0
cc_2763 N_A_4142_793#_c_3493_n N_Z_c_5208_n 7.26438e-19 $X=21.28 $Y=4.1 $X2=0
+ $Y2=0
cc_2764 N_A_4142_793#_c_3495_n N_Z_c_5223_n 0.00168443f $X=21.19 $Y=4.04 $X2=0
+ $Y2=0
cc_2765 N_A_4142_793#_c_3496_n N_Z_c_5223_n 0.00180308f $X=20.9 $Y=4.04 $X2=0
+ $Y2=0
cc_2766 N_A_4142_793#_c_3491_n N_Z_c_5223_n 0.0033343f $X=21.75 $Y=4.685 $X2=0
+ $Y2=0
cc_2767 N_A_4142_793#_M1006_g N_Z_c_5253_n 0.0040431f $X=20.81 $Y=3.365 $X2=0
+ $Y2=0
cc_2768 N_A_4142_793#_M1140_g N_Z_c_5255_n 0.00708682f $X=21.28 $Y=3.365 $X2=0
+ $Y2=0
cc_2769 N_A_4142_793#_c_3492_n N_Z_c_5255_n 0.0132841f $X=22.035 $Y=3.805 $X2=0
+ $Y2=0
cc_2770 N_A_4142_793#_c_3499_n N_Z_c_5255_n 0.0308332f $X=22.035 $Y=3.13 $X2=0
+ $Y2=0
cc_2771 N_A_4142_793#_c_3493_n N_Z_c_5255_n 9.57301e-19 $X=21.28 $Y=4.1 $X2=0
+ $Y2=0
cc_2772 N_A_4142_793#_M1006_g N_Z_c_5733_n 0.00513826f $X=20.81 $Y=3.365 $X2=0
+ $Y2=0
cc_2773 N_A_4142_793#_M1006_g N_Z_c_5707_n 2.61869e-19 $X=20.81 $Y=3.365 $X2=0
+ $Y2=0
cc_2774 N_A_4142_793#_M1006_g N_Z_c_5716_n 0.00978858f $X=20.81 $Y=3.365 $X2=0
+ $Y2=0
cc_2775 N_A_4142_793#_c_3495_n N_Z_c_5716_n 8.37785e-19 $X=21.19 $Y=4.04 $X2=0
+ $Y2=0
cc_2776 N_A_4142_793#_M1140_g N_Z_c_5716_n 0.00619657f $X=21.28 $Y=3.365 $X2=0
+ $Y2=0
cc_2777 N_A_4142_793#_M1006_g N_Z_c_5269_n 0.00455034f $X=20.81 $Y=3.365 $X2=0
+ $Y2=0
cc_2778 N_A_4142_793#_M1140_g N_Z_c_5269_n 0.00462236f $X=21.28 $Y=3.365 $X2=0
+ $Y2=0
cc_2779 N_A_4142_793#_M1006_g N_A_3891_591#_c_7450_n 0.00176121f $X=20.81
+ $Y=3.365 $X2=0 $Y2=0
cc_2780 N_A_4142_793#_M1006_g N_A_3891_591#_c_7461_n 0.00400484f $X=20.81
+ $Y=3.365 $X2=0 $Y2=0
cc_2781 N_A_4142_793#_M1140_g N_A_3891_591#_c_7447_n 0.0124482f $X=21.28
+ $Y=3.365 $X2=0 $Y2=0
cc_2782 N_A_4142_793#_c_3492_n N_A_3891_591#_c_7447_n 0.0132748f $X=22.035
+ $Y=3.805 $X2=0 $Y2=0
cc_2783 N_A_4142_793#_c_3499_n N_A_3891_591#_c_7447_n 0.0413753f $X=22.035
+ $Y=3.13 $X2=0 $Y2=0
cc_2784 N_A_4142_793#_c_3493_n N_A_3891_591#_c_7447_n 0.00133381f $X=21.28
+ $Y=4.1 $X2=0 $Y2=0
cc_2785 N_A_4142_793#_M1006_g N_A_3891_591#_c_7466_n 0.00470988f $X=20.81
+ $Y=3.365 $X2=0 $Y2=0
cc_2786 N_A_4142_793#_M1140_g N_A_3891_591#_c_7466_n 0.00334069f $X=21.28
+ $Y=3.365 $X2=0 $Y2=0
cc_2787 N_A_4142_793#_M1006_g N_A_3891_591#_c_7468_n 7.75952e-19 $X=20.81
+ $Y=3.365 $X2=0 $Y2=0
cc_2788 N_A_4142_793#_M1006_g N_A_3891_591#_c_7458_n 0.00508821f $X=20.81
+ $Y=3.365 $X2=0 $Y2=0
cc_2789 N_A_4142_793#_c_3499_n N_A_3891_591#_c_7448_n 0.00738293f $X=22.035
+ $Y=3.13 $X2=0 $Y2=0
cc_2790 N_A_4142_793#_c_3491_n N_VGND_c_7821_n 0.0173402f $X=21.75 $Y=4.685
+ $X2=0 $Y2=0
cc_2791 N_A_4142_793#_M1012_s VGND 0.00250855f $X=21.995 $Y=4.685 $X2=0 $Y2=0
cc_2792 N_A_4142_793#_c_3491_n VGND 0.0186503f $X=21.75 $Y=4.685 $X2=0 $Y2=0
cc_2793 N_A_4142_793#_c_3491_n N_A_3891_911#_c_8845_n 0.00358194f $X=21.75
+ $Y=4.685 $X2=0 $Y2=0
cc_2794 N_A_4142_793#_c_3491_n N_A_3891_911#_c_8858_n 0.0195704f $X=21.75
+ $Y=4.685 $X2=0 $Y2=0
cc_2795 N_A_4142_793#_c_3492_n N_A_3891_911#_c_8858_n 0.00285813f $X=22.035
+ $Y=3.805 $X2=0 $Y2=0
cc_2796 N_A_4142_793#_c_3493_n N_A_3891_911#_c_8858_n 0.00308807f $X=21.28
+ $Y=4.1 $X2=0 $Y2=0
cc_2797 N_S[6]_c_3579_n N_S[14]_c_3648_n 0.0130744f $X=22.27 $Y=1.41 $X2=0 $Y2=0
cc_2798 N_S[6]_c_3580_n N_S[7]_c_3703_n 0.0133556f $X=22.33 $Y=0.845 $X2=-0.19
+ $Y2=-0.24
cc_2799 N_S[6]_c_3579_n N_S[7]_c_3704_n 0.0418422f $X=22.27 $Y=1.41 $X2=0 $Y2=0
cc_2800 S[6] N_S[7]_c_3704_n 8.74983e-19 $X=22.225 $Y=1.105 $X2=0 $Y2=0
cc_2801 N_S[6]_c_3579_n S[7] 8.74983e-19 $X=22.27 $Y=1.41 $X2=0 $Y2=0
cc_2802 S[6] S[7] 0.0208489f $X=22.225 $Y=1.105 $X2=0 $Y2=0
cc_2803 N_S[6]_c_3579_n N_VPWR_c_4266_n 0.00456891f $X=22.27 $Y=1.41 $X2=0 $Y2=0
cc_2804 S[6] N_VPWR_c_4266_n 0.00569857f $X=22.225 $Y=1.105 $X2=0 $Y2=0
cc_2805 N_S[6]_c_3579_n N_VPWR_c_4276_n 0.0035837f $X=22.27 $Y=1.41 $X2=0 $Y2=0
cc_2806 N_S[6]_c_3579_n VPWR 0.00710985f $X=22.27 $Y=1.41 $X2=0 $Y2=0
cc_2807 N_S[6]_c_3571_n N_Z_c_5222_n 0.00413022f $X=20.78 $Y=0.255 $X2=0 $Y2=0
cc_2808 N_S[6]_c_3574_n N_Z_c_5222_n 0.00495983f $X=21.2 $Y=0.255 $X2=0 $Y2=0
cc_2809 N_S[6]_c_3576_n N_Z_c_5222_n 4.25992e-19 $X=21.685 $Y=0.845 $X2=0 $Y2=0
cc_2810 N_S[6]_c_3579_n N_Z_c_5254_n 0.00513674f $X=22.27 $Y=1.41 $X2=0 $Y2=0
cc_2811 S[6] N_Z_c_5254_n 0.00545567f $X=22.225 $Y=1.105 $X2=0 $Y2=0
cc_2812 N_S[6]_c_3571_n N_Z_c_5232_n 0.00199103f $X=20.78 $Y=0.255 $X2=0 $Y2=0
cc_2813 N_S[6]_c_3574_n N_Z_c_5232_n 0.00133607f $X=21.2 $Y=0.255 $X2=0 $Y2=0
cc_2814 N_S[6]_c_3580_n N_VGND_c_7803_n 0.00330937f $X=22.33 $Y=0.845 $X2=0
+ $Y2=0
cc_2815 N_S[6]_c_3573_n N_VGND_c_7819_n 0.0271255f $X=20.855 $Y=0.18 $X2=0 $Y2=0
cc_2816 N_S[6]_c_3580_n N_VGND_c_7819_n 0.00585385f $X=22.33 $Y=0.845 $X2=0
+ $Y2=0
cc_2817 N_S[6]_c_3572_n VGND 0.00642387f $X=21.125 $Y=0.18 $X2=0 $Y2=0
cc_2818 N_S[6]_c_3573_n VGND 0.00474746f $X=20.855 $Y=0.18 $X2=0 $Y2=0
cc_2819 N_S[6]_c_3575_n VGND 0.0193094f $X=21.61 $Y=0.18 $X2=0 $Y2=0
cc_2820 N_S[6]_c_3580_n VGND 0.0111218f $X=22.33 $Y=0.845 $X2=0 $Y2=0
cc_2821 N_S[6]_c_3581_n VGND 0.00366655f $X=21.2 $Y=0.18 $X2=0 $Y2=0
cc_2822 N_S[6]_c_3571_n N_A_3891_47#_c_8800_n 0.00139422f $X=20.78 $Y=0.255
+ $X2=0 $Y2=0
cc_2823 N_S[6]_c_3571_n N_A_3891_47#_c_8802_n 0.0132844f $X=20.78 $Y=0.255 $X2=0
+ $Y2=0
cc_2824 N_S[6]_c_3572_n N_A_3891_47#_c_8802_n 0.00211351f $X=21.125 $Y=0.18
+ $X2=0 $Y2=0
cc_2825 N_S[6]_c_3574_n N_A_3891_47#_c_8802_n 0.0126455f $X=21.2 $Y=0.255 $X2=0
+ $Y2=0
cc_2826 N_S[6]_c_3575_n N_A_3891_47#_c_8802_n 0.00436105f $X=21.61 $Y=0.18 $X2=0
+ $Y2=0
cc_2827 N_S[6]_c_3576_n N_A_3891_47#_c_8802_n 0.00349455f $X=21.685 $Y=0.845
+ $X2=0 $Y2=0
cc_2828 N_S[6]_c_3576_n N_A_3891_47#_c_8813_n 0.00295202f $X=21.685 $Y=0.845
+ $X2=0 $Y2=0
cc_2829 N_S[14]_c_3645_n N_S[15]_c_3766_n 0.0474978f $X=22.33 $Y=4.595 $X2=-0.19
+ $Y2=-0.24
cc_2830 S[14] N_S[15]_c_3766_n 8.74983e-19 $X=22.225 $Y=4.165 $X2=-0.19
+ $Y2=-0.24
cc_2831 N_S[14]_c_3648_n N_S[15]_c_3777_n 0.00770012f $X=22.27 $Y=4.03 $X2=0
+ $Y2=0
cc_2832 N_S[14]_c_3645_n S[15] 8.74983e-19 $X=22.33 $Y=4.595 $X2=0 $Y2=0
cc_2833 S[14] S[15] 0.0208489f $X=22.225 $Y=4.165 $X2=0 $Y2=0
cc_2834 N_S[14]_c_3648_n N_VPWR_c_4267_n 0.00362951f $X=22.27 $Y=4.03 $X2=0
+ $Y2=0
cc_2835 N_S[14]_c_3645_n N_VPWR_c_4267_n 9.39395e-19 $X=22.33 $Y=4.595 $X2=0
+ $Y2=0
cc_2836 S[14] N_VPWR_c_4267_n 0.00569857f $X=22.225 $Y=4.165 $X2=0 $Y2=0
cc_2837 N_S[14]_c_3648_n N_VPWR_c_4276_n 0.0035837f $X=22.27 $Y=4.03 $X2=0 $Y2=0
cc_2838 N_S[14]_c_3648_n VPWR 0.00710985f $X=22.27 $Y=4.03 $X2=0 $Y2=0
cc_2839 N_S[14]_c_3637_n N_Z_c_5208_n 0.00199103f $X=20.78 $Y=5.185 $X2=0 $Y2=0
cc_2840 N_S[14]_c_3640_n N_Z_c_5208_n 0.00133607f $X=21.2 $Y=5.185 $X2=0 $Y2=0
cc_2841 N_S[14]_c_3637_n N_Z_c_5223_n 0.00413022f $X=20.78 $Y=5.185 $X2=0 $Y2=0
cc_2842 N_S[14]_c_3640_n N_Z_c_5223_n 0.00495983f $X=21.2 $Y=5.185 $X2=0 $Y2=0
cc_2843 N_S[14]_c_3644_n N_Z_c_5223_n 4.25992e-19 $X=21.76 $Y=4.52 $X2=0 $Y2=0
cc_2844 N_S[14]_c_3648_n N_Z_c_5255_n 0.00477894f $X=22.27 $Y=4.03 $X2=0 $Y2=0
cc_2845 N_S[14]_c_3645_n N_Z_c_5255_n 3.57797e-19 $X=22.33 $Y=4.595 $X2=0 $Y2=0
cc_2846 S[14] N_Z_c_5255_n 0.00545567f $X=22.225 $Y=4.165 $X2=0 $Y2=0
cc_2847 N_S[14]_c_3645_n N_VGND_c_7804_n 0.00330937f $X=22.33 $Y=4.595 $X2=0
+ $Y2=0
cc_2848 N_S[14]_c_3639_n N_VGND_c_7821_n 0.0271255f $X=20.855 $Y=5.26 $X2=0
+ $Y2=0
cc_2849 N_S[14]_c_3645_n N_VGND_c_7821_n 0.00585385f $X=22.33 $Y=4.595 $X2=0
+ $Y2=0
cc_2850 N_S[14]_c_3638_n VGND 0.00642387f $X=21.125 $Y=5.26 $X2=0 $Y2=0
cc_2851 N_S[14]_c_3639_n VGND 0.00474746f $X=20.855 $Y=5.26 $X2=0 $Y2=0
cc_2852 N_S[14]_c_3641_n VGND 0.0193094f $X=21.61 $Y=5.26 $X2=0 $Y2=0
cc_2853 N_S[14]_c_3645_n VGND 0.0111218f $X=22.33 $Y=4.595 $X2=0 $Y2=0
cc_2854 N_S[14]_c_3646_n VGND 0.00366655f $X=21.2 $Y=5.26 $X2=0 $Y2=0
cc_2855 N_S[14]_c_3637_n N_A_3891_911#_c_8844_n 0.00139422f $X=20.78 $Y=5.185
+ $X2=0 $Y2=0
cc_2856 N_S[14]_c_3637_n N_A_3891_911#_c_8845_n 0.0132844f $X=20.78 $Y=5.185
+ $X2=0 $Y2=0
cc_2857 N_S[14]_c_3638_n N_A_3891_911#_c_8845_n 0.00211351f $X=21.125 $Y=5.26
+ $X2=0 $Y2=0
cc_2858 N_S[14]_c_3640_n N_A_3891_911#_c_8845_n 0.0126455f $X=21.2 $Y=5.185
+ $X2=0 $Y2=0
cc_2859 N_S[14]_c_3641_n N_A_3891_911#_c_8845_n 0.00436105f $X=21.61 $Y=5.26
+ $X2=0 $Y2=0
cc_2860 N_S[14]_c_3642_n N_A_3891_911#_c_8845_n 0.00349455f $X=21.685 $Y=5.185
+ $X2=0 $Y2=0
cc_2861 N_S[14]_c_3642_n N_A_3891_911#_c_8858_n 0.00295202f $X=21.685 $Y=5.185
+ $X2=0 $Y2=0
cc_2862 N_S[7]_c_3704_n N_S[15]_c_3777_n 0.0130744f $X=22.81 $Y=1.41 $X2=0 $Y2=0
cc_2863 N_S[7]_c_3711_n N_A_4565_47#_c_3837_n 0.00779314f $X=24.3 $Y=0.255 $X2=0
+ $Y2=0
cc_2864 N_S[7]_c_3704_n N_A_4565_47#_c_3832_n 0.00692516f $X=22.81 $Y=1.41 $X2=0
+ $Y2=0
cc_2865 N_S[7]_c_3705_n N_A_4565_47#_c_3832_n 0.00920672f $X=23.32 $Y=0.92 $X2=0
+ $Y2=0
cc_2866 N_S[7]_c_3709_n N_A_4565_47#_c_3832_n 0.00810157f $X=23.88 $Y=0.255
+ $X2=0 $Y2=0
cc_2867 S[7] N_A_4565_47#_c_3832_n 3.07062e-19 $X=22.685 $Y=1.105 $X2=0 $Y2=0
cc_2868 N_S[7]_c_3704_n N_A_4565_47#_c_3840_n 0.00861299f $X=22.81 $Y=1.41 $X2=0
+ $Y2=0
cc_2869 N_S[7]_c_3703_n N_A_4565_47#_c_3833_n 0.00149517f $X=22.75 $Y=0.845
+ $X2=0 $Y2=0
cc_2870 N_S[7]_c_3704_n N_A_4565_47#_c_3833_n 0.00205356f $X=22.81 $Y=1.41 $X2=0
+ $Y2=0
cc_2871 N_S[7]_c_3705_n N_A_4565_47#_c_3833_n 0.0135307f $X=23.32 $Y=0.92 $X2=0
+ $Y2=0
cc_2872 N_S[7]_c_3706_n N_A_4565_47#_c_3833_n 0.00267287f $X=23.395 $Y=0.845
+ $X2=0 $Y2=0
cc_2873 N_S[7]_c_3709_n N_A_4565_47#_c_3833_n 7.04048e-19 $X=23.88 $Y=0.255
+ $X2=0 $Y2=0
cc_2874 S[7] N_A_4565_47#_c_3833_n 0.0101733f $X=22.685 $Y=1.105 $X2=0 $Y2=0
cc_2875 N_S[7]_c_3704_n N_A_4565_47#_c_3834_n 0.0105766f $X=22.81 $Y=1.41 $X2=0
+ $Y2=0
cc_2876 N_S[7]_c_3706_n N_A_4565_47#_c_3834_n 0.0100587f $X=23.395 $Y=0.845
+ $X2=0 $Y2=0
cc_2877 S[7] N_A_4565_47#_c_3834_n 0.0061421f $X=22.685 $Y=1.105 $X2=0 $Y2=0
cc_2878 N_S[7]_c_3704_n N_A_4565_47#_c_3835_n 0.00828481f $X=22.81 $Y=1.41 $X2=0
+ $Y2=0
cc_2879 N_S[7]_c_3705_n N_A_4565_47#_c_3835_n 0.00785343f $X=23.32 $Y=0.92 $X2=0
+ $Y2=0
cc_2880 S[7] N_A_4565_47#_c_3835_n 0.0127184f $X=22.685 $Y=1.105 $X2=0 $Y2=0
cc_2881 N_S[7]_c_3710_n N_D[7]_M1024_g 0.0165585f $X=24.225 $Y=0.18 $X2=0 $Y2=0
cc_2882 N_S[7]_c_3704_n N_VPWR_c_4266_n 0.00456891f $X=22.81 $Y=1.41 $X2=0 $Y2=0
cc_2883 S[7] N_VPWR_c_4266_n 0.00569857f $X=22.685 $Y=1.105 $X2=0 $Y2=0
cc_2884 N_S[7]_c_3704_n VPWR 0.00710985f $X=22.81 $Y=1.41 $X2=0 $Y2=0
cc_2885 N_S[7]_c_3704_n N_VPWR_c_4293_n 0.0035837f $X=22.81 $Y=1.41 $X2=0 $Y2=0
cc_2886 N_S[7]_c_3706_n N_Z_c_5224_n 4.25992e-19 $X=23.395 $Y=0.845 $X2=0 $Y2=0
cc_2887 N_S[7]_c_3709_n N_Z_c_5224_n 0.00495983f $X=23.88 $Y=0.255 $X2=0 $Y2=0
cc_2888 N_S[7]_c_3711_n N_Z_c_5224_n 0.00413022f $X=24.3 $Y=0.255 $X2=0 $Y2=0
cc_2889 N_S[7]_c_3704_n N_Z_c_5254_n 0.00513674f $X=22.81 $Y=1.41 $X2=0 $Y2=0
cc_2890 S[7] N_Z_c_5254_n 0.00545567f $X=22.685 $Y=1.105 $X2=0 $Y2=0
cc_2891 N_S[7]_c_3709_n N_Z_c_5233_n 0.00133607f $X=23.88 $Y=0.255 $X2=0 $Y2=0
cc_2892 N_S[7]_c_3711_n N_Z_c_5233_n 0.00199103f $X=24.3 $Y=0.255 $X2=0 $Y2=0
cc_2893 N_S[7]_c_3703_n N_VGND_c_7803_n 0.00330937f $X=22.75 $Y=0.845 $X2=0
+ $Y2=0
cc_2894 N_S[7]_c_3703_n N_VGND_c_7823_n 0.00585385f $X=22.75 $Y=0.845 $X2=0
+ $Y2=0
cc_2895 N_S[7]_c_3708_n N_VGND_c_7823_n 0.0271255f $X=23.47 $Y=0.18 $X2=0 $Y2=0
cc_2896 N_S[7]_c_3703_n VGND 0.0111218f $X=22.75 $Y=0.845 $X2=0 $Y2=0
cc_2897 N_S[7]_c_3707_n VGND 0.0119932f $X=23.805 $Y=0.18 $X2=0 $Y2=0
cc_2898 N_S[7]_c_3708_n VGND 0.00731624f $X=23.47 $Y=0.18 $X2=0 $Y2=0
cc_2899 N_S[7]_c_3710_n VGND 0.0111713f $X=24.225 $Y=0.18 $X2=0 $Y2=0
cc_2900 N_S[7]_c_3712_n VGND 0.00366655f $X=23.88 $Y=0.18 $X2=0 $Y2=0
cc_2901 N_S[7]_c_3706_n N_A_4709_69#_c_8892_n 0.00295202f $X=23.395 $Y=0.845
+ $X2=0 $Y2=0
cc_2902 N_S[7]_c_3709_n N_A_4709_69#_c_8888_n 0.0126455f $X=23.88 $Y=0.255 $X2=0
+ $Y2=0
cc_2903 N_S[7]_c_3710_n N_A_4709_69#_c_8888_n 0.00211351f $X=24.225 $Y=0.18
+ $X2=0 $Y2=0
cc_2904 N_S[7]_c_3711_n N_A_4709_69#_c_8888_n 0.0132844f $X=24.3 $Y=0.255 $X2=0
+ $Y2=0
cc_2905 N_S[7]_c_3706_n N_A_4709_69#_c_8889_n 0.00349455f $X=23.395 $Y=0.845
+ $X2=0 $Y2=0
cc_2906 N_S[7]_c_3707_n N_A_4709_69#_c_8889_n 0.00436105f $X=23.805 $Y=0.18
+ $X2=0 $Y2=0
cc_2907 N_S[7]_c_3711_n N_A_4709_69#_c_8891_n 0.00139422f $X=24.3 $Y=0.255 $X2=0
+ $Y2=0
cc_2908 N_S[15]_c_3773_n N_A_4565_937#_c_3917_n 0.00779314f $X=24.3 $Y=5.185
+ $X2=0 $Y2=0
cc_2909 N_S[15]_c_3766_n N_A_4565_937#_c_3912_n 0.00543241f $X=22.75 $Y=4.595
+ $X2=0 $Y2=0
cc_2910 N_S[15]_c_3777_n N_A_4565_937#_c_3912_n 0.00149275f $X=22.81 $Y=4.03
+ $X2=0 $Y2=0
cc_2911 N_S[15]_c_3767_n N_A_4565_937#_c_3912_n 0.00920672f $X=23.32 $Y=4.52
+ $X2=0 $Y2=0
cc_2912 N_S[15]_c_3771_n N_A_4565_937#_c_3912_n 0.00810157f $X=23.88 $Y=5.185
+ $X2=0 $Y2=0
cc_2913 S[15] N_A_4565_937#_c_3912_n 3.07062e-19 $X=22.685 $Y=4.165 $X2=0 $Y2=0
cc_2914 N_S[15]_c_3777_n N_A_4565_937#_c_3920_n 0.00861299f $X=22.81 $Y=4.03
+ $X2=0 $Y2=0
cc_2915 N_S[15]_c_3766_n N_A_4565_937#_c_3913_n 0.00354873f $X=22.75 $Y=4.595
+ $X2=0 $Y2=0
cc_2916 N_S[15]_c_3767_n N_A_4565_937#_c_3913_n 0.0135307f $X=23.32 $Y=4.52
+ $X2=0 $Y2=0
cc_2917 N_S[15]_c_3768_n N_A_4565_937#_c_3913_n 0.00267287f $X=23.395 $Y=5.185
+ $X2=0 $Y2=0
cc_2918 N_S[15]_c_3771_n N_A_4565_937#_c_3913_n 7.04048e-19 $X=23.88 $Y=5.185
+ $X2=0 $Y2=0
cc_2919 S[15] N_A_4565_937#_c_3913_n 0.0101733f $X=22.685 $Y=4.165 $X2=0 $Y2=0
cc_2920 N_S[15]_c_3766_n N_A_4565_937#_c_3914_n 0.0105766f $X=22.75 $Y=4.595
+ $X2=0 $Y2=0
cc_2921 N_S[15]_c_3768_n N_A_4565_937#_c_3914_n 0.0100374f $X=23.395 $Y=5.185
+ $X2=0 $Y2=0
cc_2922 S[15] N_A_4565_937#_c_3914_n 0.0061421f $X=22.685 $Y=4.165 $X2=0 $Y2=0
cc_2923 N_S[15]_c_3766_n N_A_4565_937#_c_3915_n 0.00441664f $X=22.75 $Y=4.595
+ $X2=0 $Y2=0
cc_2924 N_S[15]_c_3777_n N_A_4565_937#_c_3915_n 0.00386817f $X=22.81 $Y=4.03
+ $X2=0 $Y2=0
cc_2925 N_S[15]_c_3767_n N_A_4565_937#_c_3915_n 0.00785343f $X=23.32 $Y=4.52
+ $X2=0 $Y2=0
cc_2926 S[15] N_A_4565_937#_c_3915_n 0.0127184f $X=22.685 $Y=4.165 $X2=0 $Y2=0
cc_2927 N_S[15]_c_3773_n N_D[15]_M1147_g 0.0165585f $X=24.3 $Y=5.185 $X2=0 $Y2=0
cc_2928 N_S[15]_c_3766_n N_VPWR_c_4267_n 9.39395e-19 $X=22.75 $Y=4.595 $X2=0
+ $Y2=0
cc_2929 N_S[15]_c_3777_n N_VPWR_c_4267_n 0.00362951f $X=22.81 $Y=4.03 $X2=0
+ $Y2=0
cc_2930 S[15] N_VPWR_c_4267_n 0.00569857f $X=22.685 $Y=4.165 $X2=0 $Y2=0
cc_2931 N_S[15]_c_3777_n VPWR 0.00710985f $X=22.81 $Y=4.03 $X2=0 $Y2=0
cc_2932 N_S[15]_c_3777_n N_VPWR_c_4293_n 0.0035837f $X=22.81 $Y=4.03 $X2=0 $Y2=0
cc_2933 N_S[15]_c_3771_n N_Z_c_5209_n 0.00133607f $X=23.88 $Y=5.185 $X2=0 $Y2=0
cc_2934 N_S[15]_c_3773_n N_Z_c_5209_n 0.00199103f $X=24.3 $Y=5.185 $X2=0 $Y2=0
cc_2935 N_S[15]_c_3767_n N_Z_c_5225_n 4.25992e-19 $X=23.32 $Y=4.52 $X2=0 $Y2=0
cc_2936 N_S[15]_c_3771_n N_Z_c_5225_n 0.00495983f $X=23.88 $Y=5.185 $X2=0 $Y2=0
cc_2937 N_S[15]_c_3773_n N_Z_c_5225_n 0.00413022f $X=24.3 $Y=5.185 $X2=0 $Y2=0
cc_2938 N_S[15]_c_3766_n N_Z_c_5255_n 3.57797e-19 $X=22.75 $Y=4.595 $X2=0 $Y2=0
cc_2939 N_S[15]_c_3777_n N_Z_c_5255_n 0.00477894f $X=22.81 $Y=4.03 $X2=0 $Y2=0
cc_2940 S[15] N_Z_c_5255_n 0.00545567f $X=22.685 $Y=4.165 $X2=0 $Y2=0
cc_2941 N_S[15]_c_3766_n N_VGND_c_7804_n 0.00330937f $X=22.75 $Y=4.595 $X2=0
+ $Y2=0
cc_2942 N_S[15]_c_3766_n N_VGND_c_7825_n 0.00585385f $X=22.75 $Y=4.595 $X2=0
+ $Y2=0
cc_2943 N_S[15]_c_3770_n N_VGND_c_7825_n 0.0271255f $X=23.47 $Y=5.26 $X2=0 $Y2=0
cc_2944 N_S[15]_c_3766_n VGND 0.0111218f $X=22.75 $Y=4.595 $X2=0 $Y2=0
cc_2945 N_S[15]_c_3769_n VGND 0.0119932f $X=23.805 $Y=5.26 $X2=0 $Y2=0
cc_2946 N_S[15]_c_3770_n VGND 0.00731624f $X=23.47 $Y=5.26 $X2=0 $Y2=0
cc_2947 N_S[15]_c_3772_n VGND 0.0111713f $X=24.225 $Y=5.26 $X2=0 $Y2=0
cc_2948 N_S[15]_c_3774_n VGND 0.00366655f $X=23.88 $Y=5.26 $X2=0 $Y2=0
cc_2949 N_S[15]_c_3768_n N_A_4709_915#_c_8938_n 0.00295202f $X=23.395 $Y=5.185
+ $X2=0 $Y2=0
cc_2950 N_S[15]_c_3771_n N_A_4709_915#_c_8934_n 0.0126455f $X=23.88 $Y=5.185
+ $X2=0 $Y2=0
cc_2951 N_S[15]_c_3772_n N_A_4709_915#_c_8934_n 0.00211351f $X=24.225 $Y=5.26
+ $X2=0 $Y2=0
cc_2952 N_S[15]_c_3773_n N_A_4709_915#_c_8934_n 0.0132844f $X=24.3 $Y=5.185
+ $X2=0 $Y2=0
cc_2953 N_S[15]_c_3768_n N_A_4709_915#_c_8935_n 0.00349455f $X=23.395 $Y=5.185
+ $X2=0 $Y2=0
cc_2954 N_S[15]_c_3769_n N_A_4709_915#_c_8935_n 0.00436105f $X=23.805 $Y=5.26
+ $X2=0 $Y2=0
cc_2955 N_S[15]_c_3773_n N_A_4709_915#_c_8936_n 0.00139422f $X=24.3 $Y=5.185
+ $X2=0 $Y2=0
cc_2956 N_A_4565_47#_M1122_g N_A_4565_937#_M1049_g 0.0130744f $X=23.8 $Y=2.075
+ $X2=0 $Y2=0
cc_2957 N_A_4565_47#_M1148_g N_A_4565_937#_M1076_g 0.0130744f $X=24.27 $Y=2.075
+ $X2=0 $Y2=0
cc_2958 N_A_4565_47#_c_3837_n N_D[7]_M1061_g 0.00671996f $X=24.18 $Y=1.4 $X2=0
+ $Y2=0
cc_2959 N_A_4565_47#_M1148_g N_D[7]_M1061_g 0.0241487f $X=24.27 $Y=2.075 $X2=0
+ $Y2=0
cc_2960 N_A_4565_47#_c_3840_n N_VPWR_c_4266_n 0.0321301f $X=23.045 $Y=2.31 $X2=0
+ $Y2=0
cc_2961 N_A_4565_47#_c_3835_n N_VPWR_c_4266_n 0.00732952f $X=23.33 $Y=1.42 $X2=0
+ $Y2=0
cc_2962 N_A_4565_47#_M1148_g N_VPWR_c_4268_n 0.00107878f $X=24.27 $Y=2.075 $X2=0
+ $Y2=0
cc_2963 N_A_4565_47#_M1129_d VPWR 0.00179197f $X=22.9 $Y=1.485 $X2=0 $Y2=0
cc_2964 N_A_4565_47#_M1122_g VPWR 0.0054792f $X=23.8 $Y=2.075 $X2=0 $Y2=0
cc_2965 N_A_4565_47#_M1148_g VPWR 0.00435072f $X=24.27 $Y=2.075 $X2=0 $Y2=0
cc_2966 N_A_4565_47#_c_3840_n VPWR 0.00594162f $X=23.045 $Y=2.31 $X2=0 $Y2=0
cc_2967 N_A_4565_47#_M1122_g N_VPWR_c_4293_n 8.06528e-19 $X=23.8 $Y=2.075 $X2=0
+ $Y2=0
cc_2968 N_A_4565_47#_c_3840_n N_VPWR_c_4293_n 0.0210596f $X=23.045 $Y=2.31 $X2=0
+ $Y2=0
cc_2969 N_A_4565_47#_c_3837_n N_Z_c_5224_n 0.00348752f $X=24.18 $Y=1.4 $X2=0
+ $Y2=0
cc_2970 N_A_4565_47#_c_3833_n N_Z_c_5224_n 0.0033343f $X=23.33 $Y=1.205 $X2=0
+ $Y2=0
cc_2971 N_A_4565_47#_M1122_g N_Z_c_5254_n 0.00708998f $X=23.8 $Y=2.075 $X2=0
+ $Y2=0
cc_2972 N_A_4565_47#_c_3832_n N_Z_c_5254_n 9.57301e-19 $X=23.89 $Y=1.4 $X2=0
+ $Y2=0
cc_2973 N_A_4565_47#_c_3840_n N_Z_c_5254_n 0.0308332f $X=23.045 $Y=2.31 $X2=0
+ $Y2=0
cc_2974 N_A_4565_47#_c_3835_n N_Z_c_5254_n 0.0132841f $X=23.33 $Y=1.42 $X2=0
+ $Y2=0
cc_2975 N_A_4565_47#_M1148_g Z 0.00635853f $X=24.27 $Y=2.075 $X2=0 $Y2=0
cc_2976 N_A_4565_47#_M1122_g N_Z_c_5777_n 0.00619657f $X=23.8 $Y=2.075 $X2=0
+ $Y2=0
cc_2977 N_A_4565_47#_c_3837_n N_Z_c_5777_n 8.37785e-19 $X=24.18 $Y=1.4 $X2=0
+ $Y2=0
cc_2978 N_A_4565_47#_M1148_g N_Z_c_5777_n 0.00978858f $X=24.27 $Y=2.075 $X2=0
+ $Y2=0
cc_2979 N_A_4565_47#_M1122_g N_Z_c_5233_n 0.00476154f $X=23.8 $Y=2.075 $X2=0
+ $Y2=0
cc_2980 N_A_4565_47#_c_3837_n N_Z_c_5233_n 0.0140957f $X=24.18 $Y=1.4 $X2=0
+ $Y2=0
cc_2981 N_A_4565_47#_c_3832_n N_Z_c_5233_n 7.26438e-19 $X=23.89 $Y=1.4 $X2=0
+ $Y2=0
cc_2982 N_A_4565_47#_M1148_g N_Z_c_5233_n 0.00268051f $X=24.27 $Y=2.075 $X2=0
+ $Y2=0
cc_2983 N_A_4565_47#_c_3833_n N_Z_c_5233_n 0.00967956f $X=23.33 $Y=1.205 $X2=0
+ $Y2=0
cc_2984 N_A_4565_47#_c_3835_n N_Z_c_5233_n 0.0117695f $X=23.33 $Y=1.42 $X2=0
+ $Y2=0
cc_2985 N_A_4565_47#_M1148_g N_Z_c_5786_n 2.61869e-19 $X=24.27 $Y=2.075 $X2=0
+ $Y2=0
cc_2986 N_A_4565_47#_M1122_g N_Z_c_5271_n 0.00462462f $X=23.8 $Y=2.075 $X2=0
+ $Y2=0
cc_2987 N_A_4565_47#_M1148_g N_Z_c_5271_n 0.00455034f $X=24.27 $Y=2.075 $X2=0
+ $Y2=0
cc_2988 N_A_4565_47#_M1148_g N_A_4688_333#_c_7542_n 0.00176121f $X=24.27
+ $Y=2.075 $X2=0 $Y2=0
cc_2989 N_A_4565_47#_M1122_g N_A_4688_333#_c_7543_n 0.00334959f $X=23.8 $Y=2.075
+ $X2=0 $Y2=0
cc_2990 N_A_4565_47#_M1148_g N_A_4688_333#_c_7543_n 0.00663284f $X=24.27
+ $Y=2.075 $X2=0 $Y2=0
cc_2991 N_A_4565_47#_c_3840_n N_A_4688_333#_c_7538_n 0.00738363f $X=23.045
+ $Y=2.31 $X2=0 $Y2=0
cc_2992 N_A_4565_47#_M1148_g N_A_4688_333#_c_7546_n 7.75952e-19 $X=24.27
+ $Y=2.075 $X2=0 $Y2=0
cc_2993 N_A_4565_47#_M1122_g N_A_4688_333#_c_7547_n 0.00692695f $X=23.8 $Y=2.075
+ $X2=0 $Y2=0
cc_2994 N_A_4565_47#_M1148_g N_A_4688_333#_c_7548_n 0.00415998f $X=24.27
+ $Y=2.075 $X2=0 $Y2=0
cc_2995 N_A_4565_47#_M1122_g N_A_4688_333#_c_7540_n 0.00550198f $X=23.8 $Y=2.075
+ $X2=0 $Y2=0
cc_2996 N_A_4565_47#_c_3832_n N_A_4688_333#_c_7540_n 0.00133381f $X=23.89 $Y=1.4
+ $X2=0 $Y2=0
cc_2997 N_A_4565_47#_c_3840_n N_A_4688_333#_c_7540_n 0.0413447f $X=23.045
+ $Y=2.31 $X2=0 $Y2=0
cc_2998 N_A_4565_47#_c_3835_n N_A_4688_333#_c_7540_n 0.0132748f $X=23.33 $Y=1.42
+ $X2=0 $Y2=0
cc_2999 N_A_4565_47#_M1148_g N_A_4688_333#_c_7553_n 0.00527462f $X=24.27
+ $Y=2.075 $X2=0 $Y2=0
cc_3000 N_A_4565_47#_c_3834_n N_VGND_c_7823_n 0.0173492f $X=22.96 $Y=0.495 $X2=0
+ $Y2=0
cc_3001 N_A_4565_47#_M1017_d VGND 0.00250855f $X=22.825 $Y=0.235 $X2=0 $Y2=0
cc_3002 N_A_4565_47#_c_3834_n VGND 0.0186564f $X=22.96 $Y=0.495 $X2=0 $Y2=0
cc_3003 N_A_4565_47#_c_3832_n N_A_4709_69#_c_8892_n 0.00308807f $X=23.89 $Y=1.4
+ $X2=0 $Y2=0
cc_3004 N_A_4565_47#_c_3833_n N_A_4709_69#_c_8892_n 0.00101918f $X=23.33
+ $Y=1.205 $X2=0 $Y2=0
cc_3005 N_A_4565_47#_c_3834_n N_A_4709_69#_c_8892_n 0.0185512f $X=22.96 $Y=0.495
+ $X2=0 $Y2=0
cc_3006 N_A_4565_47#_c_3835_n N_A_4709_69#_c_8892_n 0.00285813f $X=23.33 $Y=1.42
+ $X2=0 $Y2=0
cc_3007 N_A_4565_47#_c_3834_n N_A_4709_69#_c_8889_n 0.00358194f $X=22.96
+ $Y=0.495 $X2=0 $Y2=0
cc_3008 N_A_4565_937#_c_3917_n N_D[15]_M1068_g 0.00671996f $X=24.18 $Y=4.04
+ $X2=0 $Y2=0
cc_3009 N_A_4565_937#_M1076_g N_D[15]_M1068_g 0.0241475f $X=24.27 $Y=3.365 $X2=0
+ $Y2=0
cc_3010 N_A_4565_937#_c_3920_n N_VPWR_c_4267_n 0.0321301f $X=23.045 $Y=3.13
+ $X2=0 $Y2=0
cc_3011 N_A_4565_937#_c_3915_n N_VPWR_c_4267_n 0.00732952f $X=23.33 $Y=4.02
+ $X2=0 $Y2=0
cc_3012 N_A_4565_937#_M1076_g N_VPWR_c_4269_n 0.0012647f $X=24.27 $Y=3.365 $X2=0
+ $Y2=0
cc_3013 N_A_4565_937#_M1132_d VPWR 0.00179197f $X=22.9 $Y=2.955 $X2=0 $Y2=0
cc_3014 N_A_4565_937#_M1049_g VPWR 0.00546988f $X=23.8 $Y=3.365 $X2=0 $Y2=0
cc_3015 N_A_4565_937#_M1076_g VPWR 0.00434142f $X=24.27 $Y=3.365 $X2=0 $Y2=0
cc_3016 N_A_4565_937#_c_3920_n VPWR 0.00594162f $X=23.045 $Y=3.13 $X2=0 $Y2=0
cc_3017 N_A_4565_937#_M1049_g N_VPWR_c_4293_n 7.91347e-19 $X=23.8 $Y=3.365 $X2=0
+ $Y2=0
cc_3018 N_A_4565_937#_c_3920_n N_VPWR_c_4293_n 0.0210596f $X=23.045 $Y=3.13
+ $X2=0 $Y2=0
cc_3019 N_A_4565_937#_M1049_g N_Z_c_5209_n 0.00476154f $X=23.8 $Y=3.365 $X2=0
+ $Y2=0
cc_3020 N_A_4565_937#_c_3917_n N_Z_c_5209_n 0.0140957f $X=24.18 $Y=4.04 $X2=0
+ $Y2=0
cc_3021 N_A_4565_937#_c_3912_n N_Z_c_5209_n 7.26438e-19 $X=23.89 $Y=4.04 $X2=0
+ $Y2=0
cc_3022 N_A_4565_937#_M1076_g N_Z_c_5209_n 0.00268051f $X=24.27 $Y=3.365 $X2=0
+ $Y2=0
cc_3023 N_A_4565_937#_c_3913_n N_Z_c_5209_n 0.00967956f $X=23.33 $Y=4.685 $X2=0
+ $Y2=0
cc_3024 N_A_4565_937#_c_3915_n N_Z_c_5209_n 0.0117695f $X=23.33 $Y=4.02 $X2=0
+ $Y2=0
cc_3025 N_A_4565_937#_c_3917_n N_Z_c_5225_n 0.00348752f $X=24.18 $Y=4.04 $X2=0
+ $Y2=0
cc_3026 N_A_4565_937#_c_3913_n N_Z_c_5225_n 0.0033343f $X=23.33 $Y=4.685 $X2=0
+ $Y2=0
cc_3027 N_A_4565_937#_M1049_g N_Z_c_5255_n 0.00708682f $X=23.8 $Y=3.365 $X2=0
+ $Y2=0
cc_3028 N_A_4565_937#_c_3912_n N_Z_c_5255_n 9.57301e-19 $X=23.89 $Y=4.04 $X2=0
+ $Y2=0
cc_3029 N_A_4565_937#_c_3920_n N_Z_c_5255_n 0.0308332f $X=23.045 $Y=3.13 $X2=0
+ $Y2=0
cc_3030 N_A_4565_937#_c_3915_n N_Z_c_5255_n 0.0132841f $X=23.33 $Y=4.02 $X2=0
+ $Y2=0
cc_3031 N_A_4565_937#_M1076_g Z 0.00635853f $X=24.27 $Y=3.365 $X2=0 $Y2=0
cc_3032 N_A_4565_937#_M1076_g N_Z_c_5777_n 2.61869e-19 $X=24.27 $Y=3.365 $X2=0
+ $Y2=0
cc_3033 N_A_4565_937#_M1049_g N_Z_c_5786_n 0.00619657f $X=23.8 $Y=3.365 $X2=0
+ $Y2=0
cc_3034 N_A_4565_937#_c_3917_n N_Z_c_5786_n 8.37785e-19 $X=24.18 $Y=4.04 $X2=0
+ $Y2=0
cc_3035 N_A_4565_937#_M1076_g N_Z_c_5786_n 0.00978858f $X=24.27 $Y=3.365 $X2=0
+ $Y2=0
cc_3036 N_A_4565_937#_M1049_g N_Z_c_5271_n 0.00462236f $X=23.8 $Y=3.365 $X2=0
+ $Y2=0
cc_3037 N_A_4565_937#_M1076_g N_Z_c_5271_n 0.00455034f $X=24.27 $Y=3.365 $X2=0
+ $Y2=0
cc_3038 N_A_4565_937#_M1076_g N_A_4688_591#_c_7622_n 0.00176121f $X=24.27
+ $Y=3.365 $X2=0 $Y2=0
cc_3039 N_A_4565_937#_M1049_g N_A_4688_591#_c_7619_n 0.0124482f $X=23.8 $Y=3.365
+ $X2=0 $Y2=0
cc_3040 N_A_4565_937#_c_3912_n N_A_4688_591#_c_7619_n 0.00133381f $X=23.89
+ $Y=4.04 $X2=0 $Y2=0
cc_3041 N_A_4565_937#_c_3920_n N_A_4688_591#_c_7619_n 0.0413753f $X=23.045
+ $Y=3.13 $X2=0 $Y2=0
cc_3042 N_A_4565_937#_c_3915_n N_A_4688_591#_c_7619_n 0.0132748f $X=23.33
+ $Y=4.02 $X2=0 $Y2=0
cc_3043 N_A_4565_937#_M1076_g N_A_4688_591#_c_7627_n 0.00400484f $X=24.27
+ $Y=3.365 $X2=0 $Y2=0
cc_3044 N_A_4565_937#_M1049_g N_A_4688_591#_c_7628_n 0.00334069f $X=23.8
+ $Y=3.365 $X2=0 $Y2=0
cc_3045 N_A_4565_937#_M1076_g N_A_4688_591#_c_7628_n 0.00670811f $X=24.27
+ $Y=3.365 $X2=0 $Y2=0
cc_3046 N_A_4565_937#_c_3920_n N_A_4688_591#_c_7620_n 0.00738293f $X=23.045
+ $Y=3.13 $X2=0 $Y2=0
cc_3047 N_A_4565_937#_M1076_g N_A_4688_591#_c_7631_n 7.75952e-19 $X=24.27
+ $Y=3.365 $X2=0 $Y2=0
cc_3048 N_A_4565_937#_M1076_g N_A_4688_591#_c_7632_n 0.00527796f $X=24.27
+ $Y=3.365 $X2=0 $Y2=0
cc_3049 N_A_4565_937#_c_3914_n N_VGND_c_7825_n 0.0173402f $X=22.96 $Y=4.945
+ $X2=0 $Y2=0
cc_3050 N_A_4565_937#_M1040_d VGND 0.00250855f $X=22.825 $Y=4.685 $X2=0 $Y2=0
cc_3051 N_A_4565_937#_c_3914_n VGND 0.0186503f $X=22.96 $Y=4.945 $X2=0 $Y2=0
cc_3052 N_A_4565_937#_c_3912_n N_A_4709_915#_c_8938_n 0.00308807f $X=23.89
+ $Y=4.04 $X2=0 $Y2=0
cc_3053 N_A_4565_937#_c_3913_n N_A_4709_915#_c_8938_n 0.00101918f $X=23.33
+ $Y=4.685 $X2=0 $Y2=0
cc_3054 N_A_4565_937#_c_3914_n N_A_4709_915#_c_8938_n 0.0185512f $X=22.96
+ $Y=4.945 $X2=0 $Y2=0
cc_3055 N_A_4565_937#_c_3915_n N_A_4709_915#_c_8938_n 0.00285813f $X=23.33
+ $Y=4.02 $X2=0 $Y2=0
cc_3056 N_A_4565_937#_c_3914_n N_A_4709_915#_c_8935_n 0.00358194f $X=22.96
+ $Y=4.945 $X2=0 $Y2=0
cc_3057 N_D[7]_M1061_g N_D[15]_M1068_g 0.0129371f $X=24.795 $Y=1.985 $X2=0 $Y2=0
cc_3058 N_D[7]_M1142_g N_D[15]_M1149_g 0.0130744f $X=25.265 $Y=1.985 $X2=0 $Y2=0
cc_3059 N_D[7]_M1061_g N_VPWR_c_4268_n 0.00848021f $X=24.795 $Y=1.985 $X2=0
+ $Y2=0
cc_3060 N_D[7]_M1142_g N_VPWR_c_4268_n 0.00338721f $X=25.265 $Y=1.985 $X2=0
+ $Y2=0
cc_3061 N_D[7]_M1061_g N_VPWR_c_4634_n 0.00343746f $X=24.795 $Y=1.985 $X2=0
+ $Y2=0
cc_3062 N_D[7]_M1142_g N_VPWR_c_4634_n 0.00359955f $X=25.265 $Y=1.985 $X2=0
+ $Y2=0
cc_3063 N_D[7]_M1061_g VPWR 0.00350923f $X=24.795 $Y=1.985 $X2=0 $Y2=0
cc_3064 N_D[7]_M1142_g VPWR 0.00531592f $X=25.265 $Y=1.985 $X2=0 $Y2=0
cc_3065 N_D[7]_M1061_g N_VPWR_c_4294_n 0.00342413f $X=24.795 $Y=1.985 $X2=0
+ $Y2=0
cc_3066 N_D[7]_M1142_g N_VPWR_c_4295_n 0.0033767f $X=25.265 $Y=1.985 $X2=0 $Y2=0
cc_3067 N_D[7]_M1061_g N_Z_c_5233_n 0.00112534f $X=24.795 $Y=1.985 $X2=0 $Y2=0
cc_3068 N_D[7]_M1024_g N_Z_c_5233_n 8.13311e-19 $X=24.82 $Y=0.56 $X2=0 $Y2=0
cc_3069 D[7] N_Z_c_5233_n 0.00742792f $X=25.445 $Y=1.105 $X2=0 $Y2=0
cc_3070 N_D[7]_c_3997_n N_Z_c_5233_n 0.00583073f $X=25.35 $Y=1.16 $X2=0 $Y2=0
cc_3071 N_D[7]_M1061_g N_A_4688_333#_c_7554_n 0.0138742f $X=24.795 $Y=1.985
+ $X2=0 $Y2=0
cc_3072 N_D[7]_M1142_g N_A_4688_333#_c_7554_n 0.0111151f $X=25.265 $Y=1.985
+ $X2=0 $Y2=0
cc_3073 D[7] N_A_4688_333#_c_7554_n 0.0339353f $X=25.445 $Y=1.105 $X2=0 $Y2=0
cc_3074 N_D[7]_c_3997_n N_A_4688_333#_c_7554_n 7.13708e-19 $X=25.35 $Y=1.16
+ $X2=0 $Y2=0
cc_3075 D[7] N_A_4688_333#_c_7537_n 0.0235932f $X=25.445 $Y=1.105 $X2=0 $Y2=0
cc_3076 N_D[7]_c_3997_n N_A_4688_333#_c_7537_n 9.6385e-19 $X=25.35 $Y=1.16 $X2=0
+ $Y2=0
cc_3077 N_D[7]_M1061_g N_A_4688_333#_c_7560_n 0.00330676f $X=24.795 $Y=1.985
+ $X2=0 $Y2=0
cc_3078 N_D[7]_M1142_g N_A_4688_333#_c_7560_n 0.00332247f $X=25.265 $Y=1.985
+ $X2=0 $Y2=0
cc_3079 N_D[7]_M1142_g N_A_4688_333#_c_7539_n 0.00290175f $X=25.265 $Y=1.985
+ $X2=0 $Y2=0
cc_3080 N_D[7]_M1061_g N_A_4688_333#_c_7553_n 0.00611417f $X=24.795 $Y=1.985
+ $X2=0 $Y2=0
cc_3081 N_D[7]_M1024_g N_VGND_c_7805_n 0.00300333f $X=24.82 $Y=0.56 $X2=0 $Y2=0
cc_3082 N_D[7]_M1050_g N_VGND_c_7805_n 0.0030929f $X=25.24 $Y=0.56 $X2=0 $Y2=0
cc_3083 N_D[7]_M1024_g N_VGND_c_7823_n 0.00436487f $X=24.82 $Y=0.56 $X2=0 $Y2=0
cc_3084 N_D[7]_M1024_g VGND 0.00600262f $X=24.82 $Y=0.56 $X2=0 $Y2=0
cc_3085 N_D[7]_M1050_g VGND 0.00697949f $X=25.24 $Y=0.56 $X2=0 $Y2=0
cc_3086 N_D[7]_M1050_g N_VGND_c_7835_n 0.00430643f $X=25.24 $Y=0.56 $X2=0 $Y2=0
cc_3087 N_D[7]_M1024_g N_A_4709_69#_c_8890_n 0.0114493f $X=24.82 $Y=0.56 $X2=0
+ $Y2=0
cc_3088 N_D[7]_M1050_g N_A_4709_69#_c_8890_n 0.00931728f $X=25.24 $Y=0.56 $X2=0
+ $Y2=0
cc_3089 D[7] N_A_4709_69#_c_8890_n 0.0518587f $X=25.445 $Y=1.105 $X2=0 $Y2=0
cc_3090 N_D[7]_c_3997_n N_A_4709_69#_c_8890_n 0.00665175f $X=25.35 $Y=1.16 $X2=0
+ $Y2=0
cc_3091 N_D[7]_M1024_g N_A_4709_69#_c_8891_n 0.00114614f $X=24.82 $Y=0.56 $X2=0
+ $Y2=0
cc_3092 N_D[7]_c_3997_n N_A_4709_69#_c_8891_n 0.00120541f $X=25.35 $Y=1.16 $X2=0
+ $Y2=0
cc_3093 N_D[7]_M1024_g N_A_4709_69#_c_8910_n 5.29024e-19 $X=24.82 $Y=0.56 $X2=0
+ $Y2=0
cc_3094 N_D[7]_M1050_g N_A_4709_69#_c_8910_n 0.00633603f $X=25.24 $Y=0.56 $X2=0
+ $Y2=0
cc_3095 N_D[15]_M1068_g N_VPWR_c_4269_n 0.00847423f $X=24.795 $Y=3.455 $X2=0
+ $Y2=0
cc_3096 N_D[15]_M1149_g N_VPWR_c_4269_n 0.00338721f $X=25.265 $Y=3.455 $X2=0
+ $Y2=0
cc_3097 N_D[15]_M1068_g N_VPWR_c_4642_n 0.00343746f $X=24.795 $Y=3.455 $X2=0
+ $Y2=0
cc_3098 N_D[15]_M1149_g N_VPWR_c_4642_n 0.00359955f $X=25.265 $Y=3.455 $X2=0
+ $Y2=0
cc_3099 N_D[15]_M1068_g VPWR 0.00350923f $X=24.795 $Y=3.455 $X2=0 $Y2=0
cc_3100 N_D[15]_M1149_g VPWR 0.00531592f $X=25.265 $Y=3.455 $X2=0 $Y2=0
cc_3101 N_D[15]_M1068_g N_VPWR_c_4294_n 0.00342413f $X=24.795 $Y=3.455 $X2=0
+ $Y2=0
cc_3102 N_D[15]_M1149_g N_VPWR_c_4295_n 0.0033767f $X=25.265 $Y=3.455 $X2=0
+ $Y2=0
cc_3103 N_D[15]_M1068_g N_Z_c_5209_n 0.00112534f $X=24.795 $Y=3.455 $X2=0 $Y2=0
cc_3104 N_D[15]_M1147_g N_Z_c_5209_n 8.13311e-19 $X=24.82 $Y=4.88 $X2=0 $Y2=0
cc_3105 D[15] N_Z_c_5209_n 0.00742792f $X=25.445 $Y=4.165 $X2=0 $Y2=0
cc_3106 N_D[15]_c_4047_n N_Z_c_5209_n 0.00583073f $X=25.35 $Y=4.28 $X2=0 $Y2=0
cc_3107 N_D[15]_M1068_g N_A_4688_591#_c_7617_n 0.0138742f $X=24.795 $Y=3.455
+ $X2=0 $Y2=0
cc_3108 N_D[15]_M1149_g N_A_4688_591#_c_7617_n 0.0111151f $X=25.265 $Y=3.455
+ $X2=0 $Y2=0
cc_3109 D[15] N_A_4688_591#_c_7617_n 0.0575286f $X=25.445 $Y=4.165 $X2=0 $Y2=0
cc_3110 N_D[15]_c_4047_n N_A_4688_591#_c_7617_n 0.00167756f $X=25.35 $Y=4.28
+ $X2=0 $Y2=0
cc_3111 N_D[15]_M1068_g N_A_4688_591#_c_7637_n 0.00330232f $X=24.795 $Y=3.455
+ $X2=0 $Y2=0
cc_3112 N_D[15]_M1149_g N_A_4688_591#_c_7637_n 0.00332247f $X=25.265 $Y=3.455
+ $X2=0 $Y2=0
cc_3113 N_D[15]_M1068_g N_A_4688_591#_c_7632_n 0.00548019f $X=24.795 $Y=3.455
+ $X2=0 $Y2=0
cc_3114 N_D[15]_M1149_g N_A_4688_591#_c_7621_n 0.00290175f $X=25.265 $Y=3.455
+ $X2=0 $Y2=0
cc_3115 N_D[15]_M1147_g N_VGND_c_7806_n 0.00300333f $X=24.82 $Y=4.88 $X2=0 $Y2=0
cc_3116 N_D[15]_M1154_g N_VGND_c_7806_n 0.0030929f $X=25.24 $Y=4.88 $X2=0 $Y2=0
cc_3117 N_D[15]_M1147_g N_VGND_c_7825_n 0.00436487f $X=24.82 $Y=4.88 $X2=0 $Y2=0
cc_3118 N_D[15]_M1147_g VGND 0.00600262f $X=24.82 $Y=4.88 $X2=0 $Y2=0
cc_3119 N_D[15]_M1154_g VGND 0.00697949f $X=25.24 $Y=4.88 $X2=0 $Y2=0
cc_3120 N_D[15]_M1154_g N_VGND_c_7836_n 0.00430643f $X=25.24 $Y=4.88 $X2=0 $Y2=0
cc_3121 N_D[15]_M1147_g N_A_4709_915#_c_8936_n 0.00114614f $X=24.82 $Y=4.88
+ $X2=0 $Y2=0
cc_3122 N_D[15]_c_4047_n N_A_4709_915#_c_8936_n 0.00120541f $X=25.35 $Y=4.28
+ $X2=0 $Y2=0
cc_3123 N_D[15]_M1147_g N_A_4709_915#_c_8952_n 0.0114493f $X=24.82 $Y=4.88 $X2=0
+ $Y2=0
cc_3124 N_D[15]_M1154_g N_A_4709_915#_c_8952_n 0.0084485f $X=25.24 $Y=4.88 $X2=0
+ $Y2=0
cc_3125 D[15] N_A_4709_915#_c_8952_n 0.0274027f $X=25.445 $Y=4.165 $X2=0 $Y2=0
cc_3126 N_D[15]_c_4047_n N_A_4709_915#_c_8952_n 0.0020061f $X=25.35 $Y=4.28
+ $X2=0 $Y2=0
cc_3127 N_D[15]_M1147_g N_A_4709_915#_c_8937_n 5.29024e-19 $X=24.82 $Y=4.88
+ $X2=0 $Y2=0
cc_3128 N_D[15]_M1154_g N_A_4709_915#_c_8937_n 0.00720482f $X=25.24 $Y=4.88
+ $X2=0 $Y2=0
cc_3129 D[15] N_A_4709_915#_c_8937_n 0.024456f $X=25.445 $Y=4.165 $X2=0 $Y2=0
cc_3130 N_D[15]_c_4047_n N_A_4709_915#_c_8937_n 0.00464565f $X=25.35 $Y=4.28
+ $X2=0 $Y2=0
cc_3131 N_A_27_297#_c_4099_n N_VPWR_M1010_s 0.00346031f $X=1.115 $Y=1.58
+ $X2=-0.19 $Y2=1.305
cc_3132 N_A_27_297#_c_4103_n N_VPWR_c_4246_n 0.0174313f $X=1.055 $Y=2.225 $X2=0
+ $Y2=0
cc_3133 N_A_27_297#_c_4121_p N_VPWR_c_4246_n 0.00163482f $X=0.405 $Y=2.225 $X2=0
+ $Y2=0
cc_3134 N_A_27_297#_c_4110_n N_VPWR_c_4246_n 0.00265921f $X=1.345 $Y=2.225 $X2=0
+ $Y2=0
cc_3135 N_A_27_297#_c_4093_n N_VPWR_c_4246_n 0.0106781f $X=0.26 $Y=2.225 $X2=0
+ $Y2=0
cc_3136 N_A_27_297#_c_4111_n N_VPWR_c_4246_n 0.0177079f $X=1.2 $Y=2.225 $X2=0
+ $Y2=0
cc_3137 N_A_27_297#_c_4096_n N_VPWR_c_4246_n 0.00235484f $X=0.26 $Y=2.21 $X2=0
+ $Y2=0
cc_3138 N_A_27_297#_c_4099_n N_VPWR_c_4306_n 0.0164726f $X=1.115 $Y=1.58 $X2=0
+ $Y2=0
cc_3139 N_A_27_297#_c_4103_n N_VPWR_c_4306_n 8.54514e-19 $X=1.055 $Y=2.225 $X2=0
+ $Y2=0
cc_3140 N_A_27_297#_c_4106_n N_VPWR_c_4306_n 0.0177079f $X=1.2 $Y=1.78 $X2=0
+ $Y2=0
cc_3141 N_A_27_297#_c_4094_n N_VPWR_c_4270_n 4.83649e-19 $X=2.195 $Y=2.225 $X2=0
+ $Y2=0
cc_3142 N_A_27_297#_c_4113_n N_VPWR_c_4270_n 0.0217548f $X=2.195 $Y=2.225 $X2=0
+ $Y2=0
cc_3143 N_A_27_297#_M1010_d VPWR 0.00111289f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_3144 N_A_27_297#_M1075_d VPWR 0.00166446f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_3145 N_A_27_297#_M1031_d VPWR 0.00127816f $X=2.05 $Y=1.665 $X2=0 $Y2=0
cc_3146 N_A_27_297#_c_4103_n VPWR 0.0560119f $X=1.055 $Y=2.225 $X2=0 $Y2=0
cc_3147 N_A_27_297#_c_4121_p VPWR 0.0296407f $X=0.405 $Y=2.225 $X2=0 $Y2=0
cc_3148 N_A_27_297#_c_4108_n VPWR 0.0618665f $X=2.05 $Y=2.225 $X2=0 $Y2=0
cc_3149 N_A_27_297#_c_4110_n VPWR 0.0299024f $X=1.345 $Y=2.225 $X2=0 $Y2=0
cc_3150 N_A_27_297#_c_4093_n VPWR 0.0035565f $X=0.26 $Y=2.225 $X2=0 $Y2=0
cc_3151 N_A_27_297#_c_4111_n VPWR 0.00267234f $X=1.2 $Y=2.225 $X2=0 $Y2=0
cc_3152 N_A_27_297#_c_4094_n VPWR 0.0299832f $X=2.195 $Y=2.225 $X2=0 $Y2=0
cc_3153 N_A_27_297#_c_4113_n VPWR 0.00303374f $X=2.195 $Y=2.225 $X2=0 $Y2=0
cc_3154 N_A_27_297#_c_4103_n N_VPWR_c_4279_n 7.71354e-19 $X=1.055 $Y=2.225 $X2=0
+ $Y2=0
cc_3155 N_A_27_297#_c_4093_n N_VPWR_c_4279_n 0.020978f $X=0.26 $Y=2.225 $X2=0
+ $Y2=0
cc_3156 N_A_27_297#_c_4103_n N_VPWR_c_4280_n 7.64992e-19 $X=1.055 $Y=2.225 $X2=0
+ $Y2=0
cc_3157 N_A_27_297#_c_4110_n N_VPWR_c_4280_n 4.8162e-19 $X=1.345 $Y=2.225 $X2=0
+ $Y2=0
cc_3158 N_A_27_297#_c_4111_n N_VPWR_c_4280_n 0.0184771f $X=1.2 $Y=2.225 $X2=0
+ $Y2=0
cc_3159 N_A_27_297#_c_4108_n N_Z_M1013_s 0.00154628f $X=2.05 $Y=2.225 $X2=0
+ $Y2=0
cc_3160 N_A_27_297#_M1031_d N_Z_c_5242_n 0.00197114f $X=2.05 $Y=1.665 $X2=0
+ $Y2=0
cc_3161 N_A_27_297#_c_4108_n N_Z_c_5242_n 0.0225177f $X=2.05 $Y=2.225 $X2=0
+ $Y2=0
cc_3162 N_A_27_297#_c_4094_n N_Z_c_5242_n 0.0249588f $X=2.195 $Y=2.225 $X2=0
+ $Y2=0
cc_3163 N_A_27_297#_c_4113_n N_Z_c_5242_n 0.0016886f $X=2.195 $Y=2.225 $X2=0
+ $Y2=0
cc_3164 N_A_27_297#_c_4095_n N_Z_c_5242_n 0.0109134f $X=2.195 $Y=1.81 $X2=0
+ $Y2=0
cc_3165 N_A_27_297#_c_4108_n N_Z_c_5287_n 0.0241216f $X=2.05 $Y=2.225 $X2=0
+ $Y2=0
cc_3166 N_A_27_297#_c_4106_n N_Z_c_5287_n 0.0062686f $X=1.2 $Y=1.78 $X2=0 $Y2=0
cc_3167 N_A_27_297#_c_4095_n N_Z_c_5287_n 4.86317e-19 $X=2.195 $Y=1.81 $X2=0
+ $Y2=0
cc_3168 N_A_27_297#_c_4108_n N_Z_c_5288_n 0.00835547f $X=2.05 $Y=2.225 $X2=0
+ $Y2=0
cc_3169 N_A_27_297#_c_4110_n N_Z_c_5288_n 4.5829e-19 $X=1.345 $Y=2.225 $X2=0
+ $Y2=0
cc_3170 N_A_27_297#_c_4094_n N_Z_c_5288_n 4.48979e-19 $X=2.195 $Y=2.225 $X2=0
+ $Y2=0
cc_3171 N_A_27_297#_c_4106_n N_Z_c_5288_n 0.0233693f $X=1.2 $Y=1.78 $X2=0 $Y2=0
cc_3172 N_A_27_297#_c_4095_n N_Z_c_5288_n 0.0210951f $X=2.195 $Y=1.81 $X2=0
+ $Y2=0
cc_3173 N_A_27_297#_c_4099_n N_Z_c_5226_n 0.00930189f $X=1.115 $Y=1.58 $X2=0
+ $Y2=0
cc_3174 N_A_27_297#_c_4095_n N_Z_c_5226_n 0.00468052f $X=2.195 $Y=1.81 $X2=0
+ $Y2=0
cc_3175 N_A_27_297#_c_4108_n N_Z_c_5257_n 0.0115376f $X=2.05 $Y=2.225 $X2=0
+ $Y2=0
cc_3176 N_A_27_297#_c_4110_n N_Z_c_5257_n 2.82292e-19 $X=1.345 $Y=2.225 $X2=0
+ $Y2=0
cc_3177 N_A_27_297#_c_4094_n N_Z_c_5257_n 2.4892e-19 $X=2.195 $Y=2.225 $X2=0
+ $Y2=0
cc_3178 N_A_27_297#_c_4113_n N_Z_c_5257_n 0.0123065f $X=2.195 $Y=2.225 $X2=0
+ $Y2=0
cc_3179 N_A_27_297#_c_4106_n N_Z_c_5257_n 0.00347206f $X=1.2 $Y=1.78 $X2=0 $Y2=0
cc_3180 N_A_27_297#_c_4095_n N_Z_c_5257_n 0.00373869f $X=2.195 $Y=1.81 $X2=0
+ $Y2=0
cc_3181 N_A_27_297#_c_4099_n N_A_27_47#_c_7692_n 0.0110288f $X=1.115 $Y=1.58
+ $X2=0 $Y2=0
cc_3182 N_A_27_591#_c_4175_n N_VPWR_M1014_s 0.00346031f $X=1.115 $Y=3.86 $X2=0
+ $Y2=0
cc_3183 N_A_27_591#_c_4170_n N_VPWR_c_4247_n 0.00235484f $X=0.26 $Y=3.44 $X2=0
+ $Y2=0
cc_3184 N_A_27_591#_c_4186_n N_VPWR_c_4247_n 0.00995242f $X=1.2 $Y=3.14 $X2=0
+ $Y2=0
cc_3185 N_A_27_591#_c_4181_n N_VPWR_c_4247_n 0.0174313f $X=1.055 $Y=3.215 $X2=0
+ $Y2=0
cc_3186 N_A_27_591#_c_4200_p N_VPWR_c_4247_n 0.00163482f $X=0.405 $Y=3.215 $X2=0
+ $Y2=0
cc_3187 N_A_27_591#_c_4193_n N_VPWR_c_4247_n 0.00267717f $X=1.345 $Y=3.215 $X2=0
+ $Y2=0
cc_3188 N_A_27_591#_c_4183_n N_VPWR_c_4247_n 0.0254212f $X=1.2 $Y=3.215 $X2=0
+ $Y2=0
cc_3189 N_A_27_591#_c_4174_n N_VPWR_c_4247_n 0.0106781f $X=0.26 $Y=3.1 $X2=0
+ $Y2=0
cc_3190 N_A_27_591#_c_4175_n N_VPWR_c_4314_n 0.0164726f $X=1.115 $Y=3.86 $X2=0
+ $Y2=0
cc_3191 N_A_27_591#_c_4181_n N_VPWR_c_4314_n 8.54514e-19 $X=1.055 $Y=3.215 $X2=0
+ $Y2=0
cc_3192 N_A_27_591#_c_4172_n N_VPWR_c_4270_n 0.0218871f $X=2.195 $Y=3.14 $X2=0
+ $Y2=0
cc_3193 N_A_27_591#_c_4173_n N_VPWR_c_4270_n 4.78963e-19 $X=2.195 $Y=3.215 $X2=0
+ $Y2=0
cc_3194 N_A_27_591#_M1014_d VPWR 0.00111289f $X=0.135 $Y=2.955 $X2=0 $Y2=0
cc_3195 N_A_27_591#_M1078_d VPWR 0.00165645f $X=1.055 $Y=2.955 $X2=0 $Y2=0
cc_3196 N_A_27_591#_M1111_d VPWR 0.00127413f $X=2.05 $Y=2.955 $X2=0 $Y2=0
cc_3197 N_A_27_591#_c_4186_n VPWR 0.00247808f $X=1.2 $Y=3.14 $X2=0 $Y2=0
cc_3198 N_A_27_591#_c_4172_n VPWR 0.00305107f $X=2.195 $Y=3.14 $X2=0 $Y2=0
cc_3199 N_A_27_591#_c_4181_n VPWR 0.0560119f $X=1.055 $Y=3.215 $X2=0 $Y2=0
cc_3200 N_A_27_591#_c_4200_p VPWR 0.0296407f $X=0.405 $Y=3.215 $X2=0 $Y2=0
cc_3201 N_A_27_591#_c_4191_n VPWR 0.0621437f $X=2.05 $Y=3.215 $X2=0 $Y2=0
cc_3202 N_A_27_591#_c_4193_n VPWR 0.0298971f $X=1.345 $Y=3.215 $X2=0 $Y2=0
cc_3203 N_A_27_591#_c_4173_n VPWR 0.0299779f $X=2.195 $Y=3.215 $X2=0 $Y2=0
cc_3204 N_A_27_591#_c_4174_n VPWR 0.0035565f $X=0.26 $Y=3.1 $X2=0 $Y2=0
cc_3205 N_A_27_591#_c_4181_n N_VPWR_c_4279_n 7.71354e-19 $X=1.055 $Y=3.215 $X2=0
+ $Y2=0
cc_3206 N_A_27_591#_c_4174_n N_VPWR_c_4279_n 0.020978f $X=0.26 $Y=3.1 $X2=0
+ $Y2=0
cc_3207 N_A_27_591#_c_4186_n N_VPWR_c_4280_n 0.0173868f $X=1.2 $Y=3.14 $X2=0
+ $Y2=0
cc_3208 N_A_27_591#_c_4181_n N_VPWR_c_4280_n 7.64992e-19 $X=1.055 $Y=3.215 $X2=0
+ $Y2=0
cc_3209 N_A_27_591#_c_4193_n N_VPWR_c_4280_n 4.77412e-19 $X=1.345 $Y=3.215 $X2=0
+ $Y2=0
cc_3210 N_A_27_591#_c_4191_n N_Z_M1099_s 0.00154628f $X=2.05 $Y=3.215 $X2=0
+ $Y2=0
cc_3211 N_A_27_591#_c_4175_n N_Z_c_5202_n 0.00930189f $X=1.115 $Y=3.86 $X2=0
+ $Y2=0
cc_3212 N_A_27_591#_c_4172_n N_Z_c_5202_n 0.00468052f $X=2.195 $Y=3.14 $X2=0
+ $Y2=0
cc_3213 N_A_27_591#_M1111_d N_Z_c_5243_n 0.00197114f $X=2.05 $Y=2.955 $X2=0
+ $Y2=0
cc_3214 N_A_27_591#_c_4172_n N_Z_c_5243_n 0.0126134f $X=2.195 $Y=3.14 $X2=0
+ $Y2=0
cc_3215 N_A_27_591#_c_4191_n N_Z_c_5243_n 0.0225176f $X=2.05 $Y=3.215 $X2=0
+ $Y2=0
cc_3216 N_A_27_591#_c_4173_n N_Z_c_5243_n 0.0249588f $X=2.195 $Y=3.215 $X2=0
+ $Y2=0
cc_3217 N_A_27_591#_c_4172_n N_Z_c_5313_n 4.86317e-19 $X=2.195 $Y=3.14 $X2=0
+ $Y2=0
cc_3218 N_A_27_591#_c_4191_n N_Z_c_5313_n 0.0241216f $X=2.05 $Y=3.215 $X2=0
+ $Y2=0
cc_3219 N_A_27_591#_c_4183_n N_Z_c_5313_n 0.0062686f $X=1.2 $Y=3.215 $X2=0 $Y2=0
cc_3220 N_A_27_591#_c_4172_n N_Z_c_5297_n 0.0210951f $X=2.195 $Y=3.14 $X2=0
+ $Y2=0
cc_3221 N_A_27_591#_c_4191_n N_Z_c_5297_n 0.00835547f $X=2.05 $Y=3.215 $X2=0
+ $Y2=0
cc_3222 N_A_27_591#_c_4193_n N_Z_c_5297_n 4.5829e-19 $X=1.345 $Y=3.215 $X2=0
+ $Y2=0
cc_3223 N_A_27_591#_c_4183_n N_Z_c_5297_n 0.0233693f $X=1.2 $Y=3.215 $X2=0 $Y2=0
cc_3224 N_A_27_591#_c_4173_n N_Z_c_5297_n 4.48979e-19 $X=2.195 $Y=3.215 $X2=0
+ $Y2=0
cc_3225 N_A_27_591#_c_4172_n N_Z_c_5257_n 0.0161129f $X=2.195 $Y=3.14 $X2=0
+ $Y2=0
cc_3226 N_A_27_591#_c_4191_n N_Z_c_5257_n 0.0115376f $X=2.05 $Y=3.215 $X2=0
+ $Y2=0
cc_3227 N_A_27_591#_c_4193_n N_Z_c_5257_n 2.75404e-19 $X=1.345 $Y=3.215 $X2=0
+ $Y2=0
cc_3228 N_A_27_591#_c_4183_n N_Z_c_5257_n 0.00349107f $X=1.2 $Y=3.215 $X2=0
+ $Y2=0
cc_3229 N_A_27_591#_c_4173_n N_Z_c_5257_n 2.48349e-19 $X=2.195 $Y=3.215 $X2=0
+ $Y2=0
cc_3230 N_A_27_591#_c_4175_n N_A_27_911#_c_7737_n 0.00251701f $X=1.115 $Y=3.86
+ $X2=0 $Y2=0
cc_3231 N_A_27_591#_c_4175_n N_A_27_911#_c_7734_n 0.00851176f $X=1.115 $Y=3.86
+ $X2=0 $Y2=0
cc_3232 VPWR N_Z_M1013_s 6.43831e-19 $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3233 VPWR N_Z_M1099_s 6.43831e-19 $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3234 VPWR N_Z_M1084_s 6.43831e-19 $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3235 VPWR N_Z_M1036_d 6.43831e-19 $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3236 VPWR N_Z_M1005_d 6.43831e-19 $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3237 VPWR N_Z_M1044_s 6.43831e-19 $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3238 VPWR N_Z_M1004_d 6.43831e-19 $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3239 VPWR N_Z_M1045_s 6.43831e-19 $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3240 VPWR N_Z_M1034_s 6.43831e-19 $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3241 VPWR N_Z_M1114_s 6.43831e-19 $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3242 VPWR N_Z_M1055_s 6.43831e-19 $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3243 VPWR N_Z_M1134_s 6.43831e-19 $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3244 VPWR N_Z_M1066_s 6.43831e-19 $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3245 VPWR N_Z_M1006_d 6.43831e-19 $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3246 VPWR N_Z_M1122_s 6.43831e-19 $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3247 VPWR N_Z_M1049_s 6.43831e-19 $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3248 N_VPWR_M1023_d N_Z_c_5242_n 5.82057e-19 $X=3.04 $Y=1.485 $X2=0 $Y2=0
cc_3249 N_VPWR_c_4248_n N_Z_c_5242_n 0.0287846f $X=3.22 $Y=1.63 $X2=0 $Y2=0
cc_3250 VPWR N_Z_c_5242_n 0.083114f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3251 N_VPWR_M1027_d N_Z_c_5243_n 5.82057e-19 $X=3.04 $Y=2.955 $X2=0 $Y2=0
cc_3252 N_VPWR_c_4249_n N_Z_c_5243_n 0.0287846f $X=3.22 $Y=3.13 $X2=0 $Y2=0
cc_3253 VPWR N_Z_c_5243_n 0.083114f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3254 N_VPWR_M1052_s N_Z_c_5244_n 0.00219731f $X=5.565 $Y=1.485 $X2=0 $Y2=0
cc_3255 N_VPWR_M1003_d N_Z_c_5244_n 0.00219731f $X=7.025 $Y=1.485 $X2=0 $Y2=0
cc_3256 N_VPWR_c_4376_n N_Z_c_5244_n 0.0121265f $X=5.71 $Y=1.94 $X2=0 $Y2=0
cc_3257 N_VPWR_c_4392_n N_Z_c_5244_n 0.0121265f $X=7.17 $Y=1.94 $X2=0 $Y2=0
cc_3258 VPWR N_Z_c_5244_n 0.0120388f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3259 N_VPWR_M1056_s N_Z_c_5245_n 0.00219731f $X=5.565 $Y=2.955 $X2=0 $Y2=0
cc_3260 N_VPWR_M1009_d N_Z_c_5245_n 0.00219731f $X=7.025 $Y=2.955 $X2=0 $Y2=0
cc_3261 N_VPWR_c_4384_n N_Z_c_5245_n 0.012122f $X=5.71 $Y=3.5 $X2=0 $Y2=0
cc_3262 N_VPWR_c_4400_n N_Z_c_5245_n 0.0121243f $X=7.17 $Y=3.5 $X2=0 $Y2=0
cc_3263 VPWR N_Z_c_5245_n 0.0120388f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3264 N_VPWR_M1133_d N_Z_c_5246_n 5.82057e-19 $X=9.48 $Y=1.485 $X2=0 $Y2=0
cc_3265 N_VPWR_c_4254_n N_Z_c_5246_n 0.0287846f $X=9.66 $Y=1.63 $X2=0 $Y2=0
cc_3266 VPWR N_Z_c_5246_n 0.083114f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3267 N_VPWR_M1137_d N_Z_c_5247_n 5.82057e-19 $X=9.48 $Y=2.955 $X2=0 $Y2=0
cc_3268 N_VPWR_c_4255_n N_Z_c_5247_n 0.0287846f $X=9.66 $Y=3.13 $X2=0 $Y2=0
cc_3269 VPWR N_Z_c_5247_n 0.083114f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3270 N_VPWR_M1002_d N_Z_c_5248_n 0.00219731f $X=12.005 $Y=1.485 $X2=0 $Y2=0
cc_3271 N_VPWR_M1030_s N_Z_c_5248_n 0.00219731f $X=13.465 $Y=1.485 $X2=0 $Y2=0
cc_3272 N_VPWR_c_4462_n N_Z_c_5248_n 0.0121265f $X=12.15 $Y=1.94 $X2=0 $Y2=0
cc_3273 N_VPWR_c_4478_n N_Z_c_5248_n 0.0121265f $X=13.61 $Y=1.94 $X2=0 $Y2=0
cc_3274 VPWR N_Z_c_5248_n 0.0120388f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3275 N_VPWR_M1008_d N_Z_c_5249_n 0.00219731f $X=12.005 $Y=2.955 $X2=0 $Y2=0
cc_3276 N_VPWR_M1038_s N_Z_c_5249_n 0.00219731f $X=13.465 $Y=2.955 $X2=0 $Y2=0
cc_3277 N_VPWR_c_4470_n N_Z_c_5249_n 0.012122f $X=12.15 $Y=3.5 $X2=0 $Y2=0
cc_3278 N_VPWR_c_4486_n N_Z_c_5249_n 0.0121243f $X=13.61 $Y=3.5 $X2=0 $Y2=0
cc_3279 VPWR N_Z_c_5249_n 0.0120388f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3280 N_VPWR_M1001_d N_Z_c_5250_n 5.82057e-19 $X=15.92 $Y=1.485 $X2=0 $Y2=0
cc_3281 N_VPWR_c_4260_n N_Z_c_5250_n 0.0287846f $X=16.1 $Y=1.63 $X2=0 $Y2=0
cc_3282 VPWR N_Z_c_5250_n 0.083114f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3283 N_VPWR_M1007_d N_Z_c_5251_n 5.82057e-19 $X=15.92 $Y=2.955 $X2=0 $Y2=0
cc_3284 N_VPWR_c_4261_n N_Z_c_5251_n 0.0287846f $X=16.1 $Y=3.13 $X2=0 $Y2=0
cc_3285 VPWR N_Z_c_5251_n 0.083114f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3286 N_VPWR_M1051_s N_Z_c_5252_n 0.00219731f $X=18.445 $Y=1.485 $X2=0 $Y2=0
cc_3287 N_VPWR_M1062_s N_Z_c_5252_n 0.00219731f $X=19.905 $Y=1.485 $X2=0 $Y2=0
cc_3288 N_VPWR_c_4548_n N_Z_c_5252_n 0.0121265f $X=18.59 $Y=1.94 $X2=0 $Y2=0
cc_3289 N_VPWR_c_4564_n N_Z_c_5252_n 0.0121265f $X=20.05 $Y=1.94 $X2=0 $Y2=0
cc_3290 VPWR N_Z_c_5252_n 0.0120388f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3291 N_VPWR_M1058_s N_Z_c_5253_n 0.00219731f $X=18.445 $Y=2.955 $X2=0 $Y2=0
cc_3292 N_VPWR_M1069_s N_Z_c_5253_n 0.00219731f $X=19.905 $Y=2.955 $X2=0 $Y2=0
cc_3293 N_VPWR_c_4556_n N_Z_c_5253_n 0.012122f $X=18.59 $Y=3.5 $X2=0 $Y2=0
cc_3294 N_VPWR_c_4572_n N_Z_c_5253_n 0.0121243f $X=20.05 $Y=3.5 $X2=0 $Y2=0
cc_3295 VPWR N_Z_c_5253_n 0.0120388f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3296 N_VPWR_M1077_d N_Z_c_5254_n 5.82057e-19 $X=22.36 $Y=1.485 $X2=0 $Y2=0
cc_3297 N_VPWR_c_4266_n N_Z_c_5254_n 0.0287846f $X=22.54 $Y=1.63 $X2=0 $Y2=0
cc_3298 VPWR N_Z_c_5254_n 0.083114f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3299 N_VPWR_M1085_d N_Z_c_5255_n 5.82057e-19 $X=22.36 $Y=2.955 $X2=0 $Y2=0
cc_3300 N_VPWR_c_4267_n N_Z_c_5255_n 0.0287846f $X=22.54 $Y=3.13 $X2=0 $Y2=0
cc_3301 VPWR N_Z_c_5255_n 0.083114f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3302 N_VPWR_c_4270_n N_Z_c_5257_n 0.0121875f $X=3.055 $Y=2.72 $X2=0 $Y2=0
cc_3303 VPWR N_Z_c_5257_n 0.0388938f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3304 N_VPWR_c_4280_n N_Z_c_5257_n 0.0121875f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_3305 VPWR N_Z_c_5259_n 0.0388938f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3306 N_VPWR_c_4281_n N_Z_c_5259_n 0.0121875f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_3307 N_VPWR_c_4282_n N_Z_c_5259_n 0.0121875f $X=5.545 $Y=2.72 $X2=0 $Y2=0
cc_3308 N_VPWR_c_4272_n N_Z_c_5261_n 0.0121875f $X=9.495 $Y=2.72 $X2=0 $Y2=0
cc_3309 VPWR N_Z_c_5261_n 0.0388938f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3310 N_VPWR_c_4284_n N_Z_c_5261_n 0.0121875f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_3311 VPWR N_Z_c_5263_n 0.0388938f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3312 N_VPWR_c_4285_n N_Z_c_5263_n 0.0121875f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_3313 N_VPWR_c_4286_n N_Z_c_5263_n 0.0121875f $X=11.985 $Y=2.72 $X2=0 $Y2=0
cc_3314 N_VPWR_c_4274_n N_Z_c_5265_n 0.0121875f $X=15.935 $Y=2.72 $X2=0 $Y2=0
cc_3315 VPWR N_Z_c_5265_n 0.0388938f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3316 N_VPWR_c_4288_n N_Z_c_5265_n 0.0121875f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_3317 VPWR N_Z_c_5267_n 0.0388938f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3318 N_VPWR_c_4289_n N_Z_c_5267_n 0.0121875f $X=17.25 $Y=2.72 $X2=0 $Y2=0
cc_3319 N_VPWR_c_4290_n N_Z_c_5267_n 0.0121875f $X=18.425 $Y=2.72 $X2=0 $Y2=0
cc_3320 N_VPWR_c_4276_n N_Z_c_5269_n 0.0121875f $X=22.375 $Y=2.72 $X2=0 $Y2=0
cc_3321 VPWR N_Z_c_5269_n 0.0388938f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3322 N_VPWR_c_4292_n N_Z_c_5269_n 0.0121875f $X=20.47 $Y=2.72 $X2=0 $Y2=0
cc_3323 VPWR N_Z_c_5271_n 0.0388938f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3324 N_VPWR_c_4293_n N_Z_c_5271_n 0.0121875f $X=23.69 $Y=2.72 $X2=0 $Y2=0
cc_3325 N_VPWR_c_4294_n N_Z_c_5271_n 0.0121875f $X=24.865 $Y=2.72 $X2=0 $Y2=0
cc_3326 VPWR N_A_824_333#_M1084_d 0.00127816f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=1.305
cc_3327 VPWR N_A_824_333#_M1113_d 0.00166446f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3328 VPWR N_A_824_333#_M1097_d 0.00111289f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3329 N_VPWR_M1052_s N_A_824_333#_c_6435_n 0.00331615f $X=5.565 $Y=1.485 $X2=0
+ $Y2=0
cc_3330 N_VPWR_c_4376_n N_A_824_333#_c_6435_n 0.0158304f $X=5.71 $Y=1.94 $X2=0
+ $Y2=0
cc_3331 VPWR N_A_824_333#_c_6424_n 0.0618665f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3332 VPWR N_A_824_333#_c_6419_n 0.0299832f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3333 N_VPWR_c_4281_n N_A_824_333#_c_6419_n 4.83649e-19 $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_3334 N_VPWR_c_4250_n N_A_824_333#_c_6441_n 0.0170179f $X=5.71 $Y=2.34 $X2=0
+ $Y2=0
cc_3335 N_VPWR_c_4376_n N_A_824_333#_c_6441_n 3.68476e-19 $X=5.71 $Y=1.94 $X2=0
+ $Y2=0
cc_3336 VPWR N_A_824_333#_c_6441_n 0.0560119f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3337 N_VPWR_c_4282_n N_A_824_333#_c_6441_n 7.64992e-19 $X=5.545 $Y=2.72 $X2=0
+ $Y2=0
cc_3338 N_VPWR_c_4283_n N_A_824_333#_c_6441_n 7.71354e-19 $X=7.035 $Y=2.72 $X2=0
+ $Y2=0
cc_3339 N_VPWR_c_4250_n N_A_824_333#_c_6427_n 0.00265921f $X=5.71 $Y=2.34 $X2=0
+ $Y2=0
cc_3340 VPWR N_A_824_333#_c_6427_n 0.0299024f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3341 N_VPWR_c_4282_n N_A_824_333#_c_6427_n 4.8162e-19 $X=5.545 $Y=2.72 $X2=0
+ $Y2=0
cc_3342 VPWR N_A_824_333#_c_6428_n 0.00303374f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3343 N_VPWR_c_4281_n N_A_824_333#_c_6428_n 0.0217548f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_3344 N_VPWR_c_4250_n N_A_824_333#_c_6429_n 0.0173701f $X=5.71 $Y=2.34 $X2=0
+ $Y2=0
cc_3345 VPWR N_A_824_333#_c_6429_n 0.00267234f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3346 N_VPWR_c_4282_n N_A_824_333#_c_6429_n 0.0184771f $X=5.545 $Y=2.72 $X2=0
+ $Y2=0
cc_3347 N_VPWR_c_4250_n N_A_824_333#_c_6466_n 0.00163482f $X=5.71 $Y=2.34 $X2=0
+ $Y2=0
cc_3348 VPWR N_A_824_333#_c_6466_n 0.0296407f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3349 N_VPWR_c_4250_n N_A_824_333#_c_6420_n 0.0106781f $X=5.71 $Y=2.34 $X2=0
+ $Y2=0
cc_3350 VPWR N_A_824_333#_c_6420_n 0.00317333f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3351 N_VPWR_c_4283_n N_A_824_333#_c_6420_n 0.020978f $X=7.035 $Y=2.72 $X2=0
+ $Y2=0
cc_3352 N_VPWR_c_4376_n N_A_824_333#_c_6434_n 0.0173701f $X=5.71 $Y=1.94 $X2=0
+ $Y2=0
cc_3353 N_VPWR_c_4250_n N_A_824_333#_c_6422_n 0.00235484f $X=5.71 $Y=2.34 $X2=0
+ $Y2=0
cc_3354 N_VPWR_c_4376_n N_A_824_333#_c_6422_n 0.0115021f $X=5.71 $Y=1.94 $X2=0
+ $Y2=0
cc_3355 VPWR N_A_824_591#_M1036_s 0.00127413f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=1.305
cc_3356 VPWR N_A_824_591#_M1157_s 0.00165645f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3357 VPWR N_A_824_591#_M1101_d 0.00111289f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3358 N_VPWR_M1056_s N_A_824_591#_c_6514_n 0.00331615f $X=5.565 $Y=2.955 $X2=0
+ $Y2=0
cc_3359 N_VPWR_c_4384_n N_A_824_591#_c_6514_n 0.015867f $X=5.71 $Y=3.5 $X2=0
+ $Y2=0
cc_3360 N_VPWR_c_4251_n N_A_824_591#_c_6515_n 0.00235484f $X=5.71 $Y=3.1 $X2=0
+ $Y2=0
cc_3361 N_VPWR_c_4384_n N_A_824_591#_c_6515_n 0.0115021f $X=5.71 $Y=3.5 $X2=0
+ $Y2=0
cc_3362 VPWR N_A_824_591#_c_6516_n 0.00305107f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3363 N_VPWR_c_4281_n N_A_824_591#_c_6516_n 0.0218871f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_3364 N_VPWR_c_4251_n N_A_824_591#_c_6524_n 0.00995242f $X=5.71 $Y=3.1 $X2=0
+ $Y2=0
cc_3365 VPWR N_A_824_591#_c_6524_n 0.00247808f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3366 N_VPWR_c_4282_n N_A_824_591#_c_6524_n 0.0173868f $X=5.545 $Y=2.72 $X2=0
+ $Y2=0
cc_3367 VPWR N_A_824_591#_c_6525_n 0.0621437f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3368 VPWR N_A_824_591#_c_6517_n 0.0299779f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3369 N_VPWR_c_4281_n N_A_824_591#_c_6517_n 4.78963e-19 $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_3370 N_VPWR_c_4251_n N_A_824_591#_c_6534_n 0.0170179f $X=5.71 $Y=3.1 $X2=0
+ $Y2=0
cc_3371 N_VPWR_c_4384_n N_A_824_591#_c_6534_n 3.57652e-19 $X=5.71 $Y=3.5 $X2=0
+ $Y2=0
cc_3372 VPWR N_A_824_591#_c_6534_n 0.0560119f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3373 N_VPWR_c_4282_n N_A_824_591#_c_6534_n 7.64992e-19 $X=5.545 $Y=2.72 $X2=0
+ $Y2=0
cc_3374 N_VPWR_c_4283_n N_A_824_591#_c_6534_n 7.71354e-19 $X=7.035 $Y=2.72 $X2=0
+ $Y2=0
cc_3375 N_VPWR_c_4251_n N_A_824_591#_c_6528_n 0.00267717f $X=5.71 $Y=3.1 $X2=0
+ $Y2=0
cc_3376 VPWR N_A_824_591#_c_6528_n 0.0298971f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3377 N_VPWR_c_4282_n N_A_824_591#_c_6528_n 4.77412e-19 $X=5.545 $Y=2.72 $X2=0
+ $Y2=0
cc_3378 N_VPWR_c_4251_n N_A_824_591#_c_6529_n 0.0247455f $X=5.71 $Y=3.1 $X2=0
+ $Y2=0
cc_3379 N_VPWR_c_4251_n N_A_824_591#_c_6562_n 0.00163482f $X=5.71 $Y=3.1 $X2=0
+ $Y2=0
cc_3380 VPWR N_A_824_591#_c_6562_n 0.0296407f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3381 N_VPWR_c_4251_n N_A_824_591#_c_6518_n 0.0106781f $X=5.71 $Y=3.1 $X2=0
+ $Y2=0
cc_3382 VPWR N_A_824_591#_c_6518_n 0.00317333f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3383 N_VPWR_c_4283_n N_A_824_591#_c_6518_n 0.020978f $X=7.035 $Y=2.72 $X2=0
+ $Y2=0
cc_3384 VPWR N_A_1315_297#_M1003_s 0.00111289f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=1.305
cc_3385 VPWR N_A_1315_297#_M1120_s 0.00166446f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3386 VPWR N_A_1315_297#_M1124_s 0.00127816f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3387 N_VPWR_M1003_d N_A_1315_297#_c_6612_n 0.00331615f $X=7.025 $Y=1.485
+ $X2=0 $Y2=0
cc_3388 N_VPWR_c_4392_n N_A_1315_297#_c_6612_n 0.0158304f $X=7.17 $Y=1.94 $X2=0
+ $Y2=0
cc_3389 N_VPWR_c_4252_n N_A_1315_297#_c_6616_n 0.0170179f $X=7.17 $Y=2.34 $X2=0
+ $Y2=0
cc_3390 N_VPWR_c_4392_n N_A_1315_297#_c_6616_n 3.68476e-19 $X=7.17 $Y=1.94 $X2=0
+ $Y2=0
cc_3391 VPWR N_A_1315_297#_c_6616_n 0.0560119f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3392 N_VPWR_c_4283_n N_A_1315_297#_c_6616_n 7.71354e-19 $X=7.035 $Y=2.72
+ $X2=0 $Y2=0
cc_3393 N_VPWR_c_4284_n N_A_1315_297#_c_6616_n 7.64992e-19 $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_3394 N_VPWR_c_4252_n N_A_1315_297#_c_6642_n 0.00163482f $X=7.17 $Y=2.34 $X2=0
+ $Y2=0
cc_3395 VPWR N_A_1315_297#_c_6642_n 0.0296407f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3396 VPWR N_A_1315_297#_c_6621_n 0.0618665f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3397 N_VPWR_c_4252_n N_A_1315_297#_c_6623_n 0.00265921f $X=7.17 $Y=2.34 $X2=0
+ $Y2=0
cc_3398 VPWR N_A_1315_297#_c_6623_n 0.0299024f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3399 N_VPWR_c_4284_n N_A_1315_297#_c_6623_n 4.8162e-19 $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_3400 N_VPWR_c_4252_n N_A_1315_297#_c_6606_n 0.0106781f $X=7.17 $Y=2.34 $X2=0
+ $Y2=0
cc_3401 VPWR N_A_1315_297#_c_6606_n 0.00317333f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3402 N_VPWR_c_4283_n N_A_1315_297#_c_6606_n 0.020978f $X=7.035 $Y=2.72 $X2=0
+ $Y2=0
cc_3403 N_VPWR_c_4252_n N_A_1315_297#_c_6624_n 0.0173701f $X=7.17 $Y=2.34 $X2=0
+ $Y2=0
cc_3404 VPWR N_A_1315_297#_c_6624_n 0.00267234f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3405 N_VPWR_c_4284_n N_A_1315_297#_c_6624_n 0.0184771f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_3406 N_VPWR_c_4272_n N_A_1315_297#_c_6607_n 4.83649e-19 $X=9.495 $Y=2.72
+ $X2=0 $Y2=0
cc_3407 VPWR N_A_1315_297#_c_6607_n 0.0299832f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3408 N_VPWR_c_4272_n N_A_1315_297#_c_6626_n 0.0217548f $X=9.495 $Y=2.72 $X2=0
+ $Y2=0
cc_3409 VPWR N_A_1315_297#_c_6626_n 0.00303374f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3410 N_VPWR_c_4392_n N_A_1315_297#_c_6619_n 0.0173701f $X=7.17 $Y=1.94 $X2=0
+ $Y2=0
cc_3411 N_VPWR_c_4252_n N_A_1315_297#_c_6609_n 0.00235484f $X=7.17 $Y=2.34 $X2=0
+ $Y2=0
cc_3412 N_VPWR_c_4392_n N_A_1315_297#_c_6609_n 0.0115021f $X=7.17 $Y=1.94 $X2=0
+ $Y2=0
cc_3413 VPWR N_A_1315_591#_M1009_s 0.00111289f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=1.305
cc_3414 VPWR N_A_1315_591#_M1126_s 0.00165645f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3415 VPWR N_A_1315_591#_M1095_d 0.00127413f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3416 N_VPWR_c_4253_n N_A_1315_591#_c_6699_n 0.00235484f $X=7.17 $Y=3.1 $X2=0
+ $Y2=0
cc_3417 N_VPWR_c_4400_n N_A_1315_591#_c_6699_n 0.0115021f $X=7.17 $Y=3.5 $X2=0
+ $Y2=0
cc_3418 N_VPWR_M1009_d N_A_1315_591#_c_6704_n 0.00331615f $X=7.025 $Y=2.955
+ $X2=0 $Y2=0
cc_3419 N_VPWR_c_4400_n N_A_1315_591#_c_6704_n 0.0158304f $X=7.17 $Y=3.5 $X2=0
+ $Y2=0
cc_3420 N_VPWR_c_4253_n N_A_1315_591#_c_6715_n 0.00995242f $X=7.17 $Y=3.1 $X2=0
+ $Y2=0
cc_3421 VPWR N_A_1315_591#_c_6715_n 0.00247808f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3422 N_VPWR_c_4284_n N_A_1315_591#_c_6715_n 0.0173868f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_3423 N_VPWR_c_4272_n N_A_1315_591#_c_6701_n 0.0218871f $X=9.495 $Y=2.72 $X2=0
+ $Y2=0
cc_3424 VPWR N_A_1315_591#_c_6701_n 0.00305107f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3425 N_VPWR_c_4253_n N_A_1315_591#_c_6710_n 0.0170179f $X=7.17 $Y=3.1 $X2=0
+ $Y2=0
cc_3426 N_VPWR_c_4400_n N_A_1315_591#_c_6710_n 3.68476e-19 $X=7.17 $Y=3.5 $X2=0
+ $Y2=0
cc_3427 VPWR N_A_1315_591#_c_6710_n 0.0560119f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3428 N_VPWR_c_4283_n N_A_1315_591#_c_6710_n 7.71354e-19 $X=7.035 $Y=2.72
+ $X2=0 $Y2=0
cc_3429 N_VPWR_c_4284_n N_A_1315_591#_c_6710_n 7.64992e-19 $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_3430 N_VPWR_c_4253_n N_A_1315_591#_c_6742_n 0.00163482f $X=7.17 $Y=3.1 $X2=0
+ $Y2=0
cc_3431 VPWR N_A_1315_591#_c_6742_n 0.0296407f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3432 VPWR N_A_1315_591#_c_6720_n 0.0621437f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3433 N_VPWR_c_4253_n N_A_1315_591#_c_6722_n 0.00267717f $X=7.17 $Y=3.1 $X2=0
+ $Y2=0
cc_3434 VPWR N_A_1315_591#_c_6722_n 0.0298971f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3435 N_VPWR_c_4284_n N_A_1315_591#_c_6722_n 4.77412e-19 $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_3436 N_VPWR_c_4253_n N_A_1315_591#_c_6712_n 0.0247455f $X=7.17 $Y=3.1 $X2=0
+ $Y2=0
cc_3437 N_VPWR_c_4272_n N_A_1315_591#_c_6702_n 4.78963e-19 $X=9.495 $Y=2.72
+ $X2=0 $Y2=0
cc_3438 VPWR N_A_1315_591#_c_6702_n 0.0299779f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3439 N_VPWR_c_4253_n N_A_1315_591#_c_6703_n 0.0106781f $X=7.17 $Y=3.1 $X2=0
+ $Y2=0
cc_3440 VPWR N_A_1315_591#_c_6703_n 0.00317333f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3441 N_VPWR_c_4283_n N_A_1315_591#_c_6703_n 0.020978f $X=7.035 $Y=2.72 $X2=0
+ $Y2=0
cc_3442 VPWR N_A_2112_333#_M1004_s 0.00127816f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=1.305
cc_3443 VPWR N_A_2112_333#_M1123_s 0.00166446f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3444 VPWR N_A_2112_333#_M1135_s 0.00111289f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3445 N_VPWR_M1002_d N_A_2112_333#_c_6808_n 0.00331615f $X=12.005 $Y=1.485
+ $X2=0 $Y2=0
cc_3446 N_VPWR_c_4462_n N_A_2112_333#_c_6808_n 0.0158304f $X=12.15 $Y=1.94 $X2=0
+ $Y2=0
cc_3447 VPWR N_A_2112_333#_c_6797_n 0.0618665f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3448 VPWR N_A_2112_333#_c_6792_n 0.0299832f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3449 N_VPWR_c_4285_n N_A_2112_333#_c_6792_n 4.83649e-19 $X=10.81 $Y=2.72
+ $X2=0 $Y2=0
cc_3450 N_VPWR_c_4256_n N_A_2112_333#_c_6814_n 0.0170179f $X=12.15 $Y=2.34 $X2=0
+ $Y2=0
cc_3451 N_VPWR_c_4462_n N_A_2112_333#_c_6814_n 3.68476e-19 $X=12.15 $Y=1.94
+ $X2=0 $Y2=0
cc_3452 VPWR N_A_2112_333#_c_6814_n 0.0560119f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3453 N_VPWR_c_4286_n N_A_2112_333#_c_6814_n 7.64992e-19 $X=11.985 $Y=2.72
+ $X2=0 $Y2=0
cc_3454 N_VPWR_c_4287_n N_A_2112_333#_c_6814_n 7.71354e-19 $X=13.475 $Y=2.72
+ $X2=0 $Y2=0
cc_3455 N_VPWR_c_4256_n N_A_2112_333#_c_6800_n 0.00265921f $X=12.15 $Y=2.34
+ $X2=0 $Y2=0
cc_3456 VPWR N_A_2112_333#_c_6800_n 0.0299024f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3457 N_VPWR_c_4286_n N_A_2112_333#_c_6800_n 4.8162e-19 $X=11.985 $Y=2.72
+ $X2=0 $Y2=0
cc_3458 VPWR N_A_2112_333#_c_6801_n 0.00303374f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3459 N_VPWR_c_4285_n N_A_2112_333#_c_6801_n 0.0217548f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_3460 N_VPWR_c_4256_n N_A_2112_333#_c_6802_n 0.0173701f $X=12.15 $Y=2.34 $X2=0
+ $Y2=0
cc_3461 VPWR N_A_2112_333#_c_6802_n 0.00267234f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3462 N_VPWR_c_4286_n N_A_2112_333#_c_6802_n 0.0184771f $X=11.985 $Y=2.72
+ $X2=0 $Y2=0
cc_3463 N_VPWR_c_4256_n N_A_2112_333#_c_6839_n 0.00163482f $X=12.15 $Y=2.34
+ $X2=0 $Y2=0
cc_3464 VPWR N_A_2112_333#_c_6839_n 0.0296407f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3465 N_VPWR_c_4256_n N_A_2112_333#_c_6793_n 0.0106781f $X=12.15 $Y=2.34 $X2=0
+ $Y2=0
cc_3466 VPWR N_A_2112_333#_c_6793_n 0.00317333f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3467 N_VPWR_c_4287_n N_A_2112_333#_c_6793_n 0.020978f $X=13.475 $Y=2.72 $X2=0
+ $Y2=0
cc_3468 N_VPWR_c_4462_n N_A_2112_333#_c_6807_n 0.0173701f $X=12.15 $Y=1.94 $X2=0
+ $Y2=0
cc_3469 N_VPWR_c_4256_n N_A_2112_333#_c_6795_n 0.00235484f $X=12.15 $Y=2.34
+ $X2=0 $Y2=0
cc_3470 N_VPWR_c_4462_n N_A_2112_333#_c_6795_n 0.0115021f $X=12.15 $Y=1.94 $X2=0
+ $Y2=0
cc_3471 VPWR N_A_2112_591#_M1045_d 0.00127413f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=1.305
cc_3472 VPWR N_A_2112_591#_M1093_d 0.00165645f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3473 VPWR N_A_2112_591#_M1141_s 0.00111289f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3474 N_VPWR_M1008_d N_A_2112_591#_c_6887_n 0.00331615f $X=12.005 $Y=2.955
+ $X2=0 $Y2=0
cc_3475 N_VPWR_c_4470_n N_A_2112_591#_c_6887_n 0.015867f $X=12.15 $Y=3.5 $X2=0
+ $Y2=0
cc_3476 N_VPWR_c_4257_n N_A_2112_591#_c_6888_n 0.00235484f $X=12.15 $Y=3.1 $X2=0
+ $Y2=0
cc_3477 N_VPWR_c_4470_n N_A_2112_591#_c_6888_n 0.0115021f $X=12.15 $Y=3.5 $X2=0
+ $Y2=0
cc_3478 VPWR N_A_2112_591#_c_6889_n 0.00305107f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3479 N_VPWR_c_4285_n N_A_2112_591#_c_6889_n 0.0218871f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_3480 N_VPWR_c_4257_n N_A_2112_591#_c_6897_n 0.00995242f $X=12.15 $Y=3.1 $X2=0
+ $Y2=0
cc_3481 VPWR N_A_2112_591#_c_6897_n 0.00247808f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3482 N_VPWR_c_4286_n N_A_2112_591#_c_6897_n 0.0173868f $X=11.985 $Y=2.72
+ $X2=0 $Y2=0
cc_3483 VPWR N_A_2112_591#_c_6898_n 0.0621437f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3484 VPWR N_A_2112_591#_c_6890_n 0.0299779f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3485 N_VPWR_c_4285_n N_A_2112_591#_c_6890_n 4.78963e-19 $X=10.81 $Y=2.72
+ $X2=0 $Y2=0
cc_3486 N_VPWR_c_4257_n N_A_2112_591#_c_6907_n 0.0170179f $X=12.15 $Y=3.1 $X2=0
+ $Y2=0
cc_3487 N_VPWR_c_4470_n N_A_2112_591#_c_6907_n 3.57652e-19 $X=12.15 $Y=3.5 $X2=0
+ $Y2=0
cc_3488 VPWR N_A_2112_591#_c_6907_n 0.0560119f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3489 N_VPWR_c_4286_n N_A_2112_591#_c_6907_n 7.64992e-19 $X=11.985 $Y=2.72
+ $X2=0 $Y2=0
cc_3490 N_VPWR_c_4287_n N_A_2112_591#_c_6907_n 7.71354e-19 $X=13.475 $Y=2.72
+ $X2=0 $Y2=0
cc_3491 N_VPWR_c_4257_n N_A_2112_591#_c_6901_n 0.00267717f $X=12.15 $Y=3.1 $X2=0
+ $Y2=0
cc_3492 VPWR N_A_2112_591#_c_6901_n 0.0298971f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3493 N_VPWR_c_4286_n N_A_2112_591#_c_6901_n 4.77412e-19 $X=11.985 $Y=2.72
+ $X2=0 $Y2=0
cc_3494 N_VPWR_c_4257_n N_A_2112_591#_c_6902_n 0.0247455f $X=12.15 $Y=3.1 $X2=0
+ $Y2=0
cc_3495 N_VPWR_c_4257_n N_A_2112_591#_c_6935_n 0.00163482f $X=12.15 $Y=3.1 $X2=0
+ $Y2=0
cc_3496 VPWR N_A_2112_591#_c_6935_n 0.0296407f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3497 N_VPWR_c_4257_n N_A_2112_591#_c_6891_n 0.0106781f $X=12.15 $Y=3.1 $X2=0
+ $Y2=0
cc_3498 VPWR N_A_2112_591#_c_6891_n 0.00317333f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3499 N_VPWR_c_4287_n N_A_2112_591#_c_6891_n 0.020978f $X=13.475 $Y=2.72 $X2=0
+ $Y2=0
cc_3500 VPWR N_A_2603_297#_M1030_d 0.00111289f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=1.305
cc_3501 VPWR N_A_2603_297#_M1080_d 0.00166446f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3502 VPWR N_A_2603_297#_M1083_d 0.00127816f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3503 N_VPWR_M1030_s N_A_2603_297#_c_6985_n 0.00331615f $X=13.465 $Y=1.485
+ $X2=0 $Y2=0
cc_3504 N_VPWR_c_4478_n N_A_2603_297#_c_6985_n 0.0158304f $X=13.61 $Y=1.94 $X2=0
+ $Y2=0
cc_3505 N_VPWR_c_4258_n N_A_2603_297#_c_6989_n 0.0170179f $X=13.61 $Y=2.34 $X2=0
+ $Y2=0
cc_3506 N_VPWR_c_4478_n N_A_2603_297#_c_6989_n 3.68476e-19 $X=13.61 $Y=1.94
+ $X2=0 $Y2=0
cc_3507 VPWR N_A_2603_297#_c_6989_n 0.0560119f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3508 N_VPWR_c_4287_n N_A_2603_297#_c_6989_n 7.71354e-19 $X=13.475 $Y=2.72
+ $X2=0 $Y2=0
cc_3509 N_VPWR_c_4288_n N_A_2603_297#_c_6989_n 7.64992e-19 $X=14.03 $Y=2.72
+ $X2=0 $Y2=0
cc_3510 N_VPWR_c_4258_n N_A_2603_297#_c_7015_n 0.00163482f $X=13.61 $Y=2.34
+ $X2=0 $Y2=0
cc_3511 VPWR N_A_2603_297#_c_7015_n 0.0296407f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3512 VPWR N_A_2603_297#_c_6994_n 0.0618665f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3513 N_VPWR_c_4258_n N_A_2603_297#_c_6996_n 0.00265921f $X=13.61 $Y=2.34
+ $X2=0 $Y2=0
cc_3514 VPWR N_A_2603_297#_c_6996_n 0.0299024f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3515 N_VPWR_c_4288_n N_A_2603_297#_c_6996_n 4.8162e-19 $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_3516 N_VPWR_c_4258_n N_A_2603_297#_c_6979_n 0.0106781f $X=13.61 $Y=2.34 $X2=0
+ $Y2=0
cc_3517 VPWR N_A_2603_297#_c_6979_n 0.00317333f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3518 N_VPWR_c_4287_n N_A_2603_297#_c_6979_n 0.020978f $X=13.475 $Y=2.72 $X2=0
+ $Y2=0
cc_3519 N_VPWR_c_4258_n N_A_2603_297#_c_6997_n 0.0173701f $X=13.61 $Y=2.34 $X2=0
+ $Y2=0
cc_3520 VPWR N_A_2603_297#_c_6997_n 0.00267234f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3521 N_VPWR_c_4288_n N_A_2603_297#_c_6997_n 0.0184771f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_3522 N_VPWR_c_4274_n N_A_2603_297#_c_6980_n 4.83649e-19 $X=15.935 $Y=2.72
+ $X2=0 $Y2=0
cc_3523 VPWR N_A_2603_297#_c_6980_n 0.0299832f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3524 N_VPWR_c_4274_n N_A_2603_297#_c_6999_n 0.0217548f $X=15.935 $Y=2.72
+ $X2=0 $Y2=0
cc_3525 VPWR N_A_2603_297#_c_6999_n 0.00303374f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3526 N_VPWR_c_4478_n N_A_2603_297#_c_6992_n 0.0173701f $X=13.61 $Y=1.94 $X2=0
+ $Y2=0
cc_3527 N_VPWR_c_4258_n N_A_2603_297#_c_6982_n 0.00235484f $X=13.61 $Y=2.34
+ $X2=0 $Y2=0
cc_3528 N_VPWR_c_4478_n N_A_2603_297#_c_6982_n 0.0115021f $X=13.61 $Y=1.94 $X2=0
+ $Y2=0
cc_3529 VPWR N_A_2603_591#_M1038_d 0.00111289f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=1.305
cc_3530 VPWR N_A_2603_591#_M1088_d 0.00165645f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3531 VPWR N_A_2603_591#_M1159_d 0.00127413f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3532 N_VPWR_c_4259_n N_A_2603_591#_c_7072_n 0.00235484f $X=13.61 $Y=3.1 $X2=0
+ $Y2=0
cc_3533 N_VPWR_c_4486_n N_A_2603_591#_c_7072_n 0.0115021f $X=13.61 $Y=3.5 $X2=0
+ $Y2=0
cc_3534 N_VPWR_M1038_s N_A_2603_591#_c_7077_n 0.00331615f $X=13.465 $Y=2.955
+ $X2=0 $Y2=0
cc_3535 N_VPWR_c_4486_n N_A_2603_591#_c_7077_n 0.0158304f $X=13.61 $Y=3.5 $X2=0
+ $Y2=0
cc_3536 N_VPWR_c_4259_n N_A_2603_591#_c_7088_n 0.00995242f $X=13.61 $Y=3.1 $X2=0
+ $Y2=0
cc_3537 VPWR N_A_2603_591#_c_7088_n 0.00247808f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3538 N_VPWR_c_4288_n N_A_2603_591#_c_7088_n 0.0173868f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_3539 N_VPWR_c_4274_n N_A_2603_591#_c_7074_n 0.0218871f $X=15.935 $Y=2.72
+ $X2=0 $Y2=0
cc_3540 VPWR N_A_2603_591#_c_7074_n 0.00305107f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3541 N_VPWR_c_4259_n N_A_2603_591#_c_7083_n 0.0170179f $X=13.61 $Y=3.1 $X2=0
+ $Y2=0
cc_3542 N_VPWR_c_4486_n N_A_2603_591#_c_7083_n 3.68476e-19 $X=13.61 $Y=3.5 $X2=0
+ $Y2=0
cc_3543 VPWR N_A_2603_591#_c_7083_n 0.0560119f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3544 N_VPWR_c_4287_n N_A_2603_591#_c_7083_n 7.71354e-19 $X=13.475 $Y=2.72
+ $X2=0 $Y2=0
cc_3545 N_VPWR_c_4288_n N_A_2603_591#_c_7083_n 7.64992e-19 $X=14.03 $Y=2.72
+ $X2=0 $Y2=0
cc_3546 N_VPWR_c_4259_n N_A_2603_591#_c_7115_n 0.00163482f $X=13.61 $Y=3.1 $X2=0
+ $Y2=0
cc_3547 VPWR N_A_2603_591#_c_7115_n 0.0296407f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3548 VPWR N_A_2603_591#_c_7093_n 0.0621437f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3549 N_VPWR_c_4259_n N_A_2603_591#_c_7095_n 0.00267717f $X=13.61 $Y=3.1 $X2=0
+ $Y2=0
cc_3550 VPWR N_A_2603_591#_c_7095_n 0.0298971f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3551 N_VPWR_c_4288_n N_A_2603_591#_c_7095_n 4.77412e-19 $X=14.03 $Y=2.72
+ $X2=0 $Y2=0
cc_3552 N_VPWR_c_4259_n N_A_2603_591#_c_7085_n 0.0247455f $X=13.61 $Y=3.1 $X2=0
+ $Y2=0
cc_3553 N_VPWR_c_4274_n N_A_2603_591#_c_7075_n 4.78963e-19 $X=15.935 $Y=2.72
+ $X2=0 $Y2=0
cc_3554 VPWR N_A_2603_591#_c_7075_n 0.0299779f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3555 N_VPWR_c_4259_n N_A_2603_591#_c_7076_n 0.0106781f $X=13.61 $Y=3.1 $X2=0
+ $Y2=0
cc_3556 VPWR N_A_2603_591#_c_7076_n 0.00317333f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3557 N_VPWR_c_4287_n N_A_2603_591#_c_7076_n 0.020978f $X=13.475 $Y=2.72 $X2=0
+ $Y2=0
cc_3558 VPWR N_A_3400_333#_M1055_d 0.00127816f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=1.305
cc_3559 VPWR N_A_3400_333#_M1082_d 0.00166446f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3560 VPWR N_A_3400_333#_M1079_d 0.00111289f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3561 N_VPWR_M1051_s N_A_3400_333#_c_7181_n 0.00331615f $X=18.445 $Y=1.485
+ $X2=0 $Y2=0
cc_3562 N_VPWR_c_4548_n N_A_3400_333#_c_7181_n 0.0158304f $X=18.59 $Y=1.94 $X2=0
+ $Y2=0
cc_3563 VPWR N_A_3400_333#_c_7170_n 0.0618665f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3564 VPWR N_A_3400_333#_c_7165_n 0.0299832f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3565 N_VPWR_c_4289_n N_A_3400_333#_c_7165_n 4.83649e-19 $X=17.25 $Y=2.72
+ $X2=0 $Y2=0
cc_3566 N_VPWR_c_4262_n N_A_3400_333#_c_7187_n 0.0170179f $X=18.59 $Y=2.34 $X2=0
+ $Y2=0
cc_3567 N_VPWR_c_4548_n N_A_3400_333#_c_7187_n 3.68476e-19 $X=18.59 $Y=1.94
+ $X2=0 $Y2=0
cc_3568 VPWR N_A_3400_333#_c_7187_n 0.0560119f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3569 N_VPWR_c_4290_n N_A_3400_333#_c_7187_n 7.64992e-19 $X=18.425 $Y=2.72
+ $X2=0 $Y2=0
cc_3570 N_VPWR_c_4291_n N_A_3400_333#_c_7187_n 7.71354e-19 $X=19.915 $Y=2.72
+ $X2=0 $Y2=0
cc_3571 N_VPWR_c_4262_n N_A_3400_333#_c_7173_n 0.00265921f $X=18.59 $Y=2.34
+ $X2=0 $Y2=0
cc_3572 VPWR N_A_3400_333#_c_7173_n 0.0299024f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3573 N_VPWR_c_4290_n N_A_3400_333#_c_7173_n 4.8162e-19 $X=18.425 $Y=2.72
+ $X2=0 $Y2=0
cc_3574 VPWR N_A_3400_333#_c_7174_n 0.00303374f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3575 N_VPWR_c_4289_n N_A_3400_333#_c_7174_n 0.0217548f $X=17.25 $Y=2.72 $X2=0
+ $Y2=0
cc_3576 N_VPWR_c_4262_n N_A_3400_333#_c_7175_n 0.0173701f $X=18.59 $Y=2.34 $X2=0
+ $Y2=0
cc_3577 VPWR N_A_3400_333#_c_7175_n 0.00267234f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3578 N_VPWR_c_4290_n N_A_3400_333#_c_7175_n 0.0184771f $X=18.425 $Y=2.72
+ $X2=0 $Y2=0
cc_3579 N_VPWR_c_4262_n N_A_3400_333#_c_7212_n 0.00163482f $X=18.59 $Y=2.34
+ $X2=0 $Y2=0
cc_3580 VPWR N_A_3400_333#_c_7212_n 0.0296407f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3581 N_VPWR_c_4262_n N_A_3400_333#_c_7166_n 0.0106781f $X=18.59 $Y=2.34 $X2=0
+ $Y2=0
cc_3582 VPWR N_A_3400_333#_c_7166_n 0.00317333f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3583 N_VPWR_c_4291_n N_A_3400_333#_c_7166_n 0.020978f $X=19.915 $Y=2.72 $X2=0
+ $Y2=0
cc_3584 N_VPWR_c_4548_n N_A_3400_333#_c_7180_n 0.0173701f $X=18.59 $Y=1.94 $X2=0
+ $Y2=0
cc_3585 N_VPWR_c_4262_n N_A_3400_333#_c_7168_n 0.00235484f $X=18.59 $Y=2.34
+ $X2=0 $Y2=0
cc_3586 N_VPWR_c_4548_n N_A_3400_333#_c_7168_n 0.0115021f $X=18.59 $Y=1.94 $X2=0
+ $Y2=0
cc_3587 VPWR N_A_3400_591#_M1134_d 0.00127413f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=1.305
cc_3588 VPWR N_A_3400_591#_M1158_d 0.00165645f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3589 VPWR N_A_3400_591#_M1087_d 0.00111289f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3590 N_VPWR_M1058_s N_A_3400_591#_c_7260_n 0.00331615f $X=18.445 $Y=2.955
+ $X2=0 $Y2=0
cc_3591 N_VPWR_c_4556_n N_A_3400_591#_c_7260_n 0.015867f $X=18.59 $Y=3.5 $X2=0
+ $Y2=0
cc_3592 N_VPWR_c_4263_n N_A_3400_591#_c_7261_n 0.00235484f $X=18.59 $Y=3.1 $X2=0
+ $Y2=0
cc_3593 N_VPWR_c_4556_n N_A_3400_591#_c_7261_n 0.0115021f $X=18.59 $Y=3.5 $X2=0
+ $Y2=0
cc_3594 VPWR N_A_3400_591#_c_7262_n 0.00305107f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3595 N_VPWR_c_4289_n N_A_3400_591#_c_7262_n 0.0218871f $X=17.25 $Y=2.72 $X2=0
+ $Y2=0
cc_3596 N_VPWR_c_4263_n N_A_3400_591#_c_7270_n 0.00995242f $X=18.59 $Y=3.1 $X2=0
+ $Y2=0
cc_3597 VPWR N_A_3400_591#_c_7270_n 0.00247808f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3598 N_VPWR_c_4290_n N_A_3400_591#_c_7270_n 0.0173868f $X=18.425 $Y=2.72
+ $X2=0 $Y2=0
cc_3599 VPWR N_A_3400_591#_c_7271_n 0.0621437f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3600 VPWR N_A_3400_591#_c_7263_n 0.0299779f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3601 N_VPWR_c_4289_n N_A_3400_591#_c_7263_n 4.78963e-19 $X=17.25 $Y=2.72
+ $X2=0 $Y2=0
cc_3602 N_VPWR_c_4263_n N_A_3400_591#_c_7280_n 0.0170179f $X=18.59 $Y=3.1 $X2=0
+ $Y2=0
cc_3603 N_VPWR_c_4556_n N_A_3400_591#_c_7280_n 3.57652e-19 $X=18.59 $Y=3.5 $X2=0
+ $Y2=0
cc_3604 VPWR N_A_3400_591#_c_7280_n 0.0560119f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3605 N_VPWR_c_4290_n N_A_3400_591#_c_7280_n 7.64992e-19 $X=18.425 $Y=2.72
+ $X2=0 $Y2=0
cc_3606 N_VPWR_c_4291_n N_A_3400_591#_c_7280_n 7.71354e-19 $X=19.915 $Y=2.72
+ $X2=0 $Y2=0
cc_3607 N_VPWR_c_4263_n N_A_3400_591#_c_7274_n 0.00267717f $X=18.59 $Y=3.1 $X2=0
+ $Y2=0
cc_3608 VPWR N_A_3400_591#_c_7274_n 0.0298971f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3609 N_VPWR_c_4290_n N_A_3400_591#_c_7274_n 4.77412e-19 $X=18.425 $Y=2.72
+ $X2=0 $Y2=0
cc_3610 N_VPWR_c_4263_n N_A_3400_591#_c_7275_n 0.0247455f $X=18.59 $Y=3.1 $X2=0
+ $Y2=0
cc_3611 N_VPWR_c_4263_n N_A_3400_591#_c_7308_n 0.00163482f $X=18.59 $Y=3.1 $X2=0
+ $Y2=0
cc_3612 VPWR N_A_3400_591#_c_7308_n 0.0296407f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3613 N_VPWR_c_4263_n N_A_3400_591#_c_7264_n 0.0106781f $X=18.59 $Y=3.1 $X2=0
+ $Y2=0
cc_3614 VPWR N_A_3400_591#_c_7264_n 0.00317333f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3615 N_VPWR_c_4291_n N_A_3400_591#_c_7264_n 0.020978f $X=19.915 $Y=2.72 $X2=0
+ $Y2=0
cc_3616 VPWR N_A_3891_297#_M1062_d 0.00111289f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=1.305
cc_3617 VPWR N_A_3891_297#_M1143_d 0.00166446f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3618 VPWR N_A_3891_297#_M1091_d 0.00127816f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3619 N_VPWR_M1062_s N_A_3891_297#_c_7358_n 0.00331615f $X=19.905 $Y=1.485
+ $X2=0 $Y2=0
cc_3620 N_VPWR_c_4564_n N_A_3891_297#_c_7358_n 0.0158304f $X=20.05 $Y=1.94 $X2=0
+ $Y2=0
cc_3621 N_VPWR_c_4264_n N_A_3891_297#_c_7362_n 0.0170179f $X=20.05 $Y=2.34 $X2=0
+ $Y2=0
cc_3622 N_VPWR_c_4564_n N_A_3891_297#_c_7362_n 3.68476e-19 $X=20.05 $Y=1.94
+ $X2=0 $Y2=0
cc_3623 VPWR N_A_3891_297#_c_7362_n 0.0560119f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3624 N_VPWR_c_4291_n N_A_3891_297#_c_7362_n 7.71354e-19 $X=19.915 $Y=2.72
+ $X2=0 $Y2=0
cc_3625 N_VPWR_c_4292_n N_A_3891_297#_c_7362_n 7.64992e-19 $X=20.47 $Y=2.72
+ $X2=0 $Y2=0
cc_3626 N_VPWR_c_4264_n N_A_3891_297#_c_7388_n 0.00163482f $X=20.05 $Y=2.34
+ $X2=0 $Y2=0
cc_3627 VPWR N_A_3891_297#_c_7388_n 0.0296407f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3628 VPWR N_A_3891_297#_c_7367_n 0.0618665f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3629 N_VPWR_c_4264_n N_A_3891_297#_c_7369_n 0.00265921f $X=20.05 $Y=2.34
+ $X2=0 $Y2=0
cc_3630 VPWR N_A_3891_297#_c_7369_n 0.0299024f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3631 N_VPWR_c_4292_n N_A_3891_297#_c_7369_n 4.8162e-19 $X=20.47 $Y=2.72 $X2=0
+ $Y2=0
cc_3632 N_VPWR_c_4264_n N_A_3891_297#_c_7352_n 0.0106781f $X=20.05 $Y=2.34 $X2=0
+ $Y2=0
cc_3633 VPWR N_A_3891_297#_c_7352_n 0.00317333f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3634 N_VPWR_c_4291_n N_A_3891_297#_c_7352_n 0.020978f $X=19.915 $Y=2.72 $X2=0
+ $Y2=0
cc_3635 N_VPWR_c_4264_n N_A_3891_297#_c_7370_n 0.0173701f $X=20.05 $Y=2.34 $X2=0
+ $Y2=0
cc_3636 VPWR N_A_3891_297#_c_7370_n 0.00267234f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3637 N_VPWR_c_4292_n N_A_3891_297#_c_7370_n 0.0184771f $X=20.47 $Y=2.72 $X2=0
+ $Y2=0
cc_3638 N_VPWR_c_4276_n N_A_3891_297#_c_7353_n 4.83649e-19 $X=22.375 $Y=2.72
+ $X2=0 $Y2=0
cc_3639 VPWR N_A_3891_297#_c_7353_n 0.0299832f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3640 N_VPWR_c_4276_n N_A_3891_297#_c_7372_n 0.0217548f $X=22.375 $Y=2.72
+ $X2=0 $Y2=0
cc_3641 VPWR N_A_3891_297#_c_7372_n 0.00303374f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3642 N_VPWR_c_4564_n N_A_3891_297#_c_7365_n 0.0173701f $X=20.05 $Y=1.94 $X2=0
+ $Y2=0
cc_3643 N_VPWR_c_4264_n N_A_3891_297#_c_7355_n 0.00235484f $X=20.05 $Y=2.34
+ $X2=0 $Y2=0
cc_3644 N_VPWR_c_4564_n N_A_3891_297#_c_7355_n 0.0115021f $X=20.05 $Y=1.94 $X2=0
+ $Y2=0
cc_3645 VPWR N_A_3891_591#_M1069_d 0.00111289f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=1.305
cc_3646 VPWR N_A_3891_591#_M1152_d 0.00165645f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3647 VPWR N_A_3891_591#_M1140_s 0.00127413f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3648 N_VPWR_c_4265_n N_A_3891_591#_c_7445_n 0.00235484f $X=20.05 $Y=3.1 $X2=0
+ $Y2=0
cc_3649 N_VPWR_c_4572_n N_A_3891_591#_c_7445_n 0.0115021f $X=20.05 $Y=3.5 $X2=0
+ $Y2=0
cc_3650 N_VPWR_M1069_s N_A_3891_591#_c_7450_n 0.00331615f $X=19.905 $Y=2.955
+ $X2=0 $Y2=0
cc_3651 N_VPWR_c_4572_n N_A_3891_591#_c_7450_n 0.0158304f $X=20.05 $Y=3.5 $X2=0
+ $Y2=0
cc_3652 N_VPWR_c_4265_n N_A_3891_591#_c_7461_n 0.00995242f $X=20.05 $Y=3.1 $X2=0
+ $Y2=0
cc_3653 VPWR N_A_3891_591#_c_7461_n 0.00247808f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3654 N_VPWR_c_4292_n N_A_3891_591#_c_7461_n 0.0173868f $X=20.47 $Y=2.72 $X2=0
+ $Y2=0
cc_3655 N_VPWR_c_4276_n N_A_3891_591#_c_7447_n 0.0218871f $X=22.375 $Y=2.72
+ $X2=0 $Y2=0
cc_3656 VPWR N_A_3891_591#_c_7447_n 0.00305107f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3657 N_VPWR_c_4265_n N_A_3891_591#_c_7456_n 0.0170179f $X=20.05 $Y=3.1 $X2=0
+ $Y2=0
cc_3658 N_VPWR_c_4572_n N_A_3891_591#_c_7456_n 3.68476e-19 $X=20.05 $Y=3.5 $X2=0
+ $Y2=0
cc_3659 VPWR N_A_3891_591#_c_7456_n 0.0560119f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3660 N_VPWR_c_4291_n N_A_3891_591#_c_7456_n 7.71354e-19 $X=19.915 $Y=2.72
+ $X2=0 $Y2=0
cc_3661 N_VPWR_c_4292_n N_A_3891_591#_c_7456_n 7.64992e-19 $X=20.47 $Y=2.72
+ $X2=0 $Y2=0
cc_3662 N_VPWR_c_4265_n N_A_3891_591#_c_7488_n 0.00163482f $X=20.05 $Y=3.1 $X2=0
+ $Y2=0
cc_3663 VPWR N_A_3891_591#_c_7488_n 0.0296407f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3664 VPWR N_A_3891_591#_c_7466_n 0.0621437f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3665 N_VPWR_c_4265_n N_A_3891_591#_c_7468_n 0.00267717f $X=20.05 $Y=3.1 $X2=0
+ $Y2=0
cc_3666 VPWR N_A_3891_591#_c_7468_n 0.0298971f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3667 N_VPWR_c_4292_n N_A_3891_591#_c_7468_n 4.77412e-19 $X=20.47 $Y=2.72
+ $X2=0 $Y2=0
cc_3668 N_VPWR_c_4265_n N_A_3891_591#_c_7458_n 0.0247455f $X=20.05 $Y=3.1 $X2=0
+ $Y2=0
cc_3669 N_VPWR_c_4276_n N_A_3891_591#_c_7448_n 4.78963e-19 $X=22.375 $Y=2.72
+ $X2=0 $Y2=0
cc_3670 VPWR N_A_3891_591#_c_7448_n 0.0299779f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3671 N_VPWR_c_4265_n N_A_3891_591#_c_7449_n 0.0106781f $X=20.05 $Y=3.1 $X2=0
+ $Y2=0
cc_3672 VPWR N_A_3891_591#_c_7449_n 0.00317333f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3673 N_VPWR_c_4291_n N_A_3891_591#_c_7449_n 0.020978f $X=19.915 $Y=2.72 $X2=0
+ $Y2=0
cc_3674 VPWR N_A_4688_333#_M1122_d 0.00127816f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=1.305
cc_3675 VPWR N_A_4688_333#_M1148_d 0.00166446f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3676 VPWR N_A_4688_333#_M1142_d 0.00111289f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3677 N_VPWR_M1061_s N_A_4688_333#_c_7554_n 0.00346031f $X=24.885 $Y=1.485
+ $X2=0 $Y2=0
cc_3678 N_VPWR_c_4634_n N_A_4688_333#_c_7554_n 0.0164726f $X=25.03 $Y=1.94 $X2=0
+ $Y2=0
cc_3679 VPWR N_A_4688_333#_c_7543_n 0.0618665f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3680 VPWR N_A_4688_333#_c_7538_n 0.0299832f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3681 N_VPWR_c_4293_n N_A_4688_333#_c_7538_n 4.83649e-19 $X=23.69 $Y=2.72
+ $X2=0 $Y2=0
cc_3682 N_VPWR_c_4268_n N_A_4688_333#_c_7560_n 0.0174313f $X=25.03 $Y=2.34 $X2=0
+ $Y2=0
cc_3683 N_VPWR_c_4634_n N_A_4688_333#_c_7560_n 8.54514e-19 $X=25.03 $Y=1.94
+ $X2=0 $Y2=0
cc_3684 VPWR N_A_4688_333#_c_7560_n 0.0560119f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3685 N_VPWR_c_4294_n N_A_4688_333#_c_7560_n 7.64992e-19 $X=24.865 $Y=2.72
+ $X2=0 $Y2=0
cc_3686 N_VPWR_c_4295_n N_A_4688_333#_c_7560_n 7.71354e-19 $X=25.53 $Y=2.72
+ $X2=0 $Y2=0
cc_3687 N_VPWR_c_4268_n N_A_4688_333#_c_7546_n 0.00265921f $X=25.03 $Y=2.34
+ $X2=0 $Y2=0
cc_3688 VPWR N_A_4688_333#_c_7546_n 0.0299024f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3689 N_VPWR_c_4294_n N_A_4688_333#_c_7546_n 4.8162e-19 $X=24.865 $Y=2.72
+ $X2=0 $Y2=0
cc_3690 VPWR N_A_4688_333#_c_7547_n 0.00303374f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3691 N_VPWR_c_4293_n N_A_4688_333#_c_7547_n 0.0217548f $X=23.69 $Y=2.72 $X2=0
+ $Y2=0
cc_3692 N_VPWR_c_4268_n N_A_4688_333#_c_7548_n 0.0177079f $X=25.03 $Y=2.34 $X2=0
+ $Y2=0
cc_3693 VPWR N_A_4688_333#_c_7548_n 0.00267234f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3694 N_VPWR_c_4294_n N_A_4688_333#_c_7548_n 0.0184771f $X=24.865 $Y=2.72
+ $X2=0 $Y2=0
cc_3695 N_VPWR_c_4268_n N_A_4688_333#_c_7585_n 0.00163482f $X=25.03 $Y=2.34
+ $X2=0 $Y2=0
cc_3696 VPWR N_A_4688_333#_c_7585_n 0.0296407f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3697 N_VPWR_c_4268_n N_A_4688_333#_c_7539_n 0.0106781f $X=25.03 $Y=2.34 $X2=0
+ $Y2=0
cc_3698 VPWR N_A_4688_333#_c_7539_n 0.0035565f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3699 N_VPWR_c_4295_n N_A_4688_333#_c_7539_n 0.020978f $X=25.53 $Y=2.72 $X2=0
+ $Y2=0
cc_3700 N_VPWR_c_4634_n N_A_4688_333#_c_7553_n 0.0177079f $X=25.03 $Y=1.94 $X2=0
+ $Y2=0
cc_3701 N_VPWR_c_4268_n N_A_4688_333#_c_7541_n 0.00235484f $X=25.03 $Y=2.34
+ $X2=0 $Y2=0
cc_3702 VPWR N_A_4688_591#_M1049_d 0.00127413f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=1.305
cc_3703 VPWR N_A_4688_591#_M1076_d 0.00165645f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3704 VPWR N_A_4688_591#_M1149_d 0.00111289f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3705 N_VPWR_M1068_s N_A_4688_591#_c_7617_n 0.00346031f $X=24.885 $Y=2.955
+ $X2=0 $Y2=0
cc_3706 N_VPWR_c_4642_n N_A_4688_591#_c_7617_n 0.0164726f $X=25.03 $Y=3.5 $X2=0
+ $Y2=0
cc_3707 N_VPWR_c_4269_n N_A_4688_591#_c_7618_n 0.00235484f $X=25.03 $Y=3.1 $X2=0
+ $Y2=0
cc_3708 VPWR N_A_4688_591#_c_7619_n 0.00305107f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3709 N_VPWR_c_4293_n N_A_4688_591#_c_7619_n 0.0218871f $X=23.69 $Y=2.72 $X2=0
+ $Y2=0
cc_3710 N_VPWR_c_4269_n N_A_4688_591#_c_7627_n 0.00995242f $X=25.03 $Y=3.1 $X2=0
+ $Y2=0
cc_3711 VPWR N_A_4688_591#_c_7627_n 0.00247808f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3712 N_VPWR_c_4294_n N_A_4688_591#_c_7627_n 0.0173868f $X=24.865 $Y=2.72
+ $X2=0 $Y2=0
cc_3713 VPWR N_A_4688_591#_c_7628_n 0.0621437f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3714 VPWR N_A_4688_591#_c_7620_n 0.0299779f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3715 N_VPWR_c_4293_n N_A_4688_591#_c_7620_n 4.78963e-19 $X=23.69 $Y=2.72
+ $X2=0 $Y2=0
cc_3716 N_VPWR_c_4269_n N_A_4688_591#_c_7637_n 0.0174313f $X=25.03 $Y=3.1 $X2=0
+ $Y2=0
cc_3717 N_VPWR_c_4642_n N_A_4688_591#_c_7637_n 8.43691e-19 $X=25.03 $Y=3.5 $X2=0
+ $Y2=0
cc_3718 VPWR N_A_4688_591#_c_7637_n 0.0560119f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3719 N_VPWR_c_4294_n N_A_4688_591#_c_7637_n 7.64992e-19 $X=24.865 $Y=2.72
+ $X2=0 $Y2=0
cc_3720 N_VPWR_c_4295_n N_A_4688_591#_c_7637_n 7.71354e-19 $X=25.53 $Y=2.72
+ $X2=0 $Y2=0
cc_3721 N_VPWR_c_4269_n N_A_4688_591#_c_7631_n 0.00267717f $X=25.03 $Y=3.1 $X2=0
+ $Y2=0
cc_3722 VPWR N_A_4688_591#_c_7631_n 0.0298971f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3723 N_VPWR_c_4294_n N_A_4688_591#_c_7631_n 4.77412e-19 $X=24.865 $Y=2.72
+ $X2=0 $Y2=0
cc_3724 N_VPWR_c_4269_n N_A_4688_591#_c_7632_n 0.0254212f $X=25.03 $Y=3.1 $X2=0
+ $Y2=0
cc_3725 N_VPWR_c_4269_n N_A_4688_591#_c_7664_n 0.00163482f $X=25.03 $Y=3.1 $X2=0
+ $Y2=0
cc_3726 VPWR N_A_4688_591#_c_7664_n 0.0296407f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3727 N_VPWR_c_4269_n N_A_4688_591#_c_7621_n 0.0106781f $X=25.03 $Y=3.1 $X2=0
+ $Y2=0
cc_3728 VPWR N_A_4688_591#_c_7621_n 0.0035565f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_3729 N_VPWR_c_4295_n N_A_4688_591#_c_7621_n 0.020978f $X=25.53 $Y=2.72 $X2=0
+ $Y2=0
cc_3730 N_Z_c_5242_n N_A_824_333#_M1084_d 0.00197114f $X=4.685 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_3731 N_Z_c_5244_n N_A_824_333#_M1113_d 0.00580444f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3732 N_Z_c_5244_n N_A_824_333#_c_6435_n 0.0237468f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3733 N_Z_c_5227_n N_A_824_333#_c_6423_n 0.00930189f $X=4.76 $Y=1.755 $X2=0
+ $Y2=0
cc_3734 N_Z_M1084_s N_A_824_333#_c_6424_n 0.00154628f $X=4.57 $Y=1.665 $X2=0
+ $Y2=0
cc_3735 N_Z_c_5242_n N_A_824_333#_c_6424_n 0.0225177f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_3736 N_Z_c_5244_n N_A_824_333#_c_6424_n 0.00942629f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3737 N_Z_c_5357_n N_A_824_333#_c_6424_n 0.0241216f $X=4.975 $Y=1.87 $X2=0
+ $Y2=0
cc_3738 N_Z_c_5358_n N_A_824_333#_c_6424_n 0.00832432f $X=4.83 $Y=1.87 $X2=0
+ $Y2=0
cc_3739 N_Z_c_5259_n N_A_824_333#_c_6424_n 0.0115376f $X=4.76 $Y=3.315 $X2=0
+ $Y2=0
cc_3740 N_Z_c_5242_n N_A_824_333#_c_6419_n 0.0249588f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_3741 N_Z_c_5358_n N_A_824_333#_c_6419_n 4.48979e-19 $X=4.83 $Y=1.87 $X2=0
+ $Y2=0
cc_3742 N_Z_c_5259_n N_A_824_333#_c_6419_n 2.4892e-19 $X=4.76 $Y=3.315 $X2=0
+ $Y2=0
cc_3743 N_Z_c_5244_n N_A_824_333#_c_6441_n 0.048455f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3744 N_Z_c_5244_n N_A_824_333#_c_6427_n 0.0249366f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3745 N_Z_c_5358_n N_A_824_333#_c_6427_n 4.5829e-19 $X=4.83 $Y=1.87 $X2=0
+ $Y2=0
cc_3746 N_Z_c_5259_n N_A_824_333#_c_6427_n 2.82292e-19 $X=4.76 $Y=3.315 $X2=0
+ $Y2=0
cc_3747 N_Z_c_5242_n N_A_824_333#_c_6428_n 0.0016886f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_3748 N_Z_c_5259_n N_A_824_333#_c_6428_n 0.0123065f $X=4.76 $Y=3.315 $X2=0
+ $Y2=0
cc_3749 N_Z_c_5244_n N_A_824_333#_c_6429_n 7.67921e-19 $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3750 N_Z_c_5244_n N_A_824_333#_c_6466_n 0.0237143f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3751 N_Z_c_5242_n N_A_824_333#_c_6421_n 0.0109134f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_3752 N_Z_c_5357_n N_A_824_333#_c_6421_n 4.86317e-19 $X=4.975 $Y=1.87 $X2=0
+ $Y2=0
cc_3753 N_Z_c_5358_n N_A_824_333#_c_6421_n 0.0210951f $X=4.83 $Y=1.87 $X2=0
+ $Y2=0
cc_3754 N_Z_c_5227_n N_A_824_333#_c_6421_n 0.00468052f $X=4.76 $Y=1.755 $X2=0
+ $Y2=0
cc_3755 N_Z_c_5259_n N_A_824_333#_c_6421_n 0.00373869f $X=4.76 $Y=3.315 $X2=0
+ $Y2=0
cc_3756 N_Z_c_5244_n N_A_824_333#_c_6434_n 0.0166619f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3757 N_Z_c_5357_n N_A_824_333#_c_6434_n 0.00221246f $X=4.975 $Y=1.87 $X2=0
+ $Y2=0
cc_3758 N_Z_c_5358_n N_A_824_333#_c_6434_n 0.0240318f $X=4.83 $Y=1.87 $X2=0
+ $Y2=0
cc_3759 N_Z_c_5259_n N_A_824_333#_c_6434_n 0.00347206f $X=4.76 $Y=3.315 $X2=0
+ $Y2=0
cc_3760 N_Z_c_5244_n N_A_824_333#_c_6422_n 0.018076f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3761 N_Z_c_5243_n N_A_824_591#_M1036_s 0.00197114f $X=4.685 $Y=3.57 $X2=-0.19
+ $Y2=-0.24
cc_3762 N_Z_c_5245_n N_A_824_591#_M1157_s 0.0058104f $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3763 N_Z_c_5245_n N_A_824_591#_c_6514_n 0.0237468f $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3764 N_Z_c_5203_n N_A_824_591#_c_6519_n 0.00930189f $X=4.77 $Y=4.555 $X2=0
+ $Y2=0
cc_3765 N_Z_c_5245_n N_A_824_591#_c_6515_n 0.018076f $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3766 N_Z_c_5203_n N_A_824_591#_c_6516_n 0.00468052f $X=4.77 $Y=4.555 $X2=0
+ $Y2=0
cc_3767 N_Z_c_5243_n N_A_824_591#_c_6516_n 0.0126134f $X=4.685 $Y=3.57 $X2=0
+ $Y2=0
cc_3768 N_Z_c_5383_n N_A_824_591#_c_6516_n 4.86317e-19 $X=4.975 $Y=3.57 $X2=0
+ $Y2=0
cc_3769 N_Z_c_5367_n N_A_824_591#_c_6516_n 0.0210951f $X=4.715 $Y=3.42 $X2=0
+ $Y2=0
cc_3770 N_Z_c_5259_n N_A_824_591#_c_6516_n 0.0161129f $X=4.76 $Y=3.315 $X2=0
+ $Y2=0
cc_3771 N_Z_c_5245_n N_A_824_591#_c_6524_n 3.53114e-19 $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3772 N_Z_M1036_d N_A_824_591#_c_6525_n 0.00154628f $X=4.57 $Y=2.955 $X2=0
+ $Y2=0
cc_3773 N_Z_c_5243_n N_A_824_591#_c_6525_n 0.0225176f $X=4.685 $Y=3.57 $X2=0
+ $Y2=0
cc_3774 N_Z_c_5245_n N_A_824_591#_c_6525_n 0.0094263f $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3775 N_Z_c_5383_n N_A_824_591#_c_6525_n 0.0241216f $X=4.975 $Y=3.57 $X2=0
+ $Y2=0
cc_3776 N_Z_c_5367_n N_A_824_591#_c_6525_n 0.00832432f $X=4.715 $Y=3.42 $X2=0
+ $Y2=0
cc_3777 N_Z_c_5259_n N_A_824_591#_c_6525_n 0.0115376f $X=4.76 $Y=3.315 $X2=0
+ $Y2=0
cc_3778 N_Z_c_5243_n N_A_824_591#_c_6517_n 0.0249588f $X=4.685 $Y=3.57 $X2=0
+ $Y2=0
cc_3779 N_Z_c_5367_n N_A_824_591#_c_6517_n 4.48979e-19 $X=4.715 $Y=3.42 $X2=0
+ $Y2=0
cc_3780 N_Z_c_5259_n N_A_824_591#_c_6517_n 2.48349e-19 $X=4.76 $Y=3.315 $X2=0
+ $Y2=0
cc_3781 N_Z_c_5245_n N_A_824_591#_c_6534_n 0.048455f $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3782 N_Z_c_5245_n N_A_824_591#_c_6528_n 0.0249366f $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3783 N_Z_c_5367_n N_A_824_591#_c_6528_n 4.5829e-19 $X=4.715 $Y=3.42 $X2=0
+ $Y2=0
cc_3784 N_Z_c_5259_n N_A_824_591#_c_6528_n 2.75404e-19 $X=4.76 $Y=3.315 $X2=0
+ $Y2=0
cc_3785 N_Z_c_5245_n N_A_824_591#_c_6529_n 0.0165143f $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3786 N_Z_c_5383_n N_A_824_591#_c_6529_n 0.00221246f $X=4.975 $Y=3.57 $X2=0
+ $Y2=0
cc_3787 N_Z_c_5367_n N_A_824_591#_c_6529_n 0.0240318f $X=4.715 $Y=3.42 $X2=0
+ $Y2=0
cc_3788 N_Z_c_5259_n N_A_824_591#_c_6529_n 0.00349107f $X=4.76 $Y=3.315 $X2=0
+ $Y2=0
cc_3789 N_Z_c_5245_n N_A_824_591#_c_6562_n 0.0237143f $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3790 N_Z_c_5244_n N_A_1315_297#_M1120_s 0.00580444f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3791 N_Z_c_5246_n N_A_1315_297#_M1124_s 0.00197114f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_3792 N_Z_c_5244_n N_A_1315_297#_c_6612_n 0.0237468f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3793 N_Z_c_5228_n N_A_1315_297#_c_6612_n 0.00930189f $X=8.12 $Y=1.755 $X2=0
+ $Y2=0
cc_3794 N_Z_c_5244_n N_A_1315_297#_c_6616_n 0.048455f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3795 N_Z_c_5244_n N_A_1315_297#_c_6642_n 0.0237143f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3796 N_Z_M1005_d N_A_1315_297#_c_6621_n 0.00154628f $X=8.02 $Y=1.665 $X2=0
+ $Y2=0
cc_3797 N_Z_c_5244_n N_A_1315_297#_c_6621_n 0.00942629f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3798 N_Z_c_5246_n N_A_1315_297#_c_6621_n 0.0225177f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_3799 N_Z_c_5426_n N_A_1315_297#_c_6621_n 0.0241216f $X=8.195 $Y=1.87 $X2=0
+ $Y2=0
cc_3800 N_Z_c_5427_n N_A_1315_297#_c_6621_n 0.00835547f $X=8.05 $Y=1.87 $X2=0
+ $Y2=0
cc_3801 N_Z_c_5261_n N_A_1315_297#_c_6621_n 0.0115376f $X=8.12 $Y=3.315 $X2=0
+ $Y2=0
cc_3802 N_Z_c_5244_n N_A_1315_297#_c_6623_n 0.0249366f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3803 N_Z_c_5427_n N_A_1315_297#_c_6623_n 4.5829e-19 $X=8.05 $Y=1.87 $X2=0
+ $Y2=0
cc_3804 N_Z_c_5261_n N_A_1315_297#_c_6623_n 2.82292e-19 $X=8.12 $Y=3.315 $X2=0
+ $Y2=0
cc_3805 N_Z_c_5244_n N_A_1315_297#_c_6624_n 7.67921e-19 $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3806 N_Z_c_5246_n N_A_1315_297#_c_6607_n 0.0249588f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_3807 N_Z_c_5427_n N_A_1315_297#_c_6607_n 4.48979e-19 $X=8.05 $Y=1.87 $X2=0
+ $Y2=0
cc_3808 N_Z_c_5261_n N_A_1315_297#_c_6607_n 2.4892e-19 $X=8.12 $Y=3.315 $X2=0
+ $Y2=0
cc_3809 N_Z_c_5246_n N_A_1315_297#_c_6626_n 0.0016886f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_3810 N_Z_c_5261_n N_A_1315_297#_c_6626_n 0.0123065f $X=8.12 $Y=3.315 $X2=0
+ $Y2=0
cc_3811 N_Z_c_5244_n N_A_1315_297#_c_6619_n 0.0166619f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3812 N_Z_c_5426_n N_A_1315_297#_c_6619_n 0.00221246f $X=8.195 $Y=1.87 $X2=0
+ $Y2=0
cc_3813 N_Z_c_5427_n N_A_1315_297#_c_6619_n 0.0240318f $X=8.05 $Y=1.87 $X2=0
+ $Y2=0
cc_3814 N_Z_c_5261_n N_A_1315_297#_c_6619_n 0.00347206f $X=8.12 $Y=3.315 $X2=0
+ $Y2=0
cc_3815 N_Z_c_5246_n N_A_1315_297#_c_6608_n 0.0109134f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_3816 N_Z_c_5426_n N_A_1315_297#_c_6608_n 4.86317e-19 $X=8.195 $Y=1.87 $X2=0
+ $Y2=0
cc_3817 N_Z_c_5427_n N_A_1315_297#_c_6608_n 0.0210951f $X=8.05 $Y=1.87 $X2=0
+ $Y2=0
cc_3818 N_Z_c_5228_n N_A_1315_297#_c_6608_n 0.00468052f $X=8.12 $Y=1.755 $X2=0
+ $Y2=0
cc_3819 N_Z_c_5261_n N_A_1315_297#_c_6608_n 0.00373869f $X=8.12 $Y=3.315 $X2=0
+ $Y2=0
cc_3820 N_Z_c_5244_n N_A_1315_297#_c_6609_n 0.018076f $X=7.905 $Y=1.87 $X2=0
+ $Y2=0
cc_3821 N_Z_c_5245_n N_A_1315_591#_M1126_s 0.0058104f $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3822 N_Z_c_5247_n N_A_1315_591#_M1095_d 0.00197114f $X=11.125 $Y=3.57 $X2=0
+ $Y2=0
cc_3823 N_Z_c_5245_n N_A_1315_591#_c_6699_n 0.018076f $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3824 N_Z_c_5204_n N_A_1315_591#_c_6704_n 0.00930189f $X=8.11 $Y=4.555 $X2=0
+ $Y2=0
cc_3825 N_Z_c_5245_n N_A_1315_591#_c_6704_n 0.0237468f $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3826 N_Z_c_5245_n N_A_1315_591#_c_6715_n 3.53114e-19 $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3827 N_Z_c_5204_n N_A_1315_591#_c_6701_n 0.00468052f $X=8.11 $Y=4.555 $X2=0
+ $Y2=0
cc_3828 N_Z_c_5247_n N_A_1315_591#_c_6701_n 0.0126134f $X=11.125 $Y=3.57 $X2=0
+ $Y2=0
cc_3829 N_Z_c_5453_n N_A_1315_591#_c_6701_n 4.86317e-19 $X=8.195 $Y=3.57 $X2=0
+ $Y2=0
cc_3830 N_Z_c_5436_n N_A_1315_591#_c_6701_n 0.0210951f $X=8.165 $Y=3.42 $X2=0
+ $Y2=0
cc_3831 N_Z_c_5261_n N_A_1315_591#_c_6701_n 0.0161129f $X=8.12 $Y=3.315 $X2=0
+ $Y2=0
cc_3832 N_Z_c_5245_n N_A_1315_591#_c_6710_n 0.048455f $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3833 N_Z_c_5245_n N_A_1315_591#_c_6742_n 0.0237143f $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3834 N_Z_M1044_s N_A_1315_591#_c_6720_n 0.00154628f $X=8.02 $Y=2.955 $X2=0
+ $Y2=0
cc_3835 N_Z_c_5245_n N_A_1315_591#_c_6720_n 0.0094263f $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3836 N_Z_c_5247_n N_A_1315_591#_c_6720_n 0.0225176f $X=11.125 $Y=3.57 $X2=0
+ $Y2=0
cc_3837 N_Z_c_5453_n N_A_1315_591#_c_6720_n 0.0241216f $X=8.195 $Y=3.57 $X2=0
+ $Y2=0
cc_3838 N_Z_c_5436_n N_A_1315_591#_c_6720_n 0.00835547f $X=8.165 $Y=3.42 $X2=0
+ $Y2=0
cc_3839 N_Z_c_5261_n N_A_1315_591#_c_6720_n 0.0115376f $X=8.12 $Y=3.315 $X2=0
+ $Y2=0
cc_3840 N_Z_c_5245_n N_A_1315_591#_c_6722_n 0.0249366f $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3841 N_Z_c_5436_n N_A_1315_591#_c_6722_n 4.5829e-19 $X=8.165 $Y=3.42 $X2=0
+ $Y2=0
cc_3842 N_Z_c_5261_n N_A_1315_591#_c_6722_n 2.75404e-19 $X=8.12 $Y=3.315 $X2=0
+ $Y2=0
cc_3843 N_Z_c_5245_n N_A_1315_591#_c_6712_n 0.0165143f $X=7.905 $Y=3.57 $X2=0
+ $Y2=0
cc_3844 N_Z_c_5453_n N_A_1315_591#_c_6712_n 0.00221246f $X=8.195 $Y=3.57 $X2=0
+ $Y2=0
cc_3845 N_Z_c_5436_n N_A_1315_591#_c_6712_n 0.0240318f $X=8.165 $Y=3.42 $X2=0
+ $Y2=0
cc_3846 N_Z_c_5261_n N_A_1315_591#_c_6712_n 0.00349107f $X=8.12 $Y=3.315 $X2=0
+ $Y2=0
cc_3847 N_Z_c_5247_n N_A_1315_591#_c_6702_n 0.0249588f $X=11.125 $Y=3.57 $X2=0
+ $Y2=0
cc_3848 N_Z_c_5436_n N_A_1315_591#_c_6702_n 4.48979e-19 $X=8.165 $Y=3.42 $X2=0
+ $Y2=0
cc_3849 N_Z_c_5261_n N_A_1315_591#_c_6702_n 2.48349e-19 $X=8.12 $Y=3.315 $X2=0
+ $Y2=0
cc_3850 N_Z_c_5246_n N_A_2112_333#_M1004_s 0.00197114f $X=11.125 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_3851 N_Z_c_5248_n N_A_2112_333#_M1123_s 0.00580444f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3852 N_Z_c_5248_n N_A_2112_333#_c_6808_n 0.0237468f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3853 N_Z_c_5229_n N_A_2112_333#_c_6796_n 0.00930189f $X=11.2 $Y=1.755 $X2=0
+ $Y2=0
cc_3854 N_Z_M1004_d N_A_2112_333#_c_6797_n 0.00154628f $X=11.01 $Y=1.665 $X2=0
+ $Y2=0
cc_3855 N_Z_c_5246_n N_A_2112_333#_c_6797_n 0.0225177f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_3856 N_Z_c_5248_n N_A_2112_333#_c_6797_n 0.00942629f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3857 N_Z_c_5497_n N_A_2112_333#_c_6797_n 0.0241216f $X=11.415 $Y=1.87 $X2=0
+ $Y2=0
cc_3858 N_Z_c_5498_n N_A_2112_333#_c_6797_n 0.00832432f $X=11.27 $Y=1.87 $X2=0
+ $Y2=0
cc_3859 N_Z_c_5263_n N_A_2112_333#_c_6797_n 0.0115376f $X=11.2 $Y=3.315 $X2=0
+ $Y2=0
cc_3860 N_Z_c_5246_n N_A_2112_333#_c_6792_n 0.0249588f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_3861 N_Z_c_5498_n N_A_2112_333#_c_6792_n 4.48979e-19 $X=11.27 $Y=1.87 $X2=0
+ $Y2=0
cc_3862 N_Z_c_5263_n N_A_2112_333#_c_6792_n 2.4892e-19 $X=11.2 $Y=3.315 $X2=0
+ $Y2=0
cc_3863 N_Z_c_5248_n N_A_2112_333#_c_6814_n 0.048455f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3864 N_Z_c_5248_n N_A_2112_333#_c_6800_n 0.0249366f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3865 N_Z_c_5498_n N_A_2112_333#_c_6800_n 4.5829e-19 $X=11.27 $Y=1.87 $X2=0
+ $Y2=0
cc_3866 N_Z_c_5263_n N_A_2112_333#_c_6800_n 2.82292e-19 $X=11.2 $Y=3.315 $X2=0
+ $Y2=0
cc_3867 N_Z_c_5246_n N_A_2112_333#_c_6801_n 0.0016886f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_3868 N_Z_c_5263_n N_A_2112_333#_c_6801_n 0.0123065f $X=11.2 $Y=3.315 $X2=0
+ $Y2=0
cc_3869 N_Z_c_5248_n N_A_2112_333#_c_6802_n 7.67921e-19 $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3870 N_Z_c_5248_n N_A_2112_333#_c_6839_n 0.0237143f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3871 N_Z_c_5246_n N_A_2112_333#_c_6794_n 0.0109134f $X=11.125 $Y=1.87 $X2=0
+ $Y2=0
cc_3872 N_Z_c_5497_n N_A_2112_333#_c_6794_n 4.86317e-19 $X=11.415 $Y=1.87 $X2=0
+ $Y2=0
cc_3873 N_Z_c_5498_n N_A_2112_333#_c_6794_n 0.0210951f $X=11.27 $Y=1.87 $X2=0
+ $Y2=0
cc_3874 N_Z_c_5229_n N_A_2112_333#_c_6794_n 0.00468052f $X=11.2 $Y=1.755 $X2=0
+ $Y2=0
cc_3875 N_Z_c_5263_n N_A_2112_333#_c_6794_n 0.00373869f $X=11.2 $Y=3.315 $X2=0
+ $Y2=0
cc_3876 N_Z_c_5248_n N_A_2112_333#_c_6807_n 0.0166619f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3877 N_Z_c_5497_n N_A_2112_333#_c_6807_n 0.00221246f $X=11.415 $Y=1.87 $X2=0
+ $Y2=0
cc_3878 N_Z_c_5498_n N_A_2112_333#_c_6807_n 0.0240318f $X=11.27 $Y=1.87 $X2=0
+ $Y2=0
cc_3879 N_Z_c_5263_n N_A_2112_333#_c_6807_n 0.00347206f $X=11.2 $Y=3.315 $X2=0
+ $Y2=0
cc_3880 N_Z_c_5248_n N_A_2112_333#_c_6795_n 0.018076f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3881 N_Z_c_5247_n N_A_2112_591#_M1045_d 0.00197114f $X=11.125 $Y=3.57
+ $X2=-0.19 $Y2=-0.24
cc_3882 N_Z_c_5249_n N_A_2112_591#_M1093_d 0.0058104f $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3883 N_Z_c_5249_n N_A_2112_591#_c_6887_n 0.0237468f $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3884 N_Z_c_5205_n N_A_2112_591#_c_6892_n 0.00930189f $X=11.21 $Y=4.555 $X2=0
+ $Y2=0
cc_3885 N_Z_c_5249_n N_A_2112_591#_c_6888_n 0.018076f $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3886 N_Z_c_5205_n N_A_2112_591#_c_6889_n 0.00468052f $X=11.21 $Y=4.555 $X2=0
+ $Y2=0
cc_3887 N_Z_c_5247_n N_A_2112_591#_c_6889_n 0.0126134f $X=11.125 $Y=3.57 $X2=0
+ $Y2=0
cc_3888 N_Z_c_5523_n N_A_2112_591#_c_6889_n 4.86317e-19 $X=11.415 $Y=3.57 $X2=0
+ $Y2=0
cc_3889 N_Z_c_5507_n N_A_2112_591#_c_6889_n 0.0210951f $X=11.155 $Y=3.42 $X2=0
+ $Y2=0
cc_3890 N_Z_c_5263_n N_A_2112_591#_c_6889_n 0.0161129f $X=11.2 $Y=3.315 $X2=0
+ $Y2=0
cc_3891 N_Z_c_5249_n N_A_2112_591#_c_6897_n 3.53114e-19 $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3892 N_Z_M1045_s N_A_2112_591#_c_6898_n 0.00154628f $X=11.01 $Y=2.955 $X2=0
+ $Y2=0
cc_3893 N_Z_c_5247_n N_A_2112_591#_c_6898_n 0.0225176f $X=11.125 $Y=3.57 $X2=0
+ $Y2=0
cc_3894 N_Z_c_5249_n N_A_2112_591#_c_6898_n 0.0094263f $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3895 N_Z_c_5523_n N_A_2112_591#_c_6898_n 0.0241216f $X=11.415 $Y=3.57 $X2=0
+ $Y2=0
cc_3896 N_Z_c_5507_n N_A_2112_591#_c_6898_n 0.00832432f $X=11.155 $Y=3.42 $X2=0
+ $Y2=0
cc_3897 N_Z_c_5263_n N_A_2112_591#_c_6898_n 0.0115376f $X=11.2 $Y=3.315 $X2=0
+ $Y2=0
cc_3898 N_Z_c_5247_n N_A_2112_591#_c_6890_n 0.0249588f $X=11.125 $Y=3.57 $X2=0
+ $Y2=0
cc_3899 N_Z_c_5507_n N_A_2112_591#_c_6890_n 4.48979e-19 $X=11.155 $Y=3.42 $X2=0
+ $Y2=0
cc_3900 N_Z_c_5263_n N_A_2112_591#_c_6890_n 2.48349e-19 $X=11.2 $Y=3.315 $X2=0
+ $Y2=0
cc_3901 N_Z_c_5249_n N_A_2112_591#_c_6907_n 0.048455f $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3902 N_Z_c_5249_n N_A_2112_591#_c_6901_n 0.0249366f $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3903 N_Z_c_5507_n N_A_2112_591#_c_6901_n 4.5829e-19 $X=11.155 $Y=3.42 $X2=0
+ $Y2=0
cc_3904 N_Z_c_5263_n N_A_2112_591#_c_6901_n 2.75404e-19 $X=11.2 $Y=3.315 $X2=0
+ $Y2=0
cc_3905 N_Z_c_5249_n N_A_2112_591#_c_6902_n 0.0165143f $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3906 N_Z_c_5523_n N_A_2112_591#_c_6902_n 0.00221246f $X=11.415 $Y=3.57 $X2=0
+ $Y2=0
cc_3907 N_Z_c_5507_n N_A_2112_591#_c_6902_n 0.0240318f $X=11.155 $Y=3.42 $X2=0
+ $Y2=0
cc_3908 N_Z_c_5263_n N_A_2112_591#_c_6902_n 0.00349107f $X=11.2 $Y=3.315 $X2=0
+ $Y2=0
cc_3909 N_Z_c_5249_n N_A_2112_591#_c_6935_n 0.0237143f $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3910 N_Z_c_5248_n N_A_2603_297#_M1080_d 0.00580444f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3911 N_Z_c_5250_n N_A_2603_297#_M1083_d 0.00197114f $X=17.565 $Y=1.87 $X2=0
+ $Y2=0
cc_3912 N_Z_c_5248_n N_A_2603_297#_c_6985_n 0.0237468f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3913 N_Z_c_5230_n N_A_2603_297#_c_6985_n 0.00930189f $X=14.56 $Y=1.755 $X2=0
+ $Y2=0
cc_3914 N_Z_c_5248_n N_A_2603_297#_c_6989_n 0.048455f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3915 N_Z_c_5248_n N_A_2603_297#_c_7015_n 0.0237143f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3916 N_Z_M1034_s N_A_2603_297#_c_6994_n 0.00154628f $X=14.46 $Y=1.665 $X2=0
+ $Y2=0
cc_3917 N_Z_c_5248_n N_A_2603_297#_c_6994_n 0.00942629f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3918 N_Z_c_5250_n N_A_2603_297#_c_6994_n 0.0225177f $X=17.565 $Y=1.87 $X2=0
+ $Y2=0
cc_3919 N_Z_c_5566_n N_A_2603_297#_c_6994_n 0.0241216f $X=14.635 $Y=1.87 $X2=0
+ $Y2=0
cc_3920 N_Z_c_5567_n N_A_2603_297#_c_6994_n 0.00835547f $X=14.49 $Y=1.87 $X2=0
+ $Y2=0
cc_3921 N_Z_c_5265_n N_A_2603_297#_c_6994_n 0.0115376f $X=14.56 $Y=3.315 $X2=0
+ $Y2=0
cc_3922 N_Z_c_5248_n N_A_2603_297#_c_6996_n 0.0249366f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3923 N_Z_c_5567_n N_A_2603_297#_c_6996_n 4.5829e-19 $X=14.49 $Y=1.87 $X2=0
+ $Y2=0
cc_3924 N_Z_c_5265_n N_A_2603_297#_c_6996_n 2.82292e-19 $X=14.56 $Y=3.315 $X2=0
+ $Y2=0
cc_3925 N_Z_c_5248_n N_A_2603_297#_c_6997_n 7.67921e-19 $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3926 N_Z_c_5250_n N_A_2603_297#_c_6980_n 0.0249588f $X=17.565 $Y=1.87 $X2=0
+ $Y2=0
cc_3927 N_Z_c_5567_n N_A_2603_297#_c_6980_n 4.48979e-19 $X=14.49 $Y=1.87 $X2=0
+ $Y2=0
cc_3928 N_Z_c_5265_n N_A_2603_297#_c_6980_n 2.4892e-19 $X=14.56 $Y=3.315 $X2=0
+ $Y2=0
cc_3929 N_Z_c_5250_n N_A_2603_297#_c_6999_n 0.0016886f $X=17.565 $Y=1.87 $X2=0
+ $Y2=0
cc_3930 N_Z_c_5265_n N_A_2603_297#_c_6999_n 0.0123065f $X=14.56 $Y=3.315 $X2=0
+ $Y2=0
cc_3931 N_Z_c_5248_n N_A_2603_297#_c_6992_n 0.0166619f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3932 N_Z_c_5566_n N_A_2603_297#_c_6992_n 0.00221246f $X=14.635 $Y=1.87 $X2=0
+ $Y2=0
cc_3933 N_Z_c_5567_n N_A_2603_297#_c_6992_n 0.0240318f $X=14.49 $Y=1.87 $X2=0
+ $Y2=0
cc_3934 N_Z_c_5265_n N_A_2603_297#_c_6992_n 0.00347206f $X=14.56 $Y=3.315 $X2=0
+ $Y2=0
cc_3935 N_Z_c_5250_n N_A_2603_297#_c_6981_n 0.0109134f $X=17.565 $Y=1.87 $X2=0
+ $Y2=0
cc_3936 N_Z_c_5566_n N_A_2603_297#_c_6981_n 4.86317e-19 $X=14.635 $Y=1.87 $X2=0
+ $Y2=0
cc_3937 N_Z_c_5567_n N_A_2603_297#_c_6981_n 0.0210951f $X=14.49 $Y=1.87 $X2=0
+ $Y2=0
cc_3938 N_Z_c_5230_n N_A_2603_297#_c_6981_n 0.00468052f $X=14.56 $Y=1.755 $X2=0
+ $Y2=0
cc_3939 N_Z_c_5265_n N_A_2603_297#_c_6981_n 0.00373869f $X=14.56 $Y=3.315 $X2=0
+ $Y2=0
cc_3940 N_Z_c_5248_n N_A_2603_297#_c_6982_n 0.018076f $X=14.345 $Y=1.87 $X2=0
+ $Y2=0
cc_3941 N_Z_c_5249_n N_A_2603_591#_M1088_d 0.0058104f $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3942 N_Z_c_5251_n N_A_2603_591#_M1159_d 0.00197114f $X=17.565 $Y=3.57 $X2=0
+ $Y2=0
cc_3943 N_Z_c_5249_n N_A_2603_591#_c_7072_n 0.018076f $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3944 N_Z_c_5206_n N_A_2603_591#_c_7077_n 0.00930189f $X=14.55 $Y=4.555 $X2=0
+ $Y2=0
cc_3945 N_Z_c_5249_n N_A_2603_591#_c_7077_n 0.0237468f $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3946 N_Z_c_5249_n N_A_2603_591#_c_7088_n 3.53114e-19 $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3947 N_Z_c_5206_n N_A_2603_591#_c_7074_n 0.00468052f $X=14.55 $Y=4.555 $X2=0
+ $Y2=0
cc_3948 N_Z_c_5251_n N_A_2603_591#_c_7074_n 0.0126134f $X=17.565 $Y=3.57 $X2=0
+ $Y2=0
cc_3949 N_Z_c_5593_n N_A_2603_591#_c_7074_n 4.86317e-19 $X=14.635 $Y=3.57 $X2=0
+ $Y2=0
cc_3950 N_Z_c_5576_n N_A_2603_591#_c_7074_n 0.0210951f $X=14.605 $Y=3.42 $X2=0
+ $Y2=0
cc_3951 N_Z_c_5265_n N_A_2603_591#_c_7074_n 0.0161129f $X=14.56 $Y=3.315 $X2=0
+ $Y2=0
cc_3952 N_Z_c_5249_n N_A_2603_591#_c_7083_n 0.048455f $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3953 N_Z_c_5249_n N_A_2603_591#_c_7115_n 0.0237143f $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3954 N_Z_M1114_s N_A_2603_591#_c_7093_n 0.00154628f $X=14.46 $Y=2.955 $X2=0
+ $Y2=0
cc_3955 N_Z_c_5249_n N_A_2603_591#_c_7093_n 0.0094263f $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3956 N_Z_c_5251_n N_A_2603_591#_c_7093_n 0.0225176f $X=17.565 $Y=3.57 $X2=0
+ $Y2=0
cc_3957 N_Z_c_5593_n N_A_2603_591#_c_7093_n 0.0241216f $X=14.635 $Y=3.57 $X2=0
+ $Y2=0
cc_3958 N_Z_c_5576_n N_A_2603_591#_c_7093_n 0.00835547f $X=14.605 $Y=3.42 $X2=0
+ $Y2=0
cc_3959 N_Z_c_5265_n N_A_2603_591#_c_7093_n 0.0115376f $X=14.56 $Y=3.315 $X2=0
+ $Y2=0
cc_3960 N_Z_c_5249_n N_A_2603_591#_c_7095_n 0.0249366f $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3961 N_Z_c_5576_n N_A_2603_591#_c_7095_n 4.5829e-19 $X=14.605 $Y=3.42 $X2=0
+ $Y2=0
cc_3962 N_Z_c_5265_n N_A_2603_591#_c_7095_n 2.75404e-19 $X=14.56 $Y=3.315 $X2=0
+ $Y2=0
cc_3963 N_Z_c_5249_n N_A_2603_591#_c_7085_n 0.0165143f $X=14.345 $Y=3.57 $X2=0
+ $Y2=0
cc_3964 N_Z_c_5593_n N_A_2603_591#_c_7085_n 0.00221246f $X=14.635 $Y=3.57 $X2=0
+ $Y2=0
cc_3965 N_Z_c_5576_n N_A_2603_591#_c_7085_n 0.0240318f $X=14.605 $Y=3.42 $X2=0
+ $Y2=0
cc_3966 N_Z_c_5265_n N_A_2603_591#_c_7085_n 0.00349107f $X=14.56 $Y=3.315 $X2=0
+ $Y2=0
cc_3967 N_Z_c_5251_n N_A_2603_591#_c_7075_n 0.0249588f $X=17.565 $Y=3.57 $X2=0
+ $Y2=0
cc_3968 N_Z_c_5576_n N_A_2603_591#_c_7075_n 4.48979e-19 $X=14.605 $Y=3.42 $X2=0
+ $Y2=0
cc_3969 N_Z_c_5265_n N_A_2603_591#_c_7075_n 2.48349e-19 $X=14.56 $Y=3.315 $X2=0
+ $Y2=0
cc_3970 N_Z_c_5250_n N_A_3400_333#_M1055_d 0.00197114f $X=17.565 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_3971 N_Z_c_5252_n N_A_3400_333#_M1082_d 0.00580444f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_3972 N_Z_c_5252_n N_A_3400_333#_c_7181_n 0.0237468f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_3973 N_Z_c_5231_n N_A_3400_333#_c_7169_n 0.00930189f $X=17.64 $Y=1.755 $X2=0
+ $Y2=0
cc_3974 N_Z_M1055_s N_A_3400_333#_c_7170_n 0.00154628f $X=17.45 $Y=1.665 $X2=0
+ $Y2=0
cc_3975 N_Z_c_5250_n N_A_3400_333#_c_7170_n 0.0225177f $X=17.565 $Y=1.87 $X2=0
+ $Y2=0
cc_3976 N_Z_c_5252_n N_A_3400_333#_c_7170_n 0.00942629f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_3977 N_Z_c_5637_n N_A_3400_333#_c_7170_n 0.0241216f $X=17.855 $Y=1.87 $X2=0
+ $Y2=0
cc_3978 N_Z_c_5638_n N_A_3400_333#_c_7170_n 0.00832432f $X=17.71 $Y=1.87 $X2=0
+ $Y2=0
cc_3979 N_Z_c_5267_n N_A_3400_333#_c_7170_n 0.0115376f $X=17.64 $Y=3.315 $X2=0
+ $Y2=0
cc_3980 N_Z_c_5250_n N_A_3400_333#_c_7165_n 0.0249588f $X=17.565 $Y=1.87 $X2=0
+ $Y2=0
cc_3981 N_Z_c_5638_n N_A_3400_333#_c_7165_n 4.48979e-19 $X=17.71 $Y=1.87 $X2=0
+ $Y2=0
cc_3982 N_Z_c_5267_n N_A_3400_333#_c_7165_n 2.4892e-19 $X=17.64 $Y=3.315 $X2=0
+ $Y2=0
cc_3983 N_Z_c_5252_n N_A_3400_333#_c_7187_n 0.048455f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_3984 N_Z_c_5252_n N_A_3400_333#_c_7173_n 0.0249366f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_3985 N_Z_c_5638_n N_A_3400_333#_c_7173_n 4.5829e-19 $X=17.71 $Y=1.87 $X2=0
+ $Y2=0
cc_3986 N_Z_c_5267_n N_A_3400_333#_c_7173_n 2.82292e-19 $X=17.64 $Y=3.315 $X2=0
+ $Y2=0
cc_3987 N_Z_c_5250_n N_A_3400_333#_c_7174_n 0.0016886f $X=17.565 $Y=1.87 $X2=0
+ $Y2=0
cc_3988 N_Z_c_5267_n N_A_3400_333#_c_7174_n 0.0123065f $X=17.64 $Y=3.315 $X2=0
+ $Y2=0
cc_3989 N_Z_c_5252_n N_A_3400_333#_c_7175_n 7.67921e-19 $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_3990 N_Z_c_5252_n N_A_3400_333#_c_7212_n 0.0237143f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_3991 N_Z_c_5250_n N_A_3400_333#_c_7167_n 0.0109134f $X=17.565 $Y=1.87 $X2=0
+ $Y2=0
cc_3992 N_Z_c_5637_n N_A_3400_333#_c_7167_n 4.86317e-19 $X=17.855 $Y=1.87 $X2=0
+ $Y2=0
cc_3993 N_Z_c_5638_n N_A_3400_333#_c_7167_n 0.0210951f $X=17.71 $Y=1.87 $X2=0
+ $Y2=0
cc_3994 N_Z_c_5231_n N_A_3400_333#_c_7167_n 0.00468052f $X=17.64 $Y=1.755 $X2=0
+ $Y2=0
cc_3995 N_Z_c_5267_n N_A_3400_333#_c_7167_n 0.00373869f $X=17.64 $Y=3.315 $X2=0
+ $Y2=0
cc_3996 N_Z_c_5252_n N_A_3400_333#_c_7180_n 0.0166619f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_3997 N_Z_c_5637_n N_A_3400_333#_c_7180_n 0.00221246f $X=17.855 $Y=1.87 $X2=0
+ $Y2=0
cc_3998 N_Z_c_5638_n N_A_3400_333#_c_7180_n 0.0240318f $X=17.71 $Y=1.87 $X2=0
+ $Y2=0
cc_3999 N_Z_c_5267_n N_A_3400_333#_c_7180_n 0.00347206f $X=17.64 $Y=3.315 $X2=0
+ $Y2=0
cc_4000 N_Z_c_5252_n N_A_3400_333#_c_7168_n 0.018076f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_4001 N_Z_c_5251_n N_A_3400_591#_M1134_d 0.00197114f $X=17.565 $Y=3.57
+ $X2=-0.19 $Y2=-0.24
cc_4002 N_Z_c_5253_n N_A_3400_591#_M1158_d 0.0058104f $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4003 N_Z_c_5253_n N_A_3400_591#_c_7260_n 0.0237468f $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4004 N_Z_c_5207_n N_A_3400_591#_c_7265_n 0.00930189f $X=17.65 $Y=4.555 $X2=0
+ $Y2=0
cc_4005 N_Z_c_5253_n N_A_3400_591#_c_7261_n 0.018076f $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4006 N_Z_c_5207_n N_A_3400_591#_c_7262_n 0.00468052f $X=17.65 $Y=4.555 $X2=0
+ $Y2=0
cc_4007 N_Z_c_5251_n N_A_3400_591#_c_7262_n 0.0126134f $X=17.565 $Y=3.57 $X2=0
+ $Y2=0
cc_4008 N_Z_c_5663_n N_A_3400_591#_c_7262_n 4.86317e-19 $X=17.855 $Y=3.57 $X2=0
+ $Y2=0
cc_4009 N_Z_c_5647_n N_A_3400_591#_c_7262_n 0.0210951f $X=17.595 $Y=3.42 $X2=0
+ $Y2=0
cc_4010 N_Z_c_5267_n N_A_3400_591#_c_7262_n 0.0161129f $X=17.64 $Y=3.315 $X2=0
+ $Y2=0
cc_4011 N_Z_c_5253_n N_A_3400_591#_c_7270_n 3.53114e-19 $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4012 N_Z_M1134_s N_A_3400_591#_c_7271_n 0.00154628f $X=17.45 $Y=2.955 $X2=0
+ $Y2=0
cc_4013 N_Z_c_5251_n N_A_3400_591#_c_7271_n 0.0225176f $X=17.565 $Y=3.57 $X2=0
+ $Y2=0
cc_4014 N_Z_c_5253_n N_A_3400_591#_c_7271_n 0.0094263f $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4015 N_Z_c_5663_n N_A_3400_591#_c_7271_n 0.0241216f $X=17.855 $Y=3.57 $X2=0
+ $Y2=0
cc_4016 N_Z_c_5647_n N_A_3400_591#_c_7271_n 0.00832432f $X=17.595 $Y=3.42 $X2=0
+ $Y2=0
cc_4017 N_Z_c_5267_n N_A_3400_591#_c_7271_n 0.0115376f $X=17.64 $Y=3.315 $X2=0
+ $Y2=0
cc_4018 N_Z_c_5251_n N_A_3400_591#_c_7263_n 0.0249588f $X=17.565 $Y=3.57 $X2=0
+ $Y2=0
cc_4019 N_Z_c_5647_n N_A_3400_591#_c_7263_n 4.48979e-19 $X=17.595 $Y=3.42 $X2=0
+ $Y2=0
cc_4020 N_Z_c_5267_n N_A_3400_591#_c_7263_n 2.48349e-19 $X=17.64 $Y=3.315 $X2=0
+ $Y2=0
cc_4021 N_Z_c_5253_n N_A_3400_591#_c_7280_n 0.048455f $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4022 N_Z_c_5253_n N_A_3400_591#_c_7274_n 0.0249366f $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4023 N_Z_c_5647_n N_A_3400_591#_c_7274_n 4.5829e-19 $X=17.595 $Y=3.42 $X2=0
+ $Y2=0
cc_4024 N_Z_c_5267_n N_A_3400_591#_c_7274_n 2.75404e-19 $X=17.64 $Y=3.315 $X2=0
+ $Y2=0
cc_4025 N_Z_c_5253_n N_A_3400_591#_c_7275_n 0.0165143f $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4026 N_Z_c_5663_n N_A_3400_591#_c_7275_n 0.00221246f $X=17.855 $Y=3.57 $X2=0
+ $Y2=0
cc_4027 N_Z_c_5647_n N_A_3400_591#_c_7275_n 0.0240318f $X=17.595 $Y=3.42 $X2=0
+ $Y2=0
cc_4028 N_Z_c_5267_n N_A_3400_591#_c_7275_n 0.00349107f $X=17.64 $Y=3.315 $X2=0
+ $Y2=0
cc_4029 N_Z_c_5253_n N_A_3400_591#_c_7308_n 0.0237143f $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4030 N_Z_c_5252_n N_A_3891_297#_M1143_d 0.00580444f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_4031 N_Z_c_5254_n N_A_3891_297#_M1091_d 0.00197114f $X=24.005 $Y=1.87 $X2=0
+ $Y2=0
cc_4032 N_Z_c_5252_n N_A_3891_297#_c_7358_n 0.0237468f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_4033 N_Z_c_5232_n N_A_3891_297#_c_7358_n 0.00930189f $X=21 $Y=1.755 $X2=0
+ $Y2=0
cc_4034 N_Z_c_5252_n N_A_3891_297#_c_7362_n 0.048455f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_4035 N_Z_c_5252_n N_A_3891_297#_c_7388_n 0.0237143f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_4036 N_Z_M1066_s N_A_3891_297#_c_7367_n 0.00154628f $X=20.9 $Y=1.665 $X2=0
+ $Y2=0
cc_4037 N_Z_c_5252_n N_A_3891_297#_c_7367_n 0.00942629f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_4038 N_Z_c_5254_n N_A_3891_297#_c_7367_n 0.0225177f $X=24.005 $Y=1.87 $X2=0
+ $Y2=0
cc_4039 N_Z_c_5706_n N_A_3891_297#_c_7367_n 0.0241216f $X=21.075 $Y=1.87 $X2=0
+ $Y2=0
cc_4040 N_Z_c_5707_n N_A_3891_297#_c_7367_n 0.00835547f $X=20.93 $Y=1.87 $X2=0
+ $Y2=0
cc_4041 N_Z_c_5269_n N_A_3891_297#_c_7367_n 0.0115376f $X=21 $Y=3.315 $X2=0
+ $Y2=0
cc_4042 N_Z_c_5252_n N_A_3891_297#_c_7369_n 0.0249366f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_4043 N_Z_c_5707_n N_A_3891_297#_c_7369_n 4.5829e-19 $X=20.93 $Y=1.87 $X2=0
+ $Y2=0
cc_4044 N_Z_c_5269_n N_A_3891_297#_c_7369_n 2.82292e-19 $X=21 $Y=3.315 $X2=0
+ $Y2=0
cc_4045 N_Z_c_5252_n N_A_3891_297#_c_7370_n 7.67921e-19 $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_4046 N_Z_c_5254_n N_A_3891_297#_c_7353_n 0.0249588f $X=24.005 $Y=1.87 $X2=0
+ $Y2=0
cc_4047 N_Z_c_5707_n N_A_3891_297#_c_7353_n 4.48979e-19 $X=20.93 $Y=1.87 $X2=0
+ $Y2=0
cc_4048 N_Z_c_5269_n N_A_3891_297#_c_7353_n 2.4892e-19 $X=21 $Y=3.315 $X2=0
+ $Y2=0
cc_4049 N_Z_c_5254_n N_A_3891_297#_c_7372_n 0.0016886f $X=24.005 $Y=1.87 $X2=0
+ $Y2=0
cc_4050 N_Z_c_5269_n N_A_3891_297#_c_7372_n 0.0123065f $X=21 $Y=3.315 $X2=0
+ $Y2=0
cc_4051 N_Z_c_5252_n N_A_3891_297#_c_7365_n 0.0166619f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_4052 N_Z_c_5706_n N_A_3891_297#_c_7365_n 0.00221246f $X=21.075 $Y=1.87 $X2=0
+ $Y2=0
cc_4053 N_Z_c_5707_n N_A_3891_297#_c_7365_n 0.0240318f $X=20.93 $Y=1.87 $X2=0
+ $Y2=0
cc_4054 N_Z_c_5269_n N_A_3891_297#_c_7365_n 0.00347206f $X=21 $Y=3.315 $X2=0
+ $Y2=0
cc_4055 N_Z_c_5254_n N_A_3891_297#_c_7354_n 0.0109134f $X=24.005 $Y=1.87 $X2=0
+ $Y2=0
cc_4056 N_Z_c_5706_n N_A_3891_297#_c_7354_n 4.86317e-19 $X=21.075 $Y=1.87 $X2=0
+ $Y2=0
cc_4057 N_Z_c_5707_n N_A_3891_297#_c_7354_n 0.0210951f $X=20.93 $Y=1.87 $X2=0
+ $Y2=0
cc_4058 N_Z_c_5232_n N_A_3891_297#_c_7354_n 0.00468052f $X=21 $Y=1.755 $X2=0
+ $Y2=0
cc_4059 N_Z_c_5269_n N_A_3891_297#_c_7354_n 0.00373869f $X=21 $Y=3.315 $X2=0
+ $Y2=0
cc_4060 N_Z_c_5252_n N_A_3891_297#_c_7355_n 0.018076f $X=20.785 $Y=1.87 $X2=0
+ $Y2=0
cc_4061 N_Z_c_5253_n N_A_3891_591#_M1152_d 0.0058104f $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4062 N_Z_c_5255_n N_A_3891_591#_M1140_s 0.00197114f $X=24.005 $Y=3.57 $X2=0
+ $Y2=0
cc_4063 N_Z_c_5253_n N_A_3891_591#_c_7445_n 0.018076f $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4064 N_Z_c_5208_n N_A_3891_591#_c_7450_n 0.00930189f $X=20.99 $Y=4.555 $X2=0
+ $Y2=0
cc_4065 N_Z_c_5253_n N_A_3891_591#_c_7450_n 0.0237468f $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4066 N_Z_c_5253_n N_A_3891_591#_c_7461_n 3.53114e-19 $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4067 N_Z_c_5208_n N_A_3891_591#_c_7447_n 0.00468052f $X=20.99 $Y=4.555 $X2=0
+ $Y2=0
cc_4068 N_Z_c_5255_n N_A_3891_591#_c_7447_n 0.0126134f $X=24.005 $Y=3.57 $X2=0
+ $Y2=0
cc_4069 N_Z_c_5733_n N_A_3891_591#_c_7447_n 4.86317e-19 $X=21.075 $Y=3.57 $X2=0
+ $Y2=0
cc_4070 N_Z_c_5716_n N_A_3891_591#_c_7447_n 0.0210951f $X=21.045 $Y=3.42 $X2=0
+ $Y2=0
cc_4071 N_Z_c_5269_n N_A_3891_591#_c_7447_n 0.0161129f $X=21 $Y=3.315 $X2=0
+ $Y2=0
cc_4072 N_Z_c_5253_n N_A_3891_591#_c_7456_n 0.048455f $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4073 N_Z_c_5253_n N_A_3891_591#_c_7488_n 0.0237143f $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4074 N_Z_M1006_d N_A_3891_591#_c_7466_n 0.00154628f $X=20.9 $Y=2.955 $X2=0
+ $Y2=0
cc_4075 N_Z_c_5253_n N_A_3891_591#_c_7466_n 0.0094263f $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4076 N_Z_c_5255_n N_A_3891_591#_c_7466_n 0.0225176f $X=24.005 $Y=3.57 $X2=0
+ $Y2=0
cc_4077 N_Z_c_5733_n N_A_3891_591#_c_7466_n 0.0241216f $X=21.075 $Y=3.57 $X2=0
+ $Y2=0
cc_4078 N_Z_c_5716_n N_A_3891_591#_c_7466_n 0.00835547f $X=21.045 $Y=3.42 $X2=0
+ $Y2=0
cc_4079 N_Z_c_5269_n N_A_3891_591#_c_7466_n 0.0115376f $X=21 $Y=3.315 $X2=0
+ $Y2=0
cc_4080 N_Z_c_5253_n N_A_3891_591#_c_7468_n 0.0249366f $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4081 N_Z_c_5716_n N_A_3891_591#_c_7468_n 4.5829e-19 $X=21.045 $Y=3.42 $X2=0
+ $Y2=0
cc_4082 N_Z_c_5269_n N_A_3891_591#_c_7468_n 2.75404e-19 $X=21 $Y=3.315 $X2=0
+ $Y2=0
cc_4083 N_Z_c_5253_n N_A_3891_591#_c_7458_n 0.0165143f $X=20.785 $Y=3.57 $X2=0
+ $Y2=0
cc_4084 N_Z_c_5733_n N_A_3891_591#_c_7458_n 0.00221246f $X=21.075 $Y=3.57 $X2=0
+ $Y2=0
cc_4085 N_Z_c_5716_n N_A_3891_591#_c_7458_n 0.0240318f $X=21.045 $Y=3.42 $X2=0
+ $Y2=0
cc_4086 N_Z_c_5269_n N_A_3891_591#_c_7458_n 0.00349107f $X=21 $Y=3.315 $X2=0
+ $Y2=0
cc_4087 N_Z_c_5255_n N_A_3891_591#_c_7448_n 0.0249588f $X=24.005 $Y=3.57 $X2=0
+ $Y2=0
cc_4088 N_Z_c_5716_n N_A_3891_591#_c_7448_n 4.48979e-19 $X=21.045 $Y=3.42 $X2=0
+ $Y2=0
cc_4089 N_Z_c_5269_n N_A_3891_591#_c_7448_n 2.48349e-19 $X=21 $Y=3.315 $X2=0
+ $Y2=0
cc_4090 N_Z_c_5254_n N_A_4688_333#_M1122_d 0.00197114f $X=24.005 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_4091 N_Z_c_5233_n N_A_4688_333#_c_7542_n 0.00930189f $X=24.08 $Y=1.755 $X2=0
+ $Y2=0
cc_4092 N_Z_M1122_s N_A_4688_333#_c_7543_n 0.00154628f $X=23.89 $Y=1.665 $X2=0
+ $Y2=0
cc_4093 N_Z_c_5254_n N_A_4688_333#_c_7543_n 0.0225177f $X=24.005 $Y=1.87 $X2=0
+ $Y2=0
cc_4094 Z N_A_4688_333#_c_7543_n 0.0241216f $X=24.065 $Y=1.785 $X2=0 $Y2=0
cc_4095 N_Z_c_5777_n N_A_4688_333#_c_7543_n 0.00832432f $X=24.15 $Y=1.87 $X2=0
+ $Y2=0
cc_4096 N_Z_c_5271_n N_A_4688_333#_c_7543_n 0.0115376f $X=24.08 $Y=3.315 $X2=0
+ $Y2=0
cc_4097 N_Z_c_5254_n N_A_4688_333#_c_7538_n 0.0249588f $X=24.005 $Y=1.87 $X2=0
+ $Y2=0
cc_4098 N_Z_c_5777_n N_A_4688_333#_c_7538_n 4.48979e-19 $X=24.15 $Y=1.87 $X2=0
+ $Y2=0
cc_4099 N_Z_c_5271_n N_A_4688_333#_c_7538_n 2.4892e-19 $X=24.08 $Y=3.315 $X2=0
+ $Y2=0
cc_4100 N_Z_c_5777_n N_A_4688_333#_c_7546_n 4.5829e-19 $X=24.15 $Y=1.87 $X2=0
+ $Y2=0
cc_4101 N_Z_c_5271_n N_A_4688_333#_c_7546_n 2.82292e-19 $X=24.08 $Y=3.315 $X2=0
+ $Y2=0
cc_4102 N_Z_c_5254_n N_A_4688_333#_c_7547_n 0.0016886f $X=24.005 $Y=1.87 $X2=0
+ $Y2=0
cc_4103 N_Z_c_5271_n N_A_4688_333#_c_7547_n 0.0123065f $X=24.08 $Y=3.315 $X2=0
+ $Y2=0
cc_4104 N_Z_c_5254_n N_A_4688_333#_c_7540_n 0.0109134f $X=24.005 $Y=1.87 $X2=0
+ $Y2=0
cc_4105 Z N_A_4688_333#_c_7540_n 4.86317e-19 $X=24.065 $Y=1.785 $X2=0 $Y2=0
cc_4106 N_Z_c_5777_n N_A_4688_333#_c_7540_n 0.0210951f $X=24.15 $Y=1.87 $X2=0
+ $Y2=0
cc_4107 N_Z_c_5233_n N_A_4688_333#_c_7540_n 0.00468052f $X=24.08 $Y=1.755 $X2=0
+ $Y2=0
cc_4108 N_Z_c_5271_n N_A_4688_333#_c_7540_n 0.00373869f $X=24.08 $Y=3.315 $X2=0
+ $Y2=0
cc_4109 Z N_A_4688_333#_c_7553_n 0.0062686f $X=24.065 $Y=1.785 $X2=0 $Y2=0
cc_4110 N_Z_c_5777_n N_A_4688_333#_c_7553_n 0.0233693f $X=24.15 $Y=1.87 $X2=0
+ $Y2=0
cc_4111 N_Z_c_5271_n N_A_4688_333#_c_7553_n 0.00347206f $X=24.08 $Y=3.315 $X2=0
+ $Y2=0
cc_4112 N_Z_c_5255_n N_A_4688_591#_M1049_d 0.00197114f $X=24.005 $Y=3.57
+ $X2=-0.19 $Y2=-0.24
cc_4113 N_Z_c_5209_n N_A_4688_591#_c_7622_n 0.00930189f $X=24.09 $Y=4.555 $X2=0
+ $Y2=0
cc_4114 N_Z_c_5209_n N_A_4688_591#_c_7619_n 0.00468052f $X=24.09 $Y=4.555 $X2=0
+ $Y2=0
cc_4115 N_Z_c_5255_n N_A_4688_591#_c_7619_n 0.0126134f $X=24.005 $Y=3.57 $X2=0
+ $Y2=0
cc_4116 Z N_A_4688_591#_c_7619_n 4.86317e-19 $X=24.065 $Y=3.485 $X2=0 $Y2=0
cc_4117 N_Z_c_5786_n N_A_4688_591#_c_7619_n 0.0210951f $X=24.035 $Y=3.42 $X2=0
+ $Y2=0
cc_4118 N_Z_c_5271_n N_A_4688_591#_c_7619_n 0.0161129f $X=24.08 $Y=3.315 $X2=0
+ $Y2=0
cc_4119 N_Z_M1049_s N_A_4688_591#_c_7628_n 0.00154628f $X=23.89 $Y=2.955 $X2=0
+ $Y2=0
cc_4120 N_Z_c_5255_n N_A_4688_591#_c_7628_n 0.0225176f $X=24.005 $Y=3.57 $X2=0
+ $Y2=0
cc_4121 Z N_A_4688_591#_c_7628_n 0.0241216f $X=24.065 $Y=3.485 $X2=0 $Y2=0
cc_4122 N_Z_c_5786_n N_A_4688_591#_c_7628_n 0.00832432f $X=24.035 $Y=3.42 $X2=0
+ $Y2=0
cc_4123 N_Z_c_5271_n N_A_4688_591#_c_7628_n 0.0115376f $X=24.08 $Y=3.315 $X2=0
+ $Y2=0
cc_4124 N_Z_c_5255_n N_A_4688_591#_c_7620_n 0.0249588f $X=24.005 $Y=3.57 $X2=0
+ $Y2=0
cc_4125 N_Z_c_5786_n N_A_4688_591#_c_7620_n 4.48979e-19 $X=24.035 $Y=3.42 $X2=0
+ $Y2=0
cc_4126 N_Z_c_5271_n N_A_4688_591#_c_7620_n 2.48349e-19 $X=24.08 $Y=3.315 $X2=0
+ $Y2=0
cc_4127 N_Z_c_5786_n N_A_4688_591#_c_7631_n 4.5829e-19 $X=24.035 $Y=3.42 $X2=0
+ $Y2=0
cc_4128 N_Z_c_5271_n N_A_4688_591#_c_7631_n 2.75404e-19 $X=24.08 $Y=3.315 $X2=0
+ $Y2=0
cc_4129 Z N_A_4688_591#_c_7632_n 0.0062686f $X=24.065 $Y=3.485 $X2=0 $Y2=0
cc_4130 N_Z_c_5786_n N_A_4688_591#_c_7632_n 0.0233693f $X=24.035 $Y=3.42 $X2=0
+ $Y2=0
cc_4131 N_Z_c_5271_n N_A_4688_591#_c_7632_n 0.00349107f $X=24.08 $Y=3.315 $X2=0
+ $Y2=0
cc_4132 N_Z_c_5210_n N_A_27_47#_c_7692_n 0.00729487f $X=1.67 $Y=0.68 $X2=0 $Y2=0
cc_4133 N_Z_c_5226_n N_A_27_47#_c_7692_n 0.00238404f $X=1.68 $Y=1.755 $X2=0
+ $Y2=0
cc_4134 N_Z_M1032_s N_A_27_47#_c_7694_n 0.00165831f $X=1.535 $Y=0.345 $X2=0
+ $Y2=0
cc_4135 N_Z_c_5210_n N_A_27_47#_c_7694_n 0.0156951f $X=1.67 $Y=0.68 $X2=0 $Y2=0
cc_4136 N_Z_c_5202_n N_A_27_911#_c_7734_n 0.00238404f $X=1.67 $Y=4.555 $X2=0
+ $Y2=0
cc_4137 N_Z_c_5211_n N_A_27_911#_c_7734_n 0.00729487f $X=1.67 $Y=4.76 $X2=0
+ $Y2=0
cc_4138 N_Z_M1020_s N_A_27_911#_c_7735_n 0.00165831f $X=1.535 $Y=4.575 $X2=0
+ $Y2=0
cc_4139 N_Z_c_5211_n N_A_27_911#_c_7735_n 0.0156951f $X=1.67 $Y=4.76 $X2=0 $Y2=0
cc_4140 N_Z_M1028_s N_A_845_69#_c_8339_n 0.00165831f $X=4.635 $Y=0.345 $X2=0
+ $Y2=0
cc_4141 N_Z_c_5212_n N_A_845_69#_c_8339_n 0.0156951f $X=4.77 $Y=0.68 $X2=0 $Y2=0
cc_4142 N_Z_c_5212_n N_A_845_69#_c_8342_n 0.00729487f $X=4.77 $Y=0.68 $X2=0
+ $Y2=0
cc_4143 N_Z_c_5227_n N_A_845_69#_c_8342_n 0.00238404f $X=4.76 $Y=1.755 $X2=0
+ $Y2=0
cc_4144 N_Z_M1048_d N_A_845_915#_c_8387_n 0.00165831f $X=4.635 $Y=4.575 $X2=0
+ $Y2=0
cc_4145 N_Z_c_5213_n N_A_845_915#_c_8387_n 0.0156951f $X=4.77 $Y=4.76 $X2=0
+ $Y2=0
cc_4146 N_Z_c_5203_n N_A_845_915#_c_8389_n 0.00238404f $X=4.77 $Y=4.555 $X2=0
+ $Y2=0
cc_4147 N_Z_c_5213_n N_A_845_915#_c_8389_n 0.00729487f $X=4.77 $Y=4.76 $X2=0
+ $Y2=0
cc_4148 N_Z_c_5214_n N_A_1315_47#_c_8434_n 0.00729487f $X=8.11 $Y=0.68 $X2=0
+ $Y2=0
cc_4149 N_Z_c_5228_n N_A_1315_47#_c_8434_n 0.00238404f $X=8.12 $Y=1.755 $X2=0
+ $Y2=0
cc_4150 N_Z_M1116_d N_A_1315_47#_c_8436_n 0.00165831f $X=7.975 $Y=0.345 $X2=0
+ $Y2=0
cc_4151 N_Z_c_5214_n N_A_1315_47#_c_8436_n 0.0156951f $X=8.11 $Y=0.68 $X2=0
+ $Y2=0
cc_4152 N_Z_c_5204_n N_A_1315_911#_c_8478_n 0.00238404f $X=8.11 $Y=4.555 $X2=0
+ $Y2=0
cc_4153 N_Z_c_5215_n N_A_1315_911#_c_8478_n 0.00729487f $X=8.11 $Y=4.76 $X2=0
+ $Y2=0
cc_4154 N_Z_M1015_d N_A_1315_911#_c_8479_n 0.00165831f $X=7.975 $Y=4.575 $X2=0
+ $Y2=0
cc_4155 N_Z_c_5215_n N_A_1315_911#_c_8479_n 0.0156951f $X=8.11 $Y=4.76 $X2=0
+ $Y2=0
cc_4156 N_Z_M1102_d N_A_2133_69#_c_8522_n 0.00165831f $X=11.075 $Y=0.345 $X2=0
+ $Y2=0
cc_4157 N_Z_c_5216_n N_A_2133_69#_c_8522_n 0.0156951f $X=11.21 $Y=0.68 $X2=0
+ $Y2=0
cc_4158 N_Z_c_5216_n N_A_2133_69#_c_8525_n 0.00729487f $X=11.21 $Y=0.68 $X2=0
+ $Y2=0
cc_4159 N_Z_c_5229_n N_A_2133_69#_c_8525_n 0.00238404f $X=11.2 $Y=1.755 $X2=0
+ $Y2=0
cc_4160 N_Z_M1029_d N_A_2133_915#_c_8570_n 0.00165831f $X=11.075 $Y=4.575 $X2=0
+ $Y2=0
cc_4161 N_Z_c_5217_n N_A_2133_915#_c_8570_n 0.0156951f $X=11.21 $Y=4.76 $X2=0
+ $Y2=0
cc_4162 N_Z_c_5205_n N_A_2133_915#_c_8572_n 0.00238404f $X=11.21 $Y=4.555 $X2=0
+ $Y2=0
cc_4163 N_Z_c_5217_n N_A_2133_915#_c_8572_n 0.00729487f $X=11.21 $Y=4.76 $X2=0
+ $Y2=0
cc_4164 N_Z_c_5218_n N_A_2603_47#_c_8617_n 0.00729487f $X=14.55 $Y=0.68 $X2=0
+ $Y2=0
cc_4165 N_Z_c_5230_n N_A_2603_47#_c_8617_n 0.00238404f $X=14.56 $Y=1.755 $X2=0
+ $Y2=0
cc_4166 N_Z_M1046_d N_A_2603_47#_c_8619_n 0.00165831f $X=14.415 $Y=0.345 $X2=0
+ $Y2=0
cc_4167 N_Z_c_5218_n N_A_2603_47#_c_8619_n 0.0156951f $X=14.55 $Y=0.68 $X2=0
+ $Y2=0
cc_4168 N_Z_c_5206_n N_A_2603_911#_c_8661_n 0.00238404f $X=14.55 $Y=4.555 $X2=0
+ $Y2=0
cc_4169 N_Z_c_5219_n N_A_2603_911#_c_8661_n 0.00729487f $X=14.55 $Y=4.76 $X2=0
+ $Y2=0
cc_4170 N_Z_M1000_s N_A_2603_911#_c_8662_n 0.00165831f $X=14.415 $Y=4.575 $X2=0
+ $Y2=0
cc_4171 N_Z_c_5219_n N_A_2603_911#_c_8662_n 0.0156951f $X=14.55 $Y=4.76 $X2=0
+ $Y2=0
cc_4172 N_Z_M1022_d N_A_3421_69#_c_8705_n 0.00165831f $X=17.515 $Y=0.345 $X2=0
+ $Y2=0
cc_4173 N_Z_c_5220_n N_A_3421_69#_c_8705_n 0.0156951f $X=17.65 $Y=0.68 $X2=0
+ $Y2=0
cc_4174 N_Z_c_5220_n N_A_3421_69#_c_8708_n 0.00729487f $X=17.65 $Y=0.68 $X2=0
+ $Y2=0
cc_4175 N_Z_c_5231_n N_A_3421_69#_c_8708_n 0.00238404f $X=17.64 $Y=1.755 $X2=0
+ $Y2=0
cc_4176 N_Z_M1016_s N_A_3421_915#_c_8753_n 0.00165831f $X=17.515 $Y=4.575 $X2=0
+ $Y2=0
cc_4177 N_Z_c_5221_n N_A_3421_915#_c_8753_n 0.0156951f $X=17.65 $Y=4.76 $X2=0
+ $Y2=0
cc_4178 N_Z_c_5207_n N_A_3421_915#_c_8755_n 0.00238404f $X=17.65 $Y=4.555 $X2=0
+ $Y2=0
cc_4179 N_Z_c_5221_n N_A_3421_915#_c_8755_n 0.00729487f $X=17.65 $Y=4.76 $X2=0
+ $Y2=0
cc_4180 N_Z_c_5222_n N_A_3891_47#_c_8800_n 0.00729487f $X=20.99 $Y=0.68 $X2=0
+ $Y2=0
cc_4181 N_Z_c_5232_n N_A_3891_47#_c_8800_n 0.00238404f $X=21 $Y=1.755 $X2=0
+ $Y2=0
cc_4182 N_Z_M1112_d N_A_3891_47#_c_8802_n 0.00165831f $X=20.855 $Y=0.345 $X2=0
+ $Y2=0
cc_4183 N_Z_c_5222_n N_A_3891_47#_c_8802_n 0.0156951f $X=20.99 $Y=0.68 $X2=0
+ $Y2=0
cc_4184 N_Z_c_5208_n N_A_3891_911#_c_8844_n 0.00238404f $X=20.99 $Y=4.555 $X2=0
+ $Y2=0
cc_4185 N_Z_c_5223_n N_A_3891_911#_c_8844_n 0.00729487f $X=20.99 $Y=4.76 $X2=0
+ $Y2=0
cc_4186 N_Z_M1021_s N_A_3891_911#_c_8845_n 0.00165831f $X=20.855 $Y=4.575 $X2=0
+ $Y2=0
cc_4187 N_Z_c_5223_n N_A_3891_911#_c_8845_n 0.0156951f $X=20.99 $Y=4.76 $X2=0
+ $Y2=0
cc_4188 N_Z_M1107_d N_A_4709_69#_c_8888_n 0.00165831f $X=23.955 $Y=0.345 $X2=0
+ $Y2=0
cc_4189 N_Z_c_5224_n N_A_4709_69#_c_8888_n 0.0156951f $X=24.09 $Y=0.68 $X2=0
+ $Y2=0
cc_4190 N_Z_c_5224_n N_A_4709_69#_c_8891_n 0.00729487f $X=24.09 $Y=0.68 $X2=0
+ $Y2=0
cc_4191 N_Z_c_5233_n N_A_4709_69#_c_8891_n 0.00238404f $X=24.08 $Y=1.755 $X2=0
+ $Y2=0
cc_4192 N_Z_M1106_d N_A_4709_915#_c_8934_n 0.00165831f $X=23.955 $Y=4.575 $X2=0
+ $Y2=0
cc_4193 N_Z_c_5225_n N_A_4709_915#_c_8934_n 0.0156951f $X=24.09 $Y=4.76 $X2=0
+ $Y2=0
cc_4194 N_Z_c_5209_n N_A_4709_915#_c_8936_n 0.00238404f $X=24.09 $Y=4.555 $X2=0
+ $Y2=0
cc_4195 N_Z_c_5225_n N_A_4709_915#_c_8936_n 0.00729487f $X=24.09 $Y=4.76 $X2=0
+ $Y2=0
cc_4196 N_A_824_333#_c_6418_n N_A_1315_297#_c_6605_n 0.0147157f $X=6.195
+ $Y=1.665 $X2=0 $Y2=0
cc_4197 N_A_824_333#_c_6466_n N_A_1315_297#_c_6642_n 0.0179412f $X=6.18 $Y=2.225
+ $X2=0 $Y2=0
cc_4198 N_A_824_333#_c_6422_n N_A_1315_297#_c_6642_n 9.20345e-19 $X=6.18 $Y=2.21
+ $X2=0 $Y2=0
cc_4199 N_A_824_333#_c_6420_n N_A_1315_297#_c_6606_n 0.0277867f $X=6.18 $Y=2.225
+ $X2=0 $Y2=0
cc_4200 N_A_824_333#_c_6466_n N_A_1315_297#_c_6609_n 9.20345e-19 $X=6.18
+ $Y=2.225 $X2=0 $Y2=0
cc_4201 N_A_824_333#_c_6422_n N_A_1315_297#_c_6609_n 0.0277867f $X=6.18 $Y=2.21
+ $X2=0 $Y2=0
cc_4202 N_A_824_333#_c_6435_n N_A_845_69#_c_8341_n 0.00251701f $X=6.045 $Y=1.58
+ $X2=0 $Y2=0
cc_4203 N_A_824_333#_c_6435_n N_A_845_69#_c_8342_n 0.00200781f $X=6.045 $Y=1.58
+ $X2=0 $Y2=0
cc_4204 N_A_824_333#_c_6423_n N_A_845_69#_c_8342_n 0.00650395f $X=5.325 $Y=1.58
+ $X2=0 $Y2=0
cc_4205 N_A_824_591#_c_6515_n N_A_1315_591#_c_6699_n 0.0277867f $X=6.18 $Y=3.44
+ $X2=0 $Y2=0
cc_4206 N_A_824_591#_c_6514_n N_A_1315_591#_c_6700_n 0.0147157f $X=6.045 $Y=3.86
+ $X2=0 $Y2=0
cc_4207 N_A_824_591#_c_6562_n N_A_1315_591#_c_6742_n 0.0179412f $X=6.18 $Y=3.215
+ $X2=0 $Y2=0
cc_4208 N_A_824_591#_c_6518_n N_A_1315_591#_c_6742_n 9.20345e-19 $X=6.18 $Y=3.1
+ $X2=0 $Y2=0
cc_4209 N_A_824_591#_c_6562_n N_A_1315_591#_c_6703_n 9.20345e-19 $X=6.18
+ $Y=3.215 $X2=0 $Y2=0
cc_4210 N_A_824_591#_c_6518_n N_A_1315_591#_c_6703_n 0.0277867f $X=6.18 $Y=3.1
+ $X2=0 $Y2=0
cc_4211 N_A_824_591#_c_6514_n N_A_845_915#_c_8389_n 0.00200781f $X=6.045 $Y=3.86
+ $X2=0 $Y2=0
cc_4212 N_A_824_591#_c_6519_n N_A_845_915#_c_8389_n 0.00650395f $X=5.325 $Y=3.86
+ $X2=0 $Y2=0
cc_4213 N_A_824_591#_c_6514_n N_A_845_915#_c_8405_n 0.00251701f $X=6.045 $Y=3.86
+ $X2=0 $Y2=0
cc_4214 N_A_1315_297#_c_6612_n N_A_1315_47#_c_8434_n 0.0110288f $X=7.555 $Y=1.58
+ $X2=0 $Y2=0
cc_4215 N_A_1315_591#_c_6704_n N_A_1315_911#_c_8481_n 0.00251701f $X=7.555
+ $Y=3.86 $X2=0 $Y2=0
cc_4216 N_A_1315_591#_c_6704_n N_A_1315_911#_c_8478_n 0.00851176f $X=7.555
+ $Y=3.86 $X2=0 $Y2=0
cc_4217 N_A_2112_333#_c_6791_n N_A_2603_297#_c_6978_n 0.0147157f $X=12.635
+ $Y=1.665 $X2=0 $Y2=0
cc_4218 N_A_2112_333#_c_6839_n N_A_2603_297#_c_7015_n 0.0179412f $X=12.62
+ $Y=2.225 $X2=0 $Y2=0
cc_4219 N_A_2112_333#_c_6795_n N_A_2603_297#_c_7015_n 9.20345e-19 $X=12.62
+ $Y=2.21 $X2=0 $Y2=0
cc_4220 N_A_2112_333#_c_6793_n N_A_2603_297#_c_6979_n 0.0277867f $X=12.62
+ $Y=2.225 $X2=0 $Y2=0
cc_4221 N_A_2112_333#_c_6839_n N_A_2603_297#_c_6982_n 9.20345e-19 $X=12.62
+ $Y=2.225 $X2=0 $Y2=0
cc_4222 N_A_2112_333#_c_6795_n N_A_2603_297#_c_6982_n 0.0277867f $X=12.62
+ $Y=2.21 $X2=0 $Y2=0
cc_4223 N_A_2112_333#_c_6808_n N_A_2133_69#_c_8524_n 0.00251701f $X=12.485
+ $Y=1.58 $X2=0 $Y2=0
cc_4224 N_A_2112_333#_c_6808_n N_A_2133_69#_c_8525_n 0.00200781f $X=12.485
+ $Y=1.58 $X2=0 $Y2=0
cc_4225 N_A_2112_333#_c_6796_n N_A_2133_69#_c_8525_n 0.00650395f $X=11.765
+ $Y=1.58 $X2=0 $Y2=0
cc_4226 N_A_2112_591#_c_6888_n N_A_2603_591#_c_7072_n 0.0277867f $X=12.62
+ $Y=3.44 $X2=0 $Y2=0
cc_4227 N_A_2112_591#_c_6887_n N_A_2603_591#_c_7073_n 0.0147157f $X=12.485
+ $Y=3.86 $X2=0 $Y2=0
cc_4228 N_A_2112_591#_c_6935_n N_A_2603_591#_c_7115_n 0.0179412f $X=12.62
+ $Y=3.215 $X2=0 $Y2=0
cc_4229 N_A_2112_591#_c_6891_n N_A_2603_591#_c_7115_n 9.20345e-19 $X=12.62
+ $Y=3.1 $X2=0 $Y2=0
cc_4230 N_A_2112_591#_c_6935_n N_A_2603_591#_c_7076_n 9.20345e-19 $X=12.62
+ $Y=3.215 $X2=0 $Y2=0
cc_4231 N_A_2112_591#_c_6891_n N_A_2603_591#_c_7076_n 0.0277867f $X=12.62 $Y=3.1
+ $X2=0 $Y2=0
cc_4232 N_A_2112_591#_c_6887_n N_A_2133_915#_c_8572_n 0.00200781f $X=12.485
+ $Y=3.86 $X2=0 $Y2=0
cc_4233 N_A_2112_591#_c_6892_n N_A_2133_915#_c_8572_n 0.00650395f $X=11.765
+ $Y=3.86 $X2=0 $Y2=0
cc_4234 N_A_2112_591#_c_6887_n N_A_2133_915#_c_8588_n 0.00251701f $X=12.485
+ $Y=3.86 $X2=0 $Y2=0
cc_4235 N_A_2603_297#_c_6985_n N_A_2603_47#_c_8617_n 0.0110288f $X=13.995
+ $Y=1.58 $X2=0 $Y2=0
cc_4236 N_A_2603_591#_c_7077_n N_A_2603_911#_c_8664_n 0.00251701f $X=13.995
+ $Y=3.86 $X2=0 $Y2=0
cc_4237 N_A_2603_591#_c_7077_n N_A_2603_911#_c_8661_n 0.00851176f $X=13.995
+ $Y=3.86 $X2=0 $Y2=0
cc_4238 N_A_3400_333#_c_7164_n N_A_3891_297#_c_7351_n 0.0147157f $X=19.075
+ $Y=1.665 $X2=0 $Y2=0
cc_4239 N_A_3400_333#_c_7212_n N_A_3891_297#_c_7388_n 0.0179412f $X=19.06
+ $Y=2.225 $X2=0 $Y2=0
cc_4240 N_A_3400_333#_c_7168_n N_A_3891_297#_c_7388_n 9.20345e-19 $X=19.06
+ $Y=2.21 $X2=0 $Y2=0
cc_4241 N_A_3400_333#_c_7166_n N_A_3891_297#_c_7352_n 0.0277867f $X=19.06
+ $Y=2.225 $X2=0 $Y2=0
cc_4242 N_A_3400_333#_c_7212_n N_A_3891_297#_c_7355_n 9.20345e-19 $X=19.06
+ $Y=2.225 $X2=0 $Y2=0
cc_4243 N_A_3400_333#_c_7168_n N_A_3891_297#_c_7355_n 0.0277867f $X=19.06
+ $Y=2.21 $X2=0 $Y2=0
cc_4244 N_A_3400_333#_c_7181_n N_A_3421_69#_c_8707_n 0.00251701f $X=18.925
+ $Y=1.58 $X2=0 $Y2=0
cc_4245 N_A_3400_333#_c_7181_n N_A_3421_69#_c_8708_n 0.00200781f $X=18.925
+ $Y=1.58 $X2=0 $Y2=0
cc_4246 N_A_3400_333#_c_7169_n N_A_3421_69#_c_8708_n 0.00650395f $X=18.205
+ $Y=1.58 $X2=0 $Y2=0
cc_4247 N_A_3400_591#_c_7261_n N_A_3891_591#_c_7445_n 0.0277867f $X=19.06
+ $Y=3.44 $X2=0 $Y2=0
cc_4248 N_A_3400_591#_c_7260_n N_A_3891_591#_c_7446_n 0.0147157f $X=18.925
+ $Y=3.86 $X2=0 $Y2=0
cc_4249 N_A_3400_591#_c_7308_n N_A_3891_591#_c_7488_n 0.0179412f $X=19.06
+ $Y=3.215 $X2=0 $Y2=0
cc_4250 N_A_3400_591#_c_7264_n N_A_3891_591#_c_7488_n 9.20345e-19 $X=19.06
+ $Y=3.1 $X2=0 $Y2=0
cc_4251 N_A_3400_591#_c_7308_n N_A_3891_591#_c_7449_n 9.20345e-19 $X=19.06
+ $Y=3.215 $X2=0 $Y2=0
cc_4252 N_A_3400_591#_c_7264_n N_A_3891_591#_c_7449_n 0.0277867f $X=19.06 $Y=3.1
+ $X2=0 $Y2=0
cc_4253 N_A_3400_591#_c_7260_n N_A_3421_915#_c_8755_n 0.00200781f $X=18.925
+ $Y=3.86 $X2=0 $Y2=0
cc_4254 N_A_3400_591#_c_7265_n N_A_3421_915#_c_8755_n 0.00650395f $X=18.205
+ $Y=3.86 $X2=0 $Y2=0
cc_4255 N_A_3400_591#_c_7260_n N_A_3421_915#_c_8771_n 0.00251701f $X=18.925
+ $Y=3.86 $X2=0 $Y2=0
cc_4256 N_A_3891_297#_c_7358_n N_A_3891_47#_c_8800_n 0.0110288f $X=20.435
+ $Y=1.58 $X2=0 $Y2=0
cc_4257 N_A_3891_591#_c_7450_n N_A_3891_911#_c_8847_n 0.00251701f $X=20.435
+ $Y=3.86 $X2=0 $Y2=0
cc_4258 N_A_3891_591#_c_7450_n N_A_3891_911#_c_8844_n 0.00851176f $X=20.435
+ $Y=3.86 $X2=0 $Y2=0
cc_4259 N_A_4688_333#_c_7554_n N_A_4709_69#_c_8890_n 0.00251701f $X=25.365
+ $Y=1.58 $X2=0 $Y2=0
cc_4260 N_A_4688_333#_c_7554_n N_A_4709_69#_c_8891_n 0.00200781f $X=25.365
+ $Y=1.58 $X2=0 $Y2=0
cc_4261 N_A_4688_333#_c_7542_n N_A_4709_69#_c_8891_n 0.00650395f $X=24.645
+ $Y=1.58 $X2=0 $Y2=0
cc_4262 N_A_4688_591#_c_7617_n N_A_4709_915#_c_8936_n 0.00200781f $X=25.365
+ $Y=3.86 $X2=0 $Y2=0
cc_4263 N_A_4688_591#_c_7622_n N_A_4709_915#_c_8936_n 0.00650395f $X=24.645
+ $Y=3.86 $X2=0 $Y2=0
cc_4264 N_A_4688_591#_c_7617_n N_A_4709_915#_c_8952_n 0.00251701f $X=25.365
+ $Y=3.86 $X2=0 $Y2=0
cc_4265 N_A_27_47#_c_7692_n N_VGND_M1042_s 0.00306532f $X=1.03 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_4266 N_A_27_47#_c_7692_n N_VGND_c_7777_n 0.012179f $X=1.03 $Y=0.8 $X2=0 $Y2=0
cc_4267 N_A_27_47#_c_7692_n N_VGND_c_7807_n 0.00219745f $X=1.03 $Y=0.8 $X2=0
+ $Y2=0
cc_4268 N_A_27_47#_c_7724_p N_VGND_c_7807_n 0.0199987f $X=1.182 $Y=0.425 $X2=0
+ $Y2=0
cc_4269 N_A_27_47#_c_7694_n N_VGND_c_7807_n 0.0535945f $X=2.005 $Y=0.34 $X2=0
+ $Y2=0
cc_4270 N_A_27_47#_M1042_d VGND 0.00288496f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_4271 N_A_27_47#_M1108_d VGND 0.0024283f $X=1.015 $Y=0.235 $X2=0 $Y2=0
cc_4272 N_A_27_47#_c_7695_n VGND 0.0124017f $X=0.31 $Y=0.38 $X2=0 $Y2=0
cc_4273 N_A_27_47#_c_7692_n VGND 0.00838939f $X=1.03 $Y=0.8 $X2=0 $Y2=0
cc_4274 N_A_27_47#_c_7724_p VGND 0.0117415f $X=1.182 $Y=0.425 $X2=0 $Y2=0
cc_4275 N_A_27_47#_c_7694_n VGND 0.0279432f $X=2.005 $Y=0.34 $X2=0 $Y2=0
cc_4276 N_A_27_47#_c_7695_n N_VGND_c_7837_n 0.020879f $X=0.31 $Y=0.38 $X2=0
+ $Y2=0
cc_4277 N_A_27_47#_c_7692_n N_VGND_c_7837_n 0.0020257f $X=1.03 $Y=0.8 $X2=0
+ $Y2=0
cc_4278 N_A_27_911#_c_7737_n N_VGND_M1047_d 0.00306532f $X=1.03 $Y=4.64 $X2=0
+ $Y2=0
cc_4279 N_A_27_911#_c_7737_n N_VGND_c_7778_n 0.012179f $X=1.03 $Y=4.64 $X2=0
+ $Y2=0
cc_4280 N_A_27_911#_c_7737_n N_VGND_c_7809_n 0.00219745f $X=1.03 $Y=4.64 $X2=0
+ $Y2=0
cc_4281 N_A_27_911#_c_7735_n N_VGND_c_7809_n 0.0535945f $X=2.005 $Y=5.1 $X2=0
+ $Y2=0
cc_4282 N_A_27_911#_c_7768_p N_VGND_c_7809_n 0.0199987f $X=1.335 $Y=5.1 $X2=0
+ $Y2=0
cc_4283 N_A_27_911#_M1047_s VGND 0.00288496f $X=0.135 $Y=4.555 $X2=0 $Y2=0
cc_4284 N_A_27_911#_M1118_s VGND 0.0024283f $X=1.015 $Y=4.555 $X2=0 $Y2=0
cc_4285 N_A_27_911#_c_7737_n VGND 0.00838939f $X=1.03 $Y=4.64 $X2=0 $Y2=0
cc_4286 N_A_27_911#_c_7735_n VGND 0.0279432f $X=2.005 $Y=5.1 $X2=0 $Y2=0
cc_4287 N_A_27_911#_c_7768_p VGND 0.0117415f $X=1.335 $Y=5.1 $X2=0 $Y2=0
cc_4288 N_A_27_911#_c_7736_n VGND 0.0124017f $X=0.31 $Y=4.72 $X2=0 $Y2=0
cc_4289 N_A_27_911#_c_7737_n N_VGND_c_7838_n 0.0020257f $X=1.03 $Y=4.64 $X2=0
+ $Y2=0
cc_4290 N_A_27_911#_c_7736_n N_VGND_c_7838_n 0.020879f $X=0.31 $Y=4.72 $X2=0
+ $Y2=0
cc_4291 VGND N_A_845_69#_M1037_d 0.0024283f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4292 VGND N_A_845_69#_M1105_s 0.00288496f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4293 VGND N_A_845_69#_c_8339_n 0.0222193f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4294 N_VGND_c_7829_n N_A_845_69#_c_8339_n 0.0422314f $X=5.58 $Y=0 $X2=0 $Y2=0
cc_4295 VGND N_A_845_69#_c_8340_n 0.00572388f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4296 N_VGND_c_7829_n N_A_845_69#_c_8340_n 0.0113631f $X=5.58 $Y=0 $X2=0 $Y2=0
cc_4297 VGND N_A_845_69#_c_8376_n 0.0117415f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4298 N_VGND_c_7829_n N_A_845_69#_c_8376_n 0.0199987f $X=5.58 $Y=0 $X2=0 $Y2=0
cc_4299 N_VGND_M1074_d N_A_845_69#_c_8341_n 0.00306532f $X=5.575 $Y=0.235 $X2=0
+ $Y2=0
cc_4300 N_VGND_c_7781_n N_A_845_69#_c_8341_n 0.012179f $X=5.71 $Y=0.38 $X2=0
+ $Y2=0
cc_4301 N_VGND_c_7783_n N_A_845_69#_c_8341_n 0.0020257f $X=7.085 $Y=0 $X2=0
+ $Y2=0
cc_4302 VGND N_A_845_69#_c_8341_n 0.00838939f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4303 N_VGND_c_7829_n N_A_845_69#_c_8341_n 0.00219745f $X=5.58 $Y=0 $X2=0
+ $Y2=0
cc_4304 N_VGND_c_7783_n N_A_845_69#_c_8361_n 0.020879f $X=7.085 $Y=0 $X2=0 $Y2=0
cc_4305 VGND N_A_845_69#_c_8361_n 0.0124017f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4306 VGND N_A_845_915#_M1130_s 0.0024283f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4307 VGND N_A_845_915#_M1059_s 0.00288496f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4308 VGND N_A_845_915#_c_8387_n 0.0339608f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4309 N_VGND_c_7830_n N_A_845_915#_c_8387_n 0.0622301f $X=5.58 $Y=5.44 $X2=0
+ $Y2=0
cc_4310 VGND N_A_845_915#_c_8388_n 0.00572388f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4311 N_VGND_c_7830_n N_A_845_915#_c_8388_n 0.0113631f $X=5.58 $Y=5.44 $X2=0
+ $Y2=0
cc_4312 N_VGND_M1026_d N_A_845_915#_c_8405_n 0.00306532f $X=5.575 $Y=4.555 $X2=0
+ $Y2=0
cc_4313 N_VGND_c_7782_n N_A_845_915#_c_8405_n 0.012179f $X=5.71 $Y=5.06 $X2=0
+ $Y2=0
cc_4314 N_VGND_c_7784_n N_A_845_915#_c_8405_n 0.0020257f $X=7.085 $Y=5.44 $X2=0
+ $Y2=0
cc_4315 VGND N_A_845_915#_c_8405_n 0.00838939f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4316 N_VGND_c_7830_n N_A_845_915#_c_8405_n 0.00219745f $X=5.58 $Y=5.44 $X2=0
+ $Y2=0
cc_4317 N_VGND_c_7784_n N_A_845_915#_c_8390_n 0.020879f $X=7.085 $Y=5.44 $X2=0
+ $Y2=0
cc_4318 VGND N_A_845_915#_c_8390_n 0.0124017f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4319 VGND N_A_1315_47#_M1117_d 0.00288496f $X=25.445 $Y=-0.085 $X2=-0.19
+ $Y2=-0.24
cc_4320 VGND N_A_1315_47#_M1127_d 0.0024283f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4321 N_VGND_c_7783_n N_A_1315_47#_c_8437_n 0.020879f $X=7.085 $Y=0 $X2=0
+ $Y2=0
cc_4322 VGND N_A_1315_47#_c_8437_n 0.0124017f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4323 N_VGND_M1117_s N_A_1315_47#_c_8434_n 0.00306532f $X=7.035 $Y=0.235 $X2=0
+ $Y2=0
cc_4324 N_VGND_c_7783_n N_A_1315_47#_c_8434_n 0.0020257f $X=7.085 $Y=0 $X2=0
+ $Y2=0
cc_4325 N_VGND_c_7785_n N_A_1315_47#_c_8434_n 0.012179f $X=7.17 $Y=0.38 $X2=0
+ $Y2=0
cc_4326 N_VGND_c_7811_n N_A_1315_47#_c_8434_n 0.00219745f $X=9.535 $Y=0 $X2=0
+ $Y2=0
cc_4327 VGND N_A_1315_47#_c_8434_n 0.00838939f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4328 N_VGND_c_7811_n N_A_1315_47#_c_8472_n 0.0199987f $X=9.535 $Y=0 $X2=0
+ $Y2=0
cc_4329 VGND N_A_1315_47#_c_8472_n 0.0117415f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4330 N_VGND_c_7811_n N_A_1315_47#_c_8436_n 0.0535945f $X=9.535 $Y=0 $X2=0
+ $Y2=0
cc_4331 VGND N_A_1315_47#_c_8436_n 0.0279432f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4332 VGND N_A_1315_911#_M1035_d 0.00288496f $X=25.445 $Y=5.355 $X2=-0.19
+ $Y2=-0.24
cc_4333 VGND N_A_1315_911#_M1109_d 0.0024283f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4334 N_VGND_M1035_s N_A_1315_911#_c_8481_n 0.00306532f $X=7.035 $Y=4.555
+ $X2=0 $Y2=0
cc_4335 N_VGND_c_7784_n N_A_1315_911#_c_8481_n 0.0020257f $X=7.085 $Y=5.44 $X2=0
+ $Y2=0
cc_4336 N_VGND_c_7786_n N_A_1315_911#_c_8481_n 0.012179f $X=7.17 $Y=5.06 $X2=0
+ $Y2=0
cc_4337 N_VGND_c_7813_n N_A_1315_911#_c_8481_n 0.00219745f $X=9.535 $Y=5.44
+ $X2=0 $Y2=0
cc_4338 VGND N_A_1315_911#_c_8481_n 0.00838939f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4339 N_VGND_c_7813_n N_A_1315_911#_c_8479_n 0.0535945f $X=9.535 $Y=5.44 $X2=0
+ $Y2=0
cc_4340 VGND N_A_1315_911#_c_8479_n 0.0279432f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4341 N_VGND_c_7813_n N_A_1315_911#_c_8517_n 0.0199987f $X=9.535 $Y=5.44 $X2=0
+ $Y2=0
cc_4342 VGND N_A_1315_911#_c_8517_n 0.0117415f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4343 N_VGND_c_7784_n N_A_1315_911#_c_8480_n 0.020879f $X=7.085 $Y=5.44 $X2=0
+ $Y2=0
cc_4344 VGND N_A_1315_911#_c_8480_n 0.0124017f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4345 VGND N_A_2133_69#_M1125_s 0.0024283f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4346 VGND N_A_2133_69#_M1156_d 0.00288496f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4347 VGND N_A_2133_69#_c_8522_n 0.0222193f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4348 N_VGND_c_7831_n N_A_2133_69#_c_8522_n 0.0422314f $X=12.02 $Y=0 $X2=0
+ $Y2=0
cc_4349 VGND N_A_2133_69#_c_8523_n 0.00572388f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4350 N_VGND_c_7831_n N_A_2133_69#_c_8523_n 0.0113631f $X=12.02 $Y=0 $X2=0
+ $Y2=0
cc_4351 VGND N_A_2133_69#_c_8559_n 0.0117415f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4352 N_VGND_c_7831_n N_A_2133_69#_c_8559_n 0.0199987f $X=12.02 $Y=0 $X2=0
+ $Y2=0
cc_4353 N_VGND_M1025_s N_A_2133_69#_c_8524_n 0.00306532f $X=12.015 $Y=0.235
+ $X2=0 $Y2=0
cc_4354 N_VGND_c_7789_n N_A_2133_69#_c_8524_n 0.012179f $X=12.15 $Y=0.38 $X2=0
+ $Y2=0
cc_4355 N_VGND_c_7791_n N_A_2133_69#_c_8524_n 0.0020257f $X=13.525 $Y=0 $X2=0
+ $Y2=0
cc_4356 VGND N_A_2133_69#_c_8524_n 0.00838939f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4357 N_VGND_c_7831_n N_A_2133_69#_c_8524_n 0.00219745f $X=12.02 $Y=0 $X2=0
+ $Y2=0
cc_4358 N_VGND_c_7791_n N_A_2133_69#_c_8544_n 0.020879f $X=13.525 $Y=0 $X2=0
+ $Y2=0
cc_4359 VGND N_A_2133_69#_c_8544_n 0.0124017f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4360 VGND N_A_2133_915#_M1067_s 0.0024283f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4361 VGND N_A_2133_915#_M1136_d 0.00288496f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4362 VGND N_A_2133_915#_c_8570_n 0.0339608f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4363 N_VGND_c_7832_n N_A_2133_915#_c_8570_n 0.0622301f $X=12.02 $Y=5.44 $X2=0
+ $Y2=0
cc_4364 VGND N_A_2133_915#_c_8571_n 0.00572388f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4365 N_VGND_c_7832_n N_A_2133_915#_c_8571_n 0.0113631f $X=12.02 $Y=5.44 $X2=0
+ $Y2=0
cc_4366 N_VGND_M1011_s N_A_2133_915#_c_8588_n 0.00306532f $X=12.015 $Y=4.555
+ $X2=0 $Y2=0
cc_4367 N_VGND_c_7790_n N_A_2133_915#_c_8588_n 0.012179f $X=12.15 $Y=5.06 $X2=0
+ $Y2=0
cc_4368 N_VGND_c_7792_n N_A_2133_915#_c_8588_n 0.0020257f $X=13.525 $Y=5.44
+ $X2=0 $Y2=0
cc_4369 VGND N_A_2133_915#_c_8588_n 0.00838939f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4370 N_VGND_c_7832_n N_A_2133_915#_c_8588_n 0.00219745f $X=12.02 $Y=5.44
+ $X2=0 $Y2=0
cc_4371 N_VGND_c_7792_n N_A_2133_915#_c_8573_n 0.020879f $X=13.525 $Y=5.44 $X2=0
+ $Y2=0
cc_4372 VGND N_A_2133_915#_c_8573_n 0.0124017f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4373 VGND N_A_2603_47#_M1057_s 0.00288496f $X=25.445 $Y=-0.085 $X2=-0.19
+ $Y2=-0.24
cc_4374 VGND N_A_2603_47#_M1094_s 0.0024283f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4375 N_VGND_c_7791_n N_A_2603_47#_c_8620_n 0.020879f $X=13.525 $Y=0 $X2=0
+ $Y2=0
cc_4376 VGND N_A_2603_47#_c_8620_n 0.0124017f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4377 N_VGND_M1057_d N_A_2603_47#_c_8617_n 0.00306532f $X=13.475 $Y=0.235
+ $X2=0 $Y2=0
cc_4378 N_VGND_c_7791_n N_A_2603_47#_c_8617_n 0.0020257f $X=13.525 $Y=0 $X2=0
+ $Y2=0
cc_4379 N_VGND_c_7793_n N_A_2603_47#_c_8617_n 0.012179f $X=13.61 $Y=0.38 $X2=0
+ $Y2=0
cc_4380 N_VGND_c_7815_n N_A_2603_47#_c_8617_n 0.00219745f $X=15.975 $Y=0 $X2=0
+ $Y2=0
cc_4381 VGND N_A_2603_47#_c_8617_n 0.00838939f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4382 N_VGND_c_7815_n N_A_2603_47#_c_8655_n 0.0199987f $X=15.975 $Y=0 $X2=0
+ $Y2=0
cc_4383 VGND N_A_2603_47#_c_8655_n 0.0117415f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4384 N_VGND_c_7815_n N_A_2603_47#_c_8619_n 0.0535945f $X=15.975 $Y=0 $X2=0
+ $Y2=0
cc_4385 VGND N_A_2603_47#_c_8619_n 0.0279432f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4386 VGND N_A_2603_911#_M1073_s 0.00288496f $X=25.445 $Y=5.355 $X2=-0.19
+ $Y2=-0.24
cc_4387 VGND N_A_2603_911#_M1103_s 0.0024283f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4388 N_VGND_M1073_d N_A_2603_911#_c_8664_n 0.00306532f $X=13.475 $Y=4.555
+ $X2=0 $Y2=0
cc_4389 N_VGND_c_7792_n N_A_2603_911#_c_8664_n 0.0020257f $X=13.525 $Y=5.44
+ $X2=0 $Y2=0
cc_4390 N_VGND_c_7794_n N_A_2603_911#_c_8664_n 0.012179f $X=13.61 $Y=5.06 $X2=0
+ $Y2=0
cc_4391 N_VGND_c_7817_n N_A_2603_911#_c_8664_n 0.00219745f $X=15.975 $Y=5.44
+ $X2=0 $Y2=0
cc_4392 VGND N_A_2603_911#_c_8664_n 0.00838939f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4393 N_VGND_c_7817_n N_A_2603_911#_c_8662_n 0.0535945f $X=15.975 $Y=5.44
+ $X2=0 $Y2=0
cc_4394 VGND N_A_2603_911#_c_8662_n 0.0279432f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4395 N_VGND_c_7817_n N_A_2603_911#_c_8700_n 0.0199987f $X=15.975 $Y=5.44
+ $X2=0 $Y2=0
cc_4396 VGND N_A_2603_911#_c_8700_n 0.0117415f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4397 N_VGND_c_7792_n N_A_2603_911#_c_8663_n 0.020879f $X=13.525 $Y=5.44 $X2=0
+ $Y2=0
cc_4398 VGND N_A_2603_911#_c_8663_n 0.0124017f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4399 VGND N_A_3421_69#_M1054_s 0.0024283f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4400 VGND N_A_3421_69#_M1110_s 0.00288496f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4401 VGND N_A_3421_69#_c_8705_n 0.0222193f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4402 N_VGND_c_7833_n N_A_3421_69#_c_8705_n 0.0422314f $X=18.46 $Y=0 $X2=0
+ $Y2=0
cc_4403 VGND N_A_3421_69#_c_8706_n 0.00572388f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4404 N_VGND_c_7833_n N_A_3421_69#_c_8706_n 0.0113631f $X=18.46 $Y=0 $X2=0
+ $Y2=0
cc_4405 VGND N_A_3421_69#_c_8742_n 0.0117415f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4406 N_VGND_c_7833_n N_A_3421_69#_c_8742_n 0.0199987f $X=18.46 $Y=0 $X2=0
+ $Y2=0
cc_4407 N_VGND_M1090_d N_A_3421_69#_c_8707_n 0.00306532f $X=18.455 $Y=0.235
+ $X2=0 $Y2=0
cc_4408 N_VGND_c_7797_n N_A_3421_69#_c_8707_n 0.012179f $X=18.59 $Y=0.38 $X2=0
+ $Y2=0
cc_4409 N_VGND_c_7799_n N_A_3421_69#_c_8707_n 0.0020257f $X=19.965 $Y=0 $X2=0
+ $Y2=0
cc_4410 VGND N_A_3421_69#_c_8707_n 0.00838939f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4411 N_VGND_c_7833_n N_A_3421_69#_c_8707_n 0.00219745f $X=18.46 $Y=0 $X2=0
+ $Y2=0
cc_4412 N_VGND_c_7799_n N_A_3421_69#_c_8727_n 0.020879f $X=19.965 $Y=0 $X2=0
+ $Y2=0
cc_4413 VGND N_A_3421_69#_c_8727_n 0.0124017f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4414 VGND N_A_3421_915#_M1146_d 0.0024283f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4415 VGND N_A_3421_915#_M1121_s 0.00288496f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4416 VGND N_A_3421_915#_c_8753_n 0.0339608f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4417 N_VGND_c_7834_n N_A_3421_915#_c_8753_n 0.0622301f $X=18.46 $Y=5.44 $X2=0
+ $Y2=0
cc_4418 VGND N_A_3421_915#_c_8754_n 0.00572388f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4419 N_VGND_c_7834_n N_A_3421_915#_c_8754_n 0.0113631f $X=18.46 $Y=5.44 $X2=0
+ $Y2=0
cc_4420 N_VGND_M1100_d N_A_3421_915#_c_8771_n 0.00306532f $X=18.455 $Y=4.555
+ $X2=0 $Y2=0
cc_4421 N_VGND_c_7798_n N_A_3421_915#_c_8771_n 0.012179f $X=18.59 $Y=5.06 $X2=0
+ $Y2=0
cc_4422 N_VGND_c_7800_n N_A_3421_915#_c_8771_n 0.0020257f $X=19.965 $Y=5.44
+ $X2=0 $Y2=0
cc_4423 VGND N_A_3421_915#_c_8771_n 0.00838939f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4424 N_VGND_c_7834_n N_A_3421_915#_c_8771_n 0.00219745f $X=18.46 $Y=5.44
+ $X2=0 $Y2=0
cc_4425 N_VGND_c_7800_n N_A_3421_915#_c_8756_n 0.020879f $X=19.965 $Y=5.44 $X2=0
+ $Y2=0
cc_4426 VGND N_A_3421_915#_c_8756_n 0.0124017f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4427 VGND N_A_3891_47#_M1139_s 0.00288496f $X=25.445 $Y=-0.085 $X2=-0.19
+ $Y2=-0.24
cc_4428 VGND N_A_3891_47#_M1155_s 0.0024283f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4429 N_VGND_c_7799_n N_A_3891_47#_c_8803_n 0.020879f $X=19.965 $Y=0 $X2=0
+ $Y2=0
cc_4430 VGND N_A_3891_47#_c_8803_n 0.0124017f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4431 N_VGND_M1139_d N_A_3891_47#_c_8800_n 0.00306532f $X=19.915 $Y=0.235
+ $X2=0 $Y2=0
cc_4432 N_VGND_c_7799_n N_A_3891_47#_c_8800_n 0.0020257f $X=19.965 $Y=0 $X2=0
+ $Y2=0
cc_4433 N_VGND_c_7801_n N_A_3891_47#_c_8800_n 0.012179f $X=20.05 $Y=0.38 $X2=0
+ $Y2=0
cc_4434 N_VGND_c_7819_n N_A_3891_47#_c_8800_n 0.00219745f $X=22.415 $Y=0 $X2=0
+ $Y2=0
cc_4435 VGND N_A_3891_47#_c_8800_n 0.00838939f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4436 N_VGND_c_7819_n N_A_3891_47#_c_8838_n 0.0199987f $X=22.415 $Y=0 $X2=0
+ $Y2=0
cc_4437 VGND N_A_3891_47#_c_8838_n 0.0117415f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4438 N_VGND_c_7819_n N_A_3891_47#_c_8802_n 0.0535945f $X=22.415 $Y=0 $X2=0
+ $Y2=0
cc_4439 VGND N_A_3891_47#_c_8802_n 0.0279432f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4440 VGND N_A_3891_911#_M1018_s 0.00288496f $X=25.445 $Y=5.355 $X2=-0.19
+ $Y2=-0.24
cc_4441 VGND N_A_3891_911#_M1119_s 0.0024283f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4442 N_VGND_M1018_d N_A_3891_911#_c_8847_n 0.00306532f $X=19.915 $Y=4.555
+ $X2=0 $Y2=0
cc_4443 N_VGND_c_7800_n N_A_3891_911#_c_8847_n 0.0020257f $X=19.965 $Y=5.44
+ $X2=0 $Y2=0
cc_4444 N_VGND_c_7802_n N_A_3891_911#_c_8847_n 0.012179f $X=20.05 $Y=5.06 $X2=0
+ $Y2=0
cc_4445 N_VGND_c_7821_n N_A_3891_911#_c_8847_n 0.00219745f $X=22.415 $Y=5.44
+ $X2=0 $Y2=0
cc_4446 VGND N_A_3891_911#_c_8847_n 0.00838939f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4447 N_VGND_c_7821_n N_A_3891_911#_c_8845_n 0.0535945f $X=22.415 $Y=5.44
+ $X2=0 $Y2=0
cc_4448 VGND N_A_3891_911#_c_8845_n 0.0279432f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4449 N_VGND_c_7821_n N_A_3891_911#_c_8883_n 0.0199987f $X=22.415 $Y=5.44
+ $X2=0 $Y2=0
cc_4450 VGND N_A_3891_911#_c_8883_n 0.0117415f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4451 N_VGND_c_7800_n N_A_3891_911#_c_8846_n 0.020879f $X=19.965 $Y=5.44 $X2=0
+ $Y2=0
cc_4452 VGND N_A_3891_911#_c_8846_n 0.0124017f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4453 VGND N_A_4709_69#_M1138_s 0.0024283f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4454 VGND N_A_4709_69#_M1050_d 0.00288496f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4455 N_VGND_c_7823_n N_A_4709_69#_c_8888_n 0.0422314f $X=24.9 $Y=0 $X2=0
+ $Y2=0
cc_4456 VGND N_A_4709_69#_c_8888_n 0.0222193f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4457 N_VGND_c_7823_n N_A_4709_69#_c_8889_n 0.0113631f $X=24.9 $Y=0 $X2=0
+ $Y2=0
cc_4458 VGND N_A_4709_69#_c_8889_n 0.00572388f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4459 N_VGND_c_7823_n N_A_4709_69#_c_8925_n 0.0199987f $X=24.9 $Y=0 $X2=0
+ $Y2=0
cc_4460 VGND N_A_4709_69#_c_8925_n 0.0117415f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4461 N_VGND_M1024_s N_A_4709_69#_c_8890_n 0.00306532f $X=24.895 $Y=0.235
+ $X2=0 $Y2=0
cc_4462 N_VGND_c_7805_n N_A_4709_69#_c_8890_n 0.012179f $X=25.03 $Y=0.38 $X2=0
+ $Y2=0
cc_4463 N_VGND_c_7823_n N_A_4709_69#_c_8890_n 0.00219745f $X=24.9 $Y=0 $X2=0
+ $Y2=0
cc_4464 VGND N_A_4709_69#_c_8890_n 0.00838939f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4465 N_VGND_c_7835_n N_A_4709_69#_c_8890_n 0.0020257f $X=25.53 $Y=0 $X2=0
+ $Y2=0
cc_4466 VGND N_A_4709_69#_c_8910_n 0.0124017f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_4467 N_VGND_c_7835_n N_A_4709_69#_c_8910_n 0.020879f $X=25.53 $Y=0 $X2=0
+ $Y2=0
cc_4468 VGND N_A_4709_915#_M1131_s 0.0024283f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4469 VGND N_A_4709_915#_M1154_d 0.00288496f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4470 N_VGND_c_7825_n N_A_4709_915#_c_8934_n 0.0622301f $X=24.9 $Y=5.44 $X2=0
+ $Y2=0
cc_4471 VGND N_A_4709_915#_c_8934_n 0.0339608f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4472 N_VGND_c_7825_n N_A_4709_915#_c_8935_n 0.0113631f $X=24.9 $Y=5.44 $X2=0
+ $Y2=0
cc_4473 VGND N_A_4709_915#_c_8935_n 0.00572388f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4474 N_VGND_M1147_s N_A_4709_915#_c_8952_n 0.00306532f $X=24.895 $Y=4.555
+ $X2=0 $Y2=0
cc_4475 N_VGND_c_7806_n N_A_4709_915#_c_8952_n 0.012179f $X=25.03 $Y=5.06 $X2=0
+ $Y2=0
cc_4476 N_VGND_c_7825_n N_A_4709_915#_c_8952_n 0.00219745f $X=24.9 $Y=5.44 $X2=0
+ $Y2=0
cc_4477 VGND N_A_4709_915#_c_8952_n 0.00838939f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4478 N_VGND_c_7836_n N_A_4709_915#_c_8952_n 0.0020257f $X=25.53 $Y=5.44 $X2=0
+ $Y2=0
cc_4479 VGND N_A_4709_915#_c_8937_n 0.0124017f $X=25.445 $Y=5.355 $X2=0 $Y2=0
cc_4480 N_VGND_c_7836_n N_A_4709_915#_c_8937_n 0.020879f $X=25.53 $Y=5.44 $X2=0
+ $Y2=0
cc_4481 N_A_845_69#_c_8361_n N_A_1315_47#_c_8437_n 0.0248576f $X=6.13 $Y=0.38
+ $X2=0 $Y2=0
cc_4482 N_A_845_69#_c_8341_n N_A_1315_47#_c_8435_n 0.0103099f $X=5.965 $Y=0.8
+ $X2=0 $Y2=0
cc_4483 N_A_845_915#_c_8390_n N_A_1315_911#_c_8480_n 0.0351675f $X=6.13 $Y=4.72
+ $X2=0 $Y2=0
cc_4484 N_A_2133_69#_c_8544_n N_A_2603_47#_c_8620_n 0.0248576f $X=12.57 $Y=0.38
+ $X2=0 $Y2=0
cc_4485 N_A_2133_69#_c_8524_n N_A_2603_47#_c_8618_n 0.0103099f $X=12.405 $Y=0.8
+ $X2=0 $Y2=0
cc_4486 N_A_2133_915#_c_8573_n N_A_2603_911#_c_8663_n 0.0351675f $X=12.57
+ $Y=4.72 $X2=0 $Y2=0
cc_4487 N_A_3421_69#_c_8727_n N_A_3891_47#_c_8803_n 0.0248576f $X=19.01 $Y=0.38
+ $X2=0 $Y2=0
cc_4488 N_A_3421_69#_c_8707_n N_A_3891_47#_c_8801_n 0.0103099f $X=18.845 $Y=0.8
+ $X2=0 $Y2=0
cc_4489 N_A_3421_915#_c_8756_n N_A_3891_911#_c_8846_n 0.0351675f $X=19.01
+ $Y=4.72 $X2=0 $Y2=0
