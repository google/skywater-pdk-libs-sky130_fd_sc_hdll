* File: sky130_fd_sc_hdll__buf_4.pex.spice
* Created: Thu Aug 27 19:00:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__BUF_4%A 1 3 6 8
c30 8 0 1.35151e-19 $X=0.235 $Y=1.19
r31 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.305
+ $Y=1.16 $X2=0.305 $Y2=1.16
r32 4 11 36.8497 $w=3.87e-07 $l=2.13528e-07 $layer=POLY_cond $X=0.52 $Y=1.015
+ $X2=0.367 $Y2=1.16
r33 4 6 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.52 $Y=1.015
+ $X2=0.52 $Y2=0.56
r34 1 11 45.0358 $w=3.87e-07 $l=3.07409e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.367 $Y2=1.16
r35 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_4%A_27_47# 1 2 7 9 12 14 16 19 21 23 26 28 30
+ 33 35 37 41 43 44 45 48 50 53 58 66
c111 66 0 1.35151e-19 $X=2.375 $Y=1.217
c112 14 0 1.72053e-19 $X=1.435 $Y=1.41
r113 66 67 3.69632 $w=3.26e-07 $l=2.5e-08 $layer=POLY_cond $X=2.375 $Y=1.217
+ $X2=2.4 $Y2=1.217
r114 65 66 65.7945 $w=3.26e-07 $l=4.45e-07 $layer=POLY_cond $X=1.93 $Y=1.217
+ $X2=2.375 $Y2=1.217
r115 64 65 3.69632 $w=3.26e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.217
+ $X2=1.93 $Y2=1.217
r116 63 64 65.7945 $w=3.26e-07 $l=4.45e-07 $layer=POLY_cond $X=1.46 $Y=1.217
+ $X2=1.905 $Y2=1.217
r117 62 63 3.69632 $w=3.26e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.217
+ $X2=1.46 $Y2=1.217
r118 59 60 3.69632 $w=3.26e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.217
+ $X2=0.99 $Y2=1.217
r119 54 62 60.6196 $w=3.26e-07 $l=4.1e-07 $layer=POLY_cond $X=1.025 $Y=1.217
+ $X2=1.435 $Y2=1.217
r120 54 60 5.17485 $w=3.26e-07 $l=3.5e-08 $layer=POLY_cond $X=1.025 $Y=1.217
+ $X2=0.99 $Y2=1.217
r121 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.025
+ $Y=1.16 $X2=1.025 $Y2=1.16
r122 51 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.86 $Y=1.16
+ $X2=0.775 $Y2=1.16
r123 51 53 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=1.16
+ $X2=1.025 $Y2=1.16
r124 49 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=1.245
+ $X2=0.775 $Y2=1.16
r125 49 50 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.775 $Y=1.245
+ $X2=0.775 $Y2=1.485
r126 48 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=1.075
+ $X2=0.775 $Y2=1.16
r127 47 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.775 $Y=0.905
+ $X2=0.775 $Y2=1.075
r128 46 57 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=1.57
+ $X2=0.26 $Y2=1.57
r129 45 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.69 $Y=1.57
+ $X2=0.775 $Y2=1.485
r130 45 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.69 $Y=1.57
+ $X2=0.425 $Y2=1.57
r131 43 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.69 $Y=0.82
+ $X2=0.775 $Y2=0.905
r132 43 44 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.69 $Y=0.82
+ $X2=0.345 $Y2=0.82
r133 39 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.345 $Y2=0.82
r134 39 41 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.26 $Y2=0.56
r135 35 57 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.655
+ $X2=0.26 $Y2=1.57
r136 35 37 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=0.26 $Y=1.655
+ $X2=0.26 $Y2=2.31
r137 31 67 20.933 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.4 $Y=1.025
+ $X2=2.4 $Y2=1.217
r138 31 33 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.4 $Y=1.025
+ $X2=2.4 $Y2=0.56
r139 28 66 16.6478 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.217
r140 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r141 24 65 20.933 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=1.217
r142 24 26 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=0.56
r143 21 64 16.6478 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.217
r144 21 23 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r145 17 63 20.933 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=1.217
r146 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=0.56
r147 14 62 16.6478 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.217
r148 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r149 10 60 20.933 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=1.217
r150 10 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=0.56
r151 7 59 16.6478 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.217
r152 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r153 2 57 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.63
r154 2 37 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.31
r155 1 41 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_4%VPWR 1 2 3 12 16 20 24 26 28 33 40 41 43 45
+ 48 51
r52 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r53 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r54 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r55 43 45 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.645 $Y=2.72
+ $X2=0.765 $Y2=2.72
r56 41 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r57 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r58 38 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=2.72
+ $X2=2.585 $Y2=2.72
r59 38 40 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.775 $Y=2.72
+ $X2=2.99 $Y2=2.72
r60 37 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r61 37 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r62 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r63 34 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=2.72
+ $X2=1.645 $Y2=2.72
r64 34 36 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.835 $Y=2.72
+ $X2=2.07 $Y2=2.72
r65 33 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=2.72
+ $X2=2.585 $Y2=2.72
r66 33 36 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.395 $Y=2.72
+ $X2=2.07 $Y2=2.72
r67 32 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r68 32 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r70 29 45 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.885 $Y=2.72
+ $X2=0.765 $Y2=2.72
r71 29 31 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.885 $Y=2.72
+ $X2=1.15 $Y2=2.72
r72 28 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.645 $Y2=2.72
r73 28 31 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r74 26 46 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r75 24 43 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=0.235 $Y=2.72
+ $X2=0.645 $Y2=2.72
r76 20 23 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=2.585 $Y=1.66
+ $X2=2.585 $Y2=2.34
r77 18 51 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=2.635
+ $X2=2.585 $Y2=2.72
r78 18 23 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=2.585 $Y=2.635
+ $X2=2.585 $Y2=2.34
r79 14 48 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=2.635
+ $X2=1.645 $Y2=2.72
r80 14 16 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=1.645 $Y=2.635
+ $X2=1.645 $Y2=2
r81 10 45 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.635
+ $X2=0.765 $Y2=2.72
r82 10 12 30.4917 $w=2.38e-07 $l=6.35e-07 $layer=LI1_cond $X=0.765 $Y=2.635
+ $X2=0.765 $Y2=2
r83 3 23 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.34
r84 3 20 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.66
r85 2 16 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2
r86 1 12 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_4%X 1 2 3 4 15 19 21 22 23 24 27 29 30 31 46
c64 29 0 1.72053e-19 $X=2.08 $Y=0.85
r65 31 46 7.5855 $w=2.58e-07 $l=1.4e-07 $layer=LI1_cond $X=2.14 $Y=1.615
+ $X2=2.14 $Y2=1.755
r66 30 31 7.94868 $w=4.73e-07 $l=2.55e-07 $layer=LI1_cond $X=2.072 $Y=1.19
+ $X2=2.072 $Y2=1.445
r67 29 38 3.87901 $w=2.37e-07 $l=8.5e-08 $layer=LI1_cond $X=2.072 $Y=0.82
+ $X2=2.072 $Y2=0.905
r68 29 30 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=2.072 $Y=0.92
+ $X2=2.072 $Y2=1.19
r69 29 38 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=2.072 $Y=0.92
+ $X2=2.072 $Y2=0.905
r70 25 29 3.87901 $w=2.37e-07 $l=1.14039e-07 $layer=LI1_cond $X=2.14 $Y=0.735
+ $X2=2.072 $Y2=0.82
r71 25 27 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.14 $Y=0.735
+ $X2=2.14 $Y2=0.56
r72 23 31 2.57001 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.92 $Y=1.53
+ $X2=2.072 $Y2=1.53
r73 23 24 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.92 $Y=1.53
+ $X2=1.285 $Y2=1.53
r74 21 29 2.57001 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.92 $Y=0.82
+ $X2=2.072 $Y2=0.82
r75 21 22 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.92 $Y=0.82
+ $X2=1.285 $Y2=0.82
r76 17 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=1.285 $Y2=1.53
r77 17 19 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.2 $Y=1.615 $X2=1.2
+ $Y2=1.755
r78 13 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.2 $Y=0.735
+ $X2=1.285 $Y2=0.82
r79 13 15 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.2 $Y=0.735
+ $X2=1.2 $Y2=0.56
r80 4 46 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.755
r81 3 19 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.755
r82 2 27 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.56
r83 1 15 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_4%VGND 1 2 3 12 16 20 22 24 26 32 37 44 45 48
+ 51 54
r54 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r55 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r56 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r57 45 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r58 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r59 42 54 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.585
+ $Y2=0
r60 42 44 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.99
+ $Y2=0
r61 41 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r62 41 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r63 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r64 38 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=1.645
+ $Y2=0
r65 38 40 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=2.07
+ $Y2=0
r66 37 54 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=0 $X2=2.585
+ $Y2=0
r67 37 40 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.395 $Y=0 $X2=2.07
+ $Y2=0
r68 36 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r69 36 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r70 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r71 33 48 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.67
+ $Y2=0
r72 33 35 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=1.15
+ $Y2=0
r73 32 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.645
+ $Y2=0
r74 32 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.15
+ $Y2=0
r75 26 48 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.67
+ $Y2=0
r76 24 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r77 22 26 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=0.525
+ $Y2=0
r78 22 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r79 18 54 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=0.085
+ $X2=2.585 $Y2=0
r80 18 20 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=2.585 $Y=0.085
+ $X2=2.585 $Y2=0.38
r81 14 51 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=0.085
+ $X2=1.645 $Y2=0
r82 14 16 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=1.645 $Y=0.085
+ $X2=1.645 $Y2=0.4
r83 10 48 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0
r84 10 12 12.5179 $w=2.88e-07 $l=3.15e-07 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0.4
r85 3 20 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.475
+ $Y=0.235 $X2=2.61 $Y2=0.38
r86 2 16 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.4
r87 1 12 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.4
.ends

