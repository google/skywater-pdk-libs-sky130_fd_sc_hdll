* File: sky130_fd_sc_hdll__bufinv_8.pex.spice
* Created: Wed Sep  2 08:25:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__BUFINV_8%A 1 3 4 6 7
r22 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r23 4 10 40.2182 $w=4.3e-07 $l=2.38642e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.35 $Y2=1.16
r24 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r25 1 10 44.7166 $w=4.3e-07 $l=3.14245e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.35 $Y2=1.16
r26 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFINV_8%A_117_297# 1 2 9 11 13 16 18 20 21 23 26
+ 30 34 37 42 45 47 48 49 55
c98 42 0 1.39726e-19 $X=2.06 $Y=1.16
c99 26 0 1.25206e-19 $X=2.45 $Y=0.56
c100 21 0 1.26528e-19 $X=2.425 $Y=1.41
r101 55 56 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.425 $Y=1.217
+ $X2=2.45 $Y2=1.217
r102 52 53 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.93 $Y=1.217
+ $X2=1.955 $Y2=1.217
r103 51 52 64.997 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=1.485 $Y=1.217
+ $X2=1.93 $Y2=1.217
r104 50 51 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.46 $Y=1.217
+ $X2=1.485 $Y2=1.217
r105 47 48 6.145 $w=3.78e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.63
+ $X2=0.705 $Y2=1.545
r106 43 55 53.3121 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=2.06 $Y=1.217
+ $X2=2.425 $Y2=1.217
r107 43 53 15.3364 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=2.06 $Y=1.217
+ $X2=1.955 $Y2=1.217
r108 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.06
+ $Y=1.16 $X2=2.06 $Y2=1.16
r109 40 49 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.895 $Y=1.175
+ $X2=0.81 $Y2=1.175
r110 40 42 64.6045 $w=1.98e-07 $l=1.165e-06 $layer=LI1_cond $X=0.895 $Y=1.175
+ $X2=2.06 $Y2=1.175
r111 38 49 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.81 $Y=1.275 $X2=0.81
+ $Y2=1.175
r112 38 48 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.81 $Y=1.275
+ $X2=0.81 $Y2=1.545
r113 37 49 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.81 $Y=1.075 $X2=0.81
+ $Y2=1.175
r114 37 45 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.81 $Y=1.075
+ $X2=0.81 $Y2=0.905
r115 32 47 3.18438 $w=3.78e-07 $l=1.05e-07 $layer=LI1_cond $X=0.705 $Y=1.735
+ $X2=0.705 $Y2=1.63
r116 32 34 17.4383 $w=3.78e-07 $l=5.75e-07 $layer=LI1_cond $X=0.705 $Y=1.735
+ $X2=0.705 $Y2=2.31
r117 28 45 9.32938 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=0.705 $Y=0.715
+ $X2=0.705 $Y2=0.905
r118 28 30 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.705 $Y=0.715
+ $X2=0.705 $Y2=0.4
r119 24 56 21.2229 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.45 $Y=1.025
+ $X2=2.45 $Y2=1.217
r120 24 26 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.45 $Y=1.025
+ $X2=2.45 $Y2=0.56
r121 21 55 16.9318 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.217
r122 21 23 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.985
r123 18 53 16.9318 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.217
r124 18 20 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.985
r125 14 52 21.2229 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=1.217
r126 14 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=0.56
r127 11 51 16.9318 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.217
r128 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.985
r129 7 50 21.2229 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=1.217
r130 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=0.56
r131 2 47 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.63
r132 2 34 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.31
r133 1 30 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFINV_8%A_225_47# 1 2 3 4 15 17 19 22 24 26 29 31
+ 33 36 38 40 43 45 47 50 52 54 57 59 61 62 64 67 71 75 79 80 81 82 85 89 93 95
+ 98 100 106 109 110 111 128
c248 128 0 1.39726e-19 $X=6.185 $Y=1.217
r249 128 129 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=6.185 $Y=1.217
+ $X2=6.21 $Y2=1.217
r250 125 126 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=5.69 $Y=1.217
+ $X2=5.715 $Y2=1.217
r251 124 125 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=5.245 $Y=1.217
+ $X2=5.69 $Y2=1.217
r252 123 124 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=5.22 $Y=1.217
+ $X2=5.245 $Y2=1.217
r253 122 123 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=4.775 $Y=1.217
+ $X2=5.22 $Y2=1.217
r254 121 122 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=4.75 $Y=1.217
+ $X2=4.775 $Y2=1.217
r255 120 121 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=4.305 $Y=1.217
+ $X2=4.75 $Y2=1.217
r256 119 120 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=4.28 $Y=1.217
+ $X2=4.305 $Y2=1.217
r257 118 119 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=3.835 $Y=1.217
+ $X2=4.28 $Y2=1.217
r258 117 118 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=3.81 $Y=1.217
+ $X2=3.835 $Y2=1.217
r259 116 117 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=3.365 $Y=1.217
+ $X2=3.81 $Y2=1.217
r260 115 116 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=3.34 $Y=1.217
+ $X2=3.365 $Y2=1.217
r261 112 113 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=2.87 $Y=1.217
+ $X2=2.895 $Y2=1.217
r262 107 128 17.2143 $w=3.22e-07 $l=1.15e-07 $layer=POLY_cond $X=6.07 $Y=1.217
+ $X2=6.185 $Y2=1.217
r263 107 126 53.1398 $w=3.22e-07 $l=3.55e-07 $layer=POLY_cond $X=6.07 $Y=1.217
+ $X2=5.715 $Y2=1.217
r264 106 107 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=6.07
+ $Y=1.16 $X2=6.07 $Y2=1.16
r265 104 115 50.8944 $w=3.22e-07 $l=3.4e-07 $layer=POLY_cond $X=3 $Y=1.217
+ $X2=3.34 $Y2=1.217
r266 104 113 15.7174 $w=3.22e-07 $l=1.05e-07 $layer=POLY_cond $X=3 $Y=1.217
+ $X2=2.895 $Y2=1.217
r267 103 106 170.245 $w=1.98e-07 $l=3.07e-06 $layer=LI1_cond $X=3 $Y=1.175
+ $X2=6.07 $Y2=1.175
r268 103 104 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=3
+ $Y=1.16 $X2=3 $Y2=1.16
r269 101 111 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=1.175
+ $X2=2.66 $Y2=1.175
r270 101 103 14.1409 $w=1.98e-07 $l=2.55e-07 $layer=LI1_cond $X=2.745 $Y=1.175
+ $X2=3 $Y2=1.175
r271 99 111 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.66 $Y=1.275
+ $X2=2.66 $Y2=1.175
r272 99 100 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.66 $Y=1.275
+ $X2=2.66 $Y2=1.445
r273 98 111 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.66 $Y=1.075
+ $X2=2.66 $Y2=1.175
r274 97 98 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.66 $Y=0.905
+ $X2=2.66 $Y2=1.075
r275 96 110 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.355 $Y=1.53
+ $X2=2.165 $Y2=1.53
r276 95 100 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.575 $Y=1.53
+ $X2=2.66 $Y2=1.445
r277 95 96 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.575 $Y=1.53
+ $X2=2.355 $Y2=1.53
r278 94 109 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.355 $Y=0.82
+ $X2=2.165 $Y2=0.82
r279 93 97 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.575 $Y=0.82
+ $X2=2.66 $Y2=0.905
r280 93 94 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.575 $Y=0.82
+ $X2=2.355 $Y2=0.82
r281 89 91 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=2.165 $Y=1.63
+ $X2=2.165 $Y2=2.31
r282 87 110 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=1.615
+ $X2=2.165 $Y2=1.53
r283 87 89 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=2.165 $Y=1.615
+ $X2=2.165 $Y2=1.63
r284 83 109 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=0.735
+ $X2=2.165 $Y2=0.82
r285 83 85 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.165 $Y=0.735
+ $X2=2.165 $Y2=0.4
r286 81 110 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.975 $Y=1.53
+ $X2=2.165 $Y2=1.53
r287 81 82 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.975 $Y=1.53
+ $X2=1.415 $Y2=1.53
r288 79 109 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.975 $Y=0.82
+ $X2=2.165 $Y2=0.82
r289 79 80 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.975 $Y=0.82
+ $X2=1.415 $Y2=0.82
r290 75 77 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.25 $Y=1.63
+ $X2=1.25 $Y2=2.31
r291 73 82 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.25 $Y=1.615
+ $X2=1.415 $Y2=1.53
r292 73 75 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.25 $Y=1.615
+ $X2=1.25 $Y2=1.63
r293 69 80 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.25 $Y=0.735
+ $X2=1.415 $Y2=0.82
r294 69 71 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.25 $Y=0.735
+ $X2=1.25 $Y2=0.4
r295 65 129 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.21 $Y=1.025
+ $X2=6.21 $Y2=1.217
r296 65 67 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.21 $Y=1.025
+ $X2=6.21 $Y2=0.56
r297 62 128 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.217
r298 62 64 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.985
r299 59 126 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.217
r300 59 61 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.985
r301 55 125 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.69 $Y=1.025
+ $X2=5.69 $Y2=1.217
r302 55 57 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.69 $Y=1.025
+ $X2=5.69 $Y2=0.56
r303 52 124 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.217
r304 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.985
r305 48 123 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.22 $Y=1.025
+ $X2=5.22 $Y2=1.217
r306 48 50 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.22 $Y=1.025
+ $X2=5.22 $Y2=0.56
r307 45 122 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.217
r308 45 47 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
r309 41 121 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.75 $Y=1.025
+ $X2=4.75 $Y2=1.217
r310 41 43 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.75 $Y=1.025
+ $X2=4.75 $Y2=0.56
r311 38 120 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.217
r312 38 40 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.985
r313 34 119 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.28 $Y=1.025
+ $X2=4.28 $Y2=1.217
r314 34 36 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.28 $Y=1.025
+ $X2=4.28 $Y2=0.56
r315 31 118 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.217
r316 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.985
r317 27 117 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.81 $Y=1.025
+ $X2=3.81 $Y2=1.217
r318 27 29 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.81 $Y=1.025
+ $X2=3.81 $Y2=0.56
r319 24 116 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.217
r320 24 26 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.985
r321 20 115 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.34 $Y=1.025
+ $X2=3.34 $Y2=1.217
r322 20 22 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.34 $Y=1.025
+ $X2=3.34 $Y2=0.56
r323 17 113 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.217
r324 17 19 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.985
r325 13 112 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.87 $Y=1.025
+ $X2=2.87 $Y2=1.217
r326 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.87 $Y=1.025
+ $X2=2.87 $Y2=0.56
r327 4 91 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.485 $X2=2.19 $Y2=2.31
r328 4 89 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.485 $X2=2.19 $Y2=1.63
r329 3 77 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.25 $Y2=2.31
r330 3 75 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.25 $Y2=1.63
r331 2 85 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=2.005
+ $Y=0.235 $X2=2.19 $Y2=0.4
r332 1 71 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=1.125
+ $Y=0.235 $X2=1.25 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFINV_8%VPWR 1 2 3 4 5 6 7 22 24 30 34 38 42 46
+ 50 53 54 56 57 59 60 62 63 65 66 68 69 70 95 96
r108 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r109 93 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r110 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r111 90 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r112 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r113 87 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r114 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r115 84 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r116 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r117 81 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r118 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r119 78 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r120 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r121 75 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r122 74 77 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r123 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r124 72 99 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r125 72 74 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r126 70 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r127 70 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r128 68 92 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.335 $Y=2.72
+ $X2=6.21 $Y2=2.72
r129 68 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.335 $Y=2.72
+ $X2=6.42 $Y2=2.72
r130 67 95 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.505 $Y=2.72
+ $X2=6.67 $Y2=2.72
r131 67 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.505 $Y=2.72
+ $X2=6.42 $Y2=2.72
r132 65 89 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=5.395 $Y=2.72
+ $X2=5.29 $Y2=2.72
r133 65 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=2.72
+ $X2=5.48 $Y2=2.72
r134 64 92 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=5.565 $Y=2.72
+ $X2=6.21 $Y2=2.72
r135 64 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=2.72
+ $X2=5.48 $Y2=2.72
r136 62 86 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=2.72
+ $X2=4.37 $Y2=2.72
r137 62 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=2.72
+ $X2=4.54 $Y2=2.72
r138 61 89 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=5.29 $Y2=2.72
r139 61 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=4.54 $Y2=2.72
r140 59 83 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.515 $Y=2.72
+ $X2=3.45 $Y2=2.72
r141 59 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=2.72
+ $X2=3.6 $Y2=2.72
r142 58 86 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=4.37 $Y2=2.72
r143 58 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=3.6 $Y2=2.72
r144 56 80 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.575 $Y=2.72
+ $X2=2.53 $Y2=2.72
r145 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.575 $Y=2.72
+ $X2=2.66 $Y2=2.72
r146 55 83 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.745 $Y=2.72
+ $X2=3.45 $Y2=2.72
r147 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=2.72
+ $X2=2.66 $Y2=2.72
r148 53 77 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.635 $Y=2.72
+ $X2=1.61 $Y2=2.72
r149 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=2.72
+ $X2=1.72 $Y2=2.72
r150 52 80 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=2.53 $Y2=2.72
r151 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=1.72 $Y2=2.72
r152 48 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=2.72
r153 48 50 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=2
r154 44 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2.72
r155 44 46 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2
r156 40 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=2.635
+ $X2=4.54 $Y2=2.72
r157 40 42 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.54 $Y=2.635
+ $X2=4.54 $Y2=2
r158 36 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=2.635 $X2=3.6
+ $Y2=2.72
r159 36 38 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.6 $Y=2.635
+ $X2=3.6 $Y2=2
r160 32 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=2.635
+ $X2=2.66 $Y2=2.72
r161 32 34 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.66 $Y=2.635
+ $X2=2.66 $Y2=2
r162 28 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=2.635
+ $X2=1.72 $Y2=2.72
r163 28 30 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.72 $Y=2.635
+ $X2=1.72 $Y2=2
r164 24 27 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r165 22 99 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.172 $Y2=2.72
r166 22 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r167 7 50 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.275
+ $Y=1.485 $X2=6.42 $Y2=2
r168 6 46 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=2
r169 5 42 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.395
+ $Y=1.485 $X2=4.54 $Y2=2
r170 4 38 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.455
+ $Y=1.485 $X2=3.6 $Y2=2
r171 3 34 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.515
+ $Y=1.485 $X2=2.66 $Y2=2
r172 2 30 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.575
+ $Y=1.485 $X2=1.72 $Y2=2
r173 1 27 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r174 1 24 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFINV_8%Y 1 2 3 4 5 6 7 8 27 31 35 36 37 38 41 45
+ 49 51 55 59 63 65 69 73 77 79 81 82 83 84 85 86 88 89
c179 38 0 1.26528e-19 $X=3.295 $Y=1.53
c180 36 0 1.25206e-19 $X=3.295 $Y=0.82
r181 88 89 6.56111 $w=5.58e-07 $l=2.55e-07 $layer=LI1_cond $X=6.61 $Y=1.19
+ $X2=6.61 $Y2=1.445
r182 87 88 8.4217 $w=3.88e-07 $l=2.85e-07 $layer=LI1_cond $X=6.61 $Y=0.905
+ $X2=6.61 $Y2=1.19
r183 80 86 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.115 $Y=1.53
+ $X2=5.925 $Y2=1.53
r184 79 89 5.76906 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=6.415 $Y=1.53
+ $X2=6.61 $Y2=1.53
r185 79 80 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.415 $Y=1.53
+ $X2=6.115 $Y2=1.53
r186 78 85 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.115 $Y=0.82
+ $X2=5.925 $Y2=0.82
r187 77 87 8.28377 $w=1.7e-07 $l=2.33666e-07 $layer=LI1_cond $X=6.415 $Y=0.82
+ $X2=6.61 $Y2=0.905
r188 77 78 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.415 $Y=0.82
+ $X2=6.115 $Y2=0.82
r189 73 75 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=5.925 $Y=1.63
+ $X2=5.925 $Y2=2.31
r190 71 86 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.925 $Y=1.615
+ $X2=5.925 $Y2=1.53
r191 71 73 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=5.925 $Y=1.615
+ $X2=5.925 $Y2=1.63
r192 67 85 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.925 $Y=0.735
+ $X2=5.925 $Y2=0.82
r193 67 69 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.925 $Y=0.735
+ $X2=5.925 $Y2=0.4
r194 66 84 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.175 $Y=1.53
+ $X2=4.985 $Y2=1.53
r195 65 86 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.735 $Y=1.53
+ $X2=5.925 $Y2=1.53
r196 65 66 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.735 $Y=1.53
+ $X2=5.175 $Y2=1.53
r197 64 83 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.175 $Y=0.82
+ $X2=4.985 $Y2=0.82
r198 63 85 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.735 $Y=0.82
+ $X2=5.925 $Y2=0.82
r199 63 64 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.735 $Y=0.82
+ $X2=5.175 $Y2=0.82
r200 59 61 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=4.985 $Y=1.63
+ $X2=4.985 $Y2=2.31
r201 57 84 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.985 $Y=1.615
+ $X2=4.985 $Y2=1.53
r202 57 59 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=4.985 $Y=1.615
+ $X2=4.985 $Y2=1.63
r203 53 83 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.985 $Y=0.735
+ $X2=4.985 $Y2=0.82
r204 53 55 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.985 $Y=0.735
+ $X2=4.985 $Y2=0.4
r205 52 82 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.235 $Y=1.53
+ $X2=4.045 $Y2=1.53
r206 51 84 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.795 $Y=1.53
+ $X2=4.985 $Y2=1.53
r207 51 52 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.795 $Y=1.53
+ $X2=4.235 $Y2=1.53
r208 50 81 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.235 $Y=0.82
+ $X2=4.045 $Y2=0.82
r209 49 83 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.795 $Y=0.82
+ $X2=4.985 $Y2=0.82
r210 49 50 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.795 $Y=0.82
+ $X2=4.235 $Y2=0.82
r211 45 47 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=4.045 $Y=1.63
+ $X2=4.045 $Y2=2.31
r212 43 82 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=1.615
+ $X2=4.045 $Y2=1.53
r213 43 45 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=4.045 $Y=1.615
+ $X2=4.045 $Y2=1.63
r214 39 81 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=0.735
+ $X2=4.045 $Y2=0.82
r215 39 41 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.045 $Y=0.735
+ $X2=4.045 $Y2=0.4
r216 37 82 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.855 $Y=1.53
+ $X2=4.045 $Y2=1.53
r217 37 38 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.855 $Y=1.53
+ $X2=3.295 $Y2=1.53
r218 35 81 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.855 $Y=0.82
+ $X2=4.045 $Y2=0.82
r219 35 36 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.855 $Y=0.82
+ $X2=3.295 $Y2=0.82
r220 31 33 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=3.105 $Y=1.63
+ $X2=3.105 $Y2=2.31
r221 29 38 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=3.105 $Y=1.615
+ $X2=3.295 $Y2=1.53
r222 29 31 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=3.105 $Y=1.615
+ $X2=3.105 $Y2=1.63
r223 25 36 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=3.105 $Y=0.735
+ $X2=3.295 $Y2=0.82
r224 25 27 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.105 $Y=0.735
+ $X2=3.105 $Y2=0.4
r225 8 75 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=2.31
r226 8 73 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=1.63
r227 7 61 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=2.31
r228 7 59 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=1.63
r229 6 47 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=2.31
r230 6 45 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=1.63
r231 5 33 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=2.985
+ $Y=1.485 $X2=3.13 $Y2=2.31
r232 5 31 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.985
+ $Y=1.485 $X2=3.13 $Y2=1.63
r233 4 69 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=5.765
+ $Y=0.235 $X2=5.95 $Y2=0.4
r234 3 55 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=4.825
+ $Y=0.235 $X2=5.01 $Y2=0.4
r235 2 41 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=3.885
+ $Y=0.235 $X2=4.07 $Y2=0.4
r236 1 27 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=2.945
+ $Y=0.235 $X2=3.13 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFINV_8%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44
+ 48 51 52 54 55 57 58 60 61 63 64 66 67 68 93 94
r115 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r116 91 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r117 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r118 88 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r119 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r120 85 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r121 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r122 82 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r123 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r124 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r125 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r126 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r127 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r128 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r129 72 75 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r130 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r131 70 97 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r132 70 72 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r133 68 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r134 68 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r135 66 90 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.335 $Y=0
+ $X2=6.21 $Y2=0
r136 66 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.335 $Y=0 $X2=6.42
+ $Y2=0
r137 65 93 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.505 $Y=0
+ $X2=6.67 $Y2=0
r138 65 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.505 $Y=0 $X2=6.42
+ $Y2=0
r139 63 87 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=5.395 $Y=0
+ $X2=5.29 $Y2=0
r140 63 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=0 $X2=5.48
+ $Y2=0
r141 62 90 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=5.565 $Y=0
+ $X2=6.21 $Y2=0
r142 62 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=0 $X2=5.48
+ $Y2=0
r143 60 84 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=0 $X2=4.37
+ $Y2=0
r144 60 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=0 $X2=4.54
+ $Y2=0
r145 59 87 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.625 $Y=0 $X2=5.29
+ $Y2=0
r146 59 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=0 $X2=4.54
+ $Y2=0
r147 57 81 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.515 $Y=0 $X2=3.45
+ $Y2=0
r148 57 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=0 $X2=3.6
+ $Y2=0
r149 56 84 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.685 $Y=0
+ $X2=4.37 $Y2=0
r150 56 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.6
+ $Y2=0
r151 54 78 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.575 $Y=0 $X2=2.53
+ $Y2=0
r152 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.575 $Y=0 $X2=2.66
+ $Y2=0
r153 53 81 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.745 $Y=0
+ $X2=3.45 $Y2=0
r154 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.66
+ $Y2=0
r155 51 75 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.635 $Y=0 $X2=1.61
+ $Y2=0
r156 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=0 $X2=1.72
+ $Y2=0
r157 50 78 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.805 $Y=0
+ $X2=2.53 $Y2=0
r158 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.805 $Y=0 $X2=1.72
+ $Y2=0
r159 46 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0
r160 46 48 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0.4
r161 42 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0
r162 42 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.4
r163 38 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0
r164 38 40 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0.4
r165 34 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=0.085 $X2=3.6
+ $Y2=0
r166 34 36 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.6 $Y=0.085
+ $X2=3.6 $Y2=0.4
r167 30 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=0.085
+ $X2=2.66 $Y2=0
r168 30 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.66 $Y=0.085
+ $X2=2.66 $Y2=0.4
r169 26 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=0.085
+ $X2=1.72 $Y2=0
r170 26 28 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.72 $Y=0.085
+ $X2=1.72 $Y2=0.4
r171 22 97 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r172 22 24 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.4
r173 7 48 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=6.285
+ $Y=0.235 $X2=6.42 $Y2=0.4
r174 6 44 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=5.295
+ $Y=0.235 $X2=5.48 $Y2=0.4
r175 5 40 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=4.355
+ $Y=0.235 $X2=4.54 $Y2=0.4
r176 4 36 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.235 $X2=3.6 $Y2=0.4
r177 3 32 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.525
+ $Y=0.235 $X2=2.66 $Y2=0.4
r178 2 28 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.72 $Y2=0.4
r179 1 24 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

