* File: sky130_fd_sc_hdll__a22o_4.pex.spice
* Created: Wed Sep  2 08:18:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A22O_4%A_96_21# 1 2 3 4 13 15 16 18 19 21 22 24 25
+ 27 28 30 31 33 34 36 37 46 48 50 51 52 53 55 56 61 63 65 66 71 72 73 78 87
c169 73 0 1.39491e-19 $X=4.155 $Y=1.87
c170 66 0 1.39491e-19 $X=3.215 $Y=1.87
r171 87 88 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.99 $Y=1.202
+ $X2=2.015 $Y2=1.202
r172 84 85 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.495 $Y=1.202
+ $X2=1.52 $Y2=1.202
r173 83 84 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=1.05 $Y=1.202
+ $X2=1.495 $Y2=1.202
r174 82 83 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.025 $Y=1.202
+ $X2=1.05 $Y2=1.202
r175 79 80 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.555 $Y=1.202
+ $X2=0.58 $Y2=1.202
r176 73 76 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.155 $Y=1.87
+ $X2=4.155 $Y2=1.96
r177 72 78 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=3.905 $Y=0.82
+ $X2=5.385 $Y2=0.82
r178 66 69 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=3.215 $Y=1.87
+ $X2=3.215 $Y2=1.96
r179 61 78 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=5.515 $Y=0.775
+ $X2=5.385 $Y2=0.775
r180 61 63 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=5.515 $Y=0.775
+ $X2=5.645 $Y2=0.775
r181 56 71 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.55 $Y=0.775
+ $X2=3.42 $Y2=0.775
r182 56 58 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=3.55 $Y=0.775
+ $X2=3.685 $Y2=0.775
r183 55 72 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.775 $Y=0.775
+ $X2=3.905 $Y2=0.775
r184 55 58 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=3.775 $Y=0.775
+ $X2=3.685 $Y2=0.775
r185 54 66 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.34 $Y=1.87
+ $X2=3.215 $Y2=1.87
r186 53 73 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.03 $Y=1.87
+ $X2=4.155 $Y2=1.87
r187 53 54 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.03 $Y=1.87
+ $X2=3.34 $Y2=1.87
r188 51 66 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.09 $Y=1.87
+ $X2=3.215 $Y2=1.87
r189 51 52 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=3.09 $Y=1.87
+ $X2=2.43 $Y2=1.87
r190 50 71 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=2.43 $Y=0.82
+ $X2=3.42 $Y2=0.82
r191 48 65 3.53812 $w=3.1e-07 $l=1.09545e-07 $layer=LI1_cond $X=2.285 $Y=1.075
+ $X2=2.265 $Y2=1.175
r192 47 50 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=2.285 $Y=0.905
+ $X2=2.43 $Y2=0.82
r193 47 48 6.7557 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=2.285 $Y=0.905
+ $X2=2.285 $Y2=1.075
r194 46 52 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.265 $Y=1.785
+ $X2=2.43 $Y2=1.87
r195 45 65 3.53812 $w=3.1e-07 $l=1e-07 $layer=LI1_cond $X=2.265 $Y=1.275
+ $X2=2.265 $Y2=1.175
r196 45 46 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=2.265 $Y=1.275
+ $X2=2.265 $Y2=1.785
r197 44 87 14.9005 $w=3.72e-07 $l=1.15e-07 $layer=POLY_cond $X=1.875 $Y=1.202
+ $X2=1.99 $Y2=1.202
r198 44 85 45.9973 $w=3.72e-07 $l=3.55e-07 $layer=POLY_cond $X=1.875 $Y=1.202
+ $X2=1.52 $Y2=1.202
r199 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.875
+ $Y=1.16 $X2=1.875 $Y2=1.16
r200 40 82 41.4624 $w=3.72e-07 $l=3.2e-07 $layer=POLY_cond $X=0.705 $Y=1.202
+ $X2=1.025 $Y2=1.202
r201 40 80 16.1962 $w=3.72e-07 $l=1.25e-07 $layer=POLY_cond $X=0.705 $Y=1.202
+ $X2=0.58 $Y2=1.202
r202 39 43 64.8818 $w=1.98e-07 $l=1.17e-06 $layer=LI1_cond $X=0.705 $Y=1.175
+ $X2=1.875 $Y2=1.175
r203 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.705
+ $Y=1.16 $X2=0.705 $Y2=1.16
r204 37 65 2.95888 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.1 $Y=1.175
+ $X2=2.265 $Y2=1.175
r205 37 43 12.4773 $w=1.98e-07 $l=2.25e-07 $layer=LI1_cond $X=2.1 $Y=1.175
+ $X2=1.875 $Y2=1.175
r206 34 88 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.015 $Y=0.995
+ $X2=2.015 $Y2=1.202
r207 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.015 $Y=0.995
+ $X2=2.015 $Y2=0.56
r208 31 87 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.99 $Y=1.41
+ $X2=1.99 $Y2=1.202
r209 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.99 $Y=1.41
+ $X2=1.99 $Y2=1.985
r210 28 85 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.52 $Y=1.41
+ $X2=1.52 $Y2=1.202
r211 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.52 $Y=1.41
+ $X2=1.52 $Y2=1.985
r212 25 84 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.495 $Y=0.995
+ $X2=1.495 $Y2=1.202
r213 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.495 $Y=0.995
+ $X2=1.495 $Y2=0.56
r214 22 83 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.05 $Y=1.41
+ $X2=1.05 $Y2=1.202
r215 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.05 $Y=1.41
+ $X2=1.05 $Y2=1.985
r216 19 82 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.025 $Y=0.995
+ $X2=1.025 $Y2=1.202
r217 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.025 $Y=0.995
+ $X2=1.025 $Y2=0.56
r218 16 80 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.58 $Y=1.41
+ $X2=0.58 $Y2=1.202
r219 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.58 $Y=1.41
+ $X2=0.58 $Y2=1.985
r220 13 79 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.555 $Y=0.995
+ $X2=0.555 $Y2=1.202
r221 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.555 $Y=0.995
+ $X2=0.555 $Y2=0.56
r222 4 76 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=4.01
+ $Y=1.485 $X2=4.155 $Y2=1.96
r223 3 69 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=3.07
+ $Y=1.485 $X2=3.215 $Y2=1.96
r224 2 63 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=5.46
+ $Y=0.235 $X2=5.645 $Y2=0.73
r225 1 58 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=3.5
+ $Y=0.235 $X2=3.685 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_4%B2 1 3 4 6 7 9 10 12 13 16 21 30
c80 10 0 2.84747e-19 $X=4.39 $Y=1.41
c81 1 0 1.39491e-19 $X=2.98 $Y=1.41
r82 30 32 3.98693 $w=5.83e-07 $l=1.95e-07 $layer=LI1_cond $X=2.912 $Y=1.335
+ $X2=2.912 $Y2=1.53
r83 21 30 3.57801 $w=5.83e-07 $l=1.75e-07 $layer=LI1_cond $X=2.912 $Y=1.16
+ $X2=2.912 $Y2=1.335
r84 21 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.955
+ $Y=1.16 $X2=2.955 $Y2=1.16
r85 16 19 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=4.39 $Y=1.16
+ $X2=4.39 $Y2=1.53
r86 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.365
+ $Y=1.16 $X2=4.365 $Y2=1.16
r87 14 32 8.15384 $w=1.7e-07 $l=2.93e-07 $layer=LI1_cond $X=3.205 $Y=1.53
+ $X2=2.912 $Y2=1.53
r88 13 19 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.2 $Y=1.53 $X2=4.39
+ $Y2=1.53
r89 13 14 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=4.2 $Y=1.53
+ $X2=3.205 $Y2=1.53
r90 10 17 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=4.39 $Y=1.41
+ $X2=4.39 $Y2=1.16
r91 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.39 $Y=1.41
+ $X2=4.39 $Y2=1.985
r92 7 17 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=4.365 $Y=0.995
+ $X2=4.39 $Y2=1.16
r93 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.365 $Y=0.995
+ $X2=4.365 $Y2=0.56
r94 4 24 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=3.005 $Y=0.995
+ $X2=2.98 $Y2=1.16
r95 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.005 $Y=0.995
+ $X2=3.005 $Y2=0.56
r96 1 24 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=2.98 $Y=1.41
+ $X2=2.98 $Y2=1.16
r97 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.98 $Y=1.41 $X2=2.98
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_4%B1 1 3 4 6 7 9 10 12 13 20 25
r45 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.92 $Y=1.202
+ $X2=3.945 $Y2=1.202
r46 19 25 11.0909 $w=1.98e-07 $l=2e-07 $layer=LI1_cond $X=3.685 $Y=1.175
+ $X2=3.885 $Y2=1.175
r47 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=3.685 $Y=1.202
+ $X2=3.92 $Y2=1.202
r48 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.685
+ $Y=1.16 $X2=3.685 $Y2=1.16
r49 16 18 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=3.45 $Y=1.202
+ $X2=3.685 $Y2=1.202
r50 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.425 $Y=1.202
+ $X2=3.45 $Y2=1.202
r51 13 25 1.38636 $w=1.98e-07 $l=2.5e-08 $layer=LI1_cond $X=3.91 $Y=1.175
+ $X2=3.885 $Y2=1.175
r52 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.945 $Y=0.995
+ $X2=3.945 $Y2=1.202
r53 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.945 $Y=0.995
+ $X2=3.945 $Y2=0.56
r54 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.92 $Y=1.41
+ $X2=3.92 $Y2=1.202
r55 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.92 $Y=1.41 $X2=3.92
+ $Y2=1.985
r56 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.45 $Y=1.41
+ $X2=3.45 $Y2=1.202
r57 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.45 $Y=1.41 $X2=3.45
+ $Y2=1.985
r58 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.425 $Y=0.995
+ $X2=3.425 $Y2=1.202
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.425 $Y=0.995
+ $X2=3.425 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_4%A2 1 3 4 6 7 9 10 12 13 16 18 23 24 32
c75 10 0 8.80283e-20 $X=6.375 $Y=0.995
c76 7 0 1.89609e-19 $X=6.35 $Y=1.41
c77 1 0 1.45256e-19 $X=4.94 $Y=1.41
r78 29 32 12.4773 $w=1.98e-07 $l=2.25e-07 $layer=LI1_cond $X=6.325 $Y=1.175
+ $X2=6.55 $Y2=1.175
r79 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.325
+ $Y=1.16 $X2=6.325 $Y2=1.16
r80 24 32 6.1 $w=1.98e-07 $l=1.1e-07 $layer=LI1_cond $X=6.66 $Y=1.175 $X2=6.55
+ $Y2=1.175
r81 23 29 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=6.285 $Y=1.175
+ $X2=6.325 $Y2=1.175
r82 18 21 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=4.94 $Y=1.16
+ $X2=4.94 $Y2=1.53
r83 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.915
+ $Y=1.16 $X2=4.915 $Y2=1.16
r84 15 23 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=6.2 $Y=1.275
+ $X2=6.285 $Y2=1.175
r85 15 16 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.2 $Y=1.275 $X2=6.2
+ $Y2=1.445
r86 14 21 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.13 $Y=1.53 $X2=4.94
+ $Y2=1.53
r87 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.115 $Y=1.53
+ $X2=6.2 $Y2=1.445
r88 13 14 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=6.115 $Y=1.53
+ $X2=5.13 $Y2=1.53
r89 10 28 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=6.375 $Y=0.995
+ $X2=6.35 $Y2=1.16
r90 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.375 $Y=0.995
+ $X2=6.375 $Y2=0.56
r91 7 28 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=6.35 $Y=1.41
+ $X2=6.35 $Y2=1.16
r92 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.35 $Y=1.41 $X2=6.35
+ $Y2=1.985
r93 4 19 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=4.965 $Y=0.995
+ $X2=4.94 $Y2=1.16
r94 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.965 $Y=0.995
+ $X2=4.965 $Y2=0.56
r95 1 19 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=4.94 $Y=1.41
+ $X2=4.94 $Y2=1.16
r96 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.94 $Y=1.41 $X2=4.94
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_4%A1 1 3 4 6 7 9 10 12 13 20 25
c44 13 0 1.89609e-19 $X=5.66 $Y=1.105
c45 10 0 8.25269e-20 $X=5.905 $Y=0.995
r46 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=5.88 $Y=1.202
+ $X2=5.905 $Y2=1.202
r47 19 25 4.99091 $w=1.98e-07 $l=9e-08 $layer=LI1_cond $X=5.645 $Y=1.175
+ $X2=5.735 $Y2=1.175
r48 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=5.645 $Y=1.202
+ $X2=5.88 $Y2=1.202
r49 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.645
+ $Y=1.16 $X2=5.645 $Y2=1.16
r50 16 18 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=5.41 $Y=1.202
+ $X2=5.645 $Y2=1.202
r51 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=5.385 $Y=1.202
+ $X2=5.41 $Y2=1.202
r52 13 25 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=5.745 $Y=1.175
+ $X2=5.735 $Y2=1.175
r53 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.905 $Y=0.995
+ $X2=5.905 $Y2=1.202
r54 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.905 $Y=0.995
+ $X2=5.905 $Y2=0.56
r55 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.88 $Y=1.41
+ $X2=5.88 $Y2=1.202
r56 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.88 $Y=1.41 $X2=5.88
+ $Y2=1.985
r57 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.41 $Y=1.41
+ $X2=5.41 $Y2=1.202
r58 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.41 $Y=1.41 $X2=5.41
+ $Y2=1.985
r59 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.385 $Y=0.995
+ $X2=5.385 $Y2=1.202
r60 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.385 $Y=0.995
+ $X2=5.385 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_4%VPWR 1 2 3 4 5 16 18 22 26 30 34 37 38 40
+ 41 43 44 46 47 48 67 68
r97 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r98 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r99 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r100 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r101 61 62 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r102 59 62 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=4.83 $Y2=2.72
r103 58 61 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=4.83 $Y2=2.72
r104 58 59 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r105 56 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r106 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r107 53 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r108 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r109 50 71 3.90382 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=2.72
+ $X2=0.235 $Y2=2.72
r110 50 52 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.47 $Y=2.72
+ $X2=1.15 $Y2=2.72
r111 48 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r112 48 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r113 46 64 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.99 $Y=2.72
+ $X2=5.75 $Y2=2.72
r114 46 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.99 $Y=2.72
+ $X2=6.115 $Y2=2.72
r115 45 67 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=6.24 $Y=2.72
+ $X2=6.67 $Y2=2.72
r116 45 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.24 $Y=2.72
+ $X2=6.115 $Y2=2.72
r117 43 61 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.05 $Y=2.72
+ $X2=4.83 $Y2=2.72
r118 43 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.05 $Y=2.72
+ $X2=5.175 $Y2=2.72
r119 42 64 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.3 $Y=2.72
+ $X2=5.75 $Y2=2.72
r120 42 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.3 $Y=2.72
+ $X2=5.175 $Y2=2.72
r121 40 55 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.1 $Y=2.72 $X2=2.07
+ $Y2=2.72
r122 40 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.1 $Y=2.72
+ $X2=2.225 $Y2=2.72
r123 39 58 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.35 $Y=2.72
+ $X2=2.53 $Y2=2.72
r124 39 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.35 $Y=2.72
+ $X2=2.225 $Y2=2.72
r125 37 52 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.16 $Y=2.72
+ $X2=1.15 $Y2=2.72
r126 37 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.16 $Y=2.72
+ $X2=1.285 $Y2=2.72
r127 36 55 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=2.07 $Y2=2.72
r128 36 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=1.285 $Y2=2.72
r129 32 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.115 $Y=2.635
+ $X2=6.115 $Y2=2.72
r130 32 34 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.115 $Y=2.635
+ $X2=6.115 $Y2=2.3
r131 28 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.175 $Y=2.635
+ $X2=5.175 $Y2=2.72
r132 28 30 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.175 $Y=2.635
+ $X2=5.175 $Y2=2.3
r133 24 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.635
+ $X2=2.225 $Y2=2.72
r134 24 26 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.225 $Y=2.635
+ $X2=2.225 $Y2=2.3
r135 20 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.635
+ $X2=1.285 $Y2=2.72
r136 20 22 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=1.285 $Y=2.635
+ $X2=1.285 $Y2=1.99
r137 16 71 3.23934 $w=2.5e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.345 $Y=2.635
+ $X2=0.235 $Y2=2.72
r138 16 18 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=0.345 $Y=2.635
+ $X2=0.345 $Y2=1.99
r139 5 34 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.97
+ $Y=1.485 $X2=6.115 $Y2=2.3
r140 4 30 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.03
+ $Y=1.485 $X2=5.175 $Y2=2.3
r141 3 26 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.08
+ $Y=1.485 $X2=2.225 $Y2=2.3
r142 2 22 300 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_PDIFF $count=2 $X=1.14
+ $Y=1.485 $X2=1.285 $Y2=1.99
r143 1 18 300 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_PDIFF $count=2 $X=0.2
+ $Y=1.485 $X2=0.345 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_4%X 1 2 3 4 13 14 15 16 19 23 27 29 33 37 43
+ 44 45
r73 42 45 10.3113 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=0.227 $Y=1.445
+ $X2=0.227 $Y2=1.19
r74 41 45 11.5244 $w=2.83e-07 $l=2.85e-07 $layer=LI1_cond $X=0.227 $Y=0.905
+ $X2=0.227 $Y2=1.19
r75 37 39 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=1.755 $Y=1.62
+ $X2=1.755 $Y2=2.3
r76 35 37 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.755 $Y=1.615
+ $X2=1.755 $Y2=1.62
r77 31 33 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.73 $Y=0.725
+ $X2=1.73 $Y2=0.39
r78 30 43 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=0.98 $Y=0.815
+ $X2=0.79 $Y2=0.815
r79 29 31 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=1.54 $Y=0.815
+ $X2=1.73 $Y2=0.725
r80 29 30 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.54 $Y=0.815
+ $X2=0.98 $Y2=0.815
r81 28 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.94 $Y=1.53
+ $X2=0.815 $Y2=1.53
r82 27 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.63 $Y=1.53
+ $X2=1.755 $Y2=1.615
r83 27 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.63 $Y=1.53 $X2=0.94
+ $Y2=1.53
r84 23 25 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.815 $Y=1.62
+ $X2=0.815 $Y2=2.3
r85 21 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=1.615
+ $X2=0.815 $Y2=1.53
r86 21 23 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.815 $Y=1.615
+ $X2=0.815 $Y2=1.62
r87 17 43 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=0.79 $Y=0.725 $X2=0.79
+ $Y2=0.815
r88 17 19 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.79 $Y=0.725
+ $X2=0.79 $Y2=0.39
r89 16 42 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=0.37 $Y=1.53
+ $X2=0.227 $Y2=1.445
r90 15 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.69 $Y=1.53
+ $X2=0.815 $Y2=1.53
r91 15 16 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.69 $Y=1.53 $X2=0.37
+ $Y2=1.53
r92 14 41 7.27854 $w=1.8e-07 $l=1.82535e-07 $layer=LI1_cond $X=0.37 $Y=0.815
+ $X2=0.227 $Y2=0.905
r93 13 43 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=0.6 $Y=0.815 $X2=0.79
+ $Y2=0.815
r94 13 14 14.1717 $w=1.78e-07 $l=2.3e-07 $layer=LI1_cond $X=0.6 $Y=0.815
+ $X2=0.37 $Y2=0.815
r95 4 39 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.61
+ $Y=1.485 $X2=1.755 $Y2=2.3
r96 4 37 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.61
+ $Y=1.485 $X2=1.755 $Y2=1.62
r97 3 25 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=1.485 $X2=0.815 $Y2=2.3
r98 3 23 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=1.485 $X2=0.815 $Y2=1.62
r99 2 33 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.57
+ $Y=0.235 $X2=1.755 $Y2=0.39
r100 1 19 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.63
+ $Y=0.235 $X2=0.815 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_4%A_524_297# 1 2 3 4 5 16 18 24 25 28 30 34
+ 38 41 46 50
c59 25 0 2.90511e-19 $X=4.83 $Y=1.87
r60 46 48 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.685 $Y=2.3 $X2=3.685
+ $Y2=2.38
r61 41 43 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.745 $Y=2.3 $X2=2.745
+ $Y2=2.38
r62 36 51 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.607 $Y=1.955
+ $X2=6.607 $Y2=1.87
r63 36 38 0.27051 $w=2.03e-07 $l=5e-09 $layer=LI1_cond $X=6.607 $Y=1.955
+ $X2=6.607 $Y2=1.96
r64 32 51 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.607 $Y=1.785
+ $X2=6.607 $Y2=1.87
r65 32 34 8.92683 $w=2.03e-07 $l=1.65e-07 $layer=LI1_cond $X=6.607 $Y=1.785
+ $X2=6.607 $Y2=1.62
r66 31 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.77 $Y=1.87
+ $X2=5.645 $Y2=1.87
r67 30 51 2.0246 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=6.505 $Y=1.87
+ $X2=6.607 $Y2=1.87
r68 30 31 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=6.505 $Y=1.87
+ $X2=5.77 $Y2=1.87
r69 26 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.645 $Y=1.955
+ $X2=5.645 $Y2=1.87
r70 26 28 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=5.645 $Y=1.955
+ $X2=5.645 $Y2=1.96
r71 24 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.52 $Y=1.87
+ $X2=5.645 $Y2=1.87
r72 24 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.52 $Y=1.87 $X2=4.83
+ $Y2=1.87
r73 21 23 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.665 $Y=2.295
+ $X2=4.665 $Y2=1.96
r74 20 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.665 $Y=1.955
+ $X2=4.83 $Y2=1.87
r75 20 23 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=4.665 $Y=1.955
+ $X2=4.665 $Y2=1.96
r76 19 48 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.81 $Y=2.38
+ $X2=3.685 $Y2=2.38
r77 18 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.5 $Y=2.38
+ $X2=4.665 $Y2=2.295
r78 18 19 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.5 $Y=2.38 $X2=3.81
+ $Y2=2.38
r79 17 43 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.87 $Y=2.38
+ $X2=2.745 $Y2=2.38
r80 16 48 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.56 $Y=2.38
+ $X2=3.685 $Y2=2.38
r81 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.56 $Y=2.38 $X2=2.87
+ $Y2=2.38
r82 5 38 300 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=2 $X=6.44
+ $Y=1.485 $X2=6.59 $Y2=1.96
r83 5 34 600 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=1 $X=6.44
+ $Y=1.485 $X2=6.59 $Y2=1.62
r84 4 28 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.5
+ $Y=1.485 $X2=5.645 $Y2=1.96
r85 3 23 300 $w=1.7e-07 $l=5.57786e-07 $layer=licon1_PDIFF $count=2 $X=4.48
+ $Y=1.485 $X2=4.66 $Y2=1.96
r86 2 46 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.54
+ $Y=1.485 $X2=3.685 $Y2=2.3
r87 1 41 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=2.62
+ $Y=1.485 $X2=2.745 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_4%VGND 1 2 3 4 5 18 22 26 28 30 33 34 36 37
+ 38 40 55 70 73 76
r96 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r97 72 73 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=0.235
+ $X2=2.83 $Y2=0.235
r98 68 72 4.01808 $w=6.38e-07 $l=2.15e-07 $layer=LI1_cond $X=2.53 $Y=0.235
+ $X2=2.745 $Y2=0.235
r99 68 70 14.6218 $w=6.38e-07 $l=3.9e-07 $layer=LI1_cond $X=2.53 $Y=0.235
+ $X2=2.14 $Y2=0.235
r100 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r101 63 66 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.345 $Y2=0
r102 61 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r103 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r104 58 61 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=6.21 $Y2=0
r105 57 60 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.83 $Y=0 $X2=6.21
+ $Y2=0
r106 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r107 55 75 3.40825 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=6.5 $Y=0 $X2=6.7 $Y2=0
r108 55 60 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.5 $Y=0 $X2=6.21
+ $Y2=0
r109 54 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r110 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r111 51 54 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=4.37 $Y2=0
r112 51 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r113 50 53 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.99 $Y=0 $X2=4.37
+ $Y2=0
r114 50 73 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=2.83
+ $Y2=0
r115 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r116 47 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r117 46 70 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.14
+ $Y2=0
r118 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r119 43 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r120 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r121 40 66 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.345
+ $Y2=0
r122 40 42 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=1.15
+ $Y2=0
r123 38 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r124 38 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r125 36 53 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.585 $Y=0
+ $X2=4.37 $Y2=0
r126 36 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.585 $Y=0 $X2=4.67
+ $Y2=0
r127 35 57 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.755 $Y=0 $X2=4.83
+ $Y2=0
r128 35 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.755 $Y=0 $X2=4.67
+ $Y2=0
r129 33 42 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.15
+ $Y2=0
r130 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.285
+ $Y2=0
r131 32 46 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.37 $Y=0 $X2=2.07
+ $Y2=0
r132 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=0 $X2=1.285
+ $Y2=0
r133 28 75 3.40825 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.585 $Y=0.085
+ $X2=6.7 $Y2=0
r134 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.585 $Y=0.085
+ $X2=6.585 $Y2=0.39
r135 24 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.67 $Y=0.085
+ $X2=4.67 $Y2=0
r136 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.67 $Y=0.085
+ $X2=4.67 $Y2=0.39
r137 20 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=0.085
+ $X2=1.285 $Y2=0
r138 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.285 $Y=0.085
+ $X2=1.285 $Y2=0.39
r139 16 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=0.085
+ $X2=0.345 $Y2=0
r140 16 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.345 $Y=0.085
+ $X2=0.345 $Y2=0.39
r141 5 30 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.45
+ $Y=0.235 $X2=6.585 $Y2=0.39
r142 4 26 182 $w=1.7e-07 $l=2.97574e-07 $layer=licon1_NDIFF $count=1 $X=4.44
+ $Y=0.235 $X2=4.67 $Y2=0.39
r143 3 72 91 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_NDIFF $count=2 $X=2.09
+ $Y=0.235 $X2=2.745 $Y2=0.39
r144 2 22 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.235 $X2=1.285 $Y2=0.39
r145 1 18 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=0.2
+ $Y=0.235 $X2=0.345 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_4%A_616_47# 1 2 11
r16 8 11 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=3.215 $Y=0.365
+ $X2=4.155 $Y2=0.365
r17 2 11 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.02
+ $Y=0.235 $X2=4.155 $Y2=0.39
r18 1 8 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.08
+ $Y=0.235 $X2=3.215 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_4%A_1008_47# 1 2 7 11 13
c21 13 0 1.70555e-19 $X=6.115 $Y=0.73
r22 11 16 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=6.155 $Y=0.475
+ $X2=6.155 $Y2=0.365
r23 11 13 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=6.155 $Y=0.475
+ $X2=6.155 $Y2=0.73
r24 7 16 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=6.03 $Y=0.365
+ $X2=6.155 $Y2=0.365
r25 7 9 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=6.03 $Y=0.365
+ $X2=5.175 $Y2=0.365
r26 2 16 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.98
+ $Y=0.235 $X2=6.115 $Y2=0.39
r27 2 13 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=5.98
+ $Y=0.235 $X2=6.115 $Y2=0.73
r28 1 9 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.235 $X2=5.175 $Y2=0.39
.ends

