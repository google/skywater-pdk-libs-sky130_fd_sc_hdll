* File: sky130_fd_sc_hdll__sdlclkp_2.pxi.spice
* Created: Wed Sep  2 08:52:51 2020
* 
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_2%SCE N_SCE_c_158_n N_SCE_c_159_n N_SCE_M1007_g
+ N_SCE_M1020_g SCE SCE N_SCE_c_157_n PM_SKY130_FD_SC_HDLL__SDLCLKP_2%SCE
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_2%GATE N_GATE_c_187_n N_GATE_c_188_n
+ N_GATE_M1002_g N_GATE_M1023_g GATE GATE N_GATE_c_185_n N_GATE_c_186_n
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_2%GATE
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_269_21# N_A_269_21#_M1016_d
+ N_A_269_21#_M1001_d N_A_269_21#_M1018_g N_A_269_21#_c_237_n
+ N_A_269_21#_M1009_g N_A_269_21#_c_226_n N_A_269_21#_M1022_g
+ N_A_269_21#_M1017_g N_A_269_21#_c_228_n N_A_269_21#_c_229_n
+ N_A_269_21#_c_230_n N_A_269_21#_c_231_n N_A_269_21#_c_232_n
+ N_A_269_21#_c_241_n N_A_269_21#_c_233_n N_A_269_21#_c_234_n
+ N_A_269_21#_c_235_n N_A_269_21#_c_236_n N_A_269_21#_c_243_n
+ N_A_269_21#_c_252_n N_A_269_21#_c_244_n N_A_269_21#_c_245_n
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_269_21#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_266_243# N_A_266_243#_M1017_s
+ N_A_266_243#_M1022_s N_A_266_243#_c_411_n N_A_266_243#_c_412_n
+ N_A_266_243#_M1021_g N_A_266_243#_c_399_n N_A_266_243#_c_400_n
+ N_A_266_243#_M1008_g N_A_266_243#_c_401_n N_A_266_243#_c_402_n
+ N_A_266_243#_c_403_n N_A_266_243#_c_416_n N_A_266_243#_c_404_n
+ N_A_266_243#_c_405_n N_A_266_243#_c_406_n N_A_266_243#_c_407_n
+ N_A_266_243#_c_408_n N_A_266_243#_c_409_n N_A_266_243#_c_410_n
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_266_243#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_484_315# N_A_484_315#_M1006_d
+ N_A_484_315#_M1000_d N_A_484_315#_c_528_n N_A_484_315#_M1010_g
+ N_A_484_315#_M1015_g N_A_484_315#_c_530_n N_A_484_315#_c_531_n
+ N_A_484_315#_M1019_g N_A_484_315#_M1004_g N_A_484_315#_c_532_n
+ N_A_484_315#_c_544_n N_A_484_315#_c_525_n N_A_484_315#_c_534_n
+ N_A_484_315#_c_526_n N_A_484_315#_c_555_n N_A_484_315#_c_556_n
+ N_A_484_315#_c_527_n PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_484_315#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_299_47# N_A_299_47#_M1018_d
+ N_A_299_47#_M1021_d N_A_299_47#_c_655_n N_A_299_47#_M1000_g
+ N_A_299_47#_c_656_n N_A_299_47#_M1006_g N_A_299_47#_c_669_n
+ N_A_299_47#_c_673_n N_A_299_47#_c_663_n N_A_299_47#_c_657_n
+ N_A_299_47#_c_658_n N_A_299_47#_c_659_n N_A_299_47#_c_660_n
+ N_A_299_47#_c_661_n PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_299_47#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_2%CLK N_CLK_c_757_n N_CLK_M1016_g N_CLK_c_758_n
+ N_CLK_M1001_g N_CLK_M1005_g N_CLK_c_768_n N_CLK_c_769_n N_CLK_M1013_g
+ N_CLK_c_760_n N_CLK_c_761_n N_CLK_c_762_n CLK N_CLK_c_763_n N_CLK_c_764_n
+ N_CLK_c_765_n CLK PM_SKY130_FD_SC_HDLL__SDLCLKP_2%CLK
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_1093_47# N_A_1093_47#_M1004_s
+ N_A_1093_47#_M1019_d N_A_1093_47#_M1012_g N_A_1093_47#_c_868_n
+ N_A_1093_47#_M1003_g N_A_1093_47#_M1014_g N_A_1093_47#_c_869_n
+ N_A_1093_47#_M1011_g N_A_1093_47#_c_874_n N_A_1093_47#_c_863_n
+ N_A_1093_47#_c_864_n N_A_1093_47#_c_882_n N_A_1093_47#_c_865_n
+ N_A_1093_47#_c_870_n N_A_1093_47#_c_871_n N_A_1093_47#_c_872_n
+ N_A_1093_47#_c_866_n N_A_1093_47#_c_867_n
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_1093_47#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_2%VPWR N_VPWR_M1007_s N_VPWR_M1010_d
+ N_VPWR_M1022_d N_VPWR_M1019_s N_VPWR_M1013_d N_VPWR_M1011_d N_VPWR_c_973_n
+ N_VPWR_c_974_n N_VPWR_c_975_n N_VPWR_c_976_n N_VPWR_c_977_n N_VPWR_c_978_n
+ N_VPWR_c_979_n N_VPWR_c_980_n N_VPWR_c_981_n VPWR N_VPWR_c_982_n
+ N_VPWR_c_983_n N_VPWR_c_984_n N_VPWR_c_985_n N_VPWR_c_986_n N_VPWR_c_972_n
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_2%VPWR
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_27_47# N_A_27_47#_M1020_s N_A_27_47#_M1023_d
+ N_A_27_47#_M1002_d N_A_27_47#_c_1078_n N_A_27_47#_c_1079_n N_A_27_47#_c_1080_n
+ N_A_27_47#_c_1081_n N_A_27_47#_c_1091_n N_A_27_47#_c_1100_n
+ N_A_27_47#_c_1104_n PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_2%GCLK N_GCLK_M1012_s N_GCLK_M1003_s
+ N_GCLK_c_1140_n N_GCLK_c_1134_n N_GCLK_c_1135_n N_GCLK_c_1137_n
+ N_GCLK_c_1138_n N_GCLK_c_1157_n GCLK GCLK GCLK
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_2%GCLK
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_2%VGND N_VGND_M1020_d N_VGND_M1015_d
+ N_VGND_M1017_d N_VGND_M1005_d N_VGND_M1014_d N_VGND_c_1180_n N_VGND_c_1181_n
+ N_VGND_c_1182_n N_VGND_c_1183_n N_VGND_c_1184_n N_VGND_c_1185_n VGND
+ N_VGND_c_1186_n N_VGND_c_1187_n N_VGND_c_1188_n N_VGND_c_1189_n
+ N_VGND_c_1190_n N_VGND_c_1191_n N_VGND_c_1192_n N_VGND_c_1193_n
+ N_VGND_c_1194_n PM_SKY130_FD_SC_HDLL__SDLCLKP_2%VGND
cc_1 VNB N_SCE_M1020_g 0.035163f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB SCE 0.0151026f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_SCE_c_157_n 0.0371984f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_4 VNB N_GATE_M1023_g 0.0277666f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_5 VNB N_GATE_c_185_n 0.0265431f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_6 VNB N_GATE_c_186_n 0.00500895f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_7 VNB N_A_269_21#_M1018_g 0.0199099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_269_21#_c_226_n 0.0264962f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_9 VNB N_A_269_21#_M1017_g 0.0397281f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_269_21#_c_228_n 0.00739628f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_269_21#_c_229_n 0.0299356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_269_21#_c_230_n 0.001574f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_269_21#_c_231_n 2.06267e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_269_21#_c_232_n 0.00455116f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_269_21#_c_233_n 0.00325423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_269_21#_c_234_n 0.00472736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_269_21#_c_235_n 0.0022361f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_269_21#_c_236_n 0.00121453f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_266_243#_c_399_n 0.0157472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_266_243#_c_400_n 0.00701612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_266_243#_c_401_n 0.012193f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_22 VNB N_A_266_243#_c_402_n 0.00834345f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.16
cc_23 VNB N_A_266_243#_c_403_n 0.00748877f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_24 VNB N_A_266_243#_c_404_n 0.0101381f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_266_243#_c_405_n 0.00127289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_266_243#_c_406_n 0.00298048f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_266_243#_c_407_n 0.00716656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_266_243#_c_408_n 0.0291478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_266_243#_c_409_n 0.00249917f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_266_243#_c_410_n 0.019636f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_484_315#_M1015_g 0.0454999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_484_315#_M1004_g 0.0324637f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.16
cc_33 VNB N_A_484_315#_c_525_n 0.00841237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_484_315#_c_526_n 0.00817014f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_484_315#_c_527_n 0.0309228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_299_47#_c_655_n 0.0279771f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_37 VNB N_A_299_47#_c_656_n 0.0210956f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_38 VNB N_A_299_47#_c_657_n 0.00231901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_299_47#_c_658_n 0.00217022f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_40 VNB N_A_299_47#_c_659_n 0.001861f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_299_47#_c_660_n 0.00258328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_299_47#_c_661_n 0.00219339f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_CLK_c_757_n 0.0179045f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_44 VNB N_CLK_c_758_n 0.0680418f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.165
cc_45 VNB N_CLK_M1005_g 0.0286167f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_46 VNB N_CLK_c_760_n 0.0123945f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_47 VNB N_CLK_c_761_n 0.00270586f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_48 VNB N_CLK_c_762_n 9.64156e-19 $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.16
cc_49 VNB N_CLK_c_763_n 0.00153979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_CLK_c_764_n 0.0239107f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_CLK_c_765_n 0.00309142f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_1093_47#_M1012_g 0.0188583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_1093_47#_M1014_g 0.0213796f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_54 VNB N_A_1093_47#_c_863_n 0.00300214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_1093_47#_c_864_n 0.00292893f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_1093_47#_c_865_n 0.00151223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1093_47#_c_866_n 0.00134722f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_1093_47#_c_867_n 0.0427537f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VPWR_c_972_n 0.326667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_27_47#_c_1078_n 0.0141581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_27_47#_c_1079_n 0.0040376f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_62 VNB N_A_27_47#_c_1080_n 0.00760745f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_63 VNB N_A_27_47#_c_1081_n 0.0109602f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_GCLK_c_1134_n 0.00852041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_GCLK_c_1135_n 0.00108392f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_66 VNB GCLK 0.0203888f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1180_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_68 VNB N_VGND_c_1181_n 0.00280416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1182_n 0.00559601f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1183_n 0.00476028f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1184_n 0.0466673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1185_n 0.0064059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1186_n 0.0142754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1187_n 0.048839f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1188_n 0.0325689f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1189_n 0.0184389f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1190_n 0.00556536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1191_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1192_n 0.00507043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1193_n 0.0132544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1194_n 0.39138f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VPB N_SCE_c_158_n 0.0182203f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.67
cc_83 VPB N_SCE_c_159_n 0.0288642f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_84 VPB SCE 0.0186881f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_85 VPB N_SCE_c_157_n 0.0111298f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_86 VPB N_GATE_c_187_n 0.017984f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.67
cc_87 VPB N_GATE_c_188_n 0.0218843f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_88 VPB N_GATE_c_185_n 0.00419169f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_89 VPB N_GATE_c_186_n 0.00549189f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_90 VPB N_A_269_21#_c_237_n 0.0517349f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_91 VPB N_A_269_21#_c_226_n 0.015049f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_92 VPB N_A_269_21#_M1022_g 0.04298f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_269_21#_c_231_n 0.00364558f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_269_21#_c_241_n 0.00528567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_269_21#_c_235_n 6.69987e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_269_21#_c_243_n 0.017135f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_269_21#_c_244_n 0.00417665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_269_21#_c_245_n 7.50236e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_266_243#_c_411_n 0.0310358f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_100 VPB N_A_266_243#_c_412_n 0.0240985f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_266_243#_c_399_n 0.0175257f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_266_243#_c_400_n 0.0024724f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_266_243#_c_403_n 0.00477958f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_104 VPB N_A_266_243#_c_416_n 0.00295943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_484_315#_c_528_n 0.0570583f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_106 VPB N_A_484_315#_M1015_g 0.0168089f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_484_315#_c_530_n 0.0235157f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_108 VPB N_A_484_315#_c_531_n 0.0266486f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_109 VPB N_A_484_315#_c_532_n 0.00246621f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_484_315#_c_525_n 0.00372102f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_484_315#_c_534_n 0.0183663f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_484_315#_c_526_n 0.00860187f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_484_315#_c_527_n 0.00807999f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_299_47#_c_655_n 0.0320723f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_115 VPB N_A_299_47#_c_663_n 0.0132653f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_299_47#_c_657_n 0.00162406f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_299_47#_c_658_n 8.46875e-19 $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_118 VPB N_A_299_47#_c_660_n 0.00331303f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_299_47#_c_661_n 5.36217e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_CLK_c_758_n 0.0174416f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.165
cc_121 VPB N_CLK_M1001_g 0.0444237f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_122 VPB N_CLK_c_768_n 0.0189233f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_CLK_c_769_n 0.0216549f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_124 VPB N_CLK_c_761_n 5.24179e-19 $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_125 VPB N_CLK_c_762_n 0.00130257f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.16
cc_126 VPB N_CLK_c_764_n 0.00426725f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_CLK_c_765_n 0.00160768f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_1093_47#_c_868_n 0.0163806f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_129 VPB N_A_1093_47#_c_869_n 0.0191065f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.16
cc_130 VPB N_A_1093_47#_c_870_n 0.00159926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_1093_47#_c_871_n 0.00384171f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_1093_47#_c_872_n 0.00549668f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_1093_47#_c_867_n 0.0131067f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_973_n 0.0098838f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_135 VPB N_VPWR_c_974_n 0.0319853f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.16
cc_136 VPB N_VPWR_c_975_n 0.00505078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_976_n 0.0111306f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_977_n 0.0305996f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_978_n 0.0318994f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_979_n 0.00468713f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_980_n 0.0165457f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_981_n 0.00631443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_982_n 0.0111737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_983_n 0.0200898f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_984_n 0.0540045f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_985_n 0.0135649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_986_n 0.0201646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_972_n 0.0484934f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_27_47#_c_1079_n 0.00315748f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_150 VPB N_GCLK_c_1137_n 0.00733629f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_151 VPB N_GCLK_c_1138_n 0.00107206f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB GCLK 0.00861602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 N_SCE_c_158_n N_GATE_c_187_n 0.0155764f $X=0.495 $Y=1.67 $X2=0 $Y2=0
cc_154 N_SCE_c_159_n N_GATE_c_188_n 0.063156f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_155 N_SCE_M1020_g N_GATE_M1023_g 0.0250971f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_156 N_SCE_c_157_n N_GATE_c_185_n 0.0155764f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_157 N_SCE_M1020_g N_GATE_c_186_n 7.03241e-19 $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_158 N_SCE_c_159_n N_VPWR_c_974_n 0.00695514f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_159 SCE N_VPWR_c_974_n 0.0228425f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_160 N_SCE_c_157_n N_VPWR_c_974_n 0.0013127f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_161 N_SCE_c_159_n N_VPWR_c_984_n 0.00596194f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_162 N_SCE_c_159_n N_VPWR_c_972_n 0.0107787f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_163 N_SCE_c_158_n N_A_27_47#_c_1079_n 0.00723144f $X=0.495 $Y=1.67 $X2=0
+ $Y2=0
cc_164 N_SCE_c_159_n N_A_27_47#_c_1079_n 0.0145271f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_165 N_SCE_M1020_g N_A_27_47#_c_1079_n 0.00997848f $X=0.52 $Y=0.445 $X2=0
+ $Y2=0
cc_166 SCE N_A_27_47#_c_1079_n 0.0483698f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_167 N_SCE_c_157_n N_A_27_47#_c_1079_n 0.0088623f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_168 N_SCE_M1020_g N_A_27_47#_c_1081_n 0.0136308f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_169 SCE N_A_27_47#_c_1081_n 0.020595f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_170 N_SCE_c_157_n N_A_27_47#_c_1081_n 0.00574324f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_171 N_SCE_c_159_n N_A_27_47#_c_1091_n 0.00888327f $X=0.495 $Y=1.77 $X2=0
+ $Y2=0
cc_172 N_SCE_M1020_g N_VGND_c_1186_n 0.00196986f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_173 N_SCE_M1020_g N_VGND_c_1190_n 0.0109522f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_174 N_SCE_M1020_g N_VGND_c_1194_n 0.00356708f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_175 N_GATE_M1023_g N_A_269_21#_M1018_g 0.0192791f $X=0.945 $Y=0.445 $X2=0
+ $Y2=0
cc_176 N_GATE_M1023_g N_A_269_21#_c_228_n 9.07621e-19 $X=0.945 $Y=0.445 $X2=0
+ $Y2=0
cc_177 N_GATE_c_185_n N_A_269_21#_c_228_n 0.00101819f $X=0.975 $Y=1.16 $X2=0
+ $Y2=0
cc_178 N_GATE_c_186_n N_A_269_21#_c_228_n 0.0814955f $X=0.975 $Y=1.16 $X2=0
+ $Y2=0
cc_179 N_GATE_c_185_n N_A_269_21#_c_229_n 5.37921e-19 $X=0.975 $Y=1.16 $X2=0
+ $Y2=0
cc_180 N_GATE_c_186_n N_A_269_21#_c_229_n 4.54129e-19 $X=0.975 $Y=1.16 $X2=0
+ $Y2=0
cc_181 N_GATE_c_186_n N_A_269_21#_c_252_n 0.0014166f $X=0.975 $Y=1.16 $X2=0
+ $Y2=0
cc_182 N_GATE_c_188_n N_A_269_21#_c_244_n 2.79092e-19 $X=0.905 $Y=1.77 $X2=0
+ $Y2=0
cc_183 N_GATE_c_188_n N_A_266_243#_c_411_n 0.0147124f $X=0.905 $Y=1.77 $X2=0
+ $Y2=0
cc_184 N_GATE_c_188_n N_A_266_243#_c_412_n 0.0162039f $X=0.905 $Y=1.77 $X2=0
+ $Y2=0
cc_185 N_GATE_c_187_n N_A_266_243#_c_400_n 0.00743476f $X=0.905 $Y=1.67 $X2=0
+ $Y2=0
cc_186 N_GATE_c_185_n N_A_266_243#_c_400_n 0.00676527f $X=0.975 $Y=1.16 $X2=0
+ $Y2=0
cc_187 N_GATE_c_186_n N_A_266_243#_c_400_n 0.00662406f $X=0.975 $Y=1.16 $X2=0
+ $Y2=0
cc_188 N_GATE_c_188_n N_VPWR_c_984_n 0.00429453f $X=0.905 $Y=1.77 $X2=0 $Y2=0
cc_189 N_GATE_c_188_n N_VPWR_c_972_n 0.00613085f $X=0.905 $Y=1.77 $X2=0 $Y2=0
cc_190 N_GATE_c_186_n N_VPWR_c_972_n 0.00134766f $X=0.975 $Y=1.16 $X2=0 $Y2=0
cc_191 N_GATE_c_186_n N_A_27_47#_M1002_d 0.00263629f $X=0.975 $Y=1.16 $X2=0
+ $Y2=0
cc_192 N_GATE_c_188_n N_A_27_47#_c_1079_n 0.00501283f $X=0.905 $Y=1.77 $X2=0
+ $Y2=0
cc_193 N_GATE_M1023_g N_A_27_47#_c_1079_n 0.00395487f $X=0.945 $Y=0.445 $X2=0
+ $Y2=0
cc_194 N_GATE_c_185_n N_A_27_47#_c_1079_n 0.00474152f $X=0.975 $Y=1.16 $X2=0
+ $Y2=0
cc_195 N_GATE_c_186_n N_A_27_47#_c_1079_n 0.0771243f $X=0.975 $Y=1.16 $X2=0
+ $Y2=0
cc_196 N_GATE_M1023_g N_A_27_47#_c_1080_n 0.0119096f $X=0.945 $Y=0.445 $X2=0
+ $Y2=0
cc_197 N_GATE_c_185_n N_A_27_47#_c_1080_n 0.00315152f $X=0.975 $Y=1.16 $X2=0
+ $Y2=0
cc_198 N_GATE_c_186_n N_A_27_47#_c_1080_n 0.0342766f $X=0.975 $Y=1.16 $X2=0
+ $Y2=0
cc_199 N_GATE_c_188_n N_A_27_47#_c_1100_n 0.0196183f $X=0.905 $Y=1.77 $X2=0
+ $Y2=0
cc_200 N_GATE_c_186_n N_A_27_47#_c_1100_n 0.0268868f $X=0.975 $Y=1.16 $X2=0
+ $Y2=0
cc_201 N_GATE_M1023_g N_VGND_c_1187_n 0.0035176f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_202 N_GATE_M1023_g N_VGND_c_1190_n 0.00759201f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_203 N_GATE_M1023_g N_VGND_c_1194_n 0.00420343f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_204 N_A_269_21#_c_237_n N_A_266_243#_c_411_n 0.0213218f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_205 N_A_269_21#_c_235_n N_A_266_243#_c_411_n 0.0031061f $X=1.712 $Y=1.452
+ $X2=0 $Y2=0
cc_206 N_A_269_21#_c_244_n N_A_266_243#_c_411_n 0.0117221f $X=1.71 $Y=1.53 $X2=0
+ $Y2=0
cc_207 N_A_269_21#_c_237_n N_A_266_243#_c_412_n 0.0123925f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_208 N_A_269_21#_c_244_n N_A_266_243#_c_412_n 0.00333464f $X=1.71 $Y=1.53
+ $X2=0 $Y2=0
cc_209 N_A_269_21#_c_237_n N_A_266_243#_c_399_n 0.021863f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_210 N_A_269_21#_c_235_n N_A_266_243#_c_399_n 0.019479f $X=1.712 $Y=1.452
+ $X2=0 $Y2=0
cc_211 N_A_269_21#_c_243_n N_A_266_243#_c_399_n 0.00280811f $X=4.44 $Y=1.53
+ $X2=0 $Y2=0
cc_212 N_A_269_21#_c_229_n N_A_266_243#_c_400_n 0.0262024f $X=1.55 $Y=0.87 $X2=0
+ $Y2=0
cc_213 N_A_269_21#_c_235_n N_A_266_243#_c_400_n 0.0027111f $X=1.712 $Y=1.452
+ $X2=0 $Y2=0
cc_214 N_A_269_21#_c_235_n N_A_266_243#_c_401_n 0.00135637f $X=1.712 $Y=1.452
+ $X2=0 $Y2=0
cc_215 N_A_269_21#_M1017_g N_A_266_243#_c_402_n 0.00734457f $X=4.24 $Y=0.445
+ $X2=0 $Y2=0
cc_216 N_A_269_21#_c_233_n N_A_266_243#_c_402_n 0.00782756f $X=4.96 $Y=0.615
+ $X2=0 $Y2=0
cc_217 N_A_269_21#_c_226_n N_A_266_243#_c_403_n 0.00643314f $X=4.215 $Y=1.44
+ $X2=0 $Y2=0
cc_218 N_A_269_21#_M1022_g N_A_266_243#_c_403_n 0.00152654f $X=4.215 $Y=1.835
+ $X2=0 $Y2=0
cc_219 N_A_269_21#_M1017_g N_A_266_243#_c_403_n 0.00225643f $X=4.24 $Y=0.445
+ $X2=0 $Y2=0
cc_220 N_A_269_21#_c_230_n N_A_266_243#_c_403_n 0.0132835f $X=4.365 $Y=1.19
+ $X2=0 $Y2=0
cc_221 N_A_269_21#_c_231_n N_A_266_243#_c_403_n 0.00949266f $X=4.517 $Y=1.495
+ $X2=0 $Y2=0
cc_222 N_A_269_21#_c_232_n N_A_266_243#_c_403_n 0.00563849f $X=4.525 $Y=1.105
+ $X2=0 $Y2=0
cc_223 N_A_269_21#_c_243_n N_A_266_243#_c_403_n 0.0105724f $X=4.44 $Y=1.53 $X2=0
+ $Y2=0
cc_224 N_A_269_21#_c_245_n N_A_266_243#_c_403_n 2.64595e-19 $X=4.585 $Y=1.53
+ $X2=0 $Y2=0
cc_225 N_A_269_21#_c_226_n N_A_266_243#_c_416_n 9.91151e-19 $X=4.215 $Y=1.44
+ $X2=0 $Y2=0
cc_226 N_A_269_21#_M1022_g N_A_266_243#_c_416_n 0.00240904f $X=4.215 $Y=1.835
+ $X2=0 $Y2=0
cc_227 N_A_269_21#_c_230_n N_A_266_243#_c_416_n 0.00178751f $X=4.365 $Y=1.19
+ $X2=0 $Y2=0
cc_228 N_A_269_21#_c_231_n N_A_266_243#_c_416_n 0.0108783f $X=4.517 $Y=1.495
+ $X2=0 $Y2=0
cc_229 N_A_269_21#_c_243_n N_A_266_243#_c_416_n 0.00992705f $X=4.44 $Y=1.53
+ $X2=0 $Y2=0
cc_230 N_A_269_21#_c_245_n N_A_266_243#_c_416_n 2.76111e-19 $X=4.585 $Y=1.53
+ $X2=0 $Y2=0
cc_231 N_A_269_21#_c_243_n N_A_266_243#_c_404_n 0.0697308f $X=4.44 $Y=1.53 $X2=0
+ $Y2=0
cc_232 N_A_269_21#_c_228_n N_A_266_243#_c_405_n 0.00137702f $X=1.55 $Y=0.87
+ $X2=0 $Y2=0
cc_233 N_A_269_21#_c_243_n N_A_266_243#_c_405_n 0.0131578f $X=4.44 $Y=1.53 $X2=0
+ $Y2=0
cc_234 N_A_269_21#_c_226_n N_A_266_243#_c_406_n 0.00181472f $X=4.215 $Y=1.44
+ $X2=0 $Y2=0
cc_235 N_A_269_21#_M1017_g N_A_266_243#_c_406_n 0.00655519f $X=4.24 $Y=0.445
+ $X2=0 $Y2=0
cc_236 N_A_269_21#_c_230_n N_A_266_243#_c_406_n 0.00258532f $X=4.365 $Y=1.19
+ $X2=0 $Y2=0
cc_237 N_A_269_21#_c_232_n N_A_266_243#_c_406_n 0.00545288f $X=4.525 $Y=1.105
+ $X2=0 $Y2=0
cc_238 N_A_269_21#_c_233_n N_A_266_243#_c_406_n 0.00140104f $X=4.96 $Y=0.615
+ $X2=0 $Y2=0
cc_239 N_A_269_21#_c_243_n N_A_266_243#_c_406_n 0.0151503f $X=4.44 $Y=1.53 $X2=0
+ $Y2=0
cc_240 N_A_269_21#_c_226_n N_A_266_243#_c_407_n 0.00207242f $X=4.215 $Y=1.44
+ $X2=0 $Y2=0
cc_241 N_A_269_21#_M1017_g N_A_266_243#_c_407_n 0.00372865f $X=4.24 $Y=0.445
+ $X2=0 $Y2=0
cc_242 N_A_269_21#_c_230_n N_A_266_243#_c_407_n 0.00527536f $X=4.365 $Y=1.19
+ $X2=0 $Y2=0
cc_243 N_A_269_21#_c_232_n N_A_266_243#_c_407_n 0.00790702f $X=4.525 $Y=1.105
+ $X2=0 $Y2=0
cc_244 N_A_269_21#_c_233_n N_A_266_243#_c_407_n 0.00107367f $X=4.96 $Y=0.615
+ $X2=0 $Y2=0
cc_245 N_A_269_21#_c_243_n N_A_266_243#_c_407_n 9.62924e-19 $X=4.44 $Y=1.53
+ $X2=0 $Y2=0
cc_246 N_A_269_21#_c_228_n N_A_266_243#_c_408_n 0.00737025f $X=1.55 $Y=0.87
+ $X2=0 $Y2=0
cc_247 N_A_269_21#_c_229_n N_A_266_243#_c_408_n 0.0167295f $X=1.55 $Y=0.87 $X2=0
+ $Y2=0
cc_248 N_A_269_21#_c_237_n N_A_266_243#_c_409_n 2.78293e-19 $X=1.96 $Y=1.99
+ $X2=0 $Y2=0
cc_249 N_A_269_21#_c_228_n N_A_266_243#_c_409_n 0.0247397f $X=1.55 $Y=0.87 $X2=0
+ $Y2=0
cc_250 N_A_269_21#_c_229_n N_A_266_243#_c_409_n 2.64542e-19 $X=1.55 $Y=0.87
+ $X2=0 $Y2=0
cc_251 N_A_269_21#_c_243_n N_A_266_243#_c_409_n 0.00522235f $X=4.44 $Y=1.53
+ $X2=0 $Y2=0
cc_252 N_A_269_21#_M1018_g N_A_266_243#_c_410_n 0.0132785f $X=1.42 $Y=0.415
+ $X2=0 $Y2=0
cc_253 N_A_269_21#_c_243_n N_A_484_315#_M1000_d 8.06277e-19 $X=4.44 $Y=1.53
+ $X2=0 $Y2=0
cc_254 N_A_269_21#_c_237_n N_A_484_315#_c_528_n 0.0289443f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_255 N_A_269_21#_c_243_n N_A_484_315#_c_528_n 0.00449033f $X=4.44 $Y=1.53
+ $X2=0 $Y2=0
cc_256 N_A_269_21#_c_243_n N_A_484_315#_M1015_g 0.00420735f $X=4.44 $Y=1.53
+ $X2=0 $Y2=0
cc_257 N_A_269_21#_c_241_n N_A_484_315#_c_530_n 0.00100947f $X=5.05 $Y=1.66
+ $X2=0 $Y2=0
cc_258 N_A_269_21#_c_233_n N_A_484_315#_M1004_g 4.8685e-19 $X=4.96 $Y=0.615
+ $X2=0 $Y2=0
cc_259 N_A_269_21#_c_243_n N_A_484_315#_c_532_n 0.0222174f $X=4.44 $Y=1.53 $X2=0
+ $Y2=0
cc_260 N_A_269_21#_M1022_g N_A_484_315#_c_544_n 0.00487772f $X=4.215 $Y=1.835
+ $X2=0 $Y2=0
cc_261 N_A_269_21#_c_243_n N_A_484_315#_c_525_n 0.022258f $X=4.44 $Y=1.53 $X2=0
+ $Y2=0
cc_262 N_A_269_21#_M1001_d N_A_484_315#_c_534_n 0.00503566f $X=4.905 $Y=1.515
+ $X2=0 $Y2=0
cc_263 N_A_269_21#_c_226_n N_A_484_315#_c_534_n 9.14009e-19 $X=4.215 $Y=1.44
+ $X2=0 $Y2=0
cc_264 N_A_269_21#_M1022_g N_A_484_315#_c_534_n 0.0164643f $X=4.215 $Y=1.835
+ $X2=0 $Y2=0
cc_265 N_A_269_21#_c_230_n N_A_484_315#_c_534_n 0.0016708f $X=4.365 $Y=1.19
+ $X2=0 $Y2=0
cc_266 N_A_269_21#_c_231_n N_A_484_315#_c_534_n 0.0230625f $X=4.517 $Y=1.495
+ $X2=0 $Y2=0
cc_267 N_A_269_21#_c_241_n N_A_484_315#_c_534_n 0.0311113f $X=5.05 $Y=1.66 $X2=0
+ $Y2=0
cc_268 N_A_269_21#_c_243_n N_A_484_315#_c_534_n 0.0151471f $X=4.44 $Y=1.53 $X2=0
+ $Y2=0
cc_269 N_A_269_21#_c_245_n N_A_484_315#_c_534_n 0.00170291f $X=4.585 $Y=1.53
+ $X2=0 $Y2=0
cc_270 N_A_269_21#_c_241_n N_A_484_315#_c_526_n 0.0203634f $X=5.05 $Y=1.66 $X2=0
+ $Y2=0
cc_271 N_A_269_21#_c_243_n N_A_484_315#_c_555_n 0.007409f $X=4.44 $Y=1.53 $X2=0
+ $Y2=0
cc_272 N_A_269_21#_M1022_g N_A_484_315#_c_556_n 0.00335363f $X=4.215 $Y=1.835
+ $X2=0 $Y2=0
cc_273 N_A_269_21#_c_243_n N_A_484_315#_c_556_n 0.00302634f $X=4.44 $Y=1.53
+ $X2=0 $Y2=0
cc_274 N_A_269_21#_c_243_n N_A_299_47#_c_655_n 0.0085668f $X=4.44 $Y=1.53 $X2=0
+ $Y2=0
cc_275 N_A_269_21#_M1018_g N_A_299_47#_c_669_n 0.00807723f $X=1.42 $Y=0.415
+ $X2=0 $Y2=0
cc_276 N_A_269_21#_c_228_n N_A_299_47#_c_669_n 0.0249565f $X=1.55 $Y=0.87 $X2=0
+ $Y2=0
cc_277 N_A_269_21#_c_229_n N_A_299_47#_c_669_n 0.00135285f $X=1.55 $Y=0.87 $X2=0
+ $Y2=0
cc_278 N_A_269_21#_c_235_n N_A_299_47#_c_669_n 0.00401633f $X=1.712 $Y=1.452
+ $X2=0 $Y2=0
cc_279 N_A_269_21#_c_237_n N_A_299_47#_c_673_n 0.0152026f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_280 N_A_269_21#_c_243_n N_A_299_47#_c_673_n 0.00562701f $X=4.44 $Y=1.53 $X2=0
+ $Y2=0
cc_281 N_A_269_21#_c_252_n N_A_299_47#_c_673_n 0.00102774f $X=1.855 $Y=1.53
+ $X2=0 $Y2=0
cc_282 N_A_269_21#_c_244_n N_A_299_47#_c_673_n 0.0255421f $X=1.71 $Y=1.53 $X2=0
+ $Y2=0
cc_283 N_A_269_21#_c_237_n N_A_299_47#_c_663_n 0.0073981f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_284 N_A_269_21#_c_235_n N_A_299_47#_c_663_n 0.0438627f $X=1.712 $Y=1.452
+ $X2=0 $Y2=0
cc_285 N_A_269_21#_c_243_n N_A_299_47#_c_663_n 0.0204925f $X=4.44 $Y=1.53 $X2=0
+ $Y2=0
cc_286 N_A_269_21#_c_252_n N_A_299_47#_c_663_n 5.16817e-19 $X=1.855 $Y=1.53
+ $X2=0 $Y2=0
cc_287 N_A_269_21#_c_243_n N_A_299_47#_c_657_n 0.005814f $X=4.44 $Y=1.53 $X2=0
+ $Y2=0
cc_288 N_A_269_21#_c_235_n N_A_299_47#_c_658_n 0.0147478f $X=1.712 $Y=1.452
+ $X2=0 $Y2=0
cc_289 N_A_269_21#_c_243_n N_A_299_47#_c_660_n 0.00800313f $X=4.44 $Y=1.53 $X2=0
+ $Y2=0
cc_290 N_A_269_21#_c_228_n N_A_299_47#_c_661_n 0.00566979f $X=1.55 $Y=0.87 $X2=0
+ $Y2=0
cc_291 N_A_269_21#_c_243_n N_A_299_47#_c_661_n 0.00229606f $X=4.44 $Y=1.53 $X2=0
+ $Y2=0
cc_292 N_A_269_21#_M1017_g N_CLK_c_757_n 0.0163343f $X=4.24 $Y=0.445 $X2=-0.19
+ $Y2=-0.24
cc_293 N_A_269_21#_c_233_n N_CLK_c_757_n 0.00757408f $X=4.96 $Y=0.615 $X2=-0.19
+ $Y2=-0.24
cc_294 N_A_269_21#_c_226_n N_CLK_c_758_n 0.015573f $X=4.215 $Y=1.44 $X2=0 $Y2=0
cc_295 N_A_269_21#_M1017_g N_CLK_c_758_n 0.00391642f $X=4.24 $Y=0.445 $X2=0
+ $Y2=0
cc_296 N_A_269_21#_c_231_n N_CLK_c_758_n 0.00373288f $X=4.517 $Y=1.495 $X2=0
+ $Y2=0
cc_297 N_A_269_21#_c_232_n N_CLK_c_758_n 0.011247f $X=4.525 $Y=1.105 $X2=0 $Y2=0
cc_298 N_A_269_21#_c_241_n N_CLK_c_758_n 0.00955851f $X=5.05 $Y=1.66 $X2=0 $Y2=0
cc_299 N_A_269_21#_c_233_n N_CLK_c_758_n 0.0227137f $X=4.96 $Y=0.615 $X2=0 $Y2=0
cc_300 N_A_269_21#_c_234_n N_CLK_c_758_n 0.0014877f $X=4.92 $Y=0.465 $X2=0 $Y2=0
cc_301 N_A_269_21#_c_236_n N_CLK_c_758_n 0.00193947f $X=4.517 $Y=1.19 $X2=0
+ $Y2=0
cc_302 N_A_269_21#_c_245_n N_CLK_c_758_n 0.00292718f $X=4.585 $Y=1.53 $X2=0
+ $Y2=0
cc_303 N_A_269_21#_M1022_g N_CLK_M1001_g 0.0345002f $X=4.215 $Y=1.835 $X2=0
+ $Y2=0
cc_304 N_A_269_21#_c_231_n N_CLK_M1001_g 0.00125292f $X=4.517 $Y=1.495 $X2=0
+ $Y2=0
cc_305 N_A_269_21#_c_241_n N_CLK_M1001_g 0.018759f $X=5.05 $Y=1.66 $X2=0 $Y2=0
cc_306 N_A_269_21#_c_245_n N_CLK_M1001_g 0.00256658f $X=4.585 $Y=1.53 $X2=0
+ $Y2=0
cc_307 N_A_269_21#_c_231_n N_CLK_c_761_n 7.04183e-19 $X=4.517 $Y=1.495 $X2=0
+ $Y2=0
cc_308 N_A_269_21#_c_232_n N_CLK_c_761_n 7.02927e-19 $X=4.525 $Y=1.105 $X2=0
+ $Y2=0
cc_309 N_A_269_21#_c_241_n N_CLK_c_761_n 0.00376482f $X=5.05 $Y=1.66 $X2=0 $Y2=0
cc_310 N_A_269_21#_c_233_n N_CLK_c_761_n 0.00120125f $X=4.96 $Y=0.615 $X2=0
+ $Y2=0
cc_311 N_A_269_21#_c_236_n N_CLK_c_761_n 0.00467158f $X=4.517 $Y=1.19 $X2=0
+ $Y2=0
cc_312 N_A_269_21#_c_226_n N_CLK_c_763_n 2.87927e-19 $X=4.215 $Y=1.44 $X2=0
+ $Y2=0
cc_313 N_A_269_21#_c_231_n N_CLK_c_763_n 0.00203498f $X=4.517 $Y=1.495 $X2=0
+ $Y2=0
cc_314 N_A_269_21#_c_232_n N_CLK_c_763_n 0.0050649f $X=4.525 $Y=1.105 $X2=0
+ $Y2=0
cc_315 N_A_269_21#_c_241_n N_CLK_c_763_n 0.015439f $X=5.05 $Y=1.66 $X2=0 $Y2=0
cc_316 N_A_269_21#_c_233_n N_CLK_c_763_n 0.00653509f $X=4.96 $Y=0.615 $X2=0
+ $Y2=0
cc_317 N_A_269_21#_c_236_n N_CLK_c_763_n 0.00653299f $X=4.517 $Y=1.19 $X2=0
+ $Y2=0
cc_318 N_A_269_21#_c_234_n N_A_1093_47#_c_874_n 0.01439f $X=4.92 $Y=0.465 $X2=0
+ $Y2=0
cc_319 N_A_269_21#_c_233_n N_A_1093_47#_c_864_n 0.00807626f $X=4.96 $Y=0.615
+ $X2=0 $Y2=0
cc_320 N_A_269_21#_c_243_n N_VPWR_M1010_d 0.00203938f $X=4.44 $Y=1.53 $X2=0
+ $Y2=0
cc_321 N_A_269_21#_c_231_n N_VPWR_M1022_d 0.00773199f $X=4.517 $Y=1.495 $X2=0
+ $Y2=0
cc_322 N_A_269_21#_c_243_n N_VPWR_M1022_d 5.63848e-19 $X=4.44 $Y=1.53 $X2=0
+ $Y2=0
cc_323 N_A_269_21#_M1022_g N_VPWR_c_978_n 0.0156985f $X=4.215 $Y=1.835 $X2=0
+ $Y2=0
cc_324 N_A_269_21#_M1022_g N_VPWR_c_982_n 0.00974554f $X=4.215 $Y=1.835 $X2=0
+ $Y2=0
cc_325 N_A_269_21#_c_237_n N_VPWR_c_984_n 0.00429453f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_326 N_A_269_21#_c_237_n N_VPWR_c_985_n 0.00138786f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_327 N_A_269_21#_c_243_n N_VPWR_c_985_n 6.32368e-19 $X=4.44 $Y=1.53 $X2=0
+ $Y2=0
cc_328 N_A_269_21#_c_237_n N_VPWR_c_972_n 0.00645844f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_329 N_A_269_21#_c_244_n N_VPWR_c_972_n 0.00621311f $X=1.71 $Y=1.53 $X2=0
+ $Y2=0
cc_330 N_A_269_21#_M1018_g N_A_27_47#_c_1080_n 0.0036696f $X=1.42 $Y=0.415 $X2=0
+ $Y2=0
cc_331 N_A_269_21#_c_228_n N_A_27_47#_c_1080_n 0.00671481f $X=1.55 $Y=0.87 $X2=0
+ $Y2=0
cc_332 N_A_269_21#_M1018_g N_A_27_47#_c_1104_n 4.57344e-19 $X=1.42 $Y=0.415
+ $X2=0 $Y2=0
cc_333 N_A_269_21#_c_233_n N_VGND_M1017_d 0.0025681f $X=4.96 $Y=0.615 $X2=0
+ $Y2=0
cc_334 N_A_269_21#_c_226_n N_VGND_c_1181_n 8.44957e-19 $X=4.215 $Y=1.44 $X2=0
+ $Y2=0
cc_335 N_A_269_21#_M1017_g N_VGND_c_1181_n 0.00878261f $X=4.24 $Y=0.445 $X2=0
+ $Y2=0
cc_336 N_A_269_21#_c_230_n N_VGND_c_1181_n 0.00121818f $X=4.365 $Y=1.19 $X2=0
+ $Y2=0
cc_337 N_A_269_21#_c_233_n N_VGND_c_1181_n 0.01501f $X=4.96 $Y=0.615 $X2=0 $Y2=0
cc_338 N_A_269_21#_c_236_n N_VGND_c_1181_n 3.25845e-19 $X=4.517 $Y=1.19 $X2=0
+ $Y2=0
cc_339 N_A_269_21#_c_233_n N_VGND_c_1184_n 0.00330694f $X=4.96 $Y=0.615 $X2=0
+ $Y2=0
cc_340 N_A_269_21#_c_234_n N_VGND_c_1184_n 0.0165187f $X=4.92 $Y=0.465 $X2=0
+ $Y2=0
cc_341 N_A_269_21#_M1018_g N_VGND_c_1187_n 0.00539883f $X=1.42 $Y=0.415 $X2=0
+ $Y2=0
cc_342 N_A_269_21#_M1017_g N_VGND_c_1188_n 0.0046653f $X=4.24 $Y=0.445 $X2=0
+ $Y2=0
cc_343 N_A_269_21#_M1018_g N_VGND_c_1190_n 0.00108095f $X=1.42 $Y=0.415 $X2=0
+ $Y2=0
cc_344 N_A_269_21#_M1016_d N_VGND_c_1194_n 0.00227267f $X=4.785 $Y=0.235 $X2=0
+ $Y2=0
cc_345 N_A_269_21#_M1018_g N_VGND_c_1194_n 0.0101587f $X=1.42 $Y=0.415 $X2=0
+ $Y2=0
cc_346 N_A_269_21#_M1017_g N_VGND_c_1194_n 0.00769683f $X=4.24 $Y=0.445 $X2=0
+ $Y2=0
cc_347 N_A_269_21#_c_233_n N_VGND_c_1194_n 0.00666319f $X=4.96 $Y=0.615 $X2=0
+ $Y2=0
cc_348 N_A_269_21#_c_234_n N_VGND_c_1194_n 0.00940011f $X=4.92 $Y=0.465 $X2=0
+ $Y2=0
cc_349 N_A_266_243#_c_404_n N_A_484_315#_M1006_d 0.00127746f $X=3.93 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_350 N_A_266_243#_c_401_n N_A_484_315#_M1015_g 0.00699103f $X=2.022 $Y=1.215
+ $X2=0 $Y2=0
cc_351 N_A_266_243#_c_404_n N_A_484_315#_M1015_g 0.00341307f $X=3.93 $Y=0.85
+ $X2=0 $Y2=0
cc_352 N_A_266_243#_c_408_n N_A_484_315#_M1015_g 0.0115719f $X=2.06 $Y=0.87
+ $X2=0 $Y2=0
cc_353 N_A_266_243#_c_409_n N_A_484_315#_M1015_g 7.93707e-19 $X=2.06 $Y=0.87
+ $X2=0 $Y2=0
cc_354 N_A_266_243#_c_410_n N_A_484_315#_M1015_g 0.0121621f $X=2.082 $Y=0.705
+ $X2=0 $Y2=0
cc_355 N_A_266_243#_c_402_n N_A_484_315#_c_525_n 0.0910502f $X=3.98 $Y=0.465
+ $X2=0 $Y2=0
cc_356 N_A_266_243#_c_416_n N_A_484_315#_c_525_n 0.00406408f $X=3.98 $Y=1.66
+ $X2=0 $Y2=0
cc_357 N_A_266_243#_c_404_n N_A_484_315#_c_525_n 0.0175797f $X=3.93 $Y=0.85
+ $X2=0 $Y2=0
cc_358 N_A_266_243#_c_406_n N_A_484_315#_c_525_n 2.87915e-19 $X=4.075 $Y=0.85
+ $X2=0 $Y2=0
cc_359 N_A_266_243#_M1022_s N_A_484_315#_c_534_n 0.00535544f $X=3.855 $Y=1.515
+ $X2=0 $Y2=0
cc_360 N_A_266_243#_c_416_n N_A_484_315#_c_534_n 0.024093f $X=3.98 $Y=1.66 $X2=0
+ $Y2=0
cc_361 N_A_266_243#_c_416_n N_A_484_315#_c_556_n 0.00889198f $X=3.98 $Y=1.66
+ $X2=0 $Y2=0
cc_362 N_A_266_243#_c_416_n N_A_299_47#_c_655_n 5.9685e-19 $X=3.98 $Y=1.66 $X2=0
+ $Y2=0
cc_363 N_A_266_243#_c_404_n N_A_299_47#_c_655_n 0.00370099f $X=3.93 $Y=0.85
+ $X2=0 $Y2=0
cc_364 N_A_266_243#_c_404_n N_A_299_47#_c_656_n 0.0088114f $X=3.93 $Y=0.85 $X2=0
+ $Y2=0
cc_365 N_A_266_243#_c_400_n N_A_299_47#_c_669_n 7.38226e-19 $X=1.53 $Y=1.29
+ $X2=0 $Y2=0
cc_366 N_A_266_243#_c_404_n N_A_299_47#_c_669_n 0.00173979f $X=3.93 $Y=0.85
+ $X2=0 $Y2=0
cc_367 N_A_266_243#_c_405_n N_A_299_47#_c_669_n 0.00205588f $X=2.365 $Y=0.85
+ $X2=0 $Y2=0
cc_368 N_A_266_243#_c_408_n N_A_299_47#_c_669_n 0.00375911f $X=2.06 $Y=0.87
+ $X2=0 $Y2=0
cc_369 N_A_266_243#_c_409_n N_A_299_47#_c_669_n 0.0212161f $X=2.06 $Y=0.87 $X2=0
+ $Y2=0
cc_370 N_A_266_243#_c_410_n N_A_299_47#_c_669_n 0.0130546f $X=2.082 $Y=0.705
+ $X2=0 $Y2=0
cc_371 N_A_266_243#_c_411_n N_A_299_47#_c_663_n 6.38369e-19 $X=1.43 $Y=1.89
+ $X2=0 $Y2=0
cc_372 N_A_266_243#_c_404_n N_A_299_47#_c_657_n 0.00153861f $X=3.93 $Y=0.85
+ $X2=0 $Y2=0
cc_373 N_A_266_243#_c_405_n N_A_299_47#_c_657_n 9.40357e-19 $X=2.365 $Y=0.85
+ $X2=0 $Y2=0
cc_374 N_A_266_243#_c_409_n N_A_299_47#_c_657_n 3.1525e-19 $X=2.06 $Y=0.87 $X2=0
+ $Y2=0
cc_375 N_A_266_243#_c_401_n N_A_299_47#_c_658_n 0.00225667f $X=2.022 $Y=1.215
+ $X2=0 $Y2=0
cc_376 N_A_266_243#_c_405_n N_A_299_47#_c_658_n 7.66293e-19 $X=2.365 $Y=0.85
+ $X2=0 $Y2=0
cc_377 N_A_266_243#_c_408_n N_A_299_47#_c_658_n 0.00256252f $X=2.06 $Y=0.87
+ $X2=0 $Y2=0
cc_378 N_A_266_243#_c_409_n N_A_299_47#_c_658_n 0.0127085f $X=2.06 $Y=0.87 $X2=0
+ $Y2=0
cc_379 N_A_266_243#_c_404_n N_A_299_47#_c_659_n 0.0164716f $X=3.93 $Y=0.85 $X2=0
+ $Y2=0
cc_380 N_A_266_243#_c_405_n N_A_299_47#_c_659_n 0.00275249f $X=2.365 $Y=0.85
+ $X2=0 $Y2=0
cc_381 N_A_266_243#_c_408_n N_A_299_47#_c_659_n 7.43573e-19 $X=2.06 $Y=0.87
+ $X2=0 $Y2=0
cc_382 N_A_266_243#_c_409_n N_A_299_47#_c_659_n 0.0206686f $X=2.06 $Y=0.87 $X2=0
+ $Y2=0
cc_383 N_A_266_243#_c_410_n N_A_299_47#_c_659_n 0.00291704f $X=2.082 $Y=0.705
+ $X2=0 $Y2=0
cc_384 N_A_266_243#_c_404_n N_A_299_47#_c_660_n 0.016448f $X=3.93 $Y=0.85 $X2=0
+ $Y2=0
cc_385 N_A_266_243#_c_401_n N_A_299_47#_c_661_n 0.00188395f $X=2.022 $Y=1.215
+ $X2=0 $Y2=0
cc_386 N_A_266_243#_c_409_n N_A_299_47#_c_661_n 0.00346892f $X=2.06 $Y=0.87
+ $X2=0 $Y2=0
cc_387 N_A_266_243#_c_412_n N_VPWR_c_984_n 0.00743866f $X=1.43 $Y=1.99 $X2=0
+ $Y2=0
cc_388 N_A_266_243#_c_412_n N_VPWR_c_972_n 0.0118046f $X=1.43 $Y=1.99 $X2=0
+ $Y2=0
cc_389 N_A_266_243#_c_404_n N_VGND_M1015_d 0.00222845f $X=3.93 $Y=0.85 $X2=0
+ $Y2=0
cc_390 N_A_266_243#_c_404_n N_VGND_c_1180_n 0.00775574f $X=3.93 $Y=0.85 $X2=0
+ $Y2=0
cc_391 N_A_266_243#_c_402_n N_VGND_c_1181_n 0.012098f $X=3.98 $Y=0.465 $X2=0
+ $Y2=0
cc_392 N_A_266_243#_c_410_n N_VGND_c_1187_n 0.00357877f $X=2.082 $Y=0.705 $X2=0
+ $Y2=0
cc_393 N_A_266_243#_c_402_n N_VGND_c_1188_n 0.0232287f $X=3.98 $Y=0.465 $X2=0
+ $Y2=0
cc_394 N_A_266_243#_M1017_s N_VGND_c_1194_n 0.00233457f $X=3.855 $Y=0.235 $X2=0
+ $Y2=0
cc_395 N_A_266_243#_c_402_n N_VGND_c_1194_n 0.00590194f $X=3.98 $Y=0.465 $X2=0
+ $Y2=0
cc_396 N_A_266_243#_c_404_n N_VGND_c_1194_n 0.075561f $X=3.93 $Y=0.85 $X2=0
+ $Y2=0
cc_397 N_A_266_243#_c_405_n N_VGND_c_1194_n 0.0148704f $X=2.365 $Y=0.85 $X2=0
+ $Y2=0
cc_398 N_A_266_243#_c_406_n N_VGND_c_1194_n 0.0154936f $X=4.075 $Y=0.85 $X2=0
+ $Y2=0
cc_399 N_A_266_243#_c_407_n N_VGND_c_1194_n 6.80412e-19 $X=4.075 $Y=0.85 $X2=0
+ $Y2=0
cc_400 N_A_266_243#_c_410_n N_VGND_c_1194_n 0.00611524f $X=2.082 $Y=0.705 $X2=0
+ $Y2=0
cc_401 N_A_484_315#_c_528_n N_A_299_47#_c_655_n 0.0141627f $X=2.52 $Y=1.99 $X2=0
+ $Y2=0
cc_402 N_A_484_315#_M1015_g N_A_299_47#_c_655_n 0.033994f $X=2.655 $Y=0.445
+ $X2=0 $Y2=0
cc_403 N_A_484_315#_c_532_n N_A_299_47#_c_655_n 0.0217841f $X=3.325 $Y=1.77
+ $X2=0 $Y2=0
cc_404 N_A_484_315#_c_525_n N_A_299_47#_c_655_n 0.0079676f $X=3.46 $Y=0.42 $X2=0
+ $Y2=0
cc_405 N_A_484_315#_c_555_n N_A_299_47#_c_655_n 3.54096e-19 $X=2.665 $Y=1.74
+ $X2=0 $Y2=0
cc_406 N_A_484_315#_M1015_g N_A_299_47#_c_656_n 0.0160518f $X=2.655 $Y=0.445
+ $X2=0 $Y2=0
cc_407 N_A_484_315#_c_525_n N_A_299_47#_c_656_n 0.0207844f $X=3.46 $Y=0.42 $X2=0
+ $Y2=0
cc_408 N_A_484_315#_M1015_g N_A_299_47#_c_669_n 0.00982828f $X=2.655 $Y=0.445
+ $X2=0 $Y2=0
cc_409 N_A_484_315#_c_528_n N_A_299_47#_c_673_n 0.00307829f $X=2.52 $Y=1.99
+ $X2=0 $Y2=0
cc_410 N_A_484_315#_c_528_n N_A_299_47#_c_663_n 0.00690356f $X=2.52 $Y=1.99
+ $X2=0 $Y2=0
cc_411 N_A_484_315#_M1015_g N_A_299_47#_c_663_n 0.00512785f $X=2.655 $Y=0.445
+ $X2=0 $Y2=0
cc_412 N_A_484_315#_c_555_n N_A_299_47#_c_663_n 0.0255996f $X=2.665 $Y=1.74
+ $X2=0 $Y2=0
cc_413 N_A_484_315#_c_528_n N_A_299_47#_c_657_n 0.00169011f $X=2.52 $Y=1.99
+ $X2=0 $Y2=0
cc_414 N_A_484_315#_c_555_n N_A_299_47#_c_657_n 2.34133e-19 $X=2.665 $Y=1.74
+ $X2=0 $Y2=0
cc_415 N_A_484_315#_M1015_g N_A_299_47#_c_659_n 0.0121803f $X=2.655 $Y=0.445
+ $X2=0 $Y2=0
cc_416 N_A_484_315#_M1015_g N_A_299_47#_c_660_n 0.00997152f $X=2.655 $Y=0.445
+ $X2=0 $Y2=0
cc_417 N_A_484_315#_c_532_n N_A_299_47#_c_660_n 0.0189559f $X=3.325 $Y=1.77
+ $X2=0 $Y2=0
cc_418 N_A_484_315#_c_525_n N_A_299_47#_c_660_n 0.0302043f $X=3.46 $Y=0.42 $X2=0
+ $Y2=0
cc_419 N_A_484_315#_c_555_n N_A_299_47#_c_660_n 0.00101123f $X=2.665 $Y=1.74
+ $X2=0 $Y2=0
cc_420 N_A_484_315#_c_528_n N_A_299_47#_c_661_n 0.00197841f $X=2.52 $Y=1.99
+ $X2=0 $Y2=0
cc_421 N_A_484_315#_M1015_g N_A_299_47#_c_661_n 0.00801241f $X=2.655 $Y=0.445
+ $X2=0 $Y2=0
cc_422 N_A_484_315#_c_555_n N_A_299_47#_c_661_n 0.00960172f $X=2.665 $Y=1.74
+ $X2=0 $Y2=0
cc_423 N_A_484_315#_M1004_g N_CLK_c_758_n 0.00672564f $X=5.85 $Y=0.445 $X2=0
+ $Y2=0
cc_424 N_A_484_315#_c_526_n N_CLK_c_758_n 0.00429576f $X=5.63 $Y=1.16 $X2=0
+ $Y2=0
cc_425 N_A_484_315#_c_527_n N_CLK_c_758_n 0.0131957f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_426 N_A_484_315#_c_534_n N_CLK_M1001_g 0.0144753f $X=5.405 $Y=2 $X2=0 $Y2=0
cc_427 N_A_484_315#_c_526_n N_CLK_M1001_g 0.0051364f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_428 N_A_484_315#_M1004_g N_CLK_M1005_g 0.0389322f $X=5.85 $Y=0.445 $X2=0
+ $Y2=0
cc_429 N_A_484_315#_c_530_n N_CLK_c_768_n 0.00982937f $X=5.825 $Y=1.67 $X2=0
+ $Y2=0
cc_430 N_A_484_315#_c_526_n N_CLK_c_768_n 9.85577e-19 $X=5.63 $Y=1.16 $X2=0
+ $Y2=0
cc_431 N_A_484_315#_c_531_n N_CLK_c_769_n 0.028118f $X=5.825 $Y=1.77 $X2=0 $Y2=0
cc_432 N_A_484_315#_c_526_n N_CLK_c_760_n 0.0351863f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_433 N_A_484_315#_c_527_n N_CLK_c_760_n 0.00965113f $X=5.85 $Y=1.16 $X2=0
+ $Y2=0
cc_434 N_A_484_315#_c_534_n N_CLK_c_761_n 8.29701e-19 $X=5.405 $Y=2 $X2=0 $Y2=0
cc_435 N_A_484_315#_c_526_n N_CLK_c_761_n 0.00271044f $X=5.63 $Y=1.16 $X2=0
+ $Y2=0
cc_436 N_A_484_315#_c_526_n N_CLK_c_762_n 0.00259415f $X=5.63 $Y=1.16 $X2=0
+ $Y2=0
cc_437 N_A_484_315#_c_527_n N_CLK_c_762_n 0.00155353f $X=5.85 $Y=1.16 $X2=0
+ $Y2=0
cc_438 N_A_484_315#_c_526_n N_CLK_c_763_n 0.0181472f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_439 N_A_484_315#_c_527_n N_CLK_c_763_n 4.90794e-19 $X=5.85 $Y=1.16 $X2=0
+ $Y2=0
cc_440 N_A_484_315#_c_526_n N_CLK_c_764_n 3.15598e-19 $X=5.63 $Y=1.16 $X2=0
+ $Y2=0
cc_441 N_A_484_315#_c_527_n N_CLK_c_764_n 0.0389322f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_442 N_A_484_315#_c_526_n N_CLK_c_765_n 0.0185868f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_443 N_A_484_315#_c_527_n N_CLK_c_765_n 0.00245047f $X=5.85 $Y=1.16 $X2=0
+ $Y2=0
cc_444 N_A_484_315#_M1004_g N_A_1093_47#_c_874_n 0.00486638f $X=5.85 $Y=0.445
+ $X2=0 $Y2=0
cc_445 N_A_484_315#_M1004_g N_A_1093_47#_c_863_n 0.0122663f $X=5.85 $Y=0.445
+ $X2=0 $Y2=0
cc_446 N_A_484_315#_c_526_n N_A_1093_47#_c_863_n 0.0048853f $X=5.63 $Y=1.16
+ $X2=0 $Y2=0
cc_447 N_A_484_315#_c_527_n N_A_1093_47#_c_863_n 0.00136242f $X=5.85 $Y=1.16
+ $X2=0 $Y2=0
cc_448 N_A_484_315#_c_526_n N_A_1093_47#_c_864_n 0.0114741f $X=5.63 $Y=1.16
+ $X2=0 $Y2=0
cc_449 N_A_484_315#_c_527_n N_A_1093_47#_c_864_n 0.00127183f $X=5.85 $Y=1.16
+ $X2=0 $Y2=0
cc_450 N_A_484_315#_c_531_n N_A_1093_47#_c_882_n 0.00471521f $X=5.825 $Y=1.77
+ $X2=0 $Y2=0
cc_451 N_A_484_315#_c_530_n N_A_1093_47#_c_872_n 0.00255489f $X=5.825 $Y=1.67
+ $X2=0 $Y2=0
cc_452 N_A_484_315#_c_531_n N_A_1093_47#_c_872_n 0.00222724f $X=5.825 $Y=1.77
+ $X2=0 $Y2=0
cc_453 N_A_484_315#_c_534_n N_A_1093_47#_c_872_n 0.0120899f $X=5.405 $Y=2 $X2=0
+ $Y2=0
cc_454 N_A_484_315#_c_526_n N_A_1093_47#_c_872_n 0.0290204f $X=5.63 $Y=1.16
+ $X2=0 $Y2=0
cc_455 N_A_484_315#_c_532_n N_VPWR_M1010_d 0.00492813f $X=3.325 $Y=1.77 $X2=0
+ $Y2=0
cc_456 N_A_484_315#_c_534_n N_VPWR_M1022_d 0.00659411f $X=5.405 $Y=2 $X2=0 $Y2=0
cc_457 N_A_484_315#_c_534_n N_VPWR_M1019_s 0.00350191f $X=5.405 $Y=2 $X2=0 $Y2=0
cc_458 N_A_484_315#_c_526_n N_VPWR_M1019_s 3.81917e-19 $X=5.63 $Y=1.16 $X2=0
+ $Y2=0
cc_459 N_A_484_315#_c_534_n N_VPWR_c_978_n 0.0243816f $X=5.405 $Y=2 $X2=0 $Y2=0
cc_460 N_A_484_315#_c_531_n N_VPWR_c_979_n 0.00851749f $X=5.825 $Y=1.77 $X2=0
+ $Y2=0
cc_461 N_A_484_315#_c_531_n N_VPWR_c_980_n 0.00622633f $X=5.825 $Y=1.77 $X2=0
+ $Y2=0
cc_462 N_A_484_315#_c_544_n N_VPWR_c_982_n 0.0107733f $X=3.46 $Y=2.205 $X2=0
+ $Y2=0
cc_463 N_A_484_315#_c_534_n N_VPWR_c_982_n 0.107308f $X=5.405 $Y=2 $X2=0 $Y2=0
cc_464 N_A_484_315#_c_528_n N_VPWR_c_984_n 0.00368409f $X=2.52 $Y=1.99 $X2=0
+ $Y2=0
cc_465 N_A_484_315#_c_528_n N_VPWR_c_985_n 0.0256563f $X=2.52 $Y=1.99 $X2=0
+ $Y2=0
cc_466 N_A_484_315#_c_555_n N_VPWR_c_985_n 0.0407968f $X=2.665 $Y=1.74 $X2=0
+ $Y2=0
cc_467 N_A_484_315#_c_544_n N_VPWR_c_986_n 0.0137273f $X=3.46 $Y=2.205 $X2=0
+ $Y2=0
cc_468 N_A_484_315#_c_534_n N_VPWR_c_986_n 0.0052614f $X=5.405 $Y=2 $X2=0 $Y2=0
cc_469 N_A_484_315#_M1000_d N_VPWR_c_972_n 0.00237624f $X=3.315 $Y=1.485 $X2=0
+ $Y2=0
cc_470 N_A_484_315#_c_528_n N_VPWR_c_972_n 0.00514038f $X=2.52 $Y=1.99 $X2=0
+ $Y2=0
cc_471 N_A_484_315#_c_531_n N_VPWR_c_972_n 0.0104567f $X=5.825 $Y=1.77 $X2=0
+ $Y2=0
cc_472 N_A_484_315#_c_532_n N_VPWR_c_972_n 0.00668636f $X=3.325 $Y=1.77 $X2=0
+ $Y2=0
cc_473 N_A_484_315#_c_544_n N_VPWR_c_972_n 0.00839556f $X=3.46 $Y=2.205 $X2=0
+ $Y2=0
cc_474 N_A_484_315#_c_534_n N_VPWR_c_972_n 0.0186575f $X=5.405 $Y=2 $X2=0 $Y2=0
cc_475 N_A_484_315#_c_555_n N_VPWR_c_972_n 0.00344844f $X=2.665 $Y=1.74 $X2=0
+ $Y2=0
cc_476 N_A_484_315#_M1015_g N_VGND_c_1180_n 0.00720923f $X=2.655 $Y=0.445 $X2=0
+ $Y2=0
cc_477 N_A_484_315#_c_525_n N_VGND_c_1180_n 0.0140386f $X=3.46 $Y=0.42 $X2=0
+ $Y2=0
cc_478 N_A_484_315#_M1004_g N_VGND_c_1184_n 0.00422112f $X=5.85 $Y=0.445 $X2=0
+ $Y2=0
cc_479 N_A_484_315#_M1015_g N_VGND_c_1187_n 0.00486707f $X=2.655 $Y=0.445 $X2=0
+ $Y2=0
cc_480 N_A_484_315#_c_525_n N_VGND_c_1188_n 0.0116048f $X=3.46 $Y=0.42 $X2=0
+ $Y2=0
cc_481 N_A_484_315#_M1006_d N_VGND_c_1194_n 0.00243215f $X=3.325 $Y=0.235 $X2=0
+ $Y2=0
cc_482 N_A_484_315#_M1015_g N_VGND_c_1194_n 0.0068389f $X=2.655 $Y=0.445 $X2=0
+ $Y2=0
cc_483 N_A_484_315#_M1004_g N_VGND_c_1194_n 0.00707149f $X=5.85 $Y=0.445 $X2=0
+ $Y2=0
cc_484 N_A_484_315#_c_525_n N_VGND_c_1194_n 0.00308197f $X=3.46 $Y=0.42 $X2=0
+ $Y2=0
cc_485 N_A_299_47#_c_655_n N_VPWR_c_982_n 0.00300894f $X=3.225 $Y=1.41 $X2=0
+ $Y2=0
cc_486 N_A_299_47#_c_673_n N_VPWR_c_984_n 0.0424693f $X=2.13 $Y=2.295 $X2=0
+ $Y2=0
cc_487 N_A_299_47#_c_655_n N_VPWR_c_985_n 0.0067571f $X=3.225 $Y=1.41 $X2=0
+ $Y2=0
cc_488 N_A_299_47#_c_673_n N_VPWR_c_985_n 0.0240862f $X=2.13 $Y=2.295 $X2=0
+ $Y2=0
cc_489 N_A_299_47#_c_663_n N_VPWR_c_985_n 0.00308511f $X=2.215 $Y=2.125 $X2=0
+ $Y2=0
cc_490 N_A_299_47#_c_655_n N_VPWR_c_986_n 0.0062441f $X=3.225 $Y=1.41 $X2=0
+ $Y2=0
cc_491 N_A_299_47#_M1021_d N_VPWR_c_972_n 0.00328896f $X=1.52 $Y=2.065 $X2=0
+ $Y2=0
cc_492 N_A_299_47#_c_655_n N_VPWR_c_972_n 0.00903378f $X=3.225 $Y=1.41 $X2=0
+ $Y2=0
cc_493 N_A_299_47#_c_673_n N_VPWR_c_972_n 0.0253092f $X=2.13 $Y=2.295 $X2=0
+ $Y2=0
cc_494 N_A_299_47#_c_673_n N_A_27_47#_c_1100_n 0.0186379f $X=2.13 $Y=2.295 $X2=0
+ $Y2=0
cc_495 N_A_299_47#_c_673_n A_410_413# 0.00683749f $X=2.13 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_496 N_A_299_47#_c_663_n A_410_413# 0.0014313f $X=2.215 $Y=2.125 $X2=-0.19
+ $Y2=-0.24
cc_497 N_A_299_47#_c_655_n N_VGND_c_1180_n 0.00209689f $X=3.225 $Y=1.41 $X2=0
+ $Y2=0
cc_498 N_A_299_47#_c_656_n N_VGND_c_1180_n 0.0064755f $X=3.25 $Y=0.995 $X2=0
+ $Y2=0
cc_499 N_A_299_47#_c_669_n N_VGND_c_1180_n 0.0156107f $X=2.475 $Y=0.395 $X2=0
+ $Y2=0
cc_500 N_A_299_47#_c_659_n N_VGND_c_1180_n 0.0138859f $X=2.56 $Y=0.995 $X2=0
+ $Y2=0
cc_501 N_A_299_47#_c_660_n N_VGND_c_1180_n 0.0112879f $X=3.12 $Y=1.16 $X2=0
+ $Y2=0
cc_502 N_A_299_47#_c_669_n N_VGND_c_1187_n 0.0704643f $X=2.475 $Y=0.395 $X2=0
+ $Y2=0
cc_503 N_A_299_47#_c_656_n N_VGND_c_1188_n 0.00585385f $X=3.25 $Y=0.995 $X2=0
+ $Y2=0
cc_504 N_A_299_47#_M1018_d N_VGND_c_1194_n 0.003457f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_505 N_A_299_47#_c_656_n N_VGND_c_1194_n 0.00812028f $X=3.25 $Y=0.995 $X2=0
+ $Y2=0
cc_506 N_A_299_47#_c_669_n N_VGND_c_1194_n 0.0318035f $X=2.475 $Y=0.395 $X2=0
+ $Y2=0
cc_507 N_A_299_47#_c_669_n A_415_47# 0.0102249f $X=2.475 $Y=0.395 $X2=-0.19
+ $Y2=-0.24
cc_508 N_A_299_47#_c_659_n A_415_47# 0.00167546f $X=2.56 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_509 N_CLK_M1005_g N_A_1093_47#_M1012_g 0.0216344f $X=6.21 $Y=0.445 $X2=0
+ $Y2=0
cc_510 N_CLK_c_764_n N_A_1093_47#_M1012_g 0.015147f $X=6.27 $Y=1.16 $X2=0 $Y2=0
cc_511 N_CLK_c_765_n N_A_1093_47#_M1012_g 3.04026e-19 $X=6.27 $Y=1.16 $X2=0
+ $Y2=0
cc_512 N_CLK_c_768_n N_A_1093_47#_c_868_n 0.0125511f $X=6.295 $Y=1.67 $X2=0
+ $Y2=0
cc_513 N_CLK_c_769_n N_A_1093_47#_c_868_n 0.0187438f $X=6.295 $Y=1.77 $X2=0
+ $Y2=0
cc_514 N_CLK_M1005_g N_A_1093_47#_c_863_n 0.0121932f $X=6.21 $Y=0.445 $X2=0
+ $Y2=0
cc_515 N_CLK_c_760_n N_A_1093_47#_c_863_n 0.00646156f $X=5.94 $Y=1.19 $X2=0
+ $Y2=0
cc_516 N_CLK_c_762_n N_A_1093_47#_c_863_n 0.00300199f $X=6.085 $Y=1.19 $X2=0
+ $Y2=0
cc_517 N_CLK_c_764_n N_A_1093_47#_c_863_n 0.00483458f $X=6.27 $Y=1.16 $X2=0
+ $Y2=0
cc_518 N_CLK_c_765_n N_A_1093_47#_c_863_n 0.0260027f $X=6.27 $Y=1.16 $X2=0 $Y2=0
cc_519 N_CLK_c_758_n N_A_1093_47#_c_864_n 6.54603e-19 $X=4.815 $Y=1.44 $X2=0
+ $Y2=0
cc_520 N_CLK_c_760_n N_A_1093_47#_c_864_n 0.00108081f $X=5.94 $Y=1.19 $X2=0
+ $Y2=0
cc_521 N_CLK_c_769_n N_A_1093_47#_c_882_n 0.00479018f $X=6.295 $Y=1.77 $X2=0
+ $Y2=0
cc_522 N_CLK_M1005_g N_A_1093_47#_c_865_n 0.00398268f $X=6.21 $Y=0.445 $X2=0
+ $Y2=0
cc_523 N_CLK_c_764_n N_A_1093_47#_c_865_n 4.08409e-19 $X=6.27 $Y=1.16 $X2=0
+ $Y2=0
cc_524 N_CLK_c_765_n N_A_1093_47#_c_865_n 0.00441122f $X=6.27 $Y=1.16 $X2=0
+ $Y2=0
cc_525 N_CLK_c_768_n N_A_1093_47#_c_870_n 0.00357759f $X=6.295 $Y=1.67 $X2=0
+ $Y2=0
cc_526 N_CLK_c_765_n N_A_1093_47#_c_870_n 6.41528e-19 $X=6.27 $Y=1.16 $X2=0
+ $Y2=0
cc_527 N_CLK_c_768_n N_A_1093_47#_c_872_n 0.00998304f $X=6.295 $Y=1.67 $X2=0
+ $Y2=0
cc_528 N_CLK_c_769_n N_A_1093_47#_c_872_n 0.0197237f $X=6.295 $Y=1.77 $X2=0
+ $Y2=0
cc_529 N_CLK_c_762_n N_A_1093_47#_c_872_n 0.00202388f $X=6.085 $Y=1.19 $X2=0
+ $Y2=0
cc_530 N_CLK_c_764_n N_A_1093_47#_c_872_n 0.00402174f $X=6.27 $Y=1.16 $X2=0
+ $Y2=0
cc_531 N_CLK_c_765_n N_A_1093_47#_c_872_n 0.0333702f $X=6.27 $Y=1.16 $X2=0 $Y2=0
cc_532 N_CLK_c_762_n N_A_1093_47#_c_866_n 0.00127984f $X=6.085 $Y=1.19 $X2=0
+ $Y2=0
cc_533 N_CLK_c_764_n N_A_1093_47#_c_866_n 0.00195414f $X=6.27 $Y=1.16 $X2=0
+ $Y2=0
cc_534 N_CLK_c_765_n N_A_1093_47#_c_866_n 0.0206769f $X=6.27 $Y=1.16 $X2=0 $Y2=0
cc_535 N_CLK_c_768_n N_A_1093_47#_c_867_n 0.0028705f $X=6.295 $Y=1.67 $X2=0
+ $Y2=0
cc_536 N_CLK_c_769_n N_VPWR_c_975_n 0.00181837f $X=6.295 $Y=1.77 $X2=0 $Y2=0
cc_537 N_CLK_M1001_g N_VPWR_c_978_n 0.0274117f $X=4.815 $Y=1.835 $X2=0 $Y2=0
cc_538 N_CLK_c_769_n N_VPWR_c_979_n 5.70534e-19 $X=6.295 $Y=1.77 $X2=0 $Y2=0
cc_539 N_CLK_c_769_n N_VPWR_c_980_n 0.00510113f $X=6.295 $Y=1.77 $X2=0 $Y2=0
cc_540 N_CLK_c_769_n N_VPWR_c_972_n 0.0067498f $X=6.295 $Y=1.77 $X2=0 $Y2=0
cc_541 N_CLK_c_757_n N_VGND_c_1181_n 0.00312892f $X=4.71 $Y=0.73 $X2=0 $Y2=0
cc_542 N_CLK_M1005_g N_VGND_c_1182_n 0.00441006f $X=6.21 $Y=0.445 $X2=0 $Y2=0
cc_543 N_CLK_c_757_n N_VGND_c_1184_n 0.00422112f $X=4.71 $Y=0.73 $X2=0 $Y2=0
cc_544 N_CLK_c_758_n N_VGND_c_1184_n 0.00230382f $X=4.815 $Y=1.44 $X2=0 $Y2=0
cc_545 N_CLK_M1005_g N_VGND_c_1184_n 0.00422112f $X=6.21 $Y=0.445 $X2=0 $Y2=0
cc_546 N_CLK_c_757_n N_VGND_c_1194_n 0.00711078f $X=4.71 $Y=0.73 $X2=0 $Y2=0
cc_547 N_CLK_c_758_n N_VGND_c_1194_n 0.00262886f $X=4.815 $Y=1.44 $X2=0 $Y2=0
cc_548 N_CLK_M1005_g N_VGND_c_1194_n 0.00596584f $X=6.21 $Y=0.445 $X2=0 $Y2=0
cc_549 N_A_1093_47#_c_870_n N_VPWR_M1013_d 3.89212e-19 $X=6.665 $Y=1.495 $X2=0
+ $Y2=0
cc_550 N_A_1093_47#_c_872_n N_VPWR_M1013_d 0.00764733f $X=6.665 $Y=1.79 $X2=0
+ $Y2=0
cc_551 N_A_1093_47#_c_868_n N_VPWR_c_975_n 0.00327647f $X=6.82 $Y=1.41 $X2=0
+ $Y2=0
cc_552 N_A_1093_47#_c_872_n N_VPWR_c_975_n 0.0191719f $X=6.665 $Y=1.79 $X2=0
+ $Y2=0
cc_553 N_A_1093_47#_c_869_n N_VPWR_c_977_n 0.00726717f $X=7.29 $Y=1.41 $X2=0
+ $Y2=0
cc_554 N_A_1093_47#_c_882_n N_VPWR_c_979_n 0.013449f $X=6.06 $Y=2.085 $X2=0
+ $Y2=0
cc_555 N_A_1093_47#_c_882_n N_VPWR_c_980_n 0.0113299f $X=6.06 $Y=2.085 $X2=0
+ $Y2=0
cc_556 N_A_1093_47#_c_872_n N_VPWR_c_980_n 0.00392738f $X=6.665 $Y=1.79 $X2=0
+ $Y2=0
cc_557 N_A_1093_47#_c_868_n N_VPWR_c_983_n 0.00681089f $X=6.82 $Y=1.41 $X2=0
+ $Y2=0
cc_558 N_A_1093_47#_c_869_n N_VPWR_c_983_n 0.00673617f $X=7.29 $Y=1.41 $X2=0
+ $Y2=0
cc_559 N_A_1093_47#_c_872_n N_VPWR_c_983_n 3.86084e-19 $X=6.665 $Y=1.79 $X2=0
+ $Y2=0
cc_560 N_A_1093_47#_M1019_d N_VPWR_c_972_n 0.00462612f $X=5.915 $Y=1.845 $X2=0
+ $Y2=0
cc_561 N_A_1093_47#_c_868_n N_VPWR_c_972_n 0.0119747f $X=6.82 $Y=1.41 $X2=0
+ $Y2=0
cc_562 N_A_1093_47#_c_869_n N_VPWR_c_972_n 0.0128271f $X=7.29 $Y=1.41 $X2=0
+ $Y2=0
cc_563 N_A_1093_47#_c_882_n N_VPWR_c_972_n 0.00637602f $X=6.06 $Y=2.085 $X2=0
+ $Y2=0
cc_564 N_A_1093_47#_c_872_n N_VPWR_c_972_n 0.00878273f $X=6.665 $Y=1.79 $X2=0
+ $Y2=0
cc_565 N_A_1093_47#_M1012_g N_GCLK_c_1140_n 0.00432012f $X=6.795 $Y=0.56 $X2=0
+ $Y2=0
cc_566 N_A_1093_47#_c_863_n N_GCLK_c_1140_n 0.00647845f $X=6.58 $Y=0.7 $X2=0
+ $Y2=0
cc_567 N_A_1093_47#_M1014_g N_GCLK_c_1134_n 0.0142286f $X=7.265 $Y=0.56 $X2=0
+ $Y2=0
cc_568 N_A_1093_47#_c_871_n N_GCLK_c_1134_n 0.00632886f $X=6.75 $Y=1.185 $X2=0
+ $Y2=0
cc_569 N_A_1093_47#_M1012_g N_GCLK_c_1135_n 0.00148642f $X=6.795 $Y=0.56 $X2=0
+ $Y2=0
cc_570 N_A_1093_47#_c_863_n N_GCLK_c_1135_n 0.00502168f $X=6.58 $Y=0.7 $X2=0
+ $Y2=0
cc_571 N_A_1093_47#_c_865_n N_GCLK_c_1135_n 0.00646488f $X=6.665 $Y=1.055 $X2=0
+ $Y2=0
cc_572 N_A_1093_47#_c_871_n N_GCLK_c_1135_n 0.0141305f $X=6.75 $Y=1.185 $X2=0
+ $Y2=0
cc_573 N_A_1093_47#_c_867_n N_GCLK_c_1135_n 0.00297398f $X=7.265 $Y=1.217 $X2=0
+ $Y2=0
cc_574 N_A_1093_47#_c_869_n N_GCLK_c_1137_n 0.0164256f $X=7.29 $Y=1.41 $X2=0
+ $Y2=0
cc_575 N_A_1093_47#_c_871_n N_GCLK_c_1137_n 0.00346944f $X=6.75 $Y=1.185 $X2=0
+ $Y2=0
cc_576 N_A_1093_47#_c_868_n N_GCLK_c_1138_n 0.00144243f $X=6.82 $Y=1.41 $X2=0
+ $Y2=0
cc_577 N_A_1093_47#_c_869_n N_GCLK_c_1138_n 0.00186704f $X=7.29 $Y=1.41 $X2=0
+ $Y2=0
cc_578 N_A_1093_47#_c_870_n N_GCLK_c_1138_n 6.49246e-19 $X=6.665 $Y=1.495 $X2=0
+ $Y2=0
cc_579 N_A_1093_47#_c_871_n N_GCLK_c_1138_n 0.0185691f $X=6.75 $Y=1.185 $X2=0
+ $Y2=0
cc_580 N_A_1093_47#_c_872_n N_GCLK_c_1138_n 0.0114062f $X=6.665 $Y=1.79 $X2=0
+ $Y2=0
cc_581 N_A_1093_47#_c_867_n N_GCLK_c_1138_n 0.00150749f $X=7.265 $Y=1.217 $X2=0
+ $Y2=0
cc_582 N_A_1093_47#_M1012_g N_GCLK_c_1157_n 0.00306708f $X=6.795 $Y=0.56 $X2=0
+ $Y2=0
cc_583 N_A_1093_47#_c_871_n N_GCLK_c_1157_n 0.00260368f $X=6.75 $Y=1.185 $X2=0
+ $Y2=0
cc_584 N_A_1093_47#_c_868_n GCLK 0.00666419f $X=6.82 $Y=1.41 $X2=0 $Y2=0
cc_585 N_A_1093_47#_c_869_n GCLK 0.0162476f $X=7.29 $Y=1.41 $X2=0 $Y2=0
cc_586 N_A_1093_47#_c_872_n GCLK 0.0283421f $X=6.665 $Y=1.79 $X2=0 $Y2=0
cc_587 N_A_1093_47#_M1014_g GCLK 0.00491155f $X=7.265 $Y=0.56 $X2=0 $Y2=0
cc_588 N_A_1093_47#_c_869_n GCLK 0.00278773f $X=7.29 $Y=1.41 $X2=0 $Y2=0
cc_589 N_A_1093_47#_c_871_n GCLK 0.017086f $X=6.75 $Y=1.185 $X2=0 $Y2=0
cc_590 N_A_1093_47#_c_867_n GCLK 0.0124258f $X=7.265 $Y=1.217 $X2=0 $Y2=0
cc_591 N_A_1093_47#_c_863_n N_VGND_M1005_d 0.00973459f $X=6.58 $Y=0.7 $X2=0
+ $Y2=0
cc_592 N_A_1093_47#_c_865_n N_VGND_M1005_d 0.00126753f $X=6.665 $Y=1.055 $X2=0
+ $Y2=0
cc_593 N_A_1093_47#_M1012_g N_VGND_c_1182_n 0.00441006f $X=6.795 $Y=0.56 $X2=0
+ $Y2=0
cc_594 N_A_1093_47#_c_863_n N_VGND_c_1182_n 0.0249591f $X=6.58 $Y=0.7 $X2=0
+ $Y2=0
cc_595 N_A_1093_47#_M1014_g N_VGND_c_1183_n 0.00438629f $X=7.265 $Y=0.56 $X2=0
+ $Y2=0
cc_596 N_A_1093_47#_c_874_n N_VGND_c_1184_n 0.0116015f $X=5.59 $Y=0.46 $X2=0
+ $Y2=0
cc_597 N_A_1093_47#_c_863_n N_VGND_c_1184_n 0.009944f $X=6.58 $Y=0.7 $X2=0 $Y2=0
cc_598 N_A_1093_47#_M1012_g N_VGND_c_1189_n 0.00507199f $X=6.795 $Y=0.56 $X2=0
+ $Y2=0
cc_599 N_A_1093_47#_M1014_g N_VGND_c_1189_n 0.00436487f $X=7.265 $Y=0.56 $X2=0
+ $Y2=0
cc_600 N_A_1093_47#_c_863_n N_VGND_c_1189_n 0.00107125f $X=6.58 $Y=0.7 $X2=0
+ $Y2=0
cc_601 N_A_1093_47#_M1004_s N_VGND_c_1194_n 0.00426262f $X=5.465 $Y=0.235 $X2=0
+ $Y2=0
cc_602 N_A_1093_47#_M1012_g N_VGND_c_1194_n 0.00906461f $X=6.795 $Y=0.56 $X2=0
+ $Y2=0
cc_603 N_A_1093_47#_M1014_g N_VGND_c_1194_n 0.00701551f $X=7.265 $Y=0.56 $X2=0
+ $Y2=0
cc_604 N_A_1093_47#_c_874_n N_VGND_c_1194_n 0.00642843f $X=5.59 $Y=0.46 $X2=0
+ $Y2=0
cc_605 N_A_1093_47#_c_863_n N_VGND_c_1194_n 0.0213501f $X=6.58 $Y=0.7 $X2=0
+ $Y2=0
cc_606 N_A_1093_47#_c_863_n A_1185_47# 0.00163533f $X=6.58 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_607 N_VPWR_c_972_n A_117_369# 0.00184697f $X=7.59 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_608 N_VPWR_c_972_n N_A_27_47#_M1002_d 0.00419357f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_609 N_VPWR_c_974_n N_A_27_47#_c_1079_n 0.0213176f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_610 N_VPWR_c_974_n N_A_27_47#_c_1091_n 0.027538f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_611 N_VPWR_c_984_n N_A_27_47#_c_1091_n 0.0122125f $X=2.52 $Y=2.44 $X2=0 $Y2=0
cc_612 N_VPWR_c_972_n N_A_27_47#_c_1091_n 0.00756493f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_613 N_VPWR_c_984_n N_A_27_47#_c_1100_n 0.0332722f $X=2.52 $Y=2.44 $X2=0 $Y2=0
cc_614 N_VPWR_c_972_n N_A_27_47#_c_1100_n 0.0203569f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_615 N_VPWR_c_972_n A_410_413# 0.00736425f $X=7.59 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_616 N_VPWR_c_972_n N_GCLK_M1003_s 0.00444633f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_617 N_VPWR_M1011_d N_GCLK_c_1137_n 0.00410054f $X=7.38 $Y=1.485 $X2=0 $Y2=0
cc_618 N_VPWR_c_977_n N_GCLK_c_1137_n 0.0206716f $X=7.525 $Y=2 $X2=0 $Y2=0
cc_619 N_VPWR_c_977_n GCLK 0.039075f $X=7.525 $Y=2 $X2=0 $Y2=0
cc_620 N_VPWR_c_983_n GCLK 0.015413f $X=7.44 $Y=2.72 $X2=0 $Y2=0
cc_621 N_VPWR_c_972_n GCLK 0.00946403f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_622 A_117_369# N_A_27_47#_c_1079_n 0.0028312f $X=0.585 $Y=1.845 $X2=0 $Y2=0
cc_623 A_117_369# N_A_27_47#_c_1091_n 7.5302e-19 $X=0.585 $Y=1.845 $X2=0 $Y2=0
cc_624 A_117_369# N_A_27_47#_c_1100_n 0.00189004f $X=0.585 $Y=1.845 $X2=0.215
+ $Y2=2
cc_625 N_A_27_47#_c_1080_n N_VGND_M1020_d 9.37209e-19 $X=1.115 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_626 N_A_27_47#_c_1081_n N_VGND_M1020_d 6.9272e-19 $X=0.72 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_627 N_A_27_47#_c_1078_n N_VGND_c_1186_n 0.0173928f $X=0.26 $Y=0.43 $X2=0
+ $Y2=0
cc_628 N_A_27_47#_c_1081_n N_VGND_c_1186_n 0.00260613f $X=0.72 $Y=0.7 $X2=0
+ $Y2=0
cc_629 N_A_27_47#_c_1080_n N_VGND_c_1187_n 0.00341938f $X=1.115 $Y=0.7 $X2=0
+ $Y2=0
cc_630 N_A_27_47#_c_1104_n N_VGND_c_1187_n 0.0120906f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_631 N_A_27_47#_c_1078_n N_VGND_c_1190_n 0.0146378f $X=0.26 $Y=0.43 $X2=0
+ $Y2=0
cc_632 N_A_27_47#_c_1081_n N_VGND_c_1190_n 0.0193989f $X=0.72 $Y=0.7 $X2=0 $Y2=0
cc_633 N_A_27_47#_c_1104_n N_VGND_c_1190_n 0.0116788f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_634 N_A_27_47#_M1020_s N_VGND_c_1194_n 0.00286466f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_635 N_A_27_47#_M1023_d N_VGND_c_1194_n 0.00463742f $X=1.02 $Y=0.235 $X2=0
+ $Y2=0
cc_636 N_A_27_47#_c_1078_n N_VGND_c_1194_n 0.00977915f $X=0.26 $Y=0.43 $X2=0
+ $Y2=0
cc_637 N_A_27_47#_c_1080_n N_VGND_c_1194_n 0.00569248f $X=1.115 $Y=0.7 $X2=0
+ $Y2=0
cc_638 N_A_27_47#_c_1081_n N_VGND_c_1194_n 0.00628516f $X=0.72 $Y=0.7 $X2=0
+ $Y2=0
cc_639 N_A_27_47#_c_1104_n N_VGND_c_1194_n 0.00681108f $X=1.2 $Y=0.42 $X2=0
+ $Y2=0
cc_640 N_GCLK_c_1134_n N_VGND_M1014_d 0.00498894f $X=7.49 $Y=0.8 $X2=0 $Y2=0
cc_641 N_GCLK_c_1134_n N_VGND_c_1183_n 0.0128502f $X=7.49 $Y=0.8 $X2=0 $Y2=0
cc_642 N_GCLK_c_1134_n N_VGND_c_1189_n 0.00260889f $X=7.49 $Y=0.8 $X2=0 $Y2=0
cc_643 N_GCLK_c_1157_n N_VGND_c_1189_n 0.0183042f $X=7.005 $Y=0.36 $X2=0 $Y2=0
cc_644 N_GCLK_c_1134_n N_VGND_c_1193_n 0.00197242f $X=7.49 $Y=0.8 $X2=0 $Y2=0
cc_645 N_GCLK_M1012_s N_VGND_c_1194_n 0.00263739f $X=6.87 $Y=0.235 $X2=0 $Y2=0
cc_646 N_GCLK_c_1134_n N_VGND_c_1194_n 0.00898735f $X=7.49 $Y=0.8 $X2=0 $Y2=0
cc_647 N_GCLK_c_1157_n N_VGND_c_1194_n 0.0121135f $X=7.005 $Y=0.36 $X2=0 $Y2=0
cc_648 N_VGND_c_1194_n A_415_47# 0.00329302f $X=7.59 $Y=0 $X2=-0.19 $Y2=-0.24
cc_649 N_VGND_c_1194_n A_1185_47# 0.00239227f $X=7.59 $Y=0 $X2=-0.19 $Y2=-0.24
