* NGSPICE file created from sky130_fd_sc_hdll__mux2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__mux2_4 A0 A1 S VGND VNB VPB VPWR X
M1000 VPWR a_424_297# X VPB phighvt w=1e+06u l=180000u
+  ad=1.195e+12p pd=1.039e+07u as=5.8e+11p ps=5.16e+06u
M1001 a_424_297# A0 a_334_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.4e+11p pd=2.68e+06u as=5.4e+11p ps=5.08e+06u
M1002 X a_424_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_424_297# VGND VNB nshort w=650000u l=150000u
+  ad=4.16e+11p pd=3.88e+06u as=8.3525e+11p ps=7.77e+06u
M1004 VPWR S a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1005 VGND a_424_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_530_47# A1 a_424_297# VNB nshort w=650000u l=150000u
+  ad=5.8175e+11p pd=3.09e+06u as=2.405e+11p ps=2.04e+06u
M1007 VPWR a_424_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND S a_530_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_424_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND S a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1011 a_424_297# A0 a_226_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=5.525e+11p ps=3e+06u
M1012 VPWR S a_334_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_424_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_222_297# A1 a_424_297# VPB phighvt w=1e+06u l=180000u
+  ad=6e+11p pd=5.2e+06u as=0p ps=0u
M1015 a_226_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_222_297# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_424_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

