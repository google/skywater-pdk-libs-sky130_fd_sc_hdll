* File: sky130_fd_sc_hdll__a211o_2.spice
* Created: Thu Aug 27 18:51:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a211o_2.pex.spice"
.subckt sky130_fd_sc_hdll__a211o_2  VNB VPB A2 A1 B1 C1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_79_21#_M1008_g N_X_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.10725 PD=1.82 PS=0.98 NRD=0 NRS=8.76 M=1 R=4.33333 SA=75000.2
+ SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A_79_21#_M1011_g N_X_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.30225 AS=0.10725 PD=1.58 PS=0.98 NRD=8.304 NRS=0.456 M=1 R=4.33333
+ SA=75000.7 SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1003 A_421_47# N_A2_M1003_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.65
+ AD=0.079625 AS=0.30225 PD=0.895 PS=1.58 NRD=12.456 NRS=47.988 M=1 R=4.33333
+ SA=75001.7 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1010 N_A_79_21#_M1010_d N_A1_M1010_g A_421_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.128375 AS=0.079625 PD=1.045 PS=0.895 NRD=9.228 NRS=12.456 M=1 R=4.33333
+ SA=75002.1 SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1002_d N_B1_M1002_g N_A_79_21#_M1010_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.128375 PD=1.04 PS=1.045 NRD=15.684 NRS=11.988 M=1 R=4.33333
+ SA=75002.7 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1005 N_A_79_21#_M1005_d N_C1_M1005_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.12675 PD=1.92 PS=1.04 NRD=8.304 NRS=4.608 M=1 R=4.33333
+ SA=75003.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_79_21#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A_79_21#_M1006_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_A2_M1007_g N_A_319_297#_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.2 AS=0.32 PD=1.4 PS=2.64 NRD=13.7703 NRS=10.8153 M=1 R=5.55556 SA=90000.2
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1004 N_A_319_297#_M1004_d N_A1_M1004_g N_VPWR_M1007_d VPB PHIGHVT L=0.18 W=1
+ AD=0.18 AS=0.2 PD=1.36 PS=1.4 NRD=12.7853 NRS=9.8303 M=1 R=5.55556 SA=90000.8
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1001 A_643_297# N_B1_M1001_g N_A_319_297#_M1004_d VPB PHIGHVT L=0.18 W=1
+ AD=0.115 AS=0.18 PD=1.23 PS=1.36 NRD=11.8003 NRS=2.9353 M=1 R=5.55556
+ SA=90001.3 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1009 N_A_79_21#_M1009_d N_C1_M1009_g A_643_297# VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.115 PD=2.54 PS=1.23 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90001.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
pX13_noxref noxref_14 A2 A2 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__a211o_2.pxi.spice"
*
.ends
*
*
