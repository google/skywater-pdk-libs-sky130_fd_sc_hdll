* NGSPICE file created from sky130_fd_sc_hdll__or3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__or3_4 A B C VGND VNB VPB VPWR X
M1000 a_211_297# B a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u
M1001 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=3.77e+11p pd=3.76e+06u as=1.20575e+12p ps=8.91e+06u
M1002 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=1.48e+12p pd=8.96e+06u as=5.8e+11p ps=5.16e+06u
M1003 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_117_297# C a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1006 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1007 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND C a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A a_211_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

