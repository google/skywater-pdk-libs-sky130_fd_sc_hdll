* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__xnor3_2 A B C VGND VNB VPB VPWR X
X0 a_477_49# a_885_297# a_1003_297# VNB sky130_fd_pr__nfet_01v8 w=600000u l=150000u
X1 a_79_21# a_328_93# a_453_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 a_1286_297# B a_453_325# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X3 a_79_21# a_328_93# a_477_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X4 VGND C a_328_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_477_49# a_885_297# a_1286_297# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X6 a_1003_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VPWR B a_885_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_477_49# C a_79_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 a_453_325# a_885_297# a_1286_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_453_325# C a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X13 VPWR a_1003_297# a_1286_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 a_1003_297# B a_477_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X15 a_1003_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 VPWR C a_328_93# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X17 a_1003_297# B a_453_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 a_453_325# a_885_297# a_1003_297# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X19 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_1286_297# B a_477_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 VGND B a_885_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VGND a_1003_297# a_1286_297# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X23 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
