* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__o22ai_2 B2 B1 Y A1 A2 VPB VNB VGND VPWR
M1000 Y A2 a_515_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u
M1001 VPWR B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u
M1002 a_27_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=1.2415e+12p pd=1.032e+07u as=4.81e+11p ps=4.08e+06u
M1003 a_27_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=4.81e+11p pd=4.08e+06u as=0p ps=0u
M1007 a_27_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_515_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A1 a_515_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_515_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand2_1 Y B A VPB VNB VGND VPWR
M1000 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=5.4e+11p ps=5.08e+06u
M1001 Y A a_123_47# VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=1.755e+11p ps=1.84e+06u
M1002 a_123_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1003 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor3_4 A C B Y VPB VNB VGND VPWR
M1000 Y C VGND VNB nshort w=650000u l=150000u
+  ad=1.248e+12p pd=1.164e+07u as=1.4235e+12p ps=1.348e+07u
M1001 a_497_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=1.43e+12p ps=1.286e+07u
M1002 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1004 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y C a_497_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1007 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_497_297# C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y C a_497_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_297# B a_497_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_497_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_497_297# C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_297# B a_497_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a21bo_1 X A1 B1_N A2 VNB VPB VGND VPWR
M1000 a_326_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.65e+11p pd=5.13e+06u as=6.834e+11p ps=6.52e+06u
M1001 a_412_47# A1 a_235_297# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=1.755e+11p ps=1.84e+06u
M1002 VPWR B1_N a_27_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1003 a_235_297# a_27_413# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=9.0705e+11p ps=5.49e+06u
M1004 VGND B1_N a_27_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.323e+11p ps=1.47e+06u
M1005 X a_235_297# VGND VNB nshort w=650000u l=150000u
+  ad=2.4375e+11p pd=2.05e+06u as=0p ps=0u
M1006 VGND A2 a_412_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A1 a_326_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_326_297# a_27_413# a_235_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.75e+11p ps=2.55e+06u
M1009 X a_235_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.85e+11p pd=2.77e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand2b_2 B Y A_N VNB VPB VGND VPWR
M1000 a_215_47# a_27_93# Y VNB nshort w=650000u l=150000u
+  ad=5.135e+11p pd=5.48e+06u as=1.755e+11p ps=1.84e+06u
M1001 VPWR a_27_93# Y VPB phighvt w=1e+06u l=180000u
+  ad=1.0628e+12p pd=8.23e+06u as=6.5e+11p ps=5.3e+06u
M1002 Y a_27_93# a_215_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_215_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.172e+11p ps=3.3e+06u
M1004 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND B a_215_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A_N a_27_93# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1007 Y a_27_93# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A_N a_27_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
.ends
.subckt sky130_fd_sc_hdll__a31oi_1 VGND VPWR Y B1 A2 A1 A3 VPB VNB
M1000 VPWR A2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.95e+11p pd=5.19e+06u as=6.35e+11p ps=5.27e+06u
M1001 a_117_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_203_47# A2 a_119_47# VNB nshort w=650000u l=150000u
+  ad=2.3075e+11p pd=2.01e+06u as=1.755e+11p ps=1.84e+06u
M1003 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=5.2e+11p pd=4.2e+06u as=2.4375e+11p ps=2.05e+06u
M1004 a_117_297# A3 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_119_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1007 Y A1 a_203_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__mux2i_1 A1 S A0 Y VPB VNB VGND VPWR
M1000 Y A0 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=5.6e+11p ps=5.12e+06u
M1001 a_27_297# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.2e+11p ps=5.64e+06u
M1002 a_207_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=3.575e+11p pd=3.7e+06u as=1.755e+11p ps=1.84e+06u
M1003 VGND S a_303_205# VNB nshort w=650000u l=150000u
+  ad=3.445e+11p pd=3.66e+06u as=2.275e+11p ps=2e+06u
M1004 VPWR S a_303_205# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3e+11p ps=2.6e+06u
M1005 Y A0 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.835e+11p ps=3.78e+06u
M1006 VPWR a_303_205# a_215_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=4.5e+11p ps=2.9e+06u
M1007 a_215_297# A1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_303_205# a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_207_47# S VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__clkbuf_16 X A VNB VPB VGND VPWR
M1000 VGND a_118_297# X VNB nshort w=420000u l=150000u
+  ad=1.4679e+12p pd=1.623e+07u as=1.1298e+12p ps=1.21e+07u
M1001 VGND a_118_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 X a_118_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_118_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.4e+12p pd=2.08e+07u as=3.245e+12p ps=2.849e+07u
M1004 VPWR a_118_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_118_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_118_297# A VGND VNB nshort w=420000u l=150000u
+  ad=2.772e+11p pd=3e+06u as=0p ps=0u
M1007 VGND A a_118_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_118_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_118_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_118_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_118_297# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_118_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_118_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6e+11p pd=5.2e+06u as=0p ps=0u
M1014 a_118_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_118_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_118_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_118_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_118_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_118_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_118_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_118_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 X a_118_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A a_118_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X a_118_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_118_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 X a_118_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_118_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR a_118_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_118_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A a_118_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 X a_118_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 X a_118_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 X a_118_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR A a_118_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 X a_118_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND a_118_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 X a_118_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 X a_118_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND a_118_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o211ai_2 A1 A2 B1 Y C1 VNB VPB VGND VPWR
M1000 a_316_47# B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=6.63e+11p pd=5.94e+06u as=6.175e+11p ps=5.8e+06u
M1001 Y A2 a_527_297# VPB phighvt w=1e+06u l=180000u
+  ad=9e+11p pd=7.8e+06u as=8.5e+11p ps=7.7e+06u
M1002 a_27_47# B1 a_316_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=1.15e+12p pd=1.03e+07u as=0p ps=0u
M1004 a_316_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=6.1425e+11p ps=5.79e+06u
M1005 VPWR A1 a_527_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_47# C1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.145e+11p ps=1.96e+06u
M1008 a_527_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_316_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A1 a_316_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A2 a_316_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_527_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y C1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y C1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or2b_1 A B_N X VGND VPWR VNB VPB
M1000 VGND B_N a_27_53# VNB nshort w=420000u l=150000u
+  ad=5.7225e+11p pd=4.52e+06u as=1.302e+11p ps=1.46e+06u
M1001 X a_229_297# VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1002 a_27_53# B_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=4.241e+11p ps=4.1e+06u
M1003 a_319_297# a_27_53# a_229_297# VPB phighvt w=420000u l=180000u
+  ad=9.66e+10p pd=1.3e+06u as=1.134e+11p ps=1.38e+06u
M1004 VGND A a_229_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1005 VPWR A a_319_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_229_297# a_27_53# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_229_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__dlrtn_1 RESET_B D GATE_N Q VGND VPWR VPB VNB
M1000 VGND a_750_21# a_708_47# VNB nshort w=420000u l=150000u
+  ad=5.6425e+11p pd=6.14e+06u as=8.82e+10p ps=1.26e+06u
M1001 VPWR GATE_N a_27_363# VPB phighvt w=640000u l=180000u
+  ad=1.131e+12p pd=9.75e+06u as=1.728e+11p ps=1.82e+06u
M1002 a_203_47# a_27_363# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1003 VPWR a_750_21# a_702_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1004 a_503_369# a_319_369# VPWR VPB phighvt w=640000u l=180000u
+  ad=2.021e+11p pd=1.97e+06u as=0p ps=0u
M1005 a_708_47# a_203_47# a_604_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.58e+06u
M1006 Q a_750_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1007 VGND D a_319_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1008 VPWR D a_319_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1009 VGND RESET_B a_981_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.6575e+11p ps=1.81e+06u
M1010 a_604_47# a_27_363# a_500_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.58e+06u
M1011 Q a_750_21# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1012 VPWR RESET_B a_750_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1013 a_981_47# a_604_47# a_750_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1014 VGND GATE_N a_27_363# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1015 a_702_413# a_27_363# a_604_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1016 a_203_47# a_27_363# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1017 a_604_47# a_203_47# a_503_369# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_500_47# a_319_369# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_750_21# a_604_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__clkmux2_2 VGND VPWR S A1 A0 X VPB VNB
M1000 VPWR a_79_199# X VPB phighvt w=1e+06u l=180000u
+  ad=1.0664e+12p pd=8.08e+06u as=2.9e+11p ps=2.58e+06u
M1001 VGND a_741_21# a_570_47# VNB nshort w=420000u l=150000u
+  ad=6.32e+11p pd=5.72e+06u as=3.591e+11p ps=2.55e+06u
M1002 a_335_309# S VPWR VPB phighvt w=940000u l=180000u
+  ad=3.901e+11p pd=2.71e+06u as=0p ps=0u
M1003 X a_79_199# VGND VNB nshort w=520000u l=150000u
+  ad=1.404e+11p pd=1.58e+06u as=0p ps=0u
M1004 a_741_21# S VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1005 X a_79_199# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_691_309# A1 a_79_199# VPB phighvt w=940000u l=180000u
+  ad=2.444e+11p pd=2.4e+06u as=9.447e+11p ps=3.89e+06u
M1007 a_570_47# A0 a_79_199# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.121e+11p ps=1.85e+06u
M1008 a_337_47# S VGND VNB nshort w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=0p ps=0u
M1009 a_741_21# S VPWR VPB phighvt w=940000u l=180000u
+  ad=2.726e+11p pd=2.46e+06u as=0p ps=0u
M1010 VGND a_79_199# X VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_79_199# A0 a_335_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_741_21# a_691_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_79_199# A1 a_337_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or2_8 X A B VNB VPB VGND VPWR
M1000 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.71e+12p pd=1.542e+07u as=8.5e+11p ps=7.7e+06u
M1001 VGND A a_123_47# VNB nshort w=650000u l=150000u
+  ad=1.963e+12p pd=1.514e+07u as=3.51e+11p ps=3.68e+06u
M1002 X a_123_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=0p ps=0u
M1003 VGND a_123_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.02e+11p ps=7.36e+06u
M1004 a_123_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_123_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_297# B a_123_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1007 VPWR a_123_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_123_47# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_123_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_123_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_123_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_123_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_123_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_123_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B a_123_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_123_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_123_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_123_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_123_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_123_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 X a_123_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_123_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o21ai_2 B1 Y A2 A1 VGND VPWR VPB VNB
M1000 a_29_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=8.7425e+11p pd=7.89e+06u as=5.005e+11p ps=4.14e+06u
M1001 Y B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6e+11p pd=5.2e+06u as=9.95e+11p ps=7.99e+06u
M1002 a_120_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6.7e+11p pd=5.34e+06u as=0p ps=0u
M1003 a_120_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y B1 a_29_47# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=0p ps=0u
M1005 VPWR A1 a_120_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_29_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A2 a_120_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A1 a_29_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_29_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A2 a_29_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and3_4 A B C X VNB VPB VGND VPWR
M1000 X a_85_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6e+11p pd=5.2e+06u as=1.435e+12p ps=1.087e+07u
M1001 a_85_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6.1e+11p pd=5.22e+06u as=0p ps=0u
M1002 a_185_47# A a_85_297# VNB nshort w=650000u l=150000u
+  ad=3.2175e+11p pd=2.29e+06u as=1.9825e+11p ps=1.91e+06u
M1003 X a_85_297# VGND VNB nshort w=650000u l=150000u
+  ad=4.615e+11p pd=4.02e+06u as=7.085e+11p ps=6.08e+06u
M1004 VPWR a_85_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_85_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_314_47# B a_185_47# VNB nshort w=650000u l=150000u
+  ad=1.365e+11p pd=1.72e+06u as=0p ps=0u
M1007 VGND C a_314_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_85_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR C a_85_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_85_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_85_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_85_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A a_85_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__clkbuf_4 X A VGND VPWR VPB VNB
M1000 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=4.011e+11p pd=4.43e+06u as=1.323e+11p ps=1.47e+06u
M1001 X a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=2.982e+11p pd=3.1e+06u as=0p ps=0u
M1002 X a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=9.6e+11p pd=7.92e+06u as=2.75e+11p ps=2.55e+06u
M1004 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=6e+11p ps=5.2e+06u
M1005 VGND a_27_47# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_27_47# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__clkinv_4 A Y VNB VPB VPWR VGND
M1000 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=1.27e+12p pd=1.054e+07u as=9e+11p ps=7.8e+06u
M1001 Y A VGND VNB nshort w=420000u l=150000u
+  ad=2.772e+11p pd=3e+06u as=4.851e+11p ps=4.83e+06u
M1002 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sdfstp_4 CLK D SCD Q SCE SET_B VPWR VGND VPB VNB
M1000 VPWR SET_B a_1229_21# VPB phighvt w=420000u l=180000u
+  ad=2.3974e+12p pd=2.127e+07u as=1.722e+11p ps=1.66e+06u
M1001 VGND a_349_21# a_295_47# VNB nshort w=420000u l=150000u
+  ad=1.73245e+12p pd=1.7e+07u as=1.134e+11p ps=1.38e+06u
M1002 a_2067_47# a_1951_295# a_1995_47# VNB nshort w=420000u l=150000u
+  ad=2.016e+11p pd=1.8e+06u as=8.82e+10p ps=1.26e+06u
M1003 a_1745_329# SET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=4.746e+11p pd=4.26e+06u as=0p ps=0u
M1004 a_1951_295# a_1745_329# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1005 a_1995_47# a_693_369# a_1745_329# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.332e+11p ps=2.5e+06u
M1006 a_1891_413# a_877_369# a_1745_329# VPB phighvt w=420000u l=180000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1007 VGND SCE a_349_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1008 a_1075_413# a_877_369# a_201_47# VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=2.99e+11p ps=3.24e+06u
M1009 VGND a_2447_47# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1010 VPWR SCD a_27_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=3.456e+11p ps=3.64e+06u
M1011 a_1229_21# a_1075_413# VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Q a_2447_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1013 Q a_2447_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR SCE a_349_21# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1015 VGND SET_B a_2067_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_2447_47# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND SET_B a_1467_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1018 a_877_369# a_693_369# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1019 VGND a_1229_21# a_1177_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1020 VPWR a_1951_295# a_1891_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND CLK a_693_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1022 a_1951_295# a_1745_329# VGND VNB nshort w=420000u l=150000u
+  ad=1.596e+11p pd=1.6e+06u as=0p ps=0u
M1023 a_1654_47# a_1075_413# VGND VNB nshort w=640000u l=150000u
+  ad=5.088e+11p pd=2.87e+06u as=0p ps=0u
M1024 a_1467_47# a_1075_413# a_1229_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.512e+11p ps=1.56e+06u
M1025 Q a_2447_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_27_369# a_349_21# a_201_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_119_47# SCD VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1028 a_1177_47# a_877_369# a_1075_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1029 VPWR a_2447_47# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND a_1745_329# a_2447_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1031 a_877_369# a_693_369# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1032 a_1663_329# a_1075_413# VPWR VPB phighvt w=840000u l=180000u
+  ad=1.932e+11p pd=2.14e+06u as=0p ps=0u
M1033 a_1075_413# a_693_369# a_201_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.646e+11p ps=2.94e+06u
M1034 a_1745_329# a_693_369# a_1663_329# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_295_47# D a_201_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND a_2447_47# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_201_47# SCE a_119_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 Q a_2447_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_211_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=1.472e+11p pd=1.74e+06u as=0p ps=0u
M1040 VPWR a_1745_329# a_2447_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1041 a_201_47# D a_211_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_1169_413# a_693_369# a_1075_413# VPB phighvt w=420000u l=180000u
+  ad=1.596e+11p pd=1.6e+06u as=0p ps=0u
M1043 VPWR a_1229_21# a_1169_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VPWR CLK a_693_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1045 a_1745_329# a_877_369# a_1654_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a2bb2oi_1 A1_N Y VGND VPWR B2 B1 A2_N VPB VNB
M1000 a_521_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=2.6e+11p ps=2.1e+06u
M1001 a_119_47# A2_N a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=2.3e+11p ps=2.46e+06u
M1002 a_117_297# A1_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.7e+11p ps=5.14e+06u
M1003 VGND A2_N a_119_47# VNB nshort w=650000u l=150000u
+  ad=9.425e+11p pd=6.8e+06u as=2.145e+11p ps=1.96e+06u
M1004 Y a_119_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_409_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6.4e+11p pd=5.28e+06u as=0p ps=0u
M1006 a_409_297# a_119_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1007 a_119_47# A1_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND B1 a_521_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR B2 a_409_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor4bb_2 D_N C_N A Y B VNB VPB VGND VPWR
M1000 Y a_216_93# VGND VNB nshort w=650000u l=150000u
+  ad=9.295e+11p pd=8.06e+06u as=1.29595e+12p ps=1.29e+07u
M1001 a_823_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.65e+11p pd=7.73e+06u as=5.43625e+11p ps=5.26e+06u
M1002 a_216_93# C_N VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1003 a_433_297# a_216_93# a_343_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=8.3e+11p ps=7.66e+06u
M1004 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_27_93# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_823_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR D_N a_27_93# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1009 a_823_297# B a_433_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y a_27_93# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_343_297# a_27_93# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1012 VGND a_216_93# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_216_93# C_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1014 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_433_297# B a_823_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y a_27_93# a_343_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_343_297# a_216_93# a_433_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND D_N a_27_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
.ends
.subckt sky130_fd_sc_hdll__isobufsrc_2 A SLEEP X VPB VNB VGND VPWR
M1000 VPWR SLEEP a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=4.034e+11p pd=3.96e+06u as=8.5e+11p ps=7.7e+06u
M1001 VGND A a_271_21# VNB nshort w=420000u l=150000u
+  ad=6.5345e+11p pd=6.97e+06u as=1.092e+11p ps=1.36e+06u
M1002 a_27_297# a_271_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1003 X a_271_21# a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=4.81e+11p pd=4.08e+06u as=0p ps=0u
M1005 VGND a_271_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A a_271_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1007 a_27_297# SLEEP VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_271_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND SLEEP X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sdfxbp_1 VGND VPWR SCD Q_N D SCE CLK Q VNB VPB
M1000 VPWR a_1179_183# a_1111_413# VPB phighvt w=420000u l=180000u
+  ad=1.70555e+12p pd=1.505e+07u as=1.47e+11p ps=1.54e+06u
M1001 a_211_363# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.3638e+12p ps=1.273e+07u
M1002 Q a_1653_315# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1003 a_1179_183# a_1001_47# VGND VNB nshort w=640000u l=150000u
+  ad=1.978e+11p pd=1.99e+06u as=0p ps=0u
M1004 VPWR SCD a_698_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=2.144e+11p ps=1.95e+06u
M1005 a_1464_413# a_27_47# a_1179_183# VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=2.307e+11p ps=2.19e+06u
M1006 a_1001_47# a_27_47# a_604_369# VNB nshort w=360000u l=150000u
+  ad=1.548e+11p pd=1.58e+06u as=2.604e+11p ps=2.88e+06u
M1007 VPWR CLK a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1008 VPWR a_1653_315# a_2114_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1009 a_698_369# a_319_47# a_604_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=2.99e+11p ps=3.24e+06u
M1010 a_604_369# D a_529_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1011 VGND a_1653_315# a_2114_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1012 VPWR a_1464_413# a_1653_315# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1013 a_503_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=2.08e+11p pd=1.93e+06u as=0p ps=0u
M1014 VGND a_1179_183# a_1117_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.374e+11p ps=1.52e+06u
M1015 a_717_47# SCE a_604_369# VNB nshort w=420000u l=150000u
+  ad=9.66e+10p pd=1.3e+06u as=0p ps=0u
M1016 a_604_369# D a_503_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND SCE a_319_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1018 VPWR SCE a_319_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1019 a_1111_413# a_27_47# a_1001_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.407e+11p ps=1.51e+06u
M1020 VGND a_1653_315# a_1615_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.446e+11p ps=1.55e+06u
M1021 a_1179_183# a_1001_47# VPWR VPB phighvt w=750000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1001_47# a_211_363# a_604_369# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1024 a_1464_413# a_211_363# a_1179_183# VNB nshort w=360000u l=150000u
+  ad=1.854e+11p pd=1.75e+06u as=0p ps=0u
M1025 a_529_47# a_319_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_1653_315# a_1558_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=2.037e+11p ps=1.81e+06u
M1027 Q_N a_2114_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1028 a_211_363# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1029 a_1117_47# a_211_363# a_1001_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Q_N a_2114_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1031 a_1558_413# a_211_363# a_1464_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Q a_1653_315# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1033 VGND SCD a_717_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1615_47# a_27_47# a_1464_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND a_1464_413# a_1653_315# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
.ends
.subckt sky130_fd_sc_hdll__nor2b_1 B_N Y A VPB VNB VGND VPWR
M1000 a_253_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.3e+11p pd=2.46e+06u as=3.666e+11p ps=3e+06u
M1001 VPWR B_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1002 VGND a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=4.912e+11p pd=4.26e+06u as=1.755e+11p ps=1.84e+06u
M1003 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y a_27_47# a_253_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1005 VGND B_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
.ends
.subckt sky130_fd_sc_hdll__a21boi_4 Y A1 B1_N A2 VNB VPB VGND VPWR
M1000 a_724_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=7.8e+11p pd=7.6e+06u as=1.365e+12p ps=1.07e+07u
M1001 a_724_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=8.905e+11p ps=7.94e+06u
M1003 VPWR A2 a_227_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.465e+12p pd=1.293e+07u as=2.125e+12p ps=1.825e+07u
M1004 VGND A2 a_724_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_227_297# a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=6e+11p ps=5.2e+06u
M1006 a_227_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A1 a_724_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_227_297# a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_724_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B1_N a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.75e+11p ps=2.55e+06u
M1011 VPWR A2 a_227_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A2 a_724_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_724_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A1 a_227_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND B1_N a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.0225e+11p ps=2.23e+06u
M1016 Y a_27_47# a_227_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A1 a_227_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y A1 a_724_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_227_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y a_27_47# a_227_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_227_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_227_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand3_4 Y A B C VNB VPB VGND VPWR
M1000 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=2.25e+12p pd=2.05e+07u as=1.74e+12p ps=1.548e+07u
M1001 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_27_47# C VGND VNB nshort w=650000u l=150000u
+  ad=9.62e+11p pd=9.46e+06u as=4.16e+11p ps=3.88e+06u
M1003 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_485_47# A Y VNB nshort w=650000u l=150000u
+  ad=1.0335e+12p pd=9.68e+06u as=4.16e+11p ps=3.88e+06u
M1005 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_47# B a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_485_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_485_47# B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND C a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_47# C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_47# B a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_485_47# B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND C a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__mux2_4 X S A0 A1 VNB VPB VPWR VGND
M1000 VPWR a_424_297# X VPB phighvt w=1e+06u l=180000u
+  ad=1.195e+12p pd=1.039e+07u as=5.8e+11p ps=5.16e+06u
M1001 a_424_297# A0 a_334_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.4e+11p pd=2.68e+06u as=5.4e+11p ps=5.08e+06u
M1002 X a_424_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_424_297# VGND VNB nshort w=650000u l=150000u
+  ad=4.16e+11p pd=3.88e+06u as=8.3525e+11p ps=7.77e+06u
M1004 VPWR S a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1005 VGND a_424_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_530_47# A1 a_424_297# VNB nshort w=650000u l=150000u
+  ad=5.8175e+11p pd=3.09e+06u as=2.405e+11p ps=2.04e+06u
M1007 VPWR a_424_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND S a_530_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_424_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND S a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1011 a_424_297# A0 a_226_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=5.525e+11p ps=3e+06u
M1012 VPWR S a_334_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_424_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_222_297# A1 a_424_297# VPB phighvt w=1e+06u l=180000u
+  ad=6e+11p pd=5.2e+06u as=0p ps=0u
M1015 a_226_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_222_297# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_424_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and2b_4 B X A_N VNB VPB VGND VPWR
M1000 VPWR B a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=1.2757e+12p pd=1.065e+07u as=2.9e+11p ps=2.58e+06u
M1001 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=6.1e+11p ps=5.22e+06u
M1002 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=7.61e+11p pd=6.33e+06u as=4.615e+11p ps=4.02e+06u
M1003 VGND B a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.365e+11p ps=1.72e+06u
M1004 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_47# a_33_199# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_33_199# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1007 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_119_47# a_33_199# a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1009 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_33_199# A_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.344e+11p pd=1.48e+06u as=0p ps=0u
M1011 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o22a_2 A2 X B1 A1 B2 VNB VPB VGND VPWR
M1000 a_321_47# B2 a_83_21# VNB nshort w=650000u l=150000u
+  ad=7.02e+11p pd=6.06e+06u as=1.755e+11p ps=1.84e+06u
M1001 X a_83_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=1.38e+12p ps=8.76e+06u
M1002 a_627_297# A2 a_83_21# VPB phighvt w=1e+06u l=180000u
+  ad=2.3e+11p pd=2.46e+06u as=4.9e+11p ps=2.98e+06u
M1003 VPWR A1 a_627_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_321_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=5.655e+11p ps=5.64e+06u
M1005 a_411_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.3e+11p pd=2.46e+06u as=0p ps=0u
M1006 X a_83_21# VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=0p ps=0u
M1007 a_83_21# B2 a_411_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2 a_321_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_83_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_83_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_83_21# B1 a_321_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a221oi_2 B2 C1 A2 A1 B1 Y VNB VPB VGND VPWR
M1000 Y B1 a_413_47# VNB nshort w=650000u l=150000u
+  ad=6.89e+11p pd=6.02e+06u as=3.835e+11p ps=3.78e+06u
M1001 a_27_297# B1 a_321_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.13e+12p pd=1.026e+07u as=1.515e+12p ps=1.303e+07u
M1002 VPWR A2 a_321_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1003 a_805_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=3.835e+11p pd=3.78e+06u as=1.183e+12p ps=8.84e+06u
M1004 Y C1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=0p ps=0u
M1005 a_321_297# B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A1 a_805_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND C1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_297# B2 a_321_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_321_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B2 a_413_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_413_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A2 a_805_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A1 a_321_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_805_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_321_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y C1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_413_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_297# C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_321_297# B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sdfrtp_4 VPB VNB RESET_B VPWR VGND SCE SCD D CLK Q
M1000 a_1428_47# a_1380_303# a_1322_47# VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.518e+11p ps=1.6e+06u
M1001 Q a_1972_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6.45e+11p pd=5.29e+06u as=2.2648e+12p ps=2.094e+07u
M1002 a_213_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=1.7043e+12p ps=1.636e+07u
M1003 VPWR a_1972_21# a_1951_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
M1004 a_1972_21# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=1.344e+11p pd=1.48e+06u as=0p ps=0u
M1005 Q a_1972_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_2157_47# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=0p ps=0u
M1007 VPWR SCD a_870_389# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=1.971e+11p ps=1.81e+06u
M1008 a_700_389# D a_631_119# VNB nshort w=420000u l=150000u
+  ad=3.3215e+11p pd=3.47e+06u as=1.302e+11p ps=1.46e+06u
M1009 a_1380_303# a_1202_413# VPWR VPB phighvt w=840000u l=180000u
+  ad=2.541e+11p pd=2.37e+06u as=0p ps=0u
M1010 a_1202_413# a_27_47# a_700_389# VNB nshort w=360000u l=150000u
+  ad=1.44e+11p pd=1.52e+06u as=0p ps=0u
M1011 VPWR a_1757_47# a_1972_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1972_21# a_1757_47# a_2157_47# VNB nshort w=420000u l=150000u
+  ad=1.365e+11p pd=1.49e+06u as=0p ps=0u
M1013 VGND a_1972_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=5.265e+11p ps=4.22e+06u
M1014 VGND a_1972_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_1380_303# a_1324_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1016 VPWR CLK a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1017 a_618_389# SCE VPWR VPB phighvt w=540000u l=180000u
+  ad=1.242e+11p pd=1.54e+06u as=0p ps=0u
M1018 a_1951_413# a_213_47# a_1757_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1019 Q a_1972_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_700_389# D a_618_389# VPB phighvt w=540000u l=180000u
+  ad=5.193e+11p pd=4.01e+06u as=0p ps=0u
M1021 a_631_119# a_331_66# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND RESET_B a_1428_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1324_413# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_1972_21# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1202_413# a_213_47# a_700_389# VPB phighvt w=420000u l=180000u
+  ad=1.806e+11p pd=1.7e+06u as=0p ps=0u
M1026 a_1324_413# a_27_47# a_1202_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1866_47# a_27_47# a_1757_47# VNB nshort w=360000u l=150000u
+  ad=2.121e+11p pd=1.9e+06u as=1.422e+11p ps=1.51e+06u
M1028 a_1757_47# a_213_47# a_1380_303# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.87e+11p ps=1.93e+06u
M1029 Q a_1972_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR SCE a_331_66# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=2.214e+11p ps=1.9e+06u
M1031 VGND CLK a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1032 VGND a_1972_21# a_1866_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_213_47# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
M1034 a_899_66# SCE a_700_389# VNB nshort w=420000u l=500000u
+  ad=1.554e+11p pd=1.58e+06u as=0p ps=0u
M1035 a_1757_47# a_27_47# a_1380_303# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1322_47# a_213_47# a_1202_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR a_1972_21# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND SCD a_899_66# VNB nshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_870_389# a_331_66# a_700_389# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND SCE a_331_66# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1041 a_1380_303# a_1202_413# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and4b_1 VGND VPWR C A_N X D B VPB VNB
M1000 a_379_47# B a_307_47# VNB nshort w=420000u l=150000u
+  ad=2.1e+11p pd=1.84e+06u as=8.82e+10p ps=1.26e+06u
M1001 VPWR A_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=7.115e+11p pd=6.35e+06u as=1.134e+11p ps=1.38e+06u
M1002 a_509_47# C a_379_47# VNB nshort w=420000u l=150000u
+  ad=1.491e+11p pd=1.55e+06u as=0p ps=0u
M1003 X a_213_413# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=3.422e+11p ps=3.43e+06u
M1004 VPWR B a_213_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=3.171e+11p ps=3.19e+06u
M1005 VGND D a_509_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_213_413# a_27_47# VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_213_413# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1008 VGND A_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1009 a_213_413# C VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR D a_213_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_307_47# a_27_47# a_213_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
.ends
.subckt sky130_fd_sc_hdll__probe_p_8 X A VGND VPWR VPB VNB
M1000 a_399_297# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=1.72e+12p ps=1.544e+07u
M1001 a_27_47# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
M1002 a_27_47# A VGND VNB nshort w=650000u l=150000u
+  ad=3.77e+11p pd=3.76e+06u as=1.339e+12p ps=1.192e+07u
M1003 VPWR a_27_47# a_399_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_27_47# a_399_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.02e+11p ps=7.36e+06u
M1005 VPWR a_27_47# a_399_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_399_297# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_399_297# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_27_47# a_399_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_27_47# a_399_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_399_297# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_399_297# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_399_297# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_399_297# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
R0 a_399_297# X short w=3.02e+06u l=5000u
M1017 VPWR a_27_47# a_399_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_27_47# a_399_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_399_297# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_27_47# a_399_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o32ai_4 A1 A2 A3 B1 Y B2 VNB VPB VGND VPWR
M1000 a_27_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.425e+12p pd=1.285e+07u as=1.41e+12p ps=1.282e+07u
M1001 a_1352_297# A2 a_886_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.205e+12p pd=1.041e+07u as=1.41e+12p ps=1.282e+07u
M1002 a_27_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.16e+12p ps=1.032e+07u
M1003 a_1352_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=2.75925e+12p pd=2.279e+07u as=8.645e+11p ps=7.86e+06u
M1005 a_27_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.41375e+12p ps=1.215e+07u
M1007 VPWR B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_886_297# A2 a_1352_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A1 a_1352_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A3 a_886_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A3 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1352_297# A2 a_886_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_886_297# A2 a_1352_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_886_297# A3 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1352_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_27_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_27_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_27_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y A3 a_886_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A1 a_1352_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND A3 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_27_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND A2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Y B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_886_297# A3 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 Y B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor3_2 C Y A B VPB VNB VGND VPWR
M1000 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u
M1001 VGND C Y VNB nshort w=650000u l=150000u
+  ad=8.6125e+11p pd=9.15e+06u as=7.215e+11p ps=6.12e+06u
M1002 a_27_297# B a_309_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.3e+11p ps=7.66e+06u
M1003 a_309_297# C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1004 a_309_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y C a_309_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__xor2_4 X B A VNB VPB VGND VPWR
M1000 a_27_297# B a_112_47# VPB phighvt w=1e+06u l=180000u
+  ad=1.425e+12p pd=1.285e+07u as=5.8e+11p ps=5.16e+06u
M1001 VPWR A a_886_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.74e+12p pd=1.548e+07u as=1.9868e+12p ps=1.798e+07u
M1002 X B a_886_47# VNB nshort w=650000u l=150000u
+  ad=8.97e+11p pd=7.96e+06u as=9.295e+11p ps=9.36e+06u
M1003 a_112_47# A VGND VNB nshort w=650000u l=150000u
+  ad=8.645e+11p pd=7.86e+06u as=1.97925e+12p ps=1.909e+07u
M1004 a_886_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_112_47# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_886_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A a_886_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR B a_886_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_112_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B a_112_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A a_886_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A a_112_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_886_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_886_297# a_112_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.6245e+11p ps=7.74e+06u
M1017 X B a_886_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_886_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_112_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_886_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_886_47# B X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_297# B a_112_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X a_112_47# a_886_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_112_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND B a_112_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR B a_886_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 X a_112_47# a_886_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_112_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND A a_112_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND A a_886_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_112_47# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_886_297# a_112_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_886_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 X a_112_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_886_47# B X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND a_112_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_112_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or3b_4 A B C_N X VNB VPB VGND VPWR
M1000 VPWR a_186_21# X VPB phighvt w=1e+06u l=180000u
+  ad=8.857e+11p pd=7.87e+06u as=5.8e+11p ps=5.16e+06u
M1001 X a_186_21# VGND VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=8.635e+11p ps=7.91e+06u
M1002 a_186_21# A VGND VNB nshort w=650000u l=150000u
+  ad=3.77e+11p pd=3.76e+06u as=0p ps=0u
M1003 a_186_21# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_186_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_186_21# a_27_47# a_694_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=3.5e+11p ps=2.7e+06u
M1006 VGND B a_186_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_186_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_186_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR C_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1010 VGND C_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1011 X a_186_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_186_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_186_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_694_297# B a_600_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1015 a_600_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o21ba_4 B1_N A1 A2 X VNB VPB VGND VPWR
M1000 VPWR a_197_21# X VPB phighvt w=1e+06u l=180000u
+  ad=1.43e+12p pd=1.286e+07u as=5.8e+11p ps=5.16e+06u
M1001 a_823_297# A2 a_197_21# VPB phighvt w=1e+06u l=180000u
+  ad=8.5e+11p pd=7.7e+06u as=5.8e+11p ps=5.16e+06u
M1002 VGND A2 a_635_47# VNB nshort w=650000u l=150000u
+  ad=1.0335e+12p pd=9.68e+06u as=7.345e+11p ps=7.46e+06u
M1003 a_635_47# a_27_297# a_197_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1004 VPWR B1_N a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.9e+11p ps=2.78e+06u
M1005 a_635_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_197_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_197_21# VGND VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=0p ps=0u
M1008 a_197_21# A2 a_823_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_197_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_197_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_197_21# a_27_297# a_635_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A1 a_635_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_197_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_197_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_823_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_27_297# a_197_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND B1_N a_27_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.3075e+11p ps=2.01e+06u
M1018 VPWR A1 a_823_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_635_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_197_21# a_27_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_197_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a31o_1 A2 B1 A1 A3 X VPB VNB VGND VPWR
M1000 VGND B1 a_80_21# VNB nshort w=650000u l=150000u
+  ad=4.9075e+11p pd=4.11e+06u as=2.47e+11p ps=2.06e+06u
M1001 VPWR A2 a_225_297# VPB phighvt w=1e+06u l=180000u
+  ad=7.05e+11p pd=5.41e+06u as=7e+11p ps=5.4e+06u
M1002 a_225_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR a_80_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.75e+11p ps=2.55e+06u
M1004 VGND a_80_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u
M1005 a_225_297# A3 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_323_47# A2 a_217_47# VNB nshort w=650000u l=150000u
+  ad=2.47e+11p pd=2.06e+06u as=2.47e+11p ps=2.06e+06u
M1007 a_80_21# A1 a_323_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_217_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_80_21# B1 a_225_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.3e+11p pd=2.66e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__xnor3_1 X B C A VNB VPB VGND VPWR
M1000 VPWR a_83_21# X VPB phighvt w=1e+06u l=180000u
+  ad=1.22595e+12p pd=8.52e+06u as=2.9e+11p ps=2.58e+06u
M1001 a_901_297# a_783_297# a_375_49# VNB nshort w=600000u l=150000u
+  ad=4.4975e+11p pd=3.99e+06u as=5.4545e+11p ps=4.31e+06u
M1002 a_83_21# C a_375_49# VNB nshort w=640000u l=150000u
+  ad=2.176e+11p pd=1.96e+06u as=0p ps=0u
M1003 a_1184_297# a_901_297# VGND VNB nshort w=640000u l=150000u
+  ad=5.677e+11p pd=4.42e+06u as=9.124e+11p ps=6.76e+06u
M1004 a_783_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.2e+11p pd=2.64e+06u as=0p ps=0u
M1005 a_901_297# a_783_297# a_351_325# VPB phighvt w=840000u l=180000u
+  ad=7.226e+11p pd=5.29e+06u as=5.878e+11p ps=4.8e+06u
M1006 a_351_325# B a_901_297# VNB nshort w=640000u l=150000u
+  ad=6.091e+11p pd=4.57e+06u as=0p ps=0u
M1007 a_1184_297# a_901_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=7.998e+11p pd=5.68e+06u as=0p ps=0u
M1008 a_783_297# B VGND VNB nshort w=650000u l=150000u
+  ad=1.6515e+11p pd=1.82e+06u as=0p ps=0u
M1009 VGND A a_901_297# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_375_49# B a_901_297# VPB phighvt w=840000u l=180000u
+  ad=8.3175e+11p pd=5.4e+06u as=0p ps=0u
M1011 a_351_325# B a_1184_297# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_83_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.82e+11p ps=1.86e+06u
M1013 a_351_325# a_226_93# a_83_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A a_901_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_83_21# C a_351_325# VPB phighvt w=840000u l=180000u
+  ad=3.227e+11p pd=2.67e+06u as=0p ps=0u
M1016 a_1184_297# a_783_297# a_351_325# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_226_93# C VPWR VPB phighvt w=640000u l=180000u
+  ad=1.856e+11p pd=1.86e+06u as=0p ps=0u
M1018 a_1184_297# a_783_297# a_375_49# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_375_49# B a_1184_297# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_226_93# C VGND VNB nshort w=420000u l=150000u
+  ad=1.995e+11p pd=1.79e+06u as=0p ps=0u
M1021 a_375_49# a_226_93# a_83_21# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or4bb_4 D_N B A C_N X VNB VPB VGND VPWR
M1000 X a_335_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=1.20363e+12p ps=1.058e+07u
M1001 a_425_297# a_224_297# a_335_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.5e+11p pd=2.7e+06u as=2.7e+11p ps=2.54e+06u
M1002 VGND A a_335_297# VNB nshort w=650000u l=150000u
+  ad=1.2044e+12p pd=1.129e+07u as=4.355e+11p ps=3.94e+06u
M1003 VPWR A a_625_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1004 a_224_297# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1005 a_335_297# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_335_297# VGND VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=0p ps=0u
M1007 VPWR a_335_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND C_N a_27_410# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1009 a_625_297# B a_531_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1010 a_531_297# a_27_410# a_425_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_335_297# a_224_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_27_410# a_335_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_335_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR C_N a_27_410# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1015 X a_335_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_335_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_224_297# D_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1018 VPWR a_335_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_335_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__probec_p_8 X A VGND VPWR VPB VNB
M1000 a_399_297# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=1.72e+12p ps=1.544e+07u
M1001 a_27_47# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
M1002 a_27_47# A VGND VNB nshort w=650000u l=150000u
+  ad=3.77e+11p pd=3.76e+06u as=1.339e+12p ps=1.192e+07u
M1003 VPWR a_27_47# a_399_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
R0 X a_399_297# short w=1.6e+06u l=100000u
M1004 VGND a_27_47# a_399_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.02e+11p ps=7.36e+06u
M1005 VPWR a_27_47# a_399_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_399_297# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_399_297# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_27_47# a_399_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_27_47# a_399_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_399_297# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_399_297# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_399_297# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_399_297# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
R1 VPWR m5_872_595# short w=0u l=1.2e+06u
R2 VGND m5_872_n71# short w=0u l=1.2e+06u
M1017 VPWR a_27_47# a_399_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_27_47# a_399_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_399_297# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_27_47# a_399_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor3b_4 A C_N B Y VPB VNB VGND VPWR
M1000 VPWR A a_215_297# VPB phighvt w=1e+06u l=180000u
+  ad=8.5e+11p pd=7.7e+06u as=1.16e+12p ps=1.032e+07u
M1001 VPWR C_N a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1002 Y A VGND VNB nshort w=650000u l=150000u
+  ad=1.3455e+12p pd=1.194e+07u as=1.6575e+12p ps=1.42e+07u
M1003 a_605_297# B a_215_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.41e+12p pd=1.282e+07u as=0p ps=0u
M1004 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C_N a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.145e+11p ps=1.96e+06u
M1007 Y a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_215_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_605_297# a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1010 a_215_297# B a_605_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A a_215_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y a_27_47# a_605_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_605_297# B a_215_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_215_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_605_297# a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_215_297# B a_605_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y a_27_47# a_605_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o221ai_4 B1 B2 A2 C1 Y A1 VNB VPB VGND VPWR
M1000 Y C1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.74e+12p pd=1.548e+07u as=2.645e+12p ps=1.929e+07u
M1001 a_601_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=0p ps=0u
M1002 Y A2 a_1369_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.16e+12p ps=1.032e+07u
M1003 a_1369_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_511_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=1.976e+12p pd=1.778e+07u as=7.67e+11p ps=7.56e+06u
M1005 a_1369_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y C1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=4.16e+11p pd=3.88e+06u as=1.391e+12p ps=1.338e+07u
M1007 a_511_47# B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A1 a_511_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y B2 a_601_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_511_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y C1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR B1 a_601_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A1 a_511_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A2 a_1369_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_47# C1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A2 a_511_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_601_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_511_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y C1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_27_47# B1 a_511_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1369_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_511_47# B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_601_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR A1 a_1369_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_27_47# B2 a_511_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR B1 a_601_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_511_47# B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y B2 a_601_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_27_47# C1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_511_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_511_47# B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_601_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR A1 a_1369_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND A2 a_511_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_27_47# B1 a_511_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1369_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_27_47# B2 a_511_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or2_6 X A B VNB VPB VGND VPWR
M1000 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.42e+12p pd=1.284e+07u as=8.5e+11p ps=7.7e+06u
M1001 VGND A a_123_47# VNB nshort w=650000u l=150000u
+  ad=1.7225e+12p pd=1.31e+07u as=3.51e+11p ps=3.68e+06u
M1002 X a_123_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.7e+11p pd=7.74e+06u as=0p ps=0u
M1003 VGND a_123_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=5.265e+11p ps=5.52e+06u
M1004 a_123_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_123_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_297# B a_123_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1007 VPWR a_123_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_123_47# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_123_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_123_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_123_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_123_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND B a_123_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_123_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_123_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_123_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_123_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_123_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o31ai_4 A3 A2 A1 Y B1 VGND VPWR VPB VNB
M1000 VGND A3 a_31_47# VNB nshort w=650000u l=150000u
+  ad=1.72575e+12p pd=1.311e+07u as=1.729e+12p ps=1.702e+07u
M1001 a_497_297# A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=1.45e+12p ps=1.29e+07u
M1002 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=0p ps=0u
M1003 a_31_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_31_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1005 Y A3 a_497_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.435e+12p pd=1.287e+07u as=0p ps=0u
M1006 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_497_297# A3 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2 a_31_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 a_31_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_31_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_31_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A1 a_31_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_31_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_297# A2 a_497_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_31_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y A3 a_497_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A2 a_31_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y B1 a_31_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A3 a_31_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_497_297# A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND A1 a_31_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_31_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_497_297# A3 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_31_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_27_297# A2 a_497_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and3_2 B X A C VPWR VGND VPB VNB
M1000 VGND a_29_311# X VNB nshort w=650000u l=150000u
+  ad=5.093e+11p pd=4.31e+06u as=2.21e+11p ps=1.98e+06u
M1001 VGND C a_194_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.281e+11p ps=1.45e+06u
M1002 VPWR C a_29_311# VPB phighvt w=420000u l=180000u
+  ad=8.325e+11p pd=6.94e+06u as=2.7055e+11p ps=3.05e+06u
M1003 a_29_311# B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_194_53# B a_122_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1005 VPWR a_29_311# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1006 X a_29_311# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_29_311# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_122_53# A a_29_311# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1009 VPWR A a_29_311# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__clkbuf_2 VPB VGND VPWR VNB A X
M1000 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=2.457e+11p pd=2.85e+06u as=1.323e+11p ps=1.47e+06u
M1001 VGND a_27_47# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.554e+11p ps=1.58e+06u
M1002 VPWR A a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=6.15e+11p pd=5.23e+06u as=2.75e+11p ps=2.55e+06u
M1003 X a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1005 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__clkinv_2 Y A VNB VPB VPWR VGND
M1000 VGND A Y VNB nshort w=420000u l=150000u
+  ad=2.415e+11p pd=2.83e+06u as=1.386e+11p ps=1.5e+06u
M1001 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=5.75e+11p ps=5.15e+06u
M1002 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sdfstp_2 Q SCD D CLK SET_B SCE VGND VPWR VPB VNB
M1000 VPWR SET_B a_1229_21# VPB phighvt w=420000u l=180000u
+  ad=2.0718e+12p pd=1.868e+07u as=1.722e+11p ps=1.66e+06u
M1001 VGND a_349_21# a_295_47# VNB nshort w=420000u l=150000u
+  ad=1.50395e+12p pd=1.505e+07u as=1.134e+11p ps=1.38e+06u
M1002 a_2067_47# a_1951_295# a_1995_47# VNB nshort w=420000u l=150000u
+  ad=2.016e+11p pd=1.8e+06u as=8.82e+10p ps=1.26e+06u
M1003 a_1745_329# SET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=4.746e+11p pd=4.26e+06u as=0p ps=0u
M1004 a_1951_295# a_1745_329# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1005 a_1995_47# a_693_369# a_1745_329# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.332e+11p ps=2.5e+06u
M1006 a_1891_413# a_877_369# a_1745_329# VPB phighvt w=420000u l=180000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1007 VGND SCE a_349_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1008 a_1075_413# a_877_369# a_201_47# VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=2.99e+11p ps=3.24e+06u
M1009 VPWR SCD a_27_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=3.456e+11p ps=3.64e+06u
M1010 a_1229_21# a_1075_413# VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR SCE a_349_21# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1012 VGND SET_B a_2067_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_2447_47# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1014 VGND SET_B a_1467_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1015 a_877_369# a_693_369# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1016 VGND a_1229_21# a_1177_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1017 VPWR a_1951_295# a_1891_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND CLK a_693_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1019 a_1951_295# a_1745_329# VGND VNB nshort w=420000u l=150000u
+  ad=1.596e+11p pd=1.6e+06u as=0p ps=0u
M1020 a_1654_47# a_1075_413# VGND VNB nshort w=640000u l=150000u
+  ad=5.088e+11p pd=2.87e+06u as=0p ps=0u
M1021 a_1467_47# a_1075_413# a_1229_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.512e+11p ps=1.56e+06u
M1022 Q a_2447_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_369# a_349_21# a_201_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_119_47# SCD VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1025 a_1177_47# a_877_369# a_1075_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1026 VGND a_1745_329# a_2447_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1027 a_877_369# a_693_369# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1028 a_1663_329# a_1075_413# VPWR VPB phighvt w=840000u l=180000u
+  ad=1.932e+11p pd=2.14e+06u as=0p ps=0u
M1029 VPWR a_1745_329# a_2447_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1030 a_1075_413# a_693_369# a_201_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.646e+11p ps=2.94e+06u
M1031 a_1745_329# a_693_369# a_1663_329# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_295_47# D a_201_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND a_2447_47# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1034 a_201_47# SCE a_119_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 Q a_2447_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_211_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=1.472e+11p pd=1.74e+06u as=0p ps=0u
M1037 a_201_47# D a_211_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1169_413# a_693_369# a_1075_413# VPB phighvt w=420000u l=180000u
+  ad=1.596e+11p pd=1.6e+06u as=0p ps=0u
M1039 VPWR a_1229_21# a_1169_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VPWR CLK a_693_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1041 a_1745_329# a_877_369# a_1654_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a211o_1 VNB VPB VGND VPWR X A2 B1 A1 C1
M1000 a_80_21# C1 a_546_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.75e+11p pd=2.55e+06u as=3.5e+11p ps=2.7e+06u
M1001 VGND B1 a_80_21# VNB nshort w=650000u l=150000u
+  ad=8.32e+11p pd=5.16e+06u as=3.8675e+11p ps=3.79e+06u
M1002 VPWR a_80_21# X VPB phighvt w=1e+06u l=180000u
+  ad=7.55e+11p pd=5.51e+06u as=2.75e+11p ps=2.55e+06u
M1003 VGND a_80_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u
M1004 a_546_297# B1 a_227_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.75e+11p ps=5.15e+06u
M1005 VPWR A2 a_227_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_80_21# A1 a_320_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.315e+11p ps=2.32e+06u
M1007 a_320_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_227_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_80_21# C1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor2_8 Y A B VPB VNB VGND VPWR
M1000 Y B VGND VNB nshort w=650000u l=150000u
+  ad=1.729e+12p pd=1.572e+07u as=1.7745e+12p ps=1.716e+07u
M1001 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=2.6e+12p ps=2.32e+07u
M1002 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=0p ps=0u
M1004 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_297# B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_297# B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_297# B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_297# B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a21o_1 A2 A1 B1 X VPWR VGND VPB VNB
M1000 VGND a_81_21# X VNB nshort w=650000u l=150000u
+  ad=7.8325e+11p pd=5.01e+06u as=1.69e+11p ps=1.82e+06u
M1001 a_81_21# B1 VGND VNB nshort w=650000u l=150000u
+  ad=2.1775e+11p pd=1.97e+06u as=0p ps=0u
M1002 VPWR A1 a_317_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.7e+11p pd=5.14e+06u as=5.8e+11p ps=5.16e+06u
M1003 VPWR a_81_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1004 VGND A2 a_416_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.82e+11p ps=1.86e+06u
M1005 a_317_297# B1 a_81_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1006 a_317_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_416_47# A1 a_81_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__einvn_4 TE_B Z A VGND VPWR VPB VNB
M1000 VPWR TE_B a_222_309# VPB phighvt w=940000u l=180000u
+  ad=8.663e+11p pd=7.57e+06u as=1.3752e+12p ps=1.258e+07u
M1001 a_235_47# A Z VNB nshort w=650000u l=150000u
+  ad=1.04325e+12p pd=9.71e+06u as=4.16e+11p ps=3.88e+06u
M1002 Z A a_235_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_222_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_235_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=6.175e+11p ps=5.8e+06u
M1005 VGND a_27_47# a_235_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR TE_B a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1007 a_222_309# A Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1008 a_235_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_235_47# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Z A a_235_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Z A a_222_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_222_309# A Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_27_47# a_235_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR TE_B a_222_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_222_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND TE_B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1017 Z A a_222_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand2_16 Y A B VPB VNB VGND VPWR
M1000 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=4.89e+12p pd=4.378e+07u as=4.64e+12p ps=4.128e+07u
M1001 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=1.859e+12p pd=1.612e+07u as=3.0355e+12p ps=3.144e+07u
M1002 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.924e+12p ps=1.632e+07u
M1005 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1049 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1050 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1051 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1052 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1053 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1054 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1055 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1056 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1057 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1058 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1059 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1060 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1061 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1062 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1063 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__buf_16 A X VNB VPB VGND VPWR
M1000 VPWR a_109_47# X VPB phighvt w=1e+06u l=180000u
+  ad=3.44e+12p pd=3.088e+07u as=2.32e+12p ps=2.064e+07u
M1001 VPWR A a_109_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.7e+11p ps=7.74e+06u
M1002 VPWR a_109_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_109_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_109_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_109_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.6965e+12p pd=1.562e+07u as=2.3855e+12p ps=2.294e+07u
M1006 VGND a_109_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_109_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_109_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_109_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_109_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_109_47# A VGND VNB nshort w=650000u l=150000u
+  ad=6.565e+11p pd=5.92e+06u as=0p ps=0u
M1012 X a_109_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A a_109_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_109_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_109_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_109_47# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_109_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_109_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_109_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_109_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_109_47# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_109_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X a_109_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 X a_109_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_109_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR a_109_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND A a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND a_109_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A a_109_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR a_109_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 X a_109_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 X a_109_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND a_109_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR a_109_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_109_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_109_47# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_109_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND A a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 X a_109_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 X a_109_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 X a_109_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 X a_109_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a21boi_2 VNB VPB VPWR VGND B1_N A2 A1 Y
M1000 a_228_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.2e+12p pd=1.04e+07u as=7.055e+11p ps=6.57e+06u
M1001 VPWR A2 a_228_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_228_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_228_297# a_61_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1004 Y A1 a_529_47# VNB nshort w=650000u l=150000u
+  ad=4.225e+11p pd=3.9e+06u as=1.365e+11p ps=1.72e+06u
M1005 Y a_61_47# a_228_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_61_47# Y VNB nshort w=650000u l=150000u
+  ad=8.845e+11p pd=6.71e+06u as=0p ps=0u
M1007 a_61_47# B1_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.155e+11p pd=1.39e+06u as=0p ps=0u
M1008 VPWR A1 a_228_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_529_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B1_N a_61_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1011 a_697_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=0p ps=0u
M1012 Y a_61_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A2 a_697_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand3_2 A Y B C VNB VPB VGND VPWR
M1000 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=1.42e+12p pd=1.284e+07u as=8.7e+11p ps=7.74e+06u
M1001 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=5.785e+11p pd=5.68e+06u as=2.08e+11p ps=1.94e+06u
M1002 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND C a_307_47# VNB nshort w=650000u l=150000u
+  ad=4.03e+11p pd=3.84e+06u as=4.16e+11p ps=3.88e+06u
M1005 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_307_47# C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_47# B a_307_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_307_47# B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__einvp_1 TE A Z VPWR VGND VPB VNB
M1000 a_332_297# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=4.55e+11p pd=2.91e+06u as=8.457e+11p ps=3.79e+06u
M1001 VPWR TE a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1002 Z A a_204_47# VNB nshort w=650000u l=150000u
+  ad=2.08e+11p pd=1.94e+06u as=7.0525e+11p ps=3.47e+06u
M1003 VGND TE a_27_47# VNB nshort w=420000u l=150000u
+  ad=1.94e+11p pd=1.95e+06u as=1.092e+11p ps=1.36e+06u
M1004 Z A a_332_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1005 a_204_47# TE VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a32o_4 A3 X B1 B2 A1 A2 VNB VPB VGND VPWR
M1000 a_79_21# B1 a_493_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=2.36e+12p ps=1.672e+07u
M1001 a_485_47# A2 a_695_47# VNB nshort w=650000u l=150000u
+  ad=4.16e+11p pd=3.88e+06u as=5.785e+11p ps=5.68e+06u
M1002 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=1.7e+12p pd=1.54e+07u as=5.8e+11p ps=5.16e+06u
M1003 a_493_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=9.62e+11p ps=9.46e+06u
M1005 VPWR A3 a_493_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_1194_47# B1 a_79_21# VNB nshort w=650000u l=150000u
+  ad=6.0775e+11p pd=5.77e+06u as=4.16e+11p ps=3.88e+06u
M1008 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_493_297# B2 a_79_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_493_297# A3 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1194_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A1 a_493_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_79_21# B2 a_493_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND B2 a_1194_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_695_47# A1 a_79_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_79_21# B1 a_1194_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_493_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_695_47# A2 a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_493_297# B1 a_79_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A3 a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_485_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_79_21# A1 a_695_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR A2 a_493_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__mux2_2 VGND VPWR A1 A0 S X VPB VNB
M1000 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=7.764e+11p pd=7.11e+06u as=2.9e+11p ps=2.58e+06u
M1001 a_280_21# S VPWR VPB phighvt w=640000u l=180000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1002 a_606_369# A0 a_79_21# VPB phighvt w=640000u l=180000u
+  ad=1.472e+11p pd=1.74e+06u as=1.92e+11p ps=1.88e+06u
M1003 VPWR S a_606_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_79_21# A0 a_310_47# VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=1.386e+11p ps=1.5e+06u
M1005 VGND S a_502_47# VNB nshort w=420000u l=150000u
+  ad=5.551e+11p pd=5.47e+06u as=3.108e+11p ps=2.32e+06u
M1006 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1007 a_502_47# A1 a_79_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_318_369# a_280_21# VPWR VPB phighvt w=640000u l=180000u
+  ad=4.992e+11p pd=2.84e+06u as=0p ps=0u
M1009 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_79_21# A1 a_318_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_310_47# a_280_21# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_280_21# S VGND VNB nshort w=420000u l=150000u
+  ad=1.155e+11p pd=1.39e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and2b_2 VNB VPB VPWR VGND X B A_N
M1000 VPWR a_230_413# X VPB phighvt w=1e+06u l=180000u
+  ad=9.248e+11p pd=7.78e+06u as=4.5e+11p ps=2.9e+06u
M1001 VPWR A_N a_27_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1002 VGND B a_327_47# VNB nshort w=420000u l=150000u
+  ad=5.4195e+11p pd=5.38e+06u as=1.344e+11p ps=1.48e+06u
M1003 VPWR B a_230_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1004 VGND a_230_413# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.12e+11p ps=2.26e+06u
M1005 a_327_47# a_27_413# a_230_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1006 a_27_413# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1007 X a_230_413# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_230_413# a_27_413# VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_230_413# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sdfrtp_2 RESET_B VGND VPWR VNB VPB Q SCE SCD D CLK
M1000 a_1428_47# a_1380_303# a_1322_47# VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.518e+11p ps=1.6e+06u
M1001 a_213_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=1.6198e+12p ps=1.48e+07u
M1002 Q a_1972_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=2.0598e+12p ps=1.853e+07u
M1003 VPWR a_1972_21# a_1951_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
M1004 a_1972_21# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=1.344e+11p pd=1.48e+06u as=0p ps=0u
M1005 a_2157_47# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=0p ps=0u
M1006 VPWR SCD a_870_389# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=1.971e+11p ps=1.81e+06u
M1007 a_700_389# D a_631_119# VNB nshort w=420000u l=150000u
+  ad=3.3215e+11p pd=3.47e+06u as=1.302e+11p ps=1.46e+06u
M1008 a_1380_303# a_1202_413# VPWR VPB phighvt w=840000u l=180000u
+  ad=2.541e+11p pd=2.37e+06u as=0p ps=0u
M1009 a_1202_413# a_27_47# a_700_389# VNB nshort w=360000u l=150000u
+  ad=1.44e+11p pd=1.52e+06u as=0p ps=0u
M1010 VPWR a_1757_47# a_1972_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1972_21# a_1757_47# a_2157_47# VNB nshort w=420000u l=150000u
+  ad=1.365e+11p pd=1.49e+06u as=0p ps=0u
M1012 VPWR a_1380_303# a_1324_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1013 VPWR CLK a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1014 a_618_389# SCE VPWR VPB phighvt w=540000u l=180000u
+  ad=1.242e+11p pd=1.54e+06u as=0p ps=0u
M1015 a_1951_413# a_213_47# a_1757_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1016 VGND a_1972_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1017 a_700_389# D a_618_389# VPB phighvt w=540000u l=180000u
+  ad=5.193e+11p pd=4.01e+06u as=0p ps=0u
M1018 a_631_119# a_331_66# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Q a_1972_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND RESET_B a_1428_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1324_413# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1202_413# a_213_47# a_700_389# VPB phighvt w=420000u l=180000u
+  ad=1.806e+11p pd=1.7e+06u as=0p ps=0u
M1023 a_1324_413# a_27_47# a_1202_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1866_47# a_27_47# a_1757_47# VNB nshort w=360000u l=150000u
+  ad=2.121e+11p pd=1.9e+06u as=1.422e+11p ps=1.51e+06u
M1025 a_1757_47# a_213_47# a_1380_303# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.87e+11p ps=1.93e+06u
M1026 VPWR SCE a_331_66# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=2.214e+11p ps=1.9e+06u
M1027 VGND CLK a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1028 VGND a_1972_21# a_1866_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_213_47# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
M1030 VPWR a_1972_21# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_899_66# SCE a_700_389# VNB nshort w=420000u l=500000u
+  ad=1.554e+11p pd=1.58e+06u as=0p ps=0u
M1032 a_1757_47# a_27_47# a_1380_303# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1322_47# a_213_47# a_1202_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND SCD a_899_66# VNB nshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_870_389# a_331_66# a_700_389# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND SCE a_331_66# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1037 a_1380_303# a_1202_413# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and2_8 X B A VNB VPB VGND VPWR
M1000 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=2.01e+12p pd=1.802e+07u as=1.16e+12p ps=1.032e+07u
M1001 VGND B a_293_47# VNB nshort w=650000u l=150000u
+  ad=1.456e+12p pd=1.228e+07u as=1.82e+11p ps=1.86e+06u
M1002 VPWR A a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1003 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.02e+11p ps=7.36e+06u
M1006 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_117_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_293_47# A a_117_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1011 a_117_297# A a_131_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.56e+11p ps=1.78e+06u
M1012 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_131_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR B a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_117_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a22oi_4 A2 B2 A1 B1 Y VNB VPB VGND VPWR
M1000 a_27_297# B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=3.13e+12p pd=2.426e+07u as=1.16e+12p ps=1.032e+07u
M1001 a_883_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=9.295e+11p pd=9.36e+06u as=8.97e+11p ps=7.96e+06u
M1002 a_27_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND A2 a_883_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=0p ps=0u
M1005 a_883_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=8.645e+11p ps=7.86e+06u
M1006 Y B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=9.62e+11p ps=9.46e+06u
M1009 a_27_297# B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A1 a_883_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_883_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND A2 a_883_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_27_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_883_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_27_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y A1 a_883_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__muxb4to1_4 VPB VNB VGND VPWR Z S[0] S[1] D[1] D[2] S[2]
+ S[3] D[3] D[0]
M1000 Z a_1430_325# a_1643_311# VPB phighvt w=820000u l=180000u
+  ad=1.9024e+12p pd=1.776e+07u as=1.2606e+12p ps=1.174e+07u
M1001 a_1643_311# D[1] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.0912e+12p ps=4.808e+07u
M1002 a_2695_47# D[2] VGND VNB nshort w=650000u l=150000u
+  ad=7.618e+11p pd=8.38e+06u as=3.3176e+12p ps=3.4e+07u
M1003 VPWR D[0] a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.2606e+12p ps=1.174e+07u
M1004 VPWR S[0] a_559_265# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1005 a_2693_297# D[2] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.2606e+12p pd=1.174e+07u as=0p ps=0u
M1006 VPWR D[1] a_1643_311# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Z S[1] a_1693_66# VNB nshort w=520000u l=150000u
+  ad=1.1232e+12p pd=1.264e+07u as=7.618e+11p ps=8.38e+06u
M1008 Z S[2] a_2695_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_2695_47# S[2] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR D[3] a_4219_311# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.2606e+12p ps=1.174e+07u
M1011 Z S[3] a_4269_66# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=7.618e+11p ps=8.38e+06u
M1012 a_4269_66# S[3] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND D[3] a_4269_66# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1643_311# a_1430_325# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_119_47# S[0] Z VNB nshort w=520000u l=150000u
+  ad=7.618e+11p pd=8.38e+06u as=0p ps=0u
M1016 a_1693_66# S[1] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND D[1] a_1693_66# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_559_265# S[0] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR D[2] a_2693_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_3135_265# S[2] VPWR VPB phighvt w=820000u l=180000u
+  ad=2.378e+11p pd=2.22e+06u as=0p ps=0u
M1021 VGND D[2] a_2695_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Z S[3] a_4269_66# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Z S[0] a_119_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND D[0] a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_2693_297# a_3135_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Z S[1] a_1693_66# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_4219_311# D[3] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_119_47# S[0] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1693_66# D[1] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_2695_47# S[2] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_4269_66# S[3] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_4269_66# D[3] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1693_66# S[1] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_2695_47# D[2] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR D[3] a_4219_311# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR S[1] a_1430_325# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1037 Z S[0] a_119_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1643_311# D[1] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_4219_311# a_4006_325# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_4269_66# D[3] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_117_297# D[0] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_117_297# a_559_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 Z a_1430_325# a_1643_311# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1044 Z a_3135_265# a_2693_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_4006_325# S[3] VPWR VPB phighvt w=820000u l=180000u
+  ad=2.378e+11p pd=2.22e+06u as=0p ps=0u
M1046 a_559_265# S[0] VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1047 a_2693_297# D[2] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1048 Z a_4006_325# a_4219_311# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1049 VGND D[1] a_1693_66# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1050 a_1430_325# S[1] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1051 a_2693_297# a_3135_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1052 VGND D[2] a_2695_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1053 VGND S[0] a_559_265# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1054 VGND D[3] a_4269_66# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1055 VPWR D[0] a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1056 Z a_559_265# a_117_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1057 a_119_47# D[0] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1058 VGND S[2] a_3135_265# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1059 VGND S[3] a_4006_325# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1060 a_4219_311# a_4006_325# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1061 VGND S[1] a_1430_325# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1062 a_3135_265# S[2] VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1063 a_117_297# a_559_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1064 Z a_3135_265# a_2693_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1065 VPWR D[1] a_1643_311# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1066 a_1643_311# a_1430_325# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1067 VPWR S[3] a_4006_325# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1068 Z a_4006_325# a_4219_311# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1069 a_1430_325# S[1] VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1070 a_4219_311# D[3] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1071 a_117_297# D[0] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1072 Z a_559_265# a_117_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1073 VGND D[0] a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1074 VPWR D[2] a_2693_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1075 a_4006_325# S[3] VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1076 VPWR S[2] a_3135_265# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1077 Z S[2] a_2695_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1078 a_119_47# D[0] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1079 a_1693_66# D[1] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o32ai_2 A1 B1 A2 A3 Y B2 VPB VNB VGND VPWR
M1000 VGND A2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=1.0595e+12p pd=7.16e+06u as=1.469e+12p ps=1.232e+07u
M1001 a_27_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=8.3e+11p pd=7.66e+06u as=5.8e+11p ps=5.16e+06u
M1002 Y A3 a_525_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.7e+11p ps=7.74e+06u
M1003 a_27_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.81e+11p ps=4.08e+06u
M1004 VGND A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_807_297# VPB phighvt w=1e+06u l=180000u
+  ad=8.5e+11p pd=7.7e+06u as=5.8e+11p ps=5.16e+06u
M1007 Y B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_525_297# A2 a_807_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_807_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_807_297# A2 a_525_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_525_297# A3 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A3 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o221a_4 C1 A1 A2 B1 B2 X VNB VPB VGND VPWR
M1000 a_307_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=7.67e+11p pd=7.56e+06u as=9.945e+11p ps=9.56e+06u
M1001 VPWR C1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.22e+12p pd=1.644e+07u as=8.7e+11p ps=7.74e+06u
M1002 a_27_47# C1 a_117_297# VNB nshort w=650000u l=150000u
+  ad=8.19e+11p pd=7.72e+06u as=2.08e+11p ps=1.94e+06u
M1003 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=0p ps=0u
M1004 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1005 VPWR A1 a_785_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1006 VPWR B1 a_305_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1007 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_117_297# C1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A1 a_307_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_305_297# B2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_785_297# A2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_47# B1 a_307_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_307_47# B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_117_297# B2 a_305_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_307_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_117_297# C1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_117_297# A2 a_785_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_305_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_47# B2 a_307_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A2 a_307_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_785_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_307_47# B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or3b_2 A B C_N X VPWR VGND VPB VNB
M1000 a_448_297# A VPWR VPB phighvt w=420000u l=180000u
+  ad=1.302e+11p pd=1.46e+06u as=6.164e+11p ps=5.43e+06u
M1001 X a_186_21# VGND VNB nshort w=650000u l=150000u
+  ad=3.4125e+11p pd=2.35e+06u as=5.5575e+11p ps=5.52e+06u
M1002 VGND B a_186_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.268e+11p ps=2.76e+06u
M1003 a_186_21# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_546_297# B a_448_297# VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1005 a_186_21# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR C_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1007 VPWR a_186_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=4e+11p ps=2.8e+06u
M1008 a_186_21# a_27_47# a_546_297# VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1009 VGND C_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1010 X a_186_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_186_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__xor2_2 B VPWR VGND X A VPB VNB
M1000 X B a_510_47# VNB nshort w=650000u l=150000u
+  ad=5.1675e+11p pd=4.19e+06u as=5.785e+11p ps=5.68e+06u
M1001 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=9.25e+11p pd=7.85e+06u as=8.45e+11p ps=7.69e+06u
M1002 VGND A a_112_47# VNB nshort w=650000u l=150000u
+  ad=1.06925e+12p pd=1.109e+07u as=4.485e+11p ps=3.98e+06u
M1003 VGND A a_510_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_510_47# B X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_510_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.39e+12p pd=1.278e+07u as=0p ps=0u
M1006 a_27_297# B a_112_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1007 a_510_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_112_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_112_47# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B a_510_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_510_297# a_112_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1012 X a_112_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_112_47# a_510_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_112_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B a_112_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_112_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_510_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A a_510_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o21ba_2 B1_N A1 X A2 VNB VPB VGND VPWR
M1000 VPWR a_186_21# X VPB phighvt w=1e+06u l=180000u
+  ad=1.3807e+12p pd=8.86e+06u as=3.15e+11p ps=2.63e+06u
M1001 a_186_21# a_27_93# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.45e+11p pd=2.69e+06u as=0p ps=0u
M1002 VGND a_186_21# X VNB nshort w=650000u l=150000u
+  ad=5.66e+11p pd=5.73e+06u as=2.5675e+11p ps=2.09e+06u
M1003 X a_186_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_518_47# a_27_93# a_186_21# VNB nshort w=650000u l=150000u
+  ad=4.4525e+11p pd=3.97e+06u as=1.69e+11p ps=1.82e+06u
M1005 VPWR B1_N a_27_93# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1006 VGND A2 a_518_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_518_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_186_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_621_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.35e+11p ps=2.47e+06u
M1010 a_621_297# A2 a_186_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B1_N a_27_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
.ends
.subckt sky130_fd_sc_hdll__or4bb_2 A X B D_N C_N VPWR VGND VPB VNB
M1000 VPWR A a_614_297# VPB phighvt w=420000u l=180000u
+  ad=8.59325e+11p pd=7.99e+06u as=1.281e+11p ps=1.45e+06u
M1001 VGND C_N a_27_410# VNB nshort w=420000u l=150000u
+  ad=8.121e+11p pd=8.33e+06u as=1.302e+11p ps=1.46e+06u
M1002 a_336_413# a_216_93# VGND VNB nshort w=420000u l=150000u
+  ad=2.814e+11p pd=3.02e+06u as=0p ps=0u
M1003 a_216_93# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1004 VPWR a_336_413# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1005 X a_336_413# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_532_297# a_27_410# a_426_413# VPB phighvt w=420000u l=180000u
+  ad=9.66e+10p pd=1.3e+06u as=2.514e+11p ps=2.7e+06u
M1007 VGND A a_336_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_426_413# a_216_93# a_336_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1009 a_614_297# B a_532_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR C_N a_27_410# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1011 a_216_93# D_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
M1012 a_336_413# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_336_413# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1014 X a_336_413# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_27_410# a_336_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__dlxtn_4 D GATE_N Q VNB VPB VPWR VGND
M1000 a_709_47# a_211_363# a_609_413# VNB nshort w=360000u l=150000u
+  ad=1.32e+11p pd=1.49e+06u as=1.008e+11p ps=1.28e+06u
M1001 a_211_363# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=9.9375e+11p ps=1.015e+07u
M1002 Q a_774_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=1.3496e+12p ps=1.283e+07u
M1003 Q a_774_21# VGND VNB nshort w=650000u l=150000u
+  ad=4.16e+11p pd=3.88e+06u as=0p ps=0u
M1004 VPWR GATE_N a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1005 VGND a_774_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_503_369# a_319_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=2.042e+11p pd=1.98e+06u as=0p ps=0u
M1007 a_505_47# a_319_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.734e+11p pd=1.72e+06u as=0p ps=0u
M1008 a_609_413# a_27_47# a_505_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_774_21# a_709_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND D a_319_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1011 VPWR D a_319_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1012 Q a_774_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_774_21# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_609_413# a_774_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1015 a_703_413# a_27_47# a_609_413# VPB phighvt w=420000u l=180000u
+  ad=1.533e+11p pd=1.57e+06u as=1.218e+11p ps=1.42e+06u
M1016 VGND GATE_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1017 VPWR a_609_413# a_774_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1018 a_609_413# a_211_363# a_503_369# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_211_363# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1020 Q a_774_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_774_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_774_21# a_703_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_774_21# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand2_8 A B Y VNB VPB VGND VPWR
M1000 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=2.69e+12p pd=2.338e+07u as=2.32e+12p ps=2.064e+07u
M1001 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=1.8395e+12p pd=1.736e+07u as=8.645e+11p ps=7.86e+06u
M1006 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=8.645e+11p pd=7.86e+06u as=0p ps=0u
M1009 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o21bai_4 Y B1_N A1 A2 VNB VPB VGND VPWR
M1000 a_621_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.43e+12p pd=1.286e+07u as=1.43e+12p ps=1.286e+07u
M1001 Y a_33_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=0p ps=0u
M1002 Y A2 a_621_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A1 a_621_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_245_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=1.3455e+12p pd=1.324e+07u as=1.1115e+12p ps=9.92e+06u
M1005 VGND A1 a_245_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_245_47# a_33_297# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1007 a_245_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B1_N a_33_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1009 a_33_297# B1_N VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1010 VGND A2 a_245_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_33_297# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_621_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y a_33_297# a_245_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y a_33_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_621_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A2 a_621_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_245_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A2 a_245_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_245_47# a_33_297# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND A1 a_245_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_33_297# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR A1 a_621_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_245_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y a_33_297# a_245_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_621_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a22o_4 B1 B2 X A2 A1 VNB VPB VGND VPWR
M1000 a_1008_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=3.835e+11p pd=3.78e+06u as=1.3975e+12p ps=1.08e+07u
M1001 X a_96_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=1.43e+12p ps=1.286e+07u
M1002 VPWR A2 a_524_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.515e+12p ps=1.303e+07u
M1003 a_96_21# B1 a_524_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1004 VGND A2 a_1008_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_96_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_524_297# B1 a_96_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_96_21# VGND VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=0p ps=0u
M1008 VGND a_96_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_616_47# B1 a_96_21# VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=4.81e+11p ps=4.08e+06u
M1010 a_524_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1008_47# A1 a_96_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_96_21# B2 a_524_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_96_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND B2 a_616_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_96_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_96_21# B1 a_616_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A1 a_524_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_96_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_616_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_96_21# A1 a_1008_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_524_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_96_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_524_297# B2 a_96_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__dlygate4sd2_1 A X VPWR VGND VPB VNB
M1000 a_213_47# a_27_47# VGND VNB nshort w=420000u l=180000u
+  ad=1.092e+11p pd=1.36e+06u as=4.913e+11p ps=3.91e+06u
M1001 X a_319_93# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1002 VPWR a_213_47# a_319_93# VPB phighvt w=420000u l=180000u
+  ad=6.233e+11p pd=4.51e+06u as=1.176e+11p ps=1.4e+06u
M1003 X a_319_93# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1004 a_213_47# a_27_47# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1005 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1006 VGND a_213_47# a_319_93# VNB nshort w=420000u l=180000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1007 VPWR A a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
.ends
.subckt sky130_fd_sc_hdll__nand4bb_1 C D A_N Y B_N VNB VPB VPWR VGND
M1000 VPWR B_N a_27_93# VPB phighvt w=420000u l=180000u
+  ad=1.1325e+12p pd=8.99e+06u as=1.134e+11p ps=1.38e+06u
M1001 VPWR a_500_21# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=7e+11p ps=5.4e+06u
M1002 a_434_47# a_27_93# a_334_47# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=2.275e+11p ps=2e+06u
M1003 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_334_47# C a_218_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.795e+11p ps=2.16e+06u
M1005 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_500_21# a_434_47# VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=0p ps=0u
M1007 a_218_47# D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.372e+11p ps=3.45e+06u
M1008 a_500_21# A_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.365e+11p pd=1.49e+06u as=0p ps=0u
M1009 Y a_27_93# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_500_21# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.533e+11p pd=1.57e+06u as=0p ps=0u
M1011 VGND B_N a_27_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
.ends
.subckt sky130_fd_sc_hdll__clkbuf_12 A X VPB VNB VGND VPWR
M1000 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=2.57e+12p pd=2.314e+07u as=1.74e+12p ps=1.548e+07u
M1001 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=6.804e+11p pd=8.28e+06u as=1.3482e+12p ps=1.398e+07u
M1002 VPWR A a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1003 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A a_117_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.268e+11p ps=2.76e+06u
M1010 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_117_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_117_297# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_117_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND A a_117_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_117_297# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor3b_2 C_N Y A B VPB VNB VGND VPWR
M1000 Y a_571_21# a_309_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u
M1001 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=4.034e+11p pd=3.96e+06u as=8.7e+11p ps=7.74e+06u
M1002 VGND C_N a_571_21# VNB nshort w=420000u l=150000u
+  ad=1.0662e+12p pd=1.084e+07u as=1.092e+11p ps=1.36e+06u
M1003 a_27_297# B a_309_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_309_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_571_21# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=6.89e+11p ps=6.02e+06u
M1006 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y a_571_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR C_N a_571_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1010 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_309_297# a_571_21# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__muxb16to1_1 Z VGND VPWR VNB VPB D[0] S[12] S[13] S[8] S[9]
+ S[10] S[11] S[14] S[15] D[12] D[9] D[10] D[13] D[14] D[15] D[8] D[11] S[0] S[1]
+ D[1] D[2] S[2] S[3] D[4] S[4] S[5] D[5] D[6] S[6] S[7] D[7] D[3]
M1000 Z a_1012_793# a_945_591# VPB phighvt w=820000u l=180000u
+  ad=3.5424e+12p pd=3.488e+07u as=3.297e+11p ps=2.69e+06u
M1001 a_1765_47# D[4] VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=3.7518e+12p ps=3.424e+07u
M1002 a_937_47# D[2] VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1003 a_2593_47# D[6] VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1004 Z a_2668_793# a_2601_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=3.297e+11p ps=2.69e+06u
M1005 a_1773_297# D[4] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=6.38e+12p ps=4.876e+07u
M1006 a_1773_591# D[12] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1007 VGND S[6] a_2668_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.61e+06u
M1008 a_2390_591# a_2189_937# Z VPB phighvt w=820000u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1009 a_1361_47# S[3] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1010 VPWR D[7] a_3218_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.297e+11p ps=2.69e+06u
M1011 a_937_911# D[10] VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1012 a_1361_937# S[11] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1013 VPWR D[15] a_3218_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.297e+11p ps=2.69e+06u
M1014 Z a_1840_265# a_1773_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1574_47# S[3] Z VNB nshort w=520000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=2.1632e+12p ps=2.496e+07u
M1016 a_2402_937# S[13] Z VNB nshort w=520000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1017 a_734_333# a_533_47# Z VPB phighvt w=820000u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1018 Z S[2] a_937_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_3017_47# S[7] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1020 a_2402_47# S[5] Z VNB nshort w=520000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1021 a_3017_937# S[15] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1022 a_1562_333# a_1361_47# Z VPB phighvt w=820000u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1023 a_746_47# S[1] Z VNB nshort w=520000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1024 VGND S[12] a_1840_793# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.61e+06u
M1025 a_109_911# D[8] VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1026 VGND S[14] a_2668_793# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.61e+06u
M1027 a_117_297# D[0] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1028 VPWR D[3] a_1562_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_2601_297# D[6] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1030 Z S[4] a_1765_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_533_937# S[9] VGND VNB nshort w=520000u l=150000u
+  ad=1.482e+11p pd=1.61e+06u as=0p ps=0u
M1032 a_117_591# D[8] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1033 VPWR D[11] a_1562_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.297e+11p ps=2.69e+06u
M1034 VGND D[15] a_3230_937# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.95e+06u
M1035 a_2601_591# D[14] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Z a_184_265# a_117_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1765_911# D[12] VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1038 a_3218_591# a_3017_937# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_533_47# S[1] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1040 a_945_297# D[2] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1041 Z a_1012_265# a_945_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_533_937# S[9] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1043 VGND D[11] a_1574_937# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.95e+06u
M1044 a_945_591# D[10] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VPWR S[0] a_184_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1046 a_2189_47# S[5] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1047 a_746_937# S[9] Z VNB nshort w=520000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1048 VPWR S[8] a_184_793# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1049 a_2189_937# S[13] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1050 VPWR S[2] a_1012_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1051 Z a_2668_265# a_2601_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1052 a_1361_47# S[3] VGND VNB nshort w=520000u l=150000u
+  ad=1.482e+11p pd=1.61e+06u as=0p ps=0u
M1053 VPWR S[10] a_1012_793# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1054 a_3230_937# S[15] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1055 a_533_47# S[1] VGND VNB nshort w=520000u l=150000u
+  ad=1.482e+11p pd=1.61e+06u as=0p ps=0u
M1056 Z S[8] a_109_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1057 VGND D[9] a_746_937# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1058 VGND S[0] a_184_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.61e+06u
M1059 a_2390_333# a_2189_47# Z VPB phighvt w=820000u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1060 a_3230_47# S[7] Z VNB nshort w=520000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1061 a_1361_937# S[11] VGND VNB nshort w=520000u l=150000u
+  ad=1.482e+11p pd=1.61e+06u as=0p ps=0u
M1062 VGND D[1] a_746_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1063 Z S[6] a_2593_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1064 Z a_1840_793# a_1773_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1065 Z S[10] a_937_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1066 VPWR S[6] a_2668_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1067 VGND S[8] a_184_793# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.61e+06u
M1068 a_1574_937# S[11] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1069 Z S[12] a_1765_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1070 a_2189_937# S[13] VGND VNB nshort w=520000u l=150000u
+  ad=1.482e+11p pd=1.61e+06u as=0p ps=0u
M1071 a_734_591# a_533_937# Z VPB phighvt w=820000u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1072 VPWR S[14] a_2668_793# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1073 a_3017_937# S[15] VGND VNB nshort w=520000u l=150000u
+  ad=1.482e+11p pd=1.61e+06u as=0p ps=0u
M1074 a_1562_591# a_1361_937# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1075 VPWR D[1] a_734_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1076 VPWR D[9] a_734_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1077 VPWR D[5] a_2390_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1078 a_2189_47# S[5] VGND VNB nshort w=520000u l=150000u
+  ad=1.482e+11p pd=1.61e+06u as=0p ps=0u
M1079 VPWR D[13] a_2390_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1080 VPWR S[4] a_1840_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1081 VGND D[3] a_1574_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1082 VGND S[10] a_1012_793# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.61e+06u
M1083 a_2593_911# D[14] VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1084 Z S[14] a_2593_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1085 VPWR S[12] a_1840_793# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1086 a_109_47# D[0] VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1087 VGND D[5] a_2402_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1088 VGND S[2] a_1012_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.61e+06u
M1089 VGND D[7] a_3230_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1090 Z a_184_793# a_117_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1091 VGND D[13] a_2402_937# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1092 Z S[0] a_109_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1093 a_3218_333# a_3017_47# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1094 VGND S[4] a_1840_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.61e+06u
M1095 a_3017_47# S[7] VGND VNB nshort w=520000u l=150000u
+  ad=1.482e+11p pd=1.61e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o221ai_2 B1 B2 Y A2 A1 C1 VNB VPB VGND VPWR
M1000 VPWR B1 a_410_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.745e+12p pd=1.149e+07u as=5.8e+11p ps=5.16e+06u
M1001 VGND A2 a_320_47# VNB nshort w=650000u l=150000u
+  ad=3.835e+11p pd=3.78e+06u as=1.1115e+12p ps=9.92e+06u
M1002 Y C1 a_28_47# VNB nshort w=650000u l=150000u
+  ad=2.08e+11p pd=1.94e+06u as=7.54e+11p ps=7.52e+06u
M1003 a_28_47# B1 a_320_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_410_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.7e+11p ps=7.74e+06u
M1005 a_802_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1006 Y C1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_320_47# B2 a_28_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B2 a_410_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A1 a_320_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_410_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A1 a_802_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_320_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_28_47# C1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_320_47# B1 a_28_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_28_47# B2 a_320_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_802_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_320_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A2 a_802_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__ebufn_1 Z TE_B A VNB VPB VPWR VGND
M1000 Z a_27_47# a_543_47# VNB nshort w=650000u l=150000u
+  ad=3.055e+11p pd=2.24e+06u as=1.365e+11p ps=1.72e+06u
M1001 VPWR A a_27_47# VPB phighvt w=640000u l=180000u
+  ad=4.656e+11p pd=4.42e+06u as=1.728e+11p ps=1.82e+06u
M1002 a_543_47# a_211_369# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.6525e+11p ps=3.83e+06u
M1003 a_411_297# TE_B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.8e+11p pd=3.76e+06u as=0p ps=0u
M1004 Z a_27_47# a_411_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.95e+11p pd=2.79e+06u as=0p ps=0u
M1005 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1006 a_211_369# TE_B VGND VNB nshort w=420000u l=150000u
+  ad=2.814e+11p pd=2.18e+06u as=0p ps=0u
M1007 a_211_369# TE_B VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or2_4 X A B VNB VPB VGND VPWR
M1000 VGND a_35_297# X VNB nshort w=650000u l=150000u
+  ad=8.4175e+11p pd=7.79e+06u as=4.485e+11p ps=3.98e+06u
M1001 VPWR A a_129_297# VPB phighvt w=1e+06u l=180000u
+  ad=9.55e+11p pd=7.91e+06u as=2.3e+11p ps=2.46e+06u
M1002 X a_35_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1003 a_129_297# B a_35_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1004 VGND A a_35_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1005 X a_35_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_35_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_35_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_35_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_35_297# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_35_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_35_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a21oi_4 B1 A2 A1 Y VNB VPB VGND VPWR
M1000 VPWR A1 a_28_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.21e+12p pd=1.042e+07u as=2.075e+12p ps=1.815e+07u
M1001 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=1.014e+12p pd=9.62e+06u as=9.23e+11p ps=8.04e+06u
M1002 VPWR A2 a_28_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A1 a_28_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_502_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=8.255e+11p pd=7.74e+06u as=0p ps=0u
M1006 Y B1 a_28_297# VPB phighvt w=1e+06u l=180000u
+  ad=6e+11p pd=5.2e+06u as=0p ps=0u
M1007 a_28_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2 a_502_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 a_28_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_502_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_28_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A2 a_502_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A1 a_502_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_502_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_28_297# B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_28_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A1 a_502_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_28_297# B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_28_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR A2 a_28_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_502_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o31ai_2 A1 Y B1 A3 A2 VGND VPWR VPB VNB
M1000 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=7e+11p pd=5.4e+06u as=8.5e+11p ps=7.7e+06u
M1001 VPWR B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.5e+11p ps=7.7e+06u
M1002 a_27_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=1.01075e+12p pd=9.61e+06u as=1.0075e+12p ps=7e+06u
M1003 VGND A3 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A3 a_309_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1006 a_27_297# A2 a_309_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=2.86e+11p pd=2.18e+06u as=0p ps=0u
M1008 a_27_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_309_297# A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_309_297# A3 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o211a_4 A1 X C1 A2 B1 VNB VPB VGND VPWR
M1000 a_524_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=8.0275e+11p pd=7.67e+06u as=1.06925e+12p ps=9.79e+06u
M1001 a_80_21# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.09e+12p pd=8.18e+06u as=1.795e+12p ps=1.559e+07u
M1002 VPWR B1 a_80_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND A2 a_524_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR C1 a_80_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_80_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=6e+11p ps=5.2e+06u
M1006 a_80_21# A2 a_1010_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3e+11p ps=2.6e+06u
M1007 a_524_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_524_47# B1 a_818_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.5275e+11p ps=1.77e+06u
M1009 X a_80_21# VGND VNB nshort w=650000u l=150000u
+  ad=4.16e+11p pd=3.88e+06u as=0p ps=0u
M1010 VPWR a_80_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A1 a_1202_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3e+11p ps=2.6e+06u
M1012 X a_80_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_80_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_80_21# C1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_607_47# B1 a_524_47# VNB nshort w=650000u l=150000u
+  ad=1.365e+11p pd=1.72e+06u as=0p ps=0u
M1016 VGND A1 a_524_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_80_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1010_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_80_21# C1 a_607_47# VNB nshort w=650000u l=150000u
+  ad=3.5425e+11p pd=2.39e+06u as=0p ps=0u
M1020 a_1202_297# A2 a_80_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_80_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_80_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_818_47# C1 a_80_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__einvn_2 TE_B A Z VPWR VGND VPB VNB
M1000 VPWR TE_B a_222_309# VPB phighvt w=940000u l=180000u
+  ad=5.526e+11p pd=4.99e+06u as=5.626e+11p ps=5.04e+06u
M1001 VPWR TE_B a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1002 a_222_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_234_47# A Z VNB nshort w=650000u l=150000u
+  ad=6.5975e+11p pd=5.93e+06u as=2.08e+11p ps=1.94e+06u
M1004 VGND TE_B a_27_47# VNB nshort w=420000u l=150000u
+  ad=2.847e+11p pd=3.2e+06u as=1.302e+11p ps=1.46e+06u
M1005 a_234_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_27_47# a_234_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Z A a_222_309# VPB phighvt w=1e+06u l=180000u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
M1008 Z A a_234_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_222_309# A Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sdfsbp_1 SCD CLK Q_N D Q VPWR VGND SET_B SCE VPB VNB
M1000 VGND a_349_21# a_295_47# VNB nshort w=420000u l=150000u
+  ad=1.4601e+12p pd=1.494e+07u as=1.134e+11p ps=1.38e+06u
M1001 a_1930_295# a_1735_329# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1002 Q a_2632_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=1.9705e+12p ps=1.846e+07u
M1003 a_1930_295# a_1735_329# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1004 a_1075_413# a_877_369# a_199_47# VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=2.99e+11p ps=3.24e+06u
M1005 VGND SCE a_349_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1006 a_1735_329# a_877_369# a_1655_47# VNB nshort w=640000u l=150000u
+  ad=3.054e+11p pd=2.42e+06u as=4.736e+11p ps=2.76e+06u
M1007 VPWR SCD a_27_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=3.456e+11p ps=3.64e+06u
M1008 a_1219_21# a_1075_413# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.701e+11p pd=1.65e+06u as=0p ps=0u
M1009 a_1870_413# a_877_369# a_1735_329# VPB phighvt w=420000u l=180000u
+  ad=1.302e+11p pd=1.46e+06u as=4.305e+11p ps=4.05e+06u
M1010 a_1655_47# a_1075_413# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Q a_2632_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1012 VPWR SCE a_349_21# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1013 a_1735_329# a_693_369# a_1652_329# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=1.974e+11p ps=2.15e+06u
M1014 a_1735_329# SET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND CLK a_693_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1016 a_877_369# a_693_369# VGND VNB nshort w=420000u l=150000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
M1017 VPWR a_1930_295# a_1870_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1467_47# a_1075_413# a_1219_21# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.512e+11p ps=1.56e+06u
M1019 a_27_369# a_349_21# a_199_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR SET_B a_1219_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1177_47# a_877_369# a_1075_413# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.344e+11p ps=1.48e+06u
M1022 VGND SET_B a_1467_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_877_369# a_693_369# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1024 a_199_47# SCE a_109_47# VNB nshort w=420000u l=150000u
+  ad=2.688e+11p pd=2.96e+06u as=1.26e+11p ps=1.44e+06u
M1025 VGND a_1219_21# a_1177_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Q_N a_1735_329# VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=0p ps=0u
M1027 a_1075_413# a_693_369# a_199_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_295_47# D a_199_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1652_329# a_1075_413# VPWR VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_1735_329# a_2632_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1031 a_211_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=1.472e+11p pd=1.74e+06u as=0p ps=0u
M1032 Q_N a_1735_329# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1033 a_109_47# SCD VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_2049_47# a_1930_295# a_1977_47# VNB nshort w=420000u l=150000u
+  ad=2.688e+11p pd=2.12e+06u as=8.82e+10p ps=1.26e+06u
M1035 VGND a_1735_329# a_2632_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1036 a_199_47# D a_211_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1169_413# a_693_369# a_1075_413# VPB phighvt w=420000u l=180000u
+  ad=1.596e+11p pd=1.6e+06u as=0p ps=0u
M1038 VPWR a_1219_21# a_1169_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND SET_B a_2049_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VPWR CLK a_693_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1041 a_1977_47# a_693_369# a_1735_329# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or4_1 C A X B D VPWR VGND VPB VNB
M1000 a_27_297# D VGND VNB nshort w=420000u l=150000u
+  ad=3.15e+11p pd=3.18e+06u as=4.7985e+11p ps=4.92e+06u
M1001 X a_27_297# VGND VNB nshort w=650000u l=150000u
+  ad=2.73e+11p pd=2.14e+06u as=0p ps=0u
M1002 VGND A a_27_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_117_297# D a_27_297# VPB phighvt w=420000u l=180000u
+  ad=1.47e+11p pd=1.54e+06u as=1.134e+11p ps=1.38e+06u
M1004 VPWR A a_307_297# VPB phighvt w=420000u l=180000u
+  ad=3.107e+11p pd=2.72e+06u as=1.428e+11p ps=1.52e+06u
M1005 VGND C a_27_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_307_297# B a_223_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 a_27_297# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_27_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=4.3e+11p pd=2.86e+06u as=0p ps=0u
M1009 a_223_297# C a_117_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__inputiso0n_1 VPWR VGND X SLEEP_B A VPB VNB
M1000 X a_27_75# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.7e+11p pd=2.74e+06u as=4.691e+11p ps=4.24e+06u
M1001 X a_27_75# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=2.446e+11p ps=2.18e+06u
M1002 a_27_75# A VPWR VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
M1003 VGND SLEEP_B a_123_75# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1004 VPWR SLEEP_B a_27_75# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_123_75# A a_27_75# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
.ends
.subckt sky130_fd_sc_hdll__and4bb_1 VNB VPB VGND VPWR A_N D X C B_N
M1000 a_425_93# a_27_47# a_339_93# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.176e+11p ps=1.4e+06u
M1001 a_615_93# C a_511_93# VNB nshort w=420000u l=150000u
+  ad=1.89e+11p pd=1.74e+06u as=1.554e+11p ps=1.58e+06u
M1002 a_339_93# C VPWR VPB phighvt w=420000u l=180000u
+  ad=2.814e+11p pd=3.02e+06u as=6.779e+11p ps=7.03e+06u
M1003 a_511_93# a_225_413# a_425_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_225_413# B_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1005 VPWR a_225_413# a_339_93# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR D a_339_93# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_225_413# B_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=3.861e+11p ps=3.65e+06u
M1008 VGND A_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1009 VGND D a_615_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_339_93# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1011 VPWR A_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
M1012 a_339_93# a_27_47# VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_339_93# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__clkinvlp_4 A Y VNB VPB VPWR VGND
M1000 Y A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=5.4e+11p pd=5.08e+06u as=7.9e+11p ps=7.58e+06u
M1001 Y A a_110_47# VNB nshort w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=1.155e+11p ps=1.52e+06u
M1002 VPWR A Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_110_47# A VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=2.8875e+11p ps=3.25e+06u
M1004 VGND A a_268_47# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.52e+06u
M1005 a_268_47# A Y VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a32o_2 B2 X A2 A3 A1 B1 VNB VPB VGND VPWR
M1000 X a_21_199# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=1.01e+12p ps=8.02e+06u
M1001 VGND a_21_199# X VNB nshort w=650000u l=150000u
+  ad=8.5475e+11p pd=6.53e+06u as=2.08e+11p ps=1.94e+06u
M1002 VPWR A1 a_319_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.5e+11p ps=7.7e+06u
M1003 VPWR a_21_199# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_21_199# B1 a_382_47# VNB nshort w=650000u l=150000u
+  ad=2.47e+11p pd=2.06e+06u as=2.3075e+11p ps=2.01e+06u
M1005 a_319_297# B1 a_21_199# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1006 VPWR A3 a_319_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_589_47# A1 a_21_199# VNB nshort w=650000u l=150000u
+  ad=3.445e+11p pd=2.36e+06u as=0p ps=0u
M1008 a_21_199# B2 a_319_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_21_199# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_725_47# A2 a_589_47# VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1011 a_319_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_382_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A3 a_725_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand3b_1 B C A_N Y VPB VNB VGND VPWR
M1000 VPWR A_N a_53_93# VPB phighvt w=420000u l=180000u
+  ad=6.057e+11p pd=5.31e+06u as=1.134e+11p ps=1.38e+06u
M1001 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.9e+11p ps=5.18e+06u
M1002 a_348_47# B a_252_47# VNB nshort w=650000u l=150000u
+  ad=2.1125e+11p pd=1.95e+06u as=2.145e+11p ps=1.96e+06u
M1003 VGND A_N a_53_93# VNB nshort w=420000u l=150000u
+  ad=2.33e+11p pd=2.07e+06u as=1.302e+11p ps=1.46e+06u
M1004 Y a_53_93# a_348_47# VNB nshort w=650000u l=150000u
+  ad=1.8525e+11p pd=1.87e+06u as=0p ps=0u
M1005 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_252_47# C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y a_53_93# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and2_6 X B A VNB VPB VGND VPWR
M1000 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=1.72e+12p pd=1.544e+07u as=8.7e+11p ps=7.74e+06u
M1001 VGND B a_293_47# VNB nshort w=650000u l=150000u
+  ad=1.2155e+12p pd=1.024e+07u as=1.82e+11p ps=1.86e+06u
M1002 VPWR A a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1003 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=5.265e+11p ps=5.52e+06u
M1005 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_117_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_293_47# A a_117_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1009 a_117_297# A a_131_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.56e+11p ps=1.78e+06u
M1010 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_131_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR B a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_117_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a22oi_2 A1 A2 B1 B2 Y VPWR VGND VPB VNB
M1000 Y B2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=8.3e+11p pd=7.66e+06u as=1.51e+12p ps=1.302e+07u
M1001 a_27_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=5.46e+11p pd=5.58e+06u as=4.485e+11p ps=3.98e+06u
M1002 a_507_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=6.11e+11p pd=5.78e+06u as=4.485e+11p ps=3.98e+06u
M1003 a_117_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1004 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_507_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A1 a_507_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_117_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_117_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A2 a_507_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_117_297# B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__muxb4to1_2 VGND VPWR Z VNB VPB S[1] S[2] S[3] D[1] D[0]
+ D[2] D[3] S[0]
M1000 VPWR D[2] a_1315_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.88e+12p pd=1.576e+07u as=8.211e+11p ps=7.41e+06u
M1001 VPWR D[3] a_2112_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.211e+11p ps=7.41e+06u
M1002 a_27_297# D[0] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1003 Z a_1566_265# a_1315_297# VPB phighvt w=820000u l=180000u
+  ad=9.512e+11p pd=8.88e+06u as=0p ps=0u
M1004 Z a_1989_47# a_2112_333# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_297# a_278_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR S[0] a_278_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1007 a_1989_47# S[3] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=9.828e+11p ps=1.052e+07u
M1008 a_2133_69# D[3] VGND VNB nshort w=650000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1009 Z a_278_265# a_27_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_845_69# S[1] Z VNB nshort w=520000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=5.616e+11p ps=6.32e+06u
M1011 a_27_47# S[0] Z VNB nshort w=520000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1012 Z S[1] a_845_69# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_47# D[0] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Z S[0] a_27_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_824_333# D[1] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1016 a_1989_47# S[3] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1017 VPWR D[0] a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_701_47# S[1] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1019 VGND D[1] a_845_69# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_824_333# a_701_47# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND S[0] a_278_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1022 a_701_47# S[1] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1023 VPWR D[1] a_824_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_845_69# D[1] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Z S[3] a_2133_69# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND D[0] a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Z a_701_47# a_824_333# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1315_47# D[2] VGND VNB nshort w=650000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1029 Z S[2] a_1315_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1315_297# D[2] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1315_297# a_1566_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_2112_333# a_1989_47# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND D[2] a_1315_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_2133_69# S[3] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR S[2] a_1566_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1036 a_2112_333# D[3] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1315_47# S[2] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND S[2] a_1566_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1039 VGND D[3] a_2133_69# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sdfrbp_1 RESET_B VPWR VGND VNB VPB Q_N D CLK Q SCE SCD
M1000 a_1428_47# a_1380_303# a_1322_47# VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.518e+11p ps=1.6e+06u
M1001 a_213_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=1.5405e+12p ps=1.444e+07u
M1002 VPWR a_1972_21# a_1951_413# VPB phighvt w=420000u l=180000u
+  ad=1.88075e+12p pd=1.788e+07u as=1.386e+11p ps=1.5e+06u
M1003 a_1972_21# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=1.344e+11p pd=1.48e+06u as=0p ps=0u
M1004 Q a_1972_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.15e+11p pd=2.63e+06u as=0p ps=0u
M1005 a_2157_47# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=0p ps=0u
M1006 VPWR SCD a_870_389# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=1.971e+11p ps=1.81e+06u
M1007 a_700_389# D a_631_119# VNB nshort w=420000u l=150000u
+  ad=3.3215e+11p pd=3.47e+06u as=1.302e+11p ps=1.46e+06u
M1008 a_1380_303# a_1202_413# VPWR VPB phighvt w=840000u l=180000u
+  ad=2.541e+11p pd=2.37e+06u as=0p ps=0u
M1009 a_1202_413# a_27_47# a_700_389# VNB nshort w=360000u l=150000u
+  ad=1.44e+11p pd=1.52e+06u as=0p ps=0u
M1010 VPWR a_1757_47# a_1972_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1972_21# a_1757_47# a_2157_47# VNB nshort w=420000u l=150000u
+  ad=1.365e+11p pd=1.49e+06u as=0p ps=0u
M1012 Q a_1972_21# VGND VNB nshort w=650000u l=150000u
+  ad=1.9825e+11p pd=1.91e+06u as=0p ps=0u
M1013 VPWR a_1380_303# a_1324_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1014 VPWR a_1972_21# a_2580_47# VPB phighvt w=790000u l=180000u
+  ad=0p pd=0u as=2.133e+11p ps=2.12e+06u
M1015 VPWR CLK a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1016 a_618_389# SCE VPWR VPB phighvt w=540000u l=180000u
+  ad=1.242e+11p pd=1.54e+06u as=0p ps=0u
M1017 a_1951_413# a_213_47# a_1757_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1018 VGND a_1972_21# a_2580_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.61e+06u
M1019 a_700_389# D a_618_389# VPB phighvt w=540000u l=180000u
+  ad=5.193e+11p pd=4.01e+06u as=0p ps=0u
M1020 a_631_119# a_331_66# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND RESET_B a_1428_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1324_413# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1202_413# a_213_47# a_700_389# VPB phighvt w=420000u l=180000u
+  ad=1.806e+11p pd=1.7e+06u as=0p ps=0u
M1024 a_1324_413# a_27_47# a_1202_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1866_47# a_27_47# a_1757_47# VNB nshort w=360000u l=150000u
+  ad=2.121e+11p pd=1.9e+06u as=1.422e+11p ps=1.51e+06u
M1026 a_1757_47# a_213_47# a_1380_303# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.87e+11p ps=1.93e+06u
M1027 VPWR SCE a_331_66# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=2.214e+11p ps=1.9e+06u
M1028 VGND CLK a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1029 VGND a_1972_21# a_1866_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_213_47# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
M1031 Q_N a_2580_47# VGND VNB nshort w=520000u l=150000u
+  ad=1.456e+11p pd=1.6e+06u as=0p ps=0u
M1032 a_899_66# SCE a_700_389# VNB nshort w=420000u l=500000u
+  ad=1.554e+11p pd=1.58e+06u as=0p ps=0u
M1033 Q_N a_2580_47# VPWR VPB phighvt w=790000u l=180000u
+  ad=2.291e+11p pd=2.16e+06u as=0p ps=0u
M1034 a_1757_47# a_27_47# a_1380_303# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1322_47# a_213_47# a_1202_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND SCD a_899_66# VNB nshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_870_389# a_331_66# a_700_389# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND SCE a_331_66# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1039 a_1380_303# a_1202_413# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o221a_2 B2 A2 X B1 C1 A1 VPB VNB VGND VPWR
M1000 a_255_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.45e+11p pd=2.49e+06u as=9.7e+11p ps=7.94e+06u
M1001 a_245_47# B1 a_151_47# VNB nshort w=650000u l=150000u
+  ad=3.9325e+11p pd=3.81e+06u as=3.9975e+11p ps=3.83e+06u
M1002 a_151_47# C1 a_38_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.6975e+11p ps=2.13e+06u
M1003 a_151_47# B2 a_245_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A1 a_245_47# VNB nshort w=650000u l=150000u
+  ad=5.46e+11p pd=5.58e+06u as=0p ps=0u
M1005 VPWR A1 a_535_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.3e+11p ps=2.46e+06u
M1006 a_535_297# A2 a_38_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.13e+12p ps=6.26e+06u
M1007 VPWR C1 a_38_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_245_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_38_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1010 a_38_47# B2 a_255_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_38_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.405e+11p ps=2.04e+06u
M1012 X a_38_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_38_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__dlxtn_2 D GATE_N Q VNB VPB VPWR VGND
M1000 a_211_363# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=7.76e+11p ps=8.18e+06u
M1001 a_718_47# a_211_363# a_608_413# VNB nshort w=360000u l=150000u
+  ad=1.32e+11p pd=1.49e+06u as=1.35e+11p ps=1.47e+06u
M1002 VPWR GATE_N a_27_47# VPB phighvt w=640000u l=180000u
+  ad=1.0446e+12p pd=1.022e+07u as=1.728e+11p ps=1.82e+06u
M1003 a_503_369# a_319_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=2.021e+11p pd=1.97e+06u as=0p ps=0u
M1004 VPWR a_783_21# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1005 a_739_413# a_27_47# a_608_413# VPB phighvt w=420000u l=180000u
+  ad=9.66e+10p pd=1.3e+06u as=1.995e+11p ps=1.79e+06u
M1006 a_505_47# a_319_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.554e+11p pd=1.62e+06u as=0p ps=0u
M1007 VGND a_783_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1008 Q a_783_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND D a_319_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1010 VPWR D a_319_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1011 VGND a_783_21# a_718_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Q a_783_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_608_413# a_27_47# a_505_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_608_413# a_783_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1015 VGND GATE_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1016 a_211_363# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1017 VPWR a_608_413# a_783_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1018 a_608_413# a_211_363# a_503_369# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_783_21# a_739_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a22o_2 A1 A2 X B2 B1 VPWR VGND VPB VNB
M1000 a_27_297# B1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=6.4e+11p ps=5.28e+06u
M1001 X a_27_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=1.01e+12p ps=8.02e+06u
M1002 VGND a_27_297# X VNB nshort w=650000u l=150000u
+  ad=6.955e+11p pd=6.04e+06u as=2.08e+11p ps=1.94e+06u
M1003 VPWR A2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_27_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_117_297# B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_411_47# A1 a_27_297# VNB nshort w=650000u l=150000u
+  ad=2.47e+11p pd=2.06e+06u as=4.03e+11p ps=3.84e+06u
M1007 VGND A2 a_411_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_117_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_119_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=1.495e+11p pd=1.76e+06u as=0p ps=0u
M1010 a_27_297# B1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_27_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand2_6 Y A B VPB VNB VGND VPWR
M1000 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=1.99e+12p pd=1.798e+07u as=1.74e+12p ps=1.548e+07u
M1001 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=1.248e+12p pd=1.294e+07u as=7.215e+11p ps=6.12e+06u
M1003 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=6.89e+11p pd=6.02e+06u as=0p ps=0u
M1006 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o21bai_2 B1_N Y A2 A1 VNB VPB VGND VPWR
M1000 a_226_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=8.0925e+11p pd=7.69e+06u as=6.112e+11p ps=5.54e+06u
M1001 a_226_47# a_28_297# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1002 Y a_28_297# a_226_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_28_297# B1_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1004 VPWR B1_N a_28_297# VPB phighvt w=420000u l=180000u
+  ad=8.657e+11p pd=7.83e+06u as=1.134e+11p ps=1.38e+06u
M1005 VPWR a_28_297# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1006 a_226_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_437_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.5e+11p pd=7.7e+06u as=0p ps=0u
M1008 VGND A1 a_226_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_28_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A1 a_437_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_437_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A2 a_226_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A2 a_437_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o21a_4 A1 A2 B1 X VNB VPB VPWR VGND
M1000 X a_80_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6e+11p pd=5.2e+06u as=1.76e+12p ps=1.352e+07u
M1001 a_80_21# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6.5e+11p pd=5.3e+06u as=0p ps=0u
M1002 X a_80_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_525_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=8.84e+11p pd=7.92e+06u as=1.0075e+12p ps=9.6e+06u
M1004 a_80_21# A2 a_826_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.5e+11p ps=2.5e+06u
M1005 X a_80_21# VGND VNB nshort w=650000u l=150000u
+  ad=4.29e+11p pd=3.92e+06u as=0p ps=0u
M1006 VGND a_80_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_525_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A1 a_1008_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3e+11p ps=2.6e+06u
M1009 X a_80_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_80_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR B1 a_80_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_525_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_525_47# B1 a_80_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1014 a_826_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_80_21# B1 a_525_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A1 a_525_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_80_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_80_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1008_297# A2 a_80_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a21oi_2 B1 A2 A1 Y VNB VPB VGND VPWR
M1000 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=1.25e+12p ps=1.05e+07u
M1001 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=7.54e+11p pd=6.22e+06u as=4.55e+11p ps=4e+06u
M1003 a_123_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=0p ps=0u
M1004 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_315_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=1.365e+11p pd=1.72e+06u as=0p ps=0u
M1006 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_315_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A1 a_123_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_297# B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1010 Y B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or2_2 B X A VPWR VGND VPB VNB
M1000 VPWR A a_129_297# VPB phighvt w=420000u l=180000u
+  ad=5.957e+11p pd=5.29e+06u as=9.66e+10p ps=1.3e+06u
M1001 X a_39_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=0p ps=0u
M1002 a_129_297# B a_39_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1003 VGND A a_39_297# VNB nshort w=420000u l=150000u
+  ad=5.337e+11p pd=5.39e+06u as=1.134e+11p ps=1.38e+06u
M1004 VGND a_39_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.405e+11p ps=2.04e+06u
M1005 X a_39_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_39_297# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_39_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__decap_12 VGND VPWR VPB VNB
M1000 VPWR VGND VPWR VPB phighvt w=870000u l=4.73e+06u
+  ad=4.524e+11p pd=4.52e+06u as=0p ps=0u
M1001 VGND VPWR VGND VNB nshort w=550000u l=4.73e+06u
+  ad=2.86e+11p pd=3.24e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o211a_2 C1 B1 A2 A1 X VNB VPB VPWR VGND
M1000 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=1.12e+12p pd=8.24e+06u as=3e+11p ps=2.6e+06u
M1001 a_120_47# C1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=2.0475e+11p ps=1.93e+06u
M1002 VPWR C1 a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.055e+12p ps=6.11e+06u
M1003 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_206_47# B1 a_120_47# VNB nshort w=650000u l=150000u
+  ad=3.7375e+11p pd=3.75e+06u as=0p ps=0u
M1005 a_206_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.4425e+11p ps=6.19e+06u
M1006 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=2.34e+11p pd=2.02e+06u as=0p ps=0u
M1007 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_47# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A1 a_206_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_406_297# A2 a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=2.3e+11p pd=2.46e+06u as=0p ps=0u
M1011 VPWR A1 a_406_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor2_4 Y A B VPB VNB VGND VPWR
M1000 Y B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=1.44e+12p ps=1.288e+07u
M1001 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1002 VGND A Y VNB nshort w=650000u l=150000u
+  ad=9.425e+11p pd=9.4e+06u as=8.97e+11p ps=7.96e+06u
M1003 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_297# B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_297# B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__inputiso1p_1 SLEEP X A VPB VNB VGND VPWR
M1000 a_44_297# A VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=3.517e+11p ps=3.53e+06u
M1001 VPWR SLEEP a_134_297# VPB phighvt w=420000u l=180000u
+  ad=3.057e+11p pd=2.71e+06u as=1.218e+11p ps=1.42e+06u
M1002 X a_44_297# VGND VNB nshort w=650000u l=150000u
+  ad=2.405e+11p pd=2.04e+06u as=0p ps=0u
M1003 VGND SLEEP a_44_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_134_297# A a_44_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1005 X a_44_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=4.1e+11p pd=2.82e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__dfstp_1 D VPWR CLK VGND Q VPB VNB SET_B
M1000 VPWR SET_B a_1126_413# VPB phighvt w=420000u l=180000u
+  ad=1.3883e+12p pd=1.359e+07u as=2.856e+11p ps=3.04e+06u
M1001 a_211_363# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.18655e+12p ps=1.1e+07u
M1002 a_506_47# a_27_47# a_409_329# VNB nshort w=360000u l=150000u
+  ad=1.8e+11p pd=1.72e+06u as=1.87e+11p ps=1.93e+06u
M1003 Q a_1738_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.2e+11p pd=2.64e+06u as=0p ps=0u
M1004 a_1344_47# a_27_47# a_1126_413# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.596e+11p ps=1.6e+06u
M1005 VGND a_1126_413# a_1738_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1006 VPWR CLK a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1007 VPWR a_1126_413# a_1738_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1008 VPWR a_702_21# a_610_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.974e+11p ps=1.78e+06u
M1009 Q a_1738_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.9825e+11p pd=1.91e+06u as=0p ps=0u
M1010 VPWR a_1288_261# a_1244_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=9.66e+10p ps=1.3e+06u
M1011 a_1126_413# a_211_363# a_1156_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1012 a_1044_413# a_506_47# VPWR VPB phighvt w=420000u l=180000u
+  ad=9.66e+10p pd=1.3e+06u as=0p ps=0u
M1013 a_409_329# D VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_409_329# D VPWR VPB phighvt w=840000u l=180000u
+  ad=2.625e+11p pd=2.39e+06u as=0p ps=0u
M1015 a_1156_47# a_506_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_636_47# a_211_363# a_506_47# VNB nshort w=360000u l=150000u
+  ad=1.341e+11p pd=1.5e+06u as=0p ps=0u
M1017 VPWR a_506_47# a_702_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1018 a_1288_261# a_1126_413# VPWR VPB phighvt w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1019 a_610_413# a_27_47# a_506_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1020 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1021 a_866_47# SET_B VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1022 VGND a_702_21# a_636_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1288_261# a_1126_413# VGND VNB nshort w=540000u l=150000u
+  ad=1.404e+11p pd=1.6e+06u as=0p ps=0u
M1024 a_1244_413# a_211_363# a_1126_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_702_21# a_506_47# a_866_47# VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1026 a_702_21# SET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_211_363# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1028 a_506_47# a_211_363# a_409_329# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1416_47# a_1288_261# a_1344_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1030 a_1126_413# a_27_47# a_1044_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND SET_B a_1416_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand4b_4 C D B Y A_N VNB VPB VGND VPWR
M1000 a_225_47# B a_693_47# VNB nshort w=650000u l=150000u
+  ad=9.945e+11p pd=9.56e+06u as=8.32e+11p ps=7.76e+06u
M1001 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.32e+12p pd=2.064e+07u as=3.36e+12p ps=2.672e+07u
M1002 VGND D a_1081_47# VNB nshort w=650000u l=150000u
+  ad=5.85e+11p pd=5.7e+06u as=9.945e+11p ps=9.56e+06u
M1003 a_693_47# B a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_225_47# a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1010 Y a_27_47# a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A_N a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1012 a_1081_47# D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_225_47# a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1081_47# C a_693_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_693_47# C a_1081_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_225_47# B a_693_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A_N a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1024 VGND D a_1081_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y a_27_47# a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_693_47# B a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1081_47# D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1081_47# C a_693_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_693_47# C a_1081_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand2_12 Y A B VPB VNB VGND VPWR
M1000 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=3.73e+12p pd=3.346e+07u as=3.48e+12p ps=3.096e+07u
M1001 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=2.3335e+12p pd=2.408e+07u as=1.443e+12p ps=1.224e+07u
M1004 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=1.378e+12p pd=1.204e+07u as=0p ps=0u
M1008 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__buf_12 A X VGND VPWR VPB VNB
M1000 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=2.61e+12p pd=2.322e+07u as=1.74e+12p ps=1.548e+07u
M1001 VPWR A a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1002 VGND A a_117_297# VNB nshort w=650000u l=150000u
+  ad=1.82e+12p pd=1.73e+07u as=4.16e+11p ps=3.88e+06u
M1003 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.2805e+12p ps=1.174e+07u
M1007 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_117_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_117_297# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A a_117_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_117_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_117_297# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a21o_8 A2 A1 X B1 VNB VPB VGND VPWR
M1000 VGND A2 a_297_47# VNB nshort w=650000u l=150000u
+  ad=1.9305e+12p pd=1.504e+07u as=1.69e+11p ps=1.82e+06u
M1001 X a_213_47# VGND VNB nshort w=650000u l=150000u
+  ad=7.02e+11p pd=7.36e+06u as=0p ps=0u
M1002 VGND a_213_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.12e+12p pd=1.024e+07u as=1.99e+12p ps=1.798e+07u
M1004 a_213_47# A1 a_131_47# VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=1.69e+11p ps=1.82e+06u
M1005 X a_213_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=0p ps=0u
M1006 X a_213_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_213_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_297_47# A1 a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_297# B1 a_213_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1010 VGND a_213_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_213_47# B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_213_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_131_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_213_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_213_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_213_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_213_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_213_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_213_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 X a_213_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND B1 a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_213_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_213_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 X a_213_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sdfrtn_1 VPB VNB RESET_B VPWR VGND SCE SCD D CLK_N Q
M1000 a_1428_47# a_1380_303# a_1322_47# VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.518e+11p ps=1.6e+06u
M1001 a_213_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=1.3533e+12p ps=1.268e+07u
M1002 VPWR a_1972_21# a_1951_413# VPB phighvt w=420000u l=180000u
+  ad=1.6398e+12p pd=1.569e+07u as=1.386e+11p ps=1.5e+06u
M1003 a_1972_21# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=1.344e+11p pd=1.48e+06u as=0p ps=0u
M1004 Q a_1972_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.15e+11p pd=2.63e+06u as=0p ps=0u
M1005 a_2157_47# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=0p ps=0u
M1006 VPWR SCD a_870_389# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=1.971e+11p ps=1.81e+06u
M1007 a_700_389# D a_631_119# VNB nshort w=420000u l=150000u
+  ad=3.3215e+11p pd=3.47e+06u as=1.302e+11p ps=1.46e+06u
M1008 a_1380_303# a_1202_413# VPWR VPB phighvt w=840000u l=180000u
+  ad=2.541e+11p pd=2.37e+06u as=0p ps=0u
M1009 a_1202_413# a_213_47# a_700_389# VNB nshort w=360000u l=150000u
+  ad=1.44e+11p pd=1.52e+06u as=0p ps=0u
M1010 VPWR a_1757_47# a_1972_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1972_21# a_1757_47# a_2157_47# VNB nshort w=420000u l=150000u
+  ad=1.365e+11p pd=1.49e+06u as=0p ps=0u
M1012 Q a_1972_21# VGND VNB nshort w=650000u l=150000u
+  ad=1.9825e+11p pd=1.91e+06u as=0p ps=0u
M1013 VPWR a_1380_303# a_1324_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1014 VPWR CLK_N a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1015 a_618_389# SCE VPWR VPB phighvt w=540000u l=180000u
+  ad=1.242e+11p pd=1.54e+06u as=0p ps=0u
M1016 a_1951_413# a_27_47# a_1757_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1017 a_700_389# D a_618_389# VPB phighvt w=540000u l=180000u
+  ad=5.193e+11p pd=4.01e+06u as=0p ps=0u
M1018 a_631_119# a_331_66# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND RESET_B a_1428_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1324_413# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1202_413# a_27_47# a_700_389# VPB phighvt w=420000u l=180000u
+  ad=1.806e+11p pd=1.7e+06u as=0p ps=0u
M1022 a_1324_413# a_213_47# a_1202_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1866_47# a_213_47# a_1757_47# VNB nshort w=360000u l=150000u
+  ad=2.121e+11p pd=1.9e+06u as=1.422e+11p ps=1.51e+06u
M1024 a_1757_47# a_27_47# a_1380_303# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.87e+11p ps=1.93e+06u
M1025 VPWR SCE a_331_66# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=2.214e+11p ps=1.9e+06u
M1026 VGND CLK_N a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1027 VGND a_1972_21# a_1866_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_213_47# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
M1029 a_899_66# SCE a_700_389# VNB nshort w=420000u l=500000u
+  ad=1.554e+11p pd=1.58e+06u as=0p ps=0u
M1030 a_1757_47# a_213_47# a_1380_303# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1322_47# a_27_47# a_1202_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND SCD a_899_66# VNB nshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_870_389# a_331_66# a_700_389# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND SCE a_331_66# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1035 a_1380_303# a_1202_413# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o2bb2ai_4 A1_N B1 B2 A2_N Y VPB VNB VGND VPWR
M1000 VGND B2 a_887_47# VNB nshort w=650000u l=150000u
+  ad=1.3455e+12p pd=1.194e+07u as=1.6315e+12p ps=1.412e+07u
M1001 a_113_47# A1_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=3.08e+12p ps=2.416e+07u
M1002 a_113_47# A2_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_47# A2_N a_113_47# VNB nshort w=650000u l=150000u
+  ad=9.425e+11p pd=9.4e+06u as=4.485e+11p ps=3.98e+06u
M1004 VPWR a_113_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.16e+12p ps=1.032e+07u
M1005 VPWR B1 a_1361_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.43e+12p ps=1.286e+07u
M1006 Y a_113_47# a_887_47# VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=0p ps=0u
M1007 Y a_113_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_887_47# a_113_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B1 a_887_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A2_N a_113_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B2 a_1361_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_887_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_887_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1361_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A1_N a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B2 a_887_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_47# A1_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_113_47# A2_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_113_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR B1 a_1361_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_113_47# A2_N a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_47# A2_N a_113_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR A1_N a_113_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1361_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1361_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND B1 a_887_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_887_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_887_47# a_113_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR A2_N a_113_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y B2 a_1361_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND A1_N a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1361_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Y a_113_47# a_887_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_887_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_113_47# A1_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Y a_113_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_113_47# A2_N a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_27_47# A1_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR A1_N a_113_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor4_1 D C Y A B VPB VNB VGND VPWR
M1000 a_221_297# C a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=3.4e+11p ps=2.68e+06u
M1001 VGND C Y VNB nshort w=650000u l=150000u
+  ad=6.045e+11p pd=5.76e+06u as=4.29e+11p ps=3.92e+06u
M1002 VPWR A a_317_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=3.1e+11p ps=2.62e+06u
M1003 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_117_297# D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1005 a_317_297# B a_221_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__clkinvlp_2 VNB VPWR VGND VPB Y A
M1000 Y A a_150_67# VNB nshort w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=1.98e+11p ps=1.82e+06u
M1001 VPWR A Y VPB phighvt w=1e+06u l=250000u
+  ad=6.5e+11p pd=5.3e+06u as=2.8e+11p ps=2.56e+06u
M1002 a_150_67# A VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1003 Y A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__einvp_8 A Z TE VPWR VGND VPB VNB
M1000 Z A a_235_309# VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=2.5515e+12p ps=2.277e+07u
M1001 a_213_47# TE VGND VNB nshort w=650000u l=150000u
+  ad=1.885e+12p pd=1.75e+07u as=1.014e+12p ps=9.62e+06u
M1002 a_213_47# TE VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR a_27_47# a_235_309# VPB phighvt w=940000u l=180000u
+  ad=1.3604e+12p pd=1.238e+07u as=0p ps=0u
M1004 Z A a_235_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_235_309# A Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_27_47# a_235_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Z A a_213_47# VNB nshort w=650000u l=150000u
+  ad=8.32e+11p pd=7.76e+06u as=0p ps=0u
M1008 a_213_47# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_235_309# a_27_47# VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND TE a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Z A a_235_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_213_47# TE VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR TE a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1014 VPWR a_27_47# a_235_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_235_309# A Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND TE a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Z A a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_235_309# a_27_47# VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_213_47# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Z A a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Z A a_235_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND TE a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_213_47# TE VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_235_309# A Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND TE a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_213_47# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR a_27_47# a_235_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Z A a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_235_309# a_27_47# VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_235_309# A Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND TE a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1032 a_213_47# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_235_309# a_27_47# VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and2_4 X B A VNB VPB VGND VPWR
M1000 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6e+11p pd=5.2e+06u as=1.245e+12p ps=1.049e+07u
M1001 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=7.085e+11p pd=6.08e+06u as=4.615e+11p ps=4.02e+06u
M1002 a_120_47# A a_27_47# VNB nshort w=650000u l=150000u
+  ad=1.365e+11p pd=1.72e+06u as=2.0475e+11p ps=1.93e+06u
M1003 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_47# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1005 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B a_120_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__dfrtp_1 RESET_B VGND VPWR Q D CLK VPB VNB
M1000 a_436_413# D VPWR VPB phighvt w=420000u l=180000u
+  ad=1.428e+11p pd=1.52e+06u as=1.3145e+12p ps=1.289e+07u
M1001 VPWR a_1323_21# a_1330_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=9.66e+10p ps=1.3e+06u
M1002 a_211_363# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.1789e+12p ps=1.006e+07u
M1003 Q a_1323_21# VGND VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=0p ps=0u
M1004 a_649_413# a_27_47# a_534_47# VPB phighvt w=420000u l=180000u
+  ad=3.318e+11p pd=3.26e+06u as=1.533e+11p ps=1.57e+06u
M1005 a_805_47# a_751_289# a_642_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.748e+11p ps=2.17e+06u
M1006 VPWR CLK a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1007 VGND RESET_B a_805_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_436_413# D VGND VNB nshort w=420000u l=150000u
+  ad=1.338e+11p pd=1.5e+06u as=0p ps=0u
M1009 VGND a_1323_21# a_1237_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.698e+11p ps=1.7e+06u
M1010 VPWR a_751_289# a_649_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_751_289# a_534_47# VGND VNB nshort w=640000u l=150000u
+  ad=1.998e+11p pd=1.97e+06u as=0p ps=0u
M1012 Q a_1323_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=0p ps=0u
M1013 VPWR a_1128_47# a_1323_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1014 a_1128_47# a_211_363# a_751_289# VNB nshort w=360000u l=150000u
+  ad=1.422e+11p pd=1.51e+06u as=0p ps=0u
M1015 a_534_47# a_27_47# a_436_413# VNB nshort w=360000u l=150000u
+  ad=1.404e+11p pd=1.5e+06u as=0p ps=0u
M1016 a_751_289# a_534_47# VPWR VPB phighvt w=840000u l=180000u
+  ad=2.709e+11p pd=2.41e+06u as=0p ps=0u
M1017 a_1128_47# a_27_47# a_751_289# VPB phighvt w=420000u l=180000u
+  ad=1.512e+11p pd=1.56e+06u as=0p ps=0u
M1018 a_642_47# a_211_363# a_534_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1237_47# a_27_47# a_1128_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1542_47# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=1.596e+11p pd=1.6e+06u as=0p ps=0u
M1021 a_1323_21# a_1128_47# a_1542_47# VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1022 a_649_413# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1024 a_1323_21# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_211_363# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1026 a_534_47# a_211_363# a_436_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1330_413# a_211_363# a_1128_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sdlclkp_1 CLK VGND VPWR SCE GCLK GATE VPB VNB
M1000 a_484_315# a_299_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=1.3826e+12p ps=1.216e+07u
M1001 a_1089_47# a_484_315# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.92e+11p pd=1.88e+06u as=0p ps=0u
M1002 a_269_21# CLK VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1003 a_27_47# GATE a_117_369# VPB phighvt w=640000u l=180000u
+  ad=2.021e+11p pd=1.97e+06u as=1.472e+11p ps=1.74e+06u
M1004 a_484_315# a_299_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=7.9265e+11p ps=7.37e+06u
M1005 a_117_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_415_47# a_266_243# a_299_47# VNB nshort w=360000u l=150000u
+  ad=1.968e+11p pd=1.85e+06u as=1.548e+11p ps=1.58e+06u
M1007 a_269_21# CLK VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1008 a_1181_47# a_484_315# a_1089_47# VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=1.302e+11p ps=1.46e+06u
M1009 a_410_413# a_269_21# a_299_47# VPB phighvt w=420000u l=180000u
+  ad=1.596e+11p pd=1.6e+06u as=1.47e+11p ps=1.54e+06u
M1010 VPWR a_484_315# a_410_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_484_315# a_415_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 GCLK a_1089_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1013 VGND CLK a_1181_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_299_47# a_269_21# a_27_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=2.622e+11p ps=2.95e+06u
M1015 VGND SCE a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR CLK a_1089_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_299_47# a_266_243# a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 GCLK a_1089_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.8525e+11p pd=1.87e+06u as=0p ps=0u
M1019 VGND a_269_21# a_266_243# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1020 VPWR a_269_21# a_266_243# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1021 a_27_47# GATE VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a32oi_4 A3 A2 A1 B1 Y B2 VNB VPB VGND VPWR
M1000 a_27_297# B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=3.925e+12p pd=2.985e+07u as=1.16e+12p ps=1.032e+07u
M1001 a_27_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_27_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=9.62e+11p pd=9.46e+06u as=9.75e+11p ps=9.5e+06u
M1003 a_893_47# A2 a_1379_47# VNB nshort w=650000u l=150000u
+  ad=1.053e+12p pd=9.74e+06u as=8.97e+11p ps=7.96e+06u
M1004 Y B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.195e+12p ps=1.639e+07u
M1006 VPWR A3 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_893_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=8.645e+11p ps=7.86e+06u
M1008 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_297# B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A1 a_893_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1379_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1379_47# A2 a_893_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_893_47# A2 a_1379_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_27_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A3 a_1379_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_297# A3 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_27_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR A3 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_27_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_893_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_27_297# A3 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Y A1 a_893_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 Y B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1379_47# A2 a_893_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1379_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND A3 a_1379_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and4_1 X C A B D VGND VPWR VPB VNB
M1000 VGND D a_299_47# VNB nshort w=420000u l=150000u
+  ad=2.7525e+11p pd=2.2e+06u as=1.428e+11p ps=1.52e+06u
M1001 a_27_47# A VPWR VPB phighvt w=420000u l=180000u
+  ad=2.52e+11p pd=2.88e+06u as=5.601e+11p ps=5.56e+06u
M1002 a_203_47# B a_119_47# VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=1.134e+11p ps=1.38e+06u
M1003 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=4.6e+11p pd=2.92e+06u as=0p ps=0u
M1004 a_27_47# C VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=2.925e+11p pd=2.2e+06u as=0p ps=0u
M1006 a_299_47# C a_203_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_119_47# A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1008 VPWR B a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR D a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand2_4 Y A B VPB VNB VGND VPWR
M1000 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=1.41e+12p pd=1.282e+07u as=1.16e+12p ps=1.032e+07u
M1001 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=9.62e+11p pd=9.46e+06u as=4.16e+11p ps=3.88e+06u
M1003 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.485e+11p ps=3.98e+06u
M1006 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a21bo_4 B1_N A2 A1 X VNB VPB VGND VPWR
M1000 X a_209_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6e+11p pd=5.2e+06u as=1.47e+12p ps=1.294e+07u
M1001 X a_209_21# VGND VNB nshort w=650000u l=150000u
+  ad=4.29e+11p pd=3.92e+06u as=1.4235e+12p ps=1.088e+07u
M1002 VPWR A2 a_647_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.12e+12p ps=1.024e+07u
M1003 VPWR B1_N a_36_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.75e+11p ps=2.55e+06u
M1004 VGND a_209_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_647_297# a_36_47# a_209_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1006 VPWR a_209_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_209_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_647_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_209_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_36_47# a_209_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.485e+11p ps=3.98e+06u
M1011 a_1115_47# A1 a_209_21# VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1012 VPWR a_209_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND B1_N a_36_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.8275e+11p ps=2.17e+06u
M1014 VPWR A1 a_647_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A2 a_1115_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_209_21# a_36_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_935_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=1.495e+11p pd=1.76e+06u as=0p ps=0u
M1018 X a_209_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_209_21# a_36_47# a_647_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_647_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_209_21# A1 a_935_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o21a_2 A1 B1 A2 X VNB VPB VGND VPWR
M1000 a_79_21# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=1.365e+12p ps=8.73e+06u
M1001 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1002 a_414_47# B1 a_79_21# VNB nshort w=650000u l=150000u
+  ad=3.8675e+11p pd=3.79e+06u as=2.0475e+11p ps=1.93e+06u
M1003 a_414_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.1825e+11p ps=6.11e+06u
M1004 VGND A2 a_414_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=2.1125e+11p pd=1.95e+06u as=0p ps=0u
M1006 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_508_297# A2 a_79_21# VPB phighvt w=1e+06u l=180000u
+  ad=5e+11p pd=3e+06u as=0p ps=0u
M1008 VPWR A1 a_508_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a31oi_4 Y B1 A2 A3 A1 VNB VPB VPWR VGND
M1000 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.2e+12p pd=2.44e+07u as=1.74e+12p ps=1.548e+07u
M1001 a_27_297# A3 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_27_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=9.62e+11p pd=9.46e+06u as=8.32e+11p ps=7.76e+06u
M1003 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_297# B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1006 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=1.0335e+12p pd=9.68e+06u as=0p ps=0u
M1007 Y A1 a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=8.645e+11p ps=7.86e+06u
M1008 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_47# A2 a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A3 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_485_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_297# B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_485_47# A2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_27_297# A3 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A3 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_27_47# A2 a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y A1 a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_485_47# A2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_485_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A3 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND A3 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__mux2i_4 S A1 A0 Y VNB VPB VGND VPWR
M1000 Y A1 a_493_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.41e+12p pd=1.282e+07u as=1.215e+12p ps=1.043e+07u
M1001 VGND a_1311_21# a_109_47# VNB nshort w=650000u l=150000u
+  ad=1.03025e+12p pd=9.67e+06u as=9.3275e+11p ps=8.07e+06u
M1002 Y A0 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.16e+12p ps=1.032e+07u
M1003 VPWR a_1311_21# a_493_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.475e+12p pd=1.295e+07u as=0p ps=0u
M1004 a_109_47# a_1311_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_117_297# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND S a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=8.645e+11p ps=7.86e+06u
M1007 a_493_297# A1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_485_47# S VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR S a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_109_47# A0 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=9.295e+11p ps=9.36e+06u
M1011 Y A1 a_493_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A0 a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A1 a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_493_297# a_1311_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_117_297# A0 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND S a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_493_297# A1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_1311_21# a_493_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_485_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_117_297# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_109_47# a_1311_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y A0 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_493_297# a_1311_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_485_47# S VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y A0 a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y A1 a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_485_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND a_1311_21# a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1311_21# S VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1030 a_117_297# A0 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR S a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_109_47# A0 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1311_21# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand4_1 C B Y D A VPB VNB VPWR VGND
M1000 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=8.7e+11p pd=7.74e+06u as=6.4e+11p ps=5.28e+06u
M1001 a_213_47# C a_119_47# VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=2.08e+11p ps=1.94e+06u
M1002 Y A a_297_47# VNB nshort w=650000u l=150000u
+  ad=2.275e+11p pd=2e+06u as=2.47e+11p ps=2.06e+06u
M1003 a_297_47# B a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_119_47# D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1007 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and3b_1 A_N B X C VGND VPWR VPB VNB
M1000 a_317_53# a_117_413# a_225_311# VNB nshort w=420000u l=150000u
+  ad=1.344e+11p pd=1.48e+06u as=1.197e+11p ps=1.41e+06u
M1001 X a_225_311# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=4.7045e+11p ps=4.01e+06u
M1002 a_117_413# A_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=5.913e+11p ps=5.75e+06u
M1003 a_225_311# B VPWR VPB phighvt w=420000u l=180000u
+  ad=2.7055e+11p pd=3.05e+06u as=0p ps=0u
M1004 VPWR C a_225_311# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_117_413# a_225_311# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_117_413# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1007 a_411_53# B a_317_53# VNB nshort w=420000u l=150000u
+  ad=1.071e+11p pd=1.35e+06u as=0p ps=0u
M1008 X a_225_311# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1009 VGND C a_411_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__ebufn_8 A Z TE_B VNB VPB VGND VPWR
M1000 VPWR TE_B a_437_309# VPB phighvt w=940000u l=180000u
+  ad=1.9584e+12p pd=1.56e+07u as=3.2075e+12p ps=2.41e+07u
M1001 VPWR TE_B a_437_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_437_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_437_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_485_47# a_124_297# Z VNB nshort w=650000u l=150000u
+  ad=2.106e+12p pd=1.818e+07u as=8.645e+11p ps=7.86e+06u
M1005 VPWR A a_124_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1006 a_437_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_321_47# TE_B VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=1.417e+12p ps=1.216e+07u
M1008 a_437_309# a_124_297# Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.16e+12p ps=1.032e+07u
M1009 a_485_47# a_321_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_485_47# a_321_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_485_47# a_124_297# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR TE_B a_437_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_124_297# A VGND VNB nshort w=650000u l=150000u
+  ad=2.08e+11p pd=1.94e+06u as=0p ps=0u
M1014 a_321_47# TE_B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1015 Z a_124_297# a_437_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR TE_B a_437_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Z a_124_297# a_437_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_321_47# a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_485_47# a_321_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_437_309# a_124_297# Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_437_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_321_47# a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Z a_124_297# a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Z a_124_297# a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_485_47# a_124_297# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND A a_124_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_485_47# a_124_297# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_437_309# a_124_297# Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Z a_124_297# a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_437_309# a_124_297# Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Z a_124_297# a_437_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND a_321_47# a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_124_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND a_321_47# a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 Z a_124_297# a_437_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_485_47# a_321_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 Z a_124_297# a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor2_2 B Y A VPB VNB VGND VPWR
M1000 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=8.5e+11p ps=7.7e+06u
M1001 a_27_297# B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1002 Y B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A VGND VNB nshort w=650000u l=150000u
+  ad=4.81e+11p pd=4.08e+06u as=6.0125e+11p ps=5.75e+06u
M1004 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__dlrtn_4 RESET_B D GATE_N Q VGND VPWR VPB VNB
M1000 Q a_750_21# VGND VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=1.00625e+12p ps=1.01e+07u
M1001 VGND a_750_21# a_708_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1002 Q a_750_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=1.691e+12p ps=1.487e+07u
M1003 VPWR GATE_N a_27_363# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1004 VPWR a_750_21# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_203_47# a_27_363# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1006 VPWR a_750_21# a_702_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1007 VGND a_750_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_503_369# a_319_369# VPWR VPB phighvt w=640000u l=180000u
+  ad=2.021e+11p pd=1.97e+06u as=0p ps=0u
M1009 a_708_47# a_203_47# a_604_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.58e+06u
M1010 Q a_750_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Q a_750_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND D a_319_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1013 VPWR D a_319_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1014 VGND RESET_B a_981_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.6575e+11p ps=1.81e+06u
M1015 a_604_47# a_27_363# a_500_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.58e+06u
M1016 VPWR RESET_B a_750_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1017 a_981_47# a_604_47# a_750_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1018 VGND GATE_N a_27_363# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1019 a_702_413# a_27_363# a_604_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1020 a_203_47# a_27_363# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1021 a_604_47# a_203_47# a_503_369# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_750_21# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_500_47# a_319_369# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_750_21# a_604_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_750_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand4b_2 D C B Y A_N VNB VPB VGND VPWR
M1000 VPWR A_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=2.2234e+12p pd=1.56e+07u as=1.134e+11p ps=1.38e+06u
M1001 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.16e+12p ps=1.032e+07u
M1002 a_705_47# D VGND VNB nshort w=650000u l=150000u
+  ad=6.37e+11p pd=5.86e+06u as=3.172e+11p ps=3.3e+06u
M1003 VPWR D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_225_47# a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=5.785e+11p pd=5.68e+06u as=2.08e+11p ps=1.94e+06u
M1005 a_705_47# C a_495_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1006 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND D a_705_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_225_47# B a_495_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_495_47# B a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1012 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y a_27_47# a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_495_47# C a_705_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or2b_4 A B_N X VNB VPB VGND VPWR
M1000 VGND B_N a_27_53# VNB nshort w=420000u l=150000u
+  ad=1.11205e+12p pd=8.88e+06u as=1.302e+11p ps=1.46e+06u
M1001 a_27_53# B_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=1.0684e+12p ps=9.29e+06u
M1002 VPWR a_229_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1003 VGND A a_229_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1004 a_229_297# a_27_53# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_319_297# a_27_53# a_229_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.3e+11p pd=2.46e+06u as=2.7e+11p ps=2.54e+06u
M1006 X a_229_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_319_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_229_297# VGND VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=0p ps=0u
M1009 VGND a_229_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_229_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_229_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_229_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_229_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__xnor2_1 VGND VPWR B Y A VPB VNB
M1000 Y B a_415_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.5e+11p pd=2.7e+06u as=2.3e+11p ps=2.46e+06u
M1001 a_415_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.48e+12p ps=8.96e+06u
M1002 a_139_47# B a_47_47# VNB nshort w=650000u l=150000u
+  ad=1.365e+11p pd=1.72e+06u as=2.015e+11p ps=1.92e+06u
M1003 VPWR A a_47_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1004 a_315_47# A VGND VNB nshort w=650000u l=150000u
+  ad=3.77e+11p pd=3.76e+06u as=4.42e+11p ps=3.96e+06u
M1005 Y a_47_47# a_315_47# VNB nshort w=650000u l=150000u
+  ad=1.95e+11p pd=1.9e+06u as=0p ps=0u
M1006 a_315_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A a_139_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_47_47# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_47_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a21o_6 A2 A1 X B1 VNB VPB VGND VPWR
M1000 VGND A2 a_297_47# VNB nshort w=650000u l=150000u
+  ad=1.69e+12p pd=1.3e+07u as=1.69e+11p ps=1.82e+06u
M1001 X a_213_47# VGND VNB nshort w=650000u l=150000u
+  ad=5.265e+11p pd=5.52e+06u as=0p ps=0u
M1002 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.12e+12p pd=1.024e+07u as=1.7e+12p ps=1.54e+07u
M1003 a_213_47# A1 a_131_47# VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=1.69e+11p ps=1.82e+06u
M1004 X a_213_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.7e+11p pd=7.74e+06u as=0p ps=0u
M1005 X a_213_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_213_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_297_47# A1 a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_297# B1 a_213_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1009 VGND a_213_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_213_47# B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_131_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_213_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_213_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_213_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_213_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_213_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND B1 a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_213_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_213_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_213_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a2bb2oi_4 Y A2_N B2 A1_N B1 VNB VPB VGND VPWR
M1000 a_27_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.99e+12p pd=1.798e+07u as=1.74e+12p ps=1.548e+07u
M1001 VGND A1_N a_831_21# VNB nshort w=650000u l=150000u
+  ad=2.067e+12p pd=1.806e+07u as=8.97e+11p ps=7.96e+06u
M1002 a_27_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_831_21# A1_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_297# a_831_21# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1005 VPWR B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_831_21# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=8.97e+11p ps=7.96e+06u
M1007 a_831_21# A2_N a_1259_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=1.43e+12p ps=1.286e+07u
M1008 Y a_831_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_831_21# a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_297# B2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B1 a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.995e+11p ps=7.66e+06u
M1012 VGND B1 a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A1_N a_1259_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_109_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_831_21# A2_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1259_297# A2_N a_831_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_831_21# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A1_N a_831_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1259_297# A1_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_831_21# A2_N a_1259_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_297# a_831_21# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_831_21# A1_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A2_N a_831_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_27_297# B2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR A1_N a_1259_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1259_297# A1_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y a_831_21# a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y B2 a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_109_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_109_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Y B2 a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 Y a_831_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1259_297# A2_N a_831_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_831_21# A2_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_109_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND A2_N a_831_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__bufinv_16 A Y VNB VPB VGND VPWR
M1000 a_391_47# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.7e+11p pd=7.74e+06u as=3.75e+12p ps=3.35e+07u
M1001 a_27_47# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
M1002 Y a_391_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.32e+12p pd=2.064e+07u as=0p ps=0u
M1003 Y a_391_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_391_47# Y VNB nshort w=650000u l=150000u
+  ad=2.6e+12p pd=2.49e+07u as=1.6965e+12p ps=1.562e+07u
M1005 VPWR a_27_47# a_391_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_391_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_391_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y a_391_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_391_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y a_391_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_391_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_391_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_391_47# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_47# A VGND VNB nshort w=650000u l=150000u
+  ad=4.095e+11p pd=3.86e+06u as=0p ps=0u
M1015 VPWR a_391_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y a_391_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_391_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y a_391_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y a_391_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_391_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=6.565e+11p pd=5.92e+06u as=0p ps=0u
M1022 Y a_391_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_27_47# a_391_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_27_47# a_391_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_391_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_391_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y a_391_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y a_391_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y a_391_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_391_47# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND a_391_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Y a_391_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR a_391_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Y a_391_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR a_27_47# a_391_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_391_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 Y a_391_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 Y a_391_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR a_391_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND a_27_47# a_391_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPWR A a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_391_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VGND a_391_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VGND a_391_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 VPWR a_391_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VPWR a_391_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1048 VGND a_27_47# a_391_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or4b_1 B D_N A X C VPWR VGND VPB VNB
M1000 a_117_297# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=6.1845e+11p ps=6.42e+06u
M1001 a_225_297# a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=2.961e+11p pd=3.09e+06u as=0p ps=0u
M1002 X a_225_297# VGND VNB nshort w=650000u l=150000u
+  ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u
M1003 VGND A a_225_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_117_297# D_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=4.241e+11p ps=4.1e+06u
M1005 a_504_297# B a_416_297# VPB phighvt w=420000u l=180000u
+  ad=1.344e+11p pd=1.48e+06u as=1.092e+11p ps=1.36e+06u
M1006 a_225_297# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_504_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND C a_225_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_315_297# a_117_297# a_225_297# VPB phighvt w=420000u l=180000u
+  ad=1.365e+11p pd=1.49e+06u as=1.134e+11p ps=1.38e+06u
M1010 a_416_297# C a_315_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_225_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o2bb2ai_2 B2 Y A1_N A2_N B1 VNB VPB VGND VPWR
M1000 a_121_297# A1_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=1.96e+12p ps=1.392e+07u
M1001 a_121_297# A2_N a_123_47# VNB nshort w=650000u l=150000u
+  ad=2.405e+11p pd=2.04e+06u as=3.575e+11p ps=3.7e+06u
M1002 a_503_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=8.7425e+11p pd=7.89e+06u as=7.345e+11p ps=7.46e+06u
M1003 VPWR A1_N a_121_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A1_N a_123_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_788_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=5.8e+11p ps=5.16e+06u
M1006 a_123_47# A1_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_121_297# A2_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B2 a_788_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_121_297# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_503_47# a_121_297# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1011 a_123_47# A2_N a_121_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y a_121_297# a_503_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_503_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_788_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A2_N a_121_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y a_121_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND B2 a_503_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND B1 a_503_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR B1 a_788_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a2bb2o_1 VNB VPB VGND VPWR B1 A1_N A2_N X B2
M1000 a_525_413# a_243_47# a_79_21# VPB phighvt w=420000u l=180000u
+  ad=2.352e+11p pd=2.8e+06u as=1.134e+11p ps=1.38e+06u
M1001 a_611_47# B2 a_79_21# VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=1.134e+11p ps=1.38e+06u
M1002 a_79_21# a_243_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=7.746e+11p ps=6.34e+06u
M1003 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=4.674e+11p pd=4.32e+06u as=2.7e+11p ps=2.54e+06u
M1004 a_241_297# A1_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.029e+11p pd=1.33e+06u as=0p ps=0u
M1005 a_525_413# B1 VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2_N a_243_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1007 VGND B1 a_611_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_243_47# A1_N VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_243_47# A2_N a_241_297# VPB phighvt w=420000u l=180000u
+  ad=1.155e+11p pd=1.39e+06u as=0p ps=0u
M1010 VPWR B2 a_525_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
.ends
.subckt sky130_fd_sc_hdll__xor3_1 X C B A VNB VPB VGND VPWR
M1000 VGND A a_991_365# VNB nshort w=640000u l=150000u
+  ad=9.7095e+11p pd=6.94e+06u as=4.498e+11p ps=3.99e+06u
M1001 a_276_93# C VPWR VPB phighvt w=640000u l=180000u
+  ad=1.856e+11p pd=1.86e+06u as=1.3094e+12p ps=8.68e+06u
M1002 a_276_93# C VGND VNB nshort w=420000u l=150000u
+  ad=1.974e+11p pd=1.78e+06u as=0p ps=0u
M1003 a_875_297# B VGND VNB nshort w=650000u l=150000u
+  ad=1.653e+11p pd=1.82e+06u as=0p ps=0u
M1004 a_424_49# B a_991_365# VNB nshort w=640000u l=150000u
+  ad=5.931e+11p pd=4.52e+06u as=0p ps=0u
M1005 a_116_21# C a_406_325# VPB phighvt w=840000u l=180000u
+  ad=3.36e+11p pd=2.48e+06u as=7.824e+11p ps=5.28e+06u
M1006 a_875_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.126e+11p pd=2.64e+06u as=0p ps=0u
M1007 a_116_21# C a_424_49# VNB nshort w=640000u l=150000u
+  ad=2.88e+11p pd=2.18e+06u as=0p ps=0u
M1008 a_1276_297# a_875_297# a_424_49# VNB nshort w=420000u l=150000u
+  ad=5.677e+11p pd=4.42e+06u as=0p ps=0u
M1009 a_406_325# B a_1276_297# VNB nshort w=640000u l=150000u
+  ad=6.5745e+11p pd=4.66e+06u as=0p ps=0u
M1010 a_991_365# a_875_297# a_424_49# VPB phighvt w=840000u l=180000u
+  ad=7.234e+11p pd=5.3e+06u as=7.558e+11p ps=5.2e+06u
M1011 a_406_325# B a_991_365# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_424_49# B a_1276_297# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=7.998e+11p ps=5.68e+06u
M1013 a_1276_297# a_991_365# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_991_365# a_875_297# a_406_325# VNB nshort w=600000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1276_297# a_875_297# a_406_325# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A a_991_365# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_424_49# a_276_93# a_116_21# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_116_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.82e+11p ps=1.86e+06u
M1019 VPWR a_116_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1020 a_406_325# a_276_93# a_116_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1276_297# a_991_365# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__dlrtp_1 RESET_B D GATE Q VGND VPWR VPB VNB
M1000 VGND a_750_21# a_708_47# VNB nshort w=420000u l=150000u
+  ad=5.6425e+11p pd=6.14e+06u as=8.82e+10p ps=1.26e+06u
M1001 VPWR GATE a_27_363# VPB phighvt w=640000u l=180000u
+  ad=1.131e+12p pd=9.75e+06u as=1.728e+11p ps=1.82e+06u
M1002 a_203_47# a_27_363# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1003 VPWR a_750_21# a_702_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1004 a_503_369# a_319_369# VPWR VPB phighvt w=640000u l=180000u
+  ad=2.021e+11p pd=1.97e+06u as=0p ps=0u
M1005 a_708_47# a_27_363# a_604_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.58e+06u
M1006 Q a_750_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1007 VGND D a_319_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1008 VPWR D a_319_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1009 VGND RESET_B a_981_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.6575e+11p ps=1.81e+06u
M1010 a_604_47# a_203_47# a_500_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.58e+06u
M1011 Q a_750_21# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1012 VPWR RESET_B a_750_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1013 a_981_47# a_604_47# a_750_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1014 VGND GATE a_27_363# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1015 a_702_413# a_203_47# a_604_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1016 a_203_47# a_27_363# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1017 a_604_47# a_27_363# a_503_369# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_500_47# a_319_369# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_750_21# a_604_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor2b_4 B_N Y A VNB VPB VGND VPWR
M1000 Y a_459_21# a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=1.45e+12p ps=1.29e+07u
M1001 VGND a_459_21# Y VNB nshort w=650000u l=150000u
+  ad=1.183e+12p pd=1.144e+07u as=8.645e+11p ps=7.86e+06u
M1002 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=8.7e+11p pd=7.74e+06u as=0p ps=0u
M1003 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y a_459_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_459_21# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_297# a_459_21# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR B_N a_459_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1012 VGND B_N a_459_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.82e+11p ps=1.86e+06u
M1013 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y a_459_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y a_459_21# a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_297# a_459_21# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__buf_1 VGND VPWR X A VPB VNB
M1000 VPWR A a_27_47# VPB phighvt w=790000u l=180000u
+  ad=2.449e+11p pd=2.2e+06u as=2.133e+11p ps=2.12e+06u
M1001 X a_27_47# VPWR VPB phighvt w=790000u l=180000u
+  ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 VGND A a_27_47# VNB nshort w=520000u l=150000u
+  ad=1.768e+11p pd=1.72e+06u as=1.612e+11p ps=1.66e+06u
M1003 X a_27_47# VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__inv_1 Y A VPB VNB VGND VPWR
M1000 Y A VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=2.015e+11p ps=1.92e+06u
M1001 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=2.7e+11p ps=2.54e+06u
.ends
.subckt sky130_fd_sc_hdll__and2_2 VPWR VGND A X B VPB VNB
M1000 X a_27_75# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=4.1e+11p pd=2.82e+06u as=8.191e+11p ps=6.94e+06u
M1001 X a_27_75# VGND VNB nshort w=650000u l=150000u
+  ad=3.185e+11p pd=2.28e+06u as=4.656e+11p ps=4.16e+06u
M1002 a_27_75# A VPWR VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
M1003 VGND a_27_75# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND B a_123_75# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1005 VPWR a_27_75# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR B a_27_75# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_123_75# A a_27_75# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
.ends
.subckt sky130_fd_sc_hdll__nor4b_1 C B A D_N Y VPB VNB VGND VPWR
M1000 a_263_297# C a_169_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.5e+11p pd=2.7e+06u as=2.9e+11p ps=2.58e+06u
M1001 a_169_297# a_91_199# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.3e+11p ps=3.06e+06u
M1002 a_91_199# D_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=4.799e+11p ps=3.07e+06u
M1003 Y B VGND VNB nshort w=650000u l=150000u
+  ad=3.835e+11p pd=3.78e+06u as=8.046e+11p ps=6.45e+06u
M1004 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A a_369_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1006 Y a_91_199# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_91_199# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1009 a_369_297# B a_263_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a211oi_1 A1 C1 B1 Y A2 VPWR VGND VPB VNB
M1000 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.05e+11p pd=2.61e+06u as=6.45e+11p ps=5.29e+06u
M1001 Y C1 a_325_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.6e+11p pd=2.72e+06u as=3.15e+11p ps=2.63e+06u
M1002 a_123_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=1.8525e+11p pd=1.87e+06u as=4.3875e+11p ps=3.95e+06u
M1003 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=5.1025e+11p ps=4.17e+06u
M1005 a_325_297# B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A1 a_123_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y C1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sedfxbp_2 VPWR VGND CLK Q_N SCD DE D Q SCE VPB VNB
M1000 a_1787_159# a_1611_413# VPWR VPB phighvt w=750000u l=180000u
+  ad=2.025e+11p pd=2.04e+06u as=2.49535e+12p ps=2.217e+07u
M1001 a_211_363# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.7892e+12p ps=1.767e+07u
M1002 a_2165_413# a_1787_159# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.365e+11p pd=1.49e+06u as=0p ps=0u
M1003 a_2266_413# a_27_47# a_2165_413# VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
M1004 VGND a_851_264# a_2414_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.32e+11p ps=1.49e+06u
M1005 VPWR a_2266_413# a_851_264# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1006 VPWR DE a_455_324# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1007 VPWR CLK a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1008 VPWR a_2266_413# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1009 a_319_47# a_851_264# a_779_47# VNB nshort w=420000u l=150000u
+  ad=2.478e+11p pd=2.86e+06u as=1.932e+11p ps=1.76e+06u
M1010 a_2181_47# a_1787_159# VGND VNB nshort w=420000u l=150000u
+  ad=1.356e+11p pd=1.51e+06u as=0p ps=0u
M1011 VPWR a_851_264# Q_N VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1012 a_2266_413# a_211_363# a_2181_47# VNB nshort w=360000u l=150000u
+  ad=1.908e+11p pd=1.78e+06u as=0p ps=0u
M1013 a_1611_413# a_27_47# a_985_47# VNB nshort w=360000u l=150000u
+  ad=1.404e+11p pd=1.5e+06u as=6.015e+11p ps=4.57e+06u
M1014 a_985_47# a_955_21# a_1376_369# VPB phighvt w=640000u l=180000u
+  ad=4.837e+11p pd=4.13e+06u as=2.24e+11p ps=1.98e+06u
M1015 VGND SCE a_955_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1016 Q a_2266_413# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_851_264# Q_N VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1018 VGND a_2266_413# a_851_264# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1019 a_985_47# a_955_21# a_319_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Q_N a_851_264# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_2414_47# a_27_47# a_2266_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR SCE a_955_21# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.76e+11p ps=1.83e+06u
M1023 a_409_369# D a_319_47# VPB phighvt w=640000u l=180000u
+  ad=1.472e+11p pd=1.74e+06u as=3.84e+11p ps=3.76e+06u
M1024 a_985_47# SCE a_1373_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1025 a_787_369# DE VPWR VPB phighvt w=640000u l=180000u
+  ad=2.432e+11p pd=2.04e+06u as=0p ps=0u
M1026 a_319_47# a_851_264# a_787_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1611_413# a_211_363# a_985_47# VPB phighvt w=420000u l=180000u
+  ad=1.365e+11p pd=1.49e+06u as=0p ps=0u
M1028 VPWR a_1787_159# a_1712_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.617e+11p ps=1.61e+06u
M1029 VPWR a_455_324# a_409_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_985_47# SCE a_319_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND a_2266_413# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.405e+11p ps=2.04e+06u
M1032 a_1712_413# a_27_47# a_1611_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Q_N a_851_264# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND DE a_455_324# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1035 a_779_47# a_455_324# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1376_369# SCD VPWR VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1038 a_1373_119# SCD VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR a_851_264# a_2360_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=2.058e+11p ps=1.82e+06u
M1040 VGND a_1787_159# a_1738_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.518e+11p ps=1.6e+06u
M1041 a_211_363# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1042 a_1738_47# a_211_363# a_1611_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_413_47# D a_319_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1044 Q a_2266_413# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VGND DE a_413_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_2360_413# a_211_363# a_2266_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_1787_159# a_1611_413# VGND VNB nshort w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a32oi_2 A2 B2 A3 A1 Y B1 VNB VPB VGND VPWR
M1000 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.08e+12p pd=1.016e+07u as=1.71e+12p ps=1.542e+07u
M1001 a_27_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1002 a_27_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=5.46e+11p pd=5.58e+06u as=6.4675e+11p ps=5.89e+06u
M1003 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=4.16e+11p pd=3.88e+06u as=0p ps=0u
M1005 a_27_297# A3 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A3 a_757_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.81e+11p ps=4.08e+06u
M1007 Y B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_507_47# A2 a_757_47# VNB nshort w=650000u l=150000u
+  ad=5.135e+11p pd=5.48e+06u as=0p ps=0u
M1009 VPWR A3 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_507_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A1 a_507_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_297# B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_757_47# A2 a_507_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_757_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and4b_4 X D C B A_N VNB VPB VGND VPWR
M1000 a_184_21# a_27_47# a_814_47# VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=2.47e+11p ps=2.06e+06u
M1001 a_718_47# C a_624_47# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u
M1002 a_624_47# D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.205e+11p ps=6.17e+06u
M1003 VPWR A_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=1.6157e+12p pd=1.333e+07u as=1.134e+11p ps=1.38e+06u
M1004 a_184_21# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6.4e+11p pd=5.28e+06u as=0p ps=0u
M1005 a_814_47# B a_718_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_184_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1007 X a_184_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_184_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1009 VPWR C a_184_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_184_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_184_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_27_47# a_184_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1014 VGND a_184_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_184_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_184_21# D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_184_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand2_2 Y A B VPB VNB VGND VPWR
M1000 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=8.3e+11p pd=7.66e+06u as=5.8e+11p ps=5.16e+06u
M1001 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=5.135e+11p pd=5.48e+06u as=2.405e+11p ps=2.04e+06u
M1002 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=2.405e+11p pd=2.04e+06u as=0p ps=0u
M1003 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a31o_4 B1 A2 A3 A1 X VNB VPB VGND VPWR
M1000 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.47e+12p pd=1.294e+07u as=1.76e+12p ps=1.552e+07u
M1001 a_213_47# A2 a_119_47# VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=2.08e+11p ps=1.94e+06u
M1002 a_27_297# A3 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_297_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1004 VGND a_297_47# X VNB nshort w=650000u l=150000u
+  ad=1.404e+12p pd=1.082e+07u as=4.16e+11p ps=3.88e+06u
M1005 a_297_47# A1 a_213_47# VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=0p ps=0u
M1006 VPWR a_297_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A3 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_297_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_297# B1 a_297_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1010 VGND a_297_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND B1 a_297_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_297_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_495_47# A2 a_401_47# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u
M1015 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_119_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_401_47# A1 a_297_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_297_47# B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A3 a_495_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_297_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_297_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_297_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__xnor3_4 X B C A VNB VPB VGND VPWR
M1000 X a_101_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=1.50095e+12p ps=1.307e+07u
M1001 a_1490_297# a_1207_297# VGND VNB nshort w=640000u l=150000u
+  ad=5.677e+11p pd=4.42e+06u as=1.0748e+12p ps=9.85e+06u
M1002 a_532_93# C VPWR VPB phighvt w=640000u l=180000u
+  ad=1.856e+11p pd=1.86e+06u as=0p ps=0u
M1003 VGND A a_1207_297# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=4.44e+11p ps=3.96e+06u
M1004 a_1089_297# B VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=0p ps=0u
M1005 VGND a_101_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1006 a_657_325# B a_1207_297# VNB nshort w=640000u l=150000u
+  ad=5.835e+11p pd=4.49e+06u as=0p ps=0u
M1007 VGND a_101_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_681_49# B a_1207_297# VPB phighvt w=840000u l=180000u
+  ad=8.3175e+11p pd=5.4e+06u as=7.226e+11p ps=5.29e+06u
M1009 X a_101_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1207_297# a_1089_297# a_657_325# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=5.878e+11p ps=4.8e+06u
M1011 a_1490_297# a_1089_297# a_657_325# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_101_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1490_297# a_1207_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=7.998e+11p pd=5.68e+06u as=0p ps=0u
M1014 a_681_49# B a_1490_297# VNB nshort w=640000u l=150000u
+  ad=5.4845e+11p pd=4.32e+06u as=0p ps=0u
M1015 a_1207_297# a_1089_297# a_681_49# VNB nshort w=600000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_657_325# B a_1490_297# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_101_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A a_1207_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_101_21# C a_657_325# VPB phighvt w=840000u l=180000u
+  ad=3.227e+11p pd=2.67e+06u as=0p ps=0u
M1020 a_657_325# a_532_93# a_101_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=2.432e+11p ps=2.04e+06u
M1021 a_1490_297# a_1089_297# a_681_49# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_101_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_101_21# C a_681_49# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_101_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_681_49# a_532_93# a_101_21# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_532_93# C VGND VNB nshort w=420000u l=150000u
+  ad=1.995e+11p pd=1.79e+06u as=0p ps=0u
M1027 a_1089_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.2e+11p pd=2.64e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a21bo_2 B1_N A2 X A1 VNB VPB VGND VPWR
M1000 a_621_47# A1 a_79_21# VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=2.145e+11p ps=1.96e+06u
M1001 VPWR A1 a_523_297# VPB phighvt w=1e+06u l=180000u
+  ad=9.372e+11p pd=8.18e+06u as=5.7e+11p ps=5.14e+06u
M1002 VGND A2 a_621_47# VNB nshort w=650000u l=150000u
+  ad=7.8875e+11p pd=7.68e+06u as=0p ps=0u
M1003 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1004 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.47e+11p ps=2.06e+06u
M1005 a_523_297# a_317_93# a_79_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1006 a_317_93# B1_N VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1007 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_317_93# B1_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1009 a_523_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_79_21# a_317_93# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__mux2i_2 Y A1 A0 S VNB VPB VPWR VGND
M1000 Y A0 a_401_47# VNB nshort w=650000u l=150000u
+  ad=7.3125e+11p pd=6.15e+06u as=4.16e+11p ps=3.88e+06u
M1001 a_211_297# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=8.5e+11p ps=7.7e+06u
M1002 a_213_47# S VGND VNB nshort w=650000u l=150000u
+  ad=4.1925e+11p pd=3.89e+06u as=5.85e+11p ps=5.7e+06u
M1003 a_401_47# A0 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_211_297# A0 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.065e+12p ps=8.13e+06u
M1005 VPWR S a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1006 VPWR a_27_47# a_399_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.85e+11p ps=5.17e+06u
M1007 a_213_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_27_47# a_401_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_399_297# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y A1 a_399_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND S a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1012 a_401_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_399_297# A1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR S a_211_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A0 a_211_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND S a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y A1 a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__decap_3 VPWR VGND VPB VNB
M1000 VPWR VGND VPWR VPB phighvt w=870000u l=590000u
+  ad=4.524e+11p pd=4.52e+06u as=0p ps=0u
M1001 VGND VPWR VGND VNB nshort w=550000u l=590000u
+  ad=2.86e+11p pd=3.24e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a31oi_2 A3 B1 Y A1 A2 VNB VPB VPWR VGND
M1000 Y A1 a_297_47# VNB nshort w=650000u l=150000u
+  ad=6.37e+11p pd=5.86e+06u as=4.68e+11p ps=4.04e+06u
M1001 a_27_297# A3 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.5e+12p pd=1.3e+07u as=1.47e+12p ps=8.94e+06u
M1002 a_27_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=5.46e+11p pd=5.58e+06u as=4.68e+11p ps=4.04e+06u
M1003 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_297_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_297_47# A2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A3 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.7e+11p pd=2.74e+06u as=0p ps=0u
M1009 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_297# B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A3 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_47# A2 a_297_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__conb_1 LO HI VPB VNB VGND VPWR
R0 VGND LO short w=480000u l=45000u
R1 HI VPWR short w=480000u l=45000u
.ends
.subckt sky130_fd_sc_hdll__dlrtn_2 RESET_B D GATE_N Q VGND VPWR VPB VNB
M1000 VGND a_750_21# a_708_47# VNB nshort w=420000u l=150000u
+  ad=8.0475e+11p pd=8.18e+06u as=8.82e+10p ps=1.26e+06u
M1001 VPWR GATE_N a_27_363# VPB phighvt w=640000u l=180000u
+  ad=1.411e+12p pd=1.231e+07u as=1.728e+11p ps=1.82e+06u
M1002 VPWR a_750_21# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1003 a_203_47# a_27_363# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1004 VPWR a_750_21# a_702_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1005 VGND a_750_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1006 a_503_369# a_319_369# VPWR VPB phighvt w=640000u l=180000u
+  ad=2.021e+11p pd=1.97e+06u as=0p ps=0u
M1007 a_708_47# a_203_47# a_604_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.58e+06u
M1008 Q a_750_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Q a_750_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND D a_319_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1011 VPWR D a_319_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1012 VGND RESET_B a_981_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.6575e+11p ps=1.81e+06u
M1013 a_604_47# a_27_363# a_500_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.58e+06u
M1014 VPWR RESET_B a_750_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1015 a_981_47# a_604_47# a_750_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1016 VGND GATE_N a_27_363# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1017 a_702_413# a_27_363# a_604_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1018 a_203_47# a_27_363# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1019 a_604_47# a_203_47# a_503_369# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_500_47# a_319_369# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_750_21# a_604_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or2b_2 A B_N X VPWR VGND VNB VPB
M1000 VGND B_N a_27_53# VNB nshort w=420000u l=150000u
+  ad=7.764e+11p pd=6.48e+06u as=1.302e+11p ps=1.46e+06u
M1001 a_228_297# a_27_53# VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1002 VPWR a_228_297# X VPB phighvt w=1e+06u l=180000u
+  ad=7.191e+11p pd=6.69e+06u as=4.8e+11p ps=2.96e+06u
M1003 a_27_53# B_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1004 a_318_297# a_27_53# a_228_297# VPB phighvt w=420000u l=180000u
+  ad=9.66e+10p pd=1.3e+06u as=1.134e+11p ps=1.38e+06u
M1005 VPWR A a_318_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_228_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.315e+11p ps=2.32e+06u
M1007 X a_228_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_228_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A a_228_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__diode_8 VNB VPB VGND VPWR DIODE
D0 VNB DIODE ndiode p=1.858e+07u a=3.5464e+12p
.ends
.subckt sky130_fd_sc_hdll__sdfxtp_1 VPWR VGND CLK Q SCD D SCE VPB VNB
M1000 VPWR a_1189_21# a_1121_413# VPB phighvt w=420000u l=180000u
+  ad=1.3699e+12p pd=1.231e+07u as=1.47e+11p ps=1.54e+06u
M1001 VGND a_1474_413# a_1647_21# VNB nshort w=650000u l=150000u
+  ad=1.0782e+12p pd=1.048e+07u as=2.015e+11p ps=1.92e+06u
M1002 VPWR CLK a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1003 a_608_369# D a_507_47# VNB nshort w=420000u l=150000u
+  ad=2.604e+11p pd=2.88e+06u as=1.638e+11p ps=1.62e+06u
M1004 a_1474_413# a_27_47# a_1189_21# VPB phighvt w=420000u l=180000u
+  ad=1.26e+11p pd=1.44e+06u as=2.4195e+11p ps=2.22e+06u
M1005 VGND a_1189_21# a_1117_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.446e+11p ps=1.56e+06u
M1006 a_504_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=2.176e+11p pd=1.96e+06u as=0p ps=0u
M1007 a_203_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1008 VGND a_1647_21# a_1581_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.338e+11p ps=1.5e+06u
M1009 VPWR SCE a_319_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1010 VPWR a_1647_21# a_1570_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.659e+11p ps=1.63e+06u
M1011 a_1121_413# a_27_47# a_1011_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.407e+11p ps=1.51e+06u
M1012 a_1189_21# a_1011_47# VGND VNB nshort w=640000u l=150000u
+  ad=2.104e+11p pd=2.06e+06u as=0p ps=0u
M1013 VGND SCE a_319_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.428e+11p ps=1.52e+06u
M1014 a_1011_47# a_203_47# a_608_369# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=3.2e+11p ps=3.34e+06u
M1015 a_1570_413# a_203_47# a_1474_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Q a_1647_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1017 a_203_47# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1018 a_1474_413# a_203_47# a_1189_21# VNB nshort w=360000u l=150000u
+  ad=1.35e+11p pd=1.47e+06u as=0p ps=0u
M1019 VPWR SCD a_702_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=2.144e+11p ps=1.95e+06u
M1020 VGND SCD a_721_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=9.66e+10p ps=1.3e+06u
M1021 a_507_47# a_319_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_702_369# a_319_47# a_608_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1117_47# a_203_47# a_1011_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.368e+11p ps=1.48e+06u
M1024 VPWR a_1474_413# a_1647_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1025 a_1189_21# a_1011_47# VPWR VPB phighvt w=750000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1011_47# a_27_47# a_608_369# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1581_47# a_27_47# a_1474_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1029 a_721_47# SCE a_608_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_608_369# D a_504_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Q a_1647_21# VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a211o_4 VNB VPB VGND VPWR C1 B1 X A2 A1
M1000 VPWR A2 a_523_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.55e+12p pd=1.31e+07u as=1.25e+12p ps=1.05e+07u
M1001 X a_79_204# VGND VNB nshort w=650000u l=150000u
+  ad=4.7125e+11p pd=4.05e+06u as=1.43325e+12p ps=1.221e+07u
M1002 a_1051_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=0p ps=0u
M1003 VPWR a_79_204# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=6e+11p ps=5.2e+06u
M1004 VGND a_79_204# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_79_204# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_79_204# C1 a_613_297# VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=3e+11p ps=2.6e+06u
M1007 a_79_204# B1 VGND VNB nshort w=650000u l=150000u
+  ad=7.41e+11p pd=6.18e+06u as=0p ps=0u
M1008 VPWR A1 a_523_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_79_204# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_79_204# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_79_204# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_79_204# C1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND B1 a_79_204# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1243_47# A1 a_79_204# VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=0p ps=0u
M1015 a_523_297# B1 a_805_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.4e+11p ps=2.68e+06u
M1016 a_79_204# A1 a_1051_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_613_297# B1 a_523_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_523_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A2 a_1243_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_79_204# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_523_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_805_297# C1 a_79_204# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND C1 a_79_204# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a2bb2oi_2 A2_N A1_N Y B2 B1 VNB VPB VGND VPWR
M1000 a_27_297# B2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.12e+12p pd=1.024e+07u as=8.7e+11p ps=7.74e+06u
M1001 a_695_297# A2_N a_455_21# VPB phighvt w=1e+06u l=180000u
+  ad=8.5e+11p pd=7.7e+06u as=2.9e+11p ps=2.58e+06u
M1002 a_27_297# a_455_21# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1003 Y B2 a_119_47# VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=3.835e+11p ps=3.78e+06u
M1004 a_455_21# A1_N VGND VNB nshort w=650000u l=150000u
+  ad=4.81e+11p pd=4.08e+06u as=1.2805e+12p ps=1.044e+07u
M1005 VPWR B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2_N a_455_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y a_455_21# a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_455_21# A2_N a_695_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_119_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_695_297# A1_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A1_N a_455_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_455_21# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y a_455_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_455_21# A2_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A1_N a_695_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_119_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a21o_4 A2 A1 X B1 VNB VPB VGND VPWR
M1000 VGND B1 a_84_21# VNB nshort w=650000u l=150000u
+  ad=1.365e+12p pd=1.07e+07u as=4.81e+11p ps=4.08e+06u
M1001 a_523_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.255e+12p pd=1.051e+07u as=1.47e+12p ps=1.294e+07u
M1002 X a_84_21# VGND VNB nshort w=650000u l=150000u
+  ad=4.29e+11p pd=3.92e+06u as=0p ps=0u
M1003 VPWR a_84_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=6e+11p ps=5.2e+06u
M1004 VPWR A2 a_523_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_84_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_84_21# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_801_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=0p ps=0u
M1008 VGND a_84_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_991_47# A1 a_84_21# VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1010 VGND A2 a_991_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_523_297# B1 a_84_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1012 VPWR a_84_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_523_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_84_21# B1 a_523_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A1 a_523_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_84_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_84_21# A1 a_801_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_84_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_84_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__dlygate4sd1_1 A X VPWR VGND VPB VNB
M1000 a_213_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=5.039e+11p ps=3.97e+06u
M1001 X a_319_93# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1002 VPWR a_213_47# a_319_93# VPB phighvt w=420000u l=180000u
+  ad=6.233e+11p pd=4.51e+06u as=1.176e+11p ps=1.4e+06u
M1003 X a_319_93# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1004 a_213_47# a_27_47# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1005 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1006 VGND a_213_47# a_319_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1007 VPWR A a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
.ends
.subckt sky130_fd_sc_hdll__sdfxbp_2 VPWR VGND Q_N Q CLK SCE D SCD VNB VPB
M1000 VPWR a_1179_183# a_1111_413# VPB phighvt w=420000u l=180000u
+  ad=2.67555e+12p pd=2.099e+07u as=1.47e+11p ps=1.54e+06u
M1001 a_211_363# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.9813e+12p ps=1.723e+07u
M1002 a_1179_183# a_1001_47# VGND VNB nshort w=640000u l=150000u
+  ad=1.978e+11p pd=1.99e+06u as=0p ps=0u
M1003 VPWR a_1653_315# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1004 VGND a_2234_47# Q_N VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1005 VPWR a_2234_47# Q_N VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1006 Q_N a_2234_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR SCD a_698_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=2.144e+11p ps=1.95e+06u
M1008 a_1464_413# a_27_47# a_1179_183# VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=2.307e+11p ps=2.19e+06u
M1009 a_1001_47# a_27_47# a_604_369# VNB nshort w=360000u l=150000u
+  ad=1.548e+11p pd=1.58e+06u as=2.604e+11p ps=2.88e+06u
M1010 VPWR CLK a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1011 a_698_369# a_319_47# a_604_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=2.99e+11p ps=3.24e+06u
M1012 Q_N a_2234_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Q a_1653_315# VGND VNB nshort w=650000u l=150000u
+  ad=2.08e+11p pd=1.94e+06u as=0p ps=0u
M1014 a_604_369# D a_529_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1015 VPWR a_1464_413# a_1653_315# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1016 a_503_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=2.08e+11p pd=1.93e+06u as=0p ps=0u
M1017 VGND a_1179_183# a_1117_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.374e+11p ps=1.52e+06u
M1018 VPWR a_1653_315# a_2234_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1019 a_717_47# SCE a_604_369# VNB nshort w=420000u l=150000u
+  ad=9.66e+10p pd=1.3e+06u as=0p ps=0u
M1020 a_604_369# D a_503_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND SCE a_319_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1022 VPWR SCE a_319_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1023 a_1111_413# a_27_47# a_1001_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.407e+11p ps=1.51e+06u
M1024 VGND a_1653_315# a_1615_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.446e+11p ps=1.55e+06u
M1025 a_1179_183# a_1001_47# VPWR VPB phighvt w=750000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Q a_1653_315# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_1653_315# a_2234_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1028 a_1001_47# a_211_363# a_604_369# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1030 a_1464_413# a_211_363# a_1179_183# VNB nshort w=360000u l=150000u
+  ad=1.854e+11p pd=1.75e+06u as=0p ps=0u
M1031 a_529_47# a_319_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR a_1653_315# a_1558_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=2.037e+11p ps=1.81e+06u
M1033 a_211_363# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1034 a_1117_47# a_211_363# a_1001_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND a_1653_315# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1558_413# a_211_363# a_1464_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND SCD a_717_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1615_47# a_27_47# a_1464_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND a_1464_413# a_1653_315# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
.ends
.subckt sky130_fd_sc_hdll__nor2b_2 B_N A Y VPB VNB VGND VPWR
M1000 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=4.034e+11p pd=3.96e+06u as=8.5e+11p ps=7.7e+06u
M1001 a_27_297# a_271_21# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1002 VPWR B_N a_271_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.806e+11p ps=1.7e+06u
M1003 Y a_271_21# a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VGND VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=6.8595e+11p ps=7.07e+06u
M1005 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_271_21# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y a_271_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B_N a_271_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=1.68e+06u
.ends
.subckt sky130_fd_sc_hdll__nor4_8 A C D B Y VPB VNB VGND VPWR
M1000 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.57e+12p pd=2.314e+07u as=1.16e+12p ps=1.032e+07u
M1001 a_869_297# C a_1635_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.32e+12p pd=2.064e+07u as=2.58e+12p ps=2.316e+07u
M1002 Y B VGND VNB nshort w=650000u l=150000u
+  ad=2.808e+12p pd=2.944e+07u as=4.355e+12p ps=3.55e+07u
M1003 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_297# B a_869_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_1635_297# D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.16e+12p ps=1.032e+07u
M1007 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_869_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y D a_1635_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_869_297# C a_1635_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_869_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1635_297# C a_869_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1635_297# C a_869_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND D Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y D a_1635_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_869_297# C a_1635_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND D Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1635_297# D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND D Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_869_297# C a_1635_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_27_297# B a_869_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Y D a_1635_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1635_297# D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 Y D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_27_297# B a_869_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_1635_297# D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1045 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_869_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1048 VGND D Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 Y D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1050 a_1635_297# C a_869_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1051 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1052 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1053 a_27_297# B a_869_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1054 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1055 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1056 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1057 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1058 a_869_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1059 a_1635_297# C a_869_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1060 Y D a_1635_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1061 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1062 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1063 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__einvp_4 TE A Z VPWR VGND VPB VNB
M1000 a_213_47# TE VGND VNB nshort w=650000u l=150000u
+  ad=1.0205e+12p pd=9.64e+06u as=5.98e+11p ps=5.74e+06u
M1001 a_213_47# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1002 Z A a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR a_27_47# a_235_309# VPB phighvt w=940000u l=180000u
+  ad=8.152e+11p pd=7.46e+06u as=1.4263e+12p ps=1.269e+07u
M1004 VPWR TE a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1005 a_235_309# A Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1006 VGND TE a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_213_47# TE VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_213_47# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Z A a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND TE a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_235_309# a_27_47# VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Z A a_235_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND TE a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1014 a_235_309# A Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_27_47# a_235_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_235_309# a_27_47# VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Z A a_235_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__muxb8to1_1 VGND Z VPWR VNB VPB D[0] S[0] S[1] D[1] D[2]
+ S[2] S[3] D[4] S[4] S[5] D[5] D[6] S[6] S[7] D[7] D[3]
M1000 a_1765_47# D[4] VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=1.8759e+12p ps=1.712e+07u
M1001 a_937_47# D[2] VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1002 a_2593_47# D[6] VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1003 a_1773_297# D[4] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=3.19e+12p ps=2.438e+07u
M1004 VGND S[6] a_2668_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.61e+06u
M1005 a_1361_47# S[3] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1006 VPWR D[7] a_3218_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.297e+11p ps=2.69e+06u
M1007 Z a_1840_265# a_1773_297# VPB phighvt w=820000u l=180000u
+  ad=1.7712e+12p pd=1.744e+07u as=0p ps=0u
M1008 a_1574_47# S[3] Z VNB nshort w=520000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=1.0816e+12p ps=1.248e+07u
M1009 a_734_333# a_533_47# Z VPB phighvt w=820000u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1010 Z S[2] a_937_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_3017_47# S[7] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1012 a_2402_47# S[5] Z VNB nshort w=520000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1013 a_1562_333# a_1361_47# Z VPB phighvt w=820000u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1014 a_746_47# S[1] Z VNB nshort w=520000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1015 a_117_297# D[0] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1016 VPWR D[3] a_1562_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_2601_297# D[6] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1018 Z S[4] a_1765_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Z a_184_265# a_117_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_533_47# S[1] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1021 a_945_297# D[2] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1022 Z a_1012_265# a_945_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR S[0] a_184_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1024 a_2189_47# S[5] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1025 VPWR S[2] a_1012_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1026 Z a_2668_265# a_2601_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1361_47# S[3] VGND VNB nshort w=520000u l=150000u
+  ad=1.482e+11p pd=1.61e+06u as=0p ps=0u
M1028 a_533_47# S[1] VGND VNB nshort w=520000u l=150000u
+  ad=1.482e+11p pd=1.61e+06u as=0p ps=0u
M1029 VGND S[0] a_184_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.61e+06u
M1030 a_2390_333# a_2189_47# Z VPB phighvt w=820000u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1031 a_3230_47# S[7] Z VNB nshort w=520000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1032 VGND D[1] a_746_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Z S[6] a_2593_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR S[6] a_2668_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1035 VPWR D[1] a_734_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR D[5] a_2390_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_2189_47# S[5] VGND VNB nshort w=520000u l=150000u
+  ad=1.482e+11p pd=1.61e+06u as=0p ps=0u
M1038 VPWR S[4] a_1840_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1039 VGND D[3] a_1574_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_109_47# D[0] VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1041 VGND D[5] a_2402_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VGND S[2] a_1012_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.61e+06u
M1043 VGND D[7] a_3230_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 Z S[0] a_109_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_3218_333# a_3017_47# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1046 VGND S[4] a_1840_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.61e+06u
M1047 a_3017_47# S[7] VGND VNB nshort w=520000u l=150000u
+  ad=1.482e+11p pd=1.61e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o2bb2a_1 A1_N X A2_N B2 B1 VNB VPB VPWR VGND
M1000 VPWR A2_N a_224_369# VPB phighvt w=420000u l=180000u
+  ad=8.398e+11p pd=6.8e+06u as=2.664e+11p ps=2.4e+06u
M1001 a_225_47# A1_N VGND VNB nshort w=420000u l=150000u
+  ad=1.323e+11p pd=1.47e+06u as=3.9885e+11p ps=3.76e+06u
M1002 VPWR a_76_199# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1003 VGND B2 a_529_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.646e+11p ps=2.94e+06u
M1004 a_224_369# A2_N a_225_47# VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1005 a_633_369# B2 a_76_199# VPB phighvt w=420000u l=180000u
+  ad=1.638e+11p pd=1.62e+06u as=1.47e+11p ps=1.54e+06u
M1006 a_224_369# A1_N VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR B1 a_633_369# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_529_47# B1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_76_199# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1010 a_529_47# a_224_369# a_76_199# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1011 a_76_199# a_224_369# VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or3_1 A X B C VPWR VGND VPB VNB
M1000 X a_29_53# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=4.95e+11p pd=2.99e+06u as=3.107e+11p ps=2.72e+06u
M1001 VGND C a_29_53# VNB nshort w=420000u l=150000u
+  ad=3.4965e+11p pd=3.46e+06u as=2.856e+11p ps=3.04e+06u
M1002 a_119_297# C a_29_53# VPB phighvt w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=1.134e+11p ps=1.38e+06u
M1003 VPWR A a_203_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.428e+11p ps=1.52e+06u
M1004 X a_29_53# VGND VNB nshort w=650000u l=150000u
+  ad=3.1525e+11p pd=2.27e+06u as=0p ps=0u
M1005 VGND A a_29_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_203_297# B a_119_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_29_53# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and4b_2 VPWR VGND X A_N D C B VNB VPB
M1000 VPWR D a_211_413# VPB phighvt w=420000u l=180000u
+  ad=8.563e+11p pd=8.28e+06u as=4.683e+11p ps=3.91e+06u
M1001 VPWR A_N a_27_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1002 VGND D a_519_47# VNB nshort w=420000u l=150000u
+  ad=5.3965e+11p pd=5.38e+06u as=1.449e+11p ps=1.53e+06u
M1003 VGND a_211_413# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.3075e+11p ps=2.01e+06u
M1004 X a_211_413# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.25e+11p pd=2.65e+06u as=0p ps=0u
M1005 a_399_47# B a_317_47# VNB nshort w=420000u l=150000u
+  ad=1.89e+11p pd=1.74e+06u as=1.092e+11p ps=1.36e+06u
M1006 VPWR B a_211_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_211_413# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_413# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1009 a_211_413# C VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_317_47# a_27_413# a_211_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1011 a_211_413# a_27_413# VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_211_413# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_519_47# C a_399_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o22ai_1 B2 A1 Y B1 A2 VPB VNB VPWR VGND
M1000 VGND A2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=7.605e+11p ps=6.24e+06u
M1001 VPWR A1 a_384_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.5e+11p pd=5.1e+06u as=2.3e+11p ps=2.46e+06u
M1002 a_384_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.6e+11p ps=3.12e+06u
M1003 a_27_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.5675e+11p ps=2.09e+06u
M1004 a_117_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=4.15e+11p pd=2.83e+06u as=0p ps=0u
M1005 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a31o_2 X B1 A3 A1 A2 VNB VPB VGND VPWR
M1000 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=9.1e+11p pd=7.82e+06u as=2.9e+11p ps=2.58e+06u
M1001 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=5.46e+11p pd=5.58e+06u as=2.405e+11p ps=2.04e+06u
M1002 a_79_21# A1 a_391_47# VNB nshort w=650000u l=150000u
+  ad=3.38e+11p pd=2.34e+06u as=2.47e+11p ps=2.06e+06u
M1003 VGND B1 a_79_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_305_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6.4e+11p pd=5.28e+06u as=0p ps=0u
M1005 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A2 a_305_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_79_21# B1 a_305_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.3e+11p pd=2.66e+06u as=0p ps=0u
M1008 a_305_297# A3 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_391_47# A2 a_307_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1011 a_307_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__xnor3_2 X B C A VNB VPB VGND VPWR
M1000 a_477_49# a_328_93# a_79_21# VPB phighvt w=840000u l=180000u
+  ad=8.3175e+11p pd=5.4e+06u as=3.227e+11p ps=2.67e+06u
M1001 a_1286_297# a_885_297# a_453_325# VNB nshort w=420000u l=150000u
+  ad=7.149e+11p pd=4.88e+06u as=6.411e+11p ps=4.67e+06u
M1002 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=8.543e+11p pd=7.87e+06u as=2.405e+11p ps=2.04e+06u
M1003 a_328_93# C VPWR VPB phighvt w=640000u l=180000u
+  ad=1.856e+11p pd=1.86e+06u as=1.22095e+12p ps=1.051e+07u
M1004 a_477_49# B a_1286_297# VNB nshort w=640000u l=150000u
+  ad=5.4545e+11p pd=4.31e+06u as=0p ps=0u
M1005 a_885_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.2e+11p pd=2.64e+06u as=0p ps=0u
M1006 a_453_325# B a_1286_297# VPB phighvt w=640000u l=180000u
+  ad=6.39e+11p pd=4.96e+06u as=9.286e+11p ps=5.88e+06u
M1007 a_79_21# C a_477_49# VNB nshort w=640000u l=150000u
+  ad=1.856e+11p pd=1.86e+06u as=0p ps=0u
M1008 a_453_325# a_328_93# a_79_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_328_93# C VGND VNB nshort w=420000u l=150000u
+  ad=1.995e+11p pd=1.79e+06u as=0p ps=0u
M1010 a_477_49# B a_1003_297# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=7.226e+11p ps=5.29e+06u
M1011 a_1286_297# a_1003_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1003_297# a_885_297# a_477_49# VNB nshort w=600000u l=150000u
+  ad=4.4975e+11p pd=3.99e+06u as=0p ps=0u
M1013 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.1e+11p pd=2.62e+06u as=0p ps=0u
M1014 a_1003_297# a_885_297# a_453_325# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_453_325# B a_1003_297# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_79_21# C a_453_325# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1286_297# a_885_297# a_477_49# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A a_1003_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1286_297# a_1003_297# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A a_1003_297# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_885_297# B VGND VNB nshort w=650000u l=150000u
+  ad=1.6515e+11p pd=1.82e+06u as=0p ps=0u
M1023 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand2b_1 Y A_N B VPB VNB VGND VPWR
M1000 VPWR A_N a_27_93# VPB phighvt w=420000u l=180000u
+  ad=5.757e+11p pd=5.25e+06u as=1.134e+11p ps=1.38e+06u
M1001 VPWR a_27_93# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1002 VGND A_N a_27_93# VNB nshort w=420000u l=150000u
+  ad=2.33e+11p pd=2.07e+06u as=1.302e+11p ps=1.46e+06u
M1003 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y a_27_93# a_226_47# VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=1.755e+11p ps=1.84e+06u
M1005 a_226_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand4bb_4 B_N A_N C Y D VNB VPB VGND VPWR
M1000 a_1251_47# C a_853_47# VNB nshort w=650000u l=150000u
+  ad=1.02375e+12p pd=9.65e+06u as=8.645e+11p ps=7.86e+06u
M1001 a_206_47# B_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=4.55e+11p pd=2.91e+06u as=3.425e+12p ps=2.685e+07u
M1002 a_395_47# a_206_47# a_853_47# VNB nshort w=650000u l=150000u
+  ad=9.62e+11p pd=9.46e+06u as=0p ps=0u
M1003 Y a_206_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.32e+12p pd=2.064e+07u as=0p ps=0u
M1004 VPWR a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y a_27_47# a_395_47# VNB nshort w=650000u l=150000u
+  ad=4.16e+11p pd=3.88e+06u as=0p ps=0u
M1008 a_853_47# a_206_47# a_395_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_853_47# C a_1251_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1251_47# C a_853_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_206_47# B_N VGND VNB nshort w=650000u l=150000u
+  ad=3.12e+11p pd=2.26e+06u as=6.0125e+11p ps=5.75e+06u
M1014 VPWR A_N a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1015 VPWR a_206_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1251_47# D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND D a_1251_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y a_206_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_853_47# C a_1251_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A_N a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1022 VPWR a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_395_47# a_206_47# a_853_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1251_47# D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_853_47# a_206_47# a_395_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND D a_1251_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR a_206_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_395_47# a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Y a_27_47# a_395_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Y a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_395_47# a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o211ai_1 A1 A2 Y C1 B1 VPB VNB VGND VPWR
M1000 VGND A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=3.9325e+11p ps=3.81e+06u
M1001 a_27_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A2 a_118_297# VPB phighvt w=1e+06u l=180000u
+  ad=9.2e+11p pd=5.84e+06u as=2.3e+11p ps=2.46e+06u
M1003 VPWR B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=6.2e+11p pd=5.24e+06u as=0p ps=0u
M1004 Y C1 a_304_47# VNB nshort w=650000u l=150000u
+  ad=3.77e+11p pd=2.46e+06u as=2.4375e+11p ps=2.05e+06u
M1005 a_118_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y C1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_304_47# B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__muxb16to1_4 VGND Z VPWR VNB VPB S[6] S[10] D[12] D[13]
+ D[8] D[15] D[10] D[9] D[14] S[14] D[11] S[11] S[8] S[15] S[12] S[9] S[13] D[3] D[0]
+ D[4] D[5] D[2] D[1] D[6] S[2] S[3] S[7] S[0] S[1] S[4] S[5] D[7]
M1000 a_2693_591# a_3135_793# Z VPB phighvt w=820000u l=180000u
+  ad=1.2606e+12p pd=1.174e+07u as=7.6096e+12p ps=7.104e+07u
M1001 a_2695_47# D[2] VGND VNB nshort w=650000u l=150000u
+  ad=7.618e+11p pd=8.38e+06u as=1.32704e+13p ps=1.36e+08u
M1002 a_1643_311# D[1] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.2606e+12p pd=1.174e+07u as=2.03648e+13p ps=1.9232e+08u
M1003 a_9513_66# S[7] Z VNB nshort w=520000u l=150000u
+  ad=7.618e+11p pd=8.38e+06u as=4.4928e+12p ps=5.056e+07u
M1004 a_7939_911# D[14] VGND VNB nshort w=650000u l=150000u
+  ad=7.618e+11p pd=8.38e+06u as=0p ps=0u
M1005 a_7939_911# S[14] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_5361_591# D[12] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.2606e+12p pd=1.174e+07u as=0p ps=0u
M1007 Z a_1430_325# a_1643_311# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1430_599# S[9] VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1009 a_8379_265# S[6] VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1010 a_2695_911# S[10] Z VNB nshort w=520000u l=150000u
+  ad=7.618e+11p pd=8.38e+06u as=0p ps=0u
M1011 a_1643_613# D[9] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.2606e+12p pd=1.174e+07u as=0p ps=0u
M1012 VGND D[12] a_5363_911# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.618e+11p ps=8.38e+06u
M1013 Z a_9250_325# a_9463_311# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=1.2606e+12p ps=1.174e+07u
M1014 VPWR D[0] a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.2606e+12p ps=1.174e+07u
M1015 VPWR S[6] a_8379_265# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1016 VPWR S[4] a_5803_265# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1017 a_559_793# S[8] VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1018 VPWR S[0] a_559_265# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1019 VGND D[9] a_1693_918# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.618e+11p ps=8.38e+06u
M1020 a_2693_297# D[2] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.2606e+12p pd=1.174e+07u as=0p ps=0u
M1021 VGND D[4] a_5363_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.618e+11p ps=8.38e+06u
M1022 a_6674_325# S[5] VPWR VPB phighvt w=820000u l=180000u
+  ad=2.378e+11p pd=2.22e+06u as=0p ps=0u
M1023 VPWR D[8] a_117_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.2606e+12p ps=1.174e+07u
M1024 a_2693_591# D[10] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_7937_591# a_8379_793# Z VPB phighvt w=820000u l=180000u
+  ad=1.2606e+12p pd=1.174e+07u as=0p ps=0u
M1026 Z a_559_793# a_117_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Z S[9] a_1693_918# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_8379_793# S[14] VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1029 VGND D[5] a_6937_66# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.618e+11p ps=8.38e+06u
M1030 a_4269_66# S[3] Z VNB nshort w=520000u l=150000u
+  ad=7.618e+11p pd=8.38e+06u as=0p ps=0u
M1031 Z S[3] a_4269_66# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1693_918# S[9] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND D[10] a_2695_911# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR S[13] a_6674_599# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1035 Z S[2] a_2695_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_2695_47# S[2] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND S[4] a_5803_265# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1038 VPWR D[1] a_1643_311# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 Z S[1] a_1693_66# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=7.618e+11p ps=8.38e+06u
M1040 VPWR D[7] a_9463_311# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND D[3] a_4269_66# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPWR D[3] a_4219_311# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.2606e+12p ps=1.174e+07u
M1043 a_3135_793# S[10] VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1044 a_5363_911# S[12] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_1693_66# S[1] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 Z a_6674_325# a_6887_311# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=1.2606e+12p ps=1.174e+07u
M1047 a_4269_918# S[11] Z VNB nshort w=520000u l=150000u
+  ad=7.618e+11p pd=8.38e+06u as=0p ps=0u
M1048 a_1643_311# a_1430_325# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1049 VGND D[1] a_1693_66# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1050 a_5361_297# a_5803_265# Z VPB phighvt w=820000u l=180000u
+  ad=1.2606e+12p pd=1.174e+07u as=0p ps=0u
M1051 VPWR D[9] a_1643_613# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1052 VPWR D[11] a_4219_613# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.2606e+12p ps=1.174e+07u
M1053 a_119_47# S[0] Z VNB nshort w=520000u l=150000u
+  ad=7.618e+11p pd=8.38e+06u as=0p ps=0u
M1054 VGND S[11] a_4006_599# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1055 Z a_5803_793# a_5361_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1056 VPWR D[15] a_9463_613# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.2606e+12p ps=1.174e+07u
M1057 a_6937_66# D[5] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1058 a_9463_311# a_9250_325# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1059 Z S[3] a_4269_66# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1060 VGND S[13] a_6674_599# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1061 a_559_265# S[0] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1062 VGND D[2] a_2695_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1063 a_8379_265# S[6] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1064 Z S[14] a_7939_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1065 a_3135_265# S[2] VPWR VPB phighvt w=820000u l=180000u
+  ad=2.378e+11p pd=2.22e+06u as=0p ps=0u
M1066 VPWR S[11] a_4006_599# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1067 VPWR D[2] a_2693_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1068 VGND D[7] a_9513_66# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1069 a_7939_47# D[6] VGND VNB nshort w=650000u l=150000u
+  ad=7.618e+11p pd=8.38e+06u as=0p ps=0u
M1070 Z S[8] a_119_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=7.618e+11p ps=8.38e+06u
M1071 a_4219_613# a_4006_599# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1072 a_4006_599# S[11] VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1073 a_9513_918# D[15] VGND VNB nshort w=650000u l=150000u
+  ad=7.618e+11p pd=8.38e+06u as=0p ps=0u
M1074 Z S[0] a_119_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1075 VGND S[6] a_8379_265# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1076 VPWR D[10] a_2693_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1077 Z a_8379_793# a_7937_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1078 VGND S[8] a_559_793# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1079 a_117_591# a_559_793# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1080 Z a_3135_793# a_2693_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1081 a_7937_297# a_8379_265# Z VPB phighvt w=820000u l=180000u
+  ad=1.2606e+12p pd=1.174e+07u as=0p ps=0u
M1082 a_2693_297# a_3135_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1083 VPWR S[10] a_3135_793# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1084 VGND D[0] a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1085 VGND D[8] a_119_911# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1086 a_5803_265# S[4] VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1087 a_9463_311# D[7] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1088 VPWR D[5] a_6887_311# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1089 a_4219_311# D[3] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1090 a_119_911# D[8] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1091 a_5363_911# S[12] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1092 Z a_6674_599# a_6887_613# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=1.2606e+12p ps=1.174e+07u
M1093 Z S[1] a_1693_66# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1094 a_6887_311# a_6674_325# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1095 a_5803_265# S[4] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1096 a_1693_918# S[9] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1097 VGND S[14] a_8379_793# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1098 a_1693_66# D[1] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1099 VPWR D[6] a_7937_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1100 a_4269_66# D[3] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1101 a_4219_613# D[11] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1102 VPWR D[13] a_6887_613# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1103 a_9463_613# D[15] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1104 Z S[15] a_9513_918# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1105 a_119_47# S[0] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1106 a_4269_66# S[3] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1107 VGND S[9] a_1430_599# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1108 a_2695_47# S[2] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1109 VPWR D[14] a_7937_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1110 a_2695_47# D[2] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1111 a_1693_918# D[9] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1112 a_1643_613# a_1430_599# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1113 a_1693_66# S[1] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1114 Z a_4006_599# a_4219_613# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1115 a_9513_66# D[7] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1116 VPWR D[3] a_4219_311# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1117 a_6887_613# a_6674_599# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1118 a_5361_297# a_5803_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1119 Z a_5803_793# a_5361_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1120 VPWR S[12] a_5803_793# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1121 a_4219_311# a_4006_325# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1122 VGND D[6] a_7939_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1123 VPWR S[8] a_559_793# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1124 VPWR S[14] a_8379_793# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1125 Z S[0] a_119_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1126 VGND S[5] a_6674_325# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1127 Z a_559_793# a_117_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1128 a_5363_911# D[12] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1129 VPWR D[11] a_4219_613# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1130 a_6674_599# S[13] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1131 a_9463_311# D[7] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1132 VGND D[13] a_6937_918# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.618e+11p ps=8.38e+06u
M1133 VPWR S[1] a_1430_325# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1134 a_1643_311# D[1] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1135 a_4269_66# D[3] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1136 a_6937_918# D[13] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1137 a_117_297# a_559_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1138 Z a_3135_265# a_2693_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1139 a_559_265# S[0] VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1140 Z a_1430_325# a_1643_311# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1141 a_9250_325# S[7] VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1142 VPWR S[7] a_9250_325# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1143 a_2695_911# D[10] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1144 VGND D[15] a_9513_918# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1145 a_9463_613# D[15] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1146 a_117_297# D[0] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1147 a_7939_47# D[6] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1148 a_1643_613# D[9] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1149 a_6937_918# S[13] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1150 a_4006_325# S[3] VPWR VPB phighvt w=820000u l=180000u
+  ad=2.378e+11p pd=2.22e+06u as=0p ps=0u
M1151 VPWR D[7] a_9463_311# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1152 a_6674_325# S[5] VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1153 Z a_9250_325# a_9463_311# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1154 Z S[4] a_5363_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1155 a_117_591# D[8] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1156 VPWR D[15] a_9463_613# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1157 a_2693_297# D[2] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1158 VPWR D[4] a_5361_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1159 a_119_911# S[8] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1160 Z S[11] a_4269_918# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1161 Z a_1430_599# a_1643_613# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1162 Z S[14] a_7939_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1163 a_9463_311# a_9250_325# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1164 a_2693_591# D[10] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1165 VPWR D[12] a_5361_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1166 Z a_9250_599# a_9463_613# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1167 VGND D[1] a_1693_66# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1168 Z a_8379_265# a_7937_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1169 a_9513_918# S[15] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1170 a_8379_793# S[14] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1171 Z a_4006_325# a_4219_311# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1172 a_559_793# S[8] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1173 a_3135_793# S[10] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1174 a_9250_599# S[15] VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1175 a_6937_66# S[5] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1176 VPWR D[6] a_7937_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1177 a_5363_47# D[4] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1178 VGND D[9] a_1693_918# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1179 VGND D[14] a_7939_911# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1180 a_1430_325# S[1] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1181 a_2693_297# a_3135_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1182 VGND D[2] a_2695_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1183 a_6887_311# D[5] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1184 VPWR D[14] a_7937_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1185 a_9250_325# S[7] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1186 a_6887_613# D[13] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1187 VGND D[12] a_5363_911# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1188 a_5803_793# S[12] VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1189 VGND D[14] a_7939_911# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1190 a_9513_918# D[15] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1191 Z S[4] a_5363_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1192 VGND S[0] a_559_265# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1193 VGND D[3] a_4269_66# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1194 a_5361_297# D[4] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1195 VGND D[10] a_2695_911# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1196 Z a_6674_599# a_6887_613# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1197 Z S[15] a_9513_918# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1198 VGND S[7] a_9250_325# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1199 a_1643_613# a_1430_599# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1200 a_5361_591# a_5803_793# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1201 a_5803_793# S[12] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1202 a_7939_47# S[6] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1203 a_5361_591# D[12] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1204 a_9463_613# a_9250_599# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1205 a_5363_47# S[4] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1206 a_7937_297# a_8379_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1207 Z a_559_265# a_117_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1208 VPWR D[0] a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1209 Z S[7] a_9513_66# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1210 a_6937_66# S[5] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1211 a_6674_599# S[13] VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1212 Z S[6] a_7939_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1213 a_5363_47# S[4] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1214 Z S[10] a_2695_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1215 VGND S[10] a_3135_793# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1216 a_9513_66# D[7] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1217 VPWR D[5] a_6887_311# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1218 Z S[12] a_5363_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1219 a_119_47# D[0] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1220 Z S[5] a_6937_66# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1221 VPWR D[8] a_117_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1222 VGND S[2] a_3135_265# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1223 VGND S[15] a_9250_599# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1224 VPWR D[13] a_6887_613# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1225 VPWR S[9] a_1430_599# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1226 a_6937_918# S[13] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1227 a_7937_591# a_8379_793# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1228 Z S[5] a_6937_66# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1229 a_2693_591# a_3135_793# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1230 a_7939_911# S[14] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1231 Z a_5803_265# a_5361_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1232 VGND D[4] a_5363_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1233 VPWR S[15] a_9250_599# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1234 VGND S[3] a_4006_325# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1235 VGND D[8] a_119_911# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1236 a_119_911# S[8] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1237 a_4006_599# S[11] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1238 a_6887_613# a_6674_599# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1239 a_3135_265# S[2] VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1240 a_119_911# D[8] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1241 VGND S[1] a_1430_325# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1242 Z S[13] a_6937_918# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1243 a_4219_311# a_4006_325# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1244 a_7939_47# S[6] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1245 a_4269_918# D[11] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1246 a_7937_297# D[6] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1247 VGND D[5] a_6937_66# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1248 Z a_8379_265# a_7937_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1249 a_117_297# a_559_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1250 Z a_3135_265# a_2693_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1251 a_7937_591# D[14] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1252 a_9513_918# S[15] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1253 Z S[7] a_9513_66# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1254 Z S[6] a_7939_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1255 a_6887_311# D[5] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1256 VPWR S[5] a_6674_325# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1257 a_5361_591# a_5803_793# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1258 VGND D[6] a_7939_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1259 Z S[9] a_1693_918# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1260 a_4219_613# a_4006_599# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1261 Z a_6674_325# a_6887_311# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1262 a_6937_66# D[5] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1263 Z S[10] a_2695_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1264 a_6887_613# D[13] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1265 VPWR D[4] a_5361_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1266 a_1430_599# S[9] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1267 a_5363_911# D[12] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1268 a_2695_911# S[10] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1269 a_117_591# a_559_793# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1270 Z a_3135_793# a_2693_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1271 VPWR D[1] a_1643_311# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1272 a_9513_66# S[7] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1273 Z a_1430_599# a_1643_613# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1274 a_6937_918# D[13] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1275 a_5363_47# D[4] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1276 a_1693_918# D[9] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1277 VPWR D[12] a_5361_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1278 VGND D[15] a_9513_918# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1279 a_9250_599# S[15] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1280 VPWR S[3] a_4006_325# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1281 VGND D[7] a_9513_66# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1282 a_7937_297# D[6] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1283 VGND S[12] a_5803_793# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1284 a_1643_311# a_1430_325# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1285 VPWR D[9] a_1643_613# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1286 Z a_9250_599# a_9463_613# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1287 Z a_4006_325# a_4219_311# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1288 a_1430_325# S[1] VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1289 a_4219_311# D[3] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1290 Z S[13] a_6937_918# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1291 a_4006_325# S[3] VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1292 a_6887_311# a_6674_325# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1293 a_7937_591# D[14] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1294 a_117_297# D[0] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1295 Z a_5803_265# a_5361_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1296 VGND D[11] a_4269_918# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1297 a_4219_613# D[11] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1298 VGND D[13] a_6937_918# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1299 Z a_559_265# a_117_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1300 VGND D[0] a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1301 VPWR D[2] a_2693_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1302 Z S[8] a_119_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1303 a_9463_613# a_9250_599# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1304 a_117_591# D[8] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1305 a_7939_911# D[14] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1306 Z S[2] a_2695_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1307 a_2695_911# D[10] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1308 VPWR S[2] a_3135_265# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1309 VPWR D[10] a_2693_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1310 VGND D[11] a_4269_918# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1311 a_4269_918# D[11] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1312 Z S[12] a_5363_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1313 Z a_4006_599# a_4219_613# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1314 Z a_8379_793# a_7937_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1315 a_1693_66# D[1] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1316 Z S[11] a_4269_918# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1317 a_119_47# D[0] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1318 a_4269_918# S[11] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1319 a_5361_297# D[4] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__ebufn_4 A Z TE_B VNB VPB VGND VPWR
M1000 a_340_309# a_27_47# Z VPB phighvt w=1e+06u l=180000u
+  ad=1.9263e+12p pd=1.369e+07u as=5.8e+11p ps=5.16e+06u
M1001 Z a_27_47# a_413_47# VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=1.053e+12p ps=9.74e+06u
M1002 a_413_47# a_224_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.2475e+11p ps=6.13e+06u
M1003 a_413_47# a_27_47# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Z a_27_47# a_340_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_340_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=9.402e+11p ps=7.71e+06u
M1006 VGND a_224_47# a_413_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1008 VPWR TE_B a_340_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_224_47# TE_B VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=0p ps=0u
M1010 Z a_27_47# a_413_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_340_309# a_27_47# Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_340_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Z a_27_47# a_340_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_413_47# a_224_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_224_47# a_413_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR TE_B a_340_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_224_47# TE_B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1018 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1019 a_413_47# a_27_47# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__clkmux2_1 VGND VPWR S A1 A0 X VPB VNB
M1000 a_245_47# S VGND VNB nshort w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=4.76e+11p ps=4.08e+06u
M1001 a_478_47# A0 a_79_21# VNB nshort w=420000u l=150000u
+  ad=3.591e+11p pd=2.55e+06u as=2.121e+11p ps=1.85e+06u
M1002 a_79_21# A1 a_245_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=8.058e+11p pd=5.56e+06u as=2.7e+11p ps=2.54e+06u
M1004 a_599_309# A1 a_79_21# VPB phighvt w=940000u l=180000u
+  ad=2.444e+11p pd=2.4e+06u as=9.447e+11p ps=3.89e+06u
M1005 a_243_309# S VPWR VPB phighvt w=940000u l=180000u
+  ad=3.901e+11p pd=2.71e+06u as=0p ps=0u
M1006 a_649_21# S VPWR VPB phighvt w=940000u l=180000u
+  ad=2.726e+11p pd=2.46e+06u as=0p ps=0u
M1007 a_649_21# S VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1008 VGND a_649_21# a_478_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_79_21# A0 a_243_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_649_21# a_599_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_79_21# X VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
.ends
.subckt sky130_fd_sc_hdll__o21ai_1 VGND VPWR A2 A1 B1 Y VPB VNB
M1000 VPWR B1 Y VPB phighvt w=700000u l=180000u
+  ad=6.515e+11p pd=5.03e+06u as=3.72e+11p ps=2.84e+06u
M1001 Y A2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.3e+11p ps=2.46e+06u
M1002 a_117_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=3.8025e+11p pd=2.47e+06u as=3.77e+11p ps=3.76e+06u
M1004 a_27_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.535e+11p ps=2.08e+06u
M1005 VGND A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a222oi_1 VNB VPB VGND VPWR C2 C1 B1 A2 A1 Y B2
M1000 a_357_297# B1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=8.3e+11p pd=7.66e+06u as=5.8e+11p ps=5.16e+06u
M1001 Y C2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1002 VGND C2 a_119_47# VNB nshort w=640000u l=150000u
+  ad=9.28e+11p pd=5.46e+06u as=1.344e+11p ps=1.7e+06u
M1003 Y B1 a_449_47# VNB nshort w=640000u l=150000u
+  ad=4.416e+11p pd=3.94e+06u as=1.344e+11p ps=1.7e+06u
M1004 a_117_297# B2 a_357_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_627_47# A1 Y VNB nshort w=640000u l=150000u
+  ad=2.432e+11p pd=2.04e+06u as=0p ps=0u
M1006 a_117_297# C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_357_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.5e+11p ps=2.7e+06u
M1008 VGND A2 a_627_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_357_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_449_47# B2 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_119_47# C1 Y VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__diode_6 VNB VPB VGND VPWR DIODE
D0 VNB DIODE ndiode p=1.47e+07u a=2.2032e+12p
.ends
.subckt sky130_fd_sc_hdll__clkinv_16 Y A VGND VPWR VNB VPB
M1000 Y A VGND VNB nshort w=420000u l=150000u
+  ad=1.1739e+12p pd=1.231e+07u as=1.2285e+12p ps=1.341e+07u
M1001 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=3.895e+12p pd=3.379e+07u as=3.755e+12p ps=3.151e+07u
M1002 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a21o_2 X B1 A1 A2 VNB VPB VGND VPWR
M1000 a_444_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.7e+11p pd=5.14e+06u as=9.35e+11p ps=7.87e+06u
M1001 VPWR A1 a_444_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 X a_80_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.5e+11p pd=2.7e+06u as=0p ps=0u
M1003 X a_80_21# VGND VNB nshort w=650000u l=150000u
+  ad=2.795e+11p pd=2.16e+06u as=8.5475e+11p ps=6.53e+06u
M1004 a_444_297# B1 a_80_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.25e+11p ps=2.65e+06u
M1005 VPWR a_80_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_80_21# B1 VGND VNB nshort w=650000u l=150000u
+  ad=3.185e+11p pd=2.28e+06u as=0p ps=0u
M1007 VGND a_80_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_532_47# A1 a_80_21# VNB nshort w=650000u l=150000u
+  ad=2.3725e+11p pd=2.03e+06u as=0p ps=0u
M1009 VGND A2 a_532_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a211o_2 X A2 A1 B1 C1 VNB VPB VGND VPWR
M1000 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=9.4e+11p pd=7.88e+06u as=2.9e+11p ps=2.58e+06u
M1001 a_643_297# B1 a_319_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.3e+11p pd=2.46e+06u as=6.8e+11p ps=5.36e+06u
M1002 VGND B1 a_79_21# VNB nshort w=650000u l=150000u
+  ad=1.027e+12p pd=7.06e+06u as=4.5825e+11p ps=4.01e+06u
M1003 a_421_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=1.5925e+11p pd=1.79e+06u as=0p ps=0u
M1004 a_319_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_79_21# C1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A2 a_319_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.145e+11p ps=1.96e+06u
M1009 a_79_21# C1 a_643_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1010 a_79_21# A1 a_421_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor4bb_1 A C_N D_N B Y VNB VPB VGND VPWR
M1000 VGND C_N a_27_410# VNB nshort w=420000u l=150000u
+  ad=7.674e+11p pd=7.31e+06u as=1.302e+11p ps=1.46e+06u
M1001 Y B VGND VNB nshort w=650000u l=150000u
+  ad=3.9e+11p pd=3.8e+06u as=0p ps=0u
M1002 a_216_93# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.281e+11p pd=1.45e+06u as=0p ps=0u
M1003 Y a_216_93# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_422_297# a_216_93# Y VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=2.7e+11p ps=2.54e+06u
M1006 VGND a_27_410# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_622_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.23625e+11p pd=5.22e+06u as=2.9e+11p ps=2.58e+06u
M1008 VPWR C_N a_27_410# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1009 a_216_93# D_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1010 a_622_297# B a_518_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.4e+11p ps=2.68e+06u
M1011 a_518_297# a_27_410# a_422_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__isobufsrc_1 A X SLEEP VPB VNB VGND VPWR
M1000 VGND a_74_47# X VNB nshort w=650000u l=150000u
+  ad=4.23e+11p pd=3.99e+06u as=2.08e+11p ps=1.94e+06u
M1001 a_283_297# SLEEP VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.3e+11p pd=2.46e+06u as=3.288e+11p ps=2.82e+06u
M1002 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_74_47# a_283_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1004 VGND A a_74_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1005 VPWR A a_74_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
.ends
.subckt sky130_fd_sc_hdll__or4_4 B C A D X VNB VPB VPWR VGND
M1000 X a_32_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=9.7e+11p ps=7.94e+06u
M1001 a_332_297# B a_238_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u
M1002 X a_32_297# VGND VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=1.07575e+12p ps=9.81e+06u
M1003 VGND A a_32_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.55e+11p ps=4e+06u
M1004 VGND a_32_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_32_297# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C a_32_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_32_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_238_297# C a_122_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=4e+11p ps=2.8e+06u
M1009 VPWR a_32_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A a_332_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_32_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_32_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_32_297# D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_122_297# D a_32_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1015 VPWR a_32_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor4_6 A C D B Y VPB VNB VGND VPWR
M1000 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=8.7e+11p pd=7.74e+06u as=2.01e+12p ps=1.802e+07u
M1001 a_1263_297# C a_685_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.02e+12p pd=1.804e+07u as=1.74e+12p ps=1.548e+07u
M1002 Y D a_1263_297# VPB phighvt w=1e+06u l=180000u
+  ad=8.7e+11p pd=7.74e+06u as=0p ps=0u
M1003 VGND B Y VNB nshort w=650000u l=150000u
+  ad=3.419e+12p pd=2.742e+07u as=2.106e+12p ps=2.208e+07u
M1004 Y D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_685_297# C a_1263_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_297# B a_685_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_685_297# C a_1263_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1263_297# C a_685_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_685_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1263_297# D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND D Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_297# B a_685_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1263_297# D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y D a_1263_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y D a_1263_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Y D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_27_297# B a_685_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_685_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1263_297# D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_685_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND D Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_685_297# C a_1263_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1044 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_1263_297# C a_685_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1046 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VGND D Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and4bb_4 C A_N D X B_N VNB VPB VGND VPWR
M1000 a_606_47# D VGND VNB nshort w=650000u l=150000u
+  ad=2.6975e+11p pd=2.13e+06u as=8.552e+11p ps=7.75e+06u
M1001 a_912_21# A_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=1.9814e+12p ps=1.503e+07u
M1002 VPWR B_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1003 a_184_21# a_912_21# a_836_47# VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=2.47e+11p ps=2.06e+06u
M1004 a_184_21# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=7.35e+11p pd=5.47e+06u as=0p ps=0u
M1005 VGND a_184_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1006 VPWR C a_184_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_184_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_184_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1009 a_836_47# a_27_47# a_719_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.8275e+11p ps=2.17e+06u
M1010 X a_184_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_184_21# D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_912_21# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1013 VPWR a_184_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND B_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1015 VGND a_184_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_184_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_719_47# C a_606_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_912_21# a_184_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_184_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__einvp_2 A Z TE VGND VPWR VPB VNB
M1000 Z A a_214_47# VNB nshort w=650000u l=150000u
+  ad=2.405e+11p pd=2.04e+06u as=6.0775e+11p ps=5.77e+06u
M1001 VPWR a_27_47# a_235_309# VPB phighvt w=940000u l=180000u
+  ad=4.454e+11p pd=4.28e+06u as=9.587e+11p ps=7.84e+06u
M1002 VPWR TE a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1003 a_235_309# A Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1004 VGND TE a_214_47# VNB nshort w=650000u l=150000u
+  ad=4.1e+11p pd=3.95e+06u as=0p ps=0u
M1005 a_214_47# TE VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_214_47# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Z A a_235_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND TE a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1009 a_235_309# a_27_47# VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a221oi_1 Y C1 A1 A2 B2 B1 VGND VPWR VPB VNB
M1000 a_211_297# B2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=6.4e+11p pd=5.28e+06u as=5.6e+11p ps=5.12e+06u
M1001 VPWR A2 a_211_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
M1002 a_225_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=1.365e+11p pd=1.72e+06u as=4.3225e+11p ps=3.93e+06u
M1003 Y B1 a_225_47# VNB nshort w=650000u l=150000u
+  ad=6.045e+11p pd=5.76e+06u as=0p ps=0u
M1004 VGND A2 a_505_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.47e+11p ps=2.06e+06u
M1005 a_505_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_117_297# C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1007 a_211_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND C1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_117_297# B1 a_211_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__buf_8 A X VGND VPWR VPB VNB
M1000 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=1.72e+12p ps=1.544e+07u
M1001 a_27_47# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
M1002 a_27_47# A VGND VNB nshort w=650000u l=150000u
+  ad=4.095e+11p pd=3.86e+06u as=1.1765e+12p ps=1.142e+07u
M1003 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=8.645e+11p pd=7.86e+06u as=0p ps=0u
M1005 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__inv_8 A Y VNB VPB VGND VPWR
M1000 Y A VGND VNB nshort w=650000u l=150000u
+  ad=8.645e+11p pd=7.86e+06u as=9.62e+11p ps=9.46e+06u
M1001 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=1.41e+12p ps=1.282e+07u
M1002 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o22a_1 A2 X B1 A1 B2 VPB VNB VGND VPWR
M1000 VGND A2 a_219_47# VNB nshort w=650000u l=150000u
+  ad=3.835e+11p pd=3.78e+06u as=6.565e+11p ps=5.92e+06u
M1001 VPWR a_83_21# X VPB phighvt w=1e+06u l=180000u
+  ad=9.8e+11p pd=5.96e+06u as=2.9e+11p ps=2.58e+06u
M1002 VPWR A1 a_511_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3e+11p ps=2.6e+06u
M1003 a_83_21# B2 a_299_297# VPB phighvt w=1e+06u l=180000u
+  ad=4.1e+11p pd=2.82e+06u as=2.9e+11p ps=2.58e+06u
M1004 a_219_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_299_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_83_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.82e+11p ps=1.86e+06u
M1007 a_511_297# A2 a_83_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_83_21# B1 a_219_47# VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1009 a_219_47# B2 a_83_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__inputiso0p_1 X SLEEP A VGND VPWR VPB VNB
M1000 VGND A a_307_47# VNB nshort w=420000u l=150000u
+  ad=4.197e+11p pd=3.81e+06u as=8.82e+10p ps=1.26e+06u
M1001 VPWR SLEEP a_27_413# VPB phighvt w=420000u l=180000u
+  ad=6.233e+11p pd=5.09e+06u as=1.134e+11p ps=1.38e+06u
M1002 VPWR A a_211_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1003 X a_211_413# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1004 X a_211_413# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1005 a_27_413# SLEEP VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1006 a_211_413# a_27_413# VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_307_47# a_27_413# a_211_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
.ends
.subckt sky130_fd_sc_hdll__nand3b_4 A_N Y B C VNB VPB VGND VPWR
M1000 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.74e+12p pd=1.548e+07u as=2.61e+12p ps=2.322e+07u
M1001 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_225_47# B a_683_47# VNB nshort w=650000u l=150000u
+  ad=9.62e+11p pd=9.46e+06u as=8.645e+11p ps=7.86e+06u
M1004 a_683_47# B a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_225_47# a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1006 Y a_27_47# a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A_N a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1008 a_225_47# a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND C a_683_47# VNB nshort w=650000u l=150000u
+  ad=8.45e+11p pd=7.8e+06u as=0p ps=0u
M1012 a_683_47# C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_225_47# B a_683_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y a_27_47# a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND C a_683_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_683_47# C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A_N a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1024 a_683_47# B a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor3_1 C Y A B VPB VNB VGND VPWR
M1000 a_211_297# B a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u
M1001 Y B VGND VNB nshort w=650000u l=150000u
+  ad=3.77e+11p pd=3.76e+06u as=6.305e+11p ps=4.54e+06u
M1002 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_117_297# C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1004 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A a_211_297# VPB phighvt w=1e+06u l=180000u
+  ad=6.1e+11p pd=3.22e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand4bb_2 D C B_N A_N Y VNB VPB VGND VPWR
M1000 a_211_413# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.974e+11p pd=1.78e+06u as=3.424e+11p ps=3.42e+06u
M1001 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=2.0218e+12p ps=1.522e+07u
M1002 VPWR B_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1003 a_361_47# a_211_413# Y VNB nshort w=650000u l=150000u
+  ad=5.785e+11p pd=5.68e+06u as=2.08e+11p ps=1.94e+06u
M1004 Y a_211_413# a_361_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_841_47# D VGND VNB nshort w=650000u l=150000u
+  ad=5.59e+11p pd=5.62e+06u as=0p ps=0u
M1007 Y a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND D a_841_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_211_413# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_841_47# C a_641_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1012 VGND B_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1013 a_211_413# A_N VPWR VPB phighvt w=420000u l=180000u
+  ad=2.016e+11p pd=1.8e+06u as=0p ps=0u
M1014 Y a_211_413# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_361_47# a_27_47# a_641_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_641_47# a_27_47# a_361_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_641_47# C a_841_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__muxb16to1_2 Z VGND VPWR VNB VPB D[2] D[1] S[7] S[6] S[5]
+ D[9] D[8] S[14] S[13] S[12] S[11] S[10] S[9] S[8] D[15] D[14] D[13] D[12] D[11]
+ D[10] S[15] S[4] S[3] S[2] S[1] S[0] D[7] D[6] D[5] D[4] D[3] D[0]
M1000 a_2603_911# S[12] Z VNB nshort w=520000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=2.2464e+12p ps=2.528e+07u
M1001 VPWR S[4] a_2854_265# VPB phighvt w=1e+06u l=180000u
+  ad=7.52e+12p pd=6.304e+07u as=2.7e+11p ps=2.54e+06u
M1002 VPWR D[3] a_2112_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.211e+11p ps=7.41e+06u
M1003 VPWR D[2] a_1315_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.211e+11p ps=7.41e+06u
M1004 Z a_1989_47# a_2112_333# VPB phighvt w=820000u l=180000u
+  ad=3.8048e+12p pd=3.552e+07u as=0p ps=0u
M1005 Z a_1566_265# a_1315_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Z a_4142_793# a_3891_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=8.211e+11p ps=7.41e+06u
M1007 VPWR S[12] a_2854_793# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1008 VPWR D[11] a_2112_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.211e+11p ps=7.41e+06u
M1009 VPWR D[10] a_1315_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.211e+11p ps=7.41e+06u
M1010 a_27_297# D[0] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1011 a_2133_915# D[11] VGND VNB nshort w=650000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=3.9312e+12p ps=4.208e+07u
M1012 VGND S[14] a_4142_793# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1013 a_27_297# a_278_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_591# D[8] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1015 Z S[10] a_1315_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=5.6745e+11p ps=5.52e+06u
M1016 a_3421_915# S[13] Z VNB nshort w=520000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1017 a_4565_47# S[7] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1018 VGND D[14] a_3891_911# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=5.6745e+11p ps=5.52e+06u
M1019 a_1989_47# S[3] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1020 a_27_911# S[8] Z VNB nshort w=520000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1021 a_3891_911# S[14] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Z S[5] a_3421_69# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=5.6745e+11p ps=5.52e+06u
M1023 VPWR S[0] a_278_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1024 a_4709_69# D[7] VGND VNB nshort w=650000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1025 a_2133_69# D[3] VGND VNB nshort w=650000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1026 VGND D[9] a_845_915# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=5.6745e+11p ps=5.52e+06u
M1027 VPWR S[8] a_278_793# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1028 a_845_69# S[1] Z VNB nshort w=520000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1029 Z S[11] a_2133_915# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_2603_297# D[4] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1031 Z a_278_265# a_27_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_27_47# S[0] Z VNB nshort w=520000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1033 VGND S[10] a_1566_793# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1034 a_2603_297# a_2854_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1315_911# D[10] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Z a_701_937# a_824_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=8.211e+11p ps=7.41e+06u
M1037 Z S[1] a_845_69# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_2603_591# D[12] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1039 a_701_937# S[9] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1040 a_4565_937# S[15] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1041 Z S[0] a_27_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_27_47# D[0] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_1315_911# S[10] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_1315_591# a_1566_793# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_2112_591# a_1989_937# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1046 Z S[4] a_2603_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=5.6745e+11p ps=5.52e+06u
M1047 VGND D[8] a_27_911# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 Z S[9] a_845_915# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_4688_591# a_4565_937# Z VPB phighvt w=820000u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1050 VGND D[7] a_4709_69# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1051 a_3400_333# D[5] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1052 a_824_333# D[1] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1053 a_1989_47# S[3] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1054 a_3421_69# S[5] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1055 a_3400_333# a_3277_47# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1056 a_824_591# D[9] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1057 VGND D[4] a_2603_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1058 a_3400_591# D[13] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1059 a_845_915# D[9] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1060 a_1989_937# S[11] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1061 a_4688_333# D[7] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1062 a_3891_297# D[6] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1063 VGND S[12] a_2854_793# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1064 VGND S[4] a_2854_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1065 a_3277_47# S[5] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1066 a_3891_297# a_4142_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1067 a_2133_915# S[11] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1068 a_4688_591# D[15] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1069 a_3891_591# D[14] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1070 a_3277_937# S[13] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1071 a_1989_937# S[11] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1072 a_701_47# S[1] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1073 VGND D[12] a_2603_911# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1074 VGND D[1] a_845_69# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1075 VPWR D[0] a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1076 Z a_4565_937# a_4688_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1077 VPWR S[6] a_4142_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1078 VPWR D[8] a_27_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1079 VPWR D[5] a_3400_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1080 VPWR D[4] a_2603_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1081 VGND S[0] a_278_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1082 Z a_3277_47# a_3400_333# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1083 Z a_2854_265# a_2603_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1084 a_824_333# a_701_47# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1085 VPWR S[14] a_4142_793# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1086 a_2603_47# S[4] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1087 VPWR D[13] a_3400_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1088 VPWR D[12] a_2603_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1089 a_701_47# S[1] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1090 VGND D[5] a_3421_69# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1091 Z a_4142_265# a_3891_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1092 a_701_937# S[9] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1093 Z a_1989_937# a_2112_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1094 a_2603_47# D[4] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1095 Z a_1566_793# a_1315_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1096 a_3277_937# S[13] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1097 VPWR D[1] a_824_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1098 a_3277_47# S[5] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1099 a_27_591# a_278_793# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1100 VGND D[13] a_3421_915# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1101 VPWR D[9] a_824_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1102 Z S[3] a_2133_69# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1103 a_2603_911# D[12] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1104 Z S[8] a_27_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1105 a_845_69# D[1] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1106 Z S[15] a_4709_915# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=5.6745e+11p ps=5.52e+06u
M1107 Z S[7] a_4709_69# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1108 VGND D[0] a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1109 VGND D[10] a_1315_911# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1110 a_3421_69# D[5] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1111 Z a_278_793# a_27_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1112 Z S[6] a_3891_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=5.6745e+11p ps=5.52e+06u
M1113 Z a_701_47# a_824_333# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1114 a_2603_591# a_2854_793# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1115 VGND S[8] a_278_793# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1116 Z S[2] a_1315_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=5.6745e+11p ps=5.52e+06u
M1117 a_1315_47# D[2] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1118 a_27_911# D[8] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1119 a_3891_911# D[14] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1120 a_1315_297# D[2] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1121 a_3421_915# D[13] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1122 a_4688_333# a_4565_47# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1123 a_2112_333# a_1989_47# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1124 a_1315_297# a_1566_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1125 a_2133_69# S[3] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1126 a_1315_591# D[10] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1127 VGND D[2] a_1315_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1128 Z S[12] a_2603_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1129 a_4565_47# S[7] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1130 a_845_915# S[9] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1131 a_4709_915# S[15] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1132 a_4565_937# S[15] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1133 VPWR S[2] a_1566_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1134 a_3400_591# a_3277_937# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1135 a_2112_333# D[3] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1136 VGND D[11] a_2133_915# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1137 VPWR S[10] a_1566_793# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1138 a_4709_69# S[7] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1139 VGND D[6] a_3891_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1140 a_3891_591# a_4142_793# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1141 a_2112_591# D[11] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1142 VPWR D[7] a_4688_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1143 VPWR D[6] a_3891_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1144 VGND S[6] a_4142_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1145 a_3891_47# S[6] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1146 Z S[13] a_3421_915# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1147 a_4709_915# D[15] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1148 Z a_4565_47# a_4688_333# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1149 VPWR D[15] a_4688_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1150 VGND S[2] a_1566_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1151 a_1315_47# S[2] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1152 VPWR D[14] a_3891_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1153 Z S[14] a_3891_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1154 VGND D[15] a_4709_915# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1155 a_3891_47# D[6] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1156 VGND D[3] a_2133_69# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1157 a_824_591# a_701_937# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1158 Z a_3277_937# a_3400_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1159 Z a_2854_793# a_2603_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__ebufn_2 Z A TE_B VNB VPB VGND VPWR
M1000 VPWR A a_27_47# VPB phighvt w=640000u l=180000u
+  ad=5.254e+11p pd=4.53e+06u as=1.728e+11p ps=1.82e+06u
M1001 VGND a_224_47# a_412_47# VNB nshort w=650000u l=150000u
+  ad=3.54e+11p pd=3.53e+06u as=6.8575e+11p ps=6.01e+06u
M1002 a_224_47# TE_B VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1003 a_340_309# a_27_47# Z VPB phighvt w=1e+06u l=180000u
+  ad=1.3537e+12p pd=8.63e+06u as=2.9e+11p ps=2.58e+06u
M1004 a_412_47# a_224_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_412_47# a_27_47# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.405e+11p ps=2.04e+06u
M1006 a_224_47# TE_B VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1007 a_340_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR TE_B a_340_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Z a_27_47# a_340_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1011 Z a_27_47# a_412_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__diode_4 DIODE VGND VPWR VPB VNB
D0 VNB DIODE ndiode p=9.88e+06u a=1.0557e+12p
.ends
.subckt sky130_fd_sc_hdll__and3_1 VGND VPWR X B A C VPB VNB
M1000 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=4.548e+11p ps=4.26e+06u
M1001 a_213_47# B a_119_47# VNB nshort w=420000u l=150000u
+  ad=2.247e+11p pd=1.91e+06u as=1.344e+11p ps=1.48e+06u
M1002 VPWR A a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=3.255e+11p ps=3.23e+06u
M1003 VGND C a_213_47# VNB nshort w=420000u l=150000u
+  ad=2.58e+11p pd=2.2e+06u as=0p ps=0u
M1004 VPWR C a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1006 a_119_47# A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1007 a_27_47# B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__clkbuf_1 VGND VPWR X A VPB VNB w_233_n17#
M1000 VPWR a_75_212# X VPB phighvt w=790000u l=180000u
+  ad=5.293e+11p pd=2.92e+06u as=2.133e+11p ps=2.12e+06u
M1001 a_75_212# A VGND w_233_n17# nshort w=520000u l=150000u
+  ad=1.404e+11p pd=1.58e+06u as=3.38e+11p ps=2.34e+06u
M1002 a_75_212# A VPWR VPB phighvt w=790000u l=180000u
+  ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1003 VGND a_75_212# X w_233_n17# nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.612e+11p ps=1.66e+06u
.ends
.subckt sky130_fd_sc_hdll__clkinv_1 Y A VPB VNB VGND VPWR
M1000 VGND A Y VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.323e+11p ps=1.47e+06u
M1001 Y A VPWR VPB phighvt w=840000u l=180000u
+  ad=2.436e+11p pd=2.26e+06u as=4.704e+11p ps=4.48e+06u
M1002 VPWR A Y VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sdfstp_1 SCE SET_B VPWR VGND CLK D SCD Q VPB VNB
M1000 VPWR SET_B a_1229_21# VPB phighvt w=420000u l=180000u
+  ad=1.5997e+12p pd=1.544e+07u as=1.722e+11p ps=1.66e+06u
M1001 VGND a_349_21# a_295_47# VNB nshort w=420000u l=150000u
+  ad=1.2848e+12p pd=1.309e+07u as=1.134e+11p ps=1.38e+06u
M1002 Q a_2381_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1003 a_1955_47# a_693_369# a_1725_329# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.482e+11p ps=2.2e+06u
M1004 VPWR a_1725_329# a_2381_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1005 VGND SCE a_349_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1006 a_1075_413# a_877_369# a_201_47# VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=2.99e+11p ps=3.24e+06u
M1007 a_1725_329# a_877_369# a_1645_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=5.056e+11p ps=2.86e+06u
M1008 VPWR SCD a_27_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=3.456e+11p ps=3.64e+06u
M1009 a_1229_21# a_1075_413# VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1841_413# a_877_369# a_1725_329# VPB phighvt w=420000u l=180000u
+  ad=1.722e+11p pd=1.66e+06u as=3.906e+11p ps=3.86e+06u
M1011 a_1725_329# SET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR SCE a_349_21# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1013 a_1725_329# a_693_369# a_1643_329# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=1.932e+11p ps=2.14e+06u
M1014 a_1921_295# a_1725_329# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1015 a_877_369# a_693_369# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1016 VGND a_1229_21# a_1177_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1017 VGND CLK a_693_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1018 a_1645_47# a_1075_413# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_1921_295# a_1841_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1467_47# a_1075_413# a_1229_21# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.512e+11p ps=1.56e+06u
M1021 a_27_369# a_349_21# a_201_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_119_47# SCD VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1023 a_1177_47# a_877_369# a_1075_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1024 VGND SET_B a_1467_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_877_369# a_693_369# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1026 a_1075_413# a_693_369# a_201_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.646e+11p ps=2.94e+06u
M1027 a_2027_47# a_1921_295# a_1955_47# VNB nshort w=420000u l=150000u
+  ad=1.596e+11p pd=1.6e+06u as=0p ps=0u
M1028 a_1643_329# a_1075_413# VPWR VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_295_47# D a_201_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_201_47# SCE a_119_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND SET_B a_2027_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND a_1725_329# a_2381_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1033 a_211_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=1.472e+11p pd=1.74e+06u as=0p ps=0u
M1034 a_1921_295# a_1725_329# VGND VNB nshort w=420000u l=150000u
+  ad=1.596e+11p pd=1.6e+06u as=0p ps=0u
M1035 Q a_2381_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1036 a_201_47# D a_211_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1169_413# a_693_369# a_1075_413# VPB phighvt w=420000u l=180000u
+  ad=1.596e+11p pd=1.6e+06u as=0p ps=0u
M1038 VPWR a_1229_21# a_1169_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR CLK a_693_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
.ends
.subckt sky130_fd_sc_hdll__dfstp_4 Q D VPWR CLK VGND VPB VNB SET_B
M1000 VPWR SET_B a_1126_413# VPB phighvt w=420000u l=180000u
+  ad=1.9683e+12p pd=1.875e+07u as=2.856e+11p ps=3.04e+06u
M1001 Q a_1738_47# VGND VNB nshort w=650000u l=150000u
+  ad=5.85e+11p pd=5.7e+06u as=1.5993e+12p ps=1.487e+07u
M1002 a_211_363# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1003 a_506_47# a_27_47# a_409_329# VNB nshort w=360000u l=150000u
+  ad=1.8e+11p pd=1.72e+06u as=1.87e+11p ps=1.93e+06u
M1004 Q a_1738_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.5e+11p pd=7.7e+06u as=0p ps=0u
M1005 a_1344_47# a_27_47# a_1126_413# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.596e+11p ps=1.6e+06u
M1006 VGND a_1126_413# a_1738_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1007 VPWR CLK a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1008 VPWR a_1738_47# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_1126_413# a_1738_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1010 VPWR a_702_21# a_610_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.974e+11p ps=1.78e+06u
M1011 VPWR a_1288_261# a_1244_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=9.66e+10p ps=1.3e+06u
M1012 a_1126_413# a_211_363# a_1156_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1013 a_1044_413# a_506_47# VPWR VPB phighvt w=420000u l=180000u
+  ad=9.66e+10p pd=1.3e+06u as=0p ps=0u
M1014 Q a_1738_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_1738_47# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Q a_1738_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_409_329# D VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Q a_1738_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_409_329# D VPWR VPB phighvt w=840000u l=180000u
+  ad=2.625e+11p pd=2.39e+06u as=0p ps=0u
M1020 a_1156_47# a_506_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_636_47# a_211_363# a_506_47# VNB nshort w=360000u l=150000u
+  ad=1.341e+11p pd=1.5e+06u as=0p ps=0u
M1022 VPWR a_506_47# a_702_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1023 a_1288_261# a_1126_413# VPWR VPB phighvt w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1024 a_610_413# a_27_47# a_506_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1025 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1026 a_866_47# SET_B VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1027 VGND a_702_21# a_636_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1288_261# a_1126_413# VGND VNB nshort w=540000u l=150000u
+  ad=1.404e+11p pd=1.6e+06u as=0p ps=0u
M1029 a_1244_413# a_211_363# a_1126_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_702_21# a_506_47# a_866_47# VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1031 a_702_21# SET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_211_363# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1033 a_506_47# a_211_363# a_409_329# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1416_47# a_1288_261# a_1344_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1035 a_1126_413# a_27_47# a_1044_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR a_1738_47# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND SET_B a_1416_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 Q a_1738_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND a_1738_47# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or4_2 B C A X D VPWR VGND VPB VNB
M1000 a_27_297# D VGND VNB nshort w=420000u l=150000u
+  ad=2.94e+11p pd=3.08e+06u as=6.666e+11p ps=6.83e+06u
M1001 VGND A a_27_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 X a_27_297# VGND VNB nshort w=650000u l=150000u
+  ad=3.4775e+11p pd=2.37e+06u as=0p ps=0u
M1003 a_117_297# D a_27_297# VPB phighvt w=420000u l=180000u
+  ad=1.47e+11p pd=1.54e+06u as=1.134e+11p ps=1.38e+06u
M1004 VPWR A a_305_297# VPB phighvt w=420000u l=180000u
+  ad=6.257e+11p pd=5.35e+06u as=1.47e+11p ps=1.54e+06u
M1005 a_27_297# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C a_27_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_27_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=4.55e+11p ps=2.91e+06u
M1008 VGND a_27_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_27_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_223_297# C a_117_297# VPB phighvt w=420000u l=180000u
+  ad=9.66e+10p pd=1.3e+06u as=0p ps=0u
M1011 a_305_297# B a_223_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sdfsbp_2 Q_N Q CLK D SCD SCE SET_B VGND VPWR VPB VNB
M1000 VGND a_349_21# a_295_47# VNB nshort w=420000u l=150000u
+  ad=1.90535e+12p pd=1.891e+07u as=1.134e+11p ps=1.38e+06u
M1001 a_1930_295# a_1735_329# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1002 a_1930_295# a_1735_329# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=2.6255e+12p ps=2.377e+07u
M1003 a_1075_413# a_877_369# a_199_47# VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=2.99e+11p ps=3.24e+06u
M1004 VGND SCE a_349_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1005 a_1735_329# a_877_369# a_1655_47# VNB nshort w=640000u l=150000u
+  ad=3.054e+11p pd=2.42e+06u as=4.736e+11p ps=2.76e+06u
M1006 Q a_2739_47# VGND VNB nshort w=650000u l=150000u
+  ad=2.08e+11p pd=1.94e+06u as=0p ps=0u
M1007 VPWR SCD a_27_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=3.456e+11p ps=3.64e+06u
M1008 a_1219_21# a_1075_413# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.701e+11p pd=1.65e+06u as=0p ps=0u
M1009 a_1870_413# a_877_369# a_1735_329# VPB phighvt w=420000u l=180000u
+  ad=1.302e+11p pd=1.46e+06u as=4.305e+11p ps=4.05e+06u
M1010 a_1655_47# a_1075_413# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR SCE a_349_21# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1012 a_1735_329# a_693_369# a_1652_329# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=1.974e+11p ps=2.15e+06u
M1013 a_1735_329# SET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_2739_47# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1015 VGND a_1735_329# Q_N VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1016 VPWR a_1735_329# a_2739_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1017 VGND CLK a_693_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1018 a_877_369# a_693_369# VGND VNB nshort w=420000u l=150000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
M1019 VPWR a_1735_329# Q_N VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1020 VPWR a_1930_295# a_1870_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1467_47# a_1075_413# a_1219_21# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.512e+11p ps=1.56e+06u
M1022 a_27_369# a_349_21# a_199_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR SET_B a_1219_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1177_47# a_877_369# a_1075_413# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.344e+11p ps=1.48e+06u
M1025 VGND SET_B a_1467_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Q a_2739_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_877_369# a_693_369# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1028 a_199_47# SCE a_109_47# VNB nshort w=420000u l=150000u
+  ad=2.688e+11p pd=2.96e+06u as=1.26e+11p ps=1.44e+06u
M1029 VGND a_1219_21# a_1177_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Q_N a_1735_329# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1075_413# a_693_369# a_199_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_295_47# D a_199_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND a_1735_329# a_2739_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1034 VGND a_2739_47# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1652_329# a_1075_413# VPWR VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_211_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=1.472e+11p pd=1.74e+06u as=0p ps=0u
M1037 Q_N a_1735_329# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_109_47# SCD VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_2049_47# a_1930_295# a_1977_47# VNB nshort w=420000u l=150000u
+  ad=2.688e+11p pd=2.12e+06u as=8.82e+10p ps=1.26e+06u
M1040 a_199_47# D a_211_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1169_413# a_693_369# a_1075_413# VPB phighvt w=420000u l=180000u
+  ad=1.596e+11p pd=1.6e+06u as=0p ps=0u
M1042 VPWR a_1219_21# a_1169_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VGND SET_B a_2049_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VPWR CLK a_693_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1045 a_1977_47# a_693_369# a_1735_329# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a21boi_1 Y A1 B1_N A2 VPWR VGND VPB VNB
M1000 VPWR B1_N a_27_413# VPB phighvt w=420000u l=180000u
+  ad=5.355e+11p pd=4.23e+06u as=1.155e+11p ps=1.39e+06u
M1001 VPWR A1 a_338_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.75e+11p ps=5.15e+06u
M1002 VGND B1_N a_27_413# VNB nshort w=420000u l=150000u
+  ad=4.345e+11p pd=3.99e+06u as=1.533e+11p ps=1.57e+06u
M1003 a_434_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=2.665e+11p pd=2.12e+06u as=3.51e+11p ps=2.38e+06u
M1004 VGND A2 a_434_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y a_27_413# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_338_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_338_297# a_27_413# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.25e+11p ps=2.65e+06u
.ends
.subckt sky130_fd_sc_hdll__and4bb_2 VNB VPB VGND VPWR A_N C B_N X D
M1000 a_503_47# a_27_47# a_184_21# VNB nshort w=420000u l=150000u
+  ad=1.449e+11p pd=1.53e+06u as=1.092e+11p ps=1.36e+06u
M1001 VPWR D a_184_21# VPB phighvt w=420000u l=180000u
+  ad=1.299e+12p pd=9.38e+06u as=2.562e+11p ps=2.9e+06u
M1002 VPWR A_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1003 a_184_21# C VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_602_47# a_545_280# a_503_47# VNB nshort w=420000u l=150000u
+  ad=1.407e+11p pd=1.51e+06u as=0p ps=0u
M1005 VGND D a_699_47# VNB nshort w=420000u l=150000u
+  ad=6.1255e+11p pd=5.76e+06u as=1.134e+11p ps=1.38e+06u
M1006 a_699_47# C a_602_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_545_280# B_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1008 a_184_21# a_27_47# VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_545_280# a_184_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_184_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1011 VGND A_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1012 VGND a_184_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1013 X a_184_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_545_280# B_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1015 X a_184_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand3_1 Y A C B VPB VNB VGND VPWR
M1000 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=6.2e+11p pd=5.24e+06u as=5.6e+11p ps=5.12e+06u
M1001 a_203_47# B a_119_47# VNB nshort w=650000u l=150000u
+  ad=2.47e+11p pd=2.06e+06u as=1.755e+11p ps=1.84e+06u
M1002 Y A a_203_47# VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=0p ps=0u
M1003 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_119_47# C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
.ends
.subckt sky130_fd_sc_hdll__nor4_4 A C Y D B VPB VNB VGND VPWR
M1000 a_497_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=1.43e+12p ps=1.286e+07u
M1001 a_887_297# D Y VPB phighvt w=1e+06u l=180000u
+  ad=1.41e+12p pd=1.282e+07u as=5.8e+11p ps=5.16e+06u
M1002 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1003 VGND A Y VNB nshort w=650000u l=150000u
+  ad=2.0475e+12p pd=1.8e+07u as=1.794e+12p ps=1.592e+07u
M1004 a_497_297# C a_887_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND D Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y D a_887_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_887_297# D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_887_297# C a_497_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_297# B a_497_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_497_297# C a_887_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_497_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND D Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_887_297# C a_497_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_27_297# B a_497_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y D a_887_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__mux2_1 VGND VPWR S A1 A0 X VPB VNB
M1000 a_245_47# S VGND VNB nshort w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=4.745e+11p ps=4.06e+06u
M1001 VGND a_657_21# a_499_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.318e+11p ps=2.42e+06u
M1002 a_79_21# A0 a_243_374# VPB phighvt w=420000u l=180000u
+  ad=4.515e+11p pd=2.99e+06u as=1.743e+11p ps=1.67e+06u
M1003 a_613_374# A1 a_79_21# VPB phighvt w=420000u l=180000u
+  ad=9.66e+10p pd=1.3e+06u as=0p ps=0u
M1004 a_79_21# A1 a_245_47# VNB nshort w=420000u l=150000u
+  ad=2.562e+11p pd=2.06e+06u as=0p ps=0u
M1005 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=4.926e+11p pd=4.44e+06u as=2.7e+11p ps=2.54e+06u
M1006 VPWR a_657_21# a_613_374# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_499_47# A0 a_79_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_657_21# S VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1009 a_243_374# S VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1011 a_657_21# S VPWR VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and2b_1 X A_N B VGND VPWR VPB VNB
M1000 VPWR A_N a_27_413# VPB phighvt w=420000u l=180000u
+  ad=6.422e+11p pd=5.18e+06u as=1.134e+11p ps=1.38e+06u
M1001 VGND B a_327_47# VNB nshort w=420000u l=150000u
+  ad=3.653e+11p pd=3.54e+06u as=1.218e+11p ps=1.42e+06u
M1002 a_225_413# a_27_413# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1003 a_327_47# a_27_413# a_225_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1004 X a_225_413# VGND VNB nshort w=650000u l=150000u
+  ad=1.95e+11p pd=1.9e+06u as=0p ps=0u
M1005 X a_225_413# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.1e+11p pd=2.62e+06u as=0p ps=0u
M1006 a_27_413# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1007 VPWR B a_225_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__buf_6 VPWR VGND X A VPB VNB
M1000 VGND a_169_297# X VNB nshort w=650000u l=150000u
+  ad=9.62e+11p pd=9.46e+06u as=6.565e+11p ps=5.92e+06u
M1001 VPWR A a_169_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.41e+12p pd=1.282e+07u as=2.9e+11p ps=2.58e+06u
M1002 a_169_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR a_169_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.7e+11p ps=7.74e+06u
M1004 X a_169_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_169_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_169_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A a_169_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1008 VPWR a_169_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_169_297# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_169_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_169_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_169_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_169_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_169_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_169_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__inv_16 Y A VPB VNB VGND VPWR
M1000 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=2.57e+12p pd=2.314e+07u as=2.32e+12p ps=2.064e+07u
M1001 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VGND VNB nshort w=650000u l=150000u
+  ad=1.664e+12p pd=1.552e+07u as=1.8265e+12p ps=1.732e+07u
M1005 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__inv_6 Y A VPB VNB VPWR VGND
M1000 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=1.13e+12p pd=1.026e+07u as=8.7e+11p ps=7.74e+06u
M1001 VGND A Y VNB nshort w=650000u l=150000u
+  ad=7.605e+11p pd=7.54e+06u as=6.24e+11p ps=5.82e+06u
M1002 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand3b_2 Y C A_N B VNB VPB VGND VPWR
M1000 VGND C a_228_47# VNB nshort w=650000u l=150000u
+  ad=4.295e+11p pd=4.01e+06u as=4.485e+11p ps=3.98e+06u
M1001 Y a_27_47# a_448_47# VNB nshort w=650000u l=150000u
+  ad=2.405e+11p pd=2.04e+06u as=5.46e+11p ps=5.58e+06u
M1002 VPWR A_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=1.4657e+12p pd=1.303e+07u as=1.134e+11p ps=1.38e+06u
M1003 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.7e+11p pd=7.74e+06u as=0p ps=0u
M1004 a_448_47# B a_228_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_228_47# B a_448_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_228_47# C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_448_47# a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
.ends
.subckt sky130_fd_sc_hdll__sdfrtp_1 VPB VNB VGND VPWR RESET_B Q CLK D SCD SCE
M1000 a_1428_47# a_1380_303# a_1322_47# VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.518e+11p ps=1.6e+06u
M1001 a_213_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=1.3533e+12p ps=1.268e+07u
M1002 VPWR a_1972_21# a_1951_413# VPB phighvt w=420000u l=180000u
+  ad=1.6398e+12p pd=1.569e+07u as=1.386e+11p ps=1.5e+06u
M1003 a_1972_21# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=1.344e+11p pd=1.48e+06u as=0p ps=0u
M1004 Q a_1972_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.15e+11p pd=2.63e+06u as=0p ps=0u
M1005 a_2157_47# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=0p ps=0u
M1006 VPWR SCD a_870_389# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=1.971e+11p ps=1.81e+06u
M1007 a_700_389# D a_631_119# VNB nshort w=420000u l=150000u
+  ad=3.3215e+11p pd=3.47e+06u as=1.302e+11p ps=1.46e+06u
M1008 a_1380_303# a_1202_413# VPWR VPB phighvt w=840000u l=180000u
+  ad=2.541e+11p pd=2.37e+06u as=0p ps=0u
M1009 a_1202_413# a_27_47# a_700_389# VNB nshort w=360000u l=150000u
+  ad=1.44e+11p pd=1.52e+06u as=0p ps=0u
M1010 VPWR a_1757_47# a_1972_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1972_21# a_1757_47# a_2157_47# VNB nshort w=420000u l=150000u
+  ad=1.365e+11p pd=1.49e+06u as=0p ps=0u
M1012 Q a_1972_21# VGND VNB nshort w=650000u l=150000u
+  ad=1.9825e+11p pd=1.91e+06u as=0p ps=0u
M1013 VPWR a_1380_303# a_1324_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1014 VPWR CLK a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1015 a_618_389# SCE VPWR VPB phighvt w=540000u l=180000u
+  ad=1.242e+11p pd=1.54e+06u as=0p ps=0u
M1016 a_1951_413# a_213_47# a_1757_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1017 a_700_389# D a_618_389# VPB phighvt w=540000u l=180000u
+  ad=5.193e+11p pd=4.01e+06u as=0p ps=0u
M1018 a_631_119# a_331_66# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND RESET_B a_1428_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1324_413# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1202_413# a_213_47# a_700_389# VPB phighvt w=420000u l=180000u
+  ad=1.806e+11p pd=1.7e+06u as=0p ps=0u
M1022 a_1324_413# a_27_47# a_1202_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1866_47# a_27_47# a_1757_47# VNB nshort w=360000u l=150000u
+  ad=2.121e+11p pd=1.9e+06u as=1.422e+11p ps=1.51e+06u
M1024 a_1757_47# a_213_47# a_1380_303# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.87e+11p ps=1.93e+06u
M1025 VPWR SCE a_331_66# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=2.214e+11p ps=1.9e+06u
M1026 VGND CLK a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1027 VGND a_1972_21# a_1866_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_213_47# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
M1029 a_899_66# SCE a_700_389# VNB nshort w=420000u l=500000u
+  ad=1.554e+11p pd=1.58e+06u as=0p ps=0u
M1030 a_1757_47# a_27_47# a_1380_303# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1322_47# a_213_47# a_1202_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND SCD a_899_66# VNB nshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_870_389# a_331_66# a_700_389# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND SCE a_331_66# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1035 a_1380_303# a_1202_413# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__dfrtp_4 Q D CLK VGND VPWR RESET_B VPB VNB
M1000 a_699_413# a_27_47# a_583_47# VPB phighvt w=420000u l=180000u
+  ad=3.528e+11p pd=3.36e+06u as=1.533e+11p ps=1.57e+06u
M1001 a_865_47# a_811_289# a_689_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=3.012e+11p ps=2.3e+06u
M1002 a_211_363# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.5815e+12p ps=1.392e+07u
M1003 VGND RESET_B a_865_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR CLK a_27_47# VPB phighvt w=640000u l=180000u
+  ad=1.8817e+12p pd=1.792e+07u as=1.728e+11p ps=1.82e+06u
M1005 a_1188_47# a_211_363# a_811_289# VNB nshort w=360000u l=150000u
+  ad=1.782e+11p pd=1.71e+06u as=1.998e+11p ps=1.97e+06u
M1006 VPWR a_1403_21# a_1388_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.428e+11p ps=1.52e+06u
M1007 a_583_47# a_27_47# a_468_47# VNB nshort w=360000u l=150000u
+  ad=1.368e+11p pd=1.48e+06u as=1.71e+11p ps=1.69e+06u
M1008 VGND a_1403_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1009 a_1388_413# a_211_363# a_1188_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1010 VPWR a_1403_21# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1011 VPWR a_1188_47# a_1403_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1012 a_468_47# D VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1403_21# a_1188_47# a_1612_47# VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.491e+11p ps=1.55e+06u
M1014 a_689_47# a_211_363# a_583_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_811_289# a_699_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Q a_1403_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1403_21# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_1403_21# a_1317_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.728e+11p ps=1.7e+06u
M1019 VPWR a_1403_21# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1317_47# a_27_47# a_1188_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1022 a_811_289# a_583_47# VPWR VPB phighvt w=840000u l=180000u
+  ad=2.709e+11p pd=2.41e+06u as=0p ps=0u
M1023 Q a_1403_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_468_47# D VPWR VPB phighvt w=420000u l=180000u
+  ad=1.386e+11p pd=1.5e+06u as=0p ps=0u
M1025 a_583_47# a_211_363# a_468_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Q a_1403_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_211_363# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1028 a_1188_47# a_27_47# a_811_289# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1612_47# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND a_1403_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Q a_1403_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_811_289# a_583_47# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_699_413# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__isobufsrc_16 A X SLEEP VPB VNB VGND VPWR
M1000 X SLEEP a_585_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.32e+12p pd=2.064e+07u as=4.92e+12p ps=4.384e+07u
M1001 VPWR A a_151_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.27e+12p pd=2.854e+07u as=6.8e+11p ps=5.36e+06u
M1002 X a_151_297# VGND VNB nshort w=650000u l=150000u
+  ad=3.393e+12p pd=3.124e+07u as=4.095e+12p ps=3.73e+07u
M1003 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X SLEEP a_585_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_151_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_151_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_151_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_151_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_151_297# a_585_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_151_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_585_297# a_151_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_585_297# a_151_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_585_297# SLEEP X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_151_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_151_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_585_297# SLEEP X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_151_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND SLEEP X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_151_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND SLEEP X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_585_297# a_151_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_151_297# a_585_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_585_297# SLEEP X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X SLEEP a_585_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_151_297# a_585_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR a_151_297# a_585_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_151_297# A VGND VNB nshort w=650000u l=150000u
+  ad=5.135e+11p pd=4.18e+06u as=0p ps=0u
M1029 VGND SLEEP X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_585_297# SLEEP X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_585_297# a_151_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 X SLEEP a_585_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND SLEEP X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 X SLEEP a_585_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND a_151_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_151_297# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR a_151_297# a_585_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 X a_151_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 X a_151_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPWR a_151_297# a_585_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_585_297# SLEEP X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_585_297# SLEEP X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VGND SLEEP X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 VGND SLEEP X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VPWR A a_151_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_585_297# a_151_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1049 X SLEEP a_585_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1050 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1051 X SLEEP a_585_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1052 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1053 X a_151_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1054 a_151_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1055 VGND a_151_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1056 a_585_297# a_151_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1057 a_585_297# a_151_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1058 X SLEEP a_585_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1059 VGND A a_151_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1060 VGND a_151_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1061 VGND a_151_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1062 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1063 a_585_297# a_151_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1064 a_585_297# SLEEP X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1065 VGND SLEEP X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1066 VPWR a_151_297# a_585_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1067 VPWR a_151_297# a_585_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1068 a_585_297# SLEEP X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1069 VGND A a_151_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1070 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1071 VGND SLEEP X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sdlclkp_4 SCE GATE GCLK VGND VPWR CLK VPB VNB
M1000 a_425_47# a_277_243# a_310_47# VNB nshort w=360000u l=150000u
+  ad=2.196e+11p pd=1.96e+06u as=1.53e+11p ps=1.57e+06u
M1001 a_27_47# GATE VGND VNB nshort w=420000u l=150000u
+  ad=2.664e+11p pd=2.97e+06u as=1.3078e+12p ps=1.141e+07u
M1002 a_27_47# GATE a_117_369# VPB phighvt w=640000u l=180000u
+  ad=2.373e+11p pd=2.08e+06u as=1.472e+11p ps=1.74e+06u
M1003 GCLK a_1125_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=7.15e+11p pd=5.43e+06u as=2.2235e+12p ps=1.837e+07u
M1004 GCLK a_1125_47# VGND VNB nshort w=650000u l=150000u
+  ad=5.3625e+11p pd=4.25e+06u as=0p ps=0u
M1005 a_421_413# a_280_21# a_310_47# VPB phighvt w=420000u l=180000u
+  ad=1.806e+11p pd=1.7e+06u as=1.47e+11p ps=1.54e+06u
M1006 a_280_21# CLK VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1007 a_117_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_280_21# a_277_243# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1009 VPWR CLK a_1125_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1010 VPWR a_505_315# a_421_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1125_47# a_505_315# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_310_47# a_277_243# a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_280_21# a_277_243# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1014 VGND a_1125_47# GCLK VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_505_315# a_425_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND SCE a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 GCLK a_1125_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1217_47# a_505_315# a_1125_47# VNB nshort w=650000u l=150000u
+  ad=1.365e+11p pd=1.72e+06u as=2.015e+11p ps=1.92e+06u
M1019 a_505_315# a_310_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1020 VPWR a_1125_47# GCLK VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND CLK a_1217_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 GCLK a_1125_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_280_21# CLK VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1024 VGND a_1125_47# GCLK VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_1125_47# GCLK VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_310_47# a_280_21# a_27_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_505_315# a_310_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sdfrbp_2 VPB VNB VPWR VGND RESET_B Q_N Q SCD SCE CLK D
M1000 a_1428_47# a_1380_303# a_1322_47# VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.518e+11p ps=1.6e+06u
M1001 a_213_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=1.77805e+12p ps=1.664e+07u
M1002 VPWR a_1972_21# a_1951_413# VPB phighvt w=420000u l=180000u
+  ad=2.2692e+12p pd=2.101e+07u as=1.386e+11p ps=1.5e+06u
M1003 a_1972_21# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=1.344e+11p pd=1.48e+06u as=0p ps=0u
M1004 Q_N a_2372_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=0p ps=0u
M1005 a_2157_47# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=0p ps=0u
M1006 VPWR SCD a_870_389# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=1.971e+11p ps=1.81e+06u
M1007 a_700_389# D a_631_119# VNB nshort w=420000u l=150000u
+  ad=3.3215e+11p pd=3.47e+06u as=1.302e+11p ps=1.46e+06u
M1008 a_1380_303# a_1202_413# VPWR VPB phighvt w=840000u l=180000u
+  ad=2.541e+11p pd=2.37e+06u as=0p ps=0u
M1009 a_1202_413# a_27_47# a_700_389# VNB nshort w=360000u l=150000u
+  ad=1.44e+11p pd=1.52e+06u as=0p ps=0u
M1010 VPWR a_1757_47# a_1972_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1972_21# a_1757_47# a_2157_47# VNB nshort w=420000u l=150000u
+  ad=1.365e+11p pd=1.49e+06u as=0p ps=0u
M1012 VPWR a_1380_303# a_1324_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1013 VPWR CLK a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1014 a_618_389# SCE VPWR VPB phighvt w=540000u l=180000u
+  ad=1.242e+11p pd=1.54e+06u as=0p ps=0u
M1015 Q a_1972_21# VGND VNB nshort w=650000u l=150000u
+  ad=2.34e+11p pd=2.02e+06u as=0p ps=0u
M1016 a_1951_413# a_213_47# a_1757_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1017 a_700_389# D a_618_389# VPB phighvt w=540000u l=180000u
+  ad=5.193e+11p pd=4.01e+06u as=0p ps=0u
M1018 a_631_119# a_331_66# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_1972_21# a_2372_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1020 VGND RESET_B a_1428_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_1972_21# a_2372_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1022 a_1324_413# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1202_413# a_213_47# a_700_389# VPB phighvt w=420000u l=180000u
+  ad=1.806e+11p pd=1.7e+06u as=0p ps=0u
M1024 a_1324_413# a_27_47# a_1202_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1866_47# a_27_47# a_1757_47# VNB nshort w=360000u l=150000u
+  ad=2.121e+11p pd=1.9e+06u as=1.422e+11p ps=1.51e+06u
M1026 a_1757_47# a_213_47# a_1380_303# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.87e+11p ps=1.93e+06u
M1027 Q_N a_2372_47# VGND VNB nshort w=650000u l=150000u
+  ad=2.0475e+11p pd=1.93e+06u as=0p ps=0u
M1028 VPWR SCE a_331_66# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=2.214e+11p ps=1.9e+06u
M1029 VGND CLK a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1030 VGND a_1972_21# a_1866_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND a_1972_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Q a_1972_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.3e+11p pd=2.66e+06u as=0p ps=0u
M1033 VPWR a_1972_21# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_213_47# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
M1035 a_899_66# SCE a_700_389# VNB nshort w=420000u l=500000u
+  ad=1.554e+11p pd=1.58e+06u as=0p ps=0u
M1036 a_1757_47# a_27_47# a_1380_303# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1322_47# a_213_47# a_1202_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND a_2372_47# Q_N VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR a_2372_47# Q_N VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND SCD a_899_66# VNB nshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_870_389# a_331_66# a_700_389# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VGND SCE a_331_66# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1043 a_1380_303# a_1202_413# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or3b_1 A C_N X B VGND VPWR VPB VNB
M1000 a_225_53# B VGND VNB nshort w=420000u l=150000u
+  ad=2.835e+11p pd=3.03e+06u as=4.787e+11p ps=4.92e+06u
M1001 VGND A a_225_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND a_117_297# a_225_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_117_297# C_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=4.241e+11p ps=4.1e+06u
M1004 VPWR A a_399_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.407e+11p ps=1.51e+06u
M1005 a_399_297# B a_315_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 a_117_297# C_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1007 a_315_297# a_117_297# a_225_53# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1008 X a_225_53# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1009 X a_225_53# VGND VNB nshort w=650000u l=150000u
+  ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o32ai_1 A2 Y A1 A3 B2 B1 VPB VNB VGND VPWR
M1000 VPWR A1 a_465_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.6e+11p pd=5.12e+06u as=2.9e+11p ps=2.58e+06u
M1001 VGND A3 a_27_47# VNB nshort w=650000u l=150000u
+  ad=6.0125e+11p pd=4.45e+06u as=5.655e+11p ps=5.64e+06u
M1002 Y B2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.15e+11p pd=3.03e+06u as=2.3e+11p ps=2.46e+06u
M1003 a_117_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_465_297# A2 a_338_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=4.55e+11p ps=2.91e+06u
M1005 a_27_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.4375e+11p ps=2.05e+06u
M1006 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_338_297# A3 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__xor2_1 B X A VNB VPB VPWR VGND
M1000 VPWR A a_125_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.6e+11p pd=5.12e+06u as=3e+11p ps=2.6e+06u
M1001 X a_35_297# a_315_297# VPB phighvt w=1e+06u l=180000u
+  ad=4.5e+11p pd=2.9e+06u as=5.7e+11p ps=5.14e+06u
M1002 a_35_297# B VGND VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=7.28e+11p ps=6.14e+06u
M1003 VGND A a_35_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_35_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=5.46e+11p ps=2.98e+06u
M1005 VPWR B a_315_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_125_297# B a_35_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1007 a_317_47# A VGND VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=0p ps=0u
M1008 X B a_317_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_315_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o21ba_1 B1_N A1 X A2 VNB VPB VGND VPWR
M1000 a_79_199# a_222_93# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=9.257e+11p ps=7.95e+06u
M1001 a_222_93# B1_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
M1002 a_222_93# B1_N VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=3.76e+11p ps=3.81e+06u
M1003 a_460_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=4.29e+11p pd=3.92e+06u as=0p ps=0u
M1004 VGND A2 a_460_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_79_199# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1006 VPWR A1 a_554_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1007 VGND a_79_199# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1008 a_554_297# A2 a_79_199# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_460_47# a_222_93# a_79_199# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.95e+11p ps=1.9e+06u
.ends
.subckt sky130_fd_sc_hdll__or4bb_1 A X B D_N C_N VPWR VGND VPB VNB
M1000 X a_331_413# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.85e+11p pd=2.57e+06u as=5.64325e+11p ps=5.4e+06u
M1001 a_609_297# B a_527_297# VPB phighvt w=420000u l=180000u
+  ad=1.281e+11p pd=1.45e+06u as=9.66e+10p ps=1.3e+06u
M1002 a_421_413# a_216_93# a_331_413# VPB phighvt w=420000u l=180000u
+  ad=2.514e+11p pd=2.7e+06u as=1.134e+11p ps=1.38e+06u
M1003 a_216_93# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.281e+11p pd=1.45e+06u as=6.2055e+11p ps=6.43e+06u
M1004 a_331_413# B VGND VNB nshort w=420000u l=150000u
+  ad=2.814e+11p pd=3.02e+06u as=0p ps=0u
M1005 VGND A a_331_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C_N a_27_410# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1007 VGND a_27_410# a_331_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A a_609_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_331_413# VGND VNB nshort w=650000u l=150000u
+  ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u
M1010 a_331_413# a_216_93# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR C_N a_27_410# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1012 a_216_93# D_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
M1013 a_527_297# a_27_410# a_421_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and4_4 X C A B D VNB VPB VGND VPWR
M1000 VPWR D a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=1.51e+12p pd=1.302e+07u as=7.4e+11p ps=5.48e+06u
M1001 a_198_47# B a_119_47# VNB nshort w=650000u l=150000u
+  ad=2.47e+11p pd=2.06e+06u as=1.5925e+11p ps=1.79e+06u
M1002 VPWR B a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_47# C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=6.24e+11p pd=5.82e+06u as=4.485e+11p ps=3.98e+06u
M1005 VGND D a_304_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.1525e+11p ps=2.27e+06u
M1006 a_27_47# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1008 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_119_47# A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1013 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_304_47# C a_198_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o221ai_1 A2 Y B1 C1 A1 B2 VPB VNB VGND VPWR
M1000 Y B2 a_351_297# VPB phighvt w=1e+06u l=180000u
+  ad=7.6e+11p pd=5.52e+06u as=2.6e+11p ps=2.52e+06u
M1001 VPWR C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=1.24e+12p pd=6.48e+06u as=0p ps=0u
M1002 a_569_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=2.3e+11p pd=2.46e+06u as=0p ps=0u
M1003 VPWR A1 a_569_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_123_47# C1 Y VNB nshort w=650000u l=150000u
+  ad=3.77e+11p pd=3.76e+06u as=2.145e+11p ps=1.96e+06u
M1005 a_261_47# B2 a_123_47# VNB nshort w=650000u l=150000u
+  ad=6.695e+11p pd=5.96e+06u as=0p ps=0u
M1006 a_261_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1007 a_123_47# B1 a_261_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2 a_261_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_351_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor3b_1 C_N Y A B VPB VNB VGND VPWR
M1000 a_91_199# C_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=4.62e+11p ps=4.11e+06u
M1001 a_263_297# B a_169_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u
M1002 a_169_297# a_91_199# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.3e+11p ps=2.66e+06u
M1003 a_91_199# C_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=3.057e+11p ps=2.71e+06u
M1004 Y B VGND VNB nshort w=650000u l=150000u
+  ad=4.29e+11p pd=3.92e+06u as=0p ps=0u
M1005 VGND a_91_199# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_263_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__mux2_16 VPWR VGND VPB VNB X S A1 A0
M1000 a_119_47# S VGND VNB nshort w=650000u l=150000u
+  ad=7.02e+11p pd=7.36e+06u as=3.4515e+12p ps=3.012e+07u
M1001 VGND a_973_297# a_1163_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.02e+11p ps=7.36e+06u
M1002 a_27_47# A1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.66e+12p pd=1.532e+07u as=1.16e+12p ps=1.032e+07u
M1003 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=4.27e+12p pd=3.854e+07u as=2.32e+12p ps=2.064e+07u
M1004 a_27_47# A0 a_1163_47# VNB nshort w=650000u l=150000u
+  ad=1.287e+12p pd=1.176e+07u as=0p ps=0u
M1005 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.404e+12p ps=1.472e+07u
M1006 a_117_297# a_973_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR S a_597_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.16e+12p ps=1.032e+07u
M1008 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_597_297# A0 a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1163_47# a_973_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_47# A0 a_597_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1163_47# A0 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR S a_973_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1014 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_597_297# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_47# A1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_597_297# A0 a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND S a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_119_47# S VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_973_297# a_1163_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_117_297# A1 a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR a_973_297# a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_27_47# A0 a_597_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_973_297# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_27_47# A1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_117_297# a_973_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_973_297# S VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1043 VGND S a_973_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_119_47# A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_27_47# A0 a_1163_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 VPWR S a_597_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1048 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1049 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1050 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1051 a_1163_47# a_973_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1052 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1053 a_1163_47# A0 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1054 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1055 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1056 a_117_297# A1 a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1057 VPWR a_973_297# a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1058 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1059 a_27_47# A1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1060 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1061 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1062 VGND S a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1063 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1064 a_597_297# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1065 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1066 a_119_47# A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1067 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand4_4 A D C B Y VPWR VGND VPB VNB
M1000 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=3.15e+12p pd=2.43e+07u as=2.32e+12p ps=2.064e+07u
M1001 VPWR D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_27_47# D VGND VNB nshort w=650000u l=150000u
+  ad=9.62e+11p pd=9.46e+06u as=4.16e+11p ps=3.88e+06u
M1003 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_883_47# B a_485_47# VNB nshort w=650000u l=150000u
+  ad=1.0335e+12p pd=9.68e+06u as=8.645e+11p ps=7.86e+06u
M1006 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_485_47# B a_883_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_883_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1009 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y A a_883_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_47# C a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_883_47# B a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_485_47# C a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_485_47# B a_883_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND D a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_47# D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_883_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_27_47# C a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y A a_883_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_485_47# C a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND D a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__decap_8 VPWR VGND VPB VNB
M1000 VPWR VGND VPWR VPB phighvt w=870000u l=2.89e+06u
+  ad=4.524e+11p pd=4.52e+06u as=0p ps=0u
M1001 VGND VPWR VGND VNB nshort w=550000u l=2.89e+06u
+  ad=2.86e+11p pd=3.24e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE ndiode p=5.36e+06u a=4.347e+11p
.ends
.subckt sky130_fd_sc_hdll__o31ai_1 Y A2 A1 A3 B1 VPB VNB VPWR VGND
M1000 a_117_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=5.4e+11p ps=5.08e+06u
M1001 VGND A2 a_119_47# VNB nshort w=650000u l=150000u
+  ad=3.77e+11p pd=3.76e+06u as=5.33e+11p ps=4.24e+06u
M1002 Y B1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=2.535e+11p pd=2.08e+06u as=0p ps=0u
M1003 Y A3 a_213_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=3.16e+06u as=2.9e+11p ps=2.58e+06u
M1004 a_119_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_119_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_213_297# A2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__clkinv_12 Y A VNB VPB VGND VPWR
M1000 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=2.86e+12p pd=2.572e+07u as=2.61e+12p ps=2.322e+07u
M1001 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A VGND VNB nshort w=420000u l=150000u
+  ad=6.804e+11p pd=8.28e+06u as=1.323e+12p ps=1.218e+07u
M1003 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and3b_4 A_N X C B VNB VPB VGND VPWR
M1000 VGND C a_277_47# VNB nshort w=650000u l=150000u
+  ad=7.285e+11p pd=6.23e+06u as=1.82e+11p ps=1.86e+06u
M1001 VPWR a_56_297# X VPB phighvt w=1e+06u l=180000u
+  ad=1.3907e+12p pd=1.088e+07u as=6.1e+11p ps=5.22e+06u
M1002 X a_56_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR C a_56_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=6.6e+11p ps=5.32e+06u
M1004 X a_56_297# VGND VNB nshort w=650000u l=150000u
+  ad=4.615e+11p pd=4.02e+06u as=0p ps=0u
M1005 VPWR a_98_199# a_56_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_56_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_56_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_56_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_162_47# a_98_199# a_56_297# VNB nshort w=650000u l=150000u
+  ad=2.7625e+11p pd=2.15e+06u as=2.3075e+11p ps=2.01e+06u
M1010 VGND a_56_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_98_199# A_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.239e+11p pd=1.43e+06u as=0p ps=0u
M1012 VPWR a_56_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_98_199# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.743e+11p pd=1.67e+06u as=0p ps=0u
M1014 a_277_47# B a_162_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_56_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__einvn_1 Z A TE_B VGND VPWR VPB VNB
M1000 a_316_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=3.8025e+11p pd=2.47e+06u as=5.255e+11p ps=2.97e+06u
M1001 VPWR TE_B a_27_47# VPB phighvt w=640000u l=180000u
+  ad=3.144e+11p pd=2.69e+06u as=1.728e+11p ps=1.82e+06u
M1002 VGND TE_B a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1003 Z A a_222_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=1.065e+12p ps=4.13e+06u
M1004 a_222_297# TE_B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Z A a_316_47# VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__dfstp_2 Q VGND CLK VPWR D VPB VNB SET_B
M1000 VPWR SET_B a_1126_413# VPB phighvt w=420000u l=180000u
+  ad=1.6789e+12p pd=1.611e+07u as=2.856e+11p ps=3.04e+06u
M1001 VPWR a_1738_47# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1002 a_211_363# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.33055e+12p ps=1.269e+07u
M1003 a_506_47# a_27_47# a_409_329# VNB nshort w=360000u l=150000u
+  ad=1.8e+11p pd=1.72e+06u as=1.87e+11p ps=1.93e+06u
M1004 a_1344_47# a_27_47# a_1126_413# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.596e+11p ps=1.6e+06u
M1005 VGND a_1126_413# a_1738_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1006 VPWR CLK a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1007 VPWR a_702_21# a_610_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.974e+11p ps=1.78e+06u
M1008 Q a_1738_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_1288_261# a_1244_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=9.66e+10p ps=1.3e+06u
M1010 a_1126_413# a_211_363# a_1156_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1011 a_1044_413# a_506_47# VPWR VPB phighvt w=420000u l=180000u
+  ad=9.66e+10p pd=1.3e+06u as=0p ps=0u
M1012 VPWR a_1126_413# a_1738_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1013 a_409_329# D VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_409_329# D VPWR VPB phighvt w=840000u l=180000u
+  ad=2.625e+11p pd=2.39e+06u as=0p ps=0u
M1015 a_1156_47# a_506_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_636_47# a_211_363# a_506_47# VNB nshort w=360000u l=150000u
+  ad=1.341e+11p pd=1.5e+06u as=0p ps=0u
M1017 VPWR a_506_47# a_702_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1018 a_1288_261# a_1126_413# VPWR VPB phighvt w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1019 a_610_413# a_27_47# a_506_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1020 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1021 a_866_47# SET_B VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1022 VGND a_1738_47# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.405e+11p ps=2.04e+06u
M1023 VGND a_702_21# a_636_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1288_261# a_1126_413# VGND VNB nshort w=540000u l=150000u
+  ad=1.404e+11p pd=1.6e+06u as=0p ps=0u
M1025 a_1244_413# a_211_363# a_1126_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_702_21# a_506_47# a_866_47# VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1027 a_702_21# SET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_211_363# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1029 a_506_47# a_211_363# a_409_329# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1416_47# a_1288_261# a_1344_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1031 a_1126_413# a_27_47# a_1044_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND SET_B a_1416_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Q a_1738_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__xnor2_4 Y B A VNB VPB VGND VPWR
M1000 VPWR A a_898_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.32e+12p pd=2.064e+07u as=1.41e+12p ps=1.282e+07u
M1001 Y a_38_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.41e+12p pd=1.282e+07u as=0p ps=0u
M1002 VGND B a_980_47# VNB nshort w=650000u l=150000u
+  ad=1.378e+12p pd=1.334e+07u as=1.443e+12p ps=1.354e+07u
M1003 a_980_47# a_38_297# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.485e+11p ps=3.98e+06u
M1004 VGND A a_980_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_38_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.43e+12p pd=1.286e+07u as=0p ps=0u
M1006 Y B a_898_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_38_297# B a_38_47# VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=9.425e+11p ps=9.4e+06u
M1008 VPWR a_38_297# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_38_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_980_47# a_38_297# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_980_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR B a_38_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_898_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y a_38_297# a_980_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_38_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_38_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_38_297# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A a_898_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A a_38_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_898_297# B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_38_47# B a_38_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_980_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND B a_980_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y a_38_297# a_980_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A a_980_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_898_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_38_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y B a_898_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y a_38_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND A a_38_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_38_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND A a_38_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_980_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR B a_38_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR A a_38_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_898_297# B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_38_297# B a_38_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_38_47# B a_38_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_980_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or4b_4 D_N B C A X VNB VPB VGND VPWR
M1000 VPWR a_225_297# X VPB phighvt w=1e+06u l=180000u
+  ad=1.0734e+12p pd=9.3e+06u as=5.8e+11p ps=5.16e+06u
M1001 VPWR A a_525_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1002 X a_225_297# VGND VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=1.2023e+12p ps=1.127e+07u
M1003 a_117_413# D_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1004 X a_225_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A a_225_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.55e+11p ps=4e+06u
M1006 a_525_297# B a_431_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1007 a_225_297# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_431_297# C a_315_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=4e+11p ps=2.8e+06u
M1009 VPWR a_225_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_225_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_225_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND C a_225_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_117_413# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.0785e+11p pd=1.36e+06u as=0p ps=0u
M1014 a_225_297# a_117_413# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_225_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_225_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_315_297# a_117_413# a_225_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
.ends
.subckt sky130_fd_sc_hdll__a2bb2o_4 X B1 B2 A1_N A2_N VNB VPB VGND VPWR
M1000 a_455_21# A1_N VGND VNB nshort w=650000u l=150000u
+  ad=3.835e+11p pd=3.78e+06u as=1.716e+12p ps=1.438e+07u
M1001 a_27_297# B2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.12e+12p pd=1.024e+07u as=1.7e+12p ps=1.54e+07u
M1002 X a_203_47# VGND VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=0p ps=0u
M1003 X a_203_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1004 VPWR A1_N a_785_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1005 a_27_297# a_455_21# a_203_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1006 a_203_47# B2 a_119_47# VNB nshort w=650000u l=150000u
+  ad=4.81e+11p pd=4.08e+06u as=3.835e+11p ps=3.78e+06u
M1007 VGND a_203_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_203_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A1_N a_455_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_203_47# a_455_21# a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_203_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_785_297# A2_N a_455_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1014 VGND a_455_21# a_203_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_203_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_455_21# A2_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_119_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND B1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_455_21# A2_N a_785_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_203_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_203_47# a_455_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_203_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A2_N a_455_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_785_297# A1_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_119_47# B2 a_203_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor4_2 C D Y A B VNB VPB VGND VPWR
M1000 a_309_297# C a_515_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=8.5e+11p ps=7.7e+06u
M1001 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u
M1002 VGND C Y VNB nshort w=650000u l=150000u
+  ad=1.066e+12p pd=1.108e+07u as=9.62e+11p ps=8.16e+06u
M1003 a_27_297# B a_309_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_309_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_515_297# D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1009 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y D a_515_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND D Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_515_297# C a_309_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__xor3_4 X C B A VNB VPB VGND VPWR
M1000 VPWR a_80_207# X VPB phighvt w=1e+06u l=180000u
+  ad=1.4908e+12p pd=1.305e+07u as=5.8e+11p ps=5.16e+06u
M1001 a_658_49# a_528_297# a_80_207# VPB phighvt w=840000u l=180000u
+  ad=7.558e+11p pd=5.2e+06u as=3.36e+11p ps=2.48e+06u
M1002 VGND a_80_207# X VNB nshort w=650000u l=150000u
+  ad=1.2254e+12p pd=1.035e+07u as=4.16e+11p ps=3.88e+06u
M1003 a_658_49# B a_1225_365# VNB nshort w=640000u l=150000u
+  ad=5.931e+11p pd=4.52e+06u as=4.468e+11p ps=3.98e+06u
M1004 a_1109_297# B VGND VNB nshort w=650000u l=150000u
+  ad=1.653e+11p pd=1.82e+06u as=0p ps=0u
M1005 a_80_207# C a_658_49# VNB nshort w=640000u l=150000u
+  ad=2.88e+11p pd=2.18e+06u as=0p ps=0u
M1006 a_1225_365# a_1109_297# a_658_49# VPB phighvt w=840000u l=180000u
+  ad=7.234e+11p pd=5.3e+06u as=0p ps=0u
M1007 a_80_207# C a_652_325# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=7.32e+11p ps=5.16e+06u
M1008 a_658_49# B a_1510_297# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=7.748e+11p ps=5.63e+06u
M1009 VPWR A a_1225_365# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1510_297# a_1225_365# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_80_207# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_80_207# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_652_325# a_528_297# a_80_207# VNB nshort w=640000u l=150000u
+  ad=6.6045e+11p pd=4.67e+06u as=0p ps=0u
M1014 a_1510_297# a_1109_297# a_652_325# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A a_1225_365# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_80_207# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_80_207# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_652_325# B a_1225_365# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_80_207# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_528_297# C VPWR VPB phighvt w=640000u l=180000u
+  ad=2.112e+11p pd=1.94e+06u as=0p ps=0u
M1021 a_1510_297# a_1109_297# a_658_49# VNB nshort w=420000u l=150000u
+  ad=5.517e+11p pd=4.37e+06u as=0p ps=0u
M1022 a_1109_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.126e+11p pd=2.64e+06u as=0p ps=0u
M1023 a_528_297# C VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1024 a_1510_297# a_1225_365# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 X a_80_207# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_652_325# B a_1510_297# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1225_365# a_1109_297# a_652_325# VNB nshort w=600000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__dlrtp_4 RESET_B D GATE Q VGND VPWR VPB VNB
M1000 Q a_750_21# VGND VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=1.00625e+12p ps=1.01e+07u
M1001 VGND a_750_21# a_708_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1002 Q a_750_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=1.691e+12p ps=1.487e+07u
M1003 VPWR GATE a_27_363# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1004 VPWR a_750_21# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_203_47# a_27_363# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1006 VPWR a_750_21# a_702_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1007 VGND a_750_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_503_369# a_319_369# VPWR VPB phighvt w=640000u l=180000u
+  ad=2.021e+11p pd=1.97e+06u as=0p ps=0u
M1009 a_708_47# a_27_363# a_604_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.58e+06u
M1010 Q a_750_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Q a_750_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND D a_319_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1013 VPWR D a_319_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1014 VGND RESET_B a_981_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.6575e+11p ps=1.81e+06u
M1015 a_604_47# a_203_47# a_500_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.58e+06u
M1016 VPWR RESET_B a_750_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1017 a_981_47# a_604_47# a_750_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1018 VGND GATE a_27_363# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1019 a_702_413# a_203_47# a_604_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1020 a_203_47# a_27_363# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1021 a_604_47# a_27_363# a_503_369# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_750_21# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_500_47# a_319_369# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_750_21# a_604_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_750_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__isobufsrc_8 A X SLEEP VPB VNB VGND VPWR
M1000 VPWR a_117_297# a_345_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.76e+12p pd=1.552e+07u as=2.6e+12p ps=2.32e+07u
M1001 VPWR A a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.4e+11p ps=2.68e+06u
M1002 a_345_297# a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_345_297# SLEEP X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.16e+12p ps=1.032e+07u
M1004 a_345_297# a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_117_297# a_345_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=1.729e+12p pd=1.572e+07u as=2.249e+12p ps=1.992e+07u
M1007 X SLEEP a_345_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND SLEEP X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND SLEEP X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_117_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_345_297# a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_345_297# SLEEP X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_117_297# a_345_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A a_117_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1019 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X SLEEP a_345_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND SLEEP X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_345_297# a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_345_297# SLEEP X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_117_297# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_345_297# SLEEP X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR a_117_297# a_345_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND SLEEP X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 X SLEEP a_345_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 X SLEEP a_345_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a32o_1 X A3 B2 B1 A1 A2 VGND VPWR VPB VNB
M1000 a_276_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=1.95e+11p pd=1.9e+06u as=6.045e+11p ps=4.46e+06u
M1001 VPWR a_93_21# X VPB phighvt w=1e+06u l=180000u
+  ad=9.75e+11p pd=5.95e+06u as=3.4e+11p ps=2.68e+06u
M1002 a_93_21# B1 a_268_297# VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=1.015e+12p ps=8.03e+06u
M1003 a_93_21# A1 a_366_47# VNB nshort w=650000u l=150000u
+  ad=3.185e+11p pd=2.28e+06u as=3.575e+11p ps=2.4e+06u
M1004 a_366_47# A2 a_276_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_93_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.145e+11p ps=1.96e+06u
M1006 a_634_47# B1 a_93_21# VNB nshort w=650000u l=150000u
+  ad=1.365e+11p pd=1.72e+06u as=0p ps=0u
M1007 VPWR A2 a_268_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_268_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_268_297# A3 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_268_297# B2 a_93_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B2 a_634_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__buf_4 VPWR VGND X A VPB VNB
M1000 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=8.5e+11p ps=7.7e+06u
M1001 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=4.16e+11p pd=3.88e+06u as=5.85e+11p ps=5.7e+06u
M1002 VPWR A a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1003 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1007 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__inv_4 Y A VPB VNB VPWR VGND
M1000 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=1.075e+12p pd=8.15e+06u as=5.8e+11p ps=5.16e+06u
M1001 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A VGND VNB nshort w=650000u l=150000u
+  ad=4.16e+11p pd=3.88e+06u as=7.3775e+11p ps=6.17e+06u
M1003 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__dfrtp_2 RESET_B VPWR VGND Q CLK D VPB VNB
M1000 a_436_413# D VPWR VPB phighvt w=420000u l=180000u
+  ad=1.428e+11p pd=1.52e+06u as=1.5845e+12p ps=1.543e+07u
M1001 VPWR a_1323_21# a_1330_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=9.66e+10p ps=1.3e+06u
M1002 VPWR a_1323_21# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1003 a_211_363# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.3154e+12p ps=1.178e+07u
M1004 a_649_413# a_27_47# a_534_47# VPB phighvt w=420000u l=180000u
+  ad=3.318e+11p pd=3.26e+06u as=1.533e+11p ps=1.57e+06u
M1005 a_805_47# a_751_289# a_642_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.748e+11p ps=2.17e+06u
M1006 VPWR CLK a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1007 VGND RESET_B a_805_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_436_413# D VGND VNB nshort w=420000u l=150000u
+  ad=1.338e+11p pd=1.5e+06u as=0p ps=0u
M1009 VGND a_1323_21# a_1237_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.698e+11p ps=1.7e+06u
M1010 VPWR a_751_289# a_649_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_751_289# a_534_47# VGND VNB nshort w=640000u l=150000u
+  ad=1.998e+11p pd=1.97e+06u as=0p ps=0u
M1012 Q a_1323_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_1128_47# a_1323_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1014 a_1128_47# a_211_363# a_751_289# VNB nshort w=360000u l=150000u
+  ad=1.422e+11p pd=1.51e+06u as=0p ps=0u
M1015 a_534_47# a_27_47# a_436_413# VNB nshort w=360000u l=150000u
+  ad=1.404e+11p pd=1.5e+06u as=0p ps=0u
M1016 Q a_1323_21# VGND VNB nshort w=650000u l=150000u
+  ad=2.405e+11p pd=2.04e+06u as=0p ps=0u
M1017 a_751_289# a_534_47# VPWR VPB phighvt w=840000u l=180000u
+  ad=2.709e+11p pd=2.41e+06u as=0p ps=0u
M1018 a_1128_47# a_27_47# a_751_289# VPB phighvt w=420000u l=180000u
+  ad=1.512e+11p pd=1.56e+06u as=0p ps=0u
M1019 a_642_47# a_211_363# a_534_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1237_47# a_27_47# a_1128_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1542_47# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=1.596e+11p pd=1.6e+06u as=0p ps=0u
M1022 a_1323_21# a_1128_47# a_1542_47# VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1023 a_649_413# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1025 a_1323_21# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_1323_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_211_363# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1028 a_534_47# a_211_363# a_436_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1330_413# a_211_363# a_1128_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor4b_4 B A D_N C Y VPB VNB VGND VPWR
M1000 a_27_297# B a_493_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.41e+12p pd=1.282e+07u as=1.16e+12p ps=1.032e+07u
M1001 VGND a_1311_21# Y VNB nshort w=650000u l=150000u
+  ad=2.2815e+12p pd=2.002e+07u as=1.7615e+12p ps=1.582e+07u
M1002 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.7e+11p ps=7.74e+06u
M1003 Y a_1311_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_493_297# C a_883_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.41e+12p ps=1.282e+07u
M1005 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_493_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_883_297# C a_493_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_297# B a_493_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y a_1311_21# a_883_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1013 VPWR D_N a_1311_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1014 VGND a_1311_21# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_493_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_883_297# a_1311_21# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_493_297# C a_883_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y a_1311_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y a_1311_21# a_883_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_883_297# a_1311_21# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND D_N a_1311_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1028 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_883_297# C a_493_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a211oi_4 A2 A1 C1 Y B1 VPWR VGND VNB VPB
M1000 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.99e+12p pd=1.798e+07u as=1.16e+12p ps=1.032e+07u
M1001 VGND C1 Y VNB nshort w=650000u l=150000u
+  ad=1.404e+12p pd=1.342e+07u as=1.365e+12p ps=1.2e+07u
M1002 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND A2 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.995e+11p ps=7.66e+06u
M1004 Y C1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_869_297# C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=6.2e+11p ps=5.24e+06u
M1007 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1057_297# B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.2e+11p pd=2.64e+06u as=0p ps=0u
M1010 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A2 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_119_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND C1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y C1 a_1057_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_297# B1 a_869_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y C1 a_869_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_119_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y C1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_869_297# B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y A1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1449_297# C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=3.3e+11p pd=2.66e+06u as=0p ps=0u
M1027 a_27_297# B1 a_1449_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_119_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y A1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_119_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sdlclkp_2 CLK VPWR VGND GCLK SCE GATE VPB VNB
M1000 a_484_315# a_299_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=1.6654e+12p ps=1.474e+07u
M1001 a_269_21# CLK VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1002 a_27_47# GATE a_117_369# VPB phighvt w=640000u l=180000u
+  ad=2.021e+11p pd=1.97e+06u as=1.472e+11p ps=1.74e+06u
M1003 VPWR a_1093_47# GCLK VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1004 a_1185_47# a_484_315# a_1093_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.302e+11p ps=1.46e+06u
M1005 VGND CLK a_1185_47# VNB nshort w=420000u l=150000u
+  ad=9.4605e+11p pd=9.05e+06u as=0p ps=0u
M1006 a_484_315# a_299_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1007 a_117_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_415_47# a_266_243# a_299_47# VNB nshort w=360000u l=150000u
+  ad=1.977e+11p pd=1.85e+06u as=1.548e+11p ps=1.58e+06u
M1009 a_410_413# a_269_21# a_299_47# VPB phighvt w=420000u l=180000u
+  ad=1.596e+11p pd=1.6e+06u as=1.47e+11p ps=1.54e+06u
M1010 VPWR a_484_315# a_410_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 GCLK a_1093_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_1093_47# GCLK VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1013 VPWR CLK a_1093_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.856e+11p ps=1.86e+06u
M1014 GCLK a_1093_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_484_315# a_415_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_269_21# CLK VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1017 VGND a_269_21# a_266_243# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1018 a_299_47# a_269_21# a_27_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=2.622e+11p ps=2.95e+06u
M1019 a_1093_47# a_484_315# VPWR VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND SCE a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_299_47# a_266_243# a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_269_21# a_266_243# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1023 a_27_47# GATE VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a22oi_1 B1 A1 B2 A2 Y VPWR VGND VPB VNB
M1000 Y B1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=5.8e+11p ps=5.16e+06u
M1001 Y B1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=3.77e+11p pd=3.76e+06u as=1.755e+11p ps=1.84e+06u
M1002 a_117_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_411_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1004 VPWR A2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1005 a_117_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2 a_411_47# VNB nshort w=650000u l=150000u
+  ad=4.29e+11p pd=3.92e+06u as=0p ps=0u
M1007 a_119_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__muxb4to1_1 S[0] D[0] D[1] S[1] S[2] D[2] D[3] S[3] VPB
+ VNB VGND VPWR Z
M1000 a_937_47# D[2] VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=9.997e+11p ps=9.4e+06u
M1001 a_1361_47# S[3] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=1.69e+12p ps=1.338e+07u
M1002 a_1574_47# S[3] Z VNB nshort w=520000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=5.408e+11p ps=6.24e+06u
M1003 a_734_333# a_533_47# Z VPB phighvt w=820000u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=8.856e+11p ps=8.72e+06u
M1004 Z S[2] a_937_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_1562_333# a_1361_47# Z VPB phighvt w=820000u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1006 a_746_47# S[1] Z VNB nshort w=520000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1007 a_117_297# D[0] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1008 VPWR D[3] a_1562_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Z a_184_265# a_117_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_533_47# S[1] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1011 a_945_297# D[2] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.297e+11p pd=2.69e+06u as=0p ps=0u
M1012 Z a_1012_265# a_945_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR S[0] a_184_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1014 VPWR S[2] a_1012_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1015 a_1361_47# S[3] VGND VNB nshort w=520000u l=150000u
+  ad=1.482e+11p pd=1.61e+06u as=0p ps=0u
M1016 a_533_47# S[1] VGND VNB nshort w=520000u l=150000u
+  ad=1.482e+11p pd=1.61e+06u as=0p ps=0u
M1017 VGND S[0] a_184_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.61e+06u
M1018 VGND D[1] a_746_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR D[1] a_734_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND D[3] a_1574_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_109_47# D[0] VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.95e+06u as=0p ps=0u
M1022 VGND S[2] a_1012_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.61e+06u
M1023 Z S[0] a_109_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o221a_1 A2 X B1 C1 A1 B2 VPB VNB VGND VPWR
M1000 a_124_47# B2 a_230_47# VNB nshort w=650000u l=150000u
+  ad=4.16e+11p pd=3.88e+06u as=3.9975e+11p ps=3.83e+06u
M1001 VPWR A1 a_515_297# VPB phighvt w=1e+06u l=180000u
+  ad=7e+11p pd=5.4e+06u as=2.3e+11p ps=2.46e+06u
M1002 VGND A1 a_230_47# VNB nshort w=650000u l=150000u
+  ad=3.77e+11p pd=3.76e+06u as=0p ps=0u
M1003 a_228_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.3e+11p pd=2.46e+06u as=0p ps=0u
M1004 a_515_297# A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.14e+12p ps=6.28e+06u
M1005 a_27_297# B2 a_228_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_27_297# VGND VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=0p ps=0u
M1007 a_230_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_230_47# B1 a_124_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_27_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=0p ps=0u
M1010 a_124_47# C1 a_27_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1011 VPWR C1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__dlxtn_1 VGND VPWR Q GATE_N D VPB VNB
M1000 a_211_363# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=6.009e+11p ps=6.32e+06u
M1001 VPWR GATE_N a_27_47# VPB phighvt w=640000u l=180000u
+  ad=7.846e+11p pd=7.7e+06u as=1.728e+11p ps=1.82e+06u
M1002 VPWR a_607_47# a_760_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1003 Q a_760_21# VGND VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=0p ps=0u
M1004 a_716_413# a_27_47# a_607_47# VPB phighvt w=420000u l=180000u
+  ad=9.66e+10p pd=1.3e+06u as=1.512e+11p ps=1.56e+06u
M1005 VPWR a_760_21# a_716_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_607_47# a_760_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1007 a_503_369# a_319_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=2.021e+11p pd=1.97e+06u as=0p ps=0u
M1008 VGND D a_319_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1009 a_499_47# a_319_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.554e+11p pd=1.62e+06u as=0p ps=0u
M1010 a_695_47# a_211_363# a_607_47# VNB nshort w=360000u l=150000u
+  ad=1.32e+11p pd=1.49e+06u as=1.044e+11p ps=1.3e+06u
M1011 VPWR D a_319_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1012 VGND GATE_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1013 Q a_760_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.4e+11p pd=2.68e+06u as=0p ps=0u
M1014 a_607_47# a_27_47# a_499_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_211_363# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1016 VGND a_760_21# a_695_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_607_47# a_211_363# a_503_369# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and4_2 X C A B D VNB VPB VGND VPWR
M1000 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=5.1575e+11p pd=4.24e+06u as=2.795e+11p ps=2.16e+06u
M1001 VGND D a_301_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
M1002 a_27_47# A VPWR VPB phighvt w=420000u l=180000u
+  ad=2.478e+11p pd=2.86e+06u as=9.943e+11p ps=8.44e+06u
M1003 a_27_47# C VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.5e+11p pd=2.7e+06u as=0p ps=0u
M1005 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_203_47# B a_119_47# VNB nshort w=420000u l=150000u
+  ad=1.428e+11p pd=1.52e+06u as=1.134e+11p ps=1.38e+06u
M1007 a_119_47# A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1008 VPWR B a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_301_47# C a_203_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR D a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o21bai_1 A1 Y B1_N A2 VPB VNB VPWR VGND
M1000 VPWR A1 a_425_297# VPB phighvt w=1e+06u l=180000u
+  ad=6.607e+11p pd=5.42e+06u as=2.8e+11p ps=2.56e+06u
M1001 a_425_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.2e+11p ps=2.64e+06u
M1002 a_105_352# B1_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=3.615e+11p ps=3.5e+06u
M1003 VGND A2 a_327_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.965e+11p ps=3.82e+06u
M1004 a_327_47# a_105_352# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1005 a_327_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR B1_N a_105_352# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1007 Y a_105_352# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a22o_1 A1 A2 X B2 B1 VPWR VGND VPB VNB
M1000 a_27_297# B1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=6.3e+11p ps=5.26e+06u
M1001 VGND A2 a_411_47# VNB nshort w=650000u l=150000u
+  ad=4.355e+11p pd=3.94e+06u as=2.405e+11p ps=2.04e+06u
M1002 a_27_297# B1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=4.03e+11p pd=3.84e+06u as=1.755e+11p ps=1.84e+06u
M1003 a_117_297# B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_411_47# A1 a_27_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=6e+11p pd=5.2e+06u as=0p ps=0u
M1006 X a_27_297# VGND VNB nshort w=650000u l=150000u
+  ad=2.6e+11p pd=2.1e+06u as=0p ps=0u
M1007 X a_27_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=4.1e+11p pd=2.82e+06u as=0p ps=0u
M1008 a_117_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_119_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sdfbbp_1 SCD SCE RESET_B VGND CLK Q VPWR D Q_N SET_B VPB
+ VNB
M1000 a_2216_47# SET_B VGND VNB nshort w=420000u l=150000u
+  ad=3.931e+11p pd=3.84e+06u as=1.5247e+12p ps=1.429e+07u
M1001 a_211_363# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1002 a_2058_21# SET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=2.583e+11p pd=2.38e+06u as=2.152e+12p ps=1.881e+07u
M1003 VGND SCE a_453_315# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.365e+11p ps=1.49e+06u
M1004 a_810_413# SCE VPWR VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
M1005 Q_N a_2058_21# VGND VNB nshort w=650000u l=150000u
+  ad=2.3075e+11p pd=2.01e+06u as=0p ps=0u
M1006 a_1105_413# a_27_47# a_1003_47# VPB phighvt w=420000u l=180000u
+  ad=1.974e+11p pd=1.78e+06u as=1.218e+11p ps=1.42e+06u
M1007 a_2216_47# a_1525_21# a_2058_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=2.016e+11p ps=1.91e+06u
M1008 VPWR CLK a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1009 a_1353_47# SET_B VGND VNB nshort w=420000u l=150000u
+  ad=4.387e+11p pd=4.01e+06u as=0p ps=0u
M1010 a_1864_47# a_211_363# a_1769_47# VNB nshort w=360000u l=150000u
+  ad=1.764e+11p pd=1.7e+06u as=1.87e+11p ps=1.93e+06u
M1011 VPWR SCE a_453_315# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.449e+11p ps=1.53e+06u
M1012 a_1197_21# SET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=3.066e+11p pd=2.5e+06u as=0p ps=0u
M1013 a_1197_21# a_1003_47# a_1353_47# VNB nshort w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1014 VGND a_2058_21# a_1992_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.341e+11p ps=1.5e+06u
M1015 VPWR a_1197_21# a_1105_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Q a_2845_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1017 VPWR RESET_B a_1525_21# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1018 a_409_363# SCD VPWR VPB phighvt w=640000u l=180000u
+  ad=1.472e+11p pd=1.74e+06u as=0p ps=0u
M1019 a_1121_47# a_211_363# a_1003_47# VNB nshort w=360000u l=150000u
+  ad=1.521e+11p pd=1.6e+06u as=1.584e+11p ps=1.6e+06u
M1020 a_1003_47# a_211_363# a_483_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=3.219e+11p ps=3.37e+06u
M1021 a_1353_47# a_1525_21# a_1197_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_483_47# a_453_315# a_409_363# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_411_47# SCD VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1024 a_483_47# SCE a_411_47# VNB nshort w=420000u l=150000u
+  ad=2.805e+11p pd=3.04e+06u as=0p ps=0u
M1025 VGND a_1197_21# a_1121_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_1525_21# a_1469_329# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=2.436e+11p ps=2.26e+06u
M1027 a_1003_47# a_27_47# a_483_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND RESET_B a_1525_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1029 VPWR a_2058_21# a_1968_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.932e+11p ps=1.76e+06u
M1030 VPWR a_2058_21# a_2845_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1031 a_1469_329# a_1003_47# a_1197_21# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1968_413# a_211_363# a_1864_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1033 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1034 a_2320_329# a_1864_47# a_2058_21# VPB phighvt w=840000u l=180000u
+  ad=1.932e+11p pd=2.14e+06u as=0p ps=0u
M1035 a_483_47# D a_824_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1036 VPWR a_1525_21# a_2320_329# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1769_47# a_1197_21# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_211_363# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1039 Q_N a_2058_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.65e+11p pd=2.73e+06u as=0p ps=0u
M1040 a_2058_21# a_1864_47# a_2216_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1710_329# a_1197_21# VPWR VPB phighvt w=840000u l=180000u
+  ad=4.032e+11p pd=2.96e+06u as=0p ps=0u
M1042 a_1864_47# a_27_47# a_1710_329# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VGND a_2058_21# a_2845_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1044 a_483_47# D a_810_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_824_47# a_453_315# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_1992_47# a_27_47# a_1864_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 Q a_2845_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or2_1 A X B VPB VNB VGND VPWR
M1000 VPWR A a_128_297# VPB phighvt w=420000u l=180000u
+  ad=3.057e+11p pd=2.71e+06u as=9.66e+10p ps=1.3e+06u
M1001 a_128_297# B a_38_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1002 a_38_297# B VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=3.307e+11p ps=3.43e+06u
M1003 X a_38_297# VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=0p ps=0u
M1004 VGND A a_38_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_38_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.5e+11p pd=2.7e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a21oi_1 A1 B1 Y A2 VPWR VGND VPB VNB
M1000 a_121_297# B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=5.75e+11p pd=5.15e+06u as=2.75e+11p ps=2.55e+06u
M1001 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=4.095e+11p ps=3.86e+06u
M1002 a_219_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u
M1003 VPWR A1 a_121_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.15e+11p pd=2.63e+06u as=0p ps=0u
M1004 a_121_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A2 a_219_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand4_2 B A Y D C VNB VPB VGND VPWR
M1000 VPWR D Y VPB phighvt w=1e+06u l=180000u
+  ad=2.18e+12p pd=1.436e+07u as=1.16e+12p ps=1.032e+07u
M1001 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_27_47# D VGND VNB nshort w=650000u l=150000u
+  ad=5.59e+11p pd=5.62e+06u as=2.08e+11p ps=1.94e+06u
M1003 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_511_47# B a_297_47# VNB nshort w=650000u l=150000u
+  ad=6.89e+11p pd=6.02e+06u as=4.485e+11p ps=3.98e+06u
M1005 a_297_47# C a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_511_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1008 Y A a_511_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_297_47# B a_511_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND D a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_47# C a_297_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__decap_6 VPWR VGND VPB VNB
M1000 VPWR VGND VPWR VPB phighvt w=870000u l=1.97e+06u
+  ad=4.524e+11p pd=4.52e+06u as=0p ps=0u
M1001 VGND VPWR VGND VNB nshort w=550000u l=1.97e+06u
+  ad=2.86e+11p pd=3.24e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o211a_1 C1 B1 A2 A1 X VNB VPB VGND VPWR
M1000 a_225_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=4.875e+11p pd=4.1e+06u as=4.4525e+11p ps=3.97e+06u
M1001 a_79_21# C1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=7.7e+11p pd=5.54e+06u as=1.07e+12p ps=8.14e+06u
M1002 VPWR B1 a_79_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_540_47# B1 a_225_47# VNB nshort w=650000u l=150000u
+  ad=3.64e+11p pd=2.42e+06u as=0p ps=0u
M1004 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1005 a_79_21# A2 a_315_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.45e+11p ps=2.69e+06u
M1006 a_79_21# C1 a_540_47# VNB nshort w=650000u l=150000u
+  ad=2.275e+11p pd=2e+06u as=0p ps=0u
M1007 a_315_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1009 VGND A1 a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and3b_2 VGND VPWR B X A_N C VNB VPB
M1000 a_117_311# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=6.936e+11p ps=5.94e+06u
M1001 a_317_53# a_117_311# a_225_311# VNB nshort w=420000u l=150000u
+  ad=1.344e+11p pd=1.48e+06u as=1.218e+11p ps=1.42e+06u
M1002 a_117_311# A_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=9.409e+11p ps=8.31e+06u
M1003 a_225_311# B VPWR VPB phighvt w=420000u l=180000u
+  ad=2.7055e+11p pd=3.05e+06u as=0p ps=0u
M1004 VPWR C a_225_311# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_225_311# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1006 X a_225_311# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_117_311# a_225_311# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_225_311# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1009 a_411_53# B a_317_53# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1010 VGND C a_411_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_225_311# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__bufbuf_16 A X VNB VPB VGND VPWR
M1000 X a_589_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.32e+12p pd=2.064e+07u as=4.02e+12p ps=3.604e+07u
M1001 VGND a_589_47# X VNB nshort w=650000u l=150000u
+  ad=2.8015e+12p pd=2.682e+07u as=1.6965e+12p ps=1.562e+07u
M1002 X a_589_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_589_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_589_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_225_47# a_589_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.7e+11p ps=7.74e+06u
M1006 VGND a_589_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_589_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_225_47# a_589_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_589_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_589_47# a_225_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_589_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_589_47# a_225_47# VGND VNB nshort w=650000u l=150000u
+  ad=6.565e+11p pd=5.92e+06u as=0p ps=0u
M1013 X a_589_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_225_47# a_589_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_589_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_589_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_589_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_589_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_589_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_117_297# a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.095e+11p ps=3.86e+06u
M1021 X a_589_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_117_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1023 VGND a_225_47# a_589_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_589_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_589_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 X a_589_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR a_117_297# a_225_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.6e+11p ps=5.12e+06u
M1028 VGND a_589_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_589_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 X a_589_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_589_47# a_225_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 X a_589_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_589_47# a_225_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 X a_589_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_225_47# a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 X a_589_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_117_297# A VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1038 a_225_47# a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR a_225_47# a_589_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VPWR a_589_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPWR a_589_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPWR a_117_297# a_225_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VGND a_589_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VPWR a_589_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_589_47# a_225_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 VPWR a_589_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VGND a_225_47# a_589_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 X a_589_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_589_47# a_225_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1050 VGND a_117_297# a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1051 VGND a_589_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__xnor2_2 VGND VPWR Y A B VPB VNB
M1000 a_514_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.5e+11p pd=7.7e+06u as=1.43e+12p ps=1.286e+07u
M1001 Y a_27_297# a_600_47# VNB nshort w=650000u l=150000u
+  ad=3.38e+11p pd=3.64e+06u as=7.4425e+11p ps=6.19e+06u
M1002 a_27_47# A VGND VNB nshort w=650000u l=150000u
+  ad=5.6875e+11p pd=5.65e+06u as=7.345e+11p ps=7.46e+06u
M1003 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND B a_600_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.65e+11p ps=7.73e+06u
M1006 VPWR A a_514_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_47# B a_27_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.405e+11p ps=2.04e+06u
M1008 VPWR a_27_297# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=6.15e+11p ps=5.23e+06u
M1009 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y a_27_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A a_600_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_600_47# a_27_297# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_600_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y B a_514_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_297# B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_600_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_514_297# B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__clkbuf_8 X A VPB VNB VGND VPWR
M1000 VGND a_118_297# X VNB nshort w=420000u l=150000u
+  ad=7.791e+11p pd=8.75e+06u as=5.754e+11p ps=6.1e+06u
M1001 a_118_297# A VGND VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=0p ps=0u
M1002 VGND A a_118_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR a_118_297# X VPB phighvt w=1e+06u l=180000u
+  ad=1.75e+12p pd=1.55e+07u as=1.2e+12p ps=1.04e+07u
M1004 a_118_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1005 X a_118_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_118_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_118_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_118_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_118_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_118_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_118_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_118_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A a_118_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_118_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_118_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_118_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_118_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_118_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_118_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__clkinv_8 Y A VNB VPB VGND VPWR
M1000 VGND A Y VNB nshort w=420000u l=150000u
+  ad=7.014e+11p pd=7.54e+06u as=5.964e+11p ps=6.2e+06u
M1001 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=2.095e+12p pd=1.819e+07u as=1.79e+12p ps=1.558e+07u
M1002 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sdfxtp_4 VGND VPWR SCD D SCE CLK Q VNB VPB
M1000 VPWR a_1189_183# a_1121_413# VPB phighvt w=420000u l=180000u
+  ad=1.98115e+12p pd=1.754e+07u as=1.47e+11p ps=1.54e+06u
M1001 VPWR CLK a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1002 a_608_369# D a_517_47# VNB nshort w=420000u l=150000u
+  ad=2.604e+11p pd=2.88e+06u as=1.428e+11p ps=1.52e+06u
M1003 a_1474_413# a_27_47# a_1189_183# VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=2.307e+11p ps=2.19e+06u
M1004 VPWR a_1667_315# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1005 VGND a_1667_315# a_1625_47# VNB nshort w=420000u l=150000u
+  ad=1.48085e+12p pd=1.433e+07u as=1.32e+11p ps=1.49e+06u
M1006 VGND a_1667_315# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.485e+11p ps=3.98e+06u
M1007 VGND a_1189_183# a_1127_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.584e+11p ps=1.62e+06u
M1008 a_504_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=2.176e+11p pd=1.96e+06u as=0p ps=0u
M1009 a_203_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1010 VPWR a_1667_315# a_1568_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=2.121e+11p ps=1.85e+06u
M1011 VGND a_1667_315# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR SCE a_319_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1013 a_1121_413# a_27_47# a_1011_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.407e+11p ps=1.51e+06u
M1014 a_1474_413# a_203_47# a_1189_183# VNB nshort w=360000u l=150000u
+  ad=1.854e+11p pd=1.75e+06u as=1.978e+11p ps=1.99e+06u
M1015 Q a_1667_315# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND SCE a_319_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1017 Q a_1667_315# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_1667_315# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_1474_413# a_1667_315# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1020 a_517_47# a_319_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1127_47# a_203_47# a_1011_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.548e+11p ps=1.58e+06u
M1022 a_1189_183# a_1011_47# VPWR VPB phighvt w=750000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q a_1667_315# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1011_47# a_203_47# a_608_369# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=3.2e+11p ps=3.34e+06u
M1025 Q a_1667_315# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_203_47# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1027 a_1625_47# a_27_47# a_1474_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR SCD a_702_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=2.144e+11p ps=1.95e+06u
M1029 VGND SCD a_721_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=9.66e+10p ps=1.3e+06u
M1030 VPWR a_1474_413# a_1667_315# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1031 a_702_369# a_319_47# a_608_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1189_183# a_1011_47# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1568_413# a_203_47# a_1474_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1011_47# a_27_47# a_608_369# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1036 a_721_47# SCE a_608_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_608_369# D a_504_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or4b_2 C A X B D_N VPWR VGND VPB VNB
M1000 a_425_297# A VPWR VPB phighvt w=420000u l=180000u
+  ad=1.47e+11p pd=1.54e+06u as=7.227e+11p ps=6.17e+06u
M1001 X a_186_21# VGND VNB nshort w=650000u l=150000u
+  ad=2.08e+11p pd=1.94e+06u as=6.771e+11p ps=6.88e+06u
M1002 VGND a_27_47# a_186_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.15e+11p ps=3.18e+06u
M1003 a_186_21# a_27_47# a_615_297# VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=1.428e+11p ps=1.52e+06u
M1004 VPWR D_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1005 VPWR a_186_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1006 a_615_297# C a_531_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 VGND B a_186_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_531_297# B a_425_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_186_21# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND D_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1011 a_186_21# C VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_186_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_186_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a2bb2o_2 VNB VPB VGND VPWR B1 A1_N A2_N X B2
M1000 X a_82_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=8.49e+11p ps=7.32e+06u
M1001 a_696_47# B2 a_82_21# VNB nshort w=420000u l=150000u
+  ad=1.344e+11p pd=1.48e+06u as=1.134e+11p ps=1.38e+06u
M1002 a_343_47# A2_N a_341_297# VPB phighvt w=640000u l=180000u
+  ad=1.76e+11p pd=1.83e+06u as=1.472e+11p ps=1.74e+06u
M1003 VGND a_82_21# X VNB nshort w=650000u l=150000u
+  ad=9.0065e+11p pd=7.95e+06u as=2.08e+11p ps=1.94e+06u
M1004 a_622_369# B1 VPWR VPB phighvt w=640000u l=180000u
+  ad=3.808e+11p pd=3.75e+06u as=0p ps=0u
M1005 VGND A2_N a_343_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1006 a_343_47# A1_N VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_622_369# a_343_47# a_82_21# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1008 a_341_297# A1_N VPWR VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR B2 a_622_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_82_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_82_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND B1 a_696_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_82_21# a_343_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__xor3_2 X C B A VNB VPB VGND VPWR
M1000 VPWR A a_1050_365# VPB phighvt w=1e+06u l=180000u
+  ad=1.2694e+12p pd=1.06e+07u as=7.234e+11p ps=5.3e+06u
M1001 X a_81_21# VGND VNB nshort w=650000u l=150000u
+  ad=2.275e+11p pd=2e+06u as=8.9605e+11p ps=8e+06u
M1002 a_81_21# C a_483_49# VNB nshort w=640000u l=150000u
+  ad=2.848e+11p pd=2.17e+06u as=5.963e+11p ps=4.53e+06u
M1003 a_483_49# a_335_93# a_81_21# VPB phighvt w=840000u l=180000u
+  ad=7.558e+11p pd=5.2e+06u as=3.36e+11p ps=2.48e+06u
M1004 a_934_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.126e+11p pd=2.64e+06u as=0p ps=0u
M1005 a_465_325# B a_1335_297# VNB nshort w=640000u l=150000u
+  ad=6.6045e+11p pd=4.67e+06u as=5.517e+11p ps=4.37e+06u
M1006 VGND A a_1050_365# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=4.468e+11p ps=3.98e+06u
M1007 X a_81_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=0p ps=0u
M1008 a_335_93# C VGND VNB nshort w=420000u l=150000u
+  ad=1.974e+11p pd=1.78e+06u as=0p ps=0u
M1009 a_483_49# B a_1050_365# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1050_365# a_934_297# a_483_49# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1335_297# a_934_297# a_483_49# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_335_93# C VPWR VPB phighvt w=640000u l=180000u
+  ad=1.856e+11p pd=1.86e+06u as=0p ps=0u
M1013 a_81_21# C a_465_325# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=7.824e+11p ps=5.28e+06u
M1014 a_483_49# B a_1335_297# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=7.798e+11p ps=5.64e+06u
M1015 a_1050_365# a_934_297# a_465_325# VNB nshort w=600000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_81_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1335_297# a_934_297# a_465_325# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_934_297# B VGND VNB nshort w=650000u l=150000u
+  ad=1.978e+11p pd=1.92e+06u as=0p ps=0u
M1019 a_465_325# a_335_93# a_81_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1335_297# a_1050_365# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_465_325# B a_1050_365# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_81_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1335_297# a_1050_365# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__dlrtp_2 RESET_B D GATE Q VGND VPWR VPB VNB
M1000 VGND a_750_21# a_708_47# VNB nshort w=420000u l=150000u
+  ad=8.0475e+11p pd=8.18e+06u as=8.82e+10p ps=1.26e+06u
M1001 VPWR GATE a_27_363# VPB phighvt w=640000u l=180000u
+  ad=1.411e+12p pd=1.231e+07u as=1.728e+11p ps=1.82e+06u
M1002 VPWR a_750_21# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1003 a_203_47# a_27_363# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1004 VPWR a_750_21# a_702_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1005 VGND a_750_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1006 a_503_369# a_319_369# VPWR VPB phighvt w=640000u l=180000u
+  ad=2.021e+11p pd=1.97e+06u as=0p ps=0u
M1007 a_708_47# a_27_363# a_604_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.58e+06u
M1008 Q a_750_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Q a_750_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND D a_319_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1011 VPWR D a_319_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1012 VGND RESET_B a_981_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.6575e+11p ps=1.81e+06u
M1013 a_604_47# a_203_47# a_500_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.482e+11p ps=1.58e+06u
M1014 VPWR RESET_B a_750_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1015 a_981_47# a_604_47# a_750_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1016 VGND GATE a_27_363# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1017 a_702_413# a_203_47# a_604_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1018 a_203_47# a_27_363# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1019 a_604_47# a_27_363# a_503_369# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_500_47# a_319_369# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_750_21# a_604_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__buf_2 VPWR VGND X A VPB VNB
M1000 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=4.4425e+11p pd=4.02e+06u as=1.302e+11p ps=1.46e+06u
M1001 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=3.0875e+11p pd=2.25e+06u as=0p ps=0u
M1002 VPWR A a_27_47# VPB phighvt w=640000u l=180000u
+  ad=7.094e+11p pd=5.48e+06u as=1.728e+11p ps=1.82e+06u
M1003 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.95e+11p pd=2.79e+06u as=0p ps=0u
M1004 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__inv_12 A Y VNB VPB VGND VPWR
M1000 Y A VGND VNB nshort w=650000u l=150000u
+  ad=1.2805e+12p pd=1.174e+07u as=1.3845e+12p ps=1.336e+07u
M1001 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.74e+12p pd=1.548e+07u as=2e+12p ps=1.8e+07u
M1003 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__inv_2 A Y VPB VNB VPWR VGND
M1000 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=5.4e+11p ps=5.08e+06u
M1001 VGND A Y VNB nshort w=650000u l=150000u
+  ad=3.705e+11p pd=3.74e+06u as=2.08e+11p ps=1.94e+06u
M1002 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__dlygate4sd3_1 A X VPWR VGND VPB VNB
M1000 VPWR a_273_47# a_379_93# VPB phighvt w=420000u l=500000u
+  ad=4.491e+11p pd=4.15e+06u as=1.092e+11p ps=1.36e+06u
M1001 X a_379_93# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1002 VPWR A a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1003 a_273_47# a_27_47# VGND VNB nshort w=420000u l=500000u
+  ad=1.092e+11p pd=1.36e+06u as=3.636e+11p ps=3.51e+06u
M1004 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1005 X a_379_93# VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1006 VGND a_273_47# a_379_93# VNB nshort w=420000u l=500000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1007 a_273_47# a_27_47# VPWR VPB phighvt w=420000u l=500000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__muxb8to1_4 VGND Z VPWR VNB VPB S[6] D[3] D[0] D[4] D[5]
+ D[2] D[1] D[6] S[2] S[3] S[7] S[0] S[1] S[4] S[5] D[7]
M1000 a_1313_591# D[3] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.2606e+12p pd=1.174e+07u as=9.4224e+12p ps=8.664e+07u
M1001 VPWR S[0] a_142_325# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1002 a_3797_297# a_4239_265# Z VPB phighvt w=820000u l=180000u
+  ad=1.2606e+12p pd=1.174e+07u as=3.8048e+12p ps=3.552e+07u
M1003 a_405_66# S[0] Z VNB nshort w=520000u l=150000u
+  ad=7.618e+11p pd=8.38e+06u as=2.2464e+12p ps=2.528e+07u
M1004 Z a_2626_325# a_2839_311# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=1.2606e+12p ps=1.174e+07u
M1005 a_3799_47# D[6] VGND VNB nshort w=650000u l=150000u
+  ad=7.618e+11p pd=8.38e+06u as=6.1412e+12p ps=6.128e+07u
M1006 a_2889_66# S[4] Z VNB nshort w=520000u l=150000u
+  ad=7.618e+11p pd=8.38e+06u as=0p ps=0u
M1007 a_1755_793# S[3] VPWR VPB phighvt w=820000u l=180000u
+  ad=2.378e+11p pd=2.22e+06u as=0p ps=0u
M1008 Z S[7] a_3799_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=7.618e+11p ps=8.38e+06u
M1009 Z S[5] a_2889_918# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=7.618e+11p ps=8.38e+06u
M1010 a_355_311# a_142_325# Z VPB phighvt w=820000u l=180000u
+  ad=1.2606e+12p pd=1.174e+07u as=0p ps=0u
M1011 a_3797_591# a_4239_793# Z VPB phighvt w=820000u l=180000u
+  ad=1.2606e+12p pd=1.174e+07u as=0p ps=0u
M1012 a_355_311# D[0] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND D[2] a_1315_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.618e+11p ps=8.38e+06u
M1014 VGND D[7] a_3799_911# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1315_911# D[3] VGND VNB nshort w=650000u l=150000u
+  ad=7.618e+11p pd=8.38e+06u as=0p ps=0u
M1016 Z S[3] a_1315_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_355_613# D[1] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.2606e+12p pd=1.174e+07u as=0p ps=0u
M1018 VPWR S[5] a_2626_599# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1019 Z a_142_325# a_355_311# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1315_911# S[3] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_2839_613# a_2626_599# Z VPB phighvt w=820000u l=180000u
+  ad=1.2606e+12p pd=1.174e+07u as=0p ps=0u
M1022 Z S[4] a_2889_66# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Z a_4239_265# a_3797_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Z S[2] a_1315_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND D[7] a_3799_911# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_3799_911# D[7] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND D[4] a_2889_66# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1315_47# S[2] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_405_918# S[1] Z VNB nshort w=520000u l=150000u
+  ad=7.618e+11p pd=8.38e+06u as=0p ps=0u
M1030 a_405_918# D[1] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Z a_1755_793# a_1313_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_4239_265# S[6] VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1033 VGND D[5] a_2889_918# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_2889_66# D[4] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_2889_66# S[4] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1313_591# a_1755_793# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1315_47# D[2] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 Z S[5] a_2889_918# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_2626_599# S[5] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_142_325# S[0] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 Z a_2626_599# a_2839_613# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPWR D[4] a_2839_311# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VGND S[0] a_142_325# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1044 Z S[2] a_1315_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_2889_66# D[4] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 VPWR D[5] a_2839_613# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VGND D[3] a_1315_911# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_1315_911# S[3] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 VPWR D[0] a_355_311# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1050 Z a_1755_265# a_1313_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=1.2606e+12p ps=1.174e+07u
M1051 Z a_142_325# a_355_311# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1052 VPWR S[1] a_142_599# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1053 Z a_4239_793# a_3797_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1054 a_355_613# a_142_599# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1055 VPWR D[1] a_355_613# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1056 a_2839_613# a_2626_599# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1057 a_1315_47# S[2] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1058 Z S[1] a_405_918# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1059 VGND D[1] a_405_918# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1060 VGND S[3] a_1755_793# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1061 VGND S[6] a_4239_265# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1062 a_2839_311# D[4] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1063 a_3799_911# S[7] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1064 VPWR S[6] a_4239_265# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1065 a_405_66# D[0] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1066 Z S[4] a_2889_66# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1067 a_142_325# S[0] VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1068 a_405_918# D[1] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1069 VGND D[2] a_1315_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1070 a_2839_613# D[5] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1071 VPWR D[2] a_1313_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1072 VPWR S[2] a_1755_265# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1073 a_1313_297# a_1755_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1074 VGND S[5] a_2626_599# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1075 a_3797_591# a_4239_793# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1076 VPWR D[3] a_1313_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1077 a_2889_918# D[5] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1078 Z a_2626_599# a_2839_613# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1079 VGND D[4] a_2889_66# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1080 a_355_613# a_142_599# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1081 VGND D[6] a_3799_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1082 a_3797_297# D[6] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1083 a_405_918# S[1] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1084 a_142_599# S[1] VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1085 a_4239_265# S[6] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1086 a_355_311# D[0] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1087 a_3797_591# D[7] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1088 a_142_599# S[1] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1089 a_3799_47# S[6] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1090 a_1313_297# D[2] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1091 a_3799_911# S[7] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1092 Z a_142_599# a_355_613# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1093 a_355_613# D[1] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1094 VGND S[2] a_1755_265# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1095 a_1313_591# D[3] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1096 Z a_4239_793# a_3797_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1097 VGND D[0] a_405_66# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1098 a_3799_911# D[7] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1099 a_3797_297# a_4239_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1100 a_405_66# S[0] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1101 Z S[6] a_3799_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1102 Z S[1] a_405_918# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1103 a_1755_265# S[2] VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1104 a_1315_911# D[3] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1105 VPWR D[4] a_2839_311# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1106 VGND D[5] a_2889_918# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1107 a_2889_918# D[5] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1108 VPWR D[6] a_3797_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1109 Z S[0] a_405_66# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1110 a_2839_311# a_2626_325# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1111 a_3799_47# D[6] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1112 a_2889_918# S[5] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1113 VPWR D[5] a_2839_613# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1114 a_4239_793# S[7] VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1115 a_1755_265# S[2] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1116 Z a_1755_265# a_1313_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1117 VPWR D[7] a_3797_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1118 VPWR D[2] a_1313_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1119 VPWR S[7] a_4239_793# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1120 VPWR D[3] a_1313_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1121 VGND S[4] a_2626_325# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1122 a_3799_47# S[6] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1123 Z a_142_599# a_355_613# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1124 Z a_1755_793# a_1313_591# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1125 VPWR S[3] a_1755_793# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1126 a_1313_297# a_1755_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1127 a_2839_311# D[4] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1128 VPWR S[4] a_2626_325# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.378e+11p ps=2.22e+06u
M1129 a_2626_325# S[4] VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1130 a_3797_297# D[6] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1131 Z a_2626_325# a_2839_311# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1132 Z S[6] a_3799_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1133 Z S[0] a_405_66# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1134 a_2839_613# D[5] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1135 Z S[3] a_1315_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1136 VGND D[3] a_1315_911# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1137 VPWR D[0] a_355_311# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1138 VGND S[1] a_142_599# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1139 a_3797_591# D[7] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1140 a_1755_793# S[3] VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1141 VPWR D[1] a_355_613# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1142 a_2889_918# S[5] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1143 Z a_4239_265# a_3797_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1144 Z S[7] a_3799_911# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1145 VPWR D[6] a_3797_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1146 a_2839_311# a_2626_325# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1147 a_355_311# a_142_325# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1148 a_4239_793# S[7] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1149 VGND S[7] a_4239_793# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1150 a_1315_47# D[2] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1151 VGND D[0] a_405_66# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1152 a_1313_591# a_1755_793# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1153 VPWR D[7] a_3797_591# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1154 a_2626_599# S[5] VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1155 a_2626_325# S[4] VPWR VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1156 a_405_66# D[0] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1157 VGND D[1] a_405_918# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1158 a_1313_297# D[2] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1159 VGND D[6] a_3799_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__mux2_8 S A1 VPWR VGND VPB VNB A0 X
M1000 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=2.16e+12p pd=1.832e+07u as=1.16e+12p ps=1.032e+07u
M1001 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_870_297# A0 a_79_21# VPB phighvt w=1e+06u l=180000u
+  ad=1.385e+12p pd=6.77e+06u as=5.8e+11p ps=5.16e+06u
M1003 a_79_21# A1 a_872_47# VNB nshort w=640000u l=150000u
+  ad=4.096e+11p pd=3.84e+06u as=9.568e+11p ps=5.55e+06u
M1004 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_872_47# A1 a_79_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=8.645e+11p pd=7.86e+06u as=1.5084e+12p ps=1.374e+07u
M1007 VGND S a_872_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_1369_199# a_1422_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.0464e+12p ps=5.83e+06u
M1012 a_79_21# A0 a_870_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_1369_199# a_1420_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.675e+12p ps=7.35e+06u
M1014 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1420_297# a_1369_199# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1420_297# A1 a_79_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_79_21# A0 a_1422_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1369_199# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1020 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_870_297# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_872_47# S VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_79_21# A1 a_1420_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1422_47# a_1369_199# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1422_47# A0 a_79_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1369_199# S VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=0p ps=0u
M1033 VPWR S a_870_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o2bb2a_4 A2_N A1_N X B2 B1 VNB VPB VGND VPWR
M1000 a_787_47# A1_N VGND VNB nshort w=650000u l=150000u
+  ad=3.835e+11p pd=3.78e+06u as=1.1375e+12p ps=1.13e+07u
M1001 a_211_297# B2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=5.8e+11p ps=5.16e+06u
M1002 X a_211_297# VGND VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=0p ps=0u
M1003 X a_211_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=2.51e+12p ps=1.902e+07u
M1004 VPWR A1_N a_455_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1005 VPWR a_455_21# a_211_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=8.19e+11p pd=7.72e+06u as=0p ps=0u
M1007 VGND a_211_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_211_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_117_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A1_N a_787_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_211_297# a_455_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_211_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_455_21# A2_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR B1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_211_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_787_47# A2_N a_455_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.405e+11p ps=2.04e+06u
M1017 VGND B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A2_N a_455_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_211_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_27_47# a_455_21# a_211_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1022 a_211_297# a_455_21# a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_117_297# B2 a_211_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_211_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_455_21# A2_N a_787_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_455_21# A1_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor4b_2 D_N Y C A B VNB VPB VGND VPWR
M1000 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.3e+11p pd=7.66e+06u as=4.034e+11p ps=3.96e+06u
M1001 VGND A Y VNB nshort w=650000u l=150000u
+  ad=1.1897e+12p pd=1.252e+07u as=9.295e+11p ps=8.06e+06u
M1002 VGND D_N a_754_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1003 Y a_754_21# a_514_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=8.3e+11p ps=7.66e+06u
M1004 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR D_N a_754_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1006 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_514_297# C a_305_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1008 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_305_297# C a_514_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_297# B a_305_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_754_21# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_305_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y a_754_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_514_297# a_754_21# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a211oi_2 A2 C1 B1 Y A1 VPWR VGND VPB VNB
M1000 VPWR A2 a_320_297# VPB phighvt w=1e+06u l=180000u
+  ad=8.5e+11p pd=7.7e+06u as=9e+11p ps=7.8e+06u
M1001 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=7.085e+11p pd=6.08e+06u as=8.06e+11p ps=7.68e+06u
M1002 a_525_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=5.265e+11p pd=5.52e+06u as=0p ps=0u
M1003 a_320_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y C1 a_37_297# VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=8.5e+11p ps=7.7e+06u
M1005 a_320_297# B1 a_37_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A1 a_525_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_320_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A2 a_525_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_525_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_37_297# C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y C1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_37_297# B1 a_320_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND C1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A1 a_320_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or3_4 A X B C VPB VNB VPWR VGND
M1000 a_211_297# B a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u
M1001 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=3.77e+11p pd=3.76e+06u as=1.20575e+12p ps=8.91e+06u
M1002 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=1.48e+12p pd=8.96e+06u as=5.8e+11p ps=5.16e+06u
M1003 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_117_297# C a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1006 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1007 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND C a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A a_211_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o22ai_4 A1 Y A2 B1 B2 VNB VPB VGND VPWR
M1000 Y A2 a_123_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=1.16e+12p ps=1.032e+07u
M1001 Y B2 a_885_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.16e+12p ps=1.032e+07u
M1002 a_33_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=1.924e+12p pd=1.762e+07u as=7.995e+11p ps=7.66e+06u
M1003 a_885_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.49e+12p ps=1.298e+07u
M1004 Y B1 a_33_47# VNB nshort w=650000u l=150000u
+  ad=7.995e+11p pd=7.66e+06u as=0p ps=0u
M1005 a_33_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_33_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_123_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_885_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_33_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y B2 a_33_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A1 a_123_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A1 a_123_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y B2 a_885_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y B1 a_33_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_123_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A2 a_33_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_33_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_885_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A1 a_33_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_33_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y B2 a_33_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y A2 a_123_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR B1 a_885_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_33_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_123_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND A2 a_33_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_123_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_885_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_33_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR B1 a_885_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND A1 a_33_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__mux2_12 VPWR VGND VPB VNB X S A1 A0
M1000 a_119_47# S VGND VNB nshort w=650000u l=150000u
+  ad=7.02e+11p pd=7.36e+06u as=2.9705e+12p ps=2.604e+07u
M1001 VGND a_973_297# a_1163_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.02e+11p ps=7.36e+06u
M1002 a_27_47# A1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.66e+12p pd=1.532e+07u as=1.16e+12p ps=1.032e+07u
M1003 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=3.69e+12p pd=3.338e+07u as=1.74e+12p ps=1.548e+07u
M1004 a_27_47# A0 a_1163_47# VNB nshort w=650000u l=150000u
+  ad=1.287e+12p pd=1.176e+07u as=0p ps=0u
M1005 a_117_297# a_973_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR S a_597_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.16e+12p ps=1.032e+07u
M1007 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_597_297# A0 a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1163_47# a_973_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_47# A0 a_597_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1163_47# A0 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR S a_973_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1013 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.053e+12p pd=1.104e+07u as=0p ps=0u
M1015 a_597_297# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_47# A1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_597_297# A0 a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND S a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_119_47# S VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_973_297# a_1163_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_117_297# A1 a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_973_297# a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_27_47# A0 a_597_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_973_297# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_27_47# A1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_117_297# a_973_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_973_297# S VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1039 VGND S a_973_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_119_47# A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_27_47# A0 a_1163_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPWR S a_597_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_1163_47# a_973_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_1163_47# A0 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_117_297# A1 a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1049 VPWR a_973_297# a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1050 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1051 a_27_47# A1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1052 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1053 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1054 VGND S a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1055 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1056 a_597_297# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1057 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1058 a_119_47# A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1059 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__inputiso1n_1 A SLEEP_B X VGND VPWR VNB VPB
M1000 VGND SLEEP_B a_27_53# VNB nshort w=420000u l=150000u
+  ad=5.9745e+11p pd=4.64e+06u as=1.302e+11p ps=1.46e+06u
M1001 VPWR A a_319_297# VPB phighvt w=420000u l=180000u
+  ad=4.241e+11p pd=4.1e+06u as=1.218e+11p ps=1.42e+06u
M1002 a_27_53# SLEEP_B VPWR VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
M1003 a_319_297# a_27_53# a_229_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1004 X a_229_297# VGND VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=0p ps=0u
M1005 VGND A a_229_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1006 a_229_297# a_27_53# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_229_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o21a_1 X A1 B1 A2 VPB VNB VGND VPWR
M1000 VPWR a_83_21# X VPB phighvt w=1e+06u l=180000u
+  ad=1.255e+12p pd=6.51e+06u as=2.9e+11p ps=2.58e+06u
M1001 a_394_297# A2 a_83_21# VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=3.6e+11p ps=2.72e+06u
M1002 VGND a_83_21# X VNB nshort w=650000u l=150000u
+  ad=3.835e+11p pd=3.78e+06u as=1.82e+11p ps=1.86e+06u
M1003 a_302_47# B1 a_83_21# VNB nshort w=650000u l=150000u
+  ad=3.445e+11p pd=3.66e+06u as=1.7225e+11p ps=1.83e+06u
M1004 VGND A2 a_302_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_83_21# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_394_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_302_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand2b_4 B A_N Y VNB VPB VGND VPWR
M1000 VGND B a_225_47# VNB nshort w=650000u l=150000u
+  ad=6.175e+11p pd=5.8e+06u as=1.05625e+12p ps=9.75e+06u
M1001 a_225_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=1.825e+12p pd=1.565e+07u as=1.16e+12p ps=1.032e+07u
M1003 VPWR a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_225_47# a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1005 Y a_27_47# a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A_N a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1007 VGND B a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_225_47# a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A_N a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1014 Y a_27_47# a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_225_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__decap_4 VGND VPWR VPB VNB
M1000 VPWR VGND VPWR VPB phighvt w=870000u l=1.05e+06u
+  ad=4.524e+11p pd=4.52e+06u as=0p ps=0u
M1001 VGND VPWR VGND VNB nshort w=550000u l=1.05e+06u
+  ad=2.86e+11p pd=3.24e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o211ai_4 A1 B1 A2 C1 Y VNB VPB VGND VPWR
M1000 a_27_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=1.586e+12p pd=1.398e+07u as=8.32e+11p ps=7.76e+06u
M1001 VPWR C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=2.48e+12p pd=1.896e+07u as=1.77e+12p ps=1.554e+07u
M1002 Y A2 a_118_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.2e+12p ps=1.04e+07u
M1003 VGND A2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_886_47# C1 Y VNB nshort w=650000u l=150000u
+  ad=4.225e+11p pd=3.9e+06u as=4.485e+11p ps=3.98e+06u
M1005 Y C1 a_1088_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1006 Y B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_886_47# B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1088_47# B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_118_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_47# B1 a_886_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_118_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A1 a_118_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_47# B1 a_1464_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.47e+11p ps=2.06e+06u
M1019 Y C1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1464_47# C1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_118_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR A1 a_118_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_27_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_118_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y C1 a_886_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y A2 a_118_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND A2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y C1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor2_1 B Y A VPB VNB VGND VPWR
M1000 VPWR A a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=6.1e+11p pd=3.22e+06u as=2.9e+11p ps=2.58e+06u
M1001 VGND A Y VNB nshort w=650000u l=150000u
+  ad=5.915e+11p pd=4.42e+06u as=1.755e+11p ps=1.84e+06u
M1002 a_117_297# B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1003 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nand4b_1 Y C D A_N B VPB VNB VGND VPWR
M1000 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=1.0157e+12p ps=8.13e+06u
M1001 VGND A_N a_40_93# VNB nshort w=420000u l=150000u
+  ad=2.6875e+11p pd=2.18e+06u as=1.323e+11p ps=1.47e+06u
M1002 VPWR A_N a_40_93# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1003 VPWR a_40_93# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_431_47# B a_334_47# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=2.1775e+11p ps=1.97e+06u
M1005 Y a_40_93# a_431_47# VNB nshort w=650000u l=150000u
+  ad=2.925e+11p pd=2.2e+06u as=0p ps=0u
M1006 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_334_47# C a_251_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u
M1008 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_251_47# D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__clkmux2_4 VGND VPWR S A1 A0 X VPB VNB
M1000 VPWR a_79_199# X VPB phighvt w=1e+06u l=180000u
+  ad=1.3588e+12p pd=1.066e+07u as=5.8e+11p ps=5.16e+06u
M1001 VGND a_925_21# a_754_47# VNB nshort w=420000u l=150000u
+  ad=8.016e+11p pd=7.42e+06u as=3.591e+11p ps=2.55e+06u
M1002 a_925_21# S VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1003 X a_79_199# VGND VNB nshort w=520000u l=150000u
+  ad=2.808e+11p pd=3.16e+06u as=0p ps=0u
M1004 X a_79_199# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_79_199# A1 a_525_47# VNB nshort w=420000u l=150000u
+  ad=2.121e+11p pd=1.85e+06u as=1.428e+11p ps=1.52e+06u
M1006 a_925_21# S VPWR VPB phighvt w=940000u l=180000u
+  ad=2.726e+11p pd=2.46e+06u as=0p ps=0u
M1007 a_875_309# A1 a_79_199# VPB phighvt w=940000u l=180000u
+  ad=2.444e+11p pd=2.4e+06u as=9.447e+11p ps=3.89e+06u
M1008 X a_79_199# VGND VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_754_47# A0 a_79_199# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_79_199# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_79_199# X VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_523_309# S VPWR VPB phighvt w=940000u l=180000u
+  ad=3.713e+11p pd=2.67e+06u as=0p ps=0u
M1013 a_79_199# A0 a_523_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_79_199# X VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_79_199# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_525_47# S VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_925_21# a_875_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o21ai_4 Y B1 A2 A1 VNB VPB VPWR VGND
M1000 a_123_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=1.2e+12p pd=1.04e+07u as=1.2e+12p ps=1.04e+07u
M1001 a_32_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=1.4625e+12p pd=1.36e+07u as=8.515e+11p ps=7.82e+06u
M1002 a_32_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A1 a_123_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.49e+12p pd=1.298e+07u as=0p ps=0u
M1004 a_123_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_32_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2 a_32_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A2 a_123_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A2 a_32_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B1 a_32_47# VNB nshort w=650000u l=150000u
+  ad=4.615e+11p pd=4.02e+06u as=0p ps=0u
M1012 a_32_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A1 a_32_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A2 a_123_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A1 a_32_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y B1 a_32_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_32_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_32_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_123_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_123_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR A1 a_123_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__clkbuf_6 A X VPB VNB VGND VPWR
M1000 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=1.41e+12p pd=1.282e+07u as=8.7e+11p ps=7.74e+06u
M1001 VPWR A a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1002 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A a_117_297# VNB nshort w=420000u l=150000u
+  ad=7.245e+11p pd=7.65e+06u as=1.134e+11p ps=1.38e+06u
M1005 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=3.423e+11p pd=4.15e+06u as=0p ps=0u
M1006 a_117_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_117_297# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sdfxtp_2 VPWR VGND SCE D SCD Q CLK VNB VPB
M1000 VPWR a_1189_183# a_1121_413# VPB phighvt w=420000u l=180000u
+  ad=1.71115e+12p pd=1.5e+07u as=1.47e+11p ps=1.54e+06u
M1001 VPWR CLK a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1002 a_608_369# D a_517_47# VNB nshort w=420000u l=150000u
+  ad=2.604e+11p pd=2.88e+06u as=1.428e+11p ps=1.52e+06u
M1003 a_1474_413# a_27_47# a_1189_183# VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=2.307e+11p ps=2.19e+06u
M1004 VPWR a_1667_315# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1005 VGND a_1667_315# Q VNB nshort w=650000u l=150000u
+  ad=1.30535e+12p pd=1.249e+07u as=2.405e+11p ps=2.04e+06u
M1006 VGND a_1667_315# a_1625_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.32e+11p ps=1.49e+06u
M1007 VGND a_1189_183# a_1127_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.584e+11p ps=1.62e+06u
M1008 a_504_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=2.176e+11p pd=1.96e+06u as=0p ps=0u
M1009 a_203_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1010 VPWR a_1667_315# a_1568_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=2.121e+11p ps=1.85e+06u
M1011 VPWR SCE a_319_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1012 a_1121_413# a_27_47# a_1011_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.407e+11p ps=1.51e+06u
M1013 a_1474_413# a_203_47# a_1189_183# VNB nshort w=360000u l=150000u
+  ad=1.854e+11p pd=1.75e+06u as=1.978e+11p ps=1.99e+06u
M1014 VGND SCE a_319_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1015 Q a_1667_315# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_1474_413# a_1667_315# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1017 a_517_47# a_319_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1127_47# a_203_47# a_1011_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.548e+11p ps=1.58e+06u
M1019 a_1189_183# a_1011_47# VPWR VPB phighvt w=750000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Q a_1667_315# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1011_47# a_203_47# a_608_369# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=3.2e+11p ps=3.34e+06u
M1022 a_203_47# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1023 a_1625_47# a_27_47# a_1474_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR SCD a_702_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=2.144e+11p ps=1.95e+06u
M1025 VGND SCD a_721_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=9.66e+10p ps=1.3e+06u
M1026 VPWR a_1474_413# a_1667_315# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1027 a_702_369# a_319_47# a_608_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1189_183# a_1011_47# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1568_413# a_203_47# a_1474_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1011_47# a_27_47# a_608_369# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1032 a_721_47# SCE a_608_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_608_369# D a_504_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__einvn_8 A TE_B Z VGND VPWR VPB VNB
M1000 VPWR TE_B a_222_309# VPB phighvt w=940000u l=180000u
+  ad=1.4115e+12p pd=1.249e+07u as=2.5004e+12p ps=2.266e+07u
M1001 Z A a_222_309# VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=0p ps=0u
M1002 VPWR TE_B a_222_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Z A a_222_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_235_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.8005e+12p pd=1.724e+07u as=1.04325e+12p ps=9.71e+06u
M1005 a_222_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_222_309# A Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_27_47# a_235_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_235_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Z A a_235_47# VNB nshort w=650000u l=150000u
+  ad=8.645e+11p pd=7.86e+06u as=0p ps=0u
M1010 a_235_47# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_222_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR TE_B a_222_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Z A a_222_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR TE_B a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1015 VGND a_27_47# a_235_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_222_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_222_309# A Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_235_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Z A a_235_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_235_47# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_235_47# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Z A a_235_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Z A a_222_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND TE_B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1025 VGND a_27_47# a_235_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR TE_B a_222_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_222_309# A Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_235_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND a_27_47# a_235_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Z A a_235_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_222_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_222_309# A Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_235_47# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__nor4bb_4 D_N Y A B C_N VNB VPB VGND VPWR
M1000 Y a_207_47# a_331_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=1.41e+12p ps=1.282e+07u
M1001 a_1187_297# B a_797_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.43e+12p pd=1.286e+07u as=1.16e+12p ps=1.032e+07u
M1002 VPWR C_N a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u
M1003 a_207_47# D_N VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=2.223e+12p ps=1.984e+07u
M1004 Y a_27_297# VGND VNB nshort w=650000u l=150000u
+  ad=1.794e+12p pd=1.592e+07u as=0p ps=0u
M1005 VGND a_27_297# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C_N a_27_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.1125e+11p ps=1.95e+06u
M1007 VGND a_207_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_331_297# a_207_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_797_297# B a_1187_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_27_297# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_797_297# a_27_297# a_331_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y a_27_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y a_207_47# a_331_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1187_297# B a_797_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_331_297# a_27_297# a_797_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y a_207_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A a_1187_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_797_297# B a_1187_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_797_297# a_27_297# a_331_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1187_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_207_47# D_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=0p ps=0u
M1027 VGND a_207_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y a_207_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_331_297# a_207_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A a_1187_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1187_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_331_297# a_27_297# a_797_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o2bb2ai_1 Y A1_N A2_N B2 B1 VPB VNB VGND VPWR
M1000 a_120_297# A1_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=1.275e+12p ps=8.55e+06u
M1001 a_396_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=4.225e+11p pd=3.9e+06u as=3.8675e+11p ps=3.79e+06u
M1002 Y a_120_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.1e+11p pd=2.62e+06u as=0p ps=0u
M1003 VPWR B1 a_492_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1004 a_120_297# A2_N a_122_47# VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u
M1005 a_396_47# a_120_297# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1006 a_122_47# A1_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_492_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A2_N a_120_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B2 a_396_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__isobufsrc_4 A X SLEEP VNB VPB VGND VPWR
M1000 X a_459_21# a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=1.45e+12p ps=1.29e+07u
M1001 VPWR SLEEP a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=8.7e+11p pd=7.74e+06u as=0p ps=0u
M1002 VGND SLEEP X VNB nshort w=650000u l=150000u
+  ad=1.1505e+12p pd=1.134e+07u as=8.97e+11p ps=7.96e+06u
M1003 a_27_297# SLEEP VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_459_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_459_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR SLEEP a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND SLEEP X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_297# a_459_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A a_459_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1011 VGND A a_459_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.82e+11p ps=1.86e+06u
M1012 a_27_297# SLEEP VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_459_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_459_21# a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_459_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_297# a_459_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__bufbuf_8 A X VNB VPB VGND VPWR
M1000 VPWR a_338_47# X VPB phighvt w=1e+06u l=180000u
+  ad=2.0444e+12p pd=1.815e+07u as=1.16e+12p ps=1.032e+07u
M1001 VGND a_338_47# X VNB nshort w=650000u l=150000u
+  ad=1.4095e+12p pd=1.349e+07u as=8.645e+11p ps=7.86e+06u
M1002 VPWR a_338_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_338_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_338_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_224_297# a_338_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.095e+11p ps=3.86e+06u
M1006 X a_338_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_338_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_338_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_224_297# a_338_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.6e+11p ps=5.12e+06u
M1010 VPWR A a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1011 a_338_47# a_224_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_224_297# a_338_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_338_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_338_47# a_224_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_338_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_338_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_224_297# a_338_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1019 VPWR a_338_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_338_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_224_297# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1022 X a_338_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_338_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_224_297# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1025 X a_338_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__bufinv_8 A Y VNB VPB VGND VPWR
M1000 Y a_225_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=1.99e+12p ps=1.798e+07u
M1001 VPWR a_225_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND a_225_47# Y VNB nshort w=650000u l=150000u
+  ad=1.378e+12p pd=1.334e+07u as=8.645e+11p ps=7.86e+06u
M1003 VPWR a_225_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y a_225_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y a_225_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_225_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_117_297# a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.095e+11p ps=3.86e+06u
M1008 Y a_225_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_117_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1010 VPWR a_117_297# a_225_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.6e+11p ps=5.12e+06u
M1011 Y a_225_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y a_225_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_225_47# a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_225_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_117_297# A VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1016 a_225_47# a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_225_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_117_297# a_225_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_225_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y a_225_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_225_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y a_225_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_117_297# a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__muxb8to1_2 Z VGND VPWR VNB VPB D[2] D[1] S[7] S[6] S[5]
+ S[4] S[3] S[2] S[1] S[0] D[7] D[6] D[5] D[4] D[3] D[0]
M1000 VPWR D[2] a_1315_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.76e+12p pd=3.152e+07u as=8.211e+11p ps=7.41e+06u
M1001 VPWR D[3] a_2112_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.211e+11p ps=7.41e+06u
M1002 VPWR S[4] a_2854_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1003 a_27_297# D[0] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1004 Z a_1566_265# a_1315_297# VPB phighvt w=820000u l=180000u
+  ad=1.9024e+12p pd=1.776e+07u as=0p ps=0u
M1005 Z a_1989_47# a_2112_333# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_297# a_278_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_4565_47# S[7] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=1.9656e+12p ps=2.104e+07u
M1008 VPWR S[0] a_278_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1009 a_1989_47# S[3] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1010 Z S[5] a_3421_69# VNB nshort w=520000u l=150000u
+  ad=1.1232e+12p pd=1.264e+07u as=5.6745e+11p ps=5.52e+06u
M1011 a_4709_69# D[7] VGND VNB nshort w=650000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1012 a_2133_69# D[3] VGND VNB nshort w=650000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1013 Z a_278_265# a_27_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_2603_297# D[4] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1015 a_845_69# S[1] Z VNB nshort w=520000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1016 a_2603_297# a_2854_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_47# S[0] Z VNB nshort w=520000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1018 Z S[1] a_845_69# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_47# D[0] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Z S[0] a_27_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Z S[4] a_2603_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=5.6745e+11p ps=5.52e+06u
M1022 a_824_333# D[1] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1023 a_1989_47# S[3] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1024 a_3400_333# a_3277_47# Z VPB phighvt w=820000u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1025 a_3400_333# D[5] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_3421_69# S[5] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND D[7] a_4709_69# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_3277_47# S[5] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1029 a_3891_297# D[6] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1030 a_4688_333# D[7] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1031 VGND D[4] a_2603_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND S[4] a_2854_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1033 a_3891_297# a_4142_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR D[0] a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_701_47# S[1] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1036 VGND D[1] a_845_69# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR D[4] a_2603_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR D[5] a_3400_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR S[6] a_4142_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1040 a_824_333# a_701_47# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 Z a_2854_265# a_2603_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 Z a_3277_47# a_3400_333# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VGND S[0] a_278_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1044 a_2603_47# S[4] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_701_47# S[1] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1046 Z a_4142_265# a_3891_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VGND D[5] a_3421_69# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_2603_47# D[4] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 VPWR D[1] a_824_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1050 a_3277_47# S[5] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1051 a_845_69# D[1] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1052 Z S[3] a_2133_69# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1053 VGND D[0] a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1054 a_3421_69# D[5] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1055 Z S[7] a_4709_69# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1056 Z a_701_47# a_824_333# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1057 a_1315_47# D[2] VGND VNB nshort w=650000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1058 Z S[2] a_1315_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1059 Z S[6] a_3891_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=5.6745e+11p ps=5.52e+06u
M1060 a_1315_297# D[2] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1061 a_1315_297# a_1566_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1062 a_2112_333# a_1989_47# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1063 VGND D[2] a_1315_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1064 a_4688_333# a_4565_47# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1065 a_2133_69# S[3] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1066 a_4565_47# S[7] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1067 VPWR S[2] a_1566_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1068 a_2112_333# D[3] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1069 VPWR D[7] a_4688_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1070 VGND D[6] a_3891_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1071 a_4709_69# S[7] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1072 VPWR D[6] a_3891_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1073 Z a_4565_47# a_4688_333# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1074 a_3891_47# S[6] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1075 VGND S[6] a_4142_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1076 a_1315_47# S[2] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1077 VGND S[2] a_1566_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1078 VGND D[3] a_2133_69# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1079 a_3891_47# D[6] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__and2_1 VPWR VGND X B A VPB VNB
M1000 a_27_75# A VPWR VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=4.4565e+11p ps=4.17e+06u
M1001 X a_27_75# VGND VNB nshort w=650000u l=150000u
+  ad=2.3725e+11p pd=2.03e+06u as=2.406e+11p ps=2.11e+06u
M1002 X a_27_75# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.2e+11p pd=3.04e+06u as=0p ps=0u
M1003 VGND B a_123_75# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1004 VPWR B a_27_75# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_123_75# A a_27_75# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
.ends
.subckt sky130_fd_sc_hdll__o2bb2a_2 A1_N X A2_N B2 B1 VNB VPB VGND VPWR
M1000 a_321_369# A2_N a_313_47# VNB nshort w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=1.596e+11p ps=1.6e+06u
M1001 a_321_369# A1_N VPWR VPB phighvt w=640000u l=180000u
+  ad=3.652e+11p pd=2.86e+06u as=1.2558e+12p ps=9.86e+06u
M1002 a_627_47# B1 VGND VNB nshort w=420000u l=150000u
+  ad=2.541e+11p pd=2.89e+06u as=5.4595e+11p ps=5.41e+06u
M1003 X a_84_21# VGND VNB nshort w=650000u l=150000u
+  ad=2.08e+11p pd=1.94e+06u as=0p ps=0u
M1004 a_627_47# a_321_369# a_84_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1005 a_84_21# a_321_369# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.984e+11p pd=1.9e+06u as=0p ps=0u
M1006 VPWR B1 a_723_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=2.208e+11p ps=1.97e+06u
M1007 VPWR a_84_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1008 VPWR A2_N a_321_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_723_369# B2 a_84_21# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B2 a_627_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_84_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_313_47# A1_N VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_84_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__sedfxbp_1 VGND VPWR SCE Q D DE SCD Q_N CLK VPB VNB
M1000 a_1787_159# a_1611_413# VPWR VPB phighvt w=750000u l=180000u
+  ad=2.025e+11p pd=2.04e+06u as=1.93535e+12p ps=1.705e+07u
M1001 Q a_2266_413# VGND VNB nshort w=650000u l=150000u
+  ad=1.9825e+11p pd=1.91e+06u as=1.4487e+12p ps=1.404e+07u
M1002 a_211_363# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1003 a_2165_413# a_1787_159# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.365e+11p pd=1.49e+06u as=0p ps=0u
M1004 a_2266_413# a_27_47# a_2165_413# VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
M1005 VPWR DE a_455_324# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1006 VPWR CLK a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1007 a_319_47# a_851_264# a_779_47# VNB nshort w=420000u l=150000u
+  ad=2.478e+11p pd=2.86e+06u as=1.932e+11p ps=1.76e+06u
M1008 a_2181_47# a_1787_159# VGND VNB nshort w=420000u l=150000u
+  ad=1.356e+11p pd=1.51e+06u as=0p ps=0u
M1009 Q a_2266_413# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.15e+11p pd=2.63e+06u as=0p ps=0u
M1010 a_2266_413# a_211_363# a_2181_47# VNB nshort w=360000u l=150000u
+  ad=1.494e+11p pd=1.55e+06u as=0p ps=0u
M1011 a_1611_413# a_27_47# a_985_47# VNB nshort w=360000u l=150000u
+  ad=1.404e+11p pd=1.5e+06u as=6.015e+11p ps=4.57e+06u
M1012 a_985_47# a_955_21# a_1376_369# VPB phighvt w=640000u l=180000u
+  ad=4.837e+11p pd=4.13e+06u as=2.24e+11p ps=1.98e+06u
M1013 VGND SCE a_955_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1014 VGND a_2266_413# a_851_264# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1015 a_985_47# a_955_21# a_319_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Q_N a_851_264# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1017 VPWR SCE a_955_21# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.76e+11p ps=1.83e+06u
M1018 a_409_369# D a_319_47# VPB phighvt w=640000u l=180000u
+  ad=1.472e+11p pd=1.74e+06u as=3.84e+11p ps=3.76e+06u
M1019 a_985_47# SCE a_1373_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1020 VGND a_851_264# a_2391_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.32e+11p ps=1.49e+06u
M1021 a_787_369# DE VPWR VPB phighvt w=640000u l=180000u
+  ad=2.432e+11p pd=2.04e+06u as=0p ps=0u
M1022 a_319_47# a_851_264# a_787_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1611_413# a_211_363# a_985_47# VPB phighvt w=420000u l=180000u
+  ad=1.365e+11p pd=1.49e+06u as=0p ps=0u
M1024 VPWR a_1787_159# a_1712_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.617e+11p ps=1.61e+06u
M1025 VPWR a_455_324# a_409_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_985_47# SCE a_319_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Q_N a_851_264# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1028 a_1712_413# a_27_47# a_1611_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_2266_413# a_851_264# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1030 VGND DE a_455_324# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1031 a_779_47# a_455_324# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1376_369# SCD VPWR VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1034 a_1373_119# SCD VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR a_851_264# a_2360_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=2.058e+11p ps=1.82e+06u
M1036 VGND a_1787_159# a_1738_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.518e+11p ps=1.6e+06u
M1037 a_211_363# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1038 a_1738_47# a_211_363# a_1611_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_2391_47# a_27_47# a_2266_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_413_47# D a_319_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1041 VGND DE a_413_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_2360_413# a_211_363# a_2266_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_1787_159# a_1611_413# VGND VNB nshort w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a221oi_4 A2 Y C1 A1 B2 B1 VNB VPB VPWR VGND
M1000 a_511_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.69e+12p pd=2.338e+07u as=1.16e+12p ps=1.032e+07u
M1001 a_503_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=1.157e+12p pd=8.76e+06u as=1.48525e+12p ps=1.367e+07u
M1002 a_1375_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=7.67e+11p pd=7.56e+06u as=1.313e+12p ps=1.184e+07u
M1003 Y C1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=2.01e+12p ps=1.802e+07u
M1004 a_27_297# B1 a_511_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A2 a_511_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_1375_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y C1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A2 a_511_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1375_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_297# C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A1 a_1375_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_511_297# B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_511_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_511_297# B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND B2 a_503_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y C1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1375_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_297# B2 a_511_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A1 a_511_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND C1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_503_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y B1 a_503_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_511_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y C1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A2 a_1375_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_27_297# B1 a_511_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_503_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_27_297# C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_503_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_511_297# B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_511_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_511_297# B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND C1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_27_297# B2 a_511_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR A1 a_511_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND B2 a_503_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND A2 a_1375_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 Y B1 a_503_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 Y A1 a_1375_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__o22a_4 B2 B1 X A1 A2 VNB VPB VGND VPWR
M1000 VGND A1 a_524_47# VNB nshort w=650000u l=150000u
+  ad=9.425e+11p pd=9.4e+06u as=1.1115e+12p ps=9.92e+06u
M1001 X a_96_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=2.055e+12p ps=1.411e+07u
M1002 a_1006_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1003 a_614_297# B2 a_96_21# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=5.8e+11p ps=5.16e+06u
M1004 a_524_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_96_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_96_21# B2 a_614_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_96_21# VGND VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=0p ps=0u
M1008 VGND a_96_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_524_47# B1 a_96_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.835e+11p ps=3.78e+06u
M1010 a_96_21# B2 a_524_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A1 a_1006_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A2 a_524_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_614_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_96_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_96_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_524_47# B2 a_96_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1006_297# A2 a_96_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_96_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_96_21# B1 a_524_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_524_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_96_21# A2 a_1006_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_96_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR B1 a_614_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__a32oi_1 A2 Y A1 B2 B1 A3 VGND VPWR VPB VNB
M1000 a_27_297# B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=1.02e+12p pd=8.04e+06u as=2.9e+11p ps=2.58e+06u
M1001 Y B1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=3.445e+11p pd=2.36e+06u as=1.755e+11p ps=1.84e+06u
M1002 Y B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.6e+11p ps=5.12e+06u
M1004 a_423_47# A2 a_339_47# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=1.755e+11p ps=1.84e+06u
M1005 a_119_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.03e+11p ps=3.84e+06u
M1006 VGND A3 a_423_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A3 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_339_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__or3_2 A B X C VGND VPWR VPB VNB
M1000 VGND a_30_53# X VNB nshort w=650000u l=150000u
+  ad=6.469e+11p pd=5.71e+06u as=2.405e+11p ps=2.04e+06u
M1001 a_120_297# C a_30_53# VPB phighvt w=420000u l=180000u
+  ad=9.66e+10p pd=1.3e+06u as=1.134e+11p ps=1.38e+06u
M1002 VGND A a_30_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.646e+11p ps=2.94e+06u
M1003 VPWR a_30_53# X VPB phighvt w=1e+06u l=180000u
+  ad=8.257e+11p pd=5.75e+06u as=2.9e+11p ps=2.58e+06u
M1004 a_30_53# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_30_53# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A a_202_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1007 X a_30_53# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND C a_30_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_202_297# B a_120_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
.subckt sky130_fd_sc_hdll__tap VPWR VGND
Xsky130_fd_sc_hdll__o22ai_2_0 sky130_fd_sc_hdll__o22ai_2_0/B2 sky130_fd_sc_hdll__o22ai_2_0/B1
+ sky130_fd_sc_hdll__o22ai_2_0/Y sky130_fd_sc_hdll__o22ai_2_0/A1 sky130_fd_sc_hdll__o22ai_2_0/A2
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__o22ai_2
Xsky130_fd_sc_hdll__nand2_1_0 sky130_fd_sc_hdll__nand2_1_0/Y sky130_fd_sc_hdll__nand2_1_0/B
+ sky130_fd_sc_hdll__nand2_1_0/A VPWR VGND VGND VPWR sky130_fd_sc_hdll__nand2_1
Xsky130_fd_sc_hdll__nor3_4_0 sky130_fd_sc_hdll__nor3_4_0/A sky130_fd_sc_hdll__nor3_4_0/C
+ sky130_fd_sc_hdll__nor3_4_0/B sky130_fd_sc_hdll__nor3_4_0/Y VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__nor3_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_8 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a21bo_1_0 sky130_fd_sc_hdll__a21bo_1_0/X sky130_fd_sc_hdll__a21bo_1_0/A1
+ sky130_fd_sc_hdll__a21bo_1_0/B1_N sky130_fd_sc_hdll__a21bo_1_0/A2 VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__a21bo_1
Xsky130_fd_sc_hdll__nand2b_2_0 sky130_fd_sc_hdll__nand2b_2_0/B sky130_fd_sc_hdll__nand2b_2_0/Y
+ sky130_fd_sc_hdll__nand2b_2_0/A_N VGND VPWR VGND VPWR sky130_fd_sc_hdll__nand2b_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_305 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_316 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_19 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a31oi_1_0 VGND VPWR sky130_fd_sc_hdll__a31oi_1_0/Y sky130_fd_sc_hdll__a31oi_1_0/B1
+ sky130_fd_sc_hdll__a31oi_1_0/A2 sky130_fd_sc_hdll__a31oi_1_0/A1 sky130_fd_sc_hdll__a31oi_1_0/A3
+ VPWR VGND sky130_fd_sc_hdll__a31oi_1
Xsky130_fd_sc_hdll__mux2i_1_0 sky130_fd_sc_hdll__mux2i_1_0/A1 sky130_fd_sc_hdll__mux2i_1_0/S
+ sky130_fd_sc_hdll__mux2i_1_0/A0 sky130_fd_sc_hdll__mux2i_1_0/Y VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__mux2i_1
Xsky130_fd_sc_hdll__clkbuf_16_0 sky130_fd_sc_hdll__clkbuf_16_0/X sky130_fd_sc_hdll__clkbuf_16_0/A
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__clkbuf_16
Xsky130_fd_sc_hdll__o211ai_2_0 sky130_fd_sc_hdll__o211ai_2_0/A1 sky130_fd_sc_hdll__o211ai_2_0/A2
+ sky130_fd_sc_hdll__o211ai_2_0/B1 sky130_fd_sc_hdll__o211ai_2_0/Y sky130_fd_sc_hdll__o211ai_2_0/C1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o211ai_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_102 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_113 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_124 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_135 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_146 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_157 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_179 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_168 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__or2b_1_0 sky130_fd_sc_hdll__or2b_1_0/A sky130_fd_sc_hdll__or2b_1_0/B_N
+ sky130_fd_sc_hdll__or2b_1_0/X VGND VPWR VGND VPWR sky130_fd_sc_hdll__or2b_1
Xsky130_fd_sc_hdll__dlrtn_1_0 sky130_fd_sc_hdll__dlrtn_1_0/RESET_B sky130_fd_sc_hdll__dlrtn_1_0/D
+ sky130_fd_sc_hdll__dlrtn_1_0/GATE_N sky130_fd_sc_hdll__dlrtn_1_0/Q VGND VPWR VPWR
+ VGND sky130_fd_sc_hdll__dlrtn_1
Xsky130_fd_sc_hdll__clkmux2_2_0 VGND VPWR sky130_fd_sc_hdll__clkmux2_2_0/S sky130_fd_sc_hdll__clkmux2_2_0/A1
+ sky130_fd_sc_hdll__clkmux2_2_0/A0 sky130_fd_sc_hdll__clkmux2_2_0/X VPWR VGND sky130_fd_sc_hdll__clkmux2_2
Xsky130_fd_sc_hdll__or2_8_0 sky130_fd_sc_hdll__or2_8_0/X sky130_fd_sc_hdll__or2_8_0/A
+ sky130_fd_sc_hdll__or2_8_0/B VGND VPWR VGND VPWR sky130_fd_sc_hdll__or2_8
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_9 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o21ai_2_0 sky130_fd_sc_hdll__o21ai_2_0/B1 sky130_fd_sc_hdll__o21ai_2_0/Y
+ sky130_fd_sc_hdll__o21ai_2_0/A2 sky130_fd_sc_hdll__o21ai_2_0/A1 VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__o21ai_2
Xsky130_fd_sc_hdll__and3_4_0 sky130_fd_sc_hdll__and3_4_0/A sky130_fd_sc_hdll__and3_4_0/B
+ sky130_fd_sc_hdll__and3_4_0/C sky130_fd_sc_hdll__and3_4_0/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__and3_4
Xsky130_fd_sc_hdll__clkbuf_4_0 sky130_fd_sc_hdll__clkbuf_4_0/X sky130_fd_sc_hdll__clkbuf_4_0/A
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__clkbuf_4
Xsky130_fd_sc_hdll__clkinv_4_0 sky130_fd_sc_hdll__clkinv_4_0/A sky130_fd_sc_hdll__clkinv_4_0/Y
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__clkinv_4
Xsky130_fd_sc_hdll__sdfstp_4_0 sky130_fd_sc_hdll__sdfstp_4_0/CLK sky130_fd_sc_hdll__sdfstp_4_0/D
+ sky130_fd_sc_hdll__sdfstp_4_0/SCD sky130_fd_sc_hdll__sdfstp_4_0/Q sky130_fd_sc_hdll__sdfstp_4_0/SCE
+ sky130_fd_sc_hdll__sdfstp_4_0/SET_B VPWR VGND VPWR VGND sky130_fd_sc_hdll__sdfstp_4
Xsky130_fd_sc_hdll__a2bb2oi_1_0 sky130_fd_sc_hdll__a2bb2oi_1_0/A1_N sky130_fd_sc_hdll__a2bb2oi_1_0/Y
+ VGND VPWR sky130_fd_sc_hdll__a2bb2oi_1_0/B2 sky130_fd_sc_hdll__a2bb2oi_1_0/B1 sky130_fd_sc_hdll__a2bb2oi_1_0/A2_N
+ VPWR VGND sky130_fd_sc_hdll__a2bb2oi_1
Xsky130_fd_sc_hdll__nor4bb_2_0 sky130_fd_sc_hdll__nor4bb_2_0/D_N sky130_fd_sc_hdll__nor4bb_2_0/C_N
+ sky130_fd_sc_hdll__nor4bb_2_0/A sky130_fd_sc_hdll__nor4bb_2_0/Y sky130_fd_sc_hdll__nor4bb_2_0/B
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nor4bb_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_306 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_317 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__isobufsrc_2_0 sky130_fd_sc_hdll__isobufsrc_2_0/A sky130_fd_sc_hdll__isobufsrc_2_0/SLEEP
+ sky130_fd_sc_hdll__isobufsrc_2_0/X VPWR VGND VGND VPWR sky130_fd_sc_hdll__isobufsrc_2
Xsky130_fd_sc_hdll__sdfxbp_1_0 VGND VPWR sky130_fd_sc_hdll__sdfxbp_1_0/SCD sky130_fd_sc_hdll__sdfxbp_1_0/Q_N
+ sky130_fd_sc_hdll__sdfxbp_1_0/D sky130_fd_sc_hdll__sdfxbp_1_0/SCE sky130_fd_sc_hdll__sdfxbp_1_0/CLK
+ sky130_fd_sc_hdll__sdfxbp_1_0/Q VGND VPWR sky130_fd_sc_hdll__sdfxbp_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_103 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_114 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_125 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_136 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_147 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_158 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_169 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nor2b_1_0 sky130_fd_sc_hdll__nor2b_1_0/B_N sky130_fd_sc_hdll__nor2b_1_0/Y
+ sky130_fd_sc_hdll__nor2b_1_0/A VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor2b_1
Xsky130_fd_sc_hdll__a21boi_4_0 sky130_fd_sc_hdll__a21boi_4_0/Y sky130_fd_sc_hdll__a21boi_4_0/A1
+ sky130_fd_sc_hdll__a21boi_4_0/B1_N sky130_fd_sc_hdll__a21boi_4_0/A2 VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__a21boi_4
Xsky130_fd_sc_hdll__nand3_4_0 sky130_fd_sc_hdll__nand3_4_0/Y sky130_fd_sc_hdll__nand3_4_0/A
+ sky130_fd_sc_hdll__nand3_4_0/B sky130_fd_sc_hdll__nand3_4_0/C VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__nand3_4
Xsky130_fd_sc_hdll__mux2_4_0 sky130_fd_sc_hdll__mux2_4_0/X sky130_fd_sc_hdll__mux2_4_0/S
+ sky130_fd_sc_hdll__mux2_4_0/A0 sky130_fd_sc_hdll__mux2_4_0/A1 VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__mux2_4
Xsky130_fd_sc_hdll__and2b_4_0 sky130_fd_sc_hdll__and2b_4_0/B sky130_fd_sc_hdll__and2b_4_0/X
+ sky130_fd_sc_hdll__and2b_4_0/A_N VGND VPWR VGND VPWR sky130_fd_sc_hdll__and2b_4
Xsky130_fd_sc_hdll__o22a_2_0 sky130_fd_sc_hdll__o22a_2_0/A2 sky130_fd_sc_hdll__o22a_2_0/X
+ sky130_fd_sc_hdll__o22a_2_0/B1 sky130_fd_sc_hdll__o22a_2_0/A1 sky130_fd_sc_hdll__o22a_2_0/B2
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o22a_2
Xsky130_fd_sc_hdll__a221oi_2_0 sky130_fd_sc_hdll__a221oi_2_0/B2 sky130_fd_sc_hdll__a221oi_2_0/C1
+ sky130_fd_sc_hdll__a221oi_2_0/A2 sky130_fd_sc_hdll__a221oi_2_0/A1 sky130_fd_sc_hdll__a221oi_2_0/B1
+ sky130_fd_sc_hdll__a221oi_2_0/Y VGND VPWR VGND VPWR sky130_fd_sc_hdll__a221oi_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_307 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_318 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__sdfrtp_4_0 VPWR VGND sky130_fd_sc_hdll__sdfrtp_4_0/RESET_B VPWR
+ VGND sky130_fd_sc_hdll__sdfrtp_4_0/SCE sky130_fd_sc_hdll__sdfrtp_4_0/SCD sky130_fd_sc_hdll__sdfrtp_4_0/D
+ sky130_fd_sc_hdll__sdfrtp_4_0/CLK sky130_fd_sc_hdll__sdfrtp_4_0/Q sky130_fd_sc_hdll__sdfrtp_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_104 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_115 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_126 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_137 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_148 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_159 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__and4b_1_0 VGND VPWR sky130_fd_sc_hdll__and4b_1_0/C sky130_fd_sc_hdll__and4b_1_0/A_N
+ sky130_fd_sc_hdll__and4b_1_0/X sky130_fd_sc_hdll__and4b_1_0/D sky130_fd_sc_hdll__and4b_1_0/B
+ VPWR VGND sky130_fd_sc_hdll__and4b_1
Xsky130_fd_sc_hdll__probe_p_8_0 sky130_fd_sc_hdll__probe_p_8_0/X sky130_fd_sc_hdll__probe_p_8_0/A
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__probe_p_8
Xsky130_fd_sc_hdll__o32ai_4_0 sky130_fd_sc_hdll__o32ai_4_0/A1 sky130_fd_sc_hdll__o32ai_4_0/A2
+ sky130_fd_sc_hdll__o32ai_4_0/A3 sky130_fd_sc_hdll__o32ai_4_0/B1 sky130_fd_sc_hdll__o32ai_4_0/Y
+ sky130_fd_sc_hdll__o32ai_4_0/B2 VGND VPWR VGND VPWR sky130_fd_sc_hdll__o32ai_4
Xsky130_fd_sc_hdll__nor3_2_0 sky130_fd_sc_hdll__nor3_2_0/C sky130_fd_sc_hdll__nor3_2_0/Y
+ sky130_fd_sc_hdll__nor3_2_0/A sky130_fd_sc_hdll__nor3_2_0/B VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__nor3_2
Xsky130_fd_sc_hdll__xor2_4_0 sky130_fd_sc_hdll__xor2_4_0/X sky130_fd_sc_hdll__xor2_4_0/B
+ sky130_fd_sc_hdll__xor2_4_0/A VGND VPWR VGND VPWR sky130_fd_sc_hdll__xor2_4
Xsky130_fd_sc_hdll__or3b_4_0 sky130_fd_sc_hdll__or3b_4_0/A sky130_fd_sc_hdll__or3b_4_0/B
+ sky130_fd_sc_hdll__or3b_4_0/C_N sky130_fd_sc_hdll__or3b_4_0/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__or3b_4
Xsky130_fd_sc_hdll__o21ba_4_0 sky130_fd_sc_hdll__o21ba_4_0/B1_N sky130_fd_sc_hdll__o21ba_4_0/A1
+ sky130_fd_sc_hdll__o21ba_4_0/A2 sky130_fd_sc_hdll__o21ba_4_0/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__o21ba_4
Xsky130_fd_sc_hdll__a31o_1_0 sky130_fd_sc_hdll__a31o_1_0/A2 sky130_fd_sc_hdll__a31o_1_0/B1
+ sky130_fd_sc_hdll__a31o_1_0/A1 sky130_fd_sc_hdll__a31o_1_0/A3 sky130_fd_sc_hdll__a31o_1_0/X
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__a31o_1
Xsky130_fd_sc_hdll__xnor3_1_0 sky130_fd_sc_hdll__xnor3_1_0/X sky130_fd_sc_hdll__xnor3_1_0/B
+ sky130_fd_sc_hdll__xnor3_1_0/C sky130_fd_sc_hdll__xnor3_1_0/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__xnor3_1
Xsky130_fd_sc_hdll__or4bb_4_0 sky130_fd_sc_hdll__or4bb_4_0/D_N sky130_fd_sc_hdll__or4bb_4_0/B
+ sky130_fd_sc_hdll__or4bb_4_0/A sky130_fd_sc_hdll__or4bb_4_0/C_N sky130_fd_sc_hdll__or4bb_4_0/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__or4bb_4
Xsky130_fd_sc_hdll__probec_p_8_0 sky130_fd_sc_hdll__probec_p_8_0/X sky130_fd_sc_hdll__probec_p_8_0/A
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__probec_p_8
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_308 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_319 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_105 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_116 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_127 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_138 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_149 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nor3b_4_0 sky130_fd_sc_hdll__nor3b_4_0/A sky130_fd_sc_hdll__nor3b_4_0/C_N
+ sky130_fd_sc_hdll__nor3b_4_0/B sky130_fd_sc_hdll__nor3b_4_0/Y VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__nor3b_4
Xsky130_fd_sc_hdll__o221ai_4_0 sky130_fd_sc_hdll__o221ai_4_0/B1 sky130_fd_sc_hdll__o221ai_4_0/B2
+ sky130_fd_sc_hdll__o221ai_4_0/A2 sky130_fd_sc_hdll__o221ai_4_0/C1 sky130_fd_sc_hdll__o221ai_4_0/Y
+ sky130_fd_sc_hdll__o221ai_4_0/A1 VGND VPWR VGND VPWR sky130_fd_sc_hdll__o221ai_4
Xsky130_fd_sc_hdll__or2_6_0 sky130_fd_sc_hdll__or2_6_0/X sky130_fd_sc_hdll__or2_6_0/A
+ sky130_fd_sc_hdll__or2_6_0/B VGND VPWR VGND VPWR sky130_fd_sc_hdll__or2_6
Xsky130_fd_sc_hdll__o31ai_4_0 sky130_fd_sc_hdll__o31ai_4_0/A3 sky130_fd_sc_hdll__o31ai_4_0/A2
+ sky130_fd_sc_hdll__o31ai_4_0/A1 sky130_fd_sc_hdll__o31ai_4_0/Y sky130_fd_sc_hdll__o31ai_4_0/B1
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__o31ai_4
Xsky130_fd_sc_hdll__and3_2_0 sky130_fd_sc_hdll__and3_2_0/B sky130_fd_sc_hdll__and3_2_0/X
+ sky130_fd_sc_hdll__and3_2_0/A sky130_fd_sc_hdll__and3_2_0/C VPWR VGND VPWR VGND
+ sky130_fd_sc_hdll__and3_2
Xsky130_fd_sc_hdll__clkbuf_2_0 VPWR VGND VPWR VGND sky130_fd_sc_hdll__clkbuf_2_0/A
+ sky130_fd_sc_hdll__clkbuf_2_0/X sky130_fd_sc_hdll__clkbuf_2
Xsky130_fd_sc_hdll__clkinv_2_0 sky130_fd_sc_hdll__clkinv_2_0/Y sky130_fd_sc_hdll__clkinv_2_0/A
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__clkinv_2
Xsky130_fd_sc_hdll__sdfstp_2_0 sky130_fd_sc_hdll__sdfstp_2_0/Q sky130_fd_sc_hdll__sdfstp_2_0/SCD
+ sky130_fd_sc_hdll__sdfstp_2_0/D sky130_fd_sc_hdll__sdfstp_2_0/CLK sky130_fd_sc_hdll__sdfstp_2_0/SET_B
+ sky130_fd_sc_hdll__sdfstp_2_0/SCE VGND VPWR VPWR VGND sky130_fd_sc_hdll__sdfstp_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_309 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a211o_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a211o_1_0/X sky130_fd_sc_hdll__a211o_1_0/A2
+ sky130_fd_sc_hdll__a211o_1_0/B1 sky130_fd_sc_hdll__a211o_1_0/A1 sky130_fd_sc_hdll__a211o_1_0/C1
+ sky130_fd_sc_hdll__a211o_1
Xsky130_fd_sc_hdll__nor2_8_0 sky130_fd_sc_hdll__nor2_8_0/Y sky130_fd_sc_hdll__nor2_8_0/A
+ sky130_fd_sc_hdll__nor2_8_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor2_8
Xsky130_fd_sc_hdll__a21o_1_0 sky130_fd_sc_hdll__a21o_1_0/A2 sky130_fd_sc_hdll__a21o_1_0/A1
+ sky130_fd_sc_hdll__a21o_1_0/B1 sky130_fd_sc_hdll__a21o_1_0/X VPWR VGND VPWR VGND
+ sky130_fd_sc_hdll__a21o_1
Xsky130_fd_sc_hdll__einvn_4_0 sky130_fd_sc_hdll__einvn_4_0/TE_B sky130_fd_sc_hdll__einvn_4_0/Z
+ sky130_fd_sc_hdll__einvn_4_0/A VGND VPWR VPWR VGND sky130_fd_sc_hdll__einvn_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_106 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_117 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_128 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_139 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nand2_16_0 sky130_fd_sc_hdll__nand2_16_0/Y sky130_fd_sc_hdll__nand2_16_0/A
+ sky130_fd_sc_hdll__nand2_16_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__nand2_16
Xsky130_fd_sc_hdll__buf_16_0 sky130_fd_sc_hdll__buf_16_0/A sky130_fd_sc_hdll__buf_16_0/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__buf_16
Xsky130_fd_sc_hdll__a21boi_2_0 VGND VPWR VPWR VGND sky130_fd_sc_hdll__a21boi_2_0/B1_N
+ sky130_fd_sc_hdll__a21boi_2_0/A2 sky130_fd_sc_hdll__a21boi_2_0/A1 sky130_fd_sc_hdll__a21boi_2_0/Y
+ sky130_fd_sc_hdll__a21boi_2
Xsky130_fd_sc_hdll__nand3_2_0 sky130_fd_sc_hdll__nand3_2_0/A sky130_fd_sc_hdll__nand3_2_0/Y
+ sky130_fd_sc_hdll__nand3_2_0/B sky130_fd_sc_hdll__nand3_2_0/C VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__nand3_2
Xsky130_fd_sc_hdll__fill_4_0 VGND VPWR VPWR VGND sky130_fd_sc_hdll__fill_4
Xsky130_fd_sc_hdll__einvp_1_0 sky130_fd_sc_hdll__einvp_1_0/TE sky130_fd_sc_hdll__einvp_1_0/A
+ sky130_fd_sc_hdll__einvp_1_0/Z VPWR VGND VPWR VGND sky130_fd_sc_hdll__einvp_1
Xsky130_fd_sc_hdll__a32o_4_0 sky130_fd_sc_hdll__a32o_4_0/A3 sky130_fd_sc_hdll__a32o_4_0/X
+ sky130_fd_sc_hdll__a32o_4_0/B1 sky130_fd_sc_hdll__a32o_4_0/B2 sky130_fd_sc_hdll__a32o_4_0/A1
+ sky130_fd_sc_hdll__a32o_4_0/A2 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a32o_4
Xsky130_fd_sc_hdll__mux2_2_0 VGND VPWR sky130_fd_sc_hdll__mux2_2_0/A1 sky130_fd_sc_hdll__mux2_2_0/A0
+ sky130_fd_sc_hdll__mux2_2_0/S sky130_fd_sc_hdll__mux2_2_0/X VPWR VGND sky130_fd_sc_hdll__mux2_2
Xsky130_fd_sc_hdll__and2b_2_0 VGND VPWR VPWR VGND sky130_fd_sc_hdll__and2b_2_0/X sky130_fd_sc_hdll__and2b_2_0/B
+ sky130_fd_sc_hdll__and2b_2_0/A_N sky130_fd_sc_hdll__and2b_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_107 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_118 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_129 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__sdfrtp_2_0 sky130_fd_sc_hdll__sdfrtp_2_0/RESET_B VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__sdfrtp_2_0/Q sky130_fd_sc_hdll__sdfrtp_2_0/SCE sky130_fd_sc_hdll__sdfrtp_2_0/SCD
+ sky130_fd_sc_hdll__sdfrtp_2_0/D sky130_fd_sc_hdll__sdfrtp_2_0/CLK sky130_fd_sc_hdll__sdfrtp_2
Xsky130_fd_sc_hdll__and2_8_0 sky130_fd_sc_hdll__and2_8_0/X sky130_fd_sc_hdll__and2_8_0/B
+ sky130_fd_sc_hdll__and2_8_0/A VGND VPWR VGND VPWR sky130_fd_sc_hdll__and2_8
Xsky130_fd_sc_hdll__a22oi_4_0 sky130_fd_sc_hdll__a22oi_4_0/A2 sky130_fd_sc_hdll__a22oi_4_0/B2
+ sky130_fd_sc_hdll__a22oi_4_0/A1 sky130_fd_sc_hdll__a22oi_4_0/B1 sky130_fd_sc_hdll__a22oi_4_0/Y
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__a22oi_4
Xsky130_fd_sc_hdll__muxb4to1_4_0 VPWR VGND VGND VPWR sky130_fd_sc_hdll__muxb4to1_4_0/Z
+ sky130_fd_sc_hdll__muxb4to1_4_0/S[0] sky130_fd_sc_hdll__muxb4to1_4_0/S[1] sky130_fd_sc_hdll__muxb4to1_4_0/D[1]
+ sky130_fd_sc_hdll__muxb4to1_4_0/D[2] sky130_fd_sc_hdll__muxb4to1_4_0/S[2] sky130_fd_sc_hdll__muxb4to1_4_0/S[3]
+ sky130_fd_sc_hdll__muxb4to1_4_0/D[3] sky130_fd_sc_hdll__muxb4to1_4_0/D[0] sky130_fd_sc_hdll__muxb4to1_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_290 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o32ai_2_0 sky130_fd_sc_hdll__o32ai_2_0/A1 sky130_fd_sc_hdll__o32ai_2_0/B1
+ sky130_fd_sc_hdll__o32ai_2_0/A2 sky130_fd_sc_hdll__o32ai_2_0/A3 sky130_fd_sc_hdll__o32ai_2_0/Y
+ sky130_fd_sc_hdll__o32ai_2_0/B2 VPWR VGND VGND VPWR sky130_fd_sc_hdll__o32ai_2
Xsky130_fd_sc_hdll__o221a_4_0 sky130_fd_sc_hdll__o221a_4_0/C1 sky130_fd_sc_hdll__o221a_4_0/A1
+ sky130_fd_sc_hdll__o221a_4_0/A2 sky130_fd_sc_hdll__o221a_4_0/B1 sky130_fd_sc_hdll__o221a_4_0/B2
+ sky130_fd_sc_hdll__o221a_4_0/X VGND VPWR VGND VPWR sky130_fd_sc_hdll__o221a_4
Xsky130_fd_sc_hdll__or3b_2_0 sky130_fd_sc_hdll__or3b_2_0/A sky130_fd_sc_hdll__or3b_2_0/B
+ sky130_fd_sc_hdll__or3b_2_0/C_N sky130_fd_sc_hdll__or3b_2_0/X VPWR VGND VPWR VGND
+ sky130_fd_sc_hdll__or3b_2
Xsky130_fd_sc_hdll__xor2_2_0 sky130_fd_sc_hdll__xor2_2_0/B VPWR VGND sky130_fd_sc_hdll__xor2_2_0/X
+ sky130_fd_sc_hdll__xor2_2_0/A VPWR VGND sky130_fd_sc_hdll__xor2_2
Xsky130_fd_sc_hdll__o21ba_2_0 sky130_fd_sc_hdll__o21ba_2_0/B1_N sky130_fd_sc_hdll__o21ba_2_0/A1
+ sky130_fd_sc_hdll__o21ba_2_0/X sky130_fd_sc_hdll__o21ba_2_0/A2 VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__o21ba_2
Xsky130_fd_sc_hdll__or4bb_2_0 sky130_fd_sc_hdll__or4bb_2_0/A sky130_fd_sc_hdll__or4bb_2_0/X
+ sky130_fd_sc_hdll__or4bb_2_0/B sky130_fd_sc_hdll__or4bb_2_0/D_N sky130_fd_sc_hdll__or4bb_2_0/C_N
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__or4bb_2
Xsky130_fd_sc_hdll__dlxtn_4_0 sky130_fd_sc_hdll__dlxtn_4_0/D sky130_fd_sc_hdll__dlxtn_4_0/GATE_N
+ sky130_fd_sc_hdll__dlxtn_4_0/Q VGND VPWR VPWR VGND sky130_fd_sc_hdll__dlxtn_4
Xsky130_fd_sc_hdll__nand2_8_0 sky130_fd_sc_hdll__nand2_8_0/A sky130_fd_sc_hdll__nand2_8_0/B
+ sky130_fd_sc_hdll__nand2_8_0/Y VGND VPWR VGND VPWR sky130_fd_sc_hdll__nand2_8
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_108 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_119 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o21bai_4_0 sky130_fd_sc_hdll__o21bai_4_0/Y sky130_fd_sc_hdll__o21bai_4_0/B1_N
+ sky130_fd_sc_hdll__o21bai_4_0/A1 sky130_fd_sc_hdll__o21bai_4_0/A2 VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__o21bai_4
Xsky130_fd_sc_hdll__a22o_4_0 sky130_fd_sc_hdll__a22o_4_0/B1 sky130_fd_sc_hdll__a22o_4_0/B2
+ sky130_fd_sc_hdll__a22o_4_0/X sky130_fd_sc_hdll__a22o_4_0/A2 sky130_fd_sc_hdll__a22o_4_0/A1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__a22o_4
Xsky130_fd_sc_hdll__dlygate4sd2_1_0 sky130_fd_sc_hdll__dlygate4sd2_1_0/A sky130_fd_sc_hdll__dlygate4sd2_1_0/X
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__dlygate4sd2_1
Xsky130_fd_sc_hdll__nand4bb_1_0 sky130_fd_sc_hdll__nand4bb_1_0/C sky130_fd_sc_hdll__nand4bb_1_0/D
+ sky130_fd_sc_hdll__nand4bb_1_0/A_N sky130_fd_sc_hdll__nand4bb_1_0/Y sky130_fd_sc_hdll__nand4bb_1_0/B_N
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__nand4bb_1
Xsky130_fd_sc_hdll__clkbuf_12_0 sky130_fd_sc_hdll__clkbuf_12_0/A sky130_fd_sc_hdll__clkbuf_12_0/X
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__clkbuf_12
Xsky130_fd_sc_hdll__nor3b_2_0 sky130_fd_sc_hdll__nor3b_2_0/C_N sky130_fd_sc_hdll__nor3b_2_0/Y
+ sky130_fd_sc_hdll__nor3b_2_0/A sky130_fd_sc_hdll__nor3b_2_0/B VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__nor3b_2
Xsky130_fd_sc_hdll__muxb16to1_1_0 sky130_fd_sc_hdll__muxb16to1_1_0/Z VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__muxb16to1_1_0/D[0] sky130_fd_sc_hdll__muxb16to1_1_0/S[12]
+ sky130_fd_sc_hdll__muxb16to1_1_0/S[13] sky130_fd_sc_hdll__muxb16to1_1_0/S[8] sky130_fd_sc_hdll__muxb16to1_1_0/S[9]
+ sky130_fd_sc_hdll__muxb16to1_1_0/S[10] sky130_fd_sc_hdll__muxb16to1_1_0/S[11] sky130_fd_sc_hdll__muxb16to1_1_0/S[14]
+ sky130_fd_sc_hdll__muxb16to1_1_0/S[15] sky130_fd_sc_hdll__muxb16to1_1_0/D[12] sky130_fd_sc_hdll__muxb16to1_1_0/D[9]
+ sky130_fd_sc_hdll__muxb16to1_1_0/D[10] sky130_fd_sc_hdll__muxb16to1_1_0/D[13] sky130_fd_sc_hdll__muxb16to1_1_0/D[14]
+ sky130_fd_sc_hdll__muxb16to1_1_0/D[15] sky130_fd_sc_hdll__muxb16to1_1_0/D[8] sky130_fd_sc_hdll__muxb16to1_1_0/D[11]
+ sky130_fd_sc_hdll__muxb16to1_1_0/S[0] sky130_fd_sc_hdll__muxb16to1_1_0/S[1] sky130_fd_sc_hdll__muxb16to1_1_0/D[1]
+ sky130_fd_sc_hdll__muxb16to1_1_0/D[2] sky130_fd_sc_hdll__muxb16to1_1_0/S[2] sky130_fd_sc_hdll__muxb16to1_1_0/S[3]
+ sky130_fd_sc_hdll__muxb16to1_1_0/D[4] sky130_fd_sc_hdll__muxb16to1_1_0/S[4] sky130_fd_sc_hdll__muxb16to1_1_0/S[5]
+ sky130_fd_sc_hdll__muxb16to1_1_0/D[5] sky130_fd_sc_hdll__muxb16to1_1_0/D[6] sky130_fd_sc_hdll__muxb16to1_1_0/S[6]
+ sky130_fd_sc_hdll__muxb16to1_1_0/S[7] sky130_fd_sc_hdll__muxb16to1_1_0/D[7] sky130_fd_sc_hdll__muxb16to1_1_0/D[3]
+ sky130_fd_sc_hdll__muxb16to1_1
Xsky130_fd_sc_hdll__o221ai_2_0 sky130_fd_sc_hdll__o221ai_2_0/B1 sky130_fd_sc_hdll__o221ai_2_0/B2
+ sky130_fd_sc_hdll__o221ai_2_0/Y sky130_fd_sc_hdll__o221ai_2_0/A2 sky130_fd_sc_hdll__o221ai_2_0/A1
+ sky130_fd_sc_hdll__o221ai_2_0/C1 VGND VPWR VGND VPWR sky130_fd_sc_hdll__o221ai_2
Xsky130_fd_sc_hdll__ebufn_1_0 sky130_fd_sc_hdll__ebufn_1_0/Z sky130_fd_sc_hdll__ebufn_1_0/TE_B
+ sky130_fd_sc_hdll__ebufn_1_0/A VGND VPWR VPWR VGND sky130_fd_sc_hdll__ebufn_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_291 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_280 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__or2_4_0 sky130_fd_sc_hdll__or2_4_0/X sky130_fd_sc_hdll__or2_4_0/A
+ sky130_fd_sc_hdll__or2_4_0/B VGND VPWR VGND VPWR sky130_fd_sc_hdll__or2_4
Xsky130_fd_sc_hdll__a21oi_4_0 sky130_fd_sc_hdll__a21oi_4_0/B1 sky130_fd_sc_hdll__a21oi_4_0/A2
+ sky130_fd_sc_hdll__a21oi_4_0/A1 sky130_fd_sc_hdll__a21oi_4_0/Y VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__a21oi_4
Xsky130_fd_sc_hdll__o31ai_2_0 sky130_fd_sc_hdll__o31ai_2_0/A1 sky130_fd_sc_hdll__o31ai_2_0/Y
+ sky130_fd_sc_hdll__o31ai_2_0/B1 sky130_fd_sc_hdll__o31ai_2_0/A3 sky130_fd_sc_hdll__o31ai_2_0/A2
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__o31ai_2
Xsky130_fd_sc_hdll__o211a_4_0 sky130_fd_sc_hdll__o211a_4_0/A1 sky130_fd_sc_hdll__o211a_4_0/X
+ sky130_fd_sc_hdll__o211a_4_0/C1 sky130_fd_sc_hdll__o211a_4_0/A2 sky130_fd_sc_hdll__o211a_4_0/B1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o211a_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_109 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__einvn_2_0 sky130_fd_sc_hdll__einvn_2_0/TE_B sky130_fd_sc_hdll__einvn_2_0/A
+ sky130_fd_sc_hdll__einvn_2_0/Z VPWR VGND VPWR VGND sky130_fd_sc_hdll__einvn_2
Xsky130_fd_sc_hdll__sdfsbp_1_0 sky130_fd_sc_hdll__sdfsbp_1_0/SCD sky130_fd_sc_hdll__sdfsbp_1_0/CLK
+ sky130_fd_sc_hdll__sdfsbp_1_0/Q_N sky130_fd_sc_hdll__sdfsbp_1_0/D sky130_fd_sc_hdll__sdfsbp_1_0/Q
+ VPWR VGND sky130_fd_sc_hdll__sdfsbp_1_0/SET_B sky130_fd_sc_hdll__sdfsbp_1_0/SCE
+ VPWR VGND sky130_fd_sc_hdll__sdfsbp_1
Xsky130_fd_sc_hdll__or4_1_0 sky130_fd_sc_hdll__or4_1_0/C sky130_fd_sc_hdll__or4_1_0/A
+ sky130_fd_sc_hdll__or4_1_0/X sky130_fd_sc_hdll__or4_1_0/B sky130_fd_sc_hdll__or4_1_0/D
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__or4_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_292 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_281 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_270 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__inputiso0n_1_0 VPWR VGND sky130_fd_sc_hdll__inputiso0n_1_0/X sky130_fd_sc_hdll__inputiso0n_1_0/SLEEP_B
+ sky130_fd_sc_hdll__inputiso0n_1_0/A VPWR VGND sky130_fd_sc_hdll__inputiso0n_1
Xsky130_fd_sc_hdll__fill_2_0 VGND VPWR VPWR VGND sky130_fd_sc_hdll__fill_2
Xsky130_fd_sc_hdll__and4bb_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__and4bb_1_0/A_N
+ sky130_fd_sc_hdll__and4bb_1_0/D sky130_fd_sc_hdll__and4bb_1_0/X sky130_fd_sc_hdll__and4bb_1_0/C
+ sky130_fd_sc_hdll__and4bb_1_0/B_N sky130_fd_sc_hdll__and4bb_1
Xsky130_fd_sc_hdll__clkinvlp_4_0 sky130_fd_sc_hdll__clkinvlp_4_0/A sky130_fd_sc_hdll__clkinvlp_4_0/Y
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__clkinvlp_4
Xsky130_fd_sc_hdll__a32o_2_0 sky130_fd_sc_hdll__a32o_2_0/B2 sky130_fd_sc_hdll__a32o_2_0/X
+ sky130_fd_sc_hdll__a32o_2_0/A2 sky130_fd_sc_hdll__a32o_2_0/A3 sky130_fd_sc_hdll__a32o_2_0/A1
+ sky130_fd_sc_hdll__a32o_2_0/B1 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a32o_2
Xsky130_fd_sc_hdll__nand3b_1_0 sky130_fd_sc_hdll__nand3b_1_0/B sky130_fd_sc_hdll__nand3b_1_0/C
+ sky130_fd_sc_hdll__nand3b_1_0/A_N sky130_fd_sc_hdll__nand3b_1_0/Y VPWR VGND VGND
+ VPWR sky130_fd_sc_hdll__nand3b_1
Xsky130_fd_sc_hdll__and2_6_0 sky130_fd_sc_hdll__and2_6_0/X sky130_fd_sc_hdll__and2_6_0/B
+ sky130_fd_sc_hdll__and2_6_0/A VGND VPWR VGND VPWR sky130_fd_sc_hdll__and2_6
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_293 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_282 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_271 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_260 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a22oi_2_0 sky130_fd_sc_hdll__a22oi_2_0/A1 sky130_fd_sc_hdll__a22oi_2_0/A2
+ sky130_fd_sc_hdll__a22oi_2_0/B1 sky130_fd_sc_hdll__a22oi_2_0/B2 sky130_fd_sc_hdll__a22oi_2_0/Y
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__a22oi_2
Xsky130_fd_sc_hdll__muxb4to1_2_0 VGND VPWR sky130_fd_sc_hdll__muxb4to1_2_0/Z VGND
+ VPWR sky130_fd_sc_hdll__muxb4to1_2_0/S[1] sky130_fd_sc_hdll__muxb4to1_2_0/S[2] sky130_fd_sc_hdll__muxb4to1_2_0/S[3]
+ sky130_fd_sc_hdll__muxb4to1_2_0/D[1] sky130_fd_sc_hdll__muxb4to1_2_0/D[0] sky130_fd_sc_hdll__muxb4to1_2_0/D[2]
+ sky130_fd_sc_hdll__muxb4to1_2_0/D[3] sky130_fd_sc_hdll__muxb4to1_2_0/S[0] sky130_fd_sc_hdll__muxb4to1_2
Xsky130_fd_sc_hdll__sdfrbp_1_0 sky130_fd_sc_hdll__sdfrbp_1_0/RESET_B VPWR VGND VGND
+ VPWR sky130_fd_sc_hdll__sdfrbp_1_0/Q_N sky130_fd_sc_hdll__sdfrbp_1_0/D sky130_fd_sc_hdll__sdfrbp_1_0/CLK
+ sky130_fd_sc_hdll__sdfrbp_1_0/Q sky130_fd_sc_hdll__sdfrbp_1_0/SCE sky130_fd_sc_hdll__sdfrbp_1_0/SCD
+ sky130_fd_sc_hdll__sdfrbp_1
Xsky130_fd_sc_hdll__o221a_2_0 sky130_fd_sc_hdll__o221a_2_0/B2 sky130_fd_sc_hdll__o221a_2_0/A2
+ sky130_fd_sc_hdll__o221a_2_0/X sky130_fd_sc_hdll__o221a_2_0/B1 sky130_fd_sc_hdll__o221a_2_0/C1
+ sky130_fd_sc_hdll__o221a_2_0/A1 VPWR VGND VGND VPWR sky130_fd_sc_hdll__o221a_2
Xsky130_fd_sc_hdll__dlxtn_2_0 sky130_fd_sc_hdll__dlxtn_2_0/D sky130_fd_sc_hdll__dlxtn_2_0/GATE_N
+ sky130_fd_sc_hdll__dlxtn_2_0/Q VGND VPWR VPWR VGND sky130_fd_sc_hdll__dlxtn_2
Xsky130_fd_sc_hdll__a22o_2_0 sky130_fd_sc_hdll__a22o_2_0/A1 sky130_fd_sc_hdll__a22o_2_0/A2
+ sky130_fd_sc_hdll__a22o_2_0/X sky130_fd_sc_hdll__a22o_2_0/B2 sky130_fd_sc_hdll__a22o_2_0/B1
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__a22o_2
Xsky130_fd_sc_hdll__nand2_6_0 sky130_fd_sc_hdll__nand2_6_0/Y sky130_fd_sc_hdll__nand2_6_0/A
+ sky130_fd_sc_hdll__nand2_6_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__nand2_6
Xsky130_fd_sc_hdll__o21bai_2_0 sky130_fd_sc_hdll__o21bai_2_0/B1_N sky130_fd_sc_hdll__o21bai_2_0/Y
+ sky130_fd_sc_hdll__o21bai_2_0/A2 sky130_fd_sc_hdll__o21bai_2_0/A1 VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__o21bai_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_294 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_283 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_272 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_261 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_250 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o21a_4_0 sky130_fd_sc_hdll__o21a_4_0/A1 sky130_fd_sc_hdll__o21a_4_0/A2
+ sky130_fd_sc_hdll__o21a_4_0/B1 sky130_fd_sc_hdll__o21a_4_0/X VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__o21a_4
Xsky130_fd_sc_hdll__a21oi_2_0 sky130_fd_sc_hdll__a21oi_2_0/B1 sky130_fd_sc_hdll__a21oi_2_0/A2
+ sky130_fd_sc_hdll__a21oi_2_0/A1 sky130_fd_sc_hdll__a21oi_2_0/Y VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__a21oi_2
Xsky130_fd_sc_hdll__or2_2_0 sky130_fd_sc_hdll__or2_2_0/B sky130_fd_sc_hdll__or2_2_0/X
+ sky130_fd_sc_hdll__or2_2_0/A VPWR VGND VPWR VGND sky130_fd_sc_hdll__or2_2
Xsky130_fd_sc_hdll__decap_12_0 VGND VPWR VPWR VGND sky130_fd_sc_hdll__decap_12
Xsky130_fd_sc_hdll__o211a_2_0 sky130_fd_sc_hdll__o211a_2_0/C1 sky130_fd_sc_hdll__o211a_2_0/B1
+ sky130_fd_sc_hdll__o211a_2_0/A2 sky130_fd_sc_hdll__o211a_2_0/A1 sky130_fd_sc_hdll__o211a_2_0/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__o211a_2
Xsky130_fd_sc_hdll__tapvgnd_1_0 VPWR VGND VPWR sky130_fd_sc_hdll__tapvgnd_1
Xsky130_fd_sc_hdll__nor2_4_0 sky130_fd_sc_hdll__nor2_4_0/Y sky130_fd_sc_hdll__nor2_4_0/A
+ sky130_fd_sc_hdll__nor2_4_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor2_4
Xsky130_fd_sc_hdll__inputiso1p_1_0 sky130_fd_sc_hdll__inputiso1p_1_0/SLEEP sky130_fd_sc_hdll__inputiso1p_1_0/X
+ sky130_fd_sc_hdll__inputiso1p_1_0/A VPWR VGND VGND VPWR sky130_fd_sc_hdll__inputiso1p_1
Xsky130_fd_sc_hdll__dfstp_1_0 sky130_fd_sc_hdll__dfstp_1_0/D VPWR sky130_fd_sc_hdll__dfstp_1_0/CLK
+ VGND sky130_fd_sc_hdll__dfstp_1_0/Q VPWR VGND sky130_fd_sc_hdll__dfstp_1_0/SET_B
+ sky130_fd_sc_hdll__dfstp_1
Xsky130_fd_sc_hdll__nand4b_4_0 sky130_fd_sc_hdll__nand4b_4_0/C sky130_fd_sc_hdll__nand4b_4_0/D
+ sky130_fd_sc_hdll__nand4b_4_0/B sky130_fd_sc_hdll__nand4b_4_0/Y sky130_fd_sc_hdll__nand4b_4_0/A_N
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nand4b_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_295 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_284 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_273 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_262 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_251 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_240 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nand2_12_0 sky130_fd_sc_hdll__nand2_12_0/Y sky130_fd_sc_hdll__nand2_12_0/A
+ sky130_fd_sc_hdll__nand2_12_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__nand2_12
Xsky130_fd_sc_hdll__buf_12_0 sky130_fd_sc_hdll__buf_12_0/A sky130_fd_sc_hdll__buf_12_0/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__buf_12
Xsky130_fd_sc_hdll__a21o_8_0 sky130_fd_sc_hdll__a21o_8_0/A2 sky130_fd_sc_hdll__a21o_8_0/A1
+ sky130_fd_sc_hdll__a21o_8_0/X sky130_fd_sc_hdll__a21o_8_0/B1 VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__a21o_8
Xsky130_fd_sc_hdll__sdfrtn_1_0 VPWR VGND sky130_fd_sc_hdll__sdfrtn_1_0/RESET_B VPWR
+ VGND sky130_fd_sc_hdll__sdfrtn_1_0/SCE sky130_fd_sc_hdll__sdfrtn_1_0/SCD sky130_fd_sc_hdll__sdfrtn_1_0/D
+ sky130_fd_sc_hdll__sdfrtn_1_0/CLK_N sky130_fd_sc_hdll__sdfrtn_1_0/Q sky130_fd_sc_hdll__sdfrtn_1
Xsky130_fd_sc_hdll__o2bb2ai_4_0 sky130_fd_sc_hdll__o2bb2ai_4_0/A1_N sky130_fd_sc_hdll__o2bb2ai_4_0/B1
+ sky130_fd_sc_hdll__o2bb2ai_4_0/B2 sky130_fd_sc_hdll__o2bb2ai_4_0/A2_N sky130_fd_sc_hdll__o2bb2ai_4_0/Y
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__o2bb2ai_4
Xsky130_fd_sc_hdll__nor4_1_0 sky130_fd_sc_hdll__nor4_1_0/D sky130_fd_sc_hdll__nor4_1_0/C
+ sky130_fd_sc_hdll__nor4_1_0/Y sky130_fd_sc_hdll__nor4_1_0/A sky130_fd_sc_hdll__nor4_1_0/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor4_1
Xsky130_fd_sc_hdll__clkinvlp_2_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__clkinvlp_2_0/Y
+ sky130_fd_sc_hdll__clkinvlp_2_0/A sky130_fd_sc_hdll__clkinvlp_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_263 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_252 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_241 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_230 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__einvp_8_0 sky130_fd_sc_hdll__einvp_8_0/A sky130_fd_sc_hdll__einvp_8_0/Z
+ sky130_fd_sc_hdll__einvp_8_0/TE VPWR VGND VPWR VGND sky130_fd_sc_hdll__einvp_8
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_296 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_285 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__and2_4_0 sky130_fd_sc_hdll__and2_4_0/X sky130_fd_sc_hdll__and2_4_0/B
+ sky130_fd_sc_hdll__and2_4_0/A VGND VPWR VGND VPWR sky130_fd_sc_hdll__and2_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_274 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__dfrtp_1_0 sky130_fd_sc_hdll__dfrtp_1_0/RESET_B VGND VPWR sky130_fd_sc_hdll__dfrtp_1_0/Q
+ sky130_fd_sc_hdll__dfrtp_1_0/D sky130_fd_sc_hdll__dfrtp_1_0/CLK VPWR VGND sky130_fd_sc_hdll__dfrtp_1
Xsky130_fd_sc_hdll__sdlclkp_1_0 sky130_fd_sc_hdll__sdlclkp_1_0/CLK VGND VPWR sky130_fd_sc_hdll__sdlclkp_1_0/SCE
+ sky130_fd_sc_hdll__sdlclkp_1_0/GCLK sky130_fd_sc_hdll__sdlclkp_1_0/GATE VPWR VGND
+ sky130_fd_sc_hdll__sdlclkp_1
Xsky130_fd_sc_hdll__a32oi_4_0 sky130_fd_sc_hdll__a32oi_4_0/A3 sky130_fd_sc_hdll__a32oi_4_0/A2
+ sky130_fd_sc_hdll__a32oi_4_0/A1 sky130_fd_sc_hdll__a32oi_4_0/B1 sky130_fd_sc_hdll__a32oi_4_0/Y
+ sky130_fd_sc_hdll__a32oi_4_0/B2 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a32oi_4
Xsky130_fd_sc_hdll__and4_1_0 sky130_fd_sc_hdll__and4_1_0/X sky130_fd_sc_hdll__and4_1_0/C
+ sky130_fd_sc_hdll__and4_1_0/A sky130_fd_sc_hdll__and4_1_0/B sky130_fd_sc_hdll__and4_1_0/D
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__and4_1
Xsky130_fd_sc_hdll__nand2_4_0 sky130_fd_sc_hdll__nand2_4_0/Y sky130_fd_sc_hdll__nand2_4_0/A
+ sky130_fd_sc_hdll__nand2_4_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__nand2_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_297 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_286 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_275 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_264 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_253 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_242 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_231 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_220 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a21bo_4_0 sky130_fd_sc_hdll__a21bo_4_0/B1_N sky130_fd_sc_hdll__a21bo_4_0/A2
+ sky130_fd_sc_hdll__a21bo_4_0/A1 sky130_fd_sc_hdll__a21bo_4_0/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__a21bo_4
Xsky130_fd_sc_hdll__o21a_2_0 sky130_fd_sc_hdll__o21a_2_0/A1 sky130_fd_sc_hdll__o21a_2_0/B1
+ sky130_fd_sc_hdll__o21a_2_0/A2 sky130_fd_sc_hdll__o21a_2_0/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__o21a_2
Xsky130_fd_sc_hdll__a31oi_4_0 sky130_fd_sc_hdll__a31oi_4_0/Y sky130_fd_sc_hdll__a31oi_4_0/B1
+ sky130_fd_sc_hdll__a31oi_4_0/A2 sky130_fd_sc_hdll__a31oi_4_0/A3 sky130_fd_sc_hdll__a31oi_4_0/A1
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__a31oi_4
Xsky130_fd_sc_hdll__mux2i_4_0 sky130_fd_sc_hdll__mux2i_4_0/S sky130_fd_sc_hdll__mux2i_4_0/A1
+ sky130_fd_sc_hdll__mux2i_4_0/A0 sky130_fd_sc_hdll__mux2i_4_0/Y VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__mux2i_4
Xsky130_fd_sc_hdll__nand4_1_0 sky130_fd_sc_hdll__nand4_1_0/C sky130_fd_sc_hdll__nand4_1_0/B
+ sky130_fd_sc_hdll__nand4_1_0/Y sky130_fd_sc_hdll__nand4_1_0/D sky130_fd_sc_hdll__nand4_1_0/A
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__nand4_1
Xsky130_fd_sc_hdll__and3b_1_0 sky130_fd_sc_hdll__and3b_1_0/A_N sky130_fd_sc_hdll__and3b_1_0/B
+ sky130_fd_sc_hdll__and3b_1_0/X sky130_fd_sc_hdll__and3b_1_0/C VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__and3b_1
Xsky130_fd_sc_hdll__ebufn_8_0 sky130_fd_sc_hdll__ebufn_8_0/A sky130_fd_sc_hdll__ebufn_8_0/Z
+ sky130_fd_sc_hdll__ebufn_8_0/TE_B VGND VPWR VGND VPWR sky130_fd_sc_hdll__ebufn_8
Xsky130_fd_sc_hdll__nor2_2_0 sky130_fd_sc_hdll__nor2_2_0/B sky130_fd_sc_hdll__nor2_2_0/Y
+ sky130_fd_sc_hdll__nor2_2_0/A VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor2_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_298 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__dlrtn_4_0 sky130_fd_sc_hdll__dlrtn_4_0/RESET_B sky130_fd_sc_hdll__dlrtn_4_0/D
+ sky130_fd_sc_hdll__dlrtn_4_0/GATE_N sky130_fd_sc_hdll__dlrtn_4_0/Q VGND VPWR VPWR
+ VGND sky130_fd_sc_hdll__dlrtn_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_287 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_276 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_265 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_254 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_243 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_232 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_221 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_210 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nand4b_2_0 sky130_fd_sc_hdll__nand4b_2_0/D sky130_fd_sc_hdll__nand4b_2_0/C
+ sky130_fd_sc_hdll__nand4b_2_0/B sky130_fd_sc_hdll__nand4b_2_0/Y sky130_fd_sc_hdll__nand4b_2_0/A_N
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nand4b_2
Xsky130_fd_sc_hdll__or2b_4_0 sky130_fd_sc_hdll__or2b_4_0/A sky130_fd_sc_hdll__or2b_4_0/B_N
+ sky130_fd_sc_hdll__or2b_4_0/X VGND VPWR VGND VPWR sky130_fd_sc_hdll__or2b_4
Xsky130_fd_sc_hdll__xnor2_1_0 VGND VPWR sky130_fd_sc_hdll__xnor2_1_0/B sky130_fd_sc_hdll__xnor2_1_0/Y
+ sky130_fd_sc_hdll__xnor2_1_0/A VPWR VGND sky130_fd_sc_hdll__xnor2_1
Xsky130_fd_sc_hdll__a21o_6_0 sky130_fd_sc_hdll__a21o_6_0/A2 sky130_fd_sc_hdll__a21o_6_0/A1
+ sky130_fd_sc_hdll__a21o_6_0/X sky130_fd_sc_hdll__a21o_6_0/B1 VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__a21o_6
Xsky130_fd_sc_hdll__a2bb2oi_4_0 sky130_fd_sc_hdll__a2bb2oi_4_0/Y sky130_fd_sc_hdll__a2bb2oi_4_0/A2_N
+ sky130_fd_sc_hdll__a2bb2oi_4_0/B2 sky130_fd_sc_hdll__a2bb2oi_4_0/A1_N sky130_fd_sc_hdll__a2bb2oi_4_0/B1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__a2bb2oi_4
Xsky130_fd_sc_hdll__bufinv_16_0 sky130_fd_sc_hdll__bufinv_16_0/A sky130_fd_sc_hdll__bufinv_16_0/Y
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__bufinv_16
Xsky130_fd_sc_hdll__or4b_1_0 sky130_fd_sc_hdll__or4b_1_0/B sky130_fd_sc_hdll__or4b_1_0/D_N
+ sky130_fd_sc_hdll__or4b_1_0/A sky130_fd_sc_hdll__or4b_1_0/X sky130_fd_sc_hdll__or4b_1_0/C
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__or4b_1
Xsky130_fd_sc_hdll__o2bb2ai_2_0 sky130_fd_sc_hdll__o2bb2ai_2_0/B2 sky130_fd_sc_hdll__o2bb2ai_2_0/Y
+ sky130_fd_sc_hdll__o2bb2ai_2_0/A1_N sky130_fd_sc_hdll__o2bb2ai_2_0/A2_N sky130_fd_sc_hdll__o2bb2ai_2_0/B1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o2bb2ai_2
Xsky130_fd_sc_hdll__a2bb2o_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a2bb2o_1_0/B1
+ sky130_fd_sc_hdll__a2bb2o_1_0/A1_N sky130_fd_sc_hdll__a2bb2o_1_0/A2_N sky130_fd_sc_hdll__a2bb2o_1_0/X
+ sky130_fd_sc_hdll__a2bb2o_1_0/B2 sky130_fd_sc_hdll__a2bb2o_1
Xsky130_fd_sc_hdll__xor3_1_0 sky130_fd_sc_hdll__xor3_1_0/X sky130_fd_sc_hdll__xor3_1_0/C
+ sky130_fd_sc_hdll__xor3_1_0/B sky130_fd_sc_hdll__xor3_1_0/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__xor3_1
Xsky130_fd_sc_hdll__dlrtp_1_0 sky130_fd_sc_hdll__dlrtp_1_0/RESET_B sky130_fd_sc_hdll__dlrtp_1_0/D
+ sky130_fd_sc_hdll__dlrtp_1_0/GATE sky130_fd_sc_hdll__dlrtp_1_0/Q VGND VPWR VPWR
+ VGND sky130_fd_sc_hdll__dlrtp_1
Xsky130_fd_sc_hdll__nor2b_4_0 sky130_fd_sc_hdll__nor2b_4_0/B_N sky130_fd_sc_hdll__nor2b_4_0/Y
+ sky130_fd_sc_hdll__nor2b_4_0/A VGND VPWR VGND VPWR sky130_fd_sc_hdll__nor2b_4
Xsky130_fd_sc_hdll__buf_1_0 VGND VPWR sky130_fd_sc_hdll__buf_1_0/X sky130_fd_sc_hdll__buf_1_0/A
+ VPWR VGND sky130_fd_sc_hdll__buf_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_299 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_288 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_277 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_255 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_244 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_233 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_266 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_222 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__inv_1_0 sky130_fd_sc_hdll__inv_1_0/Y sky130_fd_sc_hdll__inv_1_0/A
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__inv_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_211 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_200 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__and2_2_0 VPWR VGND sky130_fd_sc_hdll__and2_2_0/A sky130_fd_sc_hdll__and2_2_0/X
+ sky130_fd_sc_hdll__and2_2_0/B VPWR VGND sky130_fd_sc_hdll__and2_2
Xsky130_fd_sc_hdll__nor4b_1_0 sky130_fd_sc_hdll__nor4b_1_0/C sky130_fd_sc_hdll__nor4b_1_0/B
+ sky130_fd_sc_hdll__nor4b_1_0/A sky130_fd_sc_hdll__nor4b_1_0/D_N sky130_fd_sc_hdll__nor4b_1_0/Y
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor4b_1
Xsky130_fd_sc_hdll__a211oi_1_0 sky130_fd_sc_hdll__a211oi_1_0/A1 sky130_fd_sc_hdll__a211oi_1_0/C1
+ sky130_fd_sc_hdll__a211oi_1_0/B1 sky130_fd_sc_hdll__a211oi_1_0/Y sky130_fd_sc_hdll__a211oi_1_0/A2
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__a211oi_1
Xsky130_fd_sc_hdll__sedfxbp_2_0 VPWR VGND sky130_fd_sc_hdll__sedfxbp_2_0/CLK sky130_fd_sc_hdll__sedfxbp_2_0/Q_N
+ sky130_fd_sc_hdll__sedfxbp_2_0/SCD sky130_fd_sc_hdll__sedfxbp_2_0/DE sky130_fd_sc_hdll__sedfxbp_2_0/D
+ sky130_fd_sc_hdll__sedfxbp_2_0/Q sky130_fd_sc_hdll__sedfxbp_2_0/SCE VPWR VGND sky130_fd_sc_hdll__sedfxbp_2
Xsky130_fd_sc_hdll__a32oi_2_0 sky130_fd_sc_hdll__a32oi_2_0/A2 sky130_fd_sc_hdll__a32oi_2_0/B2
+ sky130_fd_sc_hdll__a32oi_2_0/A3 sky130_fd_sc_hdll__a32oi_2_0/A1 sky130_fd_sc_hdll__a32oi_2_0/Y
+ sky130_fd_sc_hdll__a32oi_2_0/B1 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a32oi_2
Xsky130_fd_sc_hdll__and4b_4_0 sky130_fd_sc_hdll__and4b_4_0/X sky130_fd_sc_hdll__and4b_4_0/D
+ sky130_fd_sc_hdll__and4b_4_0/C sky130_fd_sc_hdll__and4b_4_0/B sky130_fd_sc_hdll__and4b_4_0/A_N
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__and4b_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_289 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_278 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_267 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_256 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_245 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_234 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_223 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_212 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_201 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nand2_2_0 sky130_fd_sc_hdll__nand2_2_0/Y sky130_fd_sc_hdll__nand2_2_0/A
+ sky130_fd_sc_hdll__nand2_2_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__nand2_2
Xsky130_fd_sc_hdll__a31o_4_0 sky130_fd_sc_hdll__a31o_4_0/B1 sky130_fd_sc_hdll__a31o_4_0/A2
+ sky130_fd_sc_hdll__a31o_4_0/A3 sky130_fd_sc_hdll__a31o_4_0/A1 sky130_fd_sc_hdll__a31o_4_0/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__a31o_4
Xsky130_fd_sc_hdll__xnor3_4_0 sky130_fd_sc_hdll__xnor3_4_0/X sky130_fd_sc_hdll__xnor3_4_0/B
+ sky130_fd_sc_hdll__xnor3_4_0/C sky130_fd_sc_hdll__xnor3_4_0/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__xnor3_4
Xsky130_fd_sc_hdll__a21bo_2_0 sky130_fd_sc_hdll__a21bo_2_0/B1_N sky130_fd_sc_hdll__a21bo_2_0/A2
+ sky130_fd_sc_hdll__a21bo_2_0/X sky130_fd_sc_hdll__a21bo_2_0/A1 VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__a21bo_2
Xsky130_fd_sc_hdll__mux2i_2_0 sky130_fd_sc_hdll__mux2i_2_0/Y sky130_fd_sc_hdll__mux2i_2_0/A1
+ sky130_fd_sc_hdll__mux2i_2_0/A0 sky130_fd_sc_hdll__mux2i_2_0/S VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__mux2i_2
Xsky130_fd_sc_hdll__decap_3_0 VPWR VGND VPWR VGND sky130_fd_sc_hdll__decap_3
Xsky130_fd_sc_hdll__a31oi_2_0 sky130_fd_sc_hdll__a31oi_2_0/A3 sky130_fd_sc_hdll__a31oi_2_0/B1
+ sky130_fd_sc_hdll__a31oi_2_0/Y sky130_fd_sc_hdll__a31oi_2_0/A1 sky130_fd_sc_hdll__a31oi_2_0/A2
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__a31oi_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_279 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_268 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_257 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_246 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_235 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_224 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_213 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_202 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__conb_1_0 sky130_fd_sc_hdll__conb_1_0/LO sky130_fd_sc_hdll__conb_1_0/HI
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__conb_1
Xsky130_fd_sc_hdll__dlrtn_2_0 sky130_fd_sc_hdll__dlrtn_2_0/RESET_B sky130_fd_sc_hdll__dlrtn_2_0/D
+ sky130_fd_sc_hdll__dlrtn_2_0/GATE_N sky130_fd_sc_hdll__dlrtn_2_0/Q VGND VPWR VPWR
+ VGND sky130_fd_sc_hdll__dlrtn_2
Xsky130_fd_sc_hdll__or2b_2_0 sky130_fd_sc_hdll__or2b_2_0/A sky130_fd_sc_hdll__or2b_2_0/B_N
+ sky130_fd_sc_hdll__or2b_2_0/X VPWR VGND VGND VPWR sky130_fd_sc_hdll__or2b_2
Xsky130_fd_sc_hdll__diode_8_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__diode_8_0/DIODE
+ sky130_fd_sc_hdll__diode_8
Xsky130_fd_sc_hdll__sdfxtp_1_0 VPWR VGND sky130_fd_sc_hdll__sdfxtp_1_0/CLK sky130_fd_sc_hdll__sdfxtp_1_0/Q
+ sky130_fd_sc_hdll__sdfxtp_1_0/SCD sky130_fd_sc_hdll__sdfxtp_1_0/D sky130_fd_sc_hdll__sdfxtp_1_0/SCE
+ VPWR VGND sky130_fd_sc_hdll__sdfxtp_1
Xsky130_fd_sc_hdll__a211o_4_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a211o_4_0/C1
+ sky130_fd_sc_hdll__a211o_4_0/B1 sky130_fd_sc_hdll__a211o_4_0/X sky130_fd_sc_hdll__a211o_4_0/A2
+ sky130_fd_sc_hdll__a211o_4_0/A1 sky130_fd_sc_hdll__a211o_4
Xsky130_fd_sc_hdll__a2bb2oi_2_0 sky130_fd_sc_hdll__a2bb2oi_2_0/A2_N sky130_fd_sc_hdll__a2bb2oi_2_0/A1_N
+ sky130_fd_sc_hdll__a2bb2oi_2_0/Y sky130_fd_sc_hdll__a2bb2oi_2_0/B2 sky130_fd_sc_hdll__a2bb2oi_2_0/B1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__a2bb2oi_2
Xsky130_fd_sc_hdll__a21o_4_0 sky130_fd_sc_hdll__a21o_4_0/A2 sky130_fd_sc_hdll__a21o_4_0/A1
+ sky130_fd_sc_hdll__a21o_4_0/X sky130_fd_sc_hdll__a21o_4_0/B1 VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__a21o_4
Xsky130_fd_sc_hdll__dlygate4sd1_1_0 sky130_fd_sc_hdll__dlygate4sd1_1_0/A sky130_fd_sc_hdll__dlygate4sd1_1_0/X
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__dlygate4sd1_1
Xsky130_fd_sc_hdll__sdfxbp_2_0 VPWR VGND sky130_fd_sc_hdll__sdfxbp_2_0/Q_N sky130_fd_sc_hdll__sdfxbp_2_0/Q
+ sky130_fd_sc_hdll__sdfxbp_2_0/CLK sky130_fd_sc_hdll__sdfxbp_2_0/SCE sky130_fd_sc_hdll__sdfxbp_2_0/D
+ sky130_fd_sc_hdll__sdfxbp_2_0/SCD VGND VPWR sky130_fd_sc_hdll__sdfxbp_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_269 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_258 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_247 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_236 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_225 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_214 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_203 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nor2b_2_0 sky130_fd_sc_hdll__nor2b_2_0/B_N sky130_fd_sc_hdll__nor2b_2_0/A
+ sky130_fd_sc_hdll__nor2b_2_0/Y VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor2b_2
Xsky130_fd_sc_hdll__nor4_8_0 sky130_fd_sc_hdll__nor4_8_0/A sky130_fd_sc_hdll__nor4_8_0/C
+ sky130_fd_sc_hdll__nor4_8_0/D sky130_fd_sc_hdll__nor4_8_0/B sky130_fd_sc_hdll__nor4_8_0/Y
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor4_8
Xsky130_fd_sc_hdll__einvp_4_0 sky130_fd_sc_hdll__einvp_4_0/TE sky130_fd_sc_hdll__einvp_4_0/A
+ sky130_fd_sc_hdll__einvp_4_0/Z VPWR VGND VPWR VGND sky130_fd_sc_hdll__einvp_4
Xsky130_fd_sc_hdll__muxb8to1_1_0 VGND sky130_fd_sc_hdll__muxb8to1_1_0/Z VPWR VGND
+ VPWR sky130_fd_sc_hdll__muxb8to1_1_0/D[0] sky130_fd_sc_hdll__muxb8to1_1_0/S[0] sky130_fd_sc_hdll__muxb8to1_1_0/S[1]
+ sky130_fd_sc_hdll__muxb8to1_1_0/D[1] sky130_fd_sc_hdll__muxb8to1_1_0/D[2] sky130_fd_sc_hdll__muxb8to1_1_0/S[2]
+ sky130_fd_sc_hdll__muxb8to1_1_0/S[3] sky130_fd_sc_hdll__muxb8to1_1_0/D[4] sky130_fd_sc_hdll__muxb8to1_1_0/S[4]
+ sky130_fd_sc_hdll__muxb8to1_1_0/S[5] sky130_fd_sc_hdll__muxb8to1_1_0/D[5] sky130_fd_sc_hdll__muxb8to1_1_0/D[6]
+ sky130_fd_sc_hdll__muxb8to1_1_0/S[6] sky130_fd_sc_hdll__muxb8to1_1_0/S[7] sky130_fd_sc_hdll__muxb8to1_1_0/D[7]
+ sky130_fd_sc_hdll__muxb8to1_1_0/D[3] sky130_fd_sc_hdll__muxb8to1_1
Xsky130_fd_sc_hdll__o2bb2a_1_0 sky130_fd_sc_hdll__o2bb2a_1_0/A1_N sky130_fd_sc_hdll__o2bb2a_1_0/X
+ sky130_fd_sc_hdll__o2bb2a_1_0/A2_N sky130_fd_sc_hdll__o2bb2a_1_0/B2 sky130_fd_sc_hdll__o2bb2a_1_0/B1
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__o2bb2a_1
Xsky130_fd_sc_hdll__or3_1_0 sky130_fd_sc_hdll__or3_1_0/A sky130_fd_sc_hdll__or3_1_0/X
+ sky130_fd_sc_hdll__or3_1_0/B sky130_fd_sc_hdll__or3_1_0/C VPWR VGND VPWR VGND sky130_fd_sc_hdll__or3_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_259 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_248 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_237 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_226 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_215 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_204 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__and4b_2_0 VPWR VGND sky130_fd_sc_hdll__and4b_2_0/X sky130_fd_sc_hdll__and4b_2_0/A_N
+ sky130_fd_sc_hdll__and4b_2_0/D sky130_fd_sc_hdll__and4b_2_0/C sky130_fd_sc_hdll__and4b_2_0/B
+ VGND VPWR sky130_fd_sc_hdll__and4b_2
Xsky130_fd_sc_hdll__o22ai_1_0 sky130_fd_sc_hdll__o22ai_1_0/B2 sky130_fd_sc_hdll__o22ai_1_0/A1
+ sky130_fd_sc_hdll__o22ai_1_0/Y sky130_fd_sc_hdll__o22ai_1_0/B1 sky130_fd_sc_hdll__o22ai_1_0/A2
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__o22ai_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_90 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a31o_2_0 sky130_fd_sc_hdll__a31o_2_0/X sky130_fd_sc_hdll__a31o_2_0/B1
+ sky130_fd_sc_hdll__a31o_2_0/A3 sky130_fd_sc_hdll__a31o_2_0/A1 sky130_fd_sc_hdll__a31o_2_0/A2
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__a31o_2
Xsky130_fd_sc_hdll__xnor3_2_0 sky130_fd_sc_hdll__xnor3_2_0/X sky130_fd_sc_hdll__xnor3_2_0/B
+ sky130_fd_sc_hdll__xnor3_2_0/C sky130_fd_sc_hdll__xnor3_2_0/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__xnor3_2
Xsky130_fd_sc_hdll__nand2b_1_0 sky130_fd_sc_hdll__nand2b_1_0/Y sky130_fd_sc_hdll__nand2b_1_0/A_N
+ sky130_fd_sc_hdll__nand2b_1_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__nand2b_1
Xsky130_fd_sc_hdll__nand4bb_4_0 sky130_fd_sc_hdll__nand4bb_4_0/B_N sky130_fd_sc_hdll__nand4bb_4_0/A_N
+ sky130_fd_sc_hdll__nand4bb_4_0/C sky130_fd_sc_hdll__nand4bb_4_0/Y sky130_fd_sc_hdll__nand4bb_4_0/D
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nand4bb_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_249 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_238 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_227 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_216 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_205 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o211ai_1_0 sky130_fd_sc_hdll__o211ai_1_0/A1 sky130_fd_sc_hdll__o211ai_1_0/A2
+ sky130_fd_sc_hdll__o211ai_1_0/Y sky130_fd_sc_hdll__o211ai_1_0/C1 sky130_fd_sc_hdll__o211ai_1_0/B1
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__o211ai_1
Xsky130_fd_sc_hdll__muxb16to1_4_0 VGND sky130_fd_sc_hdll__muxb16to1_4_0/Z VPWR VGND
+ VPWR sky130_fd_sc_hdll__muxb16to1_4_0/S[6] sky130_fd_sc_hdll__muxb16to1_4_0/S[10]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[12] sky130_fd_sc_hdll__muxb16to1_4_0/D[13] sky130_fd_sc_hdll__muxb16to1_4_0/D[8]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[15] sky130_fd_sc_hdll__muxb16to1_4_0/D[10] sky130_fd_sc_hdll__muxb16to1_4_0/D[9]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[14] sky130_fd_sc_hdll__muxb16to1_4_0/S[14] sky130_fd_sc_hdll__muxb16to1_4_0/D[11]
+ sky130_fd_sc_hdll__muxb16to1_4_0/S[11] sky130_fd_sc_hdll__muxb16to1_4_0/S[8] sky130_fd_sc_hdll__muxb16to1_4_0/S[15]
+ sky130_fd_sc_hdll__muxb16to1_4_0/S[12] sky130_fd_sc_hdll__muxb16to1_4_0/S[9] sky130_fd_sc_hdll__muxb16to1_4_0/S[13]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[3] sky130_fd_sc_hdll__muxb16to1_4_0/D[0] sky130_fd_sc_hdll__muxb16to1_4_0/D[4]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[5] sky130_fd_sc_hdll__muxb16to1_4_0/D[2] sky130_fd_sc_hdll__muxb16to1_4_0/D[1]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[6] sky130_fd_sc_hdll__muxb16to1_4_0/S[2] sky130_fd_sc_hdll__muxb16to1_4_0/S[3]
+ sky130_fd_sc_hdll__muxb16to1_4_0/S[7] sky130_fd_sc_hdll__muxb16to1_4_0/S[0] sky130_fd_sc_hdll__muxb16to1_4_0/S[1]
+ sky130_fd_sc_hdll__muxb16to1_4_0/S[4] sky130_fd_sc_hdll__muxb16to1_4_0/S[5] sky130_fd_sc_hdll__muxb16to1_4_0/D[7]
+ sky130_fd_sc_hdll__muxb16to1_4
Xsky130_fd_sc_hdll__ebufn_4_0 sky130_fd_sc_hdll__ebufn_4_0/A sky130_fd_sc_hdll__ebufn_4_0/Z
+ sky130_fd_sc_hdll__ebufn_4_0/TE_B VGND VPWR VGND VPWR sky130_fd_sc_hdll__ebufn_4
Xsky130_fd_sc_hdll__clkmux2_1_0 VGND VPWR sky130_fd_sc_hdll__clkmux2_1_0/S sky130_fd_sc_hdll__clkmux2_1_0/A1
+ sky130_fd_sc_hdll__clkmux2_1_0/A0 sky130_fd_sc_hdll__clkmux2_1_0/X VPWR VGND sky130_fd_sc_hdll__clkmux2_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_80 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_91 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o21ai_1_0 VGND VPWR sky130_fd_sc_hdll__o21ai_1_0/A2 sky130_fd_sc_hdll__o21ai_1_0/A1
+ sky130_fd_sc_hdll__o21ai_1_0/B1 sky130_fd_sc_hdll__o21ai_1_0/Y VPWR VGND sky130_fd_sc_hdll__o21ai_1
Xsky130_fd_sc_hdll__a222oi_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a222oi_1_0/C2
+ sky130_fd_sc_hdll__a222oi_1_0/C1 sky130_fd_sc_hdll__a222oi_1_0/B1 sky130_fd_sc_hdll__a222oi_1_0/A2
+ sky130_fd_sc_hdll__a222oi_1_0/A1 sky130_fd_sc_hdll__a222oi_1_0/Y sky130_fd_sc_hdll__a222oi_1_0/B2
+ sky130_fd_sc_hdll__a222oi_1
Xsky130_fd_sc_hdll__diode_6_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__diode_6_0/DIODE
+ sky130_fd_sc_hdll__diode_6
Xsky130_fd_sc_hdll__clkinv_16_0 sky130_fd_sc_hdll__clkinv_16_0/Y sky130_fd_sc_hdll__clkinv_16_0/A
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__clkinv_16
Xsky130_fd_sc_hdll__a21o_2_0 sky130_fd_sc_hdll__a21o_2_0/X sky130_fd_sc_hdll__a21o_2_0/B1
+ sky130_fd_sc_hdll__a21o_2_0/A1 sky130_fd_sc_hdll__a21o_2_0/A2 VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__a21o_2
Xsky130_fd_sc_hdll__a211o_2_0 sky130_fd_sc_hdll__a211o_2_0/X sky130_fd_sc_hdll__a211o_2_0/A2
+ sky130_fd_sc_hdll__a211o_2_0/A1 sky130_fd_sc_hdll__a211o_2_0/B1 sky130_fd_sc_hdll__a211o_2_0/C1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__a211o_2
Xsky130_fd_sc_hdll__nor4bb_1_0 sky130_fd_sc_hdll__nor4bb_1_0/A sky130_fd_sc_hdll__nor4bb_1_0/C_N
+ sky130_fd_sc_hdll__nor4bb_1_0/D_N sky130_fd_sc_hdll__nor4bb_1_0/B sky130_fd_sc_hdll__nor4bb_1_0/Y
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nor4bb_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_239 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_228 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_217 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_206 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__isobufsrc_1_0 sky130_fd_sc_hdll__isobufsrc_1_0/A sky130_fd_sc_hdll__isobufsrc_1_0/X
+ sky130_fd_sc_hdll__isobufsrc_1_0/SLEEP VPWR VGND VGND VPWR sky130_fd_sc_hdll__isobufsrc_1
Xsky130_fd_sc_hdll__or4_4_0 sky130_fd_sc_hdll__or4_4_0/B sky130_fd_sc_hdll__or4_4_0/C
+ sky130_fd_sc_hdll__or4_4_0/A sky130_fd_sc_hdll__or4_4_0/D sky130_fd_sc_hdll__or4_4_0/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__or4_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_70 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_81 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_92 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nor4_6_0 sky130_fd_sc_hdll__nor4_6_0/A sky130_fd_sc_hdll__nor4_6_0/C
+ sky130_fd_sc_hdll__nor4_6_0/D sky130_fd_sc_hdll__nor4_6_0/B sky130_fd_sc_hdll__nor4_6_0/Y
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor4_6
Xsky130_fd_sc_hdll__and4bb_4_0 sky130_fd_sc_hdll__and4bb_4_0/C sky130_fd_sc_hdll__and4bb_4_0/A_N
+ sky130_fd_sc_hdll__and4bb_4_0/D sky130_fd_sc_hdll__and4bb_4_0/X sky130_fd_sc_hdll__and4bb_4_0/B_N
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__and4bb_4
Xsky130_fd_sc_hdll__einvp_2_0 sky130_fd_sc_hdll__einvp_2_0/A sky130_fd_sc_hdll__einvp_2_0/Z
+ sky130_fd_sc_hdll__einvp_2_0/TE VGND VPWR VPWR VGND sky130_fd_sc_hdll__einvp_2
Xsky130_fd_sc_hdll__a221oi_1_0 sky130_fd_sc_hdll__a221oi_1_0/Y sky130_fd_sc_hdll__a221oi_1_0/C1
+ sky130_fd_sc_hdll__a221oi_1_0/A1 sky130_fd_sc_hdll__a221oi_1_0/A2 sky130_fd_sc_hdll__a221oi_1_0/B2
+ sky130_fd_sc_hdll__a221oi_1_0/B1 VGND VPWR VPWR VGND sky130_fd_sc_hdll__a221oi_1
Xsky130_fd_sc_hdll__buf_8_0 sky130_fd_sc_hdll__buf_8_0/A sky130_fd_sc_hdll__buf_8_0/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__buf_8
Xsky130_fd_sc_hdll__inv_8_0 sky130_fd_sc_hdll__inv_8_0/A sky130_fd_sc_hdll__inv_8_0/Y
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__inv_8
Xsky130_fd_sc_hdll__o22a_1_0 sky130_fd_sc_hdll__o22a_1_0/A2 sky130_fd_sc_hdll__o22a_1_0/X
+ sky130_fd_sc_hdll__o22a_1_0/B1 sky130_fd_sc_hdll__o22a_1_0/A1 sky130_fd_sc_hdll__o22a_1_0/B2
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__o22a_1
Xsky130_fd_sc_hdll__inputiso0p_1_0 sky130_fd_sc_hdll__inputiso0p_1_0/X sky130_fd_sc_hdll__inputiso0p_1_0/SLEEP
+ sky130_fd_sc_hdll__inputiso0p_1_0/A VGND VPWR VPWR VGND sky130_fd_sc_hdll__inputiso0p_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_229 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_218 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_207 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nand3b_4_0 sky130_fd_sc_hdll__nand3b_4_0/A_N sky130_fd_sc_hdll__nand3b_4_0/Y
+ sky130_fd_sc_hdll__nand3b_4_0/B sky130_fd_sc_hdll__nand3b_4_0/C VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__nand3b_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_60 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_71 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_82 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_93 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nor3_1_0 sky130_fd_sc_hdll__nor3_1_0/C sky130_fd_sc_hdll__nor3_1_0/Y
+ sky130_fd_sc_hdll__nor3_1_0/A sky130_fd_sc_hdll__nor3_1_0/B VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__nor3_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_219 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_208 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nand4bb_2_0 sky130_fd_sc_hdll__nand4bb_2_0/D sky130_fd_sc_hdll__nand4bb_2_0/C
+ sky130_fd_sc_hdll__nand4bb_2_0/B_N sky130_fd_sc_hdll__nand4bb_2_0/A_N sky130_fd_sc_hdll__nand4bb_2_0/Y
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nand4bb_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_50 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_61 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_72 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_83 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_94 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__muxb16to1_2_0 sky130_fd_sc_hdll__muxb16to1_2_0/Z VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__muxb16to1_2_0/D[2] sky130_fd_sc_hdll__muxb16to1_2_0/D[1]
+ sky130_fd_sc_hdll__muxb16to1_2_0/S[7] sky130_fd_sc_hdll__muxb16to1_2_0/S[6] sky130_fd_sc_hdll__muxb16to1_2_0/S[5]
+ sky130_fd_sc_hdll__muxb16to1_2_0/D[9] sky130_fd_sc_hdll__muxb16to1_2_0/D[8] sky130_fd_sc_hdll__muxb16to1_2_0/S[14]
+ sky130_fd_sc_hdll__muxb16to1_2_0/S[13] sky130_fd_sc_hdll__muxb16to1_2_0/S[12] sky130_fd_sc_hdll__muxb16to1_2_0/S[11]
+ sky130_fd_sc_hdll__muxb16to1_2_0/S[10] sky130_fd_sc_hdll__muxb16to1_2_0/S[9] sky130_fd_sc_hdll__muxb16to1_2_0/S[8]
+ sky130_fd_sc_hdll__muxb16to1_2_0/D[15] sky130_fd_sc_hdll__muxb16to1_2_0/D[14] sky130_fd_sc_hdll__muxb16to1_2_0/D[13]
+ sky130_fd_sc_hdll__muxb16to1_2_0/D[12] sky130_fd_sc_hdll__muxb16to1_2_0/D[11] sky130_fd_sc_hdll__muxb16to1_2_0/D[10]
+ sky130_fd_sc_hdll__muxb16to1_2_0/S[15] sky130_fd_sc_hdll__muxb16to1_2_0/S[4] sky130_fd_sc_hdll__muxb16to1_2_0/S[3]
+ sky130_fd_sc_hdll__muxb16to1_2_0/S[2] sky130_fd_sc_hdll__muxb16to1_2_0/S[1] sky130_fd_sc_hdll__muxb16to1_2_0/S[0]
+ sky130_fd_sc_hdll__muxb16to1_2_0/D[7] sky130_fd_sc_hdll__muxb16to1_2_0/D[6] sky130_fd_sc_hdll__muxb16to1_2_0/D[5]
+ sky130_fd_sc_hdll__muxb16to1_2_0/D[4] sky130_fd_sc_hdll__muxb16to1_2_0/D[3] sky130_fd_sc_hdll__muxb16to1_2_0/D[0]
+ sky130_fd_sc_hdll__muxb16to1_2
Xsky130_fd_sc_hdll__ebufn_2_0 sky130_fd_sc_hdll__ebufn_2_0/Z sky130_fd_sc_hdll__ebufn_2_0/A
+ sky130_fd_sc_hdll__ebufn_2_0/TE_B VGND VPWR VGND VPWR sky130_fd_sc_hdll__ebufn_2
Xsky130_fd_sc_hdll__diode_4_0 sky130_fd_sc_hdll__diode_4_0/DIODE VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__diode_4
Xsky130_fd_sc_hdll__and3_1_0 VGND VPWR sky130_fd_sc_hdll__and3_1_0/X sky130_fd_sc_hdll__and3_1_0/B
+ sky130_fd_sc_hdll__and3_1_0/A sky130_fd_sc_hdll__and3_1_0/C VPWR VGND sky130_fd_sc_hdll__and3_1
Xsky130_fd_sc_hdll__clkbuf_1_0 VGND VPWR sky130_fd_sc_hdll__clkbuf_1_0/X sky130_fd_sc_hdll__clkbuf_1_0/A
+ VPWR sky130_fd_sc_hdll__clkbuf_1_0/VNB VGND sky130_fd_sc_hdll__clkbuf_1
Xsky130_fd_sc_hdll__clkinv_1_0 sky130_fd_sc_hdll__clkinv_1_0/Y sky130_fd_sc_hdll__clkinv_1_0/A
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__clkinv_1
Xsky130_fd_sc_hdll__sdfstp_1_0 sky130_fd_sc_hdll__sdfstp_1_0/SCE sky130_fd_sc_hdll__sdfstp_1_0/SET_B
+ VPWR VGND sky130_fd_sc_hdll__sdfstp_1_0/CLK sky130_fd_sc_hdll__sdfstp_1_0/D sky130_fd_sc_hdll__sdfstp_1_0/SCD
+ sky130_fd_sc_hdll__sdfstp_1_0/Q VPWR VGND sky130_fd_sc_hdll__sdfstp_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_209 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__dfstp_4_0 sky130_fd_sc_hdll__dfstp_4_0/Q sky130_fd_sc_hdll__dfstp_4_0/D
+ VPWR sky130_fd_sc_hdll__dfstp_4_0/CLK VGND VPWR VGND sky130_fd_sc_hdll__dfstp_4_0/SET_B
+ sky130_fd_sc_hdll__dfstp_4
Xsky130_fd_sc_hdll__or4_2_0 sky130_fd_sc_hdll__or4_2_0/B sky130_fd_sc_hdll__or4_2_0/C
+ sky130_fd_sc_hdll__or4_2_0/A sky130_fd_sc_hdll__or4_2_0/X sky130_fd_sc_hdll__or4_2_0/D
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__or4_2
Xsky130_fd_sc_hdll__sdfsbp_2_0 sky130_fd_sc_hdll__sdfsbp_2_0/Q_N sky130_fd_sc_hdll__sdfsbp_2_0/Q
+ sky130_fd_sc_hdll__sdfsbp_2_0/CLK sky130_fd_sc_hdll__sdfsbp_2_0/D sky130_fd_sc_hdll__sdfsbp_2_0/SCD
+ sky130_fd_sc_hdll__sdfsbp_2_0/SCE sky130_fd_sc_hdll__sdfsbp_2_0/SET_B VGND VPWR
+ VPWR VGND sky130_fd_sc_hdll__sdfsbp_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_40 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_51 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_62 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_73 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_84 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_95 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a21boi_1_0 sky130_fd_sc_hdll__a21boi_1_0/Y sky130_fd_sc_hdll__a21boi_1_0/A1
+ sky130_fd_sc_hdll__a21boi_1_0/B1_N sky130_fd_sc_hdll__a21boi_1_0/A2 VPWR VGND VPWR
+ VGND sky130_fd_sc_hdll__a21boi_1
Xsky130_fd_sc_hdll__and4bb_2_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__and4bb_2_0/A_N
+ sky130_fd_sc_hdll__and4bb_2_0/C sky130_fd_sc_hdll__and4bb_2_0/B_N sky130_fd_sc_hdll__and4bb_2_0/X
+ sky130_fd_sc_hdll__and4bb_2_0/D sky130_fd_sc_hdll__and4bb_2
Xsky130_fd_sc_hdll__nand3_1_0 sky130_fd_sc_hdll__nand3_1_0/Y sky130_fd_sc_hdll__nand3_1_0/A
+ sky130_fd_sc_hdll__nand3_1_0/C sky130_fd_sc_hdll__nand3_1_0/B VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__nand3_1
Xsky130_fd_sc_hdll__nor4_4_0 sky130_fd_sc_hdll__nor4_4_0/A sky130_fd_sc_hdll__nor4_4_0/C
+ sky130_fd_sc_hdll__nor4_4_0/Y sky130_fd_sc_hdll__nor4_4_0/D sky130_fd_sc_hdll__nor4_4_0/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor4_4
Xsky130_fd_sc_hdll__mux2_1_0 VGND VPWR sky130_fd_sc_hdll__mux2_1_0/S sky130_fd_sc_hdll__mux2_1_0/A1
+ sky130_fd_sc_hdll__mux2_1_0/A0 sky130_fd_sc_hdll__mux2_1_0/X VPWR VGND sky130_fd_sc_hdll__mux2_1
Xsky130_fd_sc_hdll__and2b_1_0 sky130_fd_sc_hdll__and2b_1_0/X sky130_fd_sc_hdll__and2b_1_0/A_N
+ sky130_fd_sc_hdll__and2b_1_0/B VGND VPWR VPWR VGND sky130_fd_sc_hdll__and2b_1
Xsky130_fd_sc_hdll__buf_6_0 VPWR VGND sky130_fd_sc_hdll__buf_6_0/X sky130_fd_sc_hdll__buf_6_0/A
+ VPWR VGND sky130_fd_sc_hdll__buf_6
Xsky130_fd_sc_hdll__inv_16_0 sky130_fd_sc_hdll__inv_16_0/Y sky130_fd_sc_hdll__inv_16_0/A
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__inv_16
Xsky130_fd_sc_hdll__inv_6_0 sky130_fd_sc_hdll__inv_6_0/Y sky130_fd_sc_hdll__inv_6_0/A
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__inv_6
Xsky130_fd_sc_hdll__tapvgnd2_1_0 VPWR VGND VPWR sky130_fd_sc_hdll__tapvgnd2_1
Xsky130_fd_sc_hdll__nand3b_2_0 sky130_fd_sc_hdll__nand3b_2_0/Y sky130_fd_sc_hdll__nand3b_2_0/C
+ sky130_fd_sc_hdll__nand3b_2_0/A_N sky130_fd_sc_hdll__nand3b_2_0/B VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__nand3b_2
Xsky130_fd_sc_hdll__sdfrtp_1_0 VPWR VGND VGND VPWR sky130_fd_sc_hdll__sdfrtp_1_0/RESET_B
+ sky130_fd_sc_hdll__sdfrtp_1_0/Q sky130_fd_sc_hdll__sdfrtp_1_0/CLK sky130_fd_sc_hdll__sdfrtp_1_0/D
+ sky130_fd_sc_hdll__sdfrtp_1_0/SCD sky130_fd_sc_hdll__sdfrtp_1_0/SCE sky130_fd_sc_hdll__sdfrtp_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_30 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_41 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_52 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_63 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_74 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_85 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_96 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__dfrtp_4_0 sky130_fd_sc_hdll__dfrtp_4_0/Q sky130_fd_sc_hdll__dfrtp_4_0/D
+ sky130_fd_sc_hdll__dfrtp_4_0/CLK VGND VPWR sky130_fd_sc_hdll__dfrtp_4_0/RESET_B
+ VPWR VGND sky130_fd_sc_hdll__dfrtp_4
Xsky130_fd_sc_hdll__isobufsrc_16_0 sky130_fd_sc_hdll__isobufsrc_16_0/A sky130_fd_sc_hdll__isobufsrc_16_0/X
+ sky130_fd_sc_hdll__isobufsrc_16_0/SLEEP VPWR VGND VGND VPWR sky130_fd_sc_hdll__isobufsrc_16
Xsky130_fd_sc_hdll__sdlclkp_4_0 sky130_fd_sc_hdll__sdlclkp_4_0/SCE sky130_fd_sc_hdll__sdlclkp_4_0/GATE
+ sky130_fd_sc_hdll__sdlclkp_4_0/GCLK VGND VPWR sky130_fd_sc_hdll__sdlclkp_4_0/CLK
+ VPWR VGND sky130_fd_sc_hdll__sdlclkp_4
Xsky130_fd_sc_hdll__sdfrbp_2_0 VPWR VGND VPWR VGND sky130_fd_sc_hdll__sdfrbp_2_0/RESET_B
+ sky130_fd_sc_hdll__sdfrbp_2_0/Q_N sky130_fd_sc_hdll__sdfrbp_2_0/Q sky130_fd_sc_hdll__sdfrbp_2_0/SCD
+ sky130_fd_sc_hdll__sdfrbp_2_0/SCE sky130_fd_sc_hdll__sdfrbp_2_0/CLK sky130_fd_sc_hdll__sdfrbp_2_0/D
+ sky130_fd_sc_hdll__sdfrbp_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_190 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__or3b_1_0 sky130_fd_sc_hdll__or3b_1_0/A sky130_fd_sc_hdll__or3b_1_0/C_N
+ sky130_fd_sc_hdll__or3b_1_0/X sky130_fd_sc_hdll__or3b_1_0/B VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__or3b_1
Xsky130_fd_sc_hdll__o32ai_1_0 sky130_fd_sc_hdll__o32ai_1_0/A2 sky130_fd_sc_hdll__o32ai_1_0/Y
+ sky130_fd_sc_hdll__o32ai_1_0/A1 sky130_fd_sc_hdll__o32ai_1_0/A3 sky130_fd_sc_hdll__o32ai_1_0/B2
+ sky130_fd_sc_hdll__o32ai_1_0/B1 VPWR VGND VGND VPWR sky130_fd_sc_hdll__o32ai_1
Xsky130_fd_sc_hdll__xor2_1_0 sky130_fd_sc_hdll__xor2_1_0/B sky130_fd_sc_hdll__xor2_1_0/X
+ sky130_fd_sc_hdll__xor2_1_0/A VGND VPWR VPWR VGND sky130_fd_sc_hdll__xor2_1
Xsky130_fd_sc_hdll__o21ba_1_0 sky130_fd_sc_hdll__o21ba_1_0/B1_N sky130_fd_sc_hdll__o21ba_1_0/A1
+ sky130_fd_sc_hdll__o21ba_1_0/X sky130_fd_sc_hdll__o21ba_1_0/A2 VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__o21ba_1
Xsky130_fd_sc_hdll__or4bb_1_0 sky130_fd_sc_hdll__or4bb_1_0/A sky130_fd_sc_hdll__or4bb_1_0/X
+ sky130_fd_sc_hdll__or4bb_1_0/B sky130_fd_sc_hdll__or4bb_1_0/D_N sky130_fd_sc_hdll__or4bb_1_0/C_N
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__or4bb_1
Xsky130_fd_sc_hdll__and4_4_0 sky130_fd_sc_hdll__and4_4_0/X sky130_fd_sc_hdll__and4_4_0/C
+ sky130_fd_sc_hdll__and4_4_0/A sky130_fd_sc_hdll__and4_4_0/B sky130_fd_sc_hdll__and4_4_0/D
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__and4_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_31 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_42 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_53 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_64 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_75 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_86 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_97 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_20 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o221ai_1_0 sky130_fd_sc_hdll__o221ai_1_0/A2 sky130_fd_sc_hdll__o221ai_1_0/Y
+ sky130_fd_sc_hdll__o221ai_1_0/B1 sky130_fd_sc_hdll__o221ai_1_0/C1 sky130_fd_sc_hdll__o221ai_1_0/A1
+ sky130_fd_sc_hdll__o221ai_1_0/B2 VPWR VGND VGND VPWR sky130_fd_sc_hdll__o221ai_1
Xsky130_fd_sc_hdll__nor3b_1_0 sky130_fd_sc_hdll__nor3b_1_0/C_N sky130_fd_sc_hdll__nor3b_1_0/Y
+ sky130_fd_sc_hdll__nor3b_1_0/A sky130_fd_sc_hdll__nor3b_1_0/B VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__nor3b_1
Xsky130_fd_sc_hdll__mux2_16_0 VPWR VGND VPWR VGND sky130_fd_sc_hdll__mux2_16_0/X sky130_fd_sc_hdll__mux2_16_0/S
+ sky130_fd_sc_hdll__mux2_16_0/A1 sky130_fd_sc_hdll__mux2_16_0/A0 sky130_fd_sc_hdll__mux2_16
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_191 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_180 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nand4_4_0 sky130_fd_sc_hdll__nand4_4_0/A sky130_fd_sc_hdll__nand4_4_0/D
+ sky130_fd_sc_hdll__nand4_4_0/C sky130_fd_sc_hdll__nand4_4_0/B sky130_fd_sc_hdll__nand4_4_0/Y
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__nand4_4
Xsky130_fd_sc_hdll__decap_8_0 VPWR VGND VPWR VGND sky130_fd_sc_hdll__decap_8
Xsky130_fd_sc_hdll__diode_2_0 sky130_fd_sc_hdll__diode_2_0/DIODE VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__diode_2
Xsky130_fd_sc_hdll__o31ai_1_0 sky130_fd_sc_hdll__o31ai_1_0/Y sky130_fd_sc_hdll__o31ai_1_0/A2
+ sky130_fd_sc_hdll__o31ai_1_0/A1 sky130_fd_sc_hdll__o31ai_1_0/A3 sky130_fd_sc_hdll__o31ai_1_0/B1
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__o31ai_1
Xsky130_fd_sc_hdll__clkinv_12_0 sky130_fd_sc_hdll__clkinv_12_0/Y sky130_fd_sc_hdll__clkinv_12_0/A
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__clkinv_12
Xsky130_fd_sc_hdll__and3b_4_0 sky130_fd_sc_hdll__and3b_4_0/A_N sky130_fd_sc_hdll__and3b_4_0/X
+ sky130_fd_sc_hdll__and3b_4_0/C sky130_fd_sc_hdll__and3b_4_0/B VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__and3b_4
Xsky130_fd_sc_hdll__einvn_1_0 sky130_fd_sc_hdll__einvn_1_0/Z sky130_fd_sc_hdll__einvn_1_0/A
+ sky130_fd_sc_hdll__einvn_1_0/TE_B VGND VPWR VPWR VGND sky130_fd_sc_hdll__einvn_1
Xsky130_fd_sc_hdll__dfstp_2_0 sky130_fd_sc_hdll__dfstp_2_0/Q VGND sky130_fd_sc_hdll__dfstp_2_0/CLK
+ VPWR sky130_fd_sc_hdll__dfstp_2_0/D VPWR VGND sky130_fd_sc_hdll__dfstp_2_0/SET_B
+ sky130_fd_sc_hdll__dfstp_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_32 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_43 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_54 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_65 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_76 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_87 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_98 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_10 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_21 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__xnor2_4_0 sky130_fd_sc_hdll__xnor2_4_0/Y sky130_fd_sc_hdll__xnor2_4_0/B
+ sky130_fd_sc_hdll__xnor2_4_0/A VGND VPWR VGND VPWR sky130_fd_sc_hdll__xnor2_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_192 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_181 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_170 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__fill_1_0 VPWR VGND VPWR VGND sky130_fd_sc_hdll__fill_1
Xsky130_fd_sc_hdll__or4b_4_0 sky130_fd_sc_hdll__or4b_4_0/D_N sky130_fd_sc_hdll__or4b_4_0/B
+ sky130_fd_sc_hdll__or4b_4_0/C sky130_fd_sc_hdll__or4b_4_0/A sky130_fd_sc_hdll__or4b_4_0/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__or4b_4
Xsky130_fd_sc_hdll__a2bb2o_4_0 sky130_fd_sc_hdll__a2bb2o_4_0/X sky130_fd_sc_hdll__a2bb2o_4_0/B1
+ sky130_fd_sc_hdll__a2bb2o_4_0/B2 sky130_fd_sc_hdll__a2bb2o_4_0/A1_N sky130_fd_sc_hdll__a2bb2o_4_0/A2_N
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__a2bb2o_4
Xsky130_fd_sc_hdll__nor4_2_0 sky130_fd_sc_hdll__nor4_2_0/C sky130_fd_sc_hdll__nor4_2_0/D
+ sky130_fd_sc_hdll__nor4_2_0/Y sky130_fd_sc_hdll__nor4_2_0/A sky130_fd_sc_hdll__nor4_2_0/B
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nor4_2
Xsky130_fd_sc_hdll__xor3_4_0 sky130_fd_sc_hdll__xor3_4_0/X sky130_fd_sc_hdll__xor3_4_0/C
+ sky130_fd_sc_hdll__xor3_4_0/B sky130_fd_sc_hdll__xor3_4_0/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__xor3_4
Xsky130_fd_sc_hdll__dlrtp_4_0 sky130_fd_sc_hdll__dlrtp_4_0/RESET_B sky130_fd_sc_hdll__dlrtp_4_0/D
+ sky130_fd_sc_hdll__dlrtp_4_0/GATE sky130_fd_sc_hdll__dlrtp_4_0/Q VGND VPWR VPWR
+ VGND sky130_fd_sc_hdll__dlrtp_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_0 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__isobufsrc_8_0 sky130_fd_sc_hdll__isobufsrc_8_0/A sky130_fd_sc_hdll__isobufsrc_8_0/X
+ sky130_fd_sc_hdll__isobufsrc_8_0/SLEEP VPWR VGND VGND VPWR sky130_fd_sc_hdll__isobufsrc_8
Xsky130_fd_sc_hdll__a32o_1_0 sky130_fd_sc_hdll__a32o_1_0/X sky130_fd_sc_hdll__a32o_1_0/A3
+ sky130_fd_sc_hdll__a32o_1_0/B2 sky130_fd_sc_hdll__a32o_1_0/B1 sky130_fd_sc_hdll__a32o_1_0/A1
+ sky130_fd_sc_hdll__a32o_1_0/A2 VGND VPWR VPWR VGND sky130_fd_sc_hdll__a32o_1
Xsky130_fd_sc_hdll__buf_4_0 VPWR VGND sky130_fd_sc_hdll__buf_4_0/X sky130_fd_sc_hdll__buf_4_0/A
+ VPWR VGND sky130_fd_sc_hdll__buf_4
Xsky130_fd_sc_hdll__inv_4_0 sky130_fd_sc_hdll__inv_4_0/Y sky130_fd_sc_hdll__inv_4_0/A
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__inv_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_33 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_44 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_55 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_66 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_77 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_88 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_99 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_11 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_22 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__dfrtp_2_0 sky130_fd_sc_hdll__dfrtp_2_0/RESET_B VPWR VGND sky130_fd_sc_hdll__dfrtp_2_0/Q
+ sky130_fd_sc_hdll__dfrtp_2_0/CLK sky130_fd_sc_hdll__dfrtp_2_0/D VPWR VGND sky130_fd_sc_hdll__dfrtp_2
Xsky130_fd_sc_hdll__nor4b_4_0 sky130_fd_sc_hdll__nor4b_4_0/B sky130_fd_sc_hdll__nor4b_4_0/A
+ sky130_fd_sc_hdll__nor4b_4_0/D_N sky130_fd_sc_hdll__nor4b_4_0/C sky130_fd_sc_hdll__nor4b_4_0/Y
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor4b_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_160 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a211oi_4_0 sky130_fd_sc_hdll__a211oi_4_0/A2 sky130_fd_sc_hdll__a211oi_4_0/A1
+ sky130_fd_sc_hdll__a211oi_4_0/C1 sky130_fd_sc_hdll__a211oi_4_0/Y sky130_fd_sc_hdll__a211oi_4_0/B1
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__a211oi_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_193 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_182 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_171 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__sdlclkp_2_0 sky130_fd_sc_hdll__sdlclkp_2_0/CLK VPWR VGND sky130_fd_sc_hdll__sdlclkp_2_0/GCLK
+ sky130_fd_sc_hdll__sdlclkp_2_0/SCE sky130_fd_sc_hdll__sdlclkp_2_0/GATE VPWR VGND
+ sky130_fd_sc_hdll__sdlclkp_2
Xsky130_fd_sc_hdll__a22oi_1_0 sky130_fd_sc_hdll__a22oi_1_0/B1 sky130_fd_sc_hdll__a22oi_1_0/A1
+ sky130_fd_sc_hdll__a22oi_1_0/B2 sky130_fd_sc_hdll__a22oi_1_0/A2 sky130_fd_sc_hdll__a22oi_1_0/Y
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__a22oi_1
Xsky130_fd_sc_hdll__muxb4to1_1_0 sky130_fd_sc_hdll__muxb4to1_1_0/S[0] sky130_fd_sc_hdll__muxb4to1_1_0/D[0]
+ sky130_fd_sc_hdll__muxb4to1_1_0/D[1] sky130_fd_sc_hdll__muxb4to1_1_0/S[1] sky130_fd_sc_hdll__muxb4to1_1_0/S[2]
+ sky130_fd_sc_hdll__muxb4to1_1_0/D[2] sky130_fd_sc_hdll__muxb4to1_1_0/D[3] sky130_fd_sc_hdll__muxb4to1_1_0/S[3]
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__muxb4to1_1_0/Z sky130_fd_sc_hdll__muxb4to1_1
Xsky130_fd_sc_hdll__o221a_1_0 sky130_fd_sc_hdll__o221a_1_0/A2 sky130_fd_sc_hdll__o221a_1_0/X
+ sky130_fd_sc_hdll__o221a_1_0/B1 sky130_fd_sc_hdll__o221a_1_0/C1 sky130_fd_sc_hdll__o221a_1_0/A1
+ sky130_fd_sc_hdll__o221a_1_0/B2 VPWR VGND VGND VPWR sky130_fd_sc_hdll__o221a_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_1 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__dlxtn_1_0 VGND VPWR sky130_fd_sc_hdll__dlxtn_1_0/Q sky130_fd_sc_hdll__dlxtn_1_0/GATE_N
+ sky130_fd_sc_hdll__dlxtn_1_0/D VPWR VGND sky130_fd_sc_hdll__dlxtn_1
Xsky130_fd_sc_hdll__and4_2_0 sky130_fd_sc_hdll__and4_2_0/X sky130_fd_sc_hdll__and4_2_0/C
+ sky130_fd_sc_hdll__and4_2_0/A sky130_fd_sc_hdll__and4_2_0/B sky130_fd_sc_hdll__and4_2_0/D
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__and4_2
Xsky130_fd_sc_hdll__o21bai_1_0 sky130_fd_sc_hdll__o21bai_1_0/A1 sky130_fd_sc_hdll__o21bai_1_0/Y
+ sky130_fd_sc_hdll__o21bai_1_0/B1_N sky130_fd_sc_hdll__o21bai_1_0/A2 VPWR VGND VPWR
+ VGND sky130_fd_sc_hdll__o21bai_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_12 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a22o_1_0 sky130_fd_sc_hdll__a22o_1_0/A1 sky130_fd_sc_hdll__a22o_1_0/A2
+ sky130_fd_sc_hdll__a22o_1_0/X sky130_fd_sc_hdll__a22o_1_0/B2 sky130_fd_sc_hdll__a22o_1_0/B1
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__a22o_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_23 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_34 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_45 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_56 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_67 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_78 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_89 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_320 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_150 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_161 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_194 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_183 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_172 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__sdfbbp_1_0 sky130_fd_sc_hdll__sdfbbp_1_0/SCD sky130_fd_sc_hdll__sdfbbp_1_0/SCE
+ sky130_fd_sc_hdll__sdfbbp_1_0/RESET_B VGND sky130_fd_sc_hdll__sdfbbp_1_0/CLK sky130_fd_sc_hdll__sdfbbp_1_0/Q
+ VPWR sky130_fd_sc_hdll__sdfbbp_1_0/D sky130_fd_sc_hdll__sdfbbp_1_0/Q_N sky130_fd_sc_hdll__sdfbbp_1_0/SET_B
+ VPWR VGND sky130_fd_sc_hdll__sdfbbp_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_2 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__or2_1_0 sky130_fd_sc_hdll__or2_1_0/A sky130_fd_sc_hdll__or2_1_0/X
+ sky130_fd_sc_hdll__or2_1_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__or2_1
Xsky130_fd_sc_hdll__a21oi_1_0 sky130_fd_sc_hdll__a21oi_1_0/A1 sky130_fd_sc_hdll__a21oi_1_0/B1
+ sky130_fd_sc_hdll__a21oi_1_0/Y sky130_fd_sc_hdll__a21oi_1_0/A2 VPWR VGND VPWR VGND
+ sky130_fd_sc_hdll__a21oi_1
Xsky130_fd_sc_hdll__nand4_2_0 sky130_fd_sc_hdll__nand4_2_0/B sky130_fd_sc_hdll__nand4_2_0/A
+ sky130_fd_sc_hdll__nand4_2_0/Y sky130_fd_sc_hdll__nand4_2_0/D sky130_fd_sc_hdll__nand4_2_0/C
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nand4_2
Xsky130_fd_sc_hdll__decap_6_0 VPWR VGND VPWR VGND sky130_fd_sc_hdll__decap_6
Xsky130_fd_sc_hdll__o211a_1_0 sky130_fd_sc_hdll__o211a_1_0/C1 sky130_fd_sc_hdll__o211a_1_0/B1
+ sky130_fd_sc_hdll__o211a_1_0/A2 sky130_fd_sc_hdll__o211a_1_0/A1 sky130_fd_sc_hdll__o211a_1_0/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o211a_1
Xsky130_fd_sc_hdll__and3b_2_0 VGND VPWR sky130_fd_sc_hdll__and3b_2_0/B sky130_fd_sc_hdll__and3b_2_0/X
+ sky130_fd_sc_hdll__and3b_2_0/A_N sky130_fd_sc_hdll__and3b_2_0/C VGND VPWR sky130_fd_sc_hdll__and3b_2
Xsky130_fd_sc_hdll__bufbuf_16_0 sky130_fd_sc_hdll__bufbuf_16_0/A sky130_fd_sc_hdll__bufbuf_16_0/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__bufbuf_16
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_35 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_46 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_57 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_68 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_79 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_13 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_310 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_321 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_24 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_140 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_151 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_162 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_195 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_184 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_173 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__xnor2_2_0 VGND VPWR sky130_fd_sc_hdll__xnor2_2_0/Y sky130_fd_sc_hdll__xnor2_2_0/A
+ sky130_fd_sc_hdll__xnor2_2_0/B VPWR VGND sky130_fd_sc_hdll__xnor2_2
Xsky130_fd_sc_hdll__clkbuf_8_0 sky130_fd_sc_hdll__clkbuf_8_0/X sky130_fd_sc_hdll__clkbuf_8_0/A
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__clkbuf_8
Xsky130_fd_sc_hdll__clkinv_8_0 sky130_fd_sc_hdll__clkinv_8_0/Y sky130_fd_sc_hdll__clkinv_8_0/A
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__clkinv_8
Xsky130_fd_sc_hdll__sdfxtp_4_0 VGND VPWR sky130_fd_sc_hdll__sdfxtp_4_0/SCD sky130_fd_sc_hdll__sdfxtp_4_0/D
+ sky130_fd_sc_hdll__sdfxtp_4_0/SCE sky130_fd_sc_hdll__sdfxtp_4_0/CLK sky130_fd_sc_hdll__sdfxtp_4_0/Q
+ VGND VPWR sky130_fd_sc_hdll__sdfxtp_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_3 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__or4b_2_0 sky130_fd_sc_hdll__or4b_2_0/C sky130_fd_sc_hdll__or4b_2_0/A
+ sky130_fd_sc_hdll__or4b_2_0/X sky130_fd_sc_hdll__or4b_2_0/B sky130_fd_sc_hdll__or4b_2_0/D_N
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__or4b_2
Xsky130_fd_sc_hdll__a2bb2o_2_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a2bb2o_2_0/B1
+ sky130_fd_sc_hdll__a2bb2o_2_0/A1_N sky130_fd_sc_hdll__a2bb2o_2_0/A2_N sky130_fd_sc_hdll__a2bb2o_2_0/X
+ sky130_fd_sc_hdll__a2bb2o_2_0/B2 sky130_fd_sc_hdll__a2bb2o_2
Xsky130_fd_sc_hdll__xor3_2_0 sky130_fd_sc_hdll__xor3_2_0/X sky130_fd_sc_hdll__xor3_2_0/C
+ sky130_fd_sc_hdll__xor3_2_0/B sky130_fd_sc_hdll__xor3_2_0/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__xor3_2
Xsky130_fd_sc_hdll__dlrtp_2_0 sky130_fd_sc_hdll__dlrtp_2_0/RESET_B sky130_fd_sc_hdll__dlrtp_2_0/D
+ sky130_fd_sc_hdll__dlrtp_2_0/GATE sky130_fd_sc_hdll__dlrtp_2_0/Q VGND VPWR VPWR
+ VGND sky130_fd_sc_hdll__dlrtp_2
Xsky130_fd_sc_hdll__buf_2_0 VPWR VGND sky130_fd_sc_hdll__buf_2_0/X sky130_fd_sc_hdll__buf_2_0/A
+ VPWR VGND sky130_fd_sc_hdll__buf_2
Xsky130_fd_sc_hdll__inv_12_0 sky130_fd_sc_hdll__inv_12_0/A sky130_fd_sc_hdll__inv_12_0/Y
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__inv_12
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_36 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_47 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_58 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_69 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_300 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_14 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_311 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_322 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_25 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__inv_2_0 sky130_fd_sc_hdll__inv_2_0/A sky130_fd_sc_hdll__inv_2_0/Y
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__inv_2
Xsky130_fd_sc_hdll__tap_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__tap_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_130 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_141 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_152 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__dlygate4sd3_1_0 sky130_fd_sc_hdll__dlygate4sd3_1_0/A sky130_fd_sc_hdll__dlygate4sd3_1_0/X
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__dlygate4sd3_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_196 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_185 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_174 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_163 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__muxb8to1_4_0 VGND sky130_fd_sc_hdll__muxb8to1_4_0/Z VPWR VGND
+ VPWR sky130_fd_sc_hdll__muxb8to1_4_0/S[6] sky130_fd_sc_hdll__muxb8to1_4_0/D[3] sky130_fd_sc_hdll__muxb8to1_4_0/D[0]
+ sky130_fd_sc_hdll__muxb8to1_4_0/D[4] sky130_fd_sc_hdll__muxb8to1_4_0/D[5] sky130_fd_sc_hdll__muxb8to1_4_0/D[2]
+ sky130_fd_sc_hdll__muxb8to1_4_0/D[1] sky130_fd_sc_hdll__muxb8to1_4_0/D[6] sky130_fd_sc_hdll__muxb8to1_4_0/S[2]
+ sky130_fd_sc_hdll__muxb8to1_4_0/S[3] sky130_fd_sc_hdll__muxb8to1_4_0/S[7] sky130_fd_sc_hdll__muxb8to1_4_0/S[0]
+ sky130_fd_sc_hdll__muxb8to1_4_0/S[1] sky130_fd_sc_hdll__muxb8to1_4_0/S[4] sky130_fd_sc_hdll__muxb8to1_4_0/S[5]
+ sky130_fd_sc_hdll__muxb8to1_4_0/D[7] sky130_fd_sc_hdll__muxb8to1_4
Xsky130_fd_sc_hdll__mux2_8_0 sky130_fd_sc_hdll__mux2_8_0/S sky130_fd_sc_hdll__mux2_8_0/A1
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__mux2_8_0/A0 sky130_fd_sc_hdll__mux2_8_0/X
+ sky130_fd_sc_hdll__mux2_8
Xsky130_fd_sc_hdll__o2bb2a_4_0 sky130_fd_sc_hdll__o2bb2a_4_0/A2_N sky130_fd_sc_hdll__o2bb2a_4_0/A1_N
+ sky130_fd_sc_hdll__o2bb2a_4_0/X sky130_fd_sc_hdll__o2bb2a_4_0/B2 sky130_fd_sc_hdll__o2bb2a_4_0/B1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o2bb2a_4
Xsky130_fd_sc_hdll__nor4b_2_0 sky130_fd_sc_hdll__nor4b_2_0/D_N sky130_fd_sc_hdll__nor4b_2_0/Y
+ sky130_fd_sc_hdll__nor4b_2_0/C sky130_fd_sc_hdll__nor4b_2_0/A sky130_fd_sc_hdll__nor4b_2_0/B
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nor4b_2
Xsky130_fd_sc_hdll__a211oi_2_0 sky130_fd_sc_hdll__a211oi_2_0/A2 sky130_fd_sc_hdll__a211oi_2_0/C1
+ sky130_fd_sc_hdll__a211oi_2_0/B1 sky130_fd_sc_hdll__a211oi_2_0/Y sky130_fd_sc_hdll__a211oi_2_0/A1
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__a211oi_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_4 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__or3_4_0 sky130_fd_sc_hdll__or3_4_0/A sky130_fd_sc_hdll__or3_4_0/X
+ sky130_fd_sc_hdll__or3_4_0/B sky130_fd_sc_hdll__or3_4_0/C VPWR VGND VPWR VGND sky130_fd_sc_hdll__or3_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_26 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_37 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_48 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_59 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_15 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_301 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_312 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_323 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o22ai_4_0 sky130_fd_sc_hdll__o22ai_4_0/A1 sky130_fd_sc_hdll__o22ai_4_0/Y
+ sky130_fd_sc_hdll__o22ai_4_0/A2 sky130_fd_sc_hdll__o22ai_4_0/B1 sky130_fd_sc_hdll__o22ai_4_0/B2
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o22ai_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_120 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_131 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_142 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_153 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_164 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_197 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_186 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_175 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__mux2_12_0 VPWR VGND VPWR VGND sky130_fd_sc_hdll__mux2_12_0/X sky130_fd_sc_hdll__mux2_12_0/S
+ sky130_fd_sc_hdll__mux2_12_0/A1 sky130_fd_sc_hdll__mux2_12_0/A0 sky130_fd_sc_hdll__mux2_12
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_5 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__inputiso1n_1_0 sky130_fd_sc_hdll__inputiso1n_1_0/A sky130_fd_sc_hdll__inputiso1n_1_0/SLEEP_B
+ sky130_fd_sc_hdll__inputiso1n_1_0/X VGND VPWR VGND VPWR sky130_fd_sc_hdll__inputiso1n_1
Xsky130_fd_sc_hdll__o21a_1_0 sky130_fd_sc_hdll__o21a_1_0/X sky130_fd_sc_hdll__o21a_1_0/A1
+ sky130_fd_sc_hdll__o21a_1_0/B1 sky130_fd_sc_hdll__o21a_1_0/A2 VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__o21a_1
Xsky130_fd_sc_hdll__nand2b_4_0 sky130_fd_sc_hdll__nand2b_4_0/B sky130_fd_sc_hdll__nand2b_4_0/A_N
+ sky130_fd_sc_hdll__nand2b_4_0/Y VGND VPWR VGND VPWR sky130_fd_sc_hdll__nand2b_4
Xsky130_fd_sc_hdll__decap_4_0 VGND VPWR VPWR VGND sky130_fd_sc_hdll__decap_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_27 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_38 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_49 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o211ai_4_0 sky130_fd_sc_hdll__o211ai_4_0/A1 sky130_fd_sc_hdll__o211ai_4_0/B1
+ sky130_fd_sc_hdll__o211ai_4_0/A2 sky130_fd_sc_hdll__o211ai_4_0/C1 sky130_fd_sc_hdll__o211ai_4_0/Y
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o211ai_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_16 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_302 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_313 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_324 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_110 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_121 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_132 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_143 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_154 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nor2_1_0 sky130_fd_sc_hdll__nor2_1_0/B sky130_fd_sc_hdll__nor2_1_0/Y
+ sky130_fd_sc_hdll__nor2_1_0/A VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor2_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_198 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_187 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nand4b_1_0 sky130_fd_sc_hdll__nand4b_1_0/Y sky130_fd_sc_hdll__nand4b_1_0/C
+ sky130_fd_sc_hdll__nand4b_1_0/D sky130_fd_sc_hdll__nand4b_1_0/A_N sky130_fd_sc_hdll__nand4b_1_0/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__nand4b_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_176 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_165 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__clkmux2_4_0 VGND VPWR sky130_fd_sc_hdll__clkmux2_4_0/S sky130_fd_sc_hdll__clkmux2_4_0/A1
+ sky130_fd_sc_hdll__clkmux2_4_0/A0 sky130_fd_sc_hdll__clkmux2_4_0/X VPWR VGND sky130_fd_sc_hdll__clkmux2_4
Xsky130_fd_sc_hdll__o21ai_4_0 sky130_fd_sc_hdll__o21ai_4_0/Y sky130_fd_sc_hdll__o21ai_4_0/B1
+ sky130_fd_sc_hdll__o21ai_4_0/A2 sky130_fd_sc_hdll__o21ai_4_0/A1 VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__o21ai_4
Xsky130_fd_sc_hdll__clkbuf_6_0 sky130_fd_sc_hdll__clkbuf_6_0/A sky130_fd_sc_hdll__clkbuf_6_0/X
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__clkbuf_6
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_6 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__sdfxtp_2_0 VPWR VGND sky130_fd_sc_hdll__sdfxtp_2_0/SCE sky130_fd_sc_hdll__sdfxtp_2_0/D
+ sky130_fd_sc_hdll__sdfxtp_2_0/SCD sky130_fd_sc_hdll__sdfxtp_2_0/Q sky130_fd_sc_hdll__sdfxtp_2_0/CLK
+ VGND VPWR sky130_fd_sc_hdll__sdfxtp_2
Xsky130_fd_sc_hdll__einvn_8_0 sky130_fd_sc_hdll__einvn_8_0/A sky130_fd_sc_hdll__einvn_8_0/TE_B
+ sky130_fd_sc_hdll__einvn_8_0/Z VGND VPWR VPWR VGND sky130_fd_sc_hdll__einvn_8
Xsky130_fd_sc_hdll__nor4bb_4_0 sky130_fd_sc_hdll__nor4bb_4_0/D_N sky130_fd_sc_hdll__nor4bb_4_0/Y
+ sky130_fd_sc_hdll__nor4bb_4_0/A sky130_fd_sc_hdll__nor4bb_4_0/B sky130_fd_sc_hdll__nor4bb_4_0/C_N
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nor4bb_4
Xsky130_fd_sc_hdll__o2bb2ai_1_0 sky130_fd_sc_hdll__o2bb2ai_1_0/Y sky130_fd_sc_hdll__o2bb2ai_1_0/A1_N
+ sky130_fd_sc_hdll__o2bb2ai_1_0/A2_N sky130_fd_sc_hdll__o2bb2ai_1_0/B2 sky130_fd_sc_hdll__o2bb2ai_1_0/B1
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__o2bb2ai_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_28 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_39 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__isobufsrc_4_0 sky130_fd_sc_hdll__isobufsrc_4_0/A sky130_fd_sc_hdll__isobufsrc_4_0/X
+ sky130_fd_sc_hdll__isobufsrc_4_0/SLEEP VGND VPWR VGND VPWR sky130_fd_sc_hdll__isobufsrc_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_17 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_303 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_314 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_325 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__bufbuf_8_0 sky130_fd_sc_hdll__bufbuf_8_0/A sky130_fd_sc_hdll__bufbuf_8_0/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__bufbuf_8
Xsky130_fd_sc_hdll__bufinv_8_0 sky130_fd_sc_hdll__bufinv_8_0/A sky130_fd_sc_hdll__bufinv_8_0/Y
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__bufinv_8
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_100 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_111 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_122 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_133 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_144 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_155 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_199 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_188 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_177 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_166 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__fill_8_0 VGND VPWR VPWR VGND sky130_fd_sc_hdll__fill_8
Xsky130_fd_sc_hdll__muxb8to1_2_0 sky130_fd_sc_hdll__muxb8to1_2_0/Z VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__muxb8to1_2_0/D[2] sky130_fd_sc_hdll__muxb8to1_2_0/D[1] sky130_fd_sc_hdll__muxb8to1_2_0/S[7]
+ sky130_fd_sc_hdll__muxb8to1_2_0/S[6] sky130_fd_sc_hdll__muxb8to1_2_0/S[5] sky130_fd_sc_hdll__muxb8to1_2_0/S[4]
+ sky130_fd_sc_hdll__muxb8to1_2_0/S[3] sky130_fd_sc_hdll__muxb8to1_2_0/S[2] sky130_fd_sc_hdll__muxb8to1_2_0/S[1]
+ sky130_fd_sc_hdll__muxb8to1_2_0/S[0] sky130_fd_sc_hdll__muxb8to1_2_0/D[7] sky130_fd_sc_hdll__muxb8to1_2_0/D[6]
+ sky130_fd_sc_hdll__muxb8to1_2_0/D[5] sky130_fd_sc_hdll__muxb8to1_2_0/D[4] sky130_fd_sc_hdll__muxb8to1_2_0/D[3]
+ sky130_fd_sc_hdll__muxb8to1_2_0/D[0] sky130_fd_sc_hdll__muxb8to1_2
Xsky130_fd_sc_hdll__and2_1_0 VPWR VGND sky130_fd_sc_hdll__and2_1_0/X sky130_fd_sc_hdll__and2_1_0/B
+ sky130_fd_sc_hdll__and2_1_0/A VPWR VGND sky130_fd_sc_hdll__and2_1
Xsky130_fd_sc_hdll__o2bb2a_2_0 sky130_fd_sc_hdll__o2bb2a_2_0/A1_N sky130_fd_sc_hdll__o2bb2a_2_0/X
+ sky130_fd_sc_hdll__o2bb2a_2_0/A2_N sky130_fd_sc_hdll__o2bb2a_2_0/B2 sky130_fd_sc_hdll__o2bb2a_2_0/B1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o2bb2a_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_7 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__sedfxbp_1_0 VGND VPWR sky130_fd_sc_hdll__sedfxbp_1_0/SCE sky130_fd_sc_hdll__sedfxbp_1_0/Q
+ sky130_fd_sc_hdll__sedfxbp_1_0/D sky130_fd_sc_hdll__sedfxbp_1_0/DE sky130_fd_sc_hdll__sedfxbp_1_0/SCD
+ sky130_fd_sc_hdll__sedfxbp_1_0/Q_N sky130_fd_sc_hdll__sedfxbp_1_0/CLK VPWR VGND
+ sky130_fd_sc_hdll__sedfxbp_1
Xsky130_fd_sc_hdll__a221oi_4_0 sky130_fd_sc_hdll__a221oi_4_0/A2 sky130_fd_sc_hdll__a221oi_4_0/Y
+ sky130_fd_sc_hdll__a221oi_4_0/C1 sky130_fd_sc_hdll__a221oi_4_0/A1 sky130_fd_sc_hdll__a221oi_4_0/B2
+ sky130_fd_sc_hdll__a221oi_4_0/B1 VGND VPWR VPWR VGND sky130_fd_sc_hdll__a221oi_4
Xsky130_fd_sc_hdll__o22a_4_0 sky130_fd_sc_hdll__o22a_4_0/B2 sky130_fd_sc_hdll__o22a_4_0/B1
+ sky130_fd_sc_hdll__o22a_4_0/X sky130_fd_sc_hdll__o22a_4_0/A1 sky130_fd_sc_hdll__o22a_4_0/A2
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o22a_4
Xsky130_fd_sc_hdll__a32oi_1_0 sky130_fd_sc_hdll__a32oi_1_0/A2 sky130_fd_sc_hdll__a32oi_1_0/Y
+ sky130_fd_sc_hdll__a32oi_1_0/A1 sky130_fd_sc_hdll__a32oi_1_0/B2 sky130_fd_sc_hdll__a32oi_1_0/B1
+ sky130_fd_sc_hdll__a32oi_1_0/A3 VGND VPWR VPWR VGND sky130_fd_sc_hdll__a32oi_1
Xsky130_fd_sc_hdll__or3_2_0 sky130_fd_sc_hdll__or3_2_0/A sky130_fd_sc_hdll__or3_2_0/B
+ sky130_fd_sc_hdll__or3_2_0/X sky130_fd_sc_hdll__or3_2_0/C VGND VPWR VPWR VGND sky130_fd_sc_hdll__or3_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_29 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_304 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_315 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_18 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_101 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_112 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_123 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_134 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_145 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_156 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_189 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_178 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_167 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
.ends
