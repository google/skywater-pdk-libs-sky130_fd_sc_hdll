* File: sky130_fd_sc_hdll__probec_p_8.pxi.spice
* Created: Wed Sep  2 08:50:19 2020
* 
x_PM_SKY130_FD_SC_HDLL__PROBEC_P_8%A N_A_c_118_n N_A_M1001_g N_A_M1002_g
+ N_A_c_119_n N_A_M1009_g N_A_M1006_g N_A_M1015_g N_A_c_120_n N_A_M1019_g A
+ N_A_c_116_n N_A_c_117_n PM_SKY130_FD_SC_HDLL__PROBEC_P_8%A
x_PM_SKY130_FD_SC_HDLL__PROBEC_P_8%A_27_47# N_A_27_47#_M1002_d
+ N_A_27_47#_M1006_d N_A_27_47#_M1001_d N_A_27_47#_M1009_d N_A_27_47#_c_214_n
+ N_A_27_47#_M1000_g N_A_27_47#_M1004_g N_A_27_47#_M1008_g N_A_27_47#_c_215_n
+ N_A_27_47#_M1003_g N_A_27_47#_c_216_n N_A_27_47#_M1005_g N_A_27_47#_M1011_g
+ N_A_27_47#_M1013_g N_A_27_47#_c_217_n N_A_27_47#_M1007_g N_A_27_47#_c_218_n
+ N_A_27_47#_M1010_g N_A_27_47#_M1016_g N_A_27_47#_M1018_g N_A_27_47#_c_219_n
+ N_A_27_47#_M1012_g N_A_27_47#_c_220_n N_A_27_47#_M1014_g N_A_27_47#_M1020_g
+ N_A_27_47#_M1021_g N_A_27_47#_c_221_n N_A_27_47#_M1017_g N_A_27_47#_c_222_n
+ N_A_27_47#_c_430_p N_A_27_47#_c_223_n N_A_27_47#_c_224_n N_A_27_47#_c_207_n
+ N_A_27_47#_c_208_n N_A_27_47#_c_246_n N_A_27_47#_c_311_p N_A_27_47#_c_209_n
+ N_A_27_47#_c_210_n N_A_27_47#_c_211_n N_A_27_47#_c_226_n N_A_27_47#_c_212_n
+ N_A_27_47#_c_262_n N_A_27_47#_c_213_n
+ PM_SKY130_FD_SC_HDLL__PROBEC_P_8%A_27_47#
x_PM_SKY130_FD_SC_HDLL__PROBEC_P_8%VPWR N_VPWR_M1001_s N_VPWR_M1019_s
+ N_VPWR_M1003_s N_VPWR_M1007_s N_VPWR_M1012_s N_VPWR_M1017_s N_VPWR_c_490_n
+ N_VPWR_c_491_n N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_494_n N_VPWR_c_495_n
+ N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_500_n
+ N_VPWR_c_501_n VPWR VPWR N_VPWR_c_487_n N_VPWR_R1_neg N_VPWR_c_504_n
+ N_VPWR_c_505_n N_VPWR_c_506_n N_VPWR_c_507_n N_VPWR_c_508_n N_VPWR_c_509_n
+ N_VPWR_c_510_n N_VPWR_c_489_n PM_SKY130_FD_SC_HDLL__PROBEC_P_8%VPWR
x_PM_SKY130_FD_SC_HDLL__PROBEC_P_8%A_399_297# N_A_399_297#_M1004_s
+ N_A_399_297#_M1011_s N_A_399_297#_M1016_s N_A_399_297#_M1020_s
+ N_A_399_297#_M1000_d N_A_399_297#_M1005_d N_A_399_297#_M1010_d
+ N_A_399_297#_M1014_d N_A_399_297#_c_630_n N_A_399_297#_c_631_n
+ N_A_399_297#_c_612_n N_A_399_297#_c_613_n N_A_399_297#_c_620_n
+ N_A_399_297#_c_621_n N_A_399_297#_c_666_n N_A_399_297#_c_670_n
+ N_A_399_297#_c_614_n N_A_399_297#_c_622_n N_A_399_297#_c_682_n
+ N_A_399_297#_c_686_n N_A_399_297#_c_690_n N_A_399_297#_c_693_n
+ N_A_399_297#_c_615_n N_A_399_297#_c_623_n N_A_399_297#_c_704_n
+ N_A_399_297#_c_624_n N_A_399_297#_c_708_n N_A_399_297#_c_785_n
+ N_A_399_297#_c_625_n N_A_399_297#_c_616_n N_A_399_297#_c_617_n
+ N_A_399_297#_c_618_n N_A_399_297#_R0_neg N_A_399_297#_c_619_n
+ N_A_399_297#_c_629_n PM_SKY130_FD_SC_HDLL__PROBEC_P_8%A_399_297#
x_PM_SKY130_FD_SC_HDLL__PROBEC_P_8%VGND N_VGND_M1002_s N_VGND_M1015_s
+ N_VGND_M1008_d N_VGND_M1013_d N_VGND_M1018_d N_VGND_M1021_d N_VGND_c_851_n
+ N_VGND_c_852_n N_VGND_c_853_n N_VGND_c_854_n N_VGND_c_855_n N_VGND_c_856_n
+ N_VGND_c_857_n N_VGND_c_858_n N_VGND_c_859_n N_VGND_c_860_n N_VGND_c_861_n
+ VGND VGND N_VGND_c_862_n N_VGND_R2_neg N_VGND_c_864_n N_VGND_c_865_n
+ N_VGND_c_866_n N_VGND_c_867_n N_VGND_c_868_n N_VGND_c_869_n N_VGND_c_870_n
+ N_VGND_c_871_n VGND VGND N_VGND_c_872_n PM_SKY130_FD_SC_HDLL__PROBEC_P_8%VGND
x_PM_SKY130_FD_SC_HDLL__PROBEC_P_8%X X N_X_c_991_n N_X_c_992_n N_X_R0_pos
+ PM_SKY130_FD_SC_HDLL__PROBEC_P_8%X
cc_1 VNB N_A_M1002_g 0.0229771f $X=-1.26 $Y=-1.17 $X2=0.52 $Y2=0.56
cc_2 VNB N_A_M1006_g 0.0175585f $X=-1.26 $Y=-1.17 $X2=0.99 $Y2=0.56
cc_3 VNB N_A_M1015_g 0.0175958f $X=-1.26 $Y=-1.17 $X2=1.41 $Y2=0.56
cc_4 VNB N_A_c_116_n 0.00614839f $X=-1.26 $Y=-1.17 $X2=0.985 $Y2=1.16
cc_5 VNB N_A_c_117_n 0.104335f $X=-1.26 $Y=-1.17 $X2=1.41 $Y2=1.212
cc_6 VNB N_A_27_47#_M1004_g 0.0179864f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_M1008_g 0.0176972f $X=-1.26 $Y=-1.17 $X2=0.61 $Y2=1.105
cc_8 VNB N_A_27_47#_M1011_g 0.0183398f $X=-1.26 $Y=-1.17 $X2=0.985 $Y2=1.16
cc_9 VNB N_A_27_47#_M1013_g 0.0183398f $X=-1.26 $Y=-1.17 $X2=0.305 $Y2=1.175
cc_10 VNB N_A_27_47#_M1016_g 0.0183352f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_M1018_g 0.0178188f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_M1020_g 0.0173202f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_M1021_g 0.0237845f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_207_n 0.0021789f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_208_n 0.00260199f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_209_n 0.00459766f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_210_n 0.00158168f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_211_n 0.00478392f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_212_n 0.00263026f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_213_n 0.210788f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_487_n 0.0270715f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_22 VNB N_VPWR_R1_neg 0.164147f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_489_n 0.210136f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_24 VNB N_A_399_297#_c_612_n 0.00238654f $X=-1.26 $Y=-1.17 $X2=0.99 $Y2=1.212
cc_25 VNB N_A_399_297#_c_613_n 0.00156403f $X=-1.26 $Y=-1.17 $X2=1.41 $Y2=1.212
cc_26 VNB N_A_399_297#_c_614_n 0.00229857f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_27 VNB N_A_399_297#_c_615_n 0.00184854f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_28 VNB N_A_399_297#_c_616_n 0.00128963f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_29 VNB N_A_399_297#_c_617_n 0.218348f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_30 VNB N_A_399_297#_c_618_n 0.00327305f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_31 VNB N_A_399_297#_c_619_n 0.00208123f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_851_n 0.00473987f $X=-1.26 $Y=-1.17 $X2=1.435 $Y2=1.985
cc_33 VNB N_VGND_c_852_n 0.0042804f $X=-1.26 $Y=-1.17 $X2=0.305 $Y2=1.16
cc_34 VNB N_VGND_c_853_n 0.0173083f $X=-1.26 $Y=-1.17 $X2=0.495 $Y2=1.212
cc_35 VNB N_VGND_c_854_n 0.00414011f $X=-1.26 $Y=-1.17 $X2=0.985 $Y2=1.16
cc_36 VNB N_VGND_c_855_n 0.0166933f $X=-1.26 $Y=-1.17 $X2=0.99 $Y2=1.212
cc_37 VNB N_VGND_c_856_n 0.00414011f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_857_n 0.0168835f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_858_n 0.00414011f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_859_n 0.030574f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_860_n 0.0175114f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_861_n 0.00480536f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_862_n 0.0381666f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_44 VNB N_VGND_R2_neg 0.16786f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_864_n 0.0155708f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_865_n 0.0159859f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_866_n 0.0182824f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_867_n 0.00535855f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_868_n 0.00573982f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_869_n 0.00515959f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_870_n 0.00515959f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_871_n 0.00510782f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_872_n 0.255189f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_54 VNB N_X_c_991_n 0.0380493f $X=-1.26 $Y=-1.17 $X2=0.52 $Y2=1.015
cc_55 VNB N_X_c_992_n 0.028536f $X=-1.26 $Y=-1.17 $X2=0.965 $Y2=1.41
cc_56 VNB N_X_R0_pos 0.147985f $X=-1.26 $Y=-1.17 $X2=0.965 $Y2=1.985
cc_57 VNB M5_872_N71# 8.97967e-19 $X=-1.26 $Y=-1.17 $X2=0.495 $Y2=1.41
cc_58 VNB M5_872_595# 8.97967e-19 $X=-1.26 $Y=-1.17 $X2=0.495 $Y2=1.41
cc_59 VPB N_A_c_118_n 0.0198895f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_60 VPB N_A_c_119_n 0.0157272f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_61 VPB N_A_c_120_n 0.0157116f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_62 VPB N_A_c_117_n 0.0331092f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=1.212
cc_63 VPB N_A_27_47#_c_214_n 0.0159578f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_64 VPB N_A_27_47#_c_215_n 0.0156957f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.212
cc_65 VPB N_A_27_47#_c_216_n 0.0158129f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.212
cc_66 VPB N_A_27_47#_c_217_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.175
cc_67 VPB N_A_27_47#_c_218_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_27_47#_c_219_n 0.0157407f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_27_47#_c_220_n 0.0155986f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_27_47#_c_221_n 0.0207627f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_47#_c_222_n 0.0290878f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_47#_c_223_n 0.00197463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_47#_c_224_n 0.00872632f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_47#_c_210_n 0.0037956f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_47#_c_226_n 0.00263651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_47#_c_213_n 0.0521998f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_490_n 0.00466368f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_78 VPB N_VPWR_c_491_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_492_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.212
cc_80 VPB N_VPWR_c_493_n 0.017949f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.212
cc_81 VPB N_VPWR_c_494_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.212
cc_82 VPB N_VPWR_c_495_n 0.017949f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.212
cc_83 VPB N_VPWR_c_496_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_497_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_498_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_499_n 0.045966f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_500_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_501_n 0.00574121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_487_n 0.0105622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_R1_neg 0.00343944f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_504_n 0.0178692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_505_n 0.0143948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_506_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_507_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_508_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_509_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_510_n 0.00510905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_489_n 0.0430632f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_399_297#_c_620_n 0.00198493f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.212
cc_100 VPB N_A_399_297#_c_621_n 0.00181449f $X=-0.19 $Y=1.305 $X2=0.305
+ $Y2=1.175
cc_101 VPB N_A_399_297#_c_622_n 0.00147108f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_399_297#_c_623_n 0.00150412f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_399_297#_c_624_n 0.00180391f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_399_297#_c_625_n 0.0040135f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_399_297#_c_616_n 9.69885e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_399_297#_c_618_n 0.00671938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_399_297#_c_619_n 0.00159673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_399_297#_c_629_n 0.00539269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_X_c_991_n 0.0088462f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.015
cc_110 VPB N_X_c_992_n 0.00425834f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_111 VPB N_X_R0_pos 0.00880667f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_112 N_A_c_120_n N_A_27_47#_c_214_n 0.0257643f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_M1015_g N_A_27_47#_M1004_g 0.0206587f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_114 N_A_c_118_n N_A_27_47#_c_222_n 0.010616f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A_c_119_n N_A_27_47#_c_222_n 0.0013412f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A_c_118_n N_A_27_47#_c_223_n 0.012939f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A_c_119_n N_A_27_47#_c_223_n 0.0129506f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A_c_116_n N_A_27_47#_c_223_n 0.059354f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_c_117_n N_A_27_47#_c_223_n 0.00702443f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_120 N_A_c_118_n N_A_27_47#_c_224_n 0.001334f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_c_116_n N_A_27_47#_c_224_n 0.0232414f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_c_117_n N_A_27_47#_c_224_n 0.00618163f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_123 N_A_M1002_g N_A_27_47#_c_207_n 0.0099777f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_124 N_A_M1006_g N_A_27_47#_c_207_n 0.00994697f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_125 N_A_c_116_n N_A_27_47#_c_207_n 0.0580113f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A_c_117_n N_A_27_47#_c_207_n 0.00317014f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_127 N_A_M1002_g N_A_27_47#_c_208_n 3.62277e-19 $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_128 N_A_c_116_n N_A_27_47#_c_208_n 0.0244894f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A_c_117_n N_A_27_47#_c_208_n 0.00736968f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_130 N_A_c_118_n N_A_27_47#_c_246_n 0.00134387f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A_c_119_n N_A_27_47#_c_246_n 0.0106596f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A_c_120_n N_A_27_47#_c_246_n 0.01034f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A_M1006_g N_A_27_47#_c_209_n 0.0013128f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_134 N_A_M1015_g N_A_27_47#_c_209_n 0.00576719f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_135 N_A_c_117_n N_A_27_47#_c_209_n 0.00359882f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_136 N_A_c_119_n N_A_27_47#_c_210_n 3.87554e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A_c_120_n N_A_27_47#_c_210_n 0.00175411f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_c_116_n N_A_27_47#_c_210_n 0.00208972f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A_c_117_n N_A_27_47#_c_210_n 0.00899686f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_140 N_A_c_119_n N_A_27_47#_c_226_n 0.00101982f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_c_120_n N_A_27_47#_c_226_n 0.01254f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_c_117_n N_A_27_47#_c_226_n 0.00786701f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_143 N_A_M1006_g N_A_27_47#_c_212_n 2.0357e-19 $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_144 N_A_M1015_g N_A_27_47#_c_212_n 0.00958725f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_145 N_A_c_117_n N_A_27_47#_c_212_n 0.00235176f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_146 N_A_c_116_n N_A_27_47#_c_262_n 0.0133942f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_c_117_n N_A_27_47#_c_262_n 0.00585963f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_148 N_A_c_116_n N_A_27_47#_c_213_n 2.12786e-19 $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_c_117_n N_A_27_47#_c_213_n 0.0196691f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_150 N_A_c_118_n N_VPWR_c_490_n 0.00364171f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_c_119_n N_VPWR_c_490_n 0.00229017f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_c_119_n N_VPWR_c_491_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_c_120_n N_VPWR_c_491_n 0.00673617f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_c_120_n N_VPWR_c_492_n 0.00288623f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_c_118_n N_VPWR_c_504_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_c_118_n N_VPWR_c_489_n 0.0123564f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_c_119_n N_VPWR_c_489_n 0.0114449f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_c_120_n N_VPWR_c_489_n 0.0105421f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_M1015_g N_A_399_297#_c_630_n 0.00101353f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_160 N_A_c_120_n N_A_399_297#_c_631_n 0.0015039f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A_M1015_g N_A_399_297#_c_613_n 3.86822e-19 $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_162 N_A_c_120_n N_A_399_297#_c_621_n 3.99559e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A_c_120_n N_A_399_297#_c_616_n 0.0047579f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_c_116_n N_A_399_297#_c_616_n 0.00109767f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_M1015_g N_A_399_297#_c_617_n 2.53636e-19 $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_166 N_A_c_116_n N_A_399_297#_c_617_n 4.60567e-19 $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_c_117_n N_A_399_297#_c_617_n 0.00120532f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_168 N_A_c_116_n N_A_399_297#_c_618_n 0.0010351f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_M1002_g N_VGND_c_851_n 0.00308601f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_170 N_A_M1006_g N_VGND_c_851_n 0.0016661f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_171 N_A_M1015_g N_VGND_c_852_n 0.00234309f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_172 N_A_M1006_g N_VGND_c_864_n 0.00439206f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_173 N_A_M1015_g N_VGND_c_864_n 0.00439206f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_174 N_A_M1002_g N_VGND_c_866_n 0.00439206f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_175 N_A_M1002_g N_VGND_c_872_n 0.00688232f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_176 N_A_M1006_g N_VGND_c_872_n 0.00582638f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_177 N_A_M1015_g N_VGND_c_872_n 0.00916272f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_178 N_A_c_118_n N_X_c_991_n 2.38745e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_M1002_g N_X_c_991_n 7.27292e-19 $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_180 N_A_c_117_n N_X_c_991_n 5.54474e-19 $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_181 N_A_c_116_n N_X_c_992_n 0.00432327f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_c_117_n N_X_c_992_n 0.00179877f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_183 N_A_c_118_n N_X_R0_pos 0.00272812f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A_M1002_g N_X_R0_pos 0.00288293f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_185 N_A_c_119_n N_X_R0_pos 0.00255056f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_186 N_A_M1006_g N_X_R0_pos 0.00239057f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_187 N_A_c_116_n N_X_R0_pos 0.00318199f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A_c_117_n N_X_R0_pos 0.00554953f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_189 N_A_27_47#_c_223_n N_VPWR_M1001_s 0.00169388f $X=1.035 $Y=1.53 $X2=-1.26
+ $Y2=-1.17
cc_190 N_A_27_47#_c_226_n N_VPWR_M1019_s 0.00168556f $X=1.507 $Y=1.53 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_222_n N_VPWR_c_490_n 0.0304489f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_192 N_A_27_47#_c_223_n N_VPWR_c_490_n 0.0149985f $X=1.035 $Y=1.53 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_246_n N_VPWR_c_490_n 0.0304489f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_194 N_A_27_47#_c_246_n N_VPWR_c_491_n 0.0216675f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_214_n N_VPWR_c_492_n 0.00288623f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_246_n N_VPWR_c_492_n 0.0368456f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_211_n N_VPWR_c_492_n 0.00624749f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_226_n N_VPWR_c_492_n 0.00246523f $X=1.507 $Y=1.53 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_214_n N_VPWR_c_493_n 0.00673617f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_215_n N_VPWR_c_493_n 0.00673617f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_215_n N_VPWR_c_494_n 0.00288623f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_216_n N_VPWR_c_494_n 0.0028874f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A_27_47#_c_216_n N_VPWR_c_495_n 0.00673617f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_217_n N_VPWR_c_495_n 0.00673617f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_c_217_n N_VPWR_c_496_n 0.00173895f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_218_n N_VPWR_c_496_n 0.00173895f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_218_n N_VPWR_c_497_n 0.00673617f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_c_219_n N_VPWR_c_497_n 0.00673617f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_219_n N_VPWR_c_498_n 0.00173895f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_220_n N_VPWR_c_498_n 0.00233618f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_c_213_n N_VPWR_c_498_n 9.15469e-19 $X=5.17 $Y=1.217 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_221_n N_VPWR_c_499_n 0.00417286f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_220_n N_VPWR_c_500_n 0.00673617f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_c_221_n N_VPWR_c_500_n 0.00673617f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_221_n N_VPWR_c_487_n 0.00191847f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_220_n N_VPWR_R1_neg 0.00140106f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_217 N_A_27_47#_c_221_n N_VPWR_R1_neg 9.16152e-19 $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A_27_47#_c_222_n N_VPWR_c_504_n 0.0210596f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_219 N_A_27_47#_M1001_d N_VPWR_c_489_n 0.00208639f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_M1009_d N_VPWR_c_489_n 0.00660897f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_c_214_n N_VPWR_c_489_n 0.0106095f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_222 N_A_27_47#_c_215_n N_VPWR_c_489_n 0.0105843f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A_27_47#_c_216_n N_VPWR_c_489_n 0.011575f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_224 N_A_27_47#_c_217_n N_VPWR_c_489_n 0.0117593f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A_27_47#_c_218_n N_VPWR_c_489_n 0.0117593f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_226 N_A_27_47#_c_219_n N_VPWR_c_489_n 0.0117593f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_227 N_A_27_47#_c_220_n N_VPWR_c_489_n 0.0105843f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_221_n N_VPWR_c_489_n 0.0110853f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_229 N_A_27_47#_c_222_n N_VPWR_c_489_n 0.0124725f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_230 N_A_27_47#_c_246_n N_VPWR_c_489_n 0.012178f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_231 N_A_27_47#_M1004_g N_A_399_297#_c_630_n 0.00644604f $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_M1008_g N_A_399_297#_c_630_n 0.00635074f $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_M1011_g N_A_399_297#_c_630_n 0.00100159f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_311_p N_A_399_297#_c_630_n 0.00466114f $X=1.2 $Y=0.42 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_214_n N_A_399_297#_c_631_n 0.0115852f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_215_n N_A_399_297#_c_631_n 0.0115852f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_c_216_n N_A_399_297#_c_631_n 0.00151073f $X=2.845 $Y=1.41
+ $X2=0 $Y2=0
cc_238 N_A_27_47#_c_246_n N_A_399_297#_c_631_n 0.00539931f $X=1.2 $Y=1.63 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_M1008_g N_A_399_297#_c_612_n 0.00859181f $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_M1011_g N_A_399_297#_c_612_n 0.00900524f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_211_n N_A_399_297#_c_612_n 0.042103f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_213_n N_A_399_297#_c_612_n 0.00418716f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_243 N_A_27_47#_M1004_g N_A_399_297#_c_613_n 0.0028318f $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_M1008_g N_A_399_297#_c_613_n 9.9253e-19 $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_211_n N_A_399_297#_c_613_n 0.0255515f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_212_n N_A_399_297#_c_613_n 0.00742303f $X=1.507 $Y=0.82
+ $X2=0 $Y2=0
cc_247 N_A_27_47#_c_213_n N_A_399_297#_c_613_n 0.00203093f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_248 N_A_27_47#_c_215_n N_A_399_297#_c_620_n 0.0127878f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_216_n N_A_399_297#_c_620_n 0.013865f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_211_n N_A_399_297#_c_620_n 0.0351537f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_213_n N_A_399_297#_c_620_n 0.00599265f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_252 N_A_27_47#_c_214_n N_A_399_297#_c_621_n 0.00394481f $X=1.905 $Y=1.41
+ $X2=0 $Y2=0
cc_253 N_A_27_47#_c_215_n N_A_399_297#_c_621_n 0.00196108f $X=2.375 $Y=1.41
+ $X2=0 $Y2=0
cc_254 N_A_27_47#_c_211_n N_A_399_297#_c_621_n 0.0221531f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_226_n N_A_399_297#_c_621_n 0.00741886f $X=1.507 $Y=1.53
+ $X2=0 $Y2=0
cc_256 N_A_27_47#_c_213_n N_A_399_297#_c_621_n 0.0059948f $X=5.17 $Y=1.217 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_M1008_g N_A_399_297#_c_666_n 5.21968e-19 $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_M1011_g N_A_399_297#_c_666_n 0.00682312f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_M1013_g N_A_399_297#_c_666_n 0.00682312f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_M1016_g N_A_399_297#_c_666_n 5.26907e-19 $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_215_n N_A_399_297#_c_670_n 7.24675e-19 $X=2.375 $Y=1.41
+ $X2=0 $Y2=0
cc_262 N_A_27_47#_c_216_n N_A_399_297#_c_670_n 0.0125412f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_c_217_n N_A_399_297#_c_670_n 0.0125412f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_218_n N_A_399_297#_c_670_n 7.3868e-19 $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_M1013_g N_A_399_297#_c_614_n 0.00900524f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_M1016_g N_A_399_297#_c_614_n 0.00900524f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_211_n N_A_399_297#_c_614_n 0.0388885f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_213_n N_A_399_297#_c_614_n 0.00433688f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_269 N_A_27_47#_c_217_n N_A_399_297#_c_622_n 0.0138887f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_218_n N_A_399_297#_c_622_n 0.0138887f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_211_n N_A_399_297#_c_622_n 0.0311906f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_213_n N_A_399_297#_c_622_n 0.00707008f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_273 N_A_27_47#_M1013_g N_A_399_297#_c_682_n 5.26907e-19 $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_M1016_g N_A_399_297#_c_682_n 0.00682312f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_M1018_g N_A_399_297#_c_682_n 0.00682312f $X=4.23 $Y=0.56 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_M1020_g N_A_399_297#_c_682_n 5.26907e-19 $X=4.75 $Y=0.56 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_217_n N_A_399_297#_c_686_n 7.3868e-19 $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_218_n N_A_399_297#_c_686_n 0.0125412f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_219_n N_A_399_297#_c_686_n 0.0125412f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_220_n N_A_399_297#_c_686_n 7.3868e-19 $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_M1018_g N_A_399_297#_c_690_n 6.99304e-19 $X=4.23 $Y=0.56 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_M1020_g N_A_399_297#_c_690_n 0.0064517f $X=4.75 $Y=0.56 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_M1021_g N_A_399_297#_c_690_n 0.00497927f $X=5.17 $Y=0.56 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_219_n N_A_399_297#_c_693_n 9.22981e-19 $X=4.255 $Y=1.41
+ $X2=0 $Y2=0
cc_285 N_A_27_47#_c_220_n N_A_399_297#_c_693_n 0.0122206f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_221_n N_A_399_297#_c_693_n 0.0105796f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_M1011_g N_A_399_297#_c_615_n 0.00109221f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_M1013_g N_A_399_297#_c_615_n 0.00109221f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_211_n N_A_399_297#_c_615_n 0.0236973f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_213_n N_A_399_297#_c_615_n 0.00213429f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_291 N_A_27_47#_c_216_n N_A_399_297#_c_623_n 0.0020332f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_217_n N_A_399_297#_c_623_n 0.0020332f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_211_n N_A_399_297#_c_623_n 0.0193444f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_213_n N_A_399_297#_c_623_n 0.00787799f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_295 N_A_27_47#_c_211_n N_A_399_297#_c_704_n 0.0420335f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_213_n N_A_399_297#_c_704_n 0.0171962f $X=5.17 $Y=1.217 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_211_n N_A_399_297#_c_624_n 0.00469235f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_213_n N_A_399_297#_c_624_n 0.00418132f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_299 N_A_27_47#_c_211_n N_A_399_297#_c_708_n 0.00129671f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_213_n N_A_399_297#_c_708_n 0.003124f $X=5.17 $Y=1.217 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_209_n N_A_399_297#_c_625_n 4.21355e-19 $X=1.507 $Y=1.075
+ $X2=0 $Y2=0
cc_302 N_A_27_47#_c_210_n N_A_399_297#_c_625_n 0.0022543f $X=1.507 $Y=1.445
+ $X2=0 $Y2=0
cc_303 N_A_27_47#_c_211_n N_A_399_297#_c_625_n 0.0182198f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_213_n N_A_399_297#_c_625_n 0.0163619f $X=5.17 $Y=1.217 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_214_n N_A_399_297#_c_616_n 0.00267651f $X=1.905 $Y=1.41
+ $X2=0 $Y2=0
cc_306 N_A_27_47#_M1004_g N_A_399_297#_c_616_n 0.00218385f $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_M1008_g N_A_399_297#_c_616_n 2.21948e-19 $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_215_n N_A_399_297#_c_616_n 0.00183898f $X=2.375 $Y=1.41
+ $X2=0 $Y2=0
cc_309 N_A_27_47#_c_216_n N_A_399_297#_c_616_n 0.00145847f $X=2.845 $Y=1.41
+ $X2=0 $Y2=0
cc_310 N_A_27_47#_M1011_g N_A_399_297#_c_616_n 7.21245e-19 $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_246_n N_A_399_297#_c_616_n 0.00232385f $X=1.2 $Y=1.63 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_209_n N_A_399_297#_c_616_n 0.00345304f $X=1.507 $Y=1.075
+ $X2=0 $Y2=0
cc_313 N_A_27_47#_c_210_n N_A_399_297#_c_616_n 0.00408613f $X=1.507 $Y=1.445
+ $X2=0 $Y2=0
cc_314 N_A_27_47#_c_211_n N_A_399_297#_c_616_n 0.00169102f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_226_n N_A_399_297#_c_616_n 0.00322698f $X=1.507 $Y=1.53
+ $X2=0 $Y2=0
cc_316 N_A_27_47#_c_212_n N_A_399_297#_c_616_n 0.0037465f $X=1.507 $Y=0.82 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_262_n N_A_399_297#_c_616_n 0.00187497f $X=1.507 $Y=1.16
+ $X2=0 $Y2=0
cc_318 N_A_27_47#_c_213_n N_A_399_297#_c_616_n 0.00183501f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_319 N_A_27_47#_M1006_d N_A_399_297#_c_617_n 3.41926e-19 $X=1.065 $Y=0.235
+ $X2=0 $Y2=0
cc_320 N_A_27_47#_M1009_d N_A_399_297#_c_617_n 3.42017e-19 $X=1.055 $Y=1.485
+ $X2=0 $Y2=0
cc_321 N_A_27_47#_M1004_g N_A_399_297#_c_617_n 3.17501e-19 $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_216_n N_A_399_297#_c_617_n 0.0110494f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_M1011_g N_A_399_297#_c_617_n 0.00402727f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_246_n N_A_399_297#_c_617_n 0.00653266f $X=1.2 $Y=1.63 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_311_p N_A_399_297#_c_617_n 0.00616563f $X=1.2 $Y=0.42 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_209_n N_A_399_297#_c_617_n 3.62077e-19 $X=1.507 $Y=1.075
+ $X2=0 $Y2=0
cc_327 N_A_27_47#_c_210_n N_A_399_297#_c_617_n 4.01269e-19 $X=1.507 $Y=1.445
+ $X2=0 $Y2=0
cc_328 N_A_27_47#_c_211_n N_A_399_297#_c_617_n 8.57141e-19 $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_226_n N_A_399_297#_c_617_n 0.00103827f $X=1.507 $Y=1.53
+ $X2=0 $Y2=0
cc_330 N_A_27_47#_c_212_n N_A_399_297#_c_617_n 0.00129991f $X=1.507 $Y=0.82
+ $X2=0 $Y2=0
cc_331 N_A_27_47#_c_262_n N_A_399_297#_c_617_n 2.28743e-19 $X=1.507 $Y=1.16
+ $X2=0 $Y2=0
cc_332 N_A_27_47#_c_213_n N_A_399_297#_c_617_n 0.00448615f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_333 N_A_27_47#_c_209_n N_A_399_297#_c_618_n 6.76651e-19 $X=1.507 $Y=1.075
+ $X2=0 $Y2=0
cc_334 N_A_27_47#_c_210_n N_A_399_297#_c_618_n 0.00149593f $X=1.507 $Y=1.445
+ $X2=0 $Y2=0
cc_335 N_A_27_47#_c_211_n N_A_399_297#_c_618_n 0.00389039f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_213_n N_A_399_297#_c_618_n 0.0177477f $X=5.17 $Y=1.217 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_218_n N_A_399_297#_c_619_n 0.0020332f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_M1016_g N_A_399_297#_c_619_n 0.00142075f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_M1018_g N_A_399_297#_c_619_n 0.0131543f $X=4.23 $Y=0.56 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_c_219_n N_A_399_297#_c_619_n 0.0151322f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_c_220_n N_A_399_297#_c_619_n 0.013508f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_M1020_g N_A_399_297#_c_619_n 0.01178f $X=4.75 $Y=0.56 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_M1021_g N_A_399_297#_c_619_n 0.00986498f $X=5.17 $Y=0.56 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_221_n N_A_399_297#_c_619_n 0.00677208f $X=5.195 $Y=1.41
+ $X2=0 $Y2=0
cc_345 N_A_27_47#_c_211_n N_A_399_297#_c_619_n 0.0322084f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_213_n N_A_399_297#_c_619_n 0.0848407f $X=5.17 $Y=1.217 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_209_n N_A_399_297#_c_629_n 4.98958e-19 $X=1.507 $Y=1.075
+ $X2=0 $Y2=0
cc_348 N_A_27_47#_c_210_n N_A_399_297#_c_629_n 0.00172251f $X=1.507 $Y=1.445
+ $X2=0 $Y2=0
cc_349 N_A_27_47#_c_211_n N_A_399_297#_c_629_n 0.00508713f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_213_n N_A_399_297#_c_629_n 0.0177329f $X=5.17 $Y=1.217 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_207_n N_VGND_M1002_s 0.00173798f $X=1.065 $Y=0.82 $X2=-1.26
+ $Y2=-1.17
cc_352 N_A_27_47#_c_212_n N_VGND_M1015_s 0.00228583f $X=1.507 $Y=0.82 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_430_p N_VGND_c_851_n 0.0128183f $X=0.31 $Y=0.42 $X2=0 $Y2=0
cc_354 N_A_27_47#_c_207_n N_VGND_c_851_n 0.0198831f $X=1.065 $Y=0.82 $X2=0 $Y2=0
cc_355 N_A_27_47#_c_311_p N_VGND_c_851_n 0.0126144f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_356 N_A_27_47#_M1004_g N_VGND_c_852_n 0.00224944f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_357 N_A_27_47#_c_311_p N_VGND_c_852_n 0.0191661f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_358 N_A_27_47#_c_211_n N_VGND_c_852_n 0.00749407f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_359 N_A_27_47#_c_212_n N_VGND_c_852_n 0.00585571f $X=1.507 $Y=0.82 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_M1004_g N_VGND_c_853_n 0.00541359f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_361 N_A_27_47#_M1008_g N_VGND_c_853_n 0.00424416f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_362 N_A_27_47#_M1008_g N_VGND_c_854_n 0.00222387f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_363 N_A_27_47#_M1011_g N_VGND_c_854_n 0.00222387f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_364 N_A_27_47#_M1011_g N_VGND_c_855_n 0.00424416f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_365 N_A_27_47#_M1013_g N_VGND_c_855_n 0.00424416f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_366 N_A_27_47#_M1013_g N_VGND_c_856_n 0.00166854f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_367 N_A_27_47#_M1016_g N_VGND_c_856_n 0.00166854f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_368 N_A_27_47#_M1016_g N_VGND_c_857_n 0.00424416f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_369 N_A_27_47#_M1018_g N_VGND_c_857_n 0.00472104f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_370 N_A_27_47#_M1018_g N_VGND_c_858_n 0.00166854f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_371 N_A_27_47#_M1020_g N_VGND_c_858_n 0.0022161f $X=4.75 $Y=0.56 $X2=0 $Y2=0
cc_372 N_A_27_47#_c_213_n N_VGND_c_858_n 7.95874e-19 $X=5.17 $Y=1.217 $X2=0
+ $Y2=0
cc_373 N_A_27_47#_M1021_g N_VGND_c_859_n 0.0037513f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_374 N_A_27_47#_M1020_g N_VGND_c_860_n 0.00472104f $X=4.75 $Y=0.56 $X2=0 $Y2=0
cc_375 N_A_27_47#_M1021_g N_VGND_c_860_n 0.00541359f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_376 N_A_27_47#_M1021_g N_VGND_c_862_n 0.00143885f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_377 N_A_27_47#_c_213_n N_VGND_c_862_n 4.85047e-19 $X=5.17 $Y=1.217 $X2=0
+ $Y2=0
cc_378 N_A_27_47#_M1020_g N_VGND_R2_neg 0.00102843f $X=4.75 $Y=0.56 $X2=0 $Y2=0
cc_379 N_A_27_47#_M1021_g N_VGND_R2_neg 7.29361e-19 $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_380 N_A_27_47#_c_213_n N_VGND_R2_neg 4.34579e-19 $X=5.17 $Y=1.217 $X2=0 $Y2=0
cc_381 N_A_27_47#_c_207_n N_VGND_c_864_n 0.00610276f $X=1.065 $Y=0.82 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_c_311_p N_VGND_c_864_n 0.0170101f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_383 N_A_27_47#_c_430_p N_VGND_c_866_n 0.0189483f $X=0.31 $Y=0.42 $X2=0 $Y2=0
cc_384 N_A_27_47#_c_207_n N_VGND_c_866_n 0.00304253f $X=1.065 $Y=0.82 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_M1002_d N_VGND_c_872_n 0.00276728f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_M1006_d N_VGND_c_872_n 0.00624525f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_M1004_g N_VGND_c_872_n 0.009238f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_388 N_A_27_47#_M1008_g N_VGND_c_872_n 0.00919137f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_389 N_A_27_47#_M1011_g N_VGND_c_872_n 0.00597838f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_390 N_A_27_47#_M1013_g N_VGND_c_872_n 0.00597838f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_391 N_A_27_47#_M1016_g N_VGND_c_872_n 0.00597838f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_392 N_A_27_47#_M1018_g N_VGND_c_872_n 0.0075548f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_393 N_A_27_47#_M1020_g N_VGND_c_872_n 0.00922694f $X=4.75 $Y=0.56 $X2=0 $Y2=0
cc_394 N_A_27_47#_M1021_g N_VGND_c_872_n 0.00982257f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_395 N_A_27_47#_c_430_p N_VGND_c_872_n 0.0114629f $X=0.31 $Y=0.42 $X2=0 $Y2=0
cc_396 N_A_27_47#_c_207_n N_VGND_c_872_n 0.0118592f $X=1.065 $Y=0.82 $X2=0 $Y2=0
cc_397 N_A_27_47#_c_311_p N_VGND_c_872_n 0.0100577f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_398 N_A_27_47#_c_212_n N_VGND_c_872_n 0.00110273f $X=1.507 $Y=0.82 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_c_222_n N_X_c_991_n 0.00401157f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_400 N_A_27_47#_c_224_n N_X_c_991_n 0.00228854f $X=0.425 $Y=1.53 $X2=0 $Y2=0
cc_401 N_A_27_47#_c_208_n N_X_c_991_n 0.00178675f $X=0.445 $Y=0.82 $X2=0 $Y2=0
cc_402 N_A_27_47#_M1002_d N_X_R0_pos 2.2489e-19 $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_403 N_A_27_47#_c_222_n N_X_R0_pos 0.00960102f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_404 N_A_27_47#_c_430_p N_X_R0_pos 0.00544849f $X=0.31 $Y=0.42 $X2=0 $Y2=0
cc_405 N_A_27_47#_c_223_n N_X_R0_pos 0.00217275f $X=1.035 $Y=1.53 $X2=0 $Y2=0
cc_406 N_A_27_47#_c_224_n N_X_R0_pos 0.00211659f $X=0.425 $Y=1.53 $X2=0 $Y2=0
cc_407 N_A_27_47#_c_207_n N_X_R0_pos 0.0013315f $X=1.065 $Y=0.82 $X2=0 $Y2=0
cc_408 N_A_27_47#_c_208_n N_X_R0_pos 0.00158492f $X=0.445 $Y=0.82 $X2=0 $Y2=0
cc_409 N_A_27_47#_c_246_n N_X_R0_pos 0.00129226f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_410 N_VPWR_c_489_n N_A_399_297#_M1000_d 0.00915074f $X=5.68 $Y=2.72 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_489_n N_A_399_297#_M1005_d 0.00232867f $X=5.68 $Y=2.72 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_489_n N_A_399_297#_M1010_d 0.00232867f $X=5.68 $Y=2.72 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_489_n N_A_399_297#_M1014_d 0.00857341f $X=5.68 $Y=2.72 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_492_n N_A_399_297#_c_631_n 0.0368524f $X=1.67 $Y=2 $X2=0 $Y2=0
cc_415 N_VPWR_c_493_n N_A_399_297#_c_631_n 0.0235906f $X=2.475 $Y=2.72 $X2=0
+ $Y2=0
cc_416 N_VPWR_c_494_n N_A_399_297#_c_631_n 0.0368524f $X=2.61 $Y=2 $X2=0 $Y2=0
cc_417 N_VPWR_c_489_n N_A_399_297#_c_631_n 0.0121187f $X=5.68 $Y=2.72 $X2=0
+ $Y2=0
cc_418 N_VPWR_M1003_s N_A_399_297#_c_620_n 0.00160554f $X=2.465 $Y=1.485 $X2=0
+ $Y2=0
cc_419 N_VPWR_c_494_n N_A_399_297#_c_620_n 0.0149424f $X=2.61 $Y=2 $X2=0 $Y2=0
cc_420 N_VPWR_c_494_n N_A_399_297#_c_670_n 0.0365704f $X=2.61 $Y=2 $X2=0 $Y2=0
cc_421 N_VPWR_c_495_n N_A_399_297#_c_670_n 0.0190121f $X=3.415 $Y=2.72 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_489_n N_A_399_297#_c_670_n 0.0124581f $X=5.68 $Y=2.72 $X2=0
+ $Y2=0
cc_423 N_VPWR_M1007_s N_A_399_297#_c_622_n 0.00209407f $X=3.405 $Y=1.485 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_496_n N_A_399_297#_c_622_n 0.011151f $X=3.55 $Y=2 $X2=0 $Y2=0
cc_425 N_VPWR_c_497_n N_A_399_297#_c_686_n 0.0190121f $X=4.355 $Y=2.72 $X2=0
+ $Y2=0
cc_426 N_VPWR_R1_neg N_A_399_297#_c_686_n 7.9666e-19 $X=4.46 $Y=2.875 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_489_n N_A_399_297#_c_686_n 0.0124581f $X=5.68 $Y=2.72 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_498_n N_A_399_297#_c_693_n 0.0300298f $X=4.49 $Y=2 $X2=0 $Y2=0
cc_429 N_VPWR_c_499_n N_A_399_297#_c_693_n 0.0383253f $X=5.43 $Y=1.66 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_500_n N_A_399_297#_c_693_n 0.0235011f $X=5.295 $Y=2.72 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_487_n N_A_399_297#_c_693_n 0.0033778f $X=5.72 $Y=2.72 $X2=0
+ $Y2=0
cc_432 N_VPWR_R1_neg N_A_399_297#_c_693_n 0.00358352f $X=4.46 $Y=2.875 $X2=0
+ $Y2=0
cc_433 N_VPWR_c_489_n N_A_399_297#_c_693_n 0.0119808f $X=5.68 $Y=2.72 $X2=0
+ $Y2=0
cc_434 N_VPWR_c_498_n N_A_399_297#_c_708_n 0.00125393f $X=4.49 $Y=2 $X2=0 $Y2=0
cc_435 N_VPWR_R1_neg N_A_399_297#_c_785_n 0.00478002f $X=4.46 $Y=2.875 $X2=0
+ $Y2=0
cc_436 N_VPWR_M1003_s N_A_399_297#_c_616_n 0.00258481f $X=2.465 $Y=1.485 $X2=0
+ $Y2=0
cc_437 N_VPWR_c_492_n N_A_399_297#_c_616_n 0.00443932f $X=1.67 $Y=2 $X2=0 $Y2=0
cc_438 N_VPWR_c_494_n N_A_399_297#_c_616_n 0.00387397f $X=2.61 $Y=2 $X2=0 $Y2=0
cc_439 N_VPWR_c_489_n N_A_399_297#_c_616_n 0.0160911f $X=5.68 $Y=2.72 $X2=0
+ $Y2=0
cc_440 N_VPWR_c_490_n N_A_399_297#_c_617_n 0.00113136f $X=0.73 $Y=2 $X2=0 $Y2=0
cc_441 N_VPWR_c_492_n N_A_399_297#_c_617_n 0.00178229f $X=1.67 $Y=2 $X2=0 $Y2=0
cc_442 N_VPWR_c_494_n N_A_399_297#_c_617_n 0.00109478f $X=2.61 $Y=2 $X2=0 $Y2=0
cc_443 N_VPWR_c_496_n N_A_399_297#_c_617_n 3.2535e-19 $X=3.55 $Y=2 $X2=0 $Y2=0
cc_444 N_VPWR_R1_neg N_A_399_297#_c_617_n 0.102261f $X=4.46 $Y=2.875 $X2=0 $Y2=0
cc_445 N_VPWR_c_489_n N_A_399_297#_c_617_n 0.0541286f $X=5.68 $Y=2.72 $X2=0
+ $Y2=0
cc_446 N_VPWR_M1012_s N_A_399_297#_c_619_n 0.00218233f $X=4.345 $Y=1.485 $X2=0
+ $Y2=0
cc_447 N_VPWR_c_498_n N_A_399_297#_c_619_n 0.0123277f $X=4.49 $Y=2 $X2=0 $Y2=0
cc_448 N_VPWR_R1_neg N_A_399_297#_c_619_n 0.00173316f $X=4.46 $Y=2.875 $X2=0
+ $Y2=0
cc_449 N_VPWR_c_499_n N_VGND_c_859_n 0.00779664f $X=5.43 $Y=1.66 $X2=0 $Y2=0
cc_450 N_VPWR_R1_neg N_VGND_c_859_n 5.56789e-19 $X=4.46 $Y=2.875 $X2=0 $Y2=0
cc_451 N_VPWR_R1_neg N_VGND_c_862_n 0.0179445f $X=4.46 $Y=2.875 $X2=0 $Y2=0
cc_452 N_VPWR_c_499_n N_VGND_R2_neg 0.00121042f $X=5.43 $Y=1.66 $X2=0 $Y2=0
cc_453 N_VPWR_c_487_n N_VGND_R2_neg 0.0189015f $X=5.72 $Y=2.72 $X2=0 $Y2=0
cc_454 N_VPWR_R1_neg N_VGND_R2_neg 0.171054f $X=4.46 $Y=2.875 $X2=0 $Y2=0
cc_455 N_VPWR_c_489_n N_X_c_991_n 8.18796e-19 $X=5.68 $Y=2.72 $X2=0 $Y2=0
cc_456 N_VPWR_M1001_s N_X_R0_pos 3.27113e-19 $X=0.585 $Y=1.485 $X2=0 $Y2=0
cc_457 N_VPWR_c_490_n N_X_R0_pos 0.00561607f $X=0.73 $Y=2 $X2=0 $Y2=0
cc_458 N_VPWR_c_489_n N_X_R0_pos 0.0193072f $X=5.68 $Y=2.72 $X2=0 $Y2=0
cc_459 N_A_399_297#_c_616_n N_VGND_M1015_s 0.00293625f $X=2.05 $Y=1.36 $X2=0
+ $Y2=0
cc_460 N_A_399_297#_c_612_n N_VGND_M1008_d 0.00224229f $X=2.915 $Y=0.82 $X2=0
+ $Y2=0
cc_461 N_A_399_297#_c_617_n N_VGND_M1008_d 0.00679232f $X=2.05 $Y=1.36 $X2=0
+ $Y2=0
cc_462 N_A_399_297#_c_614_n N_VGND_M1013_d 0.00274103f $X=3.855 $Y=0.82 $X2=0
+ $Y2=0
cc_463 N_A_399_297#_c_619_n N_VGND_M1018_d 0.00282836f $X=4.96 $Y=1.175 $X2=0
+ $Y2=0
cc_464 N_A_399_297#_c_617_n N_VGND_c_851_n 0.00114248f $X=2.05 $Y=1.36 $X2=0
+ $Y2=0
cc_465 N_A_399_297#_c_630_n N_VGND_c_852_n 0.0182045f $X=2.14 $Y=0.42 $X2=0
+ $Y2=0
cc_466 N_A_399_297#_c_616_n N_VGND_c_852_n 0.00236269f $X=2.05 $Y=1.36 $X2=0
+ $Y2=0
cc_467 N_A_399_297#_c_617_n N_VGND_c_852_n 0.00178914f $X=2.05 $Y=1.36 $X2=0
+ $Y2=0
cc_468 N_A_399_297#_c_630_n N_VGND_c_853_n 0.023531f $X=2.14 $Y=0.42 $X2=0 $Y2=0
cc_469 N_A_399_297#_c_612_n N_VGND_c_853_n 0.00293546f $X=2.915 $Y=0.82 $X2=0
+ $Y2=0
cc_470 N_A_399_297#_c_630_n N_VGND_c_854_n 0.0181274f $X=2.14 $Y=0.42 $X2=0
+ $Y2=0
cc_471 N_A_399_297#_c_612_n N_VGND_c_854_n 0.0214278f $X=2.915 $Y=0.82 $X2=0
+ $Y2=0
cc_472 N_A_399_297#_c_666_n N_VGND_c_854_n 0.0179949f $X=3.08 $Y=0.42 $X2=0
+ $Y2=0
cc_473 N_A_399_297#_c_616_n N_VGND_c_854_n 9.3276e-19 $X=2.05 $Y=1.36 $X2=0
+ $Y2=0
cc_474 N_A_399_297#_c_617_n N_VGND_c_854_n 9.6831e-19 $X=2.05 $Y=1.36 $X2=0
+ $Y2=0
cc_475 N_A_399_297#_c_612_n N_VGND_c_855_n 0.00204707f $X=2.915 $Y=0.82 $X2=0
+ $Y2=0
cc_476 N_A_399_297#_c_666_n N_VGND_c_855_n 0.0188551f $X=3.08 $Y=0.42 $X2=0
+ $Y2=0
cc_477 N_A_399_297#_c_614_n N_VGND_c_855_n 0.00193763f $X=3.855 $Y=0.82 $X2=0
+ $Y2=0
cc_478 N_A_399_297#_c_614_n N_VGND_c_856_n 0.019437f $X=3.855 $Y=0.82 $X2=0
+ $Y2=0
cc_479 N_A_399_297#_c_617_n N_VGND_c_856_n 2.15012e-19 $X=2.05 $Y=1.36 $X2=0
+ $Y2=0
cc_480 N_A_399_297#_c_614_n N_VGND_c_857_n 0.00193763f $X=3.855 $Y=0.82 $X2=0
+ $Y2=0
cc_481 N_A_399_297#_c_682_n N_VGND_c_857_n 0.0188551f $X=4.02 $Y=0.42 $X2=0
+ $Y2=0
cc_482 N_A_399_297#_c_619_n N_VGND_c_857_n 0.00132422f $X=4.96 $Y=1.175 $X2=0
+ $Y2=0
cc_483 N_A_399_297#_c_690_n N_VGND_c_858_n 0.0180226f $X=4.96 $Y=0.42 $X2=0
+ $Y2=0
cc_484 N_A_399_297#_c_708_n N_VGND_c_858_n 0.00113435f $X=4.36 $Y=1.19 $X2=0
+ $Y2=0
cc_485 N_A_399_297#_c_619_n N_VGND_c_858_n 0.0214341f $X=4.96 $Y=1.175 $X2=0
+ $Y2=0
cc_486 N_A_399_297#_c_690_n N_VGND_c_859_n 0.0243132f $X=4.96 $Y=0.42 $X2=0
+ $Y2=0
cc_487 N_A_399_297#_c_690_n N_VGND_c_860_n 0.0235017f $X=4.96 $Y=0.42 $X2=0
+ $Y2=0
cc_488 N_A_399_297#_c_619_n N_VGND_c_860_n 0.0013974f $X=4.96 $Y=1.175 $X2=0
+ $Y2=0
cc_489 N_A_399_297#_c_690_n N_VGND_c_862_n 0.00337185f $X=4.96 $Y=0.42 $X2=0
+ $Y2=0
cc_490 N_A_399_297#_c_682_n N_VGND_R2_neg 7.9666e-19 $X=4.02 $Y=0.42 $X2=0 $Y2=0
cc_491 N_A_399_297#_c_690_n N_VGND_R2_neg 0.00359563f $X=4.96 $Y=0.42 $X2=0
+ $Y2=0
cc_492 N_A_399_297#_c_785_n N_VGND_R2_neg 0.00540571f $X=4.75 $Y=1.19 $X2=0
+ $Y2=0
cc_493 N_A_399_297#_c_617_n N_VGND_R2_neg 0.102322f $X=2.05 $Y=1.36 $X2=0 $Y2=0
cc_494 N_A_399_297#_c_619_n N_VGND_R2_neg 0.00168535f $X=4.96 $Y=1.175 $X2=0
+ $Y2=0
cc_495 N_A_399_297#_M1004_s N_VGND_c_872_n 0.00845654f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_496 N_A_399_297#_M1011_s N_VGND_c_872_n 0.00215201f $X=2.945 $Y=0.235 $X2=0
+ $Y2=0
cc_497 N_A_399_297#_M1016_s N_VGND_c_872_n 0.00215201f $X=3.885 $Y=0.235 $X2=0
+ $Y2=0
cc_498 N_A_399_297#_M1020_s N_VGND_c_872_n 0.00791551f $X=4.825 $Y=0.235 $X2=0
+ $Y2=0
cc_499 N_A_399_297#_c_630_n N_VGND_c_872_n 0.012028f $X=2.14 $Y=0.42 $X2=0 $Y2=0
cc_500 N_A_399_297#_c_612_n N_VGND_c_872_n 0.0108312f $X=2.915 $Y=0.82 $X2=0
+ $Y2=0
cc_501 N_A_399_297#_c_666_n N_VGND_c_872_n 0.0122069f $X=3.08 $Y=0.42 $X2=0
+ $Y2=0
cc_502 N_A_399_297#_c_614_n N_VGND_c_872_n 0.00863183f $X=3.855 $Y=0.82 $X2=0
+ $Y2=0
cc_503 N_A_399_297#_c_682_n N_VGND_c_872_n 0.0122069f $X=4.02 $Y=0.42 $X2=0
+ $Y2=0
cc_504 N_A_399_297#_c_690_n N_VGND_c_872_n 0.0119036f $X=4.96 $Y=0.42 $X2=0
+ $Y2=0
cc_505 N_A_399_297#_c_616_n N_VGND_c_872_n 0.0162979f $X=2.05 $Y=1.36 $X2=0
+ $Y2=0
cc_506 N_A_399_297#_c_617_n N_VGND_c_872_n 0.0541321f $X=2.05 $Y=1.36 $X2=0
+ $Y2=0
cc_507 N_A_399_297#_c_618_n N_VGND_c_872_n 0.0161149f $X=2.475 $Y=1.19 $X2=0
+ $Y2=0
cc_508 N_A_399_297#_c_619_n N_VGND_c_872_n 0.00924895f $X=4.96 $Y=1.175 $X2=0
+ $Y2=0
cc_509 N_A_399_297#_c_617_n M5_872_N71# 0.00673347f $X=2.05 $Y=1.36 $X2=-1.26
+ $Y2=-1.17
cc_510 N_A_399_297#_c_617_n M5_872_595# 0.00673347f $X=2.05 $Y=1.36 $X2=-1.26
+ $Y2=-1.17
cc_511 N_VGND_c_872_n N_X_c_991_n 8.18796e-19 $X=5.68 $Y=0 $X2=0 $Y2=0
cc_512 N_VGND_c_872_n N_X_c_992_n 0.00174134f $X=5.68 $Y=0 $X2=0 $Y2=0
cc_513 N_VGND_M1002_s N_X_R0_pos 7.36004e-19 $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_514 N_VGND_c_851_n N_X_R0_pos 0.0046429f $X=0.76 $Y=0.4 $X2=0 $Y2=0
cc_515 N_VGND_c_872_n N_X_R0_pos 0.0194743f $X=5.68 $Y=0 $X2=0 $Y2=0
