* File: sky130_fd_sc_hdll__o31ai_2.pxi.spice
* Created: Wed Sep  2 08:46:51 2020
* 
x_PM_SKY130_FD_SC_HDLL__O31AI_2%A1 N_A1_c_75_n N_A1_M1000_g N_A1_M1004_g
+ N_A1_c_76_n N_A1_M1013_g N_A1_M1015_g A1 A1 A1 N_A1_c_74_n A1 A1
+ PM_SKY130_FD_SC_HDLL__O31AI_2%A1
x_PM_SKY130_FD_SC_HDLL__O31AI_2%A2 N_A2_M1011_g N_A2_c_123_n N_A2_M1006_g
+ N_A2_c_124_n N_A2_M1009_g N_A2_M1014_g A2 A2 N_A2_c_121_n A2 A2
+ PM_SKY130_FD_SC_HDLL__O31AI_2%A2
x_PM_SKY130_FD_SC_HDLL__O31AI_2%A3 N_A3_M1002_g N_A3_c_171_n N_A3_M1005_g
+ N_A3_c_172_n N_A3_M1012_g N_A3_M1003_g A3 A3 N_A3_c_170_n
+ PM_SKY130_FD_SC_HDLL__O31AI_2%A3
x_PM_SKY130_FD_SC_HDLL__O31AI_2%B1 N_B1_c_222_n N_B1_M1007_g N_B1_c_228_n
+ N_B1_M1001_g N_B1_c_223_n N_B1_c_224_n N_B1_M1008_g N_B1_c_230_n N_B1_M1010_g
+ N_B1_c_225_n B1 B1 N_B1_c_227_n PM_SKY130_FD_SC_HDLL__O31AI_2%B1
x_PM_SKY130_FD_SC_HDLL__O31AI_2%A_27_297# N_A_27_297#_M1000_s
+ N_A_27_297#_M1013_s N_A_27_297#_M1009_d N_A_27_297#_c_275_n
+ N_A_27_297#_c_281_n N_A_27_297#_c_276_n N_A_27_297#_c_288_n
+ N_A_27_297#_c_277_n N_A_27_297#_c_278_n N_A_27_297#_c_290_n
+ PM_SKY130_FD_SC_HDLL__O31AI_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__O31AI_2%VPWR N_VPWR_M1000_d N_VPWR_M1001_d
+ N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_327_n N_VPWR_c_328_n VPWR
+ N_VPWR_c_329_n N_VPWR_c_324_n N_VPWR_c_331_n VPWR
+ PM_SKY130_FD_SC_HDLL__O31AI_2%VPWR
x_PM_SKY130_FD_SC_HDLL__O31AI_2%A_309_297# N_A_309_297#_M1006_s
+ N_A_309_297#_M1005_s N_A_309_297#_c_381_n N_A_309_297#_c_380_n
+ N_A_309_297#_c_384_n N_A_309_297#_c_387_n
+ PM_SKY130_FD_SC_HDLL__O31AI_2%A_309_297#
x_PM_SKY130_FD_SC_HDLL__O31AI_2%Y N_Y_M1007_d N_Y_M1005_d N_Y_M1012_d
+ N_Y_M1010_s N_Y_c_417_n N_Y_c_412_n N_Y_c_424_n N_Y_c_435_n N_Y_c_426_n Y Y Y
+ Y Y Y N_Y_c_413_n N_Y_c_411_n N_Y_c_415_n N_Y_c_416_n
+ PM_SKY130_FD_SC_HDLL__O31AI_2%Y
x_PM_SKY130_FD_SC_HDLL__O31AI_2%A_27_47# N_A_27_47#_M1004_s N_A_27_47#_M1015_s
+ N_A_27_47#_M1014_d N_A_27_47#_M1003_d N_A_27_47#_M1008_s N_A_27_47#_c_477_n
+ N_A_27_47#_c_483_n N_A_27_47#_c_478_n N_A_27_47#_c_489_n N_A_27_47#_c_494_n
+ N_A_27_47#_c_531_p N_A_27_47#_c_479_n N_A_27_47#_c_503_n N_A_27_47#_c_504_n
+ N_A_27_47#_c_480_n N_A_27_47#_c_481_n N_A_27_47#_c_482_n
+ PM_SKY130_FD_SC_HDLL__O31AI_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__O31AI_2%VGND N_VGND_M1004_d N_VGND_M1011_s
+ N_VGND_M1002_s N_VGND_c_559_n N_VGND_c_560_n N_VGND_c_561_n VGND
+ N_VGND_c_562_n N_VGND_c_563_n N_VGND_c_564_n N_VGND_c_565_n N_VGND_c_566_n
+ N_VGND_c_567_n VGND PM_SKY130_FD_SC_HDLL__O31AI_2%VGND
cc_1 VNB N_A1_M1004_g 0.0248455f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.56
cc_2 VNB N_A1_M1015_g 0.0182928f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.56
cc_3 VNB A1 0.0166335f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=1.105
cc_4 VNB N_A1_c_74_n 0.0528215f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.217
cc_5 VNB N_A2_M1011_g 0.0245973f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.985
cc_6 VNB N_A2_M1014_g 0.0255794f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.56
cc_7 VNB N_A2_c_121_n 0.0742763f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.217
cc_8 VNB A2 0.00206023f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_9 VNB N_A3_M1002_g 0.0204905f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.985
cc_10 VNB N_A3_M1003_g 0.0196695f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.56
cc_11 VNB A3 0.00515346f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_12 VNB N_A3_c_170_n 0.049004f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.16
cc_13 VNB N_B1_c_222_n 0.0176338f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_14 VNB N_B1_c_223_n 0.0202368f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B1_c_224_n 0.0201269f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.985
cc_16 VNB N_B1_c_225_n 0.0126284f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_17 VNB B1 0.02223f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=1.105
cc_18 VNB N_B1_c_227_n 0.0374611f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.217
cc_19 VNB N_VPWR_c_324_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.19
cc_20 VNB N_Y_c_411_n 0.00112014f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_477_n 0.0183269f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_478_n 0.00987047f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.217
cc_23 VNB N_A_27_47#_c_479_n 0.00257058f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_480_n 0.0145744f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_25 VNB N_A_27_47#_c_481_n 0.001463f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.19
cc_26 VNB N_A_27_47#_c_482_n 0.00671718f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.19
cc_27 VNB N_VGND_c_559_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_560_n 0.0183417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_561_n 0.00315697f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_30 VNB N_VGND_c_562_n 0.0429072f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.19
cc_31 VNB N_VGND_c_563_n 0.257625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_564_n 0.022381f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_33 VNB N_VGND_c_565_n 0.0191455f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.19
cc_34 VNB N_VGND_c_566_n 0.0177312f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_567_n 0.00615226f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VPB N_A1_c_75_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_37 VPB N_A1_c_76_n 0.016445f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_38 VPB A1 0.00852148f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=1.105
cc_39 VPB N_A1_c_74_n 0.015459f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.217
cc_40 VPB N_A2_c_123_n 0.016445f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.56
cc_41 VPB N_A2_c_124_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_42 VPB N_A2_c_121_n 0.0155512f $X=-0.19 $Y=1.305 $X2=0.87 $Y2=1.217
cc_43 VPB A2 0.00888956f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.19
cc_44 VPB N_A3_c_171_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.56
cc_45 VPB N_A3_c_172_n 0.0164422f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_46 VPB A3 0.00457426f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_47 VPB N_A3_c_170_n 0.0154372f $X=-0.19 $Y=1.305 $X2=0.87 $Y2=1.16
cc_48 VPB N_B1_c_228_n 0.0172936f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.025
cc_49 VPB N_B1_c_223_n 0.0117687f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_B1_c_230_n 0.0216315f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.56
cc_51 VPB N_B1_c_225_n 0.00650317f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_52 VPB B1 0.00386571f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=1.105
cc_53 VPB N_B1_c_227_n 0.018977f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.217
cc_54 VPB N_A_27_297#_c_275_n 0.0316657f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.56
cc_55 VPB N_A_27_297#_c_276_n 0.00762919f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=1.105
cc_56 VPB N_A_27_297#_c_277_n 0.00198007f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.217
cc_57 VPB N_A_27_297#_c_278_n 0.0049682f $X=-0.19 $Y=1.305 $X2=0.87 $Y2=1.16
cc_58 VPB N_VPWR_c_325_n 0.00469739f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.025
cc_59 VPB N_VPWR_c_326_n 0.00562936f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_60 VPB N_VPWR_c_327_n 0.0791518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_328_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_329_n 0.0198069f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.217
cc_63 VPB N_VPWR_c_324_n 0.0477359f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.19
cc_64 VPB N_VPWR_c_331_n 0.0230861f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.19
cc_65 VPB N_A_309_297#_c_380_n 0.0137998f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.025
cc_66 VPB N_Y_c_412_n 0.00192487f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_Y_c_413_n 0.00445247f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.19
cc_68 VPB N_Y_c_411_n 0.00160381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_Y_c_415_n 0.00822879f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_Y_c_416_n 0.0334076f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 N_A1_M1015_g N_A2_M1011_g 0.0166832f $X=1.01 $Y=0.56 $X2=0 $Y2=0
cc_72 N_A1_c_76_n N_A2_c_123_n 0.0100726f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_73 A1 N_A2_c_121_n 0.00271895f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A1_c_74_n N_A2_c_121_n 0.0166832f $X=0.985 $Y=1.217 $X2=0 $Y2=0
cc_75 A1 A2 0.0219547f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_76 N_A1_c_75_n N_A_27_297#_c_275_n 0.0106251f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A1_c_76_n N_A_27_297#_c_275_n 6.25229e-19 $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A1_c_75_n N_A_27_297#_c_281_n 0.0137916f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_79 N_A1_c_76_n N_A_27_297#_c_281_n 0.0101048f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_80 A1 N_A_27_297#_c_281_n 0.0369312f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_81 N_A1_c_74_n N_A_27_297#_c_281_n 0.00154877f $X=0.985 $Y=1.217 $X2=0 $Y2=0
cc_82 N_A1_c_75_n N_A_27_297#_c_276_n 5.79575e-19 $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_83 A1 N_A_27_297#_c_276_n 0.0276353f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_84 N_A1_c_74_n N_A_27_297#_c_276_n 5.97581e-19 $X=0.985 $Y=1.217 $X2=0 $Y2=0
cc_85 N_A1_c_75_n N_A_27_297#_c_288_n 6.48386e-19 $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A1_c_76_n N_A_27_297#_c_288_n 0.0130707f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A1_c_76_n N_A_27_297#_c_290_n 0.00210477f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_88 A1 N_A_27_297#_c_290_n 0.0228561f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_89 N_A1_c_75_n N_VPWR_c_325_n 0.0052072f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A1_c_76_n N_VPWR_c_325_n 0.004751f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_91 N_A1_c_76_n N_VPWR_c_327_n 0.00597712f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A1_c_75_n N_VPWR_c_324_n 0.0127734f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_93 N_A1_c_76_n N_VPWR_c_324_n 0.0100198f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A1_c_75_n N_VPWR_c_331_n 0.00673617f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A1_M1004_g N_A_27_47#_c_483_n 0.0103753f $X=0.54 $Y=0.56 $X2=0 $Y2=0
cc_96 N_A1_M1015_g N_A_27_47#_c_483_n 0.00600753f $X=1.01 $Y=0.56 $X2=0 $Y2=0
cc_97 A1 N_A_27_47#_c_483_n 0.0352454f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_98 N_A1_c_74_n N_A_27_47#_c_483_n 0.00312059f $X=0.985 $Y=1.217 $X2=0 $Y2=0
cc_99 A1 N_A_27_47#_c_478_n 0.0280687f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_100 N_A1_c_74_n N_A_27_47#_c_478_n 0.00300662f $X=0.985 $Y=1.217 $X2=0 $Y2=0
cc_101 N_A1_M1004_g N_A_27_47#_c_489_n 5.79378e-19 $X=0.54 $Y=0.56 $X2=0 $Y2=0
cc_102 N_A1_M1015_g N_A_27_47#_c_489_n 0.00837042f $X=1.01 $Y=0.56 $X2=0 $Y2=0
cc_103 N_A1_M1015_g N_A_27_47#_c_481_n 0.00239159f $X=1.01 $Y=0.56 $X2=0 $Y2=0
cc_104 A1 N_A_27_47#_c_481_n 0.0222628f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_105 N_A1_M1004_g N_VGND_c_559_n 0.00276126f $X=0.54 $Y=0.56 $X2=0 $Y2=0
cc_106 N_A1_M1015_g N_VGND_c_559_n 0.0035663f $X=1.01 $Y=0.56 $X2=0 $Y2=0
cc_107 N_A1_M1004_g N_VGND_c_563_n 0.00700405f $X=0.54 $Y=0.56 $X2=0 $Y2=0
cc_108 N_A1_M1015_g N_VGND_c_563_n 0.00570363f $X=1.01 $Y=0.56 $X2=0 $Y2=0
cc_109 N_A1_M1004_g N_VGND_c_564_n 0.00436487f $X=0.54 $Y=0.56 $X2=0 $Y2=0
cc_110 N_A1_M1015_g N_VGND_c_565_n 0.00395968f $X=1.01 $Y=0.56 $X2=0 $Y2=0
cc_111 N_A2_M1014_g N_A3_M1002_g 0.00965467f $X=2.34 $Y=0.56 $X2=0 $Y2=0
cc_112 N_A2_c_121_n A3 0.00121686f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_113 A2 A3 0.0176873f $X=2.075 $Y=1.19 $X2=0 $Y2=0
cc_114 N_A2_c_121_n N_A3_c_170_n 0.00965467f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_115 A2 N_A3_c_170_n 0.00109651f $X=2.075 $Y=1.19 $X2=0 $Y2=0
cc_116 N_A2_c_123_n N_A_27_297#_c_288_n 0.0106013f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A2_c_124_n N_A_27_297#_c_288_n 7.44247e-19 $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A2_c_123_n N_A_27_297#_c_277_n 0.0153694f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A2_c_124_n N_A_27_297#_c_277_n 0.0104217f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A2_c_121_n N_A_27_297#_c_277_n 0.00358321f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_121 A2 N_A_27_297#_c_277_n 0.0581455f $X=2.075 $Y=1.19 $X2=0 $Y2=0
cc_122 N_A2_c_123_n N_A_27_297#_c_278_n 6.21613e-19 $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A2_c_124_n N_A_27_297#_c_278_n 0.00870676f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A2_c_123_n N_A_27_297#_c_290_n 8.61029e-19 $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A2_c_123_n N_VPWR_c_327_n 0.00673617f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A2_c_124_n N_VPWR_c_327_n 0.00429453f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A2_c_123_n N_VPWR_c_324_n 0.0120446f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A2_c_124_n N_VPWR_c_324_n 0.00743756f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A2_c_123_n N_A_309_297#_c_381_n 0.00206455f $X=1.455 $Y=1.41 $X2=0
+ $Y2=0
cc_130 N_A2_c_124_n N_A_309_297#_c_381_n 0.0045713f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A2_c_124_n N_A_309_297#_c_380_n 0.0137146f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A2_c_123_n N_A_309_297#_c_384_n 0.00142717f $X=1.455 $Y=1.41 $X2=0
+ $Y2=0
cc_133 N_A2_M1011_g N_A_27_47#_c_489_n 0.0113393f $X=1.43 $Y=0.56 $X2=0 $Y2=0
cc_134 N_A2_M1011_g N_A_27_47#_c_494_n 0.012122f $X=1.43 $Y=0.56 $X2=0 $Y2=0
cc_135 N_A2_M1014_g N_A_27_47#_c_494_n 0.0121821f $X=2.34 $Y=0.56 $X2=0 $Y2=0
cc_136 N_A2_c_121_n N_A_27_47#_c_494_n 0.0138627f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_137 A2 N_A_27_47#_c_494_n 0.062174f $X=2.075 $Y=1.19 $X2=0 $Y2=0
cc_138 N_A2_M1011_g N_A_27_47#_c_481_n 0.00124405f $X=1.43 $Y=0.56 $X2=0 $Y2=0
cc_139 N_A2_M1014_g N_VGND_c_560_n 0.00436487f $X=2.34 $Y=0.56 $X2=0 $Y2=0
cc_140 N_A2_M1014_g N_VGND_c_561_n 9.94141e-19 $X=2.34 $Y=0.56 $X2=0 $Y2=0
cc_141 N_A2_M1011_g N_VGND_c_563_n 0.0071726f $X=1.43 $Y=0.56 $X2=0 $Y2=0
cc_142 N_A2_M1014_g N_VGND_c_563_n 0.00765965f $X=2.34 $Y=0.56 $X2=0 $Y2=0
cc_143 N_A2_M1011_g N_VGND_c_565_n 0.00422241f $X=1.43 $Y=0.56 $X2=0 $Y2=0
cc_144 N_A2_M1011_g N_VGND_c_566_n 0.00598627f $X=1.43 $Y=0.56 $X2=0 $Y2=0
cc_145 N_A2_M1014_g N_VGND_c_566_n 0.0118078f $X=2.34 $Y=0.56 $X2=0 $Y2=0
cc_146 N_A3_M1003_g N_B1_c_222_n 0.0165726f $X=3.48 $Y=0.56 $X2=-0.19 $Y2=-0.24
cc_147 N_A3_c_172_n N_B1_c_228_n 0.00975452f $X=3.455 $Y=1.41 $X2=0 $Y2=0
cc_148 A3 N_B1_c_225_n 0.00132488f $X=3.355 $Y=1.105 $X2=0 $Y2=0
cc_149 N_A3_c_170_n N_B1_c_225_n 0.0165726f $X=3.455 $Y=1.217 $X2=0 $Y2=0
cc_150 N_A3_c_171_n N_VPWR_c_327_n 0.00429453f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A3_c_172_n N_VPWR_c_327_n 0.00597712f $X=3.455 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A3_c_171_n N_VPWR_c_324_n 0.00743756f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A3_c_172_n N_VPWR_c_324_n 0.0101953f $X=3.455 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A3_c_171_n N_A_309_297#_c_380_n 0.0144317f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A3_c_172_n N_A_309_297#_c_380_n 0.0012551f $X=3.455 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A3_c_171_n N_A_309_297#_c_387_n 0.00478129f $X=2.985 $Y=1.41 $X2=0
+ $Y2=0
cc_157 N_A3_c_172_n N_A_309_297#_c_387_n 0.00173218f $X=3.455 $Y=1.41 $X2=0
+ $Y2=0
cc_158 N_A3_c_171_n N_Y_c_417_n 0.0112095f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A3_c_172_n N_Y_c_417_n 0.0101048f $X=3.455 $Y=1.41 $X2=0 $Y2=0
cc_160 A3 N_Y_c_417_n 0.0369312f $X=3.355 $Y=1.105 $X2=0 $Y2=0
cc_161 N_A3_c_170_n N_Y_c_417_n 0.00155847f $X=3.455 $Y=1.217 $X2=0 $Y2=0
cc_162 N_A3_c_171_n N_Y_c_412_n 5.6422e-19 $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_163 A3 N_Y_c_412_n 0.0155155f $X=3.355 $Y=1.105 $X2=0 $Y2=0
cc_164 N_A3_c_170_n N_Y_c_412_n 5.82211e-19 $X=3.455 $Y=1.217 $X2=0 $Y2=0
cc_165 N_A3_c_171_n N_Y_c_424_n 7.81603e-19 $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A3_c_172_n N_Y_c_424_n 0.0130518f $X=3.455 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A3_c_172_n N_Y_c_426_n 0.00210477f $X=3.455 $Y=1.41 $X2=0 $Y2=0
cc_168 A3 N_Y_c_426_n 0.0058313f $X=3.355 $Y=1.105 $X2=0 $Y2=0
cc_169 N_A3_c_171_n N_Y_c_413_n 0.00675583f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A3_c_172_n N_Y_c_413_n 5.8173e-19 $X=3.455 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A3_M1003_g N_Y_c_411_n 2.59556e-19 $X=3.48 $Y=0.56 $X2=0 $Y2=0
cc_172 A3 N_Y_c_411_n 0.00863288f $X=3.355 $Y=1.105 $X2=0 $Y2=0
cc_173 N_A3_c_170_n N_Y_c_411_n 2.39662e-19 $X=3.455 $Y=1.217 $X2=0 $Y2=0
cc_174 N_A3_M1002_g N_A_27_47#_c_479_n 0.0109298f $X=2.86 $Y=0.56 $X2=0 $Y2=0
cc_175 N_A3_M1003_g N_A_27_47#_c_479_n 0.00909694f $X=3.48 $Y=0.56 $X2=0 $Y2=0
cc_176 A3 N_A_27_47#_c_479_n 0.0528486f $X=3.355 $Y=1.105 $X2=0 $Y2=0
cc_177 N_A3_c_170_n N_A_27_47#_c_479_n 0.00673116f $X=3.455 $Y=1.217 $X2=0 $Y2=0
cc_178 N_A3_M1003_g N_A_27_47#_c_503_n 0.00307151f $X=3.48 $Y=0.56 $X2=0 $Y2=0
cc_179 N_A3_M1002_g N_A_27_47#_c_504_n 9.08184e-19 $X=2.86 $Y=0.56 $X2=0 $Y2=0
cc_180 N_A3_M1003_g N_A_27_47#_c_504_n 0.00596939f $X=3.48 $Y=0.56 $X2=0 $Y2=0
cc_181 A3 N_A_27_47#_c_482_n 0.00347323f $X=3.355 $Y=1.105 $X2=0 $Y2=0
cc_182 N_A3_M1002_g N_VGND_c_560_n 0.00406603f $X=2.86 $Y=0.56 $X2=0 $Y2=0
cc_183 N_A3_M1002_g N_VGND_c_561_n 0.0126656f $X=2.86 $Y=0.56 $X2=0 $Y2=0
cc_184 N_A3_M1003_g N_VGND_c_561_n 0.00601389f $X=3.48 $Y=0.56 $X2=0 $Y2=0
cc_185 N_A3_M1003_g N_VGND_c_562_n 0.0039445f $X=3.48 $Y=0.56 $X2=0 $Y2=0
cc_186 N_A3_M1002_g N_VGND_c_563_n 0.00495145f $X=2.86 $Y=0.56 $X2=0 $Y2=0
cc_187 N_A3_M1003_g N_VGND_c_563_n 0.00608931f $X=3.48 $Y=0.56 $X2=0 $Y2=0
cc_188 N_B1_c_228_n N_VPWR_c_326_n 0.00988612f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_189 N_B1_c_230_n N_VPWR_c_326_n 0.0032802f $X=4.515 $Y=1.41 $X2=0 $Y2=0
cc_190 N_B1_c_228_n N_VPWR_c_327_n 0.00673617f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_191 N_B1_c_230_n N_VPWR_c_329_n 0.00702461f $X=4.515 $Y=1.41 $X2=0 $Y2=0
cc_192 N_B1_c_228_n N_VPWR_c_324_n 0.0122319f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_193 N_B1_c_230_n N_VPWR_c_324_n 0.0137532f $X=4.515 $Y=1.41 $X2=0 $Y2=0
cc_194 N_B1_c_228_n N_Y_c_424_n 0.0111638f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_195 N_B1_c_230_n N_Y_c_424_n 8.75359e-19 $X=4.515 $Y=1.41 $X2=0 $Y2=0
cc_196 N_B1_c_228_n N_Y_c_435_n 0.0192631f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_197 N_B1_c_228_n N_Y_c_426_n 8.61029e-19 $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_198 N_B1_c_222_n N_Y_c_411_n 0.00584658f $X=3.9 $Y=0.995 $X2=0 $Y2=0
cc_199 N_B1_c_228_n N_Y_c_411_n 0.00250514f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_200 N_B1_c_223_n N_Y_c_411_n 0.0278401f $X=4.415 $Y=1.16 $X2=0 $Y2=0
cc_201 N_B1_c_224_n N_Y_c_411_n 0.0121445f $X=4.49 $Y=0.995 $X2=0 $Y2=0
cc_202 N_B1_c_230_n N_Y_c_411_n 0.00502455f $X=4.515 $Y=1.41 $X2=0 $Y2=0
cc_203 N_B1_c_225_n N_Y_c_411_n 0.00253459f $X=3.925 $Y=1.202 $X2=0 $Y2=0
cc_204 B1 N_Y_c_411_n 0.0430967f $X=4.74 $Y=0.765 $X2=0 $Y2=0
cc_205 N_B1_c_227_n N_Y_c_411_n 0.0111587f $X=4.515 $Y=1.202 $X2=0 $Y2=0
cc_206 N_B1_c_223_n N_Y_c_415_n 0.00164082f $X=4.415 $Y=1.16 $X2=0 $Y2=0
cc_207 N_B1_c_230_n N_Y_c_415_n 0.0216635f $X=4.515 $Y=1.41 $X2=0 $Y2=0
cc_208 B1 N_Y_c_415_n 0.0249559f $X=4.74 $Y=0.765 $X2=0 $Y2=0
cc_209 N_B1_c_227_n N_Y_c_415_n 0.0021459f $X=4.515 $Y=1.202 $X2=0 $Y2=0
cc_210 B1 N_A_27_47#_M1008_s 0.0045945f $X=4.74 $Y=0.765 $X2=0 $Y2=0
cc_211 N_B1_c_222_n N_A_27_47#_c_479_n 0.00283679f $X=3.9 $Y=0.995 $X2=0 $Y2=0
cc_212 N_B1_c_222_n N_A_27_47#_c_503_n 7.12665e-19 $X=3.9 $Y=0.995 $X2=0 $Y2=0
cc_213 N_B1_c_222_n N_A_27_47#_c_504_n 0.00501931f $X=3.9 $Y=0.995 $X2=0 $Y2=0
cc_214 N_B1_c_224_n N_A_27_47#_c_504_n 6.83284e-19 $X=4.49 $Y=0.995 $X2=0 $Y2=0
cc_215 N_B1_c_222_n N_A_27_47#_c_480_n 0.0109058f $X=3.9 $Y=0.995 $X2=0 $Y2=0
cc_216 N_B1_c_223_n N_A_27_47#_c_480_n 0.00103884f $X=4.415 $Y=1.16 $X2=0 $Y2=0
cc_217 N_B1_c_224_n N_A_27_47#_c_480_n 0.0118459f $X=4.49 $Y=0.995 $X2=0 $Y2=0
cc_218 B1 N_A_27_47#_c_480_n 0.0274186f $X=4.74 $Y=0.765 $X2=0 $Y2=0
cc_219 N_B1_c_227_n N_A_27_47#_c_480_n 0.00242205f $X=4.515 $Y=1.202 $X2=0 $Y2=0
cc_220 N_B1_c_222_n N_VGND_c_562_n 0.00357835f $X=3.9 $Y=0.995 $X2=0 $Y2=0
cc_221 N_B1_c_224_n N_VGND_c_562_n 0.00357877f $X=4.49 $Y=0.995 $X2=0 $Y2=0
cc_222 N_B1_c_222_n N_VGND_c_563_n 0.00565346f $X=3.9 $Y=0.995 $X2=0 $Y2=0
cc_223 N_B1_c_224_n N_VGND_c_563_n 0.00666354f $X=4.49 $Y=0.995 $X2=0 $Y2=0
cc_224 B1 N_VGND_c_563_n 8.05634e-19 $X=4.74 $Y=0.765 $X2=0 $Y2=0
cc_225 N_A_27_297#_c_281_n N_VPWR_M1000_d 0.00327447f $X=1.005 $Y=1.58 $X2=-0.19
+ $Y2=1.305
cc_226 N_A_27_297#_c_275_n N_VPWR_c_325_n 0.0383577f $X=0.28 $Y=1.68 $X2=0 $Y2=0
cc_227 N_A_27_297#_c_281_n N_VPWR_c_325_n 0.0136682f $X=1.005 $Y=1.58 $X2=0
+ $Y2=0
cc_228 N_A_27_297#_c_288_n N_VPWR_c_325_n 0.0470327f $X=1.22 $Y=1.68 $X2=0 $Y2=0
cc_229 N_A_27_297#_c_288_n N_VPWR_c_327_n 0.0223557f $X=1.22 $Y=1.68 $X2=0 $Y2=0
cc_230 N_A_27_297#_M1000_s N_VPWR_c_324_n 0.00233913f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_231 N_A_27_297#_M1013_s N_VPWR_c_324_n 0.00231261f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_232 N_A_27_297#_M1009_d N_VPWR_c_324_n 0.00218346f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_233 N_A_27_297#_c_275_n N_VPWR_c_324_n 0.0134353f $X=0.28 $Y=1.68 $X2=0 $Y2=0
cc_234 N_A_27_297#_c_288_n N_VPWR_c_324_n 0.0140101f $X=1.22 $Y=1.68 $X2=0 $Y2=0
cc_235 N_A_27_297#_c_275_n N_VPWR_c_331_n 0.0228244f $X=0.28 $Y=1.68 $X2=0 $Y2=0
cc_236 N_A_27_297#_c_277_n N_A_309_297#_M1006_s 0.00327447f $X=1.945 $Y=1.58
+ $X2=-0.19 $Y2=1.305
cc_237 N_A_27_297#_c_288_n N_A_309_297#_c_381_n 0.0281258f $X=1.22 $Y=1.68 $X2=0
+ $Y2=0
cc_238 N_A_27_297#_c_277_n N_A_309_297#_c_381_n 0.0135833f $X=1.945 $Y=1.58
+ $X2=0 $Y2=0
cc_239 N_A_27_297#_c_278_n N_A_309_297#_c_381_n 0.02165f $X=2.16 $Y=1.68 $X2=0
+ $Y2=0
cc_240 N_A_27_297#_M1009_d N_A_309_297#_c_380_n 0.00510164f $X=2.015 $Y=1.485
+ $X2=0 $Y2=0
cc_241 N_A_27_297#_c_277_n N_A_309_297#_c_380_n 0.00252905f $X=1.945 $Y=1.58
+ $X2=0 $Y2=0
cc_242 N_A_27_297#_c_278_n N_A_309_297#_c_380_n 0.0240558f $X=2.16 $Y=1.68 $X2=0
+ $Y2=0
cc_243 N_A_27_297#_c_288_n N_A_309_297#_c_384_n 0.0116213f $X=1.22 $Y=1.68 $X2=0
+ $Y2=0
cc_244 N_A_27_297#_c_277_n N_Y_c_412_n 0.0118151f $X=1.945 $Y=1.58 $X2=0 $Y2=0
cc_245 N_A_27_297#_c_278_n N_Y_c_413_n 0.0287439f $X=2.16 $Y=1.68 $X2=0 $Y2=0
cc_246 N_A_27_297#_c_277_n N_A_27_47#_c_494_n 0.00268167f $X=1.945 $Y=1.58 $X2=0
+ $Y2=0
cc_247 N_A_27_297#_c_290_n N_A_27_47#_c_481_n 6.95815e-19 $X=1.195 $Y=1.58 $X2=0
+ $Y2=0
cc_248 N_VPWR_c_324_n N_A_309_297#_M1006_s 0.00441167f $X=4.83 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_249 N_VPWR_c_324_n N_A_309_297#_M1005_s 0.00441167f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_250 N_VPWR_c_327_n N_A_309_297#_c_380_n 0.0911766f $X=4.075 $Y=2.72 $X2=0
+ $Y2=0
cc_251 N_VPWR_c_324_n N_A_309_297#_c_380_n 0.0555268f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_252 N_VPWR_c_327_n N_A_309_297#_c_384_n 0.0118886f $X=4.075 $Y=2.72 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_324_n N_A_309_297#_c_384_n 0.00653405f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_324_n N_Y_M1005_d 0.00234744f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_255 N_VPWR_c_324_n N_Y_M1012_d 0.00231261f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_256 N_VPWR_c_324_n N_Y_M1010_s 0.00291223f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_257 N_VPWR_c_326_n N_Y_c_424_n 0.0405335f $X=4.24 $Y=2.02 $X2=0 $Y2=0
cc_258 N_VPWR_c_327_n N_Y_c_424_n 0.0223557f $X=4.075 $Y=2.72 $X2=0 $Y2=0
cc_259 N_VPWR_c_324_n N_Y_c_424_n 0.0140101f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_260 N_VPWR_M1001_d N_Y_c_411_n 9.84633e-19 $X=4.015 $Y=1.485 $X2=0 $Y2=0
cc_261 N_VPWR_M1001_d N_Y_c_415_n 0.00420284f $X=4.015 $Y=1.485 $X2=0 $Y2=0
cc_262 N_VPWR_c_326_n N_Y_c_415_n 0.0237567f $X=4.24 $Y=2.02 $X2=0 $Y2=0
cc_263 N_VPWR_c_329_n N_Y_c_416_n 0.0226365f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_264 N_VPWR_c_324_n N_Y_c_416_n 0.013017f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_265 N_A_309_297#_c_380_n N_Y_M1005_d 0.00568807f $X=3.135 $Y=2.38 $X2=0 $Y2=0
cc_266 N_A_309_297#_M1005_s N_Y_c_417_n 0.00327447f $X=3.075 $Y=1.485 $X2=0
+ $Y2=0
cc_267 N_A_309_297#_c_380_n N_Y_c_417_n 0.00367045f $X=3.135 $Y=2.38 $X2=0 $Y2=0
cc_268 N_A_309_297#_c_387_n N_Y_c_417_n 0.0135833f $X=3.22 $Y=2.135 $X2=0 $Y2=0
cc_269 N_A_309_297#_c_380_n N_Y_c_424_n 0.0141783f $X=3.135 $Y=2.38 $X2=0 $Y2=0
cc_270 N_A_309_297#_c_387_n N_Y_c_424_n 0.034305f $X=3.22 $Y=2.135 $X2=0 $Y2=0
cc_271 N_A_309_297#_c_380_n N_Y_c_413_n 0.0204533f $X=3.135 $Y=2.38 $X2=0 $Y2=0
cc_272 N_A_309_297#_c_387_n N_Y_c_413_n 0.0175572f $X=3.22 $Y=2.135 $X2=0 $Y2=0
cc_273 N_Y_c_426_n N_A_27_47#_c_479_n 0.00638344f $X=3.665 $Y=1.58 $X2=0 $Y2=0
cc_274 N_Y_c_411_n N_A_27_47#_c_479_n 0.0115938f $X=4.24 $Y=0.755 $X2=0 $Y2=0
cc_275 N_Y_c_411_n N_A_27_47#_c_504_n 0.00777416f $X=4.24 $Y=0.755 $X2=0 $Y2=0
cc_276 N_Y_M1007_d N_A_27_47#_c_480_n 0.00799721f $X=3.975 $Y=0.235 $X2=0 $Y2=0
cc_277 N_Y_c_411_n N_A_27_47#_c_480_n 0.0242317f $X=4.24 $Y=0.755 $X2=0 $Y2=0
cc_278 N_Y_c_412_n N_A_27_47#_c_482_n 0.00395489f $X=2.915 $Y=1.58 $X2=0 $Y2=0
cc_279 N_Y_M1007_d N_VGND_c_563_n 0.00354702f $X=3.975 $Y=0.235 $X2=0 $Y2=0
cc_280 N_A_27_47#_c_483_n N_VGND_M1004_d 0.00435938f $X=1.005 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_281 N_A_27_47#_c_494_n N_VGND_M1011_s 0.0165032f $X=2.425 $Y=0.8 $X2=0 $Y2=0
cc_282 N_A_27_47#_c_479_n N_VGND_M1002_s 0.00813081f $X=3.475 $Y=0.8 $X2=0 $Y2=0
cc_283 N_A_27_47#_c_483_n N_VGND_c_559_n 0.0126475f $X=1.005 $Y=0.8 $X2=0 $Y2=0
cc_284 N_A_27_47#_c_489_n N_VGND_c_559_n 0.0216501f $X=1.22 $Y=0.36 $X2=0 $Y2=0
cc_285 N_A_27_47#_c_494_n N_VGND_c_560_n 0.00320671f $X=2.425 $Y=0.8 $X2=0 $Y2=0
cc_286 N_A_27_47#_c_531_p N_VGND_c_560_n 0.0204563f $X=2.59 $Y=0.36 $X2=0 $Y2=0
cc_287 N_A_27_47#_c_479_n N_VGND_c_560_n 0.0021402f $X=3.475 $Y=0.8 $X2=0 $Y2=0
cc_288 N_A_27_47#_c_479_n N_VGND_c_561_n 0.0250159f $X=3.475 $Y=0.8 $X2=0 $Y2=0
cc_289 N_A_27_47#_c_503_n N_VGND_c_561_n 0.0141542f $X=3.665 $Y=0.425 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_504_n N_VGND_c_561_n 0.00947726f $X=3.665 $Y=0.715 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_479_n N_VGND_c_562_n 0.00203275f $X=3.475 $Y=0.8 $X2=0 $Y2=0
cc_292 N_A_27_47#_c_503_n N_VGND_c_562_n 0.0223473f $X=3.665 $Y=0.425 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_480_n N_VGND_c_562_n 0.0660977f $X=4.63 $Y=0.34 $X2=0 $Y2=0
cc_294 N_A_27_47#_M1004_s N_VGND_c_563_n 0.00275065f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_M1015_s N_VGND_c_563_n 0.00215201f $X=1.085 $Y=0.235 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_M1014_d N_VGND_c_563_n 0.0031222f $X=2.415 $Y=0.235 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_M1003_d N_VGND_c_563_n 0.00215201f $X=3.555 $Y=0.235 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_M1008_s N_VGND_c_563_n 0.00253611f $X=4.565 $Y=0.235 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_477_n N_VGND_c_563_n 0.0135674f $X=0.28 $Y=0.36 $X2=0 $Y2=0
cc_300 N_A_27_47#_c_483_n N_VGND_c_563_n 0.00983826f $X=1.005 $Y=0.8 $X2=0 $Y2=0
cc_301 N_A_27_47#_c_489_n N_VGND_c_563_n 0.0138899f $X=1.22 $Y=0.36 $X2=0 $Y2=0
cc_302 N_A_27_47#_c_494_n N_VGND_c_563_n 0.0135107f $X=2.425 $Y=0.8 $X2=0 $Y2=0
cc_303 N_A_27_47#_c_531_p N_VGND_c_563_n 0.0126066f $X=2.59 $Y=0.36 $X2=0 $Y2=0
cc_304 N_A_27_47#_c_479_n N_VGND_c_563_n 0.0094773f $X=3.475 $Y=0.8 $X2=0 $Y2=0
cc_305 N_A_27_47#_c_503_n N_VGND_c_563_n 0.0139576f $X=3.665 $Y=0.425 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_480_n N_VGND_c_563_n 0.0401602f $X=4.63 $Y=0.34 $X2=0 $Y2=0
cc_307 N_A_27_47#_c_477_n N_VGND_c_564_n 0.0235041f $X=0.28 $Y=0.36 $X2=0 $Y2=0
cc_308 N_A_27_47#_c_483_n N_VGND_c_564_n 0.00259521f $X=1.005 $Y=0.8 $X2=0 $Y2=0
cc_309 N_A_27_47#_c_483_n N_VGND_c_565_n 0.00203275f $X=1.005 $Y=0.8 $X2=0 $Y2=0
cc_310 N_A_27_47#_c_489_n N_VGND_c_565_n 0.0222117f $X=1.22 $Y=0.36 $X2=0 $Y2=0
cc_311 N_A_27_47#_c_494_n N_VGND_c_565_n 0.00271675f $X=2.425 $Y=0.8 $X2=0 $Y2=0
cc_312 N_A_27_47#_c_489_n N_VGND_c_566_n 0.0194526f $X=1.22 $Y=0.36 $X2=0 $Y2=0
cc_313 N_A_27_47#_c_494_n N_VGND_c_566_n 0.0434928f $X=2.425 $Y=0.8 $X2=0 $Y2=0
