# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__and4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 0.765000 0.840000 1.635000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.810000 0.735000 4.190000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.330000 0.755000 3.640000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.870000 0.995000 3.120000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.030000 0.255000 1.340000 0.650000 ;
        RECT 1.030000 0.650000 2.280000 0.820000 ;
        RECT 1.030000 0.820000 1.360000 1.545000 ;
        RECT 1.030000 1.545000 2.360000 1.715000 ;
        RECT 2.110000 0.255000 2.280000 0.650000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.585000 ;
      RECT 0.085000  0.585000 0.260000 1.915000 ;
      RECT 0.085000  1.915000 4.885000 2.085000 ;
      RECT 0.085000  2.085000 0.345000 2.465000 ;
      RECT 0.515000  2.255000 0.895000 2.635000 ;
      RECT 0.565000  0.085000 0.815000 0.545000 ;
      RECT 1.510000  0.085000 1.890000 0.470000 ;
      RECT 1.510000  2.255000 1.890000 2.635000 ;
      RECT 1.530000  0.995000 2.700000 1.325000 ;
      RECT 2.450000  2.255000 2.830000 2.635000 ;
      RECT 2.530000  1.325000 2.700000 1.545000 ;
      RECT 2.530000  1.545000 4.530000 1.715000 ;
      RECT 2.535000  0.085000 2.865000 0.445000 ;
      RECT 3.510000  2.255000 3.890000 2.635000 ;
      RECT 4.360000  0.640000 4.900000 0.810000 ;
      RECT 4.360000  0.810000 4.530000 1.545000 ;
      RECT 4.570000  2.255000 4.950000 2.635000 ;
      RECT 4.715000  0.995000 4.885000 1.915000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4b_4
END LIBRARY
