* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__xor3_1 A B C VGND VNB VPB VPWR X
X0 a_991_365# B a_424_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 a_406_325# C a_116_21# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X2 a_406_325# a_875_297# a_991_365# VNB sky130_fd_pr__nfet_01v8 w=600000u l=150000u
X3 X a_116_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 a_991_365# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_406_325# a_875_297# a_1276_297# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X6 a_116_21# a_276_93# a_424_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X7 VPWR B a_875_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 a_424_49# a_875_297# a_1276_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_991_365# B a_406_325# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X10 VGND C a_276_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VGND a_991_365# a_1276_297# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 a_1276_297# B a_424_49# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X13 a_116_21# a_276_93# a_406_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X14 X a_116_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND B a_875_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_991_365# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 VPWR C a_276_93# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X18 a_424_49# a_875_297# a_991_365# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X19 a_424_49# C a_116_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 VPWR a_991_365# a_1276_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 a_1276_297# B a_406_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
