* NGSPICE file created from sky130_fd_sc_hdll__and4bb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
M1000 a_425_93# a_27_47# a_339_93# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.176e+11p ps=1.4e+06u
M1001 a_615_93# C a_511_93# VNB nshort w=420000u l=150000u
+  ad=1.89e+11p pd=1.74e+06u as=1.554e+11p ps=1.58e+06u
M1002 a_339_93# C VPWR VPB phighvt w=420000u l=180000u
+  ad=2.814e+11p pd=3.02e+06u as=6.779e+11p ps=7.03e+06u
M1003 a_511_93# a_225_413# a_425_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_225_413# B_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1005 VPWR a_225_413# a_339_93# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR D a_339_93# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_225_413# B_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=3.861e+11p ps=3.65e+06u
M1008 VGND A_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1009 VGND D a_615_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_339_93# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1011 VPWR A_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
M1012 a_339_93# a_27_47# VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_339_93# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
.ends

