* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__xnor2_1 A B VGND VNB VPB VPWR Y
X0 Y a_47_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_47_47# B a_139_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND B a_315_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR A a_415_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 VGND A a_315_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_47_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_415_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 VPWR B a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 a_315_47# a_47_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_139_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
