* File: sky130_fd_sc_hdll__nand4_2.pxi.spice
* Created: Wed Sep  2 08:38:24 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND4_2%D N_D_c_76_n N_D_M1000_g N_D_M1002_g N_D_c_77_n
+ N_D_M1009_g N_D_M1012_g D D N_D_c_74_n N_D_c_75_n
+ PM_SKY130_FD_SC_HDLL__NAND4_2%D
x_PM_SKY130_FD_SC_HDLL__NAND4_2%C N_C_M1005_g N_C_c_121_n N_C_M1011_g
+ N_C_c_122_n N_C_M1015_g N_C_M1013_g C C N_C_c_120_n
+ PM_SKY130_FD_SC_HDLL__NAND4_2%C
x_PM_SKY130_FD_SC_HDLL__NAND4_2%B N_B_c_170_n N_B_M1001_g N_B_c_171_n
+ N_B_M1006_g N_B_M1004_g N_B_M1010_g N_B_c_167_n N_B_c_168_n B B B
+ PM_SKY130_FD_SC_HDLL__NAND4_2%B
x_PM_SKY130_FD_SC_HDLL__NAND4_2%A N_A_M1007_g N_A_c_222_n N_A_M1003_g
+ N_A_M1008_g N_A_c_223_n N_A_M1014_g N_A_c_219_n A N_A_c_221_n A
+ PM_SKY130_FD_SC_HDLL__NAND4_2%A
x_PM_SKY130_FD_SC_HDLL__NAND4_2%VPWR N_VPWR_M1000_d N_VPWR_M1009_d
+ N_VPWR_M1015_d N_VPWR_M1006_d N_VPWR_M1014_s N_VPWR_c_258_n N_VPWR_c_259_n
+ N_VPWR_c_260_n N_VPWR_c_261_n N_VPWR_c_262_n N_VPWR_c_263_n N_VPWR_c_264_n
+ N_VPWR_c_265_n N_VPWR_c_266_n VPWR N_VPWR_c_267_n N_VPWR_c_268_n
+ N_VPWR_c_269_n N_VPWR_c_270_n N_VPWR_c_271_n N_VPWR_c_257_n
+ PM_SKY130_FD_SC_HDLL__NAND4_2%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND4_2%Y N_Y_M1007_s N_Y_M1000_s N_Y_M1011_s
+ N_Y_M1001_s N_Y_M1003_d N_Y_c_332_n N_Y_c_343_n N_Y_c_333_n N_Y_c_347_n
+ N_Y_c_334_n N_Y_c_357_n N_Y_c_368_n N_Y_c_384_n N_Y_c_335_n Y Y Y Y Y
+ PM_SKY130_FD_SC_HDLL__NAND4_2%Y
x_PM_SKY130_FD_SC_HDLL__NAND4_2%A_27_47# N_A_27_47#_M1002_d N_A_27_47#_M1012_d
+ N_A_27_47#_M1013_s N_A_27_47#_c_429_n N_A_27_47#_c_430_n N_A_27_47#_c_431_n
+ N_A_27_47#_c_439_n N_A_27_47#_c_440_n N_A_27_47#_c_432_n
+ PM_SKY130_FD_SC_HDLL__NAND4_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NAND4_2%VGND N_VGND_M1002_s N_VGND_c_470_n VGND
+ N_VGND_c_471_n N_VGND_c_472_n N_VGND_c_473_n
+ PM_SKY130_FD_SC_HDLL__NAND4_2%VGND
x_PM_SKY130_FD_SC_HDLL__NAND4_2%A_297_47# N_A_297_47#_M1005_d
+ N_A_297_47#_M1004_s N_A_297_47#_c_524_n
+ PM_SKY130_FD_SC_HDLL__NAND4_2%A_297_47#
x_PM_SKY130_FD_SC_HDLL__NAND4_2%A_511_47# N_A_511_47#_M1004_d
+ N_A_511_47#_M1010_d N_A_511_47#_M1008_d N_A_511_47#_c_547_n
+ N_A_511_47#_c_548_n N_A_511_47#_c_553_n N_A_511_47#_c_549_n
+ N_A_511_47#_c_550_n N_A_511_47#_c_576_n
+ PM_SKY130_FD_SC_HDLL__NAND4_2%A_511_47#
cc_1 VNB N_D_M1002_g 0.0244378f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_2 VNB N_D_M1012_g 0.0180932f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_3 VNB D 0.00806404f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_4 VNB N_D_c_74_n 0.0251778f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.217
cc_5 VNB N_D_c_75_n 0.0352518f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.217
cc_6 VNB N_C_M1005_g 0.0187386f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_7 VNB N_C_M1013_g 0.0249344f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.025
cc_8 VNB C 0.0058494f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_C_c_120_n 0.0421077f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.16
cc_10 VNB N_B_M1004_g 0.0244378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B_M1010_g 0.0183272f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.025
cc_12 VNB N_B_c_167_n 0.0443835f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_13 VNB N_B_c_168_n 0.0325603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB B 0.00223853f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.217
cc_15 VNB N_A_M1007_g 0.0177431f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_16 VNB N_A_M1008_g 0.0238147f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_17 VNB N_A_c_219_n 0.0372266f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_18 VNB A 0.00738464f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_c_221_n 0.0362156f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.217
cc_20 VNB N_VPWR_c_257_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB Y 0.00348027f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_429_n 0.0189842f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_23 VNB N_A_27_47#_c_430_n 0.00489008f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_24 VNB N_A_27_47#_c_431_n 0.00944083f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_25 VNB N_A_27_47#_c_432_n 0.00261848f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.217
cc_26 VNB N_VGND_c_470_n 0.00467885f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_27 VNB N_VGND_c_471_n 0.100042f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_28 VNB N_VGND_c_472_n 0.264202f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_29 VNB N_VGND_c_473_n 0.0219649f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.217
cc_30 VNB N_A_297_47#_c_524_n 0.020767f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_31 VNB N_A_511_47#_c_547_n 0.00247236f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_32 VNB N_A_511_47#_c_548_n 0.00214417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_511_47#_c_549_n 0.00884635f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_511_47#_c_550_n 0.0191075f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.217
cc_35 VPB N_D_c_76_n 0.0208995f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_36 VPB N_D_c_77_n 0.0160015f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_37 VPB N_D_c_74_n 0.00813297f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.217
cc_38 VPB N_D_c_75_n 0.0163834f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.217
cc_39 VPB N_C_c_121_n 0.0160015f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_40 VPB N_C_c_122_n 0.0170915f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_41 VPB N_C_c_120_n 0.0136043f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.16
cc_42 VPB N_B_c_170_n 0.0170915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_B_c_171_n 0.0195191f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_44 VPB N_B_c_167_n 0.0149219f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_45 VPB N_A_c_222_n 0.0192858f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_46 VPB N_A_c_223_n 0.0197118f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_47 VPB N_A_c_219_n 0.0161499f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_48 VPB N_A_c_221_n 0.0137398f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.217
cc_49 VPB N_VPWR_c_258_n 0.00994749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_259_n 0.0428976f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_51 VPB N_VPWR_c_260_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.217
cc_52 VPB N_VPWR_c_261_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.217
cc_53 VPB N_VPWR_c_262_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.175
cc_54 VPB N_VPWR_c_263_n 0.00559947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_264_n 0.00592343f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_265_n 0.0144238f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_266_n 0.00997332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_267_n 0.0250959f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_268_n 0.0238197f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_269_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_270_n 0.00631825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_271_n 0.00728331f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_257_n 0.0451585f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_Y_c_332_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_Y_c_333_n 0.00263714f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_Y_c_334_n 0.00678549f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.217
cc_67 VPB N_Y_c_335_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB Y 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB Y 0.00243373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB Y 0.00750013f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 N_D_M1012_g N_C_M1005_g 0.0172236f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_72 N_D_c_77_n N_C_c_121_n 0.0231619f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_73 D C 0.0167609f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_74 N_D_c_75_n C 0.00215451f $X=0.965 $Y=1.217 $X2=0 $Y2=0
cc_75 N_D_c_75_n N_C_c_120_n 0.0172236f $X=0.965 $Y=1.217 $X2=0 $Y2=0
cc_76 N_D_c_76_n N_VPWR_c_259_n 0.00777002f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_77 D N_VPWR_c_259_n 0.0153565f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_78 N_D_c_74_n N_VPWR_c_259_n 0.00533558f $X=0.495 $Y=1.217 $X2=0 $Y2=0
cc_79 N_D_c_76_n N_VPWR_c_260_n 0.00597712f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_80 N_D_c_77_n N_VPWR_c_260_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_81 N_D_c_77_n N_VPWR_c_261_n 0.0052072f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_82 N_D_c_76_n N_VPWR_c_257_n 0.010906f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_83 N_D_c_77_n N_VPWR_c_257_n 0.011869f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_84 N_D_c_76_n N_Y_c_332_n 0.0065257f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_85 N_D_c_77_n N_Y_c_332_n 0.00116723f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_86 D N_Y_c_332_n 0.0305808f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_87 N_D_c_75_n N_Y_c_332_n 0.0074788f $X=0.965 $Y=1.217 $X2=0 $Y2=0
cc_88 N_D_c_76_n N_Y_c_343_n 0.0121679f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_89 N_D_c_77_n N_Y_c_343_n 0.0106251f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_90 N_D_c_77_n N_Y_c_333_n 0.0172881f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_91 N_D_c_75_n N_Y_c_333_n 3.62694e-19 $X=0.965 $Y=1.217 $X2=0 $Y2=0
cc_92 N_D_c_77_n N_Y_c_347_n 6.48386e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_93 N_D_M1002_g N_A_27_47#_c_430_n 0.0107881f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_94 N_D_M1012_g N_A_27_47#_c_430_n 0.010458f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_95 D N_A_27_47#_c_430_n 0.0334223f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_96 N_D_c_75_n N_A_27_47#_c_430_n 0.00375198f $X=0.965 $Y=1.217 $X2=0 $Y2=0
cc_97 D N_A_27_47#_c_431_n 0.0255512f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_98 N_D_c_74_n N_A_27_47#_c_431_n 0.0076176f $X=0.495 $Y=1.217 $X2=0 $Y2=0
cc_99 N_D_M1012_g N_A_27_47#_c_439_n 0.00359564f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_100 N_D_M1002_g N_A_27_47#_c_440_n 5.85588e-19 $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_101 N_D_M1012_g N_A_27_47#_c_440_n 0.00521436f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_102 N_D_M1002_g N_VGND_c_470_n 0.00276126f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_103 N_D_M1012_g N_VGND_c_470_n 0.00356343f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_104 N_D_M1012_g N_VGND_c_471_n 0.00395719f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_105 N_D_M1002_g N_VGND_c_472_n 0.00703713f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_106 N_D_M1012_g N_VGND_c_472_n 0.00573562f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_107 N_D_M1002_g N_VGND_c_473_n 0.00439206f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_108 N_C_c_122_n N_B_c_170_n 0.0255255f $X=1.905 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_109 N_C_c_120_n N_B_c_167_n 0.0125483f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_110 C B 0.00600453f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_111 N_C_c_120_n B 0.0010017f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_112 N_C_c_121_n N_VPWR_c_261_n 0.004751f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_113 N_C_c_121_n N_VPWR_c_262_n 0.00597712f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_114 N_C_c_122_n N_VPWR_c_262_n 0.00673617f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_115 N_C_c_122_n N_VPWR_c_263_n 0.0102497f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_116 N_C_c_121_n N_VPWR_c_257_n 0.0100198f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_117 N_C_c_122_n N_VPWR_c_257_n 0.0122924f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_118 N_C_c_121_n N_Y_c_343_n 6.24674e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_119 N_C_c_121_n N_Y_c_333_n 0.0113403f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_120 C N_Y_c_333_n 0.0293961f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_121 N_C_c_120_n N_Y_c_333_n 3.10838e-19 $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_122 N_C_c_121_n N_Y_c_347_n 0.0130707f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_123 N_C_c_122_n N_Y_c_347_n 0.011306f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_124 N_C_c_122_n N_Y_c_334_n 0.0181008f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_125 C N_Y_c_334_n 0.00101487f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_126 N_C_c_120_n N_Y_c_334_n 3.62813e-19 $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_127 N_C_c_122_n N_Y_c_357_n 9.17942e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_128 N_C_c_121_n N_Y_c_335_n 0.00292783f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_129 N_C_c_122_n N_Y_c_335_n 0.00116723f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_130 C N_Y_c_335_n 0.0305808f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_131 N_C_c_120_n N_Y_c_335_n 0.00723098f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_132 C N_A_27_47#_c_430_n 0.0187199f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_133 N_C_M1005_g N_A_27_47#_c_432_n 0.0110186f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_134 N_C_M1013_g N_A_27_47#_c_432_n 0.00935436f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_135 C N_A_27_47#_c_432_n 0.00368637f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_136 N_C_M1005_g N_VGND_c_471_n 0.00357877f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_137 N_C_M1013_g N_VGND_c_471_n 0.00357877f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_138 N_C_M1005_g N_VGND_c_472_n 0.005504f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_139 N_C_M1013_g N_VGND_c_472_n 0.00680287f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_140 N_C_M1005_g N_A_297_47#_c_524_n 0.00389235f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_141 N_C_M1013_g N_A_297_47#_c_524_n 0.0164699f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_142 C N_A_297_47#_c_524_n 0.0295549f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_143 N_C_c_120_n N_A_297_47#_c_524_n 0.00438872f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_144 N_B_M1010_g N_A_M1007_g 0.0133074f $X=3.48 $Y=0.56 $X2=0 $Y2=0
cc_145 N_B_c_167_n N_A_c_219_n 0.00120824f $X=3.105 $Y=1.16 $X2=0 $Y2=0
cc_146 N_B_c_168_n N_A_c_219_n 0.0133074f $X=3.405 $Y=1.16 $X2=0 $Y2=0
cc_147 N_B_c_170_n N_VPWR_c_263_n 0.00971824f $X=2.535 $Y=1.41 $X2=0 $Y2=0
cc_148 N_B_c_171_n N_VPWR_c_264_n 0.0180703f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_149 N_B_c_170_n N_VPWR_c_267_n 0.00597712f $X=2.535 $Y=1.41 $X2=0 $Y2=0
cc_150 N_B_c_171_n N_VPWR_c_267_n 0.00673617f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_151 N_B_c_170_n N_VPWR_c_257_n 0.0104431f $X=2.535 $Y=1.41 $X2=0 $Y2=0
cc_152 N_B_c_171_n N_VPWR_c_257_n 0.013351f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_153 N_B_c_170_n N_Y_c_347_n 8.7249e-19 $X=2.535 $Y=1.41 $X2=0 $Y2=0
cc_154 N_B_c_170_n N_Y_c_334_n 0.0123232f $X=2.535 $Y=1.41 $X2=0 $Y2=0
cc_155 N_B_c_167_n N_Y_c_334_n 2.73568e-19 $X=3.105 $Y=1.16 $X2=0 $Y2=0
cc_156 B N_Y_c_334_n 0.00840447f $X=3.21 $Y=1.105 $X2=0 $Y2=0
cc_157 N_B_c_170_n N_Y_c_357_n 0.0137562f $X=2.535 $Y=1.41 $X2=0 $Y2=0
cc_158 N_B_c_171_n N_Y_c_357_n 0.0176136f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_159 N_B_M1010_g N_Y_c_368_n 8.9525e-19 $X=3.48 $Y=0.56 $X2=0 $Y2=0
cc_160 N_B_c_170_n Y 0.00292783f $X=2.535 $Y=1.41 $X2=0 $Y2=0
cc_161 N_B_c_171_n Y 0.00116723f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_162 N_B_c_167_n Y 0.00675985f $X=3.105 $Y=1.16 $X2=0 $Y2=0
cc_163 B Y 0.0305808f $X=3.21 $Y=1.105 $X2=0 $Y2=0
cc_164 N_B_c_171_n Y 0.00131833f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_165 N_B_c_167_n Y 0.00210946f $X=3.105 $Y=1.16 $X2=0 $Y2=0
cc_166 N_B_c_168_n Y 0.00319209f $X=3.405 $Y=1.16 $X2=0 $Y2=0
cc_167 B Y 0.0103636f $X=3.21 $Y=1.105 $X2=0 $Y2=0
cc_168 N_B_c_171_n Y 0.0178161f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_169 N_B_c_167_n Y 3.10838e-19 $X=3.105 $Y=1.16 $X2=0 $Y2=0
cc_170 N_B_c_168_n Y 0.0142667f $X=3.405 $Y=1.16 $X2=0 $Y2=0
cc_171 B Y 0.0321882f $X=3.21 $Y=1.105 $X2=0 $Y2=0
cc_172 N_B_M1004_g N_A_27_47#_c_432_n 7.1971e-19 $X=3.01 $Y=0.56 $X2=0 $Y2=0
cc_173 N_B_M1004_g N_VGND_c_471_n 0.00357877f $X=3.01 $Y=0.56 $X2=0 $Y2=0
cc_174 N_B_M1010_g N_VGND_c_471_n 0.00357877f $X=3.48 $Y=0.56 $X2=0 $Y2=0
cc_175 N_B_M1004_g N_VGND_c_472_n 0.00677297f $X=3.01 $Y=0.56 $X2=0 $Y2=0
cc_176 N_B_M1010_g N_VGND_c_472_n 0.00538422f $X=3.48 $Y=0.56 $X2=0 $Y2=0
cc_177 N_B_M1004_g N_A_297_47#_c_524_n 0.0145739f $X=3.01 $Y=0.56 $X2=0 $Y2=0
cc_178 N_B_M1010_g N_A_297_47#_c_524_n 3.04133e-19 $X=3.48 $Y=0.56 $X2=0 $Y2=0
cc_179 N_B_c_167_n N_A_297_47#_c_524_n 0.0126239f $X=3.105 $Y=1.16 $X2=0 $Y2=0
cc_180 N_B_c_168_n N_A_297_47#_c_524_n 0.00323379f $X=3.405 $Y=1.16 $X2=0 $Y2=0
cc_181 B N_A_297_47#_c_524_n 0.0703552f $X=3.21 $Y=1.105 $X2=0 $Y2=0
cc_182 N_B_M1004_g N_A_511_47#_c_547_n 0.0135941f $X=3.01 $Y=0.56 $X2=0 $Y2=0
cc_183 N_B_M1010_g N_A_511_47#_c_547_n 0.0137288f $X=3.48 $Y=0.56 $X2=0 $Y2=0
cc_184 N_A_c_222_n N_VPWR_c_264_n 0.0183448f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A_c_223_n N_VPWR_c_266_n 0.0297054f $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_186 A N_VPWR_c_266_n 0.0211194f $X=4.735 $Y=1.105 $X2=0 $Y2=0
cc_187 N_A_c_221_n N_VPWR_c_266_n 0.00805837f $X=4.78 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A_c_222_n N_VPWR_c_268_n 0.00597712f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A_c_223_n N_VPWR_c_268_n 0.00673617f $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_190 N_A_c_222_n N_VPWR_c_257_n 0.0115018f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_191 N_A_c_223_n N_VPWR_c_257_n 0.0129968f $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_192 N_A_M1007_g N_Y_c_368_n 0.00745156f $X=3.9 $Y=0.56 $X2=0 $Y2=0
cc_193 N_A_M1008_g N_Y_c_368_n 0.010862f $X=4.37 $Y=0.56 $X2=0 $Y2=0
cc_194 N_A_c_219_n N_Y_c_368_n 0.00584162f $X=4.495 $Y=1.165 $X2=0 $Y2=0
cc_195 N_A_c_222_n N_Y_c_384_n 0.0194822f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A_c_223_n N_Y_c_384_n 0.0100147f $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A_c_222_n Y 0.0150179f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_c_223_n Y 0.00517802f $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A_c_219_n Y 0.0412385f $X=4.495 $Y=1.165 $X2=0 $Y2=0
cc_200 A Y 0.0101989f $X=4.735 $Y=1.105 $X2=0 $Y2=0
cc_201 N_A_c_222_n Y 0.00135015f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A_M1007_g N_VGND_c_471_n 0.00357877f $X=3.9 $Y=0.56 $X2=0 $Y2=0
cc_203 N_A_M1008_g N_VGND_c_471_n 0.00357877f $X=4.37 $Y=0.56 $X2=0 $Y2=0
cc_204 N_A_M1007_g N_VGND_c_472_n 0.00538422f $X=3.9 $Y=0.56 $X2=0 $Y2=0
cc_205 N_A_M1008_g N_VGND_c_472_n 0.00654724f $X=4.37 $Y=0.56 $X2=0 $Y2=0
cc_206 N_A_M1007_g N_A_511_47#_c_553_n 0.0106231f $X=3.9 $Y=0.56 $X2=0 $Y2=0
cc_207 N_A_M1008_g N_A_511_47#_c_553_n 0.0174287f $X=4.37 $Y=0.56 $X2=0 $Y2=0
cc_208 N_A_c_219_n N_A_511_47#_c_553_n 0.00237535f $X=4.495 $Y=1.165 $X2=0 $Y2=0
cc_209 N_A_M1008_g N_A_511_47#_c_550_n 0.0127115f $X=4.37 $Y=0.56 $X2=0 $Y2=0
cc_210 A N_A_511_47#_c_550_n 0.0210372f $X=4.735 $Y=1.105 $X2=0 $Y2=0
cc_211 N_A_c_221_n N_A_511_47#_c_550_n 0.00822743f $X=4.78 $Y=1.16 $X2=0 $Y2=0
cc_212 N_VPWR_c_257_n N_Y_M1000_s 0.00231261f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_213 N_VPWR_c_257_n N_Y_M1011_s 0.00231261f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_214 N_VPWR_c_257_n N_Y_M1001_s 0.00231261f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_215 N_VPWR_c_257_n N_Y_M1003_d 0.00231261f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_216 N_VPWR_c_259_n N_Y_c_332_n 0.0137498f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_217 N_VPWR_c_259_n N_Y_c_343_n 0.0615045f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_218 N_VPWR_c_260_n N_Y_c_343_n 0.0223557f $X=1.115 $Y=2.72 $X2=0 $Y2=0
cc_219 N_VPWR_c_261_n N_Y_c_343_n 0.0385613f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_220 N_VPWR_c_257_n N_Y_c_343_n 0.0140101f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_221 N_VPWR_M1009_d N_Y_c_333_n 0.00180012f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_222 N_VPWR_c_261_n N_Y_c_333_n 0.0139097f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_223 N_VPWR_c_261_n N_Y_c_347_n 0.0470327f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_224 N_VPWR_c_262_n N_Y_c_347_n 0.0223557f $X=2.055 $Y=2.72 $X2=0 $Y2=0
cc_225 N_VPWR_c_263_n N_Y_c_347_n 0.0405335f $X=2.22 $Y=2 $X2=0 $Y2=0
cc_226 N_VPWR_c_257_n N_Y_c_347_n 0.0140101f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_227 N_VPWR_M1015_d N_Y_c_334_n 0.00440622f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_228 N_VPWR_c_263_n N_Y_c_334_n 0.027157f $X=2.22 $Y=2 $X2=0 $Y2=0
cc_229 N_VPWR_c_263_n N_Y_c_357_n 0.0494193f $X=2.22 $Y=2 $X2=0 $Y2=0
cc_230 N_VPWR_c_264_n N_Y_c_357_n 0.0280788f $X=3.46 $Y=2 $X2=0 $Y2=0
cc_231 N_VPWR_c_267_n N_Y_c_357_n 0.0223557f $X=3.295 $Y=2.72 $X2=0 $Y2=0
cc_232 N_VPWR_c_257_n N_Y_c_357_n 0.0140101f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_233 N_VPWR_c_264_n N_Y_c_384_n 0.035042f $X=3.46 $Y=2 $X2=0 $Y2=0
cc_234 N_VPWR_c_268_n N_Y_c_384_n 0.0223557f $X=4.545 $Y=2.72 $X2=0 $Y2=0
cc_235 N_VPWR_c_257_n N_Y_c_384_n 0.0140101f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_236 N_VPWR_M1006_d Y 0.0030349f $X=3.095 $Y=1.485 $X2=0 $Y2=0
cc_237 N_VPWR_c_266_n Y 0.0661633f $X=4.71 $Y=1.66 $X2=0 $Y2=0
cc_238 N_VPWR_M1006_d Y 0.0156626f $X=3.095 $Y=1.485 $X2=0 $Y2=0
cc_239 N_VPWR_c_264_n Y 0.0312967f $X=3.46 $Y=2 $X2=0 $Y2=0
cc_240 N_VPWR_c_259_n N_A_27_47#_c_431_n 7.42972e-19 $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_241 N_VPWR_c_266_n N_A_511_47#_c_550_n 0.0028454f $X=4.71 $Y=1.66 $X2=0 $Y2=0
cc_242 N_Y_c_333_n N_A_27_47#_c_430_n 0.004887f $X=1.455 $Y=1.555 $X2=0 $Y2=0
cc_243 N_Y_M1007_s N_VGND_c_472_n 0.00256987f $X=3.975 $Y=0.235 $X2=0 $Y2=0
cc_244 N_Y_c_334_n N_A_297_47#_c_524_n 0.019717f $X=2.555 $Y=1.555 $X2=0 $Y2=0
cc_245 N_Y_c_368_n N_A_297_47#_c_524_n 6.34677e-19 $X=4.16 $Y=0.72 $X2=0 $Y2=0
cc_246 Y N_A_511_47#_c_548_n 0.0045377f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_247 Y N_A_511_47#_c_548_n 0.00392188f $X=3.72 $Y=1.445 $X2=0 $Y2=0
cc_248 N_Y_M1007_s N_A_511_47#_c_553_n 0.00400901f $X=3.975 $Y=0.235 $X2=0 $Y2=0
cc_249 N_Y_c_368_n N_A_511_47#_c_553_n 0.020229f $X=4.16 $Y=0.72 $X2=0 $Y2=0
cc_250 Y N_A_511_47#_c_553_n 0.00423076f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_251 N_Y_c_368_n N_A_511_47#_c_550_n 0.0174035f $X=4.16 $Y=0.72 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_430_n N_VGND_M1002_s 0.00259473f $X=0.985 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_253 N_A_27_47#_c_430_n N_VGND_c_470_n 0.0115453f $X=0.985 $Y=0.82 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_439_n N_VGND_c_470_n 0.0165057f $X=1.135 $Y=0.465 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_440_n N_VGND_c_470_n 0.00582645f $X=1.2 $Y=0.72 $X2=0 $Y2=0
cc_256 N_A_27_47#_c_430_n N_VGND_c_471_n 0.00194552f $X=0.985 $Y=0.82 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_439_n N_VGND_c_471_n 0.0186086f $X=1.135 $Y=0.465 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_c_432_n N_VGND_c_471_n 0.0598688f $X=2.16 $Y=0.38 $X2=0 $Y2=0
cc_259 N_A_27_47#_M1002_d N_VGND_c_472_n 0.00259235f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_M1012_d N_VGND_c_472_n 0.00215206f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_M1013_s N_VGND_c_472_n 0.00225742f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_429_n N_VGND_c_472_n 0.0128092f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_430_n N_VGND_c_472_n 0.00969159f $X=0.985 $Y=0.82 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_439_n N_VGND_c_472_n 0.0111017f $X=1.135 $Y=0.465 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_432_n N_VGND_c_472_n 0.0374007f $X=2.16 $Y=0.38 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_429_n N_VGND_c_473_n 0.0221535f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_267 N_A_27_47#_c_430_n N_VGND_c_473_n 0.00248202f $X=0.985 $Y=0.82 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_432_n N_A_297_47#_M1005_d 0.00508685f $X=2.16 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_269 N_A_27_47#_M1013_s N_A_297_47#_c_524_n 0.00369694f $X=2.005 $Y=0.235
+ $X2=0 $Y2=0
cc_270 N_A_27_47#_c_430_n N_A_297_47#_c_524_n 0.00799569f $X=0.985 $Y=0.82 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_432_n N_A_297_47#_c_524_n 0.0497861f $X=2.16 $Y=0.38 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_432_n N_A_511_47#_c_547_n 0.0180053f $X=2.16 $Y=0.38 $X2=0
+ $Y2=0
cc_273 N_VGND_c_472_n N_A_297_47#_M1005_d 0.00297142f $X=4.83 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_274 N_VGND_c_472_n N_A_297_47#_M1004_s 0.00256987f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_275 N_VGND_c_471_n N_A_297_47#_c_524_n 0.00358979f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_276 N_VGND_c_472_n N_A_297_47#_c_524_n 0.00905523f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_277 N_VGND_c_472_n N_A_511_47#_M1004_d 0.00308534f $X=4.83 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_278 N_VGND_c_472_n N_A_511_47#_M1010_d 0.0021521f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_279 N_VGND_c_472_n N_A_511_47#_M1008_d 0.00333101f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_280 N_VGND_c_471_n N_A_511_47#_c_547_n 0.0631108f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_281 N_VGND_c_472_n N_A_511_47#_c_547_n 0.0393417f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_282 N_VGND_c_471_n N_A_511_47#_c_553_n 0.0424633f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_283 N_VGND_c_472_n N_A_511_47#_c_553_n 0.0273648f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_284 N_VGND_c_471_n N_A_511_47#_c_549_n 0.0231569f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_285 N_VGND_c_472_n N_A_511_47#_c_549_n 0.0126939f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_286 N_VGND_c_471_n N_A_511_47#_c_576_n 0.0114055f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_287 N_VGND_c_472_n N_A_511_47#_c_576_n 0.00653405f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_288 N_A_297_47#_c_524_n N_A_511_47#_M1004_d 0.00611495f $X=3.22 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_289 N_A_297_47#_M1004_s N_A_511_47#_c_547_n 0.00401386f $X=3.085 $Y=0.235
+ $X2=0 $Y2=0
cc_290 N_A_297_47#_c_524_n N_A_511_47#_c_547_n 0.0514451f $X=3.22 $Y=0.72 $X2=0
+ $Y2=0
