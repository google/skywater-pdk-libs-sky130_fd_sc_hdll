* File: sky130_fd_sc_hdll__nand4_4.pex.spice
* Created: Thu Aug 27 19:14:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND4_4%D 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 37 51 57 60 65
c81 65 0 1.74465e-19 $X=1.615 $Y=1.19
c82 27 0 1.09605e-19 $X=1.93 $Y=0.56
r83 51 52 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.217
+ $X2=1.93 $Y2=1.217
r84 49 51 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=1.67 $Y=1.217
+ $X2=1.905 $Y2=1.217
r85 49 65 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.67
+ $Y=1.16 $X2=1.67 $Y2=1.16
r86 47 49 30.9541 $w=3.27e-07 $l=2.1e-07 $layer=POLY_cond $X=1.46 $Y=1.217
+ $X2=1.67 $Y2=1.217
r87 46 47 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.217
+ $X2=1.46 $Y2=1.217
r88 45 46 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=0.99 $Y=1.217
+ $X2=1.435 $Y2=1.217
r89 44 45 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.217
+ $X2=0.99 $Y2=1.217
r90 43 44 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=0.52 $Y=1.217
+ $X2=0.965 $Y2=1.217
r91 42 43 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.217
+ $X2=0.52 $Y2=1.217
r92 37 42 15.8716 $w=3.27e-07 $l=1.23288e-07 $layer=POLY_cond $X=0.395 $Y=1.165
+ $X2=0.495 $Y2=1.217
r93 37 39 25.7087 $w=2.8e-07 $l=1.2e-07 $layer=POLY_cond $X=0.395 $Y=1.165
+ $X2=0.275 $Y2=1.165
r94 32 65 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=1.595 $Y=1.175
+ $X2=1.615 $Y2=1.175
r95 31 32 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=1.255 $Y=1.175
+ $X2=1.595 $Y2=1.175
r96 31 60 5.54545 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=1.255 $Y=1.175
+ $X2=1.155 $Y2=1.175
r97 30 60 22.7364 $w=1.98e-07 $l=4.1e-07 $layer=LI1_cond $X=0.745 $Y=1.175
+ $X2=1.155 $Y2=1.175
r98 30 57 2.77273 $w=1.98e-07 $l=5e-08 $layer=LI1_cond $X=0.745 $Y=1.175
+ $X2=0.695 $Y2=1.175
r99 29 57 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.695 $Y2=1.175
r100 29 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r101 25 52 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=1.217
r102 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=0.56
r103 22 51 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.217
r104 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r105 18 47 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=1.217
r106 18 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=0.56
r107 15 46 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.217
r108 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r109 11 45 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=1.217
r110 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=0.56
r111 8 44 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.217
r112 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r113 4 43 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=1.217
r114 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=0.56
r115 1 42 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.217
r116 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_4%C 3 5 7 10 12 14 17 19 21 22 24 27 29 30
+ 31 32 49 54 58 60 64
c78 49 0 1.74465e-19 $X=3.785 $Y=1.217
r79 58 60 28.2818 $w=1.98e-07 $l=5.1e-07 $layer=LI1_cond $X=2.825 $Y=1.175
+ $X2=3.335 $Y2=1.175
r80 49 50 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=3.785 $Y=1.217
+ $X2=3.81 $Y2=1.217
r81 48 64 13.5864 $w=1.98e-07 $l=2.45e-07 $layer=LI1_cond $X=3.55 $Y=1.175
+ $X2=3.795 $Y2=1.175
r82 47 49 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=3.55 $Y=1.217
+ $X2=3.785 $Y2=1.217
r83 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.16 $X2=3.55 $Y2=1.16
r84 45 47 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=3.315 $Y=1.217
+ $X2=3.55 $Y2=1.217
r85 44 45 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.217
+ $X2=3.315 $Y2=1.217
r86 43 44 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=2.845 $Y=1.217
+ $X2=3.29 $Y2=1.217
r87 42 43 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.217
+ $X2=2.845 $Y2=1.217
r88 41 54 17.4682 $w=1.98e-07 $l=3.15e-07 $layer=LI1_cond $X=2.605 $Y=1.175
+ $X2=2.29 $Y2=1.175
r89 40 42 31.6911 $w=3.27e-07 $l=2.15e-07 $layer=POLY_cond $X=2.605 $Y=1.217
+ $X2=2.82 $Y2=1.217
r90 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.605
+ $Y=1.16 $X2=2.605 $Y2=1.16
r91 38 40 33.9021 $w=3.27e-07 $l=2.3e-07 $layer=POLY_cond $X=2.375 $Y=1.217
+ $X2=2.605 $Y2=1.217
r92 37 38 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.217
+ $X2=2.375 $Y2=1.217
r93 32 64 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=3.805 $Y=1.175
+ $X2=3.795 $Y2=1.175
r94 31 48 11.3682 $w=1.98e-07 $l=2.05e-07 $layer=LI1_cond $X=3.345 $Y=1.175
+ $X2=3.55 $Y2=1.175
r95 31 60 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=3.345 $Y=1.175
+ $X2=3.335 $Y2=1.175
r96 30 58 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=2.785 $Y=1.175
+ $X2=2.825 $Y2=1.175
r97 30 41 9.98182 $w=1.98e-07 $l=1.8e-07 $layer=LI1_cond $X=2.785 $Y=1.175
+ $X2=2.605 $Y2=1.175
r98 29 54 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=2.275 $Y=1.175
+ $X2=2.29 $Y2=1.175
r99 25 50 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.81 $Y=1.025
+ $X2=3.81 $Y2=1.217
r100 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.81 $Y=1.025
+ $X2=3.81 $Y2=0.56
r101 22 49 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.217
r102 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r103 19 45 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.217
r104 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r105 15 44 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=1.217
r106 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=0.56
r107 12 43 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.217
r108 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r109 8 42 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.82 $Y=1.025
+ $X2=2.82 $Y2=1.217
r110 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.82 $Y=1.025
+ $X2=2.82 $Y2=0.56
r111 5 38 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.217
r112 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r113 1 37 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=1.217
r114 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_4%B 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 37 50 51 56 60 63 66
c79 50 0 1.79329e-19 $X=5.95 $Y=1.16
r80 51 52 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=6.185 $Y=1.217
+ $X2=6.21 $Y2=1.217
r81 50 66 5.54545 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=5.95 $Y=1.175 $X2=5.85
+ $Y2=1.175
r82 49 51 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=5.95 $Y=1.217
+ $X2=6.185 $Y2=1.217
r83 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.95
+ $Y=1.16 $X2=5.95 $Y2=1.16
r84 47 49 30.9541 $w=3.27e-07 $l=2.1e-07 $layer=POLY_cond $X=5.74 $Y=1.217
+ $X2=5.95 $Y2=1.217
r85 46 47 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=5.715 $Y=1.217
+ $X2=5.74 $Y2=1.217
r86 45 46 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=5.27 $Y=1.217
+ $X2=5.715 $Y2=1.217
r87 44 45 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=5.245 $Y=1.217
+ $X2=5.27 $Y2=1.217
r88 43 44 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=4.8 $Y=1.217
+ $X2=5.245 $Y2=1.217
r89 42 43 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=4.775 $Y=1.217
+ $X2=4.8 $Y2=1.217
r90 40 56 6.37727 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=4.51 $Y=1.175
+ $X2=4.395 $Y2=1.175
r91 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.51
+ $Y=1.16 $X2=4.51 $Y2=1.16
r92 37 42 16.3472 $w=3.27e-07 $l=1.253e-07 $layer=POLY_cond $X=4.675 $Y=1.16
+ $X2=4.775 $Y2=1.217
r93 37 39 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.675 $Y=1.16
+ $X2=4.51 $Y2=1.16
r94 32 66 1.83 $w=1.98e-07 $l=3.3e-08 $layer=LI1_cond $X=5.817 $Y=1.175 $X2=5.85
+ $Y2=1.175
r95 32 63 27.8382 $w=1.98e-07 $l=5.02e-07 $layer=LI1_cond $X=5.817 $Y=1.175
+ $X2=5.315 $Y2=1.175
r96 31 63 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=5.305 $Y=1.175
+ $X2=5.315 $Y2=1.175
r97 31 60 24.9545 $w=1.98e-07 $l=4.5e-07 $layer=LI1_cond $X=5.305 $Y=1.175
+ $X2=4.855 $Y2=1.175
r98 30 60 3.32727 $w=1.98e-07 $l=6e-08 $layer=LI1_cond $X=4.795 $Y=1.175
+ $X2=4.855 $Y2=1.175
r99 30 40 15.8045 $w=1.98e-07 $l=2.85e-07 $layer=LI1_cond $X=4.795 $Y=1.175
+ $X2=4.51 $Y2=1.175
r100 29 56 3.32727 $w=1.98e-07 $l=6e-08 $layer=LI1_cond $X=4.335 $Y=1.175
+ $X2=4.395 $Y2=1.175
r101 25 52 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.21 $Y=1.025
+ $X2=6.21 $Y2=1.217
r102 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.21 $Y=1.025
+ $X2=6.21 $Y2=0.56
r103 22 51 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.217
r104 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.985
r105 18 47 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.74 $Y=1.025
+ $X2=5.74 $Y2=1.217
r106 18 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.74 $Y=1.025
+ $X2=5.74 $Y2=0.56
r107 15 46 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.217
r108 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.985
r109 11 45 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.27 $Y=1.025
+ $X2=5.27 $Y2=1.217
r110 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.27 $Y=1.025
+ $X2=5.27 $Y2=0.56
r111 8 44 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.217
r112 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.985
r113 4 43 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.8 $Y=1.025
+ $X2=4.8 $Y2=1.217
r114 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.8 $Y=1.025 $X2=4.8
+ $Y2=0.56
r115 1 42 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.217
r116 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_4%A 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 35 37 54 56 59
c77 35 0 1.79329e-19 $X=8.225 $Y=1.165
r78 54 56 29.9455 $w=1.98e-07 $l=5.4e-07 $layer=LI1_cond $X=7.325 $Y=1.175
+ $X2=7.865 $Y2=1.175
r79 49 50 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=8.1 $Y=1.217
+ $X2=8.125 $Y2=1.217
r80 48 49 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=7.655 $Y=1.217
+ $X2=8.1 $Y2=1.217
r81 47 48 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=7.63 $Y=1.217
+ $X2=7.655 $Y2=1.217
r82 45 47 51.5902 $w=3.27e-07 $l=3.5e-07 $layer=POLY_cond $X=7.28 $Y=1.217
+ $X2=7.63 $Y2=1.217
r83 43 45 14.0031 $w=3.27e-07 $l=9.5e-08 $layer=POLY_cond $X=7.185 $Y=1.217
+ $X2=7.28 $Y2=1.217
r84 42 43 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=7.16 $Y=1.217
+ $X2=7.185 $Y2=1.217
r85 41 42 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=6.715 $Y=1.217
+ $X2=7.16 $Y2=1.217
r86 40 41 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=6.69 $Y=1.217
+ $X2=6.715 $Y2=1.217
r87 37 59 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.345
+ $Y=1.16 $X2=8.345 $Y2=1.16
r88 35 50 15.8716 $w=3.27e-07 $l=1.23288e-07 $layer=POLY_cond $X=8.225 $Y=1.165
+ $X2=8.125 $Y2=1.217
r89 35 37 25.7087 $w=2.8e-07 $l=1.2e-07 $layer=POLY_cond $X=8.225 $Y=1.165
+ $X2=8.345 $Y2=1.165
r90 31 59 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=8.385 $Y=1.175
+ $X2=8.345 $Y2=1.175
r91 30 59 26.0636 $w=1.98e-07 $l=4.7e-07 $layer=LI1_cond $X=7.875 $Y=1.175
+ $X2=8.345 $Y2=1.175
r92 30 56 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=7.875 $Y=1.175
+ $X2=7.865 $Y2=1.175
r93 29 54 2.49545 $w=1.98e-07 $l=4.5e-08 $layer=LI1_cond $X=7.28 $Y=1.175
+ $X2=7.325 $Y2=1.175
r94 29 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.28
+ $Y=1.16 $X2=7.28 $Y2=1.16
r95 26 50 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=8.125 $Y=1.41
+ $X2=8.125 $Y2=1.217
r96 26 28 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.125 $Y=1.41
+ $X2=8.125 $Y2=1.985
r97 22 49 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=8.1 $Y=1.025
+ $X2=8.1 $Y2=1.217
r98 22 24 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.1 $Y=1.025
+ $X2=8.1 $Y2=0.56
r99 19 48 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.655 $Y=1.41
+ $X2=7.655 $Y2=1.217
r100 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.655 $Y=1.41
+ $X2=7.655 $Y2=1.985
r101 15 47 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.63 $Y=1.025
+ $X2=7.63 $Y2=1.217
r102 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.63 $Y=1.025
+ $X2=7.63 $Y2=0.56
r103 12 43 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.185 $Y=1.41
+ $X2=7.185 $Y2=1.217
r104 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.185 $Y=1.41
+ $X2=7.185 $Y2=1.985
r105 8 42 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.16 $Y=1.025
+ $X2=7.16 $Y2=1.217
r106 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.16 $Y=1.025
+ $X2=7.16 $Y2=0.56
r107 5 41 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.715 $Y=1.41
+ $X2=6.715 $Y2=1.217
r108 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.715 $Y=1.41
+ $X2=6.715 $Y2=1.985
r109 1 40 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.69 $Y=1.025
+ $X2=6.69 $Y2=1.217
r110 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.69 $Y=1.025
+ $X2=6.69 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_4%VPWR 1 2 3 4 5 6 7 8 9 28 30 34 38 40 44
+ 48 52 56 60 64 66 68 73 74 76 77 79 80 82 83 84 90 104 112 115 118 122
r139 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r140 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r141 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r142 113 116 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r143 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r144 107 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.51 $Y2=2.72
r145 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r146 104 121 3.9934 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=8.275 $Y=2.72
+ $X2=8.507 $Y2=2.72
r147 104 106 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=8.275 $Y=2.72
+ $X2=8.05 $Y2=2.72
r148 103 107 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r149 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r150 100 103 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r151 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r152 97 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r153 97 119 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.37 $Y2=2.72
r154 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r155 94 118 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=4.28 $Y2=2.72
r156 94 96 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=5.29 $Y2=2.72
r157 93 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r158 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r159 90 118 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=3.935 $Y=2.72
+ $X2=4.28 $Y2=2.72
r160 90 92 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.935 $Y=2.72
+ $X2=3.91 $Y2=2.72
r161 89 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r162 89 116 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r163 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r164 86 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.14 $Y2=2.72
r165 86 88 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.99 $Y2=2.72
r166 84 113 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r167 84 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r168 82 102 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.335 $Y=2.72
+ $X2=7.13 $Y2=2.72
r169 82 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.335 $Y=2.72
+ $X2=7.42 $Y2=2.72
r170 81 106 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=7.505 $Y=2.72
+ $X2=8.05 $Y2=2.72
r171 81 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.505 $Y=2.72
+ $X2=7.42 $Y2=2.72
r172 79 99 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=6.37 $Y=2.72
+ $X2=6.21 $Y2=2.72
r173 79 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.37 $Y=2.72
+ $X2=6.455 $Y2=2.72
r174 78 102 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.54 $Y=2.72
+ $X2=7.13 $Y2=2.72
r175 78 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.54 $Y=2.72
+ $X2=6.455 $Y2=2.72
r176 76 96 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=5.395 $Y=2.72
+ $X2=5.29 $Y2=2.72
r177 76 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=2.72
+ $X2=5.48 $Y2=2.72
r178 75 99 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=5.565 $Y=2.72
+ $X2=6.21 $Y2=2.72
r179 75 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=2.72
+ $X2=5.48 $Y2=2.72
r180 73 88 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.995 $Y=2.72
+ $X2=2.99 $Y2=2.72
r181 73 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=2.72
+ $X2=3.08 $Y2=2.72
r182 72 92 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3.165 $Y=2.72
+ $X2=3.91 $Y2=2.72
r183 72 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=2.72
+ $X2=3.08 $Y2=2.72
r184 68 71 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=8.405 $Y=1.66
+ $X2=8.405 $Y2=2.34
r185 66 121 3.21882 $w=2.6e-07 $l=1.38109e-07 $layer=LI1_cond $X=8.405 $Y=2.635
+ $X2=8.507 $Y2=2.72
r186 66 71 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=8.405 $Y=2.635
+ $X2=8.405 $Y2=2.34
r187 62 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.42 $Y=2.635
+ $X2=7.42 $Y2=2.72
r188 62 64 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.42 $Y=2.635
+ $X2=7.42 $Y2=2
r189 58 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.455 $Y=2.635
+ $X2=6.455 $Y2=2.72
r190 58 60 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.455 $Y=2.635
+ $X2=6.455 $Y2=2
r191 54 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2.72
r192 54 56 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2
r193 50 118 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.28 $Y=2.635
+ $X2=4.28 $Y2=2.72
r194 50 52 11.0074 $w=6.88e-07 $l=6.35e-07 $layer=LI1_cond $X=4.28 $Y=2.635
+ $X2=4.28 $Y2=2
r195 46 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2.72
r196 46 48 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2
r197 42 115 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.72
r198 42 44 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2
r199 41 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=1.2 $Y2=2.72
r200 40 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=2.14 $Y2=2.72
r201 40 41 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=1.285 $Y2=2.72
r202 36 112 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.72
r203 36 38 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r204 35 109 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r205 34 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=1.2 $Y2=2.72
r206 34 35 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=0.345 $Y2=2.72
r207 30 33 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.34
r208 28 109 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r209 28 33 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.34
r210 9 71 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=8.215
+ $Y=1.485 $X2=8.36 $Y2=2.34
r211 9 68 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=8.215
+ $Y=1.485 $X2=8.36 $Y2=1.66
r212 8 64 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=7.275
+ $Y=1.485 $X2=7.42 $Y2=2
r213 7 60 300 $w=1.7e-07 $l=5.98268e-07 $layer=licon1_PDIFF $count=2 $X=6.275
+ $Y=1.485 $X2=6.455 $Y2=2
r214 6 56 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=2
r215 5 52 150 $w=1.7e-07 $l=8.85833e-07 $layer=licon1_PDIFF $count=4 $X=3.875
+ $Y=1.485 $X2=4.54 $Y2=2
r216 4 48 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2
r217 3 44 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r218 2 38 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r219 1 33 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r220 1 30 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_4%Y 1 2 3 4 5 6 7 8 9 10 31 33 35 39 41 45
+ 47 51 53 57 59 63 65 69 71 75 77 79 81 86 88 90 92 94 98 101
c192 71 0 1.70629e-19 $X=6.825 $Y=0.78
r193 96 101 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=6.685 $Y=1.445
+ $X2=6.685 $Y2=1.19
r194 96 98 1.91251 $w=2.8e-07 $l=1.92289e-07 $layer=LI1_cond $X=6.685 $Y=1.445
+ $X2=6.83 $Y2=1.555
r195 95 101 11.7302 $w=2.78e-07 $l=2.85e-07 $layer=LI1_cond $X=6.685 $Y=0.905
+ $X2=6.685 $Y2=1.19
r196 79 100 2.73777 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=7.865 $Y=1.665
+ $X2=7.865 $Y2=1.555
r197 79 81 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=7.865 $Y=1.665
+ $X2=7.865 $Y2=2.34
r198 78 98 4.36787 $w=2.2e-07 $l=2.85e-07 $layer=LI1_cond $X=7.115 $Y=1.555
+ $X2=6.83 $Y2=1.555
r199 77 100 4.72888 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=7.675 $Y=1.555
+ $X2=7.865 $Y2=1.555
r200 77 78 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=7.675 $Y=1.555
+ $X2=7.115 $Y2=1.555
r201 73 75 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=6.95 $Y=0.78
+ $X2=7.89 $Y2=0.78
r202 71 95 6.84494 $w=2.5e-07 $l=1.92614e-07 $layer=LI1_cond $X=6.825 $Y=0.78
+ $X2=6.685 $Y2=0.905
r203 71 73 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.825 $Y=0.78
+ $X2=6.95 $Y2=0.78
r204 67 98 1.91251 $w=3.8e-07 $l=1.50167e-07 $layer=LI1_cond $X=6.925 $Y=1.665
+ $X2=6.83 $Y2=1.555
r205 67 69 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=6.925 $Y=1.665
+ $X2=6.925 $Y2=2.34
r206 66 94 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=6.115 $Y=1.555
+ $X2=5.925 $Y2=1.555
r207 65 98 4.36787 $w=2.2e-07 $l=2.85e-07 $layer=LI1_cond $X=6.545 $Y=1.555
+ $X2=6.83 $Y2=1.555
r208 65 66 22.525 $w=2.18e-07 $l=4.3e-07 $layer=LI1_cond $X=6.545 $Y=1.555
+ $X2=6.115 $Y2=1.555
r209 61 94 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=5.925 $Y=1.665
+ $X2=5.925 $Y2=1.555
r210 61 63 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=5.925 $Y=1.665
+ $X2=5.925 $Y2=2.34
r211 60 92 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=5.175 $Y=1.555
+ $X2=4.985 $Y2=1.555
r212 59 94 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=5.735 $Y=1.555
+ $X2=5.925 $Y2=1.555
r213 59 60 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=5.735 $Y=1.555
+ $X2=5.175 $Y2=1.555
r214 55 92 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=4.985 $Y=1.665
+ $X2=4.985 $Y2=1.555
r215 55 57 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=4.985 $Y=1.665
+ $X2=4.985 $Y2=2.34
r216 54 90 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=3.715 $Y=1.555
+ $X2=3.525 $Y2=1.555
r217 53 92 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=4.795 $Y=1.555
+ $X2=4.985 $Y2=1.555
r218 53 54 56.5745 $w=2.18e-07 $l=1.08e-06 $layer=LI1_cond $X=4.795 $Y=1.555
+ $X2=3.715 $Y2=1.555
r219 49 90 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=3.525 $Y=1.665
+ $X2=3.525 $Y2=1.555
r220 49 51 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=3.525 $Y=1.665
+ $X2=3.525 $Y2=2.34
r221 48 88 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=1.555
+ $X2=2.585 $Y2=1.555
r222 47 90 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=3.335 $Y=1.555
+ $X2=3.525 $Y2=1.555
r223 47 48 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=3.335 $Y=1.555
+ $X2=2.775 $Y2=1.555
r224 43 88 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=2.585 $Y=1.665
+ $X2=2.585 $Y2=1.555
r225 43 45 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=2.585 $Y=1.665
+ $X2=2.585 $Y2=2.34
r226 42 86 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=1.555
+ $X2=1.645 $Y2=1.555
r227 41 88 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=1.555
+ $X2=2.585 $Y2=1.555
r228 41 42 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=2.395 $Y=1.555
+ $X2=1.835 $Y2=1.555
r229 37 86 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.645 $Y2=1.555
r230 37 39 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.645 $Y2=2.34
r231 36 84 4.72888 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=1.555
+ $X2=0.705 $Y2=1.555
r232 35 86 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=1.555
+ $X2=1.645 $Y2=1.555
r233 35 36 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=1.455 $Y=1.555
+ $X2=0.895 $Y2=1.555
r234 31 84 2.73777 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=1.555
r235 31 33 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=2.34
r236 10 100 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=7.745
+ $Y=1.485 $X2=7.89 $Y2=1.66
r237 10 81 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.745
+ $Y=1.485 $X2=7.89 $Y2=2.34
r238 9 98 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=6.805
+ $Y=1.485 $X2=6.95 $Y2=1.66
r239 9 69 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.805
+ $Y=1.485 $X2=6.95 $Y2=2.34
r240 8 94 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=1.66
r241 8 63 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=2.34
r242 7 92 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=1.66
r243 7 57 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=2.34
r244 6 90 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.66
r245 6 51 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2.34
r246 5 88 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.66
r247 5 45 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.34
r248 4 86 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r249 4 39 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
r250 3 84 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r251 3 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r252 2 75 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=7.705
+ $Y=0.235 $X2=7.89 $Y2=0.74
r253 1 73 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=6.765
+ $Y=0.235 $X2=6.95 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_4%A_27_47# 1 2 3 4 5 16 19 20 21 24 30 34 36
r62 32 34 47.0998 $w=2.28e-07 $l=9.4e-07 $layer=LI1_cond $X=3.08 $Y=0.37
+ $X2=4.02 $Y2=0.37
r63 30 32 42.8408 $w=2.28e-07 $l=8.55e-07 $layer=LI1_cond $X=2.225 $Y=0.37
+ $X2=3.08 $Y2=0.37
r64 27 29 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.14 $Y=0.655 $X2=2.14
+ $Y2=0.625
r65 26 30 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.14 $Y=0.485
+ $X2=2.225 $Y2=0.37
r66 26 29 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.14 $Y=0.485
+ $X2=2.14 $Y2=0.625
r67 25 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=0.78 $X2=1.2
+ $Y2=0.78
r68 24 27 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.055 $Y=0.78
+ $X2=2.14 $Y2=0.655
r69 24 25 35.4952 $w=2.48e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=0.78
+ $X2=1.285 $Y2=0.78
r70 21 36 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.2 $Y=0.655 $X2=1.2
+ $Y2=0.78
r71 21 23 2.15294 $w=1.7e-07 $l=3e-08 $layer=LI1_cond $X=1.2 $Y=0.655 $X2=1.2
+ $Y2=0.625
r72 19 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0.78 $X2=1.2
+ $Y2=0.78
r73 19 20 35.4952 $w=2.48e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=0.78
+ $X2=0.345 $Y2=0.78
r74 16 20 6.81736 $w=2.5e-07 $l=1.79956e-07 $layer=LI1_cond $X=0.217 $Y=0.655
+ $X2=0.345 $Y2=0.78
r75 16 18 1.43529 $w=2.55e-07 $l=3e-08 $layer=LI1_cond $X=0.217 $Y=0.655
+ $X2=0.217 $Y2=0.625
r76 5 34 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.235 $X2=4.02 $Y2=0.4
r77 4 32 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.4
r78 3 29 182 $w=1.7e-07 $l=4.52493e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.625
r79 2 23 182 $w=1.7e-07 $l=4.52493e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.625
r80 1 18 182 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_4%VGND 1 2 9 13 15 17 22 32 33 36 39
r87 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r88 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r89 32 33 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r90 30 33 1.83245 $w=4.8e-07 $l=6.44e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=8.51
+ $Y2=0
r91 30 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r92 29 32 420.15 $w=1.68e-07 $l=6.44e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=8.51
+ $Y2=0
r93 29 30 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r94 27 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=1.645
+ $Y2=0
r95 27 29 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=2.07
+ $Y2=0
r96 26 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r97 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r98 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r99 23 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r100 23 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r101 22 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.645
+ $Y2=0
r102 22 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r103 17 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r104 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r105 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r106 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r107 11 39 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=0.085
+ $X2=1.645 $Y2=0
r108 11 13 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=1.645 $Y=0.085
+ $X2=1.645 $Y2=0.4
r109 7 36 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r110 7 9 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.4
r111 2 13 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.4
r112 1 9 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_4%A_485_47# 1 2 3 4 21
c33 21 0 1.09605e-19 $X=5.95 $Y=0.74
r34 19 21 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=5.01 $Y=0.78
+ $X2=5.95 $Y2=0.78
r35 17 19 67.3027 $w=2.48e-07 $l=1.46e-06 $layer=LI1_cond $X=3.55 $Y=0.78
+ $X2=5.01 $Y2=0.78
r36 14 17 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=2.61 $Y=0.78
+ $X2=3.55 $Y2=0.78
r37 4 21 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=5.815
+ $Y=0.235 $X2=5.95 $Y2=0.74
r38 3 19 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.875
+ $Y=0.235 $X2=5.01 $Y2=0.74
r39 2 17 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.74
r40 1 14 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_4%A_883_47# 1 2 3 4 5 16 26 28
r39 26 31 3.25045 $w=2.55e-07 $l=1.15e-07 $layer=LI1_cond $X=8.402 $Y=0.485
+ $X2=8.402 $Y2=0.37
r40 26 28 11.5244 $w=2.53e-07 $l=2.55e-07 $layer=LI1_cond $X=8.402 $Y=0.485
+ $X2=8.402 $Y2=0.74
r41 23 25 48.3525 $w=2.28e-07 $l=9.65e-07 $layer=LI1_cond $X=6.455 $Y=0.37
+ $X2=7.42 $Y2=0.37
r42 21 23 48.8536 $w=2.28e-07 $l=9.75e-07 $layer=LI1_cond $X=5.48 $Y=0.37
+ $X2=6.455 $Y2=0.37
r43 18 21 47.0998 $w=2.28e-07 $l=9.4e-07 $layer=LI1_cond $X=4.54 $Y=0.37
+ $X2=5.48 $Y2=0.37
r44 16 31 3.58963 $w=2.3e-07 $l=1.27e-07 $layer=LI1_cond $X=8.275 $Y=0.37
+ $X2=8.402 $Y2=0.37
r45 16 25 42.8408 $w=2.28e-07 $l=8.55e-07 $layer=LI1_cond $X=8.275 $Y=0.37
+ $X2=7.42 $Y2=0.37
r46 5 31 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=8.175
+ $Y=0.235 $X2=8.36 $Y2=0.4
r47 5 28 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=8.175
+ $Y=0.235 $X2=8.36 $Y2=0.74
r48 4 25 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=7.235
+ $Y=0.235 $X2=7.42 $Y2=0.4
r49 3 23 182 $w=1.7e-07 $l=2.38642e-07 $layer=licon1_NDIFF $count=1 $X=6.285
+ $Y=0.235 $X2=6.455 $Y2=0.4
r50 2 21 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.345
+ $Y=0.235 $X2=5.48 $Y2=0.4
r51 1 18 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=4.415
+ $Y=0.235 $X2=4.54 $Y2=0.4
.ends

