# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__mux2_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  10.58000 BY  2.720000 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.580000 0.645000 7.495000 0.815000 ;
        RECT 5.580000 0.815000 5.800000 1.325000 ;
        RECT 5.755000 0.425000 6.390000 0.645000 ;
        RECT 7.325000 0.815000 7.495000 0.995000 ;
        RECT 7.325000 0.995000 7.845000 1.165000 ;
        RECT 7.625000 1.165000 7.845000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.620000 1.075000 4.960000 1.120000 ;
        RECT 4.620000 1.120000 9.115000 1.260000 ;
        RECT 4.620000 1.260000 4.960000 1.305000 ;
        RECT 8.765000 1.075000 9.115000 1.120000 ;
        RECT 8.765000 1.260000 9.115000 1.305000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 6.110000 1.415000  6.400000 1.460000 ;
        RECT 6.110000 1.460000 10.035000 1.600000 ;
        RECT 6.110000 1.600000  6.400000 1.645000 ;
        RECT 9.745000 1.415000 10.035000 1.460000 ;
        RECT 9.745000 1.600000 10.035000 1.645000 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  2.024500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.255000 0.815000 0.635000 ;
        RECT 0.605000 0.635000 3.635000 0.805000 ;
        RECT 0.605000 0.805000 0.865000 1.575000 ;
        RECT 0.605000 1.575000 3.635000 1.745000 ;
        RECT 0.605000 1.745000 0.815000 2.465000 ;
        RECT 1.585000 0.295000 1.755000 0.635000 ;
        RECT 1.585000 1.745000 1.755000 2.465000 ;
        RECT 2.525000 0.255000 2.695000 0.635000 ;
        RECT 2.525000 1.745000 2.695000 2.465000 ;
        RECT 3.465000 0.295000 3.635000 0.635000 ;
        RECT 3.465000 1.745000 3.635000 2.465000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.580000 0.085000 ;
      RECT  0.000000  2.635000 10.580000 2.805000 ;
      RECT  0.090000  0.085000  0.425000 0.465000 ;
      RECT  0.090000  1.915000  0.425000 2.635000 ;
      RECT  0.985000  0.085000  1.365000 0.465000 ;
      RECT  0.985000  1.915000  1.365000 2.635000 ;
      RECT  1.085000  1.075000  3.975000 1.245000 ;
      RECT  1.925000  0.085000  2.305000 0.465000 ;
      RECT  1.925000  1.915000  2.305000 2.635000 ;
      RECT  2.865000  0.085000  3.245000 0.465000 ;
      RECT  2.865000  1.915000  3.245000 2.635000 ;
      RECT  3.805000  0.085000  4.185000 0.465000 ;
      RECT  3.805000  0.635000  5.340000 0.805000 ;
      RECT  3.805000  0.805000  3.975000 1.075000 ;
      RECT  3.805000  1.245000  3.975000 1.835000 ;
      RECT  3.805000  1.835000  8.975000 2.005000 ;
      RECT  3.805000  2.255000  4.185000 2.635000 ;
      RECT  4.145000  0.995000  4.365000 1.495000 ;
      RECT  4.145000  1.495000  6.585000 1.665000 ;
      RECT  4.355000  0.295000  5.525000 0.465000 ;
      RECT  4.630000  2.255000  6.405000 2.425000 ;
      RECT  4.690000  1.105000  4.925000 1.275000 ;
      RECT  4.705000  0.995000  4.925000 1.105000 ;
      RECT  4.705000  1.275000  4.925000 1.325000 ;
      RECT  5.170000  0.805000  5.340000 0.935000 ;
      RECT  6.170000  0.995000  6.585000 1.495000 ;
      RECT  6.660000  0.085000  6.990000 0.465000 ;
      RECT  6.675000  2.175000  6.845000 2.635000 ;
      RECT  6.895000  0.995000  7.115000 1.495000 ;
      RECT  6.895000  1.495000  9.635000 1.665000 ;
      RECT  7.030000  2.255000  9.445000 2.425000 ;
      RECT  7.175000  0.295000  8.565000 0.465000 ;
      RECT  7.715000  0.635000  8.370000 0.805000 ;
      RECT  8.150000  0.805000  8.370000 0.935000 ;
      RECT  8.885000  0.995000  9.170000 1.325000 ;
      RECT  9.415000  0.645000 10.385000 0.815000 ;
      RECT  9.415000  0.815000  9.635000 1.495000 ;
      RECT  9.415000  1.665000  9.635000 1.915000 ;
      RECT  9.415000  1.915000 10.385000 2.085000 ;
      RECT  9.665000  0.085000 10.045000 0.465000 ;
      RECT  9.665000  2.255000 10.045000 2.635000 ;
      RECT  9.805000  0.995000 10.235000 1.615000 ;
      RECT 10.215000  0.295000 10.385000 0.645000 ;
      RECT 10.215000  1.795000 10.385000 1.915000 ;
      RECT 10.215000  2.085000 10.385000 2.465000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.690000  1.105000  4.860000 1.275000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.170000  0.765000  5.340000 0.935000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.170000  1.445000  6.340000 1.615000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.150000  0.765000  8.320000 0.935000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  1.105000  9.055000 1.275000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  1.445000  9.975000 1.615000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
    LAYER met1 ;
      RECT 5.110000 0.735000 5.400000 0.780000 ;
      RECT 5.110000 0.780000 8.430000 0.920000 ;
      RECT 5.110000 0.920000 5.400000 0.965000 ;
      RECT 8.090000 0.735000 8.430000 0.780000 ;
      RECT 8.090000 0.920000 8.430000 0.965000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2_8
END LIBRARY
