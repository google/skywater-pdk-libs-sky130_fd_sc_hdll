* File: sky130_fd_sc_hdll__o32ai_2.pxi.spice
* Created: Thu Aug 27 19:22:53 2020
* 
x_PM_SKY130_FD_SC_HDLL__O32AI_2%B2 N_B2_c_87_n N_B2_M1003_g N_B2_c_91_n
+ N_B2_M1001_g N_B2_c_92_n N_B2_M1007_g N_B2_c_88_n N_B2_M1019_g B2 B2
+ N_B2_c_89_n B2 PM_SKY130_FD_SC_HDLL__O32AI_2%B2
x_PM_SKY130_FD_SC_HDLL__O32AI_2%B1 N_B1_c_125_n N_B1_M1005_g N_B1_c_129_n
+ N_B1_M1012_g N_B1_c_130_n N_B1_M1018_g N_B1_c_126_n N_B1_M1013_g B1 B1
+ N_B1_c_128_n B1 PM_SKY130_FD_SC_HDLL__O32AI_2%B1
x_PM_SKY130_FD_SC_HDLL__O32AI_2%A3 N_A3_M1014_g N_A3_c_178_n N_A3_c_179_n
+ N_A3_c_183_n N_A3_M1002_g N_A3_c_180_n N_A3_M1016_g N_A3_c_184_n N_A3_M1015_g
+ A3 N_A3_c_181_n N_A3_c_182_n A3 PM_SKY130_FD_SC_HDLL__O32AI_2%A3
x_PM_SKY130_FD_SC_HDLL__O32AI_2%A2 N_A2_c_234_n N_A2_M1000_g N_A2_c_238_n
+ N_A2_M1009_g N_A2_c_235_n N_A2_M1008_g N_A2_c_239_n N_A2_M1011_g A2 A2
+ N_A2_c_236_n A2 PM_SKY130_FD_SC_HDLL__O32AI_2%A2
x_PM_SKY130_FD_SC_HDLL__O32AI_2%A1 N_A1_c_280_n N_A1_M1004_g N_A1_c_284_n
+ N_A1_M1006_g N_A1_c_281_n N_A1_M1017_g N_A1_c_285_n N_A1_M1010_g A1 A1 A1
+ N_A1_c_283_n A1 A1 PM_SKY130_FD_SC_HDLL__O32AI_2%A1
x_PM_SKY130_FD_SC_HDLL__O32AI_2%A_27_297# N_A_27_297#_M1001_d
+ N_A_27_297#_M1007_d N_A_27_297#_M1018_d N_A_27_297#_c_319_n
+ N_A_27_297#_c_320_n N_A_27_297#_c_323_n N_A_27_297#_c_326_n
+ N_A_27_297#_c_327_n N_A_27_297#_c_329_n N_A_27_297#_c_321_n
+ PM_SKY130_FD_SC_HDLL__O32AI_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__O32AI_2%Y N_Y_M1003_s N_Y_M1005_d N_Y_M1001_s
+ N_Y_M1002_d N_Y_c_364_n N_Y_c_372_n N_Y_c_366_n N_Y_c_373_n N_Y_c_398_n Y Y
+ PM_SKY130_FD_SC_HDLL__O32AI_2%Y
x_PM_SKY130_FD_SC_HDLL__O32AI_2%VPWR N_VPWR_M1012_s N_VPWR_M1006_d
+ N_VPWR_M1010_d N_VPWR_c_443_n N_VPWR_c_444_n N_VPWR_c_445_n N_VPWR_c_446_n
+ N_VPWR_c_447_n N_VPWR_c_448_n VPWR N_VPWR_c_449_n N_VPWR_c_450_n
+ N_VPWR_c_451_n N_VPWR_c_442_n PM_SKY130_FD_SC_HDLL__O32AI_2%VPWR
x_PM_SKY130_FD_SC_HDLL__O32AI_2%A_525_297# N_A_525_297#_M1002_s
+ N_A_525_297#_M1015_s N_A_525_297#_M1011_d N_A_525_297#_c_523_n
+ N_A_525_297#_c_524_n N_A_525_297#_c_527_n N_A_525_297#_c_529_n
+ N_A_525_297#_c_531_n N_A_525_297#_c_525_n N_A_525_297#_c_526_n
+ N_A_525_297#_c_555_n PM_SKY130_FD_SC_HDLL__O32AI_2%A_525_297#
x_PM_SKY130_FD_SC_HDLL__O32AI_2%A_807_297# N_A_807_297#_M1009_s
+ N_A_807_297#_M1006_s N_A_807_297#_c_565_n N_A_807_297#_c_575_n
+ N_A_807_297#_c_579_n N_A_807_297#_c_568_n
+ PM_SKY130_FD_SC_HDLL__O32AI_2%A_807_297#
x_PM_SKY130_FD_SC_HDLL__O32AI_2%A_27_47# N_A_27_47#_M1003_d N_A_27_47#_M1019_d
+ N_A_27_47#_M1013_s N_A_27_47#_M1016_d N_A_27_47#_M1008_s N_A_27_47#_M1017_s
+ N_A_27_47#_c_598_n N_A_27_47#_c_599_n N_A_27_47#_c_609_n N_A_27_47#_c_615_n
+ N_A_27_47#_c_600_n N_A_27_47#_c_601_n N_A_27_47#_c_622_n N_A_27_47#_c_602_n
+ N_A_27_47#_c_603_n N_A_27_47#_c_604_n N_A_27_47#_c_605_n N_A_27_47#_c_606_n
+ PM_SKY130_FD_SC_HDLL__O32AI_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__O32AI_2%VGND N_VGND_M1014_s N_VGND_M1000_d
+ N_VGND_M1004_d N_VGND_c_691_n N_VGND_c_692_n N_VGND_c_693_n N_VGND_c_694_n
+ N_VGND_c_695_n N_VGND_c_696_n N_VGND_c_697_n VGND N_VGND_c_698_n
+ N_VGND_c_699_n N_VGND_c_700_n N_VGND_c_701_n
+ PM_SKY130_FD_SC_HDLL__O32AI_2%VGND
cc_1 VNB N_B2_c_87_n 0.02229f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_B2_c_88_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB N_B2_c_89_n 0.0419878f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_4 VNB B2 0.0135148f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_5 VNB N_B1_c_125_n 0.0169097f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_6 VNB N_B1_c_126_n 0.0163996f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_7 VNB B1 0.00315088f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_8 VNB N_B1_c_128_n 0.0355875f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_9 VNB N_A3_M1014_g 0.0287142f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_10 VNB N_A3_c_178_n 0.0328699f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_11 VNB N_A3_c_179_n 0.00849829f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_12 VNB N_A3_c_180_n 0.0217006f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_13 VNB N_A3_c_181_n 0.00301463f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.16
cc_14 VNB N_A3_c_182_n 0.0437797f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_15 VNB N_A2_c_234_n 0.0169324f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_16 VNB N_A2_c_235_n 0.0224149f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_17 VNB N_A2_c_236_n 0.0446644f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_18 VNB A2 0.00999544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A1_c_280_n 0.0216895f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_20 VNB N_A1_c_281_n 0.0218012f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_21 VNB A1 0.0156584f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A1_c_283_n 0.053288f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.2
cc_23 VNB N_Y_c_364_n 0.00851249f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_24 VNB Y 0.00266127f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_442_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_598_n 0.0100703f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.202
cc_27 VNB N_A_27_47#_c_599_n 0.0183982f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.16
cc_28 VNB N_A_27_47#_c_600_n 0.00445219f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_27_47#_c_601_n 0.00194411f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_27_47#_c_602_n 0.0153368f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_603_n 0.0180521f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_27_47#_c_604_n 0.00484878f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_27_47#_c_605_n 0.00305374f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_27_47#_c_606_n 0.00822315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_691_n 0.00592343f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_36 VNB N_VGND_c_692_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_693_n 4.89699e-19 $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.16
cc_38 VNB N_VGND_c_694_n 0.0195627f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.202
cc_39 VNB N_VGND_c_695_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.2
cc_40 VNB N_VGND_c_696_n 0.0273833f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_697_n 0.00503156f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.2
cc_42 VNB N_VGND_c_698_n 0.0678694f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_699_n 0.0195271f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_700_n 0.316851f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_701_n 0.00728035f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VPB N_B2_c_91_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_47 VPB N_B2_c_92_n 0.016445f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_48 VPB N_B2_c_89_n 0.0224377f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_49 VPB B2 0.00503392f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.19
cc_50 VPB N_B1_c_129_n 0.0164409f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_51 VPB N_B1_c_130_n 0.0196266f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_52 VPB B1 0.00252951f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_53 VPB N_B1_c_128_n 0.0204811f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_54 VPB N_A3_c_183_n 0.0197335f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_55 VPB N_A3_c_184_n 0.016445f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_56 VPB N_A3_c_181_n 0.00249044f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.16
cc_57 VPB N_A3_c_182_n 0.020726f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_58 VPB N_A2_c_238_n 0.016445f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_59 VPB N_A2_c_239_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_60 VPB N_A2_c_236_n 0.0255797f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_61 VPB A2 0.00489897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A1_c_284_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_63 VPB N_A1_c_285_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_64 VPB A1 0.00641694f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A1_c_283_n 0.0276468f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.2
cc_66 VPB N_A_27_297#_c_319_n 0.00753428f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_67 VPB N_A_27_297#_c_320_n 0.0305647f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_68 VPB N_A_27_297#_c_321_n 0.00718079f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.2
cc_69 VPB N_Y_c_366_n 0.0118291f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.202
cc_70 VPB Y 0.0065524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_443_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_72 VPB N_VPWR_c_444_n 0.0049401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_445_n 0.011989f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_74 VPB N_VPWR_c_446_n 0.00502493f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.16
cc_75 VPB N_VPWR_c_447_n 0.0809579f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_448_n 0.00391723f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_449_n 0.0393666f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.19
cc_78 VPB N_VPWR_c_450_n 0.0212818f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_451_n 0.0032427f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_442_n 0.0692154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_525_297#_c_523_n 0.00230104f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_82 VPB N_A_525_297#_c_524_n 0.0046399f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_83 VPB N_A_525_297#_c_525_n 0.00212461f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_84 VPB N_A_525_297#_c_526_n 0.00433313f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.2
cc_85 VPB N_A_807_297#_c_565_n 0.0133368f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_86 N_B2_c_88_n N_B1_c_125_n 0.0247014f $X=0.99 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_87 N_B2_c_92_n N_B1_c_129_n 0.0243056f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_88 N_B2_c_89_n B1 0.00267209f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_89 B2 B1 0.0209934f $X=0.695 $Y=1.19 $X2=0 $Y2=0
cc_90 N_B2_c_89_n N_B1_c_128_n 0.0247014f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_91 B2 N_A_27_297#_c_320_n 0.0215753f $X=0.695 $Y=1.19 $X2=0 $Y2=0
cc_92 N_B2_c_91_n N_A_27_297#_c_323_n 0.0123313f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_93 N_B2_c_92_n N_A_27_297#_c_323_n 0.0111735f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_94 N_B2_c_87_n N_Y_c_364_n 0.0038241f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_95 N_B2_c_88_n N_Y_c_364_n 0.0125545f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_96 N_B2_c_89_n N_Y_c_364_n 0.00472855f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_97 B2 N_Y_c_364_n 0.0287109f $X=0.695 $Y=1.19 $X2=0 $Y2=0
cc_98 N_B2_c_92_n N_Y_c_372_n 0.0131951f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_99 N_B2_c_91_n N_Y_c_373_n 0.0107257f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_100 N_B2_c_92_n N_Y_c_373_n 0.00707269f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_101 N_B2_c_89_n N_Y_c_373_n 0.00629709f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_102 B2 N_Y_c_373_n 0.0251217f $X=0.695 $Y=1.19 $X2=0 $Y2=0
cc_103 N_B2_c_91_n N_VPWR_c_449_n 0.00429453f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_104 N_B2_c_92_n N_VPWR_c_449_n 0.00429453f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_105 N_B2_c_91_n N_VPWR_c_442_n 0.00697643f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_106 N_B2_c_92_n N_VPWR_c_442_n 0.00609021f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_107 N_B2_c_87_n N_A_27_47#_c_599_n 4.62114e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_108 B2 N_A_27_47#_c_599_n 0.0218655f $X=0.695 $Y=1.19 $X2=0 $Y2=0
cc_109 N_B2_c_87_n N_A_27_47#_c_609_n 0.0115551f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_110 N_B2_c_88_n N_A_27_47#_c_609_n 0.00994068f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_111 B2 N_A_27_47#_c_609_n 0.00389697f $X=0.695 $Y=1.19 $X2=0 $Y2=0
cc_112 N_B2_c_87_n N_VGND_c_698_n 0.00357877f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_113 N_B2_c_88_n N_VGND_c_698_n 0.00357877f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_114 N_B2_c_87_n N_VGND_c_700_n 0.006431f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_115 N_B2_c_88_n N_VGND_c_700_n 0.005504f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_116 N_B1_c_126_n N_A3_M1014_g 0.01859f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_117 N_B1_c_128_n N_A3_c_179_n 0.01859f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_118 N_B1_c_128_n N_A3_c_181_n 3.12012e-19 $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_119 N_B1_c_129_n N_A_27_297#_c_323_n 0.00215639f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_120 N_B1_c_129_n N_A_27_297#_c_326_n 5.78668e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_121 N_B1_c_129_n N_A_27_297#_c_327_n 0.00450227f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_122 N_B1_c_130_n N_A_27_297#_c_327_n 4.63737e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_123 N_B1_c_129_n N_A_27_297#_c_329_n 0.0107484f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_124 N_B1_c_130_n N_A_27_297#_c_329_n 0.00797545f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_125 N_B1_c_129_n N_A_27_297#_c_321_n 5.48372e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_126 N_B1_c_130_n N_A_27_297#_c_321_n 0.0102842f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_127 N_B1_c_125_n N_Y_c_364_n 0.0106952f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_128 N_B1_c_126_n N_Y_c_364_n 0.011473f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_129 B1 N_Y_c_364_n 0.0573809f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_130 N_B1_c_128_n N_Y_c_364_n 0.00472855f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_131 N_B1_c_129_n N_Y_c_372_n 0.0118662f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_132 N_B1_c_130_n N_Y_c_372_n 0.0115212f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_133 B1 N_Y_c_372_n 0.0469226f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_134 N_B1_c_128_n N_Y_c_372_n 0.00616252f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_135 N_B1_c_129_n N_Y_c_373_n 7.20922e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_136 N_B1_c_125_n Y 4.11928e-19 $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_137 N_B1_c_126_n Y 0.00245966f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_138 B1 Y 0.0198794f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_139 N_B1_c_128_n Y 0.0107911f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_140 N_B1_c_129_n Y 3.79936e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_141 N_B1_c_130_n Y 0.00768207f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_142 N_B1_c_128_n Y 0.00495892f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_143 N_B1_c_129_n N_VPWR_c_443_n 0.00402381f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_144 N_B1_c_130_n N_VPWR_c_443_n 0.00398422f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_145 N_B1_c_130_n N_VPWR_c_447_n 0.00489481f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_146 N_B1_c_129_n N_VPWR_c_449_n 0.00513275f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_147 N_B1_c_129_n N_VPWR_c_442_n 0.00680962f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_148 N_B1_c_130_n N_VPWR_c_442_n 0.00778876f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_149 N_B1_c_125_n N_A_27_47#_c_609_n 0.00994068f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_150 N_B1_c_126_n N_A_27_47#_c_609_n 0.00993988f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_151 N_B1_c_125_n N_VGND_c_698_n 0.00357877f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_152 N_B1_c_126_n N_VGND_c_698_n 0.00357877f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_153 N_B1_c_125_n N_VGND_c_700_n 0.005504f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_154 N_B1_c_126_n N_VGND_c_700_n 0.005504f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A3_c_180_n N_A2_c_234_n 0.0124239f $X=3.44 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_156 N_A3_c_184_n N_A2_c_238_n 0.0100726f $X=3.475 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A3_c_181_n N_A2_c_236_n 2.09263e-19 $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A3_c_182_n N_A2_c_236_n 0.0278816f $X=3.44 $Y=1.202 $X2=0 $Y2=0
cc_159 N_A3_c_181_n A2 0.012753f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A3_c_182_n A2 0.0024903f $X=3.44 $Y=1.202 $X2=0 $Y2=0
cc_161 N_A3_M1014_g N_Y_c_364_n 0.00118111f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_162 N_A3_c_178_n N_Y_c_366_n 0.00142437f $X=2.905 $Y=1.19 $X2=0 $Y2=0
cc_163 N_A3_c_179_n N_Y_c_366_n 0.00770918f $X=2.425 $Y=1.19 $X2=0 $Y2=0
cc_164 N_A3_c_183_n N_Y_c_366_n 0.0102325f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A3_c_181_n N_Y_c_366_n 0.0253615f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A3_c_183_n N_Y_c_398_n 0.01493f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A3_c_184_n N_Y_c_398_n 0.00765949f $X=3.475 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A3_c_181_n N_Y_c_398_n 0.0228639f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A3_c_182_n N_Y_c_398_n 0.00601902f $X=3.44 $Y=1.202 $X2=0 $Y2=0
cc_170 N_A3_M1014_g Y 0.00786068f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_171 N_A3_c_179_n Y 0.0078945f $X=2.425 $Y=1.19 $X2=0 $Y2=0
cc_172 N_A3_c_181_n Y 0.01359f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A3_c_182_n Y 2.59064e-19 $X=3.44 $Y=1.202 $X2=0 $Y2=0
cc_174 N_A3_c_183_n Y 0.00218873f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A3_c_182_n Y 0.00229257f $X=3.44 $Y=1.202 $X2=0 $Y2=0
cc_176 N_A3_c_183_n N_VPWR_c_447_n 0.00434439f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A3_c_184_n N_VPWR_c_447_n 0.00434439f $X=3.475 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A3_c_183_n N_VPWR_c_442_n 0.00735385f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A3_c_184_n N_VPWR_c_442_n 0.00609671f $X=3.475 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A3_c_183_n N_A_525_297#_c_527_n 0.0110966f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A3_c_184_n N_A_525_297#_c_527_n 0.0146153f $X=3.475 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A3_M1014_g N_A_27_47#_c_609_n 0.0139835f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_183 N_A3_M1014_g N_A_27_47#_c_615_n 0.00790593f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_184 N_A3_c_178_n N_A_27_47#_c_600_n 0.00160685f $X=2.905 $Y=1.19 $X2=0 $Y2=0
cc_185 N_A3_c_180_n N_A_27_47#_c_600_n 0.00980487f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A3_c_181_n N_A_27_47#_c_600_n 0.0536568f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A3_c_182_n N_A_27_47#_c_600_n 0.0121659f $X=3.44 $Y=1.202 $X2=0 $Y2=0
cc_188 N_A3_M1014_g N_A_27_47#_c_601_n 0.00461232f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_189 N_A3_c_178_n N_A_27_47#_c_601_n 0.0041434f $X=2.905 $Y=1.19 $X2=0 $Y2=0
cc_190 N_A3_c_180_n N_A_27_47#_c_622_n 0.0131252f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A3_c_180_n N_A_27_47#_c_604_n 0.00571033f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A3_c_182_n N_A_27_47#_c_604_n 0.0030994f $X=3.44 $Y=1.202 $X2=0 $Y2=0
cc_193 N_A3_M1014_g N_VGND_c_691_n 0.00397473f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_194 N_A3_c_180_n N_VGND_c_691_n 0.0109709f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A3_c_180_n N_VGND_c_694_n 0.00395968f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A3_M1014_g N_VGND_c_698_n 0.00357877f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_197 N_A3_M1014_g N_VGND_c_700_n 0.00662944f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_198 N_A3_c_180_n N_VGND_c_700_n 0.00699801f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A2_c_236_n A1 8.76878e-19 $X=4.38 $Y=1.202 $X2=0 $Y2=0
cc_200 A2 A1 0.0167879f $X=4.375 $Y=1.19 $X2=0 $Y2=0
cc_201 A2 N_A1_c_283_n 0.00167207f $X=4.375 $Y=1.19 $X2=0 $Y2=0
cc_202 N_A2_c_239_n N_VPWR_c_444_n 0.00225336f $X=4.415 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A2_c_238_n N_VPWR_c_447_n 0.00434439f $X=3.945 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A2_c_239_n N_VPWR_c_447_n 0.00434439f $X=4.415 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A2_c_238_n N_VPWR_c_442_n 0.00609671f $X=3.945 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A2_c_239_n N_VPWR_c_442_n 0.00735385f $X=4.415 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A2_c_236_n N_A_525_297#_c_529_n 2.45159e-19 $X=4.38 $Y=1.202 $X2=0
+ $Y2=0
cc_208 A2 N_A_525_297#_c_529_n 0.00625213f $X=4.375 $Y=1.19 $X2=0 $Y2=0
cc_209 N_A2_c_238_n N_A_525_297#_c_531_n 0.0146153f $X=3.945 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A2_c_239_n N_A_525_297#_c_531_n 0.0117706f $X=4.415 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A2_c_239_n N_A_807_297#_c_565_n 0.0130606f $X=4.415 $Y=1.41 $X2=0 $Y2=0
cc_212 A2 N_A_807_297#_c_565_n 0.0416135f $X=4.375 $Y=1.19 $X2=0 $Y2=0
cc_213 N_A2_c_238_n N_A_807_297#_c_568_n 0.00740338f $X=3.945 $Y=1.41 $X2=0
+ $Y2=0
cc_214 N_A2_c_239_n N_A_807_297#_c_568_n 0.0113557f $X=4.415 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A2_c_236_n N_A_807_297#_c_568_n 0.006374f $X=4.38 $Y=1.202 $X2=0 $Y2=0
cc_216 A2 N_A_807_297#_c_568_n 0.0212256f $X=4.375 $Y=1.19 $X2=0 $Y2=0
cc_217 N_A2_c_234_n N_A_27_47#_c_622_n 0.00707713f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A2_c_235_n N_A_27_47#_c_622_n 8.10277e-19 $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A2_c_234_n N_A_27_47#_c_604_n 0.00115517f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_220 A2 N_A_27_47#_c_604_n 0.0079569f $X=4.375 $Y=1.19 $X2=0 $Y2=0
cc_221 N_A2_c_234_n N_A_27_47#_c_605_n 0.00952594f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A2_c_235_n N_A_27_47#_c_605_n 0.0158078f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A2_c_236_n N_A_27_47#_c_605_n 0.00646614f $X=4.38 $Y=1.202 $X2=0 $Y2=0
cc_224 A2 N_A_27_47#_c_605_n 0.0866535f $X=4.375 $Y=1.19 $X2=0 $Y2=0
cc_225 N_A2_c_234_n N_VGND_c_692_n 0.00382269f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A2_c_235_n N_VGND_c_692_n 0.00412745f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A2_c_234_n N_VGND_c_694_n 0.00422241f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A2_c_235_n N_VGND_c_696_n 0.00436487f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A2_c_234_n N_VGND_c_700_n 0.00608884f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A2_c_235_n N_VGND_c_700_n 0.00764859f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A1_c_284_n N_VPWR_c_444_n 0.00713502f $X=5.425 $Y=1.41 $X2=0 $Y2=0
cc_232 N_A1_c_285_n N_VPWR_c_446_n 0.00844976f $X=5.895 $Y=1.41 $X2=0 $Y2=0
cc_233 A1 N_VPWR_c_446_n 0.0185234f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_234 N_A1_c_284_n N_VPWR_c_450_n 0.0067375f $X=5.425 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A1_c_285_n N_VPWR_c_450_n 0.0067375f $X=5.895 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A1_c_284_n N_VPWR_c_442_n 0.0131263f $X=5.425 $Y=1.41 $X2=0 $Y2=0
cc_237 N_A1_c_285_n N_VPWR_c_442_n 0.0127987f $X=5.895 $Y=1.41 $X2=0 $Y2=0
cc_238 N_A1_c_284_n N_A_807_297#_c_565_n 0.0157914f $X=5.425 $Y=1.41 $X2=0 $Y2=0
cc_239 A1 N_A_807_297#_c_565_n 0.0190075f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_240 N_A1_c_283_n N_A_807_297#_c_565_n 0.00200573f $X=5.79 $Y=1.202 $X2=0
+ $Y2=0
cc_241 N_A1_c_284_n N_A_807_297#_c_575_n 5.79575e-19 $X=5.425 $Y=1.41 $X2=0
+ $Y2=0
cc_242 N_A1_c_285_n N_A_807_297#_c_575_n 0.00238098f $X=5.895 $Y=1.41 $X2=0
+ $Y2=0
cc_243 A1 N_A_807_297#_c_575_n 0.0214226f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_244 N_A1_c_283_n N_A_807_297#_c_575_n 0.00667391f $X=5.79 $Y=1.202 $X2=0
+ $Y2=0
cc_245 N_A1_c_284_n N_A_807_297#_c_579_n 0.0151916f $X=5.425 $Y=1.41 $X2=0 $Y2=0
cc_246 N_A1_c_285_n N_A_807_297#_c_579_n 0.00995715f $X=5.895 $Y=1.41 $X2=0
+ $Y2=0
cc_247 N_A1_c_280_n N_A_27_47#_c_602_n 0.0150457f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A1_c_281_n N_A_27_47#_c_602_n 0.014871f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_249 A1 N_A_27_47#_c_602_n 0.0841107f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_250 N_A1_c_283_n N_A_27_47#_c_602_n 0.00735634f $X=5.79 $Y=1.202 $X2=0 $Y2=0
cc_251 N_A1_c_281_n N_A_27_47#_c_603_n 0.0130837f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A1_c_280_n N_A_27_47#_c_606_n 0.0142899f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A1_c_280_n N_VGND_c_693_n 0.0102068f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A1_c_281_n N_VGND_c_693_n 0.00935559f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A1_c_280_n N_VGND_c_696_n 0.00319306f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_256 N_A1_c_281_n N_VGND_c_699_n 0.00377504f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_257 N_A1_c_280_n N_VGND_c_700_n 0.00522424f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_258 N_A1_c_281_n N_VGND_c_700_n 0.00557352f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A_27_297#_c_323_n N_Y_M1001_s 0.003659f $X=1.115 $Y=2.38 $X2=0 $Y2=0
cc_260 N_A_27_297#_M1007_d N_Y_c_372_n 0.0037145f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_261 N_A_27_297#_c_323_n N_Y_c_372_n 0.00367045f $X=1.115 $Y=2.38 $X2=0 $Y2=0
cc_262 N_A_27_297#_c_326_n N_Y_c_372_n 0.0154597f $X=1.24 $Y=2.005 $X2=0 $Y2=0
cc_263 N_A_27_297#_c_329_n N_Y_c_372_n 0.0310164f $X=1.925 $Y=1.92 $X2=0 $Y2=0
cc_264 N_A_27_297#_c_321_n N_Y_c_372_n 0.00450177f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_265 N_A_27_297#_c_320_n N_Y_c_373_n 0.0467908f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_266 N_A_27_297#_c_323_n N_Y_c_373_n 0.0168436f $X=1.115 $Y=2.38 $X2=0 $Y2=0
cc_267 N_A_27_297#_c_326_n N_Y_c_373_n 0.0116213f $X=1.24 $Y=2.005 $X2=0 $Y2=0
cc_268 N_A_27_297#_c_327_n N_Y_c_373_n 0.00563756f $X=1.24 $Y=2.295 $X2=0 $Y2=0
cc_269 N_A_27_297#_M1018_d Y 0.00315008f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_270 N_A_27_297#_c_321_n Y 0.0234735f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_271 N_A_27_297#_c_329_n N_VPWR_M1012_s 0.00341225f $X=1.925 $Y=1.92 $X2=-0.19
+ $Y2=1.305
cc_272 N_A_27_297#_c_323_n N_VPWR_c_443_n 0.0109394f $X=1.115 $Y=2.38 $X2=0
+ $Y2=0
cc_273 N_A_27_297#_c_327_n N_VPWR_c_443_n 0.00708316f $X=1.24 $Y=2.295 $X2=0
+ $Y2=0
cc_274 N_A_27_297#_c_329_n N_VPWR_c_443_n 0.0131159f $X=1.925 $Y=1.92 $X2=0
+ $Y2=0
cc_275 N_A_27_297#_c_321_n N_VPWR_c_443_n 0.0209034f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_276 N_A_27_297#_c_329_n N_VPWR_c_447_n 0.00198891f $X=1.925 $Y=1.92 $X2=0
+ $Y2=0
cc_277 N_A_27_297#_c_321_n N_VPWR_c_447_n 0.0228567f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_278 N_A_27_297#_c_319_n N_VPWR_c_449_n 0.0179936f $X=0.217 $Y=2.295 $X2=0
+ $Y2=0
cc_279 N_A_27_297#_c_323_n N_VPWR_c_449_n 0.056947f $X=1.115 $Y=2.38 $X2=0 $Y2=0
cc_280 N_A_27_297#_c_329_n N_VPWR_c_449_n 0.00267292f $X=1.925 $Y=1.92 $X2=0
+ $Y2=0
cc_281 N_A_27_297#_M1001_d N_VPWR_c_442_n 0.00217523f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_282 N_A_27_297#_M1007_d N_VPWR_c_442_n 0.00231266f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_283 N_A_27_297#_M1018_d N_VPWR_c_442_n 0.00217852f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_284 N_A_27_297#_c_319_n N_VPWR_c_442_n 0.0098205f $X=0.217 $Y=2.295 $X2=0
+ $Y2=0
cc_285 N_A_27_297#_c_323_n N_VPWR_c_442_n 0.036323f $X=1.115 $Y=2.38 $X2=0 $Y2=0
cc_286 N_A_27_297#_c_329_n N_VPWR_c_442_n 0.00968081f $X=1.925 $Y=1.92 $X2=0
+ $Y2=0
cc_287 N_A_27_297#_c_321_n N_VPWR_c_442_n 0.0140629f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_288 N_A_27_297#_c_321_n N_A_525_297#_c_523_n 0.0119856f $X=2.14 $Y=2 $X2=0
+ $Y2=0
cc_289 N_A_27_297#_c_321_n N_A_525_297#_c_524_n 0.0249272f $X=2.14 $Y=2 $X2=0
+ $Y2=0
cc_290 N_Y_c_372_n N_VPWR_M1012_s 0.00326319f $X=1.985 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_291 N_Y_M1001_s N_VPWR_c_442_n 0.00232895f $X=0.585 $Y=1.485 $X2=0 $Y2=0
cc_292 N_Y_M1002_d N_VPWR_c_442_n 0.00233833f $X=3.095 $Y=1.485 $X2=0 $Y2=0
cc_293 N_Y_c_366_n N_A_525_297#_M1002_s 0.00586325f $X=3.025 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_294 N_Y_c_366_n N_A_525_297#_c_524_n 0.0201185f $X=3.025 $Y=1.58 $X2=0 $Y2=0
cc_295 N_Y_c_398_n N_A_525_297#_c_524_n 0.0176241f $X=3.24 $Y=1.66 $X2=0 $Y2=0
cc_296 N_Y_M1002_d N_A_525_297#_c_527_n 0.00361015f $X=3.095 $Y=1.485 $X2=0
+ $Y2=0
cc_297 N_Y_c_366_n N_A_525_297#_c_527_n 0.00331741f $X=3.025 $Y=1.58 $X2=0 $Y2=0
cc_298 N_Y_c_398_n N_A_525_297#_c_527_n 0.0197169f $X=3.24 $Y=1.66 $X2=0 $Y2=0
cc_299 N_Y_c_398_n N_A_525_297#_c_529_n 0.0366157f $X=3.24 $Y=1.66 $X2=0 $Y2=0
cc_300 N_Y_c_364_n N_A_27_47#_M1019_d 0.00162409f $X=1.985 $Y=0.78 $X2=0 $Y2=0
cc_301 N_Y_c_364_n N_A_27_47#_M1013_s 0.00207431f $X=1.985 $Y=0.78 $X2=0 $Y2=0
cc_302 N_Y_c_364_n N_A_27_47#_c_599_n 0.01117f $X=1.985 $Y=0.78 $X2=0 $Y2=0
cc_303 N_Y_M1003_s N_A_27_47#_c_609_n 0.00508491f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_304 N_Y_M1005_d N_A_27_47#_c_609_n 0.00508491f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_305 N_Y_c_364_n N_A_27_47#_c_609_n 0.0934304f $X=1.985 $Y=0.78 $X2=0 $Y2=0
cc_306 Y N_A_27_47#_c_609_n 0.00299102f $X=2 $Y=1.105 $X2=0 $Y2=0
cc_307 N_Y_c_398_n N_A_27_47#_c_600_n 7.74003e-19 $X=3.24 $Y=1.66 $X2=0 $Y2=0
cc_308 N_Y_c_364_n N_A_27_47#_c_601_n 0.00735544f $X=1.985 $Y=0.78 $X2=0 $Y2=0
cc_309 N_Y_c_366_n N_A_27_47#_c_601_n 0.00590606f $X=3.025 $Y=1.58 $X2=0 $Y2=0
cc_310 N_Y_M1003_s N_VGND_c_700_n 0.00297142f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_311 N_Y_M1005_d N_VGND_c_700_n 0.00297142f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_312 N_VPWR_c_442_n N_A_525_297#_M1002_s 0.00234829f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_313 N_VPWR_c_442_n N_A_525_297#_M1015_s 0.00232182f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_314 N_VPWR_c_442_n N_A_525_297#_M1011_d 0.00234829f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_447_n N_A_525_297#_c_523_n 0.0155085f $X=5.07 $Y=2.72 $X2=0
+ $Y2=0
cc_316 N_VPWR_c_442_n N_A_525_297#_c_523_n 0.00950669f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_317 N_VPWR_c_447_n N_A_525_297#_c_527_n 0.038255f $X=5.07 $Y=2.72 $X2=0 $Y2=0
cc_318 N_VPWR_c_442_n N_A_525_297#_c_527_n 0.0273315f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_319 N_VPWR_c_447_n N_A_525_297#_c_531_n 0.038255f $X=5.07 $Y=2.72 $X2=0 $Y2=0
cc_320 N_VPWR_c_442_n N_A_525_297#_c_531_n 0.0273315f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_321 N_VPWR_c_444_n N_A_525_297#_c_525_n 0.0126677f $X=5.19 $Y=2 $X2=0 $Y2=0
cc_322 N_VPWR_c_447_n N_A_525_297#_c_525_n 0.0155085f $X=5.07 $Y=2.72 $X2=0
+ $Y2=0
cc_323 N_VPWR_c_442_n N_A_525_297#_c_525_n 0.00950669f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_324 N_VPWR_c_444_n N_A_525_297#_c_526_n 0.0256957f $X=5.19 $Y=2 $X2=0 $Y2=0
cc_325 N_VPWR_c_447_n N_A_525_297#_c_555_n 0.0105923f $X=5.07 $Y=2.72 $X2=0
+ $Y2=0
cc_326 N_VPWR_c_442_n N_A_525_297#_c_555_n 0.00648411f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_327 N_VPWR_c_442_n N_A_807_297#_M1009_s 0.00233833f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_328 N_VPWR_c_442_n N_A_807_297#_M1006_s 0.00231418f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_329 N_VPWR_M1006_d N_A_807_297#_c_565_n 0.00660326f $X=5.065 $Y=1.485 $X2=0
+ $Y2=0
cc_330 N_VPWR_c_444_n N_A_807_297#_c_565_n 0.0165158f $X=5.19 $Y=2 $X2=0 $Y2=0
cc_331 N_VPWR_c_446_n N_A_807_297#_c_575_n 0.0111411f $X=6.15 $Y=1.66 $X2=0
+ $Y2=0
cc_332 N_VPWR_c_444_n N_A_807_297#_c_579_n 0.0383726f $X=5.19 $Y=2 $X2=0 $Y2=0
cc_333 N_VPWR_c_446_n N_A_807_297#_c_579_n 0.0490403f $X=6.15 $Y=1.66 $X2=0
+ $Y2=0
cc_334 N_VPWR_c_450_n N_A_807_297#_c_579_n 0.0183657f $X=6.045 $Y=2.72 $X2=0
+ $Y2=0
cc_335 N_VPWR_c_442_n N_A_807_297#_c_579_n 0.0122834f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_336 N_A_525_297#_c_531_n N_A_807_297#_M1009_s 0.00361015f $X=4.585 $Y=2.35
+ $X2=-0.19 $Y2=1.305
cc_337 N_A_525_297#_M1011_d N_A_807_297#_c_565_n 0.00617683f $X=4.505 $Y=1.485
+ $X2=0 $Y2=0
cc_338 N_A_525_297#_c_531_n N_A_807_297#_c_565_n 0.0045407f $X=4.585 $Y=2.35
+ $X2=0 $Y2=0
cc_339 N_A_525_297#_c_526_n N_A_807_297#_c_565_n 0.0201185f $X=4.67 $Y=2 $X2=0
+ $Y2=0
cc_340 N_A_525_297#_c_529_n N_A_807_297#_c_568_n 0.0363365f $X=3.71 $Y=1.66
+ $X2=0 $Y2=0
cc_341 N_A_525_297#_c_531_n N_A_807_297#_c_568_n 0.0161319f $X=4.585 $Y=2.35
+ $X2=0 $Y2=0
cc_342 N_A_525_297#_c_526_n N_A_807_297#_c_568_n 0.0145781f $X=4.67 $Y=2 $X2=0
+ $Y2=0
cc_343 N_A_525_297#_c_529_n N_A_27_47#_c_604_n 0.00349481f $X=3.71 $Y=1.66 $X2=0
+ $Y2=0
cc_344 N_A_807_297#_c_565_n N_A_27_47#_c_606_n 0.0092242f $X=5.495 $Y=1.58 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_609_n N_VGND_M1014_s 0.00512461f $X=2.485 $Y=0.37 $X2=-0.19
+ $Y2=-0.24
cc_346 N_A_27_47#_c_615_n N_VGND_M1014_s 0.0105002f $X=2.57 $Y=0.715 $X2=-0.19
+ $Y2=-0.24
cc_347 N_A_27_47#_c_600_n N_VGND_M1014_s 0.0140685f $X=3.435 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_348 N_A_27_47#_c_601_n N_VGND_M1014_s 0.0032492f $X=2.655 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_349 N_A_27_47#_c_605_n N_VGND_M1000_d 0.00348106f $X=4.505 $Y=0.58 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_602_n N_VGND_M1004_d 0.00214118f $X=5.975 $Y=0.81 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_609_n N_VGND_c_691_n 0.0166143f $X=2.485 $Y=0.37 $X2=0 $Y2=0
cc_352 N_A_27_47#_c_615_n N_VGND_c_691_n 0.00386676f $X=2.57 $Y=0.715 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_600_n N_VGND_c_691_n 0.029725f $X=3.435 $Y=0.81 $X2=0 $Y2=0
cc_354 N_A_27_47#_c_622_n N_VGND_c_691_n 0.0215442f $X=3.65 $Y=0.38 $X2=0 $Y2=0
cc_355 N_A_27_47#_c_622_n N_VGND_c_692_n 0.0177507f $X=3.65 $Y=0.38 $X2=0 $Y2=0
cc_356 N_A_27_47#_c_605_n N_VGND_c_692_n 0.0132111f $X=4.505 $Y=0.58 $X2=0 $Y2=0
cc_357 N_A_27_47#_c_602_n N_VGND_c_693_n 0.0203868f $X=5.975 $Y=0.81 $X2=0 $Y2=0
cc_358 N_A_27_47#_c_603_n N_VGND_c_693_n 0.0174574f $X=6.14 $Y=0.38 $X2=0 $Y2=0
cc_359 N_A_27_47#_c_606_n N_VGND_c_693_n 0.0230311f $X=5.175 $Y=0.58 $X2=0 $Y2=0
cc_360 N_A_27_47#_c_600_n N_VGND_c_694_n 0.00226786f $X=3.435 $Y=0.81 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_622_n N_VGND_c_694_n 0.0222529f $X=3.65 $Y=0.38 $X2=0 $Y2=0
cc_362 N_A_27_47#_c_605_n N_VGND_c_694_n 0.00273345f $X=4.505 $Y=0.58 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_602_n N_VGND_c_696_n 0.00214783f $X=5.975 $Y=0.81 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_605_n N_VGND_c_696_n 0.00355041f $X=4.505 $Y=0.58 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_606_n N_VGND_c_696_n 0.0464092f $X=5.175 $Y=0.58 $X2=0 $Y2=0
cc_366 N_A_27_47#_c_598_n N_VGND_c_698_n 0.0176918f $X=0.217 $Y=0.485 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_609_n N_VGND_c_698_n 0.132122f $X=2.485 $Y=0.37 $X2=0 $Y2=0
cc_368 N_A_27_47#_c_600_n N_VGND_c_698_n 0.00318662f $X=3.435 $Y=0.81 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_602_n N_VGND_c_699_n 0.00301904f $X=5.975 $Y=0.81 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_c_603_n N_VGND_c_699_n 0.0230421f $X=6.14 $Y=0.38 $X2=0 $Y2=0
cc_371 N_A_27_47#_M1003_d N_VGND_c_700_n 0.00209324f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_372 N_A_27_47#_M1019_d N_VGND_c_700_n 0.00215227f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_373 N_A_27_47#_M1013_s N_VGND_c_700_n 0.00215227f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_M1016_d N_VGND_c_700_n 0.00215201f $X=3.515 $Y=0.235 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_M1008_s N_VGND_c_700_n 0.00699525f $X=4.455 $Y=0.235 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_M1017_s N_VGND_c_700_n 0.00377139f $X=5.865 $Y=0.235 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_c_598_n N_VGND_c_700_n 0.00980895f $X=0.217 $Y=0.485 $X2=0
+ $Y2=0
cc_378 N_A_27_47#_c_609_n N_VGND_c_700_n 0.0829814f $X=2.485 $Y=0.37 $X2=0 $Y2=0
cc_379 N_A_27_47#_c_600_n N_VGND_c_700_n 0.0118937f $X=3.435 $Y=0.81 $X2=0 $Y2=0
cc_380 N_A_27_47#_c_622_n N_VGND_c_700_n 0.0139016f $X=3.65 $Y=0.38 $X2=0 $Y2=0
cc_381 N_A_27_47#_c_602_n N_VGND_c_700_n 0.0115433f $X=5.975 $Y=0.81 $X2=0 $Y2=0
cc_382 N_A_27_47#_c_603_n N_VGND_c_700_n 0.0126169f $X=6.14 $Y=0.38 $X2=0 $Y2=0
cc_383 N_A_27_47#_c_605_n N_VGND_c_700_n 0.0132079f $X=4.505 $Y=0.58 $X2=0 $Y2=0
cc_384 N_A_27_47#_c_606_n N_VGND_c_700_n 0.0257581f $X=5.175 $Y=0.58 $X2=0 $Y2=0
