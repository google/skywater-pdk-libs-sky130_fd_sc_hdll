* File: sky130_fd_sc_hdll__a31o_1.pex.spice
* Created: Wed Sep  2 08:19:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A31O_1%A_80_21# 1 2 7 9 10 12 14 15 16 17 27 30 35
+ 36
r78 35 36 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=1.91
+ $X2=2.92 $Y2=1.825
r79 30 32 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=2.315 $Y=0.4
+ $X2=2.315 $Y2=0.74
r80 24 27 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=0.54 $Y=1.16
+ $X2=0.73 $Y2=1.16
r81 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.54
+ $Y=1.16 $X2=0.54 $Y2=1.16
r82 21 36 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=3 $Y=0.825 $X2=3
+ $Y2=1.825
r83 18 32 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.505 $Y=0.74
+ $X2=2.315 $Y2=0.74
r84 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.915 $Y=0.74
+ $X2=3 $Y2=0.825
r85 17 18 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.915 $Y=0.74
+ $X2=2.505 $Y2=0.74
r86 15 32 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.125 $Y=0.74
+ $X2=2.315 $Y2=0.74
r87 15 16 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=2.125 $Y=0.74
+ $X2=0.815 $Y2=0.74
r88 14 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=0.995
+ $X2=0.73 $Y2=1.16
r89 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.73 $Y=0.825
+ $X2=0.815 $Y2=0.74
r90 13 14 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.73 $Y=0.825
+ $X2=0.73 $Y2=0.995
r91 10 25 47.8775 $w=2.99e-07 $l=2.79285e-07 $layer=POLY_cond $X=0.5 $Y=1.41
+ $X2=0.562 $Y2=1.16
r92 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.985
r93 7 25 38.5562 $w=2.99e-07 $l=2.03912e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.562 $Y2=1.16
r94 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=0.56
r95 2 35 300 $w=1.7e-07 $l=5.17446e-07 $layer=licon1_PDIFF $count=2 $X=2.715
+ $Y=1.485 $X2=2.92 $Y2=1.91
r96 1 30 91 $w=1.7e-07 $l=2.64953e-07 $layer=licon1_NDIFF $count=2 $X=2.145
+ $Y=0.235 $X2=2.34 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_1%A3 1 3 4 6 7 8
c32 7 0 1.20528e-19 $X=1.155 $Y=1.19
c33 1 0 1.13706e-19 $X=1.01 $Y=0.995
r34 8 21 8.91512 $w=2.63e-07 $l=2.05e-07 $layer=LI1_cond $X=1.207 $Y=1.53
+ $X2=1.207 $Y2=1.325
r35 7 21 6.12224 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=1.162 $Y=1.16
+ $X2=1.162 $Y2=1.325
r36 7 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.07
+ $Y=1.16 $X2=1.07 $Y2=1.16
r37 4 12 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=1.035 $Y=1.41
+ $X2=1.095 $Y2=1.16
r38 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.035 $Y=1.41
+ $X2=1.035 $Y2=1.985
r39 1 12 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.095 $Y2=1.16
r40 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.01 $Y=0.995 $X2=1.01
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_1%A2 1 3 4 6 7 8
r28 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6 $Y=1.16
+ $X2=1.6 $Y2=1.16
r29 7 8 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.665 $Y=1.53
+ $X2=1.665 $Y2=1.16
r30 4 12 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=1.565 $Y=1.41
+ $X2=1.625 $Y2=1.16
r31 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.565 $Y=1.41
+ $X2=1.565 $Y2=1.985
r32 1 12 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.54 $Y=0.995
+ $X2=1.625 $Y2=1.16
r33 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.54 $Y=0.995 $X2=1.54
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_1%A1 1 3 4 6 7 8
r29 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.16 $X2=2.13 $Y2=1.16
r30 7 8 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.13 $Y=1.53 $X2=2.13
+ $Y2=1.16
r31 4 12 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.095 $Y=1.41
+ $X2=2.155 $Y2=1.16
r32 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.095 $Y=1.41
+ $X2=2.095 $Y2=1.985
r33 1 12 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.07 $Y=0.995
+ $X2=2.155 $Y2=1.16
r34 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.07 $Y=0.995 $X2=2.07
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_1%B1 1 3 4 6 7 8 13
r25 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.66
+ $Y=1.16 $X2=2.66 $Y2=1.16
r26 7 8 13.061 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=2.595 $Y=1.19 $X2=2.595
+ $Y2=1.53
r27 7 13 1.15244 $w=2.98e-07 $l=3e-08 $layer=LI1_cond $X=2.595 $Y=1.19 $X2=2.595
+ $Y2=1.16
r28 4 12 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.625 $Y=1.41
+ $X2=2.685 $Y2=1.16
r29 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.625 $Y=1.41
+ $X2=2.625 $Y2=1.985
r30 1 12 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.6 $Y=0.995
+ $X2=2.685 $Y2=1.16
r31 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.6 $Y=0.995 $X2=2.6
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_1%X 1 2 10 13 14 15 16 17 22
c22 10 0 1.13706e-19 $X=0.26 $Y=0.81
r23 17 31 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.26 $Y=2.21
+ $X2=0.26 $Y2=2.34
r24 16 17 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.26 $Y=1.87
+ $X2=0.26 $Y2=2.21
r25 15 22 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.51
+ $X2=0.26 $Y2=0.385
r26 13 14 5.02519 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=1.575
r27 11 16 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.26 $Y=1.74
+ $X2=0.26 $Y2=1.87
r28 11 13 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.26 $Y=1.74 $X2=0.26
+ $Y2=1.66
r29 10 14 44.6555 $w=1.88e-07 $l=7.65e-07 $layer=LI1_cond $X=0.19 $Y=0.81
+ $X2=0.19 $Y2=1.575
r30 9 15 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.26 $Y=0.645
+ $X2=0.26 $Y2=0.51
r31 9 10 7.81899 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.26 $Y=0.645
+ $X2=0.26 $Y2=0.81
r32 2 31 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r33 2 13 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r34 1 22 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_1%VPWR 1 2 11 17 20 21 22 32 33 36 39
r42 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r44 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 29 32 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r46 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r47 27 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r48 27 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r49 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r50 24 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.77 $Y2=2.72
r51 24 26 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r52 22 37 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r53 22 39 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r54 20 26 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.665 $Y=2.72
+ $X2=1.61 $Y2=2.72
r55 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.665 $Y=2.72
+ $X2=1.83 $Y2=2.72
r56 19 29 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=1.995 $Y=2.72
+ $X2=2.07 $Y2=2.72
r57 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.995 $Y=2.72
+ $X2=1.83 $Y2=2.72
r58 15 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.83 $Y=2.635
+ $X2=1.83 $Y2=2.72
r59 15 17 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=1.83 $Y=2.635
+ $X2=1.83 $Y2=2.25
r60 11 14 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.77 $Y=1.66
+ $X2=0.77 $Y2=2.34
r61 9 36 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=2.635
+ $X2=0.77 $Y2=2.72
r62 9 14 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.77 $Y=2.635
+ $X2=0.77 $Y2=2.34
r63 2 17 600 $w=1.7e-07 $l=8.47998e-07 $layer=licon1_PDIFF $count=1 $X=1.655
+ $Y=1.485 $X2=1.83 $Y2=2.25
r64 1 14 400 $w=1.7e-07 $l=9.40705e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.485 $X2=0.77 $Y2=2.34
r65 1 11 400 $w=1.7e-07 $l=2.52785e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.485 $X2=0.77 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_1%A_225_297# 1 2 7 9 11 13 15
r23 13 20 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.4 $Y=1.995 $X2=2.4
+ $Y2=1.91
r24 13 15 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=2.4 $Y=1.995
+ $X2=2.4 $Y2=2.25
r25 12 18 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.385 $Y=1.91
+ $X2=1.235 $Y2=1.91
r26 11 20 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.275 $Y=1.91
+ $X2=2.4 $Y2=1.91
r27 11 12 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=2.275 $Y=1.91
+ $X2=1.385 $Y2=1.91
r28 7 18 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=1.995 $X2=1.235
+ $Y2=1.91
r29 7 9 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=1.235 $Y=1.995
+ $X2=1.235 $Y2=2.25
r30 2 20 600 $w=1.7e-07 $l=5.04975e-07 $layer=licon1_PDIFF $count=1 $X=2.185
+ $Y=1.485 $X2=2.36 $Y2=1.91
r31 2 15 600 $w=1.7e-07 $l=8.47998e-07 $layer=licon1_PDIFF $count=1 $X=2.185
+ $Y=1.485 $X2=2.36 $Y2=2.25
r32 1 18 600 $w=1.7e-07 $l=5.04975e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.3 $Y2=1.91
r33 1 9 600 $w=1.7e-07 $l=8.47998e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.3 $Y2=2.25
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_1%VGND 1 2 9 11 13 15 17 22 31 35
r44 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r45 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r46 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r47 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r48 26 29 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r49 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r50 25 28 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r51 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r52 23 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.77
+ $Y2=0
r53 23 25 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.15
+ $Y2=0
r54 22 34 4.63344 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.972
+ $Y2=0
r55 22 28 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.53
+ $Y2=0
r56 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.77
+ $Y2=0
r57 17 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.23
+ $Y2=0
r58 15 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r59 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r60 11 34 3.13273 $w=3.3e-07 $l=1.19143e-07 $layer=LI1_cond $X=2.89 $Y=0.085
+ $X2=2.972 $Y2=0
r61 11 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.89 $Y=0.085
+ $X2=2.89 $Y2=0.4
r62 7 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=0.085 $X2=0.77
+ $Y2=0
r63 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.77 $Y=0.085
+ $X2=0.77 $Y2=0.4
r64 2 13 182 $w=1.7e-07 $l=2.85832e-07 $layer=licon1_NDIFF $count=1 $X=2.675
+ $Y=0.235 $X2=2.89 $Y2=0.4
r65 1 9 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.77 $Y2=0.4
.ends

