* File: sky130_fd_sc_hdll__inputiso0p_1.pxi.spice
* Created: Thu Aug 27 19:08:36 2020
* 
x_PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%SLEEP N_SLEEP_c_57_n N_SLEEP_c_58_n
+ N_SLEEP_M1001_g N_SLEEP_M1005_g SLEEP SLEEP SLEEP N_SLEEP_c_56_n
+ PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%SLEEP
x_PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%A_27_413# N_A_27_413#_M1005_d
+ N_A_27_413#_M1001_s N_A_27_413#_c_87_n N_A_27_413#_c_95_n N_A_27_413#_M1006_g
+ N_A_27_413#_c_88_n N_A_27_413#_M1007_g N_A_27_413#_c_96_n N_A_27_413#_c_97_n
+ N_A_27_413#_c_98_n N_A_27_413#_c_90_n N_A_27_413#_c_91_n N_A_27_413#_c_92_n
+ N_A_27_413#_c_93_n PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%A_27_413#
x_PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%A N_A_c_159_n N_A_M1002_g N_A_M1000_g A
+ N_A_c_162_n A PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%A
x_PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%A_211_413# N_A_211_413#_M1007_s
+ N_A_211_413#_M1006_d N_A_211_413#_c_196_n N_A_211_413#_M1004_g
+ N_A_211_413#_c_197_n N_A_211_413#_M1003_g N_A_211_413#_c_202_n
+ N_A_211_413#_c_198_n N_A_211_413#_c_199_n N_A_211_413#_c_200_n
+ N_A_211_413#_c_218_n PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%A_211_413#
x_PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%VPWR N_VPWR_M1001_d N_VPWR_M1002_d
+ N_VPWR_c_253_n VPWR N_VPWR_c_254_n N_VPWR_c_255_n N_VPWR_c_252_n
+ N_VPWR_c_257_n N_VPWR_c_258_n N_VPWR_c_259_n
+ PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%VPWR
x_PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%X N_X_M1003_d N_X_M1004_d X X X N_X_c_292_n
+ PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%X
x_PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%VGND N_VGND_M1005_s N_VGND_M1000_d
+ N_VGND_c_307_n N_VGND_c_308_n N_VGND_c_309_n VGND N_VGND_c_310_n
+ N_VGND_c_311_n N_VGND_c_312_n N_VGND_c_313_n
+ PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%VGND
cc_1 VNB N_SLEEP_M1005_g 0.0380335f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB SLEEP 0.0246847f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_SLEEP_c_56_n 0.0350009f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_4 VNB N_A_27_413#_c_87_n 0.0108642f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_5 VNB N_A_27_413#_c_88_n 0.0237194f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_6 VNB N_A_27_413#_M1007_g 0.0210777f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.16
cc_7 VNB N_A_27_413#_c_90_n 0.0075685f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_413#_c_91_n 0.00191082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_413#_c_92_n 0.00550201f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_413#_c_93_n 0.0302858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_M1000_g 0.0484972f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_12 VNB N_A_211_413#_c_196_n 0.0292536f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_13 VNB N_A_211_413#_c_197_n 0.0208714f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_14 VNB N_A_211_413#_c_198_n 0.00495488f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_15 VNB N_A_211_413#_c_199_n 0.0131351f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=0.995
cc_16 VNB N_A_211_413#_c_200_n 0.0116189f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=0.85
cc_17 VNB N_VPWR_c_252_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB X 0.0297395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_X_c_292_n 0.0265499f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_307_n 0.0114894f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_21 VNB N_VGND_c_308_n 0.0211579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_309_n 0.00562936f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_310_n 0.0468447f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_24 VNB N_VGND_c_311_n 0.0239286f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.16
cc_25 VNB N_VGND_c_312_n 0.187736f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.19
cc_26 VNB N_VGND_c_313_n 0.00632082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VPB N_SLEEP_c_57_n 0.041336f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_28 VPB N_SLEEP_c_58_n 0.0256797f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_29 VPB SLEEP 0.0149437f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_30 VPB N_SLEEP_c_56_n 0.007518f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_31 VPB N_A_27_413#_c_87_n 0.0328248f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_32 VPB N_A_27_413#_c_95_n 0.0223898f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A_27_413#_c_96_n 0.00219961f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.325
cc_34 VPB N_A_27_413#_c_97_n 0.00539927f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_27_413#_c_98_n 0.0110178f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_27_413#_c_91_n 0.00393863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_c_159_n 0.0213926f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_38 VPB N_A_M1000_g 0.0173323f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_39 VPB A 0.0034319f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_40 VPB N_A_c_162_n 0.0622039f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_41 VPB N_A_211_413#_c_196_n 0.0370091f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_42 VPB N_A_211_413#_c_202_n 0.0137569f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_211_413#_c_199_n 0.00965832f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=0.995
cc_44 VPB N_A_211_413#_c_200_n 0.0136504f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=0.85
cc_45 VPB N_VPWR_c_253_n 4.21319e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_254_n 0.015299f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_255_n 0.0261914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_252_n 0.0492213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_257_n 0.00503094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_258_n 0.0178886f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_259_n 0.0221134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB X 0.0437541f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_53 VPB N_X_c_292_n 0.0139685f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 SLEEP N_A_27_413#_c_87_n 3.52543e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_55 N_SLEEP_c_56_n N_A_27_413#_c_87_n 0.0174017f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_56 N_SLEEP_c_57_n N_A_27_413#_c_95_n 0.0174017f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_57 N_SLEEP_c_58_n N_A_27_413#_c_95_n 0.009997f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_58 N_SLEEP_c_58_n N_A_27_413#_c_96_n 0.00550801f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_59 N_SLEEP_c_57_n N_A_27_413#_c_97_n 0.0126367f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_60 N_SLEEP_c_58_n N_A_27_413#_c_97_n 0.00996415f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_61 SLEEP N_A_27_413#_c_97_n 0.00808417f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_62 SLEEP N_A_27_413#_c_98_n 0.0158932f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_63 N_SLEEP_c_56_n N_A_27_413#_c_98_n 6.27406e-19 $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_64 N_SLEEP_M1005_g N_A_27_413#_c_90_n 0.00565159f $X=0.52 $Y=0.445 $X2=0
+ $Y2=0
cc_65 SLEEP N_A_27_413#_c_90_n 0.00287744f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_66 SLEEP N_A_27_413#_c_91_n 0.0326308f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_67 N_SLEEP_c_56_n N_A_27_413#_c_91_n 0.0083556f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_68 N_SLEEP_M1005_g N_A_27_413#_c_92_n 0.00288066f $X=0.52 $Y=0.445 $X2=0
+ $Y2=0
cc_69 SLEEP N_A_27_413#_c_92_n 0.0246147f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_70 N_SLEEP_M1005_g N_A_27_413#_c_93_n 0.0174017f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_71 N_SLEEP_c_58_n N_VPWR_c_253_n 0.0129428f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_72 N_SLEEP_c_58_n N_VPWR_c_254_n 0.00321743f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_73 N_SLEEP_c_58_n N_VPWR_c_252_n 0.00482954f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_74 N_SLEEP_M1005_g N_VGND_c_308_n 0.00511692f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_75 SLEEP N_VGND_c_308_n 0.0225521f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_76 N_SLEEP_c_56_n N_VGND_c_308_n 0.0010017f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_77 N_SLEEP_M1005_g N_VGND_c_310_n 0.00585385f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_78 N_SLEEP_M1005_g N_VGND_c_312_n 0.0130277f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_79 SLEEP N_VGND_c_312_n 0.00193939f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_80 N_A_27_413#_c_95_n N_A_c_159_n 0.0106594f $X=0.965 $Y=1.99 $X2=-0.19
+ $Y2=-0.24
cc_81 N_A_27_413#_c_87_n N_A_M1000_g 0.00436452f $X=0.965 $Y=1.89 $X2=0 $Y2=0
cc_82 N_A_27_413#_M1007_g N_A_M1000_g 0.0516569f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_83 N_A_27_413#_c_92_n N_A_M1000_g 3.6021e-19 $X=1 $Y=0.97 $X2=0 $Y2=0
cc_84 N_A_27_413#_c_93_n N_A_M1000_g 0.00237117f $X=1 $Y=0.88 $X2=0 $Y2=0
cc_85 N_A_27_413#_c_87_n N_A_c_162_n 0.0155964f $X=0.965 $Y=1.89 $X2=0 $Y2=0
cc_86 N_A_27_413#_c_88_n N_A_c_162_n 0.00236694f $X=1.385 $Y=0.88 $X2=0 $Y2=0
cc_87 N_A_27_413#_c_87_n N_A_211_413#_c_202_n 0.00491629f $X=0.965 $Y=1.89 $X2=0
+ $Y2=0
cc_88 N_A_27_413#_c_95_n N_A_211_413#_c_202_n 0.00160047f $X=0.965 $Y=1.99 $X2=0
+ $Y2=0
cc_89 N_A_27_413#_c_97_n N_A_211_413#_c_202_n 0.0190097f $X=0.645 $Y=1.9 $X2=0
+ $Y2=0
cc_90 N_A_27_413#_c_91_n N_A_211_413#_c_202_n 0.0235825f $X=0.77 $Y=1.785 $X2=0
+ $Y2=0
cc_91 N_A_27_413#_c_88_n N_A_211_413#_c_198_n 0.0054228f $X=1.385 $Y=0.88 $X2=0
+ $Y2=0
cc_92 N_A_27_413#_M1007_g N_A_211_413#_c_198_n 0.00569078f $X=1.46 $Y=0.445
+ $X2=0 $Y2=0
cc_93 N_A_27_413#_c_90_n N_A_211_413#_c_198_n 0.00680547f $X=0.73 $Y=0.445 $X2=0
+ $Y2=0
cc_94 N_A_27_413#_c_92_n N_A_211_413#_c_198_n 0.0106003f $X=1 $Y=0.97 $X2=0
+ $Y2=0
cc_95 N_A_27_413#_c_87_n N_A_211_413#_c_199_n 0.00452546f $X=0.965 $Y=1.89 $X2=0
+ $Y2=0
cc_96 N_A_27_413#_c_88_n N_A_211_413#_c_199_n 0.00976362f $X=1.385 $Y=0.88 $X2=0
+ $Y2=0
cc_97 N_A_27_413#_c_91_n N_A_211_413#_c_199_n 0.0200374f $X=0.77 $Y=1.785 $X2=0
+ $Y2=0
cc_98 N_A_27_413#_c_92_n N_A_211_413#_c_199_n 0.0271875f $X=1 $Y=0.97 $X2=0
+ $Y2=0
cc_99 N_A_27_413#_c_93_n N_A_211_413#_c_199_n 0.00240816f $X=1 $Y=0.88 $X2=0
+ $Y2=0
cc_100 N_A_27_413#_c_88_n N_A_211_413#_c_218_n 0.00602472f $X=1.385 $Y=0.88
+ $X2=0 $Y2=0
cc_101 N_A_27_413#_M1007_g N_A_211_413#_c_218_n 0.00560284f $X=1.46 $Y=0.445
+ $X2=0 $Y2=0
cc_102 N_A_27_413#_c_90_n N_A_211_413#_c_218_n 0.0183359f $X=0.73 $Y=0.445 $X2=0
+ $Y2=0
cc_103 N_A_27_413#_c_92_n N_A_211_413#_c_218_n 0.00101452f $X=1 $Y=0.97 $X2=0
+ $Y2=0
cc_104 N_A_27_413#_c_95_n N_VPWR_c_253_n 0.00817078f $X=0.965 $Y=1.99 $X2=0
+ $Y2=0
cc_105 N_A_27_413#_c_96_n N_VPWR_c_253_n 0.0194103f $X=0.26 $Y=2.225 $X2=0 $Y2=0
cc_106 N_A_27_413#_c_97_n N_VPWR_c_253_n 0.0264502f $X=0.645 $Y=1.9 $X2=0 $Y2=0
cc_107 N_A_27_413#_c_96_n N_VPWR_c_254_n 0.010445f $X=0.26 $Y=2.225 $X2=0 $Y2=0
cc_108 N_A_27_413#_c_97_n N_VPWR_c_254_n 0.00252438f $X=0.645 $Y=1.9 $X2=0 $Y2=0
cc_109 N_A_27_413#_M1001_s N_VPWR_c_252_n 0.00388418f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_110 N_A_27_413#_c_95_n N_VPWR_c_252_n 0.0108251f $X=0.965 $Y=1.99 $X2=0 $Y2=0
cc_111 N_A_27_413#_c_96_n N_VPWR_c_252_n 0.00640243f $X=0.26 $Y=2.225 $X2=0
+ $Y2=0
cc_112 N_A_27_413#_c_97_n N_VPWR_c_252_n 0.00568986f $X=0.645 $Y=1.9 $X2=0 $Y2=0
cc_113 N_A_27_413#_c_95_n N_VPWR_c_258_n 0.00643335f $X=0.965 $Y=1.99 $X2=0
+ $Y2=0
cc_114 N_A_27_413#_M1007_g N_VGND_c_310_n 0.00388886f $X=1.46 $Y=0.445 $X2=0
+ $Y2=0
cc_115 N_A_27_413#_c_90_n N_VGND_c_310_n 0.0140172f $X=0.73 $Y=0.445 $X2=0 $Y2=0
cc_116 N_A_27_413#_M1005_d N_VGND_c_312_n 0.0038379f $X=0.595 $Y=0.235 $X2=0
+ $Y2=0
cc_117 N_A_27_413#_M1007_g N_VGND_c_312_n 0.00665486f $X=1.46 $Y=0.445 $X2=0
+ $Y2=0
cc_118 N_A_27_413#_c_90_n N_VGND_c_312_n 0.00898926f $X=0.73 $Y=0.445 $X2=0
+ $Y2=0
cc_119 N_A_27_413#_c_92_n N_VGND_c_312_n 0.00958879f $X=1 $Y=0.97 $X2=0 $Y2=0
cc_120 N_A_27_413#_c_93_n N_VGND_c_312_n 0.00692832f $X=1 $Y=0.88 $X2=0 $Y2=0
cc_121 N_A_M1000_g N_A_211_413#_c_196_n 0.0258936f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_122 A N_A_211_413#_c_196_n 0.00185434f $X=1.605 $Y=1.785 $X2=0 $Y2=0
cc_123 N_A_M1000_g N_A_211_413#_c_197_n 0.0156991f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_124 N_A_c_159_n N_A_211_413#_c_202_n 0.00203711f $X=1.455 $Y=1.99 $X2=0 $Y2=0
cc_125 N_A_M1000_g N_A_211_413#_c_202_n 0.00174203f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_126 A N_A_211_413#_c_202_n 0.0241053f $X=1.605 $Y=1.785 $X2=0 $Y2=0
cc_127 N_A_c_162_n N_A_211_413#_c_202_n 0.00621711f $X=1.67 $Y=1.73 $X2=0 $Y2=0
cc_128 N_A_M1000_g N_A_211_413#_c_198_n 0.00638307f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_129 N_A_M1000_g N_A_211_413#_c_199_n 0.0301133f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_130 A N_A_211_413#_c_199_n 0.0268966f $X=1.605 $Y=1.785 $X2=0 $Y2=0
cc_131 N_A_c_162_n N_A_211_413#_c_199_n 0.011394f $X=1.67 $Y=1.73 $X2=0 $Y2=0
cc_132 N_A_M1000_g N_A_211_413#_c_200_n 0.00669547f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_133 N_A_c_159_n N_VPWR_c_253_n 6.79847e-19 $X=1.455 $Y=1.99 $X2=0 $Y2=0
cc_134 N_A_c_159_n N_VPWR_c_252_n 0.0126424f $X=1.455 $Y=1.99 $X2=0 $Y2=0
cc_135 A N_VPWR_c_252_n 0.0030545f $X=1.605 $Y=1.785 $X2=0 $Y2=0
cc_136 N_A_c_162_n N_VPWR_c_252_n 4.86259e-19 $X=1.67 $Y=1.73 $X2=0 $Y2=0
cc_137 N_A_c_159_n N_VPWR_c_258_n 0.00702461f $X=1.455 $Y=1.99 $X2=0 $Y2=0
cc_138 N_A_c_162_n N_VPWR_c_258_n 3.80525e-19 $X=1.67 $Y=1.73 $X2=0 $Y2=0
cc_139 N_A_c_159_n N_VPWR_c_259_n 0.00363135f $X=1.455 $Y=1.99 $X2=0 $Y2=0
cc_140 A N_VPWR_c_259_n 0.017383f $X=1.605 $Y=1.785 $X2=0 $Y2=0
cc_141 N_A_c_162_n N_VPWR_c_259_n 0.00424172f $X=1.67 $Y=1.73 $X2=0 $Y2=0
cc_142 A X 0.00791941f $X=1.605 $Y=1.785 $X2=0 $Y2=0
cc_143 N_A_c_162_n X 0.00132493f $X=1.67 $Y=1.73 $X2=0 $Y2=0
cc_144 N_A_M1000_g N_VGND_c_309_n 0.00907f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_145 N_A_M1000_g N_VGND_c_310_n 0.00585385f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_146 N_A_M1000_g N_VGND_c_312_n 0.0112294f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_147 N_A_211_413#_c_196_n N_VPWR_c_255_n 0.00627701f $X=2.47 $Y=1.41 $X2=0
+ $Y2=0
cc_148 N_A_211_413#_M1006_d N_VPWR_c_252_n 0.00346822f $X=1.055 $Y=2.065 $X2=0
+ $Y2=0
cc_149 N_A_211_413#_c_196_n N_VPWR_c_252_n 0.0131269f $X=2.47 $Y=1.41 $X2=0
+ $Y2=0
cc_150 N_A_211_413#_c_202_n N_VPWR_c_252_n 0.0100902f $X=1.21 $Y=2.225 $X2=0
+ $Y2=0
cc_151 N_A_211_413#_c_202_n N_VPWR_c_258_n 0.0127054f $X=1.21 $Y=2.225 $X2=0
+ $Y2=0
cc_152 N_A_211_413#_c_196_n N_VPWR_c_259_n 0.0111983f $X=2.47 $Y=1.41 $X2=0
+ $Y2=0
cc_153 N_A_211_413#_c_196_n X 0.0269696f $X=2.47 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_211_413#_c_196_n N_X_c_292_n 0.00347882f $X=2.47 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_211_413#_c_197_n N_X_c_292_n 0.0136803f $X=2.495 $Y=0.985 $X2=0 $Y2=0
cc_156 N_A_211_413#_c_200_n N_X_c_292_n 0.0150073f $X=2.39 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A_211_413#_c_196_n N_VGND_c_309_n 8.08257e-19 $X=2.47 $Y=1.41 $X2=0
+ $Y2=0
cc_158 N_A_211_413#_c_197_n N_VGND_c_309_n 0.00372187f $X=2.495 $Y=0.985 $X2=0
+ $Y2=0
cc_159 N_A_211_413#_c_200_n N_VGND_c_309_n 0.0156725f $X=2.39 $Y=1.16 $X2=0
+ $Y2=0
cc_160 N_A_211_413#_c_218_n N_VGND_c_310_n 0.0169914f $X=1.25 $Y=0.445 $X2=0
+ $Y2=0
cc_161 N_A_211_413#_c_197_n N_VGND_c_311_n 0.00585385f $X=2.495 $Y=0.985 $X2=0
+ $Y2=0
cc_162 N_A_211_413#_M1007_s N_VGND_c_312_n 0.00239557f $X=1.125 $Y=0.235 $X2=0
+ $Y2=0
cc_163 N_A_211_413#_c_197_n N_VGND_c_312_n 0.012334f $X=2.495 $Y=0.985 $X2=0
+ $Y2=0
cc_164 N_A_211_413#_c_218_n N_VGND_c_312_n 0.01456f $X=1.25 $Y=0.445 $X2=0 $Y2=0
cc_165 N_VPWR_c_252_n N_X_M1004_d 0.00228914f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_166 N_VPWR_c_255_n X 0.0234486f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_167 N_VPWR_c_252_n X 0.0206322f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_168 X N_VGND_c_311_n 0.0319568f $X=2.65 $Y=0.425 $X2=0 $Y2=0
cc_169 N_X_M1003_d N_VGND_c_312_n 0.00387172f $X=2.57 $Y=0.235 $X2=0 $Y2=0
cc_170 X N_VGND_c_312_n 0.0175629f $X=2.65 $Y=0.425 $X2=0 $Y2=0
cc_171 N_VGND_c_312_n A_307_47# 0.00711569f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
