# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__clkbuf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkbuf_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.972000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.400000 1.325000 ;
    END
  END A
  PIN VGND
    ANTENNADIFFAREA  1.467900 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  3.245000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  3.529800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.530000 0.280000  2.790000 0.735000 ;
        RECT 2.530000 0.735000 10.025000 0.905000 ;
        RECT 2.530000 1.495000 10.025000 1.720000 ;
        RECT 2.530000 1.720000  8.535000 1.735000 ;
        RECT 2.530000 1.735000  2.790000 2.460000 ;
        RECT 3.490000 0.280000  3.750000 0.735000 ;
        RECT 3.490000 1.735000  3.750000 2.460000 ;
        RECT 4.450000 0.280000  4.710000 0.735000 ;
        RECT 4.450000 1.735000  4.710000 2.460000 ;
        RECT 5.345000 0.280000  5.670000 0.735000 ;
        RECT 5.410000 1.735000  5.670000 2.460000 ;
        RECT 6.355000 0.280000  6.615000 0.735000 ;
        RECT 6.355000 1.735000  6.615000 2.460000 ;
        RECT 7.315000 0.280000  7.575000 0.735000 ;
        RECT 7.315000 1.735000  7.575000 2.460000 ;
        RECT 8.275000 0.280000  8.535000 0.735000 ;
        RECT 8.275000 1.735000  8.535000 2.460000 ;
        RECT 8.760000 0.905000 10.025000 1.495000 ;
        RECT 9.245000 0.280000  9.505000 0.735000 ;
        RECT 9.245000 1.720000  9.535000 2.460000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.085000  0.085000  0.390000 0.595000 ;
      RECT 0.095000  1.825000  0.390000 2.635000 ;
      RECT 0.620000  0.265000  0.870000 1.075000 ;
      RECT 0.620000  1.075000  8.540000 1.325000 ;
      RECT 0.620000  1.325000  0.865000 2.465000 ;
      RECT 1.090000  0.085000  1.350000 0.610000 ;
      RECT 1.090000  1.825000  1.350000 2.635000 ;
      RECT 1.580000  0.265000  1.830000 1.075000 ;
      RECT 1.580000  1.325000  1.830000 2.460000 ;
      RECT 2.050000  0.085000  2.310000 0.645000 ;
      RECT 2.050000  1.835000  2.310000 2.630000 ;
      RECT 2.050000  2.630000  9.025000 2.635000 ;
      RECT 3.010000  0.085000  3.270000 0.565000 ;
      RECT 3.010000  1.905000  3.270000 2.630000 ;
      RECT 3.970000  0.085000  4.230000 0.565000 ;
      RECT 3.970000  1.905000  4.230000 2.630000 ;
      RECT 4.930000  0.085000  5.175000 0.565000 ;
      RECT 4.930000  1.905000  5.190000 2.630000 ;
      RECT 5.890000  0.085000  6.135000 0.565000 ;
      RECT 5.890000  1.905000  6.135000 2.630000 ;
      RECT 6.845000  0.085000  7.095000 0.565000 ;
      RECT 6.850000  1.905000  7.095000 2.630000 ;
      RECT 7.805000  0.085000  8.055000 0.565000 ;
      RECT 7.810000  1.905000  8.055000 2.630000 ;
      RECT 8.765000  0.085000  9.025000 0.565000 ;
      RECT 8.770000  1.905000  9.025000 2.630000 ;
      RECT 9.725000  0.085000 10.025000 0.565000 ;
      RECT 9.755000  1.890000 10.025000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkbuf_16
END LIBRARY
