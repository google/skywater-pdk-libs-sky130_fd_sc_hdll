* File: sky130_fd_sc_hdll__isobufsrc_16.pex.spice
* Created: Wed Sep  2 08:33:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_16%A 3 5 6 8 9 11 12 14 15 17 18 20 21
+ 23 24 26 29 32 33 40
r78 40 41 39.1708 $w=3.63e-07 $l=2.95e-07 $layer=POLY_cond $X=2.225 $Y=1.202
+ $X2=2.52 $Y2=1.202
r79 39 40 36.5152 $w=3.63e-07 $l=2.75e-07 $layer=POLY_cond $X=1.95 $Y=1.202
+ $X2=2.225 $Y2=1.202
r80 38 39 32.5317 $w=3.63e-07 $l=2.45e-07 $layer=POLY_cond $X=1.705 $Y=1.202
+ $X2=1.95 $Y2=1.202
r81 37 38 36.5152 $w=3.63e-07 $l=2.75e-07 $layer=POLY_cond $X=1.43 $Y=1.202
+ $X2=1.705 $Y2=1.202
r82 36 37 32.5317 $w=3.63e-07 $l=2.45e-07 $layer=POLY_cond $X=1.185 $Y=1.202
+ $X2=1.43 $Y2=1.202
r83 35 36 36.5152 $w=3.63e-07 $l=2.75e-07 $layer=POLY_cond $X=0.91 $Y=1.202
+ $X2=1.185 $Y2=1.202
r84 34 35 32.5317 $w=3.63e-07 $l=2.45e-07 $layer=POLY_cond $X=0.665 $Y=1.202
+ $X2=0.91 $Y2=1.202
r85 32 34 11.2865 $w=3.63e-07 $l=8.5e-08 $layer=POLY_cond $X=0.58 $Y=1.202
+ $X2=0.665 $Y2=1.202
r86 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.58
+ $Y=1.16 $X2=0.58 $Y2=1.16
r87 29 33 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.38 $Y=1.16 $X2=0.58
+ $Y2=1.16
r88 24 41 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.52 $Y=0.995
+ $X2=2.52 $Y2=1.202
r89 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.52 $Y=0.995
+ $X2=2.52 $Y2=0.56
r90 21 40 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.225 $Y=1.41
+ $X2=2.225 $Y2=1.202
r91 21 23 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.225 $Y=1.41
+ $X2=2.225 $Y2=1.985
r92 18 39 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=1.202
r93 18 20 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=0.56
r94 15 38 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.705 $Y=1.41
+ $X2=1.705 $Y2=1.202
r95 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.705 $Y=1.41
+ $X2=1.705 $Y2=1.985
r96 12 37 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=1.202
r97 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=0.56
r98 9 36 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.185 $Y=1.41
+ $X2=1.185 $Y2=1.202
r99 9 11 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.185 $Y=1.41
+ $X2=1.185 $Y2=1.985
r100 6 35 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.202
r101 6 8 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=0.56
r102 3 34 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.665 $Y=1.41
+ $X2=0.665 $Y2=1.202
r103 3 5 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.665 $Y=1.41
+ $X2=0.665 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_16%A_151_297# 1 2 3 4 13 15 16 18 19 21
+ 22 24 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 51 52 54 55 57 58 60
+ 61 63 64 66 67 69 70 72 73 75 76 78 79 81 82 84 85 87 88 90 91 93 94 96 97 99
+ 100 102 103 105 106 108 111 117 119 120 123 129 136 140 141 145 178
r335 178 179 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=10.355 $Y=1.202
+ $X2=10.38 $Y2=1.202
r336 175 176 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=9.86 $Y=1.202
+ $X2=9.885 $Y2=1.202
r337 174 175 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=9.415 $Y=1.202
+ $X2=9.86 $Y2=1.202
r338 173 174 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=9.39 $Y=1.202
+ $X2=9.415 $Y2=1.202
r339 172 173 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=8.945 $Y=1.202
+ $X2=9.39 $Y2=1.202
r340 171 172 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=8.92 $Y=1.202
+ $X2=8.945 $Y2=1.202
r341 170 171 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=8.475 $Y=1.202
+ $X2=8.92 $Y2=1.202
r342 169 170 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=8.45 $Y=1.202
+ $X2=8.475 $Y2=1.202
r343 168 169 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=8.005 $Y=1.202
+ $X2=8.45 $Y2=1.202
r344 167 168 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=7.98 $Y=1.202
+ $X2=8.005 $Y2=1.202
r345 166 167 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=7.535 $Y=1.202
+ $X2=7.98 $Y2=1.202
r346 165 166 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=7.51 $Y=1.202
+ $X2=7.535 $Y2=1.202
r347 164 165 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=7.065 $Y=1.202
+ $X2=7.51 $Y2=1.202
r348 163 164 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=7.04 $Y=1.202
+ $X2=7.065 $Y2=1.202
r349 162 163 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=6.595 $Y=1.202
+ $X2=7.04 $Y2=1.202
r350 161 162 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=6.57 $Y=1.202
+ $X2=6.595 $Y2=1.202
r351 160 161 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=6.125 $Y=1.202
+ $X2=6.57 $Y2=1.202
r352 159 160 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=6.1 $Y=1.202
+ $X2=6.125 $Y2=1.202
r353 158 159 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=5.655 $Y=1.202
+ $X2=6.1 $Y2=1.202
r354 157 158 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=5.63 $Y=1.202
+ $X2=5.655 $Y2=1.202
r355 156 157 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=5.185 $Y=1.202
+ $X2=5.63 $Y2=1.202
r356 155 156 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=5.16 $Y=1.202
+ $X2=5.185 $Y2=1.202
r357 154 155 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=4.715 $Y=1.202
+ $X2=5.16 $Y2=1.202
r358 153 154 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=4.69 $Y=1.202
+ $X2=4.715 $Y2=1.202
r359 152 153 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=4.245 $Y=1.202
+ $X2=4.69 $Y2=1.202
r360 151 152 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=4.22 $Y=1.202
+ $X2=4.245 $Y2=1.202
r361 150 151 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=3.775 $Y=1.202
+ $X2=4.22 $Y2=1.202
r362 149 150 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=3.75 $Y=1.202
+ $X2=3.775 $Y2=1.202
r363 146 147 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=3.28 $Y=1.202
+ $X2=3.305 $Y2=1.202
r364 140 141 5.82817 $w=4.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.9 $Y=1.62
+ $X2=0.9 $Y2=1.495
r365 137 178 15.1035 $w=3.67e-07 $l=1.15e-07 $layer=POLY_cond $X=10.24 $Y=1.202
+ $X2=10.355 $Y2=1.202
r366 137 176 46.624 $w=3.67e-07 $l=3.55e-07 $layer=POLY_cond $X=10.24 $Y=1.202
+ $X2=9.885 $Y2=1.202
r367 136 137 15.2926 $w=1.7e-07 $l=1.615e-06 $layer=licon1_POLY $count=9
+ $X=10.24 $Y=1.16 $X2=10.24 $Y2=1.16
r368 134 149 49.9074 $w=3.67e-07 $l=3.8e-07 $layer=POLY_cond $X=3.37 $Y=1.202
+ $X2=3.75 $Y2=1.202
r369 134 147 8.53679 $w=3.67e-07 $l=6.5e-08 $layer=POLY_cond $X=3.37 $Y=1.202
+ $X2=3.305 $Y2=1.202
r370 133 136 362.831 $w=2.08e-07 $l=6.87e-06 $layer=LI1_cond $X=3.37 $Y=1.18
+ $X2=10.24 $Y2=1.18
r371 133 134 15.2926 $w=1.7e-07 $l=1.615e-06 $layer=licon1_POLY $count=9 $X=3.37
+ $Y=1.16 $X2=3.37 $Y2=1.16
r372 131 145 4.79724 $w=2.1e-07 $l=3.32491e-07 $layer=LI1_cond $X=2.385 $Y=1.18
+ $X2=2.055 $Y2=1.175
r373 131 133 52.0216 $w=2.08e-07 $l=9.85e-07 $layer=LI1_cond $X=2.385 $Y=1.18
+ $X2=3.37 $Y2=1.18
r374 127 145 1.60795 $w=3e-07 $l=2.28473e-07 $layer=LI1_cond $X=2.235 $Y=1.065
+ $X2=2.055 $Y2=1.175
r375 127 129 24.7775 $w=2.98e-07 $l=6.45e-07 $layer=LI1_cond $X=2.235 $Y=1.065
+ $X2=2.235 $Y2=0.42
r376 123 125 18.2247 $w=4.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.94 $Y=1.62
+ $X2=1.94 $Y2=2.3
r377 121 145 1.60795 $w=4.3e-07 $l=1.60857e-07 $layer=LI1_cond $X=1.94 $Y=1.285
+ $X2=2.055 $Y2=1.175
r378 121 123 8.97834 $w=4.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.94 $Y=1.285
+ $X2=1.94 $Y2=1.62
r379 119 145 4.79724 $w=2.2e-07 $l=3.3e-07 $layer=LI1_cond $X=1.725 $Y=1.175
+ $X2=2.055 $Y2=1.175
r380 119 120 19.9058 $w=2.18e-07 $l=3.8e-07 $layer=LI1_cond $X=1.725 $Y=1.175
+ $X2=1.345 $Y2=1.175
r381 115 120 6.80989 $w=2.18e-07 $l=1.3e-07 $layer=LI1_cond $X=1.215 $Y=1.175
+ $X2=1.345 $Y2=1.175
r382 115 142 11.2625 $w=2.18e-07 $l=2.15e-07 $layer=LI1_cond $X=1.215 $Y=1.175
+ $X2=1 $Y2=1.175
r383 115 117 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=1.215 $Y=1.065
+ $X2=1.215 $Y2=0.42
r384 113 142 0.443598 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=1 $Y=1.285 $X2=1
+ $Y2=1.175
r385 113 141 10.5223 $w=2.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1 $Y=1.285 $X2=1
+ $Y2=1.495
r386 109 140 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=0.9 $Y=1.71 $X2=0.9
+ $Y2=1.62
r387 109 111 15.8126 $w=4.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.9 $Y=1.71
+ $X2=0.9 $Y2=2.3
r388 106 179 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.38 $Y=0.995
+ $X2=10.38 $Y2=1.202
r389 106 108 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.38 $Y=0.995
+ $X2=10.38 $Y2=0.56
r390 103 178 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.355 $Y=1.41
+ $X2=10.355 $Y2=1.202
r391 103 105 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.355 $Y=1.41
+ $X2=10.355 $Y2=1.985
r392 100 176 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.885 $Y=1.41
+ $X2=9.885 $Y2=1.202
r393 100 102 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.885 $Y=1.41
+ $X2=9.885 $Y2=1.985
r394 97 175 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.86 $Y=0.995
+ $X2=9.86 $Y2=1.202
r395 97 99 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.86 $Y=0.995
+ $X2=9.86 $Y2=0.56
r396 94 174 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.415 $Y=1.41
+ $X2=9.415 $Y2=1.202
r397 94 96 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.415 $Y=1.41
+ $X2=9.415 $Y2=1.985
r398 91 173 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.39 $Y=0.995
+ $X2=9.39 $Y2=1.202
r399 91 93 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.39 $Y=0.995
+ $X2=9.39 $Y2=0.56
r400 88 172 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.945 $Y=1.41
+ $X2=8.945 $Y2=1.202
r401 88 90 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.945 $Y=1.41
+ $X2=8.945 $Y2=1.985
r402 85 171 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.92 $Y=0.995
+ $X2=8.92 $Y2=1.202
r403 85 87 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.92 $Y=0.995
+ $X2=8.92 $Y2=0.56
r404 82 170 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.475 $Y=1.41
+ $X2=8.475 $Y2=1.202
r405 82 84 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.475 $Y=1.41
+ $X2=8.475 $Y2=1.985
r406 79 169 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.45 $Y=0.995
+ $X2=8.45 $Y2=1.202
r407 79 81 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.45 $Y=0.995
+ $X2=8.45 $Y2=0.56
r408 76 168 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.005 $Y=1.41
+ $X2=8.005 $Y2=1.202
r409 76 78 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.005 $Y=1.41
+ $X2=8.005 $Y2=1.985
r410 73 167 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.98 $Y=0.995
+ $X2=7.98 $Y2=1.202
r411 73 75 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.98 $Y=0.995
+ $X2=7.98 $Y2=0.56
r412 70 166 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.535 $Y=1.41
+ $X2=7.535 $Y2=1.202
r413 70 72 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.535 $Y=1.41
+ $X2=7.535 $Y2=1.985
r414 67 165 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.51 $Y=0.995
+ $X2=7.51 $Y2=1.202
r415 67 69 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.51 $Y=0.995
+ $X2=7.51 $Y2=0.56
r416 64 164 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.065 $Y=1.41
+ $X2=7.065 $Y2=1.202
r417 64 66 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.065 $Y=1.41
+ $X2=7.065 $Y2=1.985
r418 61 163 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.04 $Y=0.995
+ $X2=7.04 $Y2=1.202
r419 61 63 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.04 $Y=0.995
+ $X2=7.04 $Y2=0.56
r420 58 162 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.595 $Y=1.41
+ $X2=6.595 $Y2=1.202
r421 58 60 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.595 $Y=1.41
+ $X2=6.595 $Y2=1.985
r422 55 161 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.57 $Y=0.995
+ $X2=6.57 $Y2=1.202
r423 55 57 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.57 $Y=0.995
+ $X2=6.57 $Y2=0.56
r424 52 160 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.125 $Y=1.41
+ $X2=6.125 $Y2=1.202
r425 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.125 $Y=1.41
+ $X2=6.125 $Y2=1.985
r426 49 159 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.1 $Y=0.995
+ $X2=6.1 $Y2=1.202
r427 49 51 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.1 $Y=0.995
+ $X2=6.1 $Y2=0.56
r428 46 158 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.655 $Y=1.41
+ $X2=5.655 $Y2=1.202
r429 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.655 $Y=1.41
+ $X2=5.655 $Y2=1.985
r430 43 157 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.63 $Y=0.995
+ $X2=5.63 $Y2=1.202
r431 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.63 $Y=0.995
+ $X2=5.63 $Y2=0.56
r432 40 156 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.185 $Y=1.41
+ $X2=5.185 $Y2=1.202
r433 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.185 $Y=1.41
+ $X2=5.185 $Y2=1.985
r434 37 155 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.16 $Y=0.995
+ $X2=5.16 $Y2=1.202
r435 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.16 $Y=0.995
+ $X2=5.16 $Y2=0.56
r436 34 154 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.715 $Y=1.41
+ $X2=4.715 $Y2=1.202
r437 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.715 $Y=1.41
+ $X2=4.715 $Y2=1.985
r438 31 153 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.69 $Y=0.995
+ $X2=4.69 $Y2=1.202
r439 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.69 $Y=0.995
+ $X2=4.69 $Y2=0.56
r440 28 152 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.245 $Y=1.41
+ $X2=4.245 $Y2=1.202
r441 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.245 $Y=1.41
+ $X2=4.245 $Y2=1.985
r442 25 151 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.22 $Y=0.995
+ $X2=4.22 $Y2=1.202
r443 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.22 $Y=0.995
+ $X2=4.22 $Y2=0.56
r444 22 150 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.775 $Y=1.41
+ $X2=3.775 $Y2=1.202
r445 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.775 $Y=1.41
+ $X2=3.775 $Y2=1.985
r446 19 149 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.75 $Y=0.995
+ $X2=3.75 $Y2=1.202
r447 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.75 $Y=0.995
+ $X2=3.75 $Y2=0.56
r448 16 147 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.305 $Y=1.41
+ $X2=3.305 $Y2=1.202
r449 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.305 $Y=1.41
+ $X2=3.305 $Y2=1.985
r450 13 146 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.28 $Y=0.995
+ $X2=3.28 $Y2=1.202
r451 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.28 $Y=0.995
+ $X2=3.28 $Y2=0.56
r452 4 125 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.795
+ $Y=1.485 $X2=1.94 $Y2=2.3
r453 4 123 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.795
+ $Y=1.485 $X2=1.94 $Y2=1.62
r454 3 140 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.755
+ $Y=1.485 $X2=0.9 $Y2=1.62
r455 3 111 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.755
+ $Y=1.485 $X2=0.9 $Y2=2.3
r456 2 129 91 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=2 $X=2.025
+ $Y=0.235 $X2=2.21 $Y2=0.42
r457 1 117 91 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=2 $X=0.985
+ $Y=0.235 $X2=1.17 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_16%SLEEP 1 3 4 6 7 9 10 12 13 15 16 18
+ 19 21 22 24 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 51 52 54 55 57
+ 58 60 61 63 64 66 67 69 70 72 73 75 76 78 79 81 82 84 85 87 88 90 91 93 94 96
+ 97 132 135 140
r277 135 136 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=17.875 $Y=1.202
+ $X2=17.9 $Y2=1.202
r278 134 135 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=17.405 $Y=1.202
+ $X2=17.875 $Y2=1.202
r279 133 134 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=17.38 $Y=1.202
+ $X2=17.405 $Y2=1.202
r280 131 133 1.31335 $w=3.67e-07 $l=1e-08 $layer=POLY_cond $X=17.37 $Y=1.202
+ $X2=17.38 $Y2=1.202
r281 131 132 16.1422 $w=1.7e-07 $l=1.53e-06 $layer=licon1_POLY $count=9 $X=17.37
+ $Y=1.16 $X2=17.37 $Y2=1.16
r282 129 131 57.1308 $w=3.67e-07 $l=4.35e-07 $layer=POLY_cond $X=16.935 $Y=1.202
+ $X2=17.37 $Y2=1.202
r283 128 129 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=16.91 $Y=1.202
+ $X2=16.935 $Y2=1.202
r284 127 128 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=16.465 $Y=1.202
+ $X2=16.91 $Y2=1.202
r285 126 127 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=16.44 $Y=1.202
+ $X2=16.465 $Y2=1.202
r286 125 126 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=15.995 $Y=1.202
+ $X2=16.44 $Y2=1.202
r287 124 125 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=15.97 $Y=1.202
+ $X2=15.995 $Y2=1.202
r288 123 124 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=15.525 $Y=1.202
+ $X2=15.97 $Y2=1.202
r289 122 123 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=15.5 $Y=1.202
+ $X2=15.525 $Y2=1.202
r290 121 122 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=15.055 $Y=1.202
+ $X2=15.5 $Y2=1.202
r291 120 121 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=15.03 $Y=1.202
+ $X2=15.055 $Y2=1.202
r292 119 120 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=14.585 $Y=1.202
+ $X2=15.03 $Y2=1.202
r293 118 119 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=14.56 $Y=1.202
+ $X2=14.585 $Y2=1.202
r294 117 118 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=14.115 $Y=1.202
+ $X2=14.56 $Y2=1.202
r295 116 117 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=14.09 $Y=1.202
+ $X2=14.115 $Y2=1.202
r296 115 116 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=13.645 $Y=1.202
+ $X2=14.09 $Y2=1.202
r297 114 115 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=13.62 $Y=1.202
+ $X2=13.645 $Y2=1.202
r298 113 114 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=13.175 $Y=1.202
+ $X2=13.62 $Y2=1.202
r299 112 113 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=13.15 $Y=1.202
+ $X2=13.175 $Y2=1.202
r300 111 112 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=12.705 $Y=1.202
+ $X2=13.15 $Y2=1.202
r301 110 111 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=12.68 $Y=1.202
+ $X2=12.705 $Y2=1.202
r302 109 110 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=12.235 $Y=1.202
+ $X2=12.68 $Y2=1.202
r303 108 109 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=12.21 $Y=1.202
+ $X2=12.235 $Y2=1.202
r304 107 108 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=11.765 $Y=1.202
+ $X2=12.21 $Y2=1.202
r305 106 107 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=11.74 $Y=1.202
+ $X2=11.765 $Y2=1.202
r306 105 106 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=11.295 $Y=1.202
+ $X2=11.74 $Y2=1.202
r307 104 105 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=11.27 $Y=1.202
+ $X2=11.295 $Y2=1.202
r308 103 140 89.2554 $w=2.08e-07 $l=1.69e-06 $layer=LI1_cond $X=10.89 $Y=1.18
+ $X2=12.58 $Y2=1.18
r309 102 104 49.9074 $w=3.67e-07 $l=3.8e-07 $layer=POLY_cond $X=10.89 $Y=1.202
+ $X2=11.27 $Y2=1.202
r310 102 103 16.1422 $w=1.7e-07 $l=1.53e-06 $layer=licon1_POLY $count=9 $X=10.89
+ $Y=1.16 $X2=10.89 $Y2=1.16
r311 100 102 8.53679 $w=3.67e-07 $l=6.5e-08 $layer=POLY_cond $X=10.825 $Y=1.202
+ $X2=10.89 $Y2=1.202
r312 99 100 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=10.8 $Y=1.202
+ $X2=10.825 $Y2=1.202
r313 97 132 171.117 $w=2.08e-07 $l=3.24e-06 $layer=LI1_cond $X=14.13 $Y=1.18
+ $X2=17.37 $Y2=1.18
r314 97 140 81.8615 $w=2.08e-07 $l=1.55e-06 $layer=LI1_cond $X=14.13 $Y=1.18
+ $X2=12.58 $Y2=1.18
r315 94 136 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=17.9 $Y=0.995
+ $X2=17.9 $Y2=1.202
r316 94 96 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=17.9 $Y=0.995
+ $X2=17.9 $Y2=0.56
r317 91 135 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=17.875 $Y=1.41
+ $X2=17.875 $Y2=1.202
r318 91 93 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=17.875 $Y=1.41
+ $X2=17.875 $Y2=1.985
r319 88 134 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=17.405 $Y=1.41
+ $X2=17.405 $Y2=1.202
r320 88 90 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=17.405 $Y=1.41
+ $X2=17.405 $Y2=1.985
r321 85 133 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=17.38 $Y=0.995
+ $X2=17.38 $Y2=1.202
r322 85 87 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=17.38 $Y=0.995
+ $X2=17.38 $Y2=0.56
r323 82 129 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=16.935 $Y=1.41
+ $X2=16.935 $Y2=1.202
r324 82 84 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=16.935 $Y=1.41
+ $X2=16.935 $Y2=1.985
r325 79 128 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=16.91 $Y=0.995
+ $X2=16.91 $Y2=1.202
r326 79 81 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=16.91 $Y=0.995
+ $X2=16.91 $Y2=0.56
r327 76 127 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=16.465 $Y=1.41
+ $X2=16.465 $Y2=1.202
r328 76 78 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=16.465 $Y=1.41
+ $X2=16.465 $Y2=1.985
r329 73 126 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=16.44 $Y=0.995
+ $X2=16.44 $Y2=1.202
r330 73 75 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=16.44 $Y=0.995
+ $X2=16.44 $Y2=0.56
r331 70 125 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=15.995 $Y=1.41
+ $X2=15.995 $Y2=1.202
r332 70 72 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.995 $Y=1.41
+ $X2=15.995 $Y2=1.985
r333 67 124 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=15.97 $Y=0.995
+ $X2=15.97 $Y2=1.202
r334 67 69 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=15.97 $Y=0.995
+ $X2=15.97 $Y2=0.56
r335 64 123 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=15.525 $Y=1.41
+ $X2=15.525 $Y2=1.202
r336 64 66 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.525 $Y=1.41
+ $X2=15.525 $Y2=1.985
r337 61 122 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=15.5 $Y=0.995
+ $X2=15.5 $Y2=1.202
r338 61 63 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=15.5 $Y=0.995
+ $X2=15.5 $Y2=0.56
r339 58 121 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=15.055 $Y=1.41
+ $X2=15.055 $Y2=1.202
r340 58 60 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.055 $Y=1.41
+ $X2=15.055 $Y2=1.985
r341 55 120 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=15.03 $Y=0.995
+ $X2=15.03 $Y2=1.202
r342 55 57 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=15.03 $Y=0.995
+ $X2=15.03 $Y2=0.56
r343 52 119 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=14.585 $Y=1.41
+ $X2=14.585 $Y2=1.202
r344 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=14.585 $Y=1.41
+ $X2=14.585 $Y2=1.985
r345 49 118 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=14.56 $Y=0.995
+ $X2=14.56 $Y2=1.202
r346 49 51 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=14.56 $Y=0.995
+ $X2=14.56 $Y2=0.56
r347 46 117 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=14.115 $Y=1.41
+ $X2=14.115 $Y2=1.202
r348 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=14.115 $Y=1.41
+ $X2=14.115 $Y2=1.985
r349 43 116 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=14.09 $Y=0.995
+ $X2=14.09 $Y2=1.202
r350 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=14.09 $Y=0.995
+ $X2=14.09 $Y2=0.56
r351 40 115 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=13.645 $Y=1.41
+ $X2=13.645 $Y2=1.202
r352 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=13.645 $Y=1.41
+ $X2=13.645 $Y2=1.985
r353 37 114 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=13.62 $Y=0.995
+ $X2=13.62 $Y2=1.202
r354 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.62 $Y=0.995
+ $X2=13.62 $Y2=0.56
r355 34 113 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=13.175 $Y=1.41
+ $X2=13.175 $Y2=1.202
r356 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=13.175 $Y=1.41
+ $X2=13.175 $Y2=1.985
r357 31 112 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=13.15 $Y=0.995
+ $X2=13.15 $Y2=1.202
r358 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.15 $Y=0.995
+ $X2=13.15 $Y2=0.56
r359 28 111 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=12.705 $Y=1.41
+ $X2=12.705 $Y2=1.202
r360 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.705 $Y=1.41
+ $X2=12.705 $Y2=1.985
r361 25 110 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=12.68 $Y=0.995
+ $X2=12.68 $Y2=1.202
r362 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.68 $Y=0.995
+ $X2=12.68 $Y2=0.56
r363 22 109 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=12.235 $Y=1.41
+ $X2=12.235 $Y2=1.202
r364 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.235 $Y=1.41
+ $X2=12.235 $Y2=1.985
r365 19 108 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=12.21 $Y=0.995
+ $X2=12.21 $Y2=1.202
r366 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.21 $Y=0.995
+ $X2=12.21 $Y2=0.56
r367 16 107 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=11.765 $Y=1.41
+ $X2=11.765 $Y2=1.202
r368 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.765 $Y=1.41
+ $X2=11.765 $Y2=1.985
r369 13 106 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.74 $Y=0.995
+ $X2=11.74 $Y2=1.202
r370 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.74 $Y=0.995
+ $X2=11.74 $Y2=0.56
r371 10 105 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=11.295 $Y=1.41
+ $X2=11.295 $Y2=1.202
r372 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.295 $Y=1.41
+ $X2=11.295 $Y2=1.985
r373 7 104 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.27 $Y=0.995
+ $X2=11.27 $Y2=1.202
r374 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.27 $Y=0.995
+ $X2=11.27 $Y2=0.56
r375 4 100 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.825 $Y=1.41
+ $X2=10.825 $Y2=1.202
r376 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.825 $Y=1.41
+ $X2=10.825 $Y2=1.985
r377 1 99 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.8 $Y=0.995
+ $X2=10.8 $Y2=1.202
r378 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.8 $Y=0.995
+ $X2=10.8 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 36 42 48
+ 52 56 58 62 66 70 74 78 82 86 89 90 92 93 95 96 98 99 101 102 104 105 107 108
+ 110 111 112 121 148 149 152 155 158
r237 158 159 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r238 156 159 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r239 155 156 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r240 153 156 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r241 152 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r242 148 149 1.03333 $w=1.7e-07 $l=1.53e-06 $layer=mcon $count=9 $X=18.17
+ $Y=2.72 $X2=18.17 $Y2=2.72
r243 146 149 2.22512 $w=4.8e-07 $l=7.82e-06 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=18.17 $Y2=2.72
r244 145 148 510.182 $w=1.68e-07 $l=7.82e-06 $layer=LI1_cond $X=10.35 $Y=2.72
+ $X2=18.17 $Y2=2.72
r245 145 146 1.03333 $w=1.7e-07 $l=1.53e-06 $layer=mcon $count=9 $X=10.35
+ $Y=2.72 $X2=10.35 $Y2=2.72
r246 143 146 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.35 $Y2=2.72
r247 142 143 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r248 140 143 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r249 139 140 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r250 137 140 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r251 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r252 134 137 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r253 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r254 131 134 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r255 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r256 128 131 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r257 128 159 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.37 $Y2=2.72
r258 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r259 125 158 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.605 $Y=2.72
+ $X2=4.48 $Y2=2.72
r260 125 127 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=4.605 $Y=2.72
+ $X2=5.29 $Y2=2.72
r261 124 153 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r262 123 124 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r263 121 152 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=2.375 $Y=2.72
+ $X2=2.522 $Y2=2.72
r264 121 123 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.375 $Y=2.72
+ $X2=2.07 $Y2=2.72
r265 120 124 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r266 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r267 112 120 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r268 112 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r269 110 142 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=9.995 $Y=2.72
+ $X2=9.89 $Y2=2.72
r270 110 111 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.995 $Y=2.72
+ $X2=10.12 $Y2=2.72
r271 109 145 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=10.245 $Y=2.72
+ $X2=10.35 $Y2=2.72
r272 109 111 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.245 $Y=2.72
+ $X2=10.12 $Y2=2.72
r273 107 139 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=9.055 $Y=2.72
+ $X2=8.97 $Y2=2.72
r274 107 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.055 $Y=2.72
+ $X2=9.18 $Y2=2.72
r275 106 142 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=9.305 $Y=2.72
+ $X2=9.89 $Y2=2.72
r276 106 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.305 $Y=2.72
+ $X2=9.18 $Y2=2.72
r277 104 136 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=8.115 $Y=2.72
+ $X2=8.05 $Y2=2.72
r278 104 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.115 $Y=2.72
+ $X2=8.24 $Y2=2.72
r279 103 139 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=8.365 $Y=2.72
+ $X2=8.97 $Y2=2.72
r280 103 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.365 $Y=2.72
+ $X2=8.24 $Y2=2.72
r281 101 133 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=7.175 $Y=2.72
+ $X2=7.13 $Y2=2.72
r282 101 102 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.175 $Y=2.72
+ $X2=7.3 $Y2=2.72
r283 100 136 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=7.425 $Y=2.72
+ $X2=8.05 $Y2=2.72
r284 100 102 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.425 $Y=2.72
+ $X2=7.3 $Y2=2.72
r285 98 130 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=6.235 $Y=2.72
+ $X2=6.21 $Y2=2.72
r286 98 99 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.235 $Y=2.72
+ $X2=6.36 $Y2=2.72
r287 97 133 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=6.485 $Y=2.72
+ $X2=7.13 $Y2=2.72
r288 97 99 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.485 $Y=2.72
+ $X2=6.36 $Y2=2.72
r289 95 127 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.295 $Y=2.72
+ $X2=5.29 $Y2=2.72
r290 95 96 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.295 $Y=2.72
+ $X2=5.42 $Y2=2.72
r291 94 130 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=5.545 $Y=2.72
+ $X2=6.21 $Y2=2.72
r292 94 96 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.545 $Y=2.72
+ $X2=5.42 $Y2=2.72
r293 92 119 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.15 $Y2=2.72
r294 92 93 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.445 $Y2=2.72
r295 91 123 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=1.555 $Y=2.72
+ $X2=2.07 $Y2=2.72
r296 91 93 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.555 $Y=2.72
+ $X2=1.445 $Y2=2.72
r297 89 115 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=0.3 $Y=2.72 $X2=0.23
+ $Y2=2.72
r298 89 90 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=0.3 $Y=2.72
+ $X2=0.407 $Y2=2.72
r299 88 119 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=1.15 $Y2=2.72
r300 88 90 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.407 $Y2=2.72
r301 84 111 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.12 $Y=2.635
+ $X2=10.12 $Y2=2.72
r302 84 86 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=10.12 $Y=2.635
+ $X2=10.12 $Y2=2
r303 80 108 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.18 $Y=2.635
+ $X2=9.18 $Y2=2.72
r304 80 82 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=9.18 $Y=2.635
+ $X2=9.18 $Y2=2
r305 76 105 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.24 $Y=2.635
+ $X2=8.24 $Y2=2.72
r306 76 78 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=8.24 $Y=2.635
+ $X2=8.24 $Y2=2
r307 72 102 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.3 $Y=2.635
+ $X2=7.3 $Y2=2.72
r308 72 74 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=7.3 $Y=2.635
+ $X2=7.3 $Y2=2
r309 68 99 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.36 $Y=2.635
+ $X2=6.36 $Y2=2.72
r310 68 70 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=6.36 $Y=2.635
+ $X2=6.36 $Y2=2
r311 64 96 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.42 $Y=2.635
+ $X2=5.42 $Y2=2.72
r312 64 66 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=5.42 $Y=2.635
+ $X2=5.42 $Y2=2
r313 60 158 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.48 $Y=2.635
+ $X2=4.48 $Y2=2.72
r314 60 62 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=4.48 $Y=2.635
+ $X2=4.48 $Y2=2
r315 59 155 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.665 $Y=2.72
+ $X2=3.54 $Y2=2.72
r316 58 158 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.355 $Y=2.72
+ $X2=4.48 $Y2=2.72
r317 58 59 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.355 $Y=2.72
+ $X2=3.665 $Y2=2.72
r318 54 155 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=2.635
+ $X2=3.54 $Y2=2.72
r319 54 56 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=3.54 $Y=2.635
+ $X2=3.54 $Y2=2
r320 53 152 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=2.67 $Y=2.72
+ $X2=2.522 $Y2=2.72
r321 52 155 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.415 $Y=2.72
+ $X2=3.54 $Y2=2.72
r322 52 53 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3.415 $Y=2.72
+ $X2=2.67 $Y2=2.72
r323 48 51 27.3461 $w=2.93e-07 $l=7e-07 $layer=LI1_cond $X=2.522 $Y=1.64
+ $X2=2.522 $Y2=2.34
r324 46 152 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.522 $Y=2.635
+ $X2=2.522 $Y2=2.72
r325 46 51 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=2.522 $Y=2.635
+ $X2=2.522 $Y2=2.34
r326 42 45 36.6686 $w=2.18e-07 $l=7e-07 $layer=LI1_cond $X=1.445 $Y=1.64
+ $X2=1.445 $Y2=2.34
r327 40 93 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.445 $Y=2.635
+ $X2=1.445 $Y2=2.72
r328 40 45 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=1.445 $Y=2.635
+ $X2=1.445 $Y2=2.34
r329 36 39 36.4494 $w=2.13e-07 $l=6.8e-07 $layer=LI1_cond $X=0.407 $Y=1.66
+ $X2=0.407 $Y2=2.34
r330 34 90 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.407 $Y=2.635
+ $X2=0.407 $Y2=2.72
r331 34 39 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=0.407 $Y=2.635
+ $X2=0.407 $Y2=2.34
r332 11 86 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=9.975
+ $Y=1.485 $X2=10.12 $Y2=2
r333 10 82 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=9.035
+ $Y=1.485 $X2=9.18 $Y2=2
r334 9 78 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=8.095
+ $Y=1.485 $X2=8.24 $Y2=2
r335 8 74 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=7.155
+ $Y=1.485 $X2=7.3 $Y2=2
r336 7 70 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.215
+ $Y=1.485 $X2=6.36 $Y2=2
r337 6 66 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.275
+ $Y=1.485 $X2=5.42 $Y2=2
r338 5 62 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.335
+ $Y=1.485 $X2=4.48 $Y2=2
r339 4 56 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.395
+ $Y=1.485 $X2=3.54 $Y2=2
r340 3 51 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=1.485 $X2=2.46 $Y2=2.34
r341 3 48 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=1.485 $X2=2.46 $Y2=1.64
r342 2 45 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.275
+ $Y=1.485 $X2=1.42 $Y2=2.34
r343 2 42 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=1.275
+ $Y=1.485 $X2=1.42 $Y2=1.64
r344 1 39 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.305
+ $Y=1.485 $X2=0.43 $Y2=2.34
r345 1 36 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.305
+ $Y=1.485 $X2=0.43 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_16%A_585_297# 1 2 3 4 5 6 7 8 9 10 11 12
+ 13 14 15 16 17 52 54 56 60 62 66 68 72 74 78 80 84 86 90 92 96 98 100 101 102
+ 106 108 112 114 118 120 124 126 130 132 136 138 142 144 148 153 155 157 159
+ 161 163 165 170 171 172 173 174 175 176
r215 146 148 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=18.11 $Y=2.295
+ $X2=18.11 $Y2=1.96
r216 145 176 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=17.295 $Y=2.38
+ $X2=17.17 $Y2=2.38
r217 144 146 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=17.985 $Y=2.38
+ $X2=18.11 $Y2=2.295
r218 144 145 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=17.985 $Y=2.38
+ $X2=17.295 $Y2=2.38
r219 140 176 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=17.17 $Y=2.295
+ $X2=17.17 $Y2=2.38
r220 140 142 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=17.17 $Y=2.295
+ $X2=17.17 $Y2=1.96
r221 139 175 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.355 $Y=2.38
+ $X2=16.23 $Y2=2.38
r222 138 176 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=17.045 $Y=2.38
+ $X2=17.17 $Y2=2.38
r223 138 139 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=17.045 $Y=2.38
+ $X2=16.355 $Y2=2.38
r224 134 175 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.23 $Y=2.295
+ $X2=16.23 $Y2=2.38
r225 134 136 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=16.23 $Y=2.295
+ $X2=16.23 $Y2=1.96
r226 133 174 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.415 $Y=2.38
+ $X2=15.29 $Y2=2.38
r227 132 175 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.105 $Y=2.38
+ $X2=16.23 $Y2=2.38
r228 132 133 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=16.105 $Y=2.38
+ $X2=15.415 $Y2=2.38
r229 128 174 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=15.29 $Y=2.295
+ $X2=15.29 $Y2=2.38
r230 128 130 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=15.29 $Y=2.295
+ $X2=15.29 $Y2=1.96
r231 127 173 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.475 $Y=2.38
+ $X2=14.35 $Y2=2.38
r232 126 174 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.165 $Y=2.38
+ $X2=15.29 $Y2=2.38
r233 126 127 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=15.165 $Y=2.38
+ $X2=14.475 $Y2=2.38
r234 122 173 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=14.35 $Y=2.295
+ $X2=14.35 $Y2=2.38
r235 122 124 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=14.35 $Y=2.295
+ $X2=14.35 $Y2=1.96
r236 121 172 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.535 $Y=2.38
+ $X2=13.41 $Y2=2.38
r237 120 173 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.225 $Y=2.38
+ $X2=14.35 $Y2=2.38
r238 120 121 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=14.225 $Y=2.38
+ $X2=13.535 $Y2=2.38
r239 116 172 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.41 $Y=2.295
+ $X2=13.41 $Y2=2.38
r240 116 118 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=13.41 $Y=2.295
+ $X2=13.41 $Y2=1.96
r241 115 171 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.595 $Y=2.38
+ $X2=12.47 $Y2=2.38
r242 114 172 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.285 $Y=2.38
+ $X2=13.41 $Y2=2.38
r243 114 115 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=13.285 $Y=2.38
+ $X2=12.595 $Y2=2.38
r244 110 171 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.47 $Y=2.295
+ $X2=12.47 $Y2=2.38
r245 110 112 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=12.47 $Y=2.295
+ $X2=12.47 $Y2=1.96
r246 109 170 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.655 $Y=2.38
+ $X2=11.53 $Y2=2.38
r247 108 171 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.345 $Y=2.38
+ $X2=12.47 $Y2=2.38
r248 108 109 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=12.345 $Y=2.38
+ $X2=11.655 $Y2=2.38
r249 104 170 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.53 $Y=2.295
+ $X2=11.53 $Y2=2.38
r250 104 106 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=11.53 $Y=2.295
+ $X2=11.53 $Y2=1.96
r251 103 169 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.715 $Y=2.38
+ $X2=10.59 $Y2=2.38
r252 102 170 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.405 $Y=2.38
+ $X2=11.53 $Y2=2.38
r253 102 103 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.405 $Y=2.38
+ $X2=10.715 $Y2=2.38
r254 101 169 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.59 $Y=2.295
+ $X2=10.59 $Y2=2.38
r255 100 167 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=10.59 $Y=1.665
+ $X2=10.59 $Y2=1.56
r256 100 101 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=10.59 $Y=1.665
+ $X2=10.59 $Y2=2.295
r257 99 165 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=9.775 $Y=1.56
+ $X2=9.65 $Y2=1.56
r258 98 167 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=10.465 $Y=1.56
+ $X2=10.59 $Y2=1.56
r259 98 99 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=10.465 $Y=1.56
+ $X2=9.775 $Y2=1.56
r260 94 165 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=9.65 $Y=1.665
+ $X2=9.65 $Y2=1.56
r261 94 96 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=9.65 $Y=1.665
+ $X2=9.65 $Y2=2.3
r262 93 163 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=8.835 $Y=1.56
+ $X2=8.71 $Y2=1.56
r263 92 165 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=9.525 $Y=1.56
+ $X2=9.65 $Y2=1.56
r264 92 93 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=9.525 $Y=1.56
+ $X2=8.835 $Y2=1.56
r265 88 163 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=8.71 $Y=1.665
+ $X2=8.71 $Y2=1.56
r266 88 90 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=8.71 $Y=1.665
+ $X2=8.71 $Y2=2.3
r267 87 161 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=7.895 $Y=1.56
+ $X2=7.77 $Y2=1.56
r268 86 163 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=8.585 $Y=1.56
+ $X2=8.71 $Y2=1.56
r269 86 87 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=8.585 $Y=1.56
+ $X2=7.895 $Y2=1.56
r270 82 161 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=7.77 $Y=1.665
+ $X2=7.77 $Y2=1.56
r271 82 84 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=7.77 $Y=1.665
+ $X2=7.77 $Y2=2.3
r272 81 159 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=6.955 $Y=1.56
+ $X2=6.83 $Y2=1.56
r273 80 161 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=7.645 $Y=1.56
+ $X2=7.77 $Y2=1.56
r274 80 81 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=7.645 $Y=1.56
+ $X2=6.955 $Y2=1.56
r275 76 159 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=6.83 $Y=1.665
+ $X2=6.83 $Y2=1.56
r276 76 78 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=6.83 $Y=1.665
+ $X2=6.83 $Y2=2.3
r277 75 157 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=6.015 $Y=1.56
+ $X2=5.89 $Y2=1.56
r278 74 159 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=6.705 $Y=1.56
+ $X2=6.83 $Y2=1.56
r279 74 75 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=6.705 $Y=1.56
+ $X2=6.015 $Y2=1.56
r280 70 157 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=5.89 $Y=1.665
+ $X2=5.89 $Y2=1.56
r281 70 72 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=5.89 $Y=1.665
+ $X2=5.89 $Y2=2.3
r282 69 155 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=5.075 $Y=1.56
+ $X2=4.95 $Y2=1.56
r283 68 157 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=5.765 $Y=1.56
+ $X2=5.89 $Y2=1.56
r284 68 69 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=5.765 $Y=1.56
+ $X2=5.075 $Y2=1.56
r285 64 155 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=4.95 $Y=1.665
+ $X2=4.95 $Y2=1.56
r286 64 66 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=4.95 $Y=1.665
+ $X2=4.95 $Y2=2.3
r287 63 153 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=4.135 $Y=1.56
+ $X2=4.01 $Y2=1.56
r288 62 155 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=4.825 $Y=1.56
+ $X2=4.95 $Y2=1.56
r289 62 63 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=4.825 $Y=1.56
+ $X2=4.135 $Y2=1.56
r290 58 153 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=4.01 $Y=1.665
+ $X2=4.01 $Y2=1.56
r291 58 60 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=4.01 $Y=1.665
+ $X2=4.01 $Y2=2.3
r292 57 151 4.35048 $w=2.1e-07 $l=1.6e-07 $layer=LI1_cond $X=3.195 $Y=1.56
+ $X2=3.035 $Y2=1.56
r293 56 153 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=3.885 $Y=1.56
+ $X2=4.01 $Y2=1.56
r294 56 57 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=3.885 $Y=1.56
+ $X2=3.195 $Y2=1.56
r295 52 151 2.855 $w=3.2e-07 $l=1.05e-07 $layer=LI1_cond $X=3.035 $Y=1.665
+ $X2=3.035 $Y2=1.56
r296 52 54 22.8688 $w=3.18e-07 $l=6.35e-07 $layer=LI1_cond $X=3.035 $Y=1.665
+ $X2=3.035 $Y2=2.3
r297 17 148 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=17.965
+ $Y=1.485 $X2=18.11 $Y2=1.96
r298 16 142 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=17.025
+ $Y=1.485 $X2=17.17 $Y2=1.96
r299 15 136 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=16.085
+ $Y=1.485 $X2=16.23 $Y2=1.96
r300 14 130 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=15.145
+ $Y=1.485 $X2=15.29 $Y2=1.96
r301 13 124 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=14.205
+ $Y=1.485 $X2=14.35 $Y2=1.96
r302 12 118 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=13.265
+ $Y=1.485 $X2=13.41 $Y2=1.96
r303 11 112 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=12.325
+ $Y=1.485 $X2=12.47 $Y2=1.96
r304 10 106 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=11.385
+ $Y=1.485 $X2=11.53 $Y2=1.96
r305 9 169 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=10.445
+ $Y=1.485 $X2=10.59 $Y2=2.3
r306 9 167 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.445
+ $Y=1.485 $X2=10.59 $Y2=1.62
r307 8 165 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.505
+ $Y=1.485 $X2=9.65 $Y2=1.62
r308 8 96 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=9.505
+ $Y=1.485 $X2=9.65 $Y2=2.3
r309 7 163 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.565
+ $Y=1.485 $X2=8.71 $Y2=1.62
r310 7 90 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=8.565
+ $Y=1.485 $X2=8.71 $Y2=2.3
r311 6 161 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.625
+ $Y=1.485 $X2=7.77 $Y2=1.62
r312 6 84 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=7.625
+ $Y=1.485 $X2=7.77 $Y2=2.3
r313 5 159 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.685
+ $Y=1.485 $X2=6.83 $Y2=1.62
r314 5 78 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=6.685
+ $Y=1.485 $X2=6.83 $Y2=2.3
r315 4 157 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.745
+ $Y=1.485 $X2=5.89 $Y2=1.62
r316 4 72 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.745
+ $Y=1.485 $X2=5.89 $Y2=2.3
r317 3 155 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.805
+ $Y=1.485 $X2=4.95 $Y2=1.62
r318 3 66 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.805
+ $Y=1.485 $X2=4.95 $Y2=2.3
r319 2 153 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.865
+ $Y=1.485 $X2=4.01 $Y2=1.62
r320 2 60 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.865
+ $Y=1.485 $X2=4.01 $Y2=2.3
r321 1 151 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.485 $X2=3.07 $Y2=1.62
r322 1 54 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.485 $X2=3.07 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
+ 16 17 18 19 20 21 22 23 24 75 77 78 81 83 87 89 93 95 99 101 105 107 111 113
+ 117 119 123 127 129 133 137 139 143 147 149 153 157 159 163 167 169 173 177
+ 179 183 187 189 193 194 195 196 197 198 199 200 202 203 205 206 208 209 211
+ 212 214 215 217 218 220 222 225
c472 222 0 1.70671e-19 $X=17.64 $Y=0.39
r473 225 228 2.46131 $w=3.92e-07 $l=1.64085e-07 $layer=LI1_cond $X=17.91 $Y=1.54
+ $X2=18.037 $Y2=1.455
r474 225 228 0.111783 $w=5.33e-07 $l=5e-09 $layer=LI1_cond $X=18.037 $Y=1.45
+ $X2=18.037 $Y2=1.455
r475 224 225 12.1844 $w=5.33e-07 $l=5.45e-07 $layer=LI1_cond $X=18.037 $Y=0.905
+ $X2=18.037 $Y2=1.45
r476 222 224 12.6791 $w=3.82e-07 $l=5.805e-07 $layer=LI1_cond $X=17.64 $Y=0.49
+ $X2=18.037 $Y2=0.905
r477 190 218 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=16.865 $Y=0.815
+ $X2=16.675 $Y2=0.815
r478 189 222 10.2989 $w=3.82e-07 $l=4.18927e-07 $layer=LI1_cond $X=17.425
+ $Y=0.815 $X2=17.64 $Y2=0.49
r479 189 190 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=17.425 $Y=0.815
+ $X2=16.865 $Y2=0.815
r480 188 220 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.825 $Y=1.54
+ $X2=16.7 $Y2=1.54
r481 187 225 4.47094 $w=1.7e-07 $l=3.95e-07 $layer=LI1_cond $X=17.515 $Y=1.54
+ $X2=17.91 $Y2=1.54
r482 187 188 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=17.515 $Y=1.54
+ $X2=16.825 $Y2=1.54
r483 181 218 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=16.675 $Y=0.725
+ $X2=16.675 $Y2=0.815
r484 181 183 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=16.675 $Y=0.725
+ $X2=16.675 $Y2=0.39
r485 180 215 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=15.925 $Y=0.815
+ $X2=15.735 $Y2=0.815
r486 179 218 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=16.485 $Y=0.815
+ $X2=16.675 $Y2=0.815
r487 179 180 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=16.485 $Y=0.815
+ $X2=15.925 $Y2=0.815
r488 178 217 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.885 $Y=1.54
+ $X2=15.76 $Y2=1.54
r489 177 220 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.575 $Y=1.54
+ $X2=16.7 $Y2=1.54
r490 177 178 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=16.575 $Y=1.54
+ $X2=15.885 $Y2=1.54
r491 171 215 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=15.735 $Y=0.725
+ $X2=15.735 $Y2=0.815
r492 171 173 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=15.735 $Y=0.725
+ $X2=15.735 $Y2=0.39
r493 170 212 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=14.985 $Y=0.815
+ $X2=14.795 $Y2=0.815
r494 169 215 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=15.545 $Y=0.815
+ $X2=15.735 $Y2=0.815
r495 169 170 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=15.545 $Y=0.815
+ $X2=14.985 $Y2=0.815
r496 168 214 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.945 $Y=1.54
+ $X2=14.82 $Y2=1.54
r497 167 217 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.635 $Y=1.54
+ $X2=15.76 $Y2=1.54
r498 167 168 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=15.635 $Y=1.54
+ $X2=14.945 $Y2=1.54
r499 161 212 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=14.795 $Y=0.725
+ $X2=14.795 $Y2=0.815
r500 161 163 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=14.795 $Y=0.725
+ $X2=14.795 $Y2=0.39
r501 160 209 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=14.045 $Y=0.815
+ $X2=13.855 $Y2=0.815
r502 159 212 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=14.605 $Y=0.815
+ $X2=14.795 $Y2=0.815
r503 159 160 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=14.605 $Y=0.815
+ $X2=14.045 $Y2=0.815
r504 158 211 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.005 $Y=1.54
+ $X2=13.88 $Y2=1.54
r505 157 214 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.695 $Y=1.54
+ $X2=14.82 $Y2=1.54
r506 157 158 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=14.695 $Y=1.54
+ $X2=14.005 $Y2=1.54
r507 151 209 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=13.855 $Y=0.725
+ $X2=13.855 $Y2=0.815
r508 151 153 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=13.855 $Y=0.725
+ $X2=13.855 $Y2=0.39
r509 150 206 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=13.105 $Y=0.815
+ $X2=12.915 $Y2=0.815
r510 149 209 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=13.665 $Y=0.815
+ $X2=13.855 $Y2=0.815
r511 149 150 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=13.665 $Y=0.815
+ $X2=13.105 $Y2=0.815
r512 148 208 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.065 $Y=1.54
+ $X2=12.94 $Y2=1.54
r513 147 211 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.755 $Y=1.54
+ $X2=13.88 $Y2=1.54
r514 147 148 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=13.755 $Y=1.54
+ $X2=13.065 $Y2=1.54
r515 141 206 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=12.915 $Y=0.725
+ $X2=12.915 $Y2=0.815
r516 141 143 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=12.915 $Y=0.725
+ $X2=12.915 $Y2=0.39
r517 140 203 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=12.165 $Y=0.815
+ $X2=11.975 $Y2=0.815
r518 139 206 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=12.725 $Y=0.815
+ $X2=12.915 $Y2=0.815
r519 139 140 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=12.725 $Y=0.815
+ $X2=12.165 $Y2=0.815
r520 138 205 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.125 $Y=1.54
+ $X2=12 $Y2=1.54
r521 137 208 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.815 $Y=1.54
+ $X2=12.94 $Y2=1.54
r522 137 138 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=12.815 $Y=1.54
+ $X2=12.125 $Y2=1.54
r523 131 203 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=11.975 $Y=0.725
+ $X2=11.975 $Y2=0.815
r524 131 133 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=11.975 $Y=0.725
+ $X2=11.975 $Y2=0.39
r525 130 200 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=11.225 $Y=0.815
+ $X2=11.035 $Y2=0.815
r526 129 203 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=11.785 $Y=0.815
+ $X2=11.975 $Y2=0.815
r527 129 130 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=11.785 $Y=0.815
+ $X2=11.225 $Y2=0.815
r528 128 202 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.185 $Y=1.54
+ $X2=11.06 $Y2=1.54
r529 127 205 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.875 $Y=1.54
+ $X2=12 $Y2=1.54
r530 127 128 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.875 $Y=1.54
+ $X2=11.185 $Y2=1.54
r531 121 200 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=11.035 $Y=0.725
+ $X2=11.035 $Y2=0.815
r532 121 123 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=11.035 $Y=0.725
+ $X2=11.035 $Y2=0.39
r533 120 199 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=10.285 $Y=0.815
+ $X2=10.095 $Y2=0.815
r534 119 200 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=10.845 $Y=0.815
+ $X2=11.035 $Y2=0.815
r535 119 120 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=10.845 $Y=0.815
+ $X2=10.285 $Y2=0.815
r536 115 199 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=10.095 $Y=0.725
+ $X2=10.095 $Y2=0.815
r537 115 117 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=10.095 $Y=0.725
+ $X2=10.095 $Y2=0.39
r538 114 198 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=9.345 $Y=0.815
+ $X2=9.155 $Y2=0.815
r539 113 199 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=9.905 $Y=0.815
+ $X2=10.095 $Y2=0.815
r540 113 114 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=9.905 $Y=0.815
+ $X2=9.345 $Y2=0.815
r541 109 198 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=9.155 $Y=0.725
+ $X2=9.155 $Y2=0.815
r542 109 111 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=9.155 $Y=0.725
+ $X2=9.155 $Y2=0.39
r543 108 197 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=8.405 $Y=0.815
+ $X2=8.215 $Y2=0.815
r544 107 198 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=8.965 $Y=0.815
+ $X2=9.155 $Y2=0.815
r545 107 108 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=8.965 $Y=0.815
+ $X2=8.405 $Y2=0.815
r546 103 197 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=8.215 $Y=0.725
+ $X2=8.215 $Y2=0.815
r547 103 105 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=8.215 $Y=0.725
+ $X2=8.215 $Y2=0.39
r548 102 196 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=7.465 $Y=0.815
+ $X2=7.275 $Y2=0.815
r549 101 197 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=8.025 $Y=0.815
+ $X2=8.215 $Y2=0.815
r550 101 102 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=8.025 $Y=0.815
+ $X2=7.465 $Y2=0.815
r551 97 196 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=7.275 $Y=0.725
+ $X2=7.275 $Y2=0.815
r552 97 99 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.275 $Y=0.725
+ $X2=7.275 $Y2=0.39
r553 96 195 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.525 $Y=0.815
+ $X2=6.335 $Y2=0.815
r554 95 196 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=7.085 $Y=0.815
+ $X2=7.275 $Y2=0.815
r555 95 96 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=7.085 $Y=0.815
+ $X2=6.525 $Y2=0.815
r556 91 195 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=6.335 $Y=0.725
+ $X2=6.335 $Y2=0.815
r557 91 93 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.335 $Y=0.725
+ $X2=6.335 $Y2=0.39
r558 90 194 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.585 $Y=0.815
+ $X2=5.395 $Y2=0.815
r559 89 195 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.145 $Y=0.815
+ $X2=6.335 $Y2=0.815
r560 89 90 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=6.145 $Y=0.815
+ $X2=5.585 $Y2=0.815
r561 85 194 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=5.395 $Y=0.725
+ $X2=5.395 $Y2=0.815
r562 85 87 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.395 $Y=0.725
+ $X2=5.395 $Y2=0.39
r563 84 193 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.645 $Y=0.815
+ $X2=4.455 $Y2=0.815
r564 83 194 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.205 $Y=0.815
+ $X2=5.395 $Y2=0.815
r565 83 84 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=5.205 $Y=0.815
+ $X2=4.645 $Y2=0.815
r566 79 193 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=4.455 $Y=0.725
+ $X2=4.455 $Y2=0.815
r567 79 81 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.455 $Y=0.725
+ $X2=4.455 $Y2=0.39
r568 77 193 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.265 $Y=0.815
+ $X2=4.455 $Y2=0.815
r569 77 78 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.265 $Y=0.815
+ $X2=3.705 $Y2=0.815
r570 73 78 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=3.515 $Y=0.725
+ $X2=3.705 $Y2=0.815
r571 73 75 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.515 $Y=0.725
+ $X2=3.515 $Y2=0.39
r572 24 225 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=17.495
+ $Y=1.485 $X2=17.64 $Y2=1.62
r573 23 220 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=16.555
+ $Y=1.485 $X2=16.7 $Y2=1.62
r574 22 217 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=15.615
+ $Y=1.485 $X2=15.76 $Y2=1.62
r575 21 214 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=14.675
+ $Y=1.485 $X2=14.82 $Y2=1.62
r576 20 211 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=13.735
+ $Y=1.485 $X2=13.88 $Y2=1.62
r577 19 208 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=12.795
+ $Y=1.485 $X2=12.94 $Y2=1.62
r578 18 205 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=11.855
+ $Y=1.485 $X2=12 $Y2=1.62
r579 17 202 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=10.915
+ $Y=1.485 $X2=11.06 $Y2=1.62
r580 16 222 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=17.455
+ $Y=0.235 $X2=17.64 $Y2=0.39
r581 15 183 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=16.515
+ $Y=0.235 $X2=16.7 $Y2=0.39
r582 14 173 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=15.575
+ $Y=0.235 $X2=15.76 $Y2=0.39
r583 13 163 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=14.635
+ $Y=0.235 $X2=14.82 $Y2=0.39
r584 12 153 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=13.695
+ $Y=0.235 $X2=13.88 $Y2=0.39
r585 11 143 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=12.755
+ $Y=0.235 $X2=12.94 $Y2=0.39
r586 10 133 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=11.815
+ $Y=0.235 $X2=12 $Y2=0.39
r587 9 123 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=10.875
+ $Y=0.235 $X2=11.06 $Y2=0.39
r588 8 117 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=9.935
+ $Y=0.235 $X2=10.12 $Y2=0.39
r589 7 111 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=8.995
+ $Y=0.235 $X2=9.18 $Y2=0.39
r590 6 105 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=8.055
+ $Y=0.235 $X2=8.24 $Y2=0.39
r591 5 99 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=7.115
+ $Y=0.235 $X2=7.3 $Y2=0.39
r592 4 93 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=6.175
+ $Y=0.235 $X2=6.36 $Y2=0.39
r593 3 87 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=5.235
+ $Y=0.235 $X2=5.42 $Y2=0.39
r594 2 81 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.295
+ $Y=0.235 $X2=4.48 $Y2=0.39
r595 1 75 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.355
+ $Y=0.235 $X2=3.54 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 18 19 60 62 66 70 74 78 82 86 90 94 98 102 106 110 114 118 122 126
+ 130 132 134 137 138 140 141 143 144 146 147 149 150 152 153 155 156 158 159
+ 161 162 164 165 167 168 170 171 173 174 176 177 179 180 181 183 188 239 244
+ 247 250 254
c327 132 0 1.70671e-19 $X=18.16 $Y=0.085
r328 253 254 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.17 $Y=0
+ $X2=18.17 $Y2=0
r329 250 251 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r330 247 248 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r331 245 248 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.61 $Y2=0
r332 244 245 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r333 242 254 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=17.71 $Y=0
+ $X2=18.17 $Y2=0
r334 241 242 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=17.71 $Y=0
+ $X2=17.71 $Y2=0
r335 239 253 4.20444 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=18.025 $Y=0
+ $X2=18.212 $Y2=0
r336 239 241 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=18.025 $Y=0
+ $X2=17.71 $Y2=0
r337 238 242 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=16.79 $Y=0
+ $X2=17.71 $Y2=0
r338 237 238 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.79 $Y=0
+ $X2=16.79 $Y2=0
r339 235 238 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=15.87 $Y=0
+ $X2=16.79 $Y2=0
r340 234 235 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.87 $Y=0
+ $X2=15.87 $Y2=0
r341 232 235 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=14.95 $Y=0
+ $X2=15.87 $Y2=0
r342 231 232 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.95 $Y=0
+ $X2=14.95 $Y2=0
r343 229 232 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=14.03 $Y=0
+ $X2=14.95 $Y2=0
r344 228 229 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.03 $Y=0
+ $X2=14.03 $Y2=0
r345 226 229 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.11 $Y=0
+ $X2=14.03 $Y2=0
r346 225 226 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r347 223 226 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.19 $Y=0
+ $X2=13.11 $Y2=0
r348 222 223 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r349 220 223 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=12.19 $Y2=0
r350 219 220 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r351 217 220 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=11.27 $Y2=0
r352 216 217 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r353 214 217 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.35 $Y2=0
r354 213 214 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r355 211 214 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=9.43 $Y2=0
r356 210 211 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r357 208 211 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.51 $Y2=0
r358 207 208 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r359 205 208 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r360 204 205 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r361 202 205 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r362 201 202 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r363 199 202 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r364 198 199 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r365 196 199 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.83 $Y2=0
r366 196 251 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=2.99 $Y2=0
r367 195 196 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r368 193 250 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.155 $Y=0
+ $X2=2.88 $Y2=0
r369 193 195 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=3.155 $Y=0
+ $X2=3.91 $Y2=0
r370 192 251 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=2.99 $Y2=0
r371 192 248 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=1.61 $Y2=0
r372 191 192 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r373 189 247 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.865 $Y=0
+ $X2=1.715 $Y2=0
r374 189 191 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.865 $Y=0
+ $X2=2.53 $Y2=0
r375 188 250 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=2.605 $Y=0
+ $X2=2.88 $Y2=0
r376 188 191 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.605 $Y=0
+ $X2=2.53 $Y2=0
r377 183 244 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.485 $Y=0
+ $X2=0.675 $Y2=0
r378 183 185 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.485 $Y=0
+ $X2=0.23 $Y2=0
r379 181 245 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r380 181 185 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r381 179 237 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=17.085 $Y=0
+ $X2=16.79 $Y2=0
r382 179 180 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=17.085 $Y=0
+ $X2=17.17 $Y2=0
r383 178 241 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=17.255 $Y=0
+ $X2=17.71 $Y2=0
r384 178 180 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=17.255 $Y=0
+ $X2=17.17 $Y2=0
r385 176 234 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=16.145 $Y=0
+ $X2=15.87 $Y2=0
r386 176 177 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.145 $Y=0
+ $X2=16.23 $Y2=0
r387 175 237 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=16.315 $Y=0
+ $X2=16.79 $Y2=0
r388 175 177 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.315 $Y=0
+ $X2=16.23 $Y2=0
r389 173 231 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=15.205 $Y=0
+ $X2=14.95 $Y2=0
r390 173 174 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.205 $Y=0
+ $X2=15.29 $Y2=0
r391 172 234 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=15.375 $Y=0
+ $X2=15.87 $Y2=0
r392 172 174 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.375 $Y=0
+ $X2=15.29 $Y2=0
r393 170 228 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=14.265 $Y=0
+ $X2=14.03 $Y2=0
r394 170 171 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.265 $Y=0
+ $X2=14.35 $Y2=0
r395 169 231 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=14.435 $Y=0
+ $X2=14.95 $Y2=0
r396 169 171 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.435 $Y=0
+ $X2=14.35 $Y2=0
r397 167 225 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=13.325 $Y=0
+ $X2=13.11 $Y2=0
r398 167 168 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.325 $Y=0
+ $X2=13.41 $Y2=0
r399 166 228 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=13.495 $Y=0
+ $X2=14.03 $Y2=0
r400 166 168 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.495 $Y=0
+ $X2=13.41 $Y2=0
r401 164 222 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=12.385 $Y=0
+ $X2=12.19 $Y2=0
r402 164 165 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.385 $Y=0
+ $X2=12.47 $Y2=0
r403 163 225 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=12.555 $Y=0
+ $X2=13.11 $Y2=0
r404 163 165 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.555 $Y=0
+ $X2=12.47 $Y2=0
r405 161 219 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=11.445 $Y=0
+ $X2=11.27 $Y2=0
r406 161 162 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.445 $Y=0
+ $X2=11.53 $Y2=0
r407 160 222 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=11.615 $Y=0
+ $X2=12.19 $Y2=0
r408 160 162 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.615 $Y=0
+ $X2=11.53 $Y2=0
r409 158 216 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=10.505 $Y=0
+ $X2=10.35 $Y2=0
r410 158 159 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.505 $Y=0
+ $X2=10.59 $Y2=0
r411 157 219 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=10.675 $Y=0
+ $X2=11.27 $Y2=0
r412 157 159 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.675 $Y=0
+ $X2=10.59 $Y2=0
r413 155 213 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=9.565 $Y=0
+ $X2=9.43 $Y2=0
r414 155 156 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.565 $Y=0
+ $X2=9.65 $Y2=0
r415 154 216 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=9.735 $Y=0
+ $X2=10.35 $Y2=0
r416 154 156 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.735 $Y=0
+ $X2=9.65 $Y2=0
r417 152 210 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=8.625 $Y=0
+ $X2=8.51 $Y2=0
r418 152 153 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.625 $Y=0
+ $X2=8.71 $Y2=0
r419 151 213 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.795 $Y=0
+ $X2=9.43 $Y2=0
r420 151 153 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.795 $Y=0
+ $X2=8.71 $Y2=0
r421 149 207 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.685 $Y=0
+ $X2=7.59 $Y2=0
r422 149 150 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.685 $Y=0
+ $X2=7.77 $Y2=0
r423 148 210 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=7.855 $Y=0
+ $X2=8.51 $Y2=0
r424 148 150 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.855 $Y=0
+ $X2=7.77 $Y2=0
r425 146 204 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.745 $Y=0
+ $X2=6.67 $Y2=0
r426 146 147 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.745 $Y=0
+ $X2=6.83 $Y2=0
r427 145 207 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=6.915 $Y=0
+ $X2=7.59 $Y2=0
r428 145 147 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.915 $Y=0
+ $X2=6.83 $Y2=0
r429 143 201 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=5.805 $Y=0
+ $X2=5.75 $Y2=0
r430 143 144 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.805 $Y=0
+ $X2=5.89 $Y2=0
r431 142 204 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=5.975 $Y=0
+ $X2=6.67 $Y2=0
r432 142 144 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.975 $Y=0
+ $X2=5.89 $Y2=0
r433 140 198 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.865 $Y=0
+ $X2=4.83 $Y2=0
r434 140 141 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.865 $Y=0
+ $X2=4.95 $Y2=0
r435 139 201 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=5.035 $Y=0
+ $X2=5.75 $Y2=0
r436 139 141 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.035 $Y=0
+ $X2=4.95 $Y2=0
r437 137 195 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.925 $Y=0
+ $X2=3.91 $Y2=0
r438 137 138 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=0
+ $X2=4.01 $Y2=0
r439 136 198 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=4.095 $Y=0
+ $X2=4.83 $Y2=0
r440 136 138 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.095 $Y=0
+ $X2=4.01 $Y2=0
r441 132 253 3.08026 $w=2.7e-07 $l=1.07912e-07 $layer=LI1_cond $X=18.16 $Y=0.085
+ $X2=18.212 $Y2=0
r442 132 134 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=18.16 $Y=0.085
+ $X2=18.16 $Y2=0.39
r443 128 180 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=17.17 $Y=0.085
+ $X2=17.17 $Y2=0
r444 128 130 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=17.17 $Y=0.085
+ $X2=17.17 $Y2=0.39
r445 124 177 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.23 $Y=0.085
+ $X2=16.23 $Y2=0
r446 124 126 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=16.23 $Y=0.085
+ $X2=16.23 $Y2=0.39
r447 120 174 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.29 $Y=0.085
+ $X2=15.29 $Y2=0
r448 120 122 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=15.29 $Y=0.085
+ $X2=15.29 $Y2=0.39
r449 116 171 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.35 $Y=0.085
+ $X2=14.35 $Y2=0
r450 116 118 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=14.35 $Y=0.085
+ $X2=14.35 $Y2=0.39
r451 112 168 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.41 $Y=0.085
+ $X2=13.41 $Y2=0
r452 112 114 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=13.41 $Y=0.085
+ $X2=13.41 $Y2=0.39
r453 108 165 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.47 $Y=0.085
+ $X2=12.47 $Y2=0
r454 108 110 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=12.47 $Y=0.085
+ $X2=12.47 $Y2=0.39
r455 104 162 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.53 $Y=0.085
+ $X2=11.53 $Y2=0
r456 104 106 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=11.53 $Y=0.085
+ $X2=11.53 $Y2=0.39
r457 100 159 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.59 $Y=0.085
+ $X2=10.59 $Y2=0
r458 100 102 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.59 $Y=0.085
+ $X2=10.59 $Y2=0.39
r459 96 156 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.65 $Y=0.085
+ $X2=9.65 $Y2=0
r460 96 98 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.65 $Y=0.085
+ $X2=9.65 $Y2=0.39
r461 92 153 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.71 $Y=0.085
+ $X2=8.71 $Y2=0
r462 92 94 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.71 $Y=0.085
+ $X2=8.71 $Y2=0.39
r463 88 150 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.77 $Y=0.085
+ $X2=7.77 $Y2=0
r464 88 90 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.77 $Y=0.085
+ $X2=7.77 $Y2=0.39
r465 84 147 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.83 $Y=0.085
+ $X2=6.83 $Y2=0
r466 84 86 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.83 $Y=0.085
+ $X2=6.83 $Y2=0.39
r467 80 144 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.89 $Y=0.085
+ $X2=5.89 $Y2=0
r468 80 82 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.89 $Y=0.085
+ $X2=5.89 $Y2=0.39
r469 76 141 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.95 $Y=0.085
+ $X2=4.95 $Y2=0
r470 76 78 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.95 $Y=0.085
+ $X2=4.95 $Y2=0.39
r471 72 138 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.01 $Y=0.085
+ $X2=4.01 $Y2=0
r472 72 74 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.01 $Y=0.085
+ $X2=4.01 $Y2=0.39
r473 68 250 2.31338 $w=5.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=0.085
+ $X2=2.88 $Y2=0
r474 68 70 6.6328 $w=5.48e-07 $l=3.05e-07 $layer=LI1_cond $X=2.88 $Y=0.085
+ $X2=2.88 $Y2=0.39
r475 64 247 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.715 $Y=0.085
+ $X2=1.715 $Y2=0
r476 64 66 11.7165 $w=2.98e-07 $l=3.05e-07 $layer=LI1_cond $X=1.715 $Y=0.085
+ $X2=1.715 $Y2=0.39
r477 63 244 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.865 $Y=0
+ $X2=0.675 $Y2=0
r478 62 247 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.565 $Y=0
+ $X2=1.715 $Y2=0
r479 62 63 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.565 $Y=0 $X2=0.865
+ $Y2=0
r480 58 244 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.675 $Y=0.085
+ $X2=0.675 $Y2=0
r481 58 60 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=0.675 $Y=0.085
+ $X2=0.675 $Y2=0.39
r482 19 134 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=17.975
+ $Y=0.235 $X2=18.11 $Y2=0.39
r483 18 130 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=16.985
+ $Y=0.235 $X2=17.17 $Y2=0.39
r484 17 126 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=16.045
+ $Y=0.235 $X2=16.23 $Y2=0.39
r485 16 122 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=15.105
+ $Y=0.235 $X2=15.29 $Y2=0.39
r486 15 118 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=14.165
+ $Y=0.235 $X2=14.35 $Y2=0.39
r487 14 114 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=13.225
+ $Y=0.235 $X2=13.41 $Y2=0.39
r488 13 110 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=12.285
+ $Y=0.235 $X2=12.47 $Y2=0.39
r489 12 106 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=11.345
+ $Y=0.235 $X2=11.53 $Y2=0.39
r490 11 102 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=10.455
+ $Y=0.235 $X2=10.59 $Y2=0.39
r491 10 98 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=9.465
+ $Y=0.235 $X2=9.65 $Y2=0.39
r492 9 94 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=8.525
+ $Y=0.235 $X2=8.71 $Y2=0.39
r493 8 90 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=7.585
+ $Y=0.235 $X2=7.77 $Y2=0.39
r494 7 86 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=6.645
+ $Y=0.235 $X2=6.83 $Y2=0.39
r495 6 82 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=5.705
+ $Y=0.235 $X2=5.89 $Y2=0.39
r496 5 78 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.765
+ $Y=0.235 $X2=4.95 $Y2=0.39
r497 4 74 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=3.825
+ $Y=0.235 $X2=4.01 $Y2=0.39
r498 3 70 45.5 $w=1.7e-07 $l=5.47037e-07 $layer=licon1_NDIFF $count=4 $X=2.595
+ $Y=0.235 $X2=3.07 $Y2=0.39
r499 2 66 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.505
+ $Y=0.235 $X2=1.69 $Y2=0.39
r500 1 60 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.525
+ $Y=0.235 $X2=0.65 $Y2=0.39
.ends

