* File: sky130_fd_sc_hdll__nand3b_1.pxi.spice
* Created: Thu Aug 27 19:13:58 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND3B_1%A_N N_A_N_c_44_n N_A_N_M1000_g N_A_N_c_45_n
+ N_A_N_M1003_g A_N PM_SKY130_FD_SC_HDLL__NAND3B_1%A_N
x_PM_SKY130_FD_SC_HDLL__NAND3B_1%C N_C_c_70_n N_C_M1005_g N_C_c_71_n N_C_M1006_g
+ C C PM_SKY130_FD_SC_HDLL__NAND3B_1%C
x_PM_SKY130_FD_SC_HDLL__NAND3B_1%B N_B_c_97_n N_B_M1001_g N_B_c_98_n N_B_M1002_g
+ B B PM_SKY130_FD_SC_HDLL__NAND3B_1%B
x_PM_SKY130_FD_SC_HDLL__NAND3B_1%A_53_93# N_A_53_93#_M1003_s N_A_53_93#_M1000_s
+ N_A_53_93#_c_128_n N_A_53_93#_M1007_g N_A_53_93#_c_129_n N_A_53_93#_M1004_g
+ N_A_53_93#_c_130_n N_A_53_93#_c_139_n N_A_53_93#_c_131_n N_A_53_93#_c_132_n
+ N_A_53_93#_c_135_n PM_SKY130_FD_SC_HDLL__NAND3B_1%A_53_93#
x_PM_SKY130_FD_SC_HDLL__NAND3B_1%VPWR N_VPWR_M1000_d N_VPWR_M1001_d
+ N_VPWR_c_190_n N_VPWR_c_191_n N_VPWR_c_192_n N_VPWR_c_193_n N_VPWR_c_194_n
+ N_VPWR_c_195_n VPWR N_VPWR_c_196_n N_VPWR_c_189_n
+ PM_SKY130_FD_SC_HDLL__NAND3B_1%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND3B_1%Y N_Y_M1004_d N_Y_M1005_d N_Y_M1007_d
+ N_Y_c_231_n N_Y_c_233_n N_Y_c_237_n N_Y_c_239_n Y Y Y Y Y Y N_Y_c_226_n Y
+ PM_SKY130_FD_SC_HDLL__NAND3B_1%Y
x_PM_SKY130_FD_SC_HDLL__NAND3B_1%VGND N_VGND_M1003_d N_VGND_c_271_n
+ N_VGND_c_272_n N_VGND_c_273_n VGND N_VGND_c_274_n N_VGND_c_275_n
+ PM_SKY130_FD_SC_HDLL__NAND3B_1%VGND
cc_1 VNB N_A_N_c_44_n 0.0286128f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.41
cc_2 VNB N_A_N_c_45_n 0.0216557f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=0.995
cc_3 VNB A_N 0.00282637f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_4 VNB N_C_c_70_n 0.0232617f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.41
cc_5 VNB N_C_c_71_n 0.020135f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=0.995
cc_6 VNB C 0.00258765f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_7 VNB N_B_c_97_n 0.0201021f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.41
cc_8 VNB N_B_c_98_n 0.0175095f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=0.995
cc_9 VNB B 0.00247822f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_10 VNB N_A_53_93#_c_128_n 0.0244367f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_11 VNB N_A_53_93#_c_129_n 0.02003f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_12 VNB N_A_53_93#_c_130_n 0.0234199f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.16
cc_13 VNB N_A_53_93#_c_131_n 0.00221371f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_53_93#_c_132_n 0.0228672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VPWR_c_189_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_Y_c_226_n 0.011802f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB Y 0.039017f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_271_n 0.0107731f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=0.675
cc_19 VNB N_VGND_c_272_n 0.0225153f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.16
cc_20 VNB N_VGND_c_273_n 0.00631563f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_21 VNB N_VGND_c_274_n 0.0455953f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_275_n 0.168737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VPB N_A_N_c_44_n 0.0355147f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.41
cc_24 VPB A_N 0.00205187f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_25 VPB N_C_c_70_n 0.0310531f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.41
cc_26 VPB C 8.11817e-19 $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_27 VPB N_B_c_97_n 0.0251308f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.41
cc_28 VPB B 6.32037e-19 $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_29 VPB N_A_53_93#_c_128_n 0.0285551f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_30 VPB N_A_53_93#_c_130_n 0.0150052f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.16
cc_31 VPB N_A_53_93#_c_135_n 0.023627f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_190_n 0.0232531f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=1.16
cc_33 VPB N_VPWR_c_191_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_192_n 0.026328f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_193_n 0.00477947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_194_n 0.0209591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_195_n 0.0031889f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_196_n 0.02235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_189_n 0.0559351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB Y 0.00802402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB Y 0.0380712f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB Y 0.0104363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 N_A_N_c_44_n N_C_c_70_n 0.0344709f $X=0.625 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_44 A_N N_C_c_70_n 0.00222602f $X=0.605 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_45 N_A_N_c_45_n N_C_c_71_n 0.0174573f $X=0.65 $Y=0.995 $X2=0 $Y2=0
cc_46 N_A_N_c_44_n C 2.99721e-19 $X=0.625 $Y=1.41 $X2=0 $Y2=0
cc_47 A_N C 0.0244095f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_48 N_A_N_c_44_n N_A_53_93#_c_130_n 0.0152894f $X=0.625 $Y=1.41 $X2=0 $Y2=0
cc_49 N_A_N_c_45_n N_A_53_93#_c_130_n 0.0049454f $X=0.65 $Y=0.995 $X2=0 $Y2=0
cc_50 A_N N_A_53_93#_c_130_n 0.0251381f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_51 N_A_N_c_45_n N_A_53_93#_c_139_n 0.0104712f $X=0.65 $Y=0.995 $X2=0 $Y2=0
cc_52 N_A_N_c_44_n N_A_53_93#_c_132_n 0.00672937f $X=0.625 $Y=1.41 $X2=0 $Y2=0
cc_53 N_A_N_c_45_n N_A_53_93#_c_132_n 0.00463471f $X=0.65 $Y=0.995 $X2=0 $Y2=0
cc_54 A_N N_A_53_93#_c_132_n 0.0258008f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_55 N_A_N_c_44_n N_A_53_93#_c_135_n 0.00510605f $X=0.625 $Y=1.41 $X2=0 $Y2=0
cc_56 A_N N_A_53_93#_c_135_n 0.00371578f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_57 N_A_N_c_44_n N_VPWR_c_190_n 0.00545995f $X=0.625 $Y=1.41 $X2=0 $Y2=0
cc_58 A_N N_VPWR_c_190_n 0.00505451f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_59 N_A_N_c_44_n N_VPWR_c_192_n 0.00393512f $X=0.625 $Y=1.41 $X2=0 $Y2=0
cc_60 N_A_N_c_44_n N_VPWR_c_189_n 0.00500987f $X=0.625 $Y=1.41 $X2=0 $Y2=0
cc_61 N_A_N_c_45_n N_VGND_c_271_n 0.00354897f $X=0.65 $Y=0.995 $X2=0 $Y2=0
cc_62 N_A_N_c_45_n N_VGND_c_272_n 0.00393318f $X=0.65 $Y=0.995 $X2=0 $Y2=0
cc_63 N_A_N_c_45_n N_VGND_c_275_n 0.00512902f $X=0.65 $Y=0.995 $X2=0 $Y2=0
cc_64 N_C_c_70_n N_B_c_97_n 0.0344916f $X=1.16 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_65 C N_B_c_97_n 0.00199566f $X=1.115 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_66 N_C_c_71_n N_B_c_98_n 0.0362361f $X=1.185 $Y=0.995 $X2=0 $Y2=0
cc_67 N_C_c_70_n B 3.28206e-19 $X=1.16 $Y=1.41 $X2=0 $Y2=0
cc_68 C B 0.0242038f $X=1.115 $Y=1.105 $X2=0 $Y2=0
cc_69 N_C_c_70_n N_A_53_93#_c_139_n 0.00442168f $X=1.16 $Y=1.41 $X2=0 $Y2=0
cc_70 N_C_c_71_n N_A_53_93#_c_139_n 0.0126873f $X=1.185 $Y=0.995 $X2=0 $Y2=0
cc_71 C N_A_53_93#_c_139_n 0.0194328f $X=1.115 $Y=1.105 $X2=0 $Y2=0
cc_72 N_C_c_70_n N_VPWR_c_190_n 0.00998255f $X=1.16 $Y=1.41 $X2=0 $Y2=0
cc_73 N_C_c_70_n N_VPWR_c_194_n 0.00597712f $X=1.16 $Y=1.41 $X2=0 $Y2=0
cc_74 N_C_c_70_n N_VPWR_c_189_n 0.0113258f $X=1.16 $Y=1.41 $X2=0 $Y2=0
cc_75 N_C_c_70_n N_Y_c_231_n 0.00339981f $X=1.16 $Y=1.41 $X2=0 $Y2=0
cc_76 C N_Y_c_231_n 0.010315f $X=1.115 $Y=1.105 $X2=0 $Y2=0
cc_77 N_C_c_70_n N_Y_c_233_n 0.0120097f $X=1.16 $Y=1.41 $X2=0 $Y2=0
cc_78 N_C_c_71_n N_VGND_c_271_n 0.00482545f $X=1.185 $Y=0.995 $X2=0 $Y2=0
cc_79 N_C_c_71_n N_VGND_c_274_n 0.00428022f $X=1.185 $Y=0.995 $X2=0 $Y2=0
cc_80 N_C_c_71_n N_VGND_c_275_n 0.0071845f $X=1.185 $Y=0.995 $X2=0 $Y2=0
cc_81 N_B_c_97_n N_A_53_93#_c_128_n 0.0468945f $X=1.64 $Y=1.41 $X2=0 $Y2=0
cc_82 B N_A_53_93#_c_128_n 0.00197866f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_83 N_B_c_98_n N_A_53_93#_c_129_n 0.0342921f $X=1.665 $Y=0.995 $X2=0 $Y2=0
cc_84 N_B_c_97_n N_A_53_93#_c_139_n 0.00297968f $X=1.64 $Y=1.41 $X2=0 $Y2=0
cc_85 N_B_c_98_n N_A_53_93#_c_139_n 0.0123947f $X=1.665 $Y=0.995 $X2=0 $Y2=0
cc_86 B N_A_53_93#_c_139_n 0.0161005f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_87 N_B_c_97_n N_A_53_93#_c_131_n 3.45136e-19 $X=1.64 $Y=1.41 $X2=0 $Y2=0
cc_88 N_B_c_98_n N_A_53_93#_c_131_n 0.00336667f $X=1.665 $Y=0.995 $X2=0 $Y2=0
cc_89 B N_A_53_93#_c_131_n 0.0216895f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_90 N_B_c_97_n N_VPWR_c_191_n 0.0053108f $X=1.64 $Y=1.41 $X2=0 $Y2=0
cc_91 N_B_c_97_n N_VPWR_c_194_n 0.00688798f $X=1.64 $Y=1.41 $X2=0 $Y2=0
cc_92 N_B_c_97_n N_VPWR_c_189_n 0.0123115f $X=1.64 $Y=1.41 $X2=0 $Y2=0
cc_93 N_B_c_97_n N_Y_c_231_n 0.00192027f $X=1.64 $Y=1.41 $X2=0 $Y2=0
cc_94 B N_Y_c_231_n 0.00188714f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_95 N_B_c_97_n N_Y_c_233_n 0.0101748f $X=1.64 $Y=1.41 $X2=0 $Y2=0
cc_96 N_B_c_97_n N_Y_c_237_n 0.0145431f $X=1.64 $Y=1.41 $X2=0 $Y2=0
cc_97 B N_Y_c_237_n 0.0150619f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_98 N_B_c_98_n N_Y_c_239_n 0.00121092f $X=1.665 $Y=0.995 $X2=0 $Y2=0
cc_99 N_B_c_97_n Y 6.57811e-19 $X=1.64 $Y=1.41 $X2=0 $Y2=0
cc_100 N_B_c_98_n N_VGND_c_274_n 0.00428022f $X=1.665 $Y=0.995 $X2=0 $Y2=0
cc_101 N_B_c_98_n N_VGND_c_275_n 0.00626245f $X=1.665 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A_53_93#_c_139_n N_VPWR_c_190_n 0.00529132f $X=2 $Y=0.74 $X2=0 $Y2=0
cc_103 N_A_53_93#_c_135_n N_VPWR_c_190_n 0.00114603f $X=0.39 $Y=1.76 $X2=0 $Y2=0
cc_104 N_A_53_93#_c_128_n N_VPWR_c_191_n 0.00467386f $X=2.12 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A_53_93#_c_128_n N_VPWR_c_196_n 0.00582531f $X=2.12 $Y=1.41 $X2=0 $Y2=0
cc_106 N_A_53_93#_c_128_n N_VPWR_c_189_n 0.0107197f $X=2.12 $Y=1.41 $X2=0 $Y2=0
cc_107 N_A_53_93#_c_135_n N_VPWR_c_189_n 0.0161088f $X=0.39 $Y=1.76 $X2=0 $Y2=0
cc_108 N_A_53_93#_c_139_n N_Y_c_231_n 0.00490078f $X=2 $Y=0.74 $X2=0 $Y2=0
cc_109 N_A_53_93#_c_128_n N_Y_c_233_n 6.17548e-19 $X=2.12 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A_53_93#_c_128_n N_Y_c_237_n 0.0105727f $X=2.12 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A_53_93#_c_139_n N_Y_c_237_n 0.00490308f $X=2 $Y=0.74 $X2=0 $Y2=0
cc_112 N_A_53_93#_c_131_n N_Y_c_237_n 0.00879284f $X=2.085 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_53_93#_c_129_n N_Y_c_239_n 0.0074527f $X=2.14 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A_53_93#_c_139_n N_Y_c_239_n 0.00623159f $X=2 $Y=0.74 $X2=0 $Y2=0
cc_115 N_A_53_93#_c_128_n Y 0.00240634f $X=2.12 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A_53_93#_c_131_n Y 0.00710219f $X=2.085 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A_53_93#_c_128_n Y 0.0137405f $X=2.12 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A_53_93#_c_128_n Y 0.0130166f $X=2.12 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_53_93#_c_129_n Y 0.00690756f $X=2.14 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A_53_93#_c_131_n Y 0.0331145f $X=2.085 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_53_93#_c_139_n N_VGND_M1003_d 0.00726083f $X=2 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_122 N_A_53_93#_c_139_n N_VGND_c_271_n 0.020804f $X=2 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A_53_93#_c_132_n N_VGND_c_271_n 0.00183174f $X=0.51 $Y=0.635 $X2=0
+ $Y2=0
cc_124 N_A_53_93#_c_139_n N_VGND_c_272_n 0.00330937f $X=2 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A_53_93#_c_132_n N_VGND_c_272_n 0.01312f $X=0.51 $Y=0.635 $X2=0 $Y2=0
cc_126 N_A_53_93#_c_129_n N_VGND_c_274_n 0.0038821f $X=2.14 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_53_93#_c_139_n N_VGND_c_274_n 0.015259f $X=2 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A_53_93#_c_129_n N_VGND_c_275_n 0.00674365f $X=2.14 $Y=0.995 $X2=0
+ $Y2=0
cc_129 N_A_53_93#_c_139_n N_VGND_c_275_n 0.0357816f $X=2 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_53_93#_c_132_n N_VGND_c_275_n 0.0143027f $X=0.51 $Y=0.635 $X2=0 $Y2=0
cc_131 N_A_53_93#_c_139_n A_252_47# 0.00773946f $X=2 $Y=0.74 $X2=-0.19 $Y2=-0.24
cc_132 N_A_53_93#_c_139_n A_348_47# 0.00768771f $X=2 $Y=0.74 $X2=-0.19 $Y2=-0.24
cc_133 N_A_53_93#_c_131_n A_348_47# 7.56176e-19 $X=2.085 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_134 N_VPWR_c_189_n N_Y_M1005_d 0.00239291f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_135 N_VPWR_c_189_n N_Y_M1007_d 0.00233913f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_136 N_VPWR_c_190_n N_Y_c_231_n 0.0137304f $X=0.925 $Y=1.66 $X2=0 $Y2=0
cc_137 N_VPWR_c_190_n N_Y_c_233_n 0.0614133f $X=0.925 $Y=1.66 $X2=0 $Y2=0
cc_138 N_VPWR_c_191_n N_Y_c_233_n 0.0372693f $X=1.875 $Y=2 $X2=0 $Y2=0
cc_139 N_VPWR_c_194_n N_Y_c_233_n 0.0223771f $X=1.79 $Y=2.72 $X2=0 $Y2=0
cc_140 N_VPWR_c_189_n N_Y_c_233_n 0.0140558f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_141 N_VPWR_M1001_d N_Y_c_237_n 0.00601623f $X=1.73 $Y=1.485 $X2=0 $Y2=0
cc_142 N_VPWR_c_191_n N_Y_c_237_n 0.0136682f $X=1.875 $Y=2 $X2=0 $Y2=0
cc_143 N_VPWR_c_191_n Y 0.0484016f $X=1.875 $Y=2 $X2=0 $Y2=0
cc_144 N_VPWR_c_196_n Y 0.0362356f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_145 N_VPWR_c_189_n Y 0.0204782f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_146 N_Y_c_239_n N_VGND_c_274_n 0.0162164f $X=2.41 $Y=0.37 $X2=0 $Y2=0
cc_147 N_Y_c_226_n N_VGND_c_274_n 0.0188755f $X=2.542 $Y=0.485 $X2=0 $Y2=0
cc_148 N_Y_M1004_d N_VGND_c_275_n 0.0022662f $X=2.215 $Y=0.235 $X2=0 $Y2=0
cc_149 N_Y_c_239_n N_VGND_c_275_n 0.0100352f $X=2.41 $Y=0.37 $X2=0 $Y2=0
cc_150 N_Y_c_226_n N_VGND_c_275_n 0.0102056f $X=2.542 $Y=0.485 $X2=0 $Y2=0
cc_151 N_VGND_c_275_n A_252_47# 0.00394943f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24
cc_152 N_VGND_c_275_n A_348_47# 0.00388865f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24
