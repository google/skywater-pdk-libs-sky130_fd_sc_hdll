* File: sky130_fd_sc_hdll__clkmux2_4.pex.spice
* Created: Thu Aug 27 19:03:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_4%A_79_199# 1 2 7 9 12 16 18 20 21 23 26
+ 30 32 34 37 40 41 43 46 48 52 54 62
c133 54 0 1.9931e-19 $X=2.902 $Y=0.54
c134 52 0 1.80039e-19 $X=4.05 $Y=2.04
r135 61 62 4.57182 $w=3.69e-07 $l=3.5e-08 $layer=POLY_cond $X=1.87 $Y=1.202
+ $X2=1.905 $Y2=1.202
r136 60 61 54.8618 $w=3.69e-07 $l=4.2e-07 $layer=POLY_cond $X=1.45 $Y=1.202
+ $X2=1.87 $Y2=1.202
r137 59 60 1.95935 $w=3.69e-07 $l=1.5e-08 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.45 $Y2=1.202
r138 58 59 61.393 $w=3.69e-07 $l=4.7e-07 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=1.435 $Y2=1.202
r139 57 58 4.57182 $w=3.69e-07 $l=3.5e-08 $layer=POLY_cond $X=0.93 $Y=1.202
+ $X2=0.965 $Y2=1.202
r140 56 57 54.8618 $w=3.69e-07 $l=4.2e-07 $layer=POLY_cond $X=0.51 $Y=1.202
+ $X2=0.93 $Y2=1.202
r141 55 56 1.95935 $w=3.69e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.51 $Y2=1.202
r142 50 52 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=3.335 $Y=2.04
+ $X2=4.05 $Y2=2.04
r143 48 50 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.99 $Y=2.04
+ $X2=3.335 $Y2=2.04
r144 44 54 3.49088 $w=2.67e-07 $l=1.4026e-07 $layer=LI1_cond $X=2.99 $Y=0.437
+ $X2=2.902 $Y2=0.54
r145 44 46 13.4189 $w=3.63e-07 $l=4.25e-07 $layer=LI1_cond $X=2.99 $Y=0.437
+ $X2=3.415 $Y2=0.437
r146 43 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.905 $Y=1.955
+ $X2=2.99 $Y2=2.04
r147 42 54 3.01551 $w=1.7e-07 $l=2.86496e-07 $layer=LI1_cond $X=2.905 $Y=0.825
+ $X2=2.902 $Y2=0.54
r148 42 43 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=2.905 $Y=0.825
+ $X2=2.905 $Y2=1.955
r149 40 54 3.49088 $w=2.67e-07 $l=2.39583e-07 $layer=LI1_cond $X=2.815 $Y=0.74
+ $X2=2.902 $Y2=0.54
r150 40 41 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.815 $Y=0.74
+ $X2=2.085 $Y2=0.74
r151 38 62 12.4092 $w=3.69e-07 $l=9.5e-08 $layer=POLY_cond $X=2 $Y=1.202
+ $X2=1.905 $Y2=1.202
r152 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2 $Y=1.16
+ $X2=2 $Y2=1.16
r153 35 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2 $Y=0.825
+ $X2=2.085 $Y2=0.74
r154 35 37 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2 $Y=0.825 $X2=2
+ $Y2=1.16
r155 32 62 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r156 32 34 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r157 28 61 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.87 $Y=0.995
+ $X2=1.87 $Y2=1.202
r158 28 30 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=1.87 $Y=0.995
+ $X2=1.87 $Y2=0.495
r159 24 60 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.45 $Y=0.995
+ $X2=1.45 $Y2=1.202
r160 24 26 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=1.45 $Y=0.995
+ $X2=1.45 $Y2=0.495
r161 21 59 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r162 21 23 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r163 18 58 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r164 18 20 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r165 14 57 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.93 $Y=0.995
+ $X2=0.93 $Y2=1.202
r166 14 16 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.93 $Y=0.995
+ $X2=0.93 $Y2=0.495
r167 10 56 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.51 $Y=0.995
+ $X2=0.51 $Y2=1.202
r168 10 12 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.51 $Y=0.995
+ $X2=0.51 $Y2=0.495
r169 7 55 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r170 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r171 2 52 400 $w=1.7e-07 $l=1.07949e-06 $layer=licon1_PDIFF $count=1 $X=3.19
+ $Y=1.545 $X2=4.05 $Y2=2.04
r172 2 50 400 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=1 $X=3.19
+ $Y=1.545 $X2=3.335 $Y2=2.04
r173 1 46 182 $w=1.7e-07 $l=3.94968e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.235 $X2=3.415 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_4%S 1 3 6 8 10 13 16 17 18 19 20 21 23 27
+ 31 32
c95 16 0 1.20693e-19 $X=2.55 $Y=2.295
r96 31 32 13.2166 $w=3.58e-07 $l=3.33e-07 $layer=LI1_cond $X=4.852 $Y=1.535
+ $X2=5.185 $Y2=1.535
r97 27 30 7.79239 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=2.512 $Y=1.16
+ $X2=2.512 $Y2=1.325
r98 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.48
+ $Y=1.16 $X2=2.48 $Y2=1.16
r99 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.27
+ $Y=1.22 $X2=5.27 $Y2=1.22
r100 21 32 3.40825 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=5.28 $Y=1.44
+ $X2=5.28 $Y2=1.535
r101 21 23 12.8421 $w=1.88e-07 $l=2.2e-07 $layer=LI1_cond $X=5.28 $Y=1.44
+ $X2=5.28 $Y2=1.22
r102 19 31 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.71 $Y=1.63
+ $X2=4.71 $Y2=1.535
r103 19 20 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.71 $Y=1.63
+ $X2=4.71 $Y2=2.295
r104 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.625 $Y=2.38
+ $X2=4.71 $Y2=2.295
r105 17 18 128.85 $w=1.68e-07 $l=1.975e-06 $layer=LI1_cond $X=4.625 $Y=2.38
+ $X2=2.65 $Y2=2.38
r106 16 18 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.55 $Y=2.295
+ $X2=2.65 $Y2=2.38
r107 16 30 53.7909 $w=1.98e-07 $l=9.7e-07 $layer=LI1_cond $X=2.55 $Y=2.295
+ $X2=2.55 $Y2=1.325
r108 11 24 39.2931 $w=2.55e-07 $l=1.88348e-07 $layer=POLY_cond $X=5.32 $Y=1.055
+ $X2=5.27 $Y2=1.22
r109 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.32 $Y=1.055
+ $X2=5.32 $Y2=0.495
r110 8 24 51.486 $w=2.55e-07 $l=2.62202e-07 $layer=POLY_cond $X=5.295 $Y=1.47
+ $X2=5.27 $Y2=1.22
r111 8 10 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=5.295 $Y=1.47
+ $X2=5.295 $Y2=2.015
r112 4 28 39.2931 $w=2.55e-07 $l=1.94808e-07 $layer=POLY_cond $X=2.55 $Y=0.995
+ $X2=2.485 $Y2=1.16
r113 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.55 $Y=0.995
+ $X2=2.55 $Y2=0.445
r114 1 28 62.8272 $w=2.55e-07 $l=3.29393e-07 $layer=POLY_cond $X=2.525 $Y=1.47
+ $X2=2.485 $Y2=1.16
r115 1 3 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.525 $Y=1.47
+ $X2=2.525 $Y2=2.015
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_4%A1 3 5 7 10 11 13 14 16 17
c69 5 0 1.3232e-19 $X=4.285 $Y=1.47
r70 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.25
+ $Y=1.22 $X2=4.25 $Y2=1.22
r71 17 26 1.19218 $w=2.88e-07 $l=3e-08 $layer=LI1_cond $X=4.31 $Y=1.19 $X2=4.31
+ $Y2=1.22
r72 16 17 13.5114 $w=2.88e-07 $l=3.4e-07 $layer=LI1_cond $X=4.31 $Y=0.85
+ $X2=4.31 $Y2=1.19
r73 15 26 15.6971 $w=2.88e-07 $l=3.95e-07 $layer=LI1_cond $X=4.31 $Y=1.615
+ $X2=4.31 $Y2=1.22
r74 13 15 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=4.165 $Y=1.7
+ $X2=4.31 $Y2=1.615
r75 13 14 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=4.165 $Y=1.7
+ $X2=3.33 $Y2=1.7
r76 11 20 45.5456 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=3.245 $Y=0.975
+ $X2=3.04 $Y2=0.975
r77 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.245
+ $Y=0.975 $X2=3.245 $Y2=0.975
r78 8 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.245 $Y=1.615
+ $X2=3.33 $Y2=1.7
r79 8 10 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.245 $Y=1.615
+ $X2=3.245 $Y2=0.975
r80 5 25 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=4.285 $Y=1.47
+ $X2=4.25 $Y2=1.22
r81 5 7 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=4.285 $Y=1.47
+ $X2=4.285 $Y2=2.015
r82 1 20 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.04 $Y=0.84
+ $X2=3.04 $Y2=0.975
r83 1 3 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.04 $Y=0.84 $X2=3.04
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_4%A0 1 3 4 5 8 11 12 15 16
c50 1 0 1.20693e-19 $X=3.1 $Y=1.47
r51 15 18 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.755 $Y=0.98
+ $X2=3.755 $Y2=1.145
r52 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.755 $Y=0.98
+ $X2=3.755 $Y2=0.815
r53 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.755
+ $Y=0.98 $X2=3.755 $Y2=0.98
r54 12 16 7.44655 $w=3.23e-07 $l=2.1e-07 $layer=LI1_cond $X=3.832 $Y=1.19
+ $X2=3.832 $Y2=0.98
r55 11 18 58.026 $w=2e-07 $l=1.75e-07 $layer=POLY_cond $X=3.72 $Y=1.32 $X2=3.72
+ $Y2=1.145
r56 8 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.695 $Y=0.445
+ $X2=3.695 $Y2=0.815
r57 4 11 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=3.62 $Y=1.395
+ $X2=3.72 $Y2=1.32
r58 4 5 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.62 $Y=1.395 $X2=3.19
+ $Y2=1.395
r59 1 5 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.1 $Y=1.47
+ $X2=3.19 $Y2=1.395
r60 1 3 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=3.1 $Y=1.47 $X2=3.1
+ $Y2=2.015
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_4%A_925_21# 1 2 9 12 13 15 18 19 21 22 27
+ 32 33 34
c68 18 0 1.3232e-19 $X=4.79 $Y=1.02
c69 13 0 1.80039e-19 $X=4.725 $Y=1.47
c70 9 0 1.95128e-19 $X=4.7 $Y=0.445
r71 32 33 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=5.565 $Y=2
+ $X2=5.565 $Y2=1.835
r72 29 34 4.36305 $w=2.07e-07 $l=1.25499e-07 $layer=LI1_cond $X=5.68 $Y=0.865
+ $X2=5.59 $Y2=0.78
r73 29 33 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=5.68 $Y=0.865
+ $X2=5.68 $Y2=1.835
r74 25 34 4.36305 $w=2.07e-07 $l=1.08305e-07 $layer=LI1_cond $X=5.537 $Y=0.695
+ $X2=5.59 $Y2=0.78
r75 25 27 11.2892 $w=2.43e-07 $l=2.4e-07 $layer=LI1_cond $X=5.537 $Y=0.695
+ $X2=5.537 $Y2=0.455
r76 21 34 2.06925 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.415 $Y=0.78
+ $X2=5.59 $Y2=0.78
r77 21 22 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=5.415 $Y=0.78
+ $X2=4.875 $Y2=0.78
r78 19 37 39.6736 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.775 $Y=1.02
+ $X2=4.775 $Y2=1.185
r79 19 36 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.775 $Y=1.02
+ $X2=4.775 $Y2=0.855
r80 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.79
+ $Y=1.02 $X2=4.79 $Y2=1.02
r81 16 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.79 $Y=0.865
+ $X2=4.875 $Y2=0.78
r82 16 18 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.79 $Y=0.865
+ $X2=4.79 $Y2=1.02
r83 13 15 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=4.725 $Y=1.47
+ $X2=4.725 $Y2=2.015
r84 12 13 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.725 $Y=1.37 $X2=4.725
+ $Y2=1.47
r85 12 37 61.3418 $w=2e-07 $l=1.85e-07 $layer=POLY_cond $X=4.725 $Y=1.37
+ $X2=4.725 $Y2=1.185
r86 9 36 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=4.7 $Y=0.445 $X2=4.7
+ $Y2=0.855
r87 2 32 300 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=2 $X=5.385
+ $Y=1.545 $X2=5.53 $Y2=2
r88 1 27 182 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_NDIFF $count=1 $X=5.395
+ $Y=0.235 $X2=5.53 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_4%VPWR 1 2 3 4 13 15 21 25 29 35 38 39 40
+ 42 55 56 62 65
r66 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r67 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r68 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r69 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r70 53 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r71 52 53 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r72 50 53 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=4.83 $Y2=2.72
r73 50 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r74 49 52 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=4.83 $Y2=2.72
r75 49 50 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r76 47 65 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=2.28 $Y=2.72
+ $X2=2.142 $Y2=2.72
r77 47 49 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.28 $Y=2.72
+ $X2=2.53 $Y2=2.72
r78 46 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r79 46 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r80 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r81 43 59 4.06843 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r82 43 45 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.69 $Y2=2.72
r83 42 62 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=1.185 $Y2=2.72
r84 42 45 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=0.69 $Y2=2.72
r85 40 66 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=1.615 $Y=2.72
+ $X2=2.07 $Y2=2.72
r86 40 63 0.132312 $w=4.8e-07 $l=4.65e-07 $layer=MET1_cond $X=1.615 $Y=2.72
+ $X2=1.15 $Y2=2.72
r87 38 52 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.965 $Y=2.72
+ $X2=4.83 $Y2=2.72
r88 38 39 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.965 $Y=2.72
+ $X2=5.08 $Y2=2.72
r89 37 55 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=5.195 $Y=2.72
+ $X2=5.75 $Y2=2.72
r90 37 39 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.195 $Y=2.72
+ $X2=5.08 $Y2=2.72
r91 33 39 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.08 $Y=2.635
+ $X2=5.08 $Y2=2.72
r92 33 35 31.8174 $w=2.28e-07 $l=6.35e-07 $layer=LI1_cond $X=5.08 $Y=2.635
+ $X2=5.08 $Y2=2
r93 29 32 28.4968 $w=2.73e-07 $l=6.8e-07 $layer=LI1_cond $X=2.142 $Y=1.66
+ $X2=2.142 $Y2=2.34
r94 27 65 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.142 $Y=2.635
+ $X2=2.142 $Y2=2.72
r95 27 32 12.3626 $w=2.73e-07 $l=2.95e-07 $layer=LI1_cond $X=2.142 $Y=2.635
+ $X2=2.142 $Y2=2.34
r96 26 62 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.305 $Y=2.72
+ $X2=1.185 $Y2=2.72
r97 25 65 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=2.142 $Y2=2.72
r98 25 26 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=1.305 $Y2=2.72
r99 21 24 32.6526 $w=2.38e-07 $l=6.8e-07 $layer=LI1_cond $X=1.185 $Y=1.66
+ $X2=1.185 $Y2=2.34
r100 19 62 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.635
+ $X2=1.185 $Y2=2.72
r101 19 24 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=1.185 $Y=2.635
+ $X2=1.185 $Y2=2.34
r102 15 18 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=0.265 $Y=1.66
+ $X2=0.265 $Y2=2.34
r103 13 59 3.14379 $w=2.6e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.197 $Y2=2.72
r104 13 18 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.265 $Y2=2.34
r105 4 35 300 $w=1.7e-07 $l=5.60312e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=1.545 $X2=5.05 $Y2=2
r106 3 32 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2.34
r107 3 29 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.66
r108 2 24 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.34
r109 2 21 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.66
r110 1 18 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r111 1 15 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_4%X 1 2 3 4 15 17 21 25 29 30 32 35 36 37
+ 38 39
r48 39 52 4.1616 $w=3.58e-07 $l=1.3e-07 $layer=LI1_cond $X=1.655 $Y=2.21
+ $X2=1.655 $Y2=2.34
r49 38 39 10.8842 $w=3.58e-07 $l=3.4e-07 $layer=LI1_cond $X=1.655 $Y=1.87
+ $X2=1.655 $Y2=2.21
r50 35 36 6.02816 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.655 $Y=1.66
+ $X2=1.655 $Y2=1.495
r51 33 38 6.2424 $w=3.58e-07 $l=1.95e-07 $layer=LI1_cond $X=1.655 $Y=1.675
+ $X2=1.655 $Y2=1.87
r52 33 35 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=1.655 $Y=1.675
+ $X2=1.655 $Y2=1.66
r53 31 37 25.183 $w=2.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.61 $Y=1.065
+ $X2=1.61 $Y2=0.475
r54 31 32 5.00572 $w=2.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.61 $Y=1.065
+ $X2=1.61 $Y2=1.195
r55 27 32 5.00572 $w=2.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.61 $Y=1.325
+ $X2=1.61 $Y2=1.195
r56 27 36 7.25612 $w=2.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.61 $Y=1.325
+ $X2=1.61 $Y2=1.495
r57 26 30 1.34256 $w=2.6e-07 $l=1.3e-07 $layer=LI1_cond $X=0.85 $Y=1.195
+ $X2=0.72 $Y2=1.195
r58 25 32 1.47881 $w=2.6e-07 $l=1.35e-07 $layer=LI1_cond $X=1.475 $Y=1.195
+ $X2=1.61 $Y2=1.195
r59 25 26 27.703 $w=2.58e-07 $l=6.25e-07 $layer=LI1_cond $X=1.475 $Y=1.195
+ $X2=0.85 $Y2=1.195
r60 23 30 5.16603 $w=2.6e-07 $l=1.3e-07 $layer=LI1_cond $X=0.72 $Y=1.325
+ $X2=0.72 $Y2=1.195
r61 23 29 7.5352 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=0.72 $Y=1.325
+ $X2=0.72 $Y2=1.495
r62 19 30 5.16603 $w=2.6e-07 $l=1.3e-07 $layer=LI1_cond $X=0.72 $Y=1.065
+ $X2=0.72 $Y2=1.195
r63 19 21 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=0.72 $Y=1.065
+ $X2=0.72 $Y2=0.49
r64 15 29 6.08339 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=1.66
+ $X2=0.73 $Y2=1.495
r65 15 17 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.73 $Y=1.66
+ $X2=0.73 $Y2=2.34
r66 4 52 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
r67 4 35 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r68 3 17 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r69 3 15 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r70 2 37 182 $w=1.7e-07 $l=3e-07 $layer=licon1_NDIFF $count=1 $X=1.525 $Y=0.235
+ $X2=1.66 $Y2=0.475
r71 1 21 182 $w=1.7e-07 $l=3.15357e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.235 $X2=0.72 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_4%VGND 1 2 3 4 13 15 19 23 25 27 32 37 47
+ 48 54 57
c77 37 0 1.95128e-19 $X=4.63 $Y=0
r78 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r79 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r80 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r81 48 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=4.83
+ $Y2=0
r82 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r83 45 47 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=5.145 $Y=0 $X2=5.75
+ $Y2=0
r84 44 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r85 43 44 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r86 41 44 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.53 $Y=0 $X2=4.37
+ $Y2=0
r87 41 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r88 40 43 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=4.37
+ $Y2=0
r89 40 41 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r90 38 57 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.095
+ $Y2=0
r91 38 40 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.53
+ $Y2=0
r92 37 64 8.36094 $w=5.13e-07 $l=3.6e-07 $layer=LI1_cond $X=4.887 $Y=0 $X2=4.887
+ $Y2=0.36
r93 37 45 7.34265 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=4.887 $Y=0 $X2=5.145
+ $Y2=0
r94 37 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r95 37 43 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=4.63 $Y=0 $X2=4.37
+ $Y2=0
r96 33 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.18
+ $Y2=0
r97 33 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.61
+ $Y2=0
r98 32 57 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.915 $Y=0 $X2=2.095
+ $Y2=0
r99 32 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.915 $Y=0 $X2=1.61
+ $Y2=0
r100 31 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r101 31 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r102 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r103 28 51 3.9087 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=0.42 $Y=0 $X2=0.21
+ $Y2=0
r104 28 30 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.42 $Y=0 $X2=0.69
+ $Y2=0
r105 27 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.18
+ $Y2=0
r106 27 30 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.69 $Y2=0
r107 25 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r108 25 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r109 25 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r110 21 57 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=0.085
+ $X2=2.095 $Y2=0
r111 21 23 9.44363 $w=3.58e-07 $l=2.95e-07 $layer=LI1_cond $X=2.095 $Y=0.085
+ $X2=2.095 $Y2=0.38
r112 17 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0
r113 17 19 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0.49
r114 13 51 3.20141 $w=2.45e-07 $l=1.22327e-07 $layer=LI1_cond $X=0.297 $Y=0.085
+ $X2=0.21 $Y2=0
r115 13 15 19.0506 $w=2.43e-07 $l=4.05e-07 $layer=LI1_cond $X=0.297 $Y=0.085
+ $X2=0.297 $Y2=0.49
r116 4 64 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.235 $X2=5.01 $Y2=0.36
r117 3 23 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=1.945
+ $Y=0.235 $X2=2.11 $Y2=0.38
r118 2 19 182 $w=1.7e-07 $l=3.31134e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.235 $X2=1.18 $Y2=0.49
r119 1 15 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.235 $X2=0.3 $Y2=0.49
.ends

