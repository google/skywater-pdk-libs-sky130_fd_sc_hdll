* File: sky130_fd_sc_hdll__or4b_4.spice
* Created: Wed Sep  2 08:49:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or4b_4.pex.spice"
.subckt sky130_fd_sc_hdll__or4b_4  VNB VPB D_N C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1013 N_A_117_413#_M1013_d N_D_N_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15
+ W=0.42 AD=0.10785 AS=0.1302 PD=1.36 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 N_A_225_297#_M1014_d N_A_117_413#_M1014_g N_VGND_M1014_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.13975 AS=0.19785 PD=1.08 PS=1.92 NRD=13.836 NRS=8.304 M=1
+ R=4.33333 SA=75000.2 SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_C_M1012_g N_A_225_297#_M1014_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.13975 PD=0.97 PS=1.08 NRD=0 NRS=13.836 M=1 R=4.33333 SA=75000.8
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1007 N_A_225_297#_M1007_d N_B_M1007_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.3
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g N_A_225_297#_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.13975 AS=0.08775 PD=1.08 PS=0.92 NRD=26.76 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1002 N_X_M1002_d N_A_225_297#_M1002_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.13975 PD=0.97 PS=1.08 NRD=8.304 NRS=0.912 M=1 R=4.33333
+ SA=75002.3 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1010 N_X_M1002_d N_A_225_297#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1015 N_X_M1015_d N_A_225_297#_M1015_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1016 N_X_M1015_d N_A_225_297#_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.17875 PD=1.02 PS=1.85 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_A_117_413#_M1003_d N_D_N_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.1134 PD=1.38 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1017 A_315_297# N_A_117_413#_M1017_g N_A_225_297#_M1017_s VPB PHIGHVT L=0.18
+ W=1 AD=0.2 AS=0.27 PD=1.4 PS=2.54 NRD=28.5453 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.7 A=0.18 P=2.36 MULT=1
MM1008 A_431_297# N_C_M1008_g A_315_297# VPB PHIGHVT L=0.18 W=1 AD=0.145 AS=0.2
+ PD=1.29 PS=1.4 NRD=17.7103 NRS=28.5453 M=1 R=5.55556 SA=90000.8 SB=90003.1
+ A=0.18 P=2.36 MULT=1
MM1006 A_525_297# N_B_M1006_g A_431_297# VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=17.7103 NRS=17.7103 M=1 R=5.55556 SA=90001.2
+ SB=90002.6 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g A_525_297# VPB PHIGHVT L=0.18 W=1 AD=0.2
+ AS=0.145 PD=1.4 PS=1.29 NRD=11.8003 NRS=17.7103 M=1 R=5.55556 SA=90001.7
+ SB=90002.2 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1001_d N_A_225_297#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.2 AS=0.145 PD=1.4 PS=1.29 NRD=11.8003 NRS=0.9653 M=1 R=5.55556 SA=90002.3
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A_225_297#_M1004_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.7 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1004_d N_A_225_297#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_A_225_297#_M1011_g N_X_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.7 SB=90000.2 A=0.18 P=2.36 MULT=1
DX18_noxref VNB VPB NWDIODE A=9.4695 P=15.01
pX19_noxref noxref_15 A A PROBETYPE=1
*
.include "sky130_fd_sc_hdll__or4b_4.pxi.spice"
*
.ends
*
*
