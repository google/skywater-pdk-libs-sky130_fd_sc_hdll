* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__clkmux2_1 A0 A1 S VGND VNB VPB VPWR X
M1000 a_245_47# S VGND VNB nshort w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=4.76e+11p ps=4.08e+06u
M1001 a_478_47# A0 a_79_21# VNB nshort w=420000u l=150000u
+  ad=3.591e+11p pd=2.55e+06u as=2.121e+11p ps=1.85e+06u
M1002 a_79_21# A1 a_245_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=8.058e+11p pd=5.56e+06u as=2.7e+11p ps=2.54e+06u
M1004 a_599_309# A1 a_79_21# VPB phighvt w=940000u l=180000u
+  ad=2.444e+11p pd=2.4e+06u as=9.447e+11p ps=3.89e+06u
M1005 a_243_309# S VPWR VPB phighvt w=940000u l=180000u
+  ad=3.901e+11p pd=2.71e+06u as=0p ps=0u
M1006 a_649_21# S VPWR VPB phighvt w=940000u l=180000u
+  ad=2.726e+11p pd=2.46e+06u as=0p ps=0u
M1007 a_649_21# S VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1008 VGND a_649_21# a_478_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_79_21# A0 a_243_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_649_21# a_599_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_79_21# X VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
.ends
