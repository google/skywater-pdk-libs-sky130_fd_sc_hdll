* File: sky130_fd_sc_hdll__inv_1.pxi.spice
* Created: Wed Sep  2 08:32:57 2020
* 
x_PM_SKY130_FD_SC_HDLL__INV_1%A N_A_c_22_n N_A_M1001_g N_A_c_23_n N_A_M1000_g A
+ N_A_c_24_n A PM_SKY130_FD_SC_HDLL__INV_1%A
x_PM_SKY130_FD_SC_HDLL__INV_1%VPWR N_VPWR_M1001_s N_VPWR_c_43_n N_VPWR_c_44_n
+ N_VPWR_c_45_n VPWR N_VPWR_c_46_n N_VPWR_c_42_n
+ PM_SKY130_FD_SC_HDLL__INV_1%VPWR
x_PM_SKY130_FD_SC_HDLL__INV_1%Y N_Y_M1000_d N_Y_M1001_d N_Y_c_58_n N_Y_c_56_n Y
+ Y Y PM_SKY130_FD_SC_HDLL__INV_1%Y
x_PM_SKY130_FD_SC_HDLL__INV_1%VGND N_VGND_M1000_s N_VGND_c_75_n N_VGND_c_76_n
+ N_VGND_c_77_n VGND N_VGND_c_78_n N_VGND_c_79_n
+ PM_SKY130_FD_SC_HDLL__INV_1%VGND
cc_1 VNB N_A_c_22_n 0.0451735f $X=-0.19 $Y=-0.24 $X2=0.7 $Y2=1.41
cc_2 VNB N_A_c_23_n 0.0259537f $X=-0.19 $Y=-0.24 $X2=0.725 $Y2=0.995
cc_3 VNB N_A_c_24_n 0.0175443f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.16
cc_4 VNB N_VPWR_c_42_n 0.0609879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_Y_c_56_n 0.0335947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB Y 0.0232935f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.195
cc_7 VNB N_VGND_c_75_n 0.0309566f $X=-0.19 $Y=-0.24 $X2=0.725 $Y2=0.56
cc_8 VNB N_VGND_c_76_n 0.0123263f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=1.16
cc_9 VNB N_VGND_c_77_n 0.00442399f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.16
cc_10 VNB N_VGND_c_78_n 0.0236003f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_VGND_c_79_n 0.115195f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VPB N_A_c_22_n 0.0450154f $X=-0.19 $Y=1.305 $X2=0.7 $Y2=1.41
cc_13 VPB N_A_c_24_n 0.00843691f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.16
cc_14 VPB N_VPWR_c_43_n 0.00496839f $X=-0.19 $Y=1.305 $X2=0.725 $Y2=0.56
cc_15 VPB N_VPWR_c_44_n 0.0129628f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.16
cc_16 VPB N_VPWR_c_45_n 0.00401341f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.195
cc_17 VPB N_VPWR_c_46_n 0.0236036f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_18 VPB N_VPWR_c_42_n 0.0550088f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_19 VPB N_Y_c_58_n 0.0360264f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.16
cc_20 VPB Y 0.0100058f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.195
cc_21 VPB Y 0.0143357f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_22 N_A_c_22_n N_VPWR_c_43_n 0.0131923f $X=0.7 $Y=1.41 $X2=0 $Y2=0
cc_23 N_A_c_24_n N_VPWR_c_43_n 0.0160759f $X=0.485 $Y=1.16 $X2=0 $Y2=0
cc_24 N_A_c_22_n N_VPWR_c_46_n 0.00673617f $X=0.7 $Y=1.41 $X2=0 $Y2=0
cc_25 N_A_c_22_n N_VPWR_c_42_n 0.0139414f $X=0.7 $Y=1.41 $X2=0 $Y2=0
cc_26 N_A_c_22_n N_Y_c_58_n 0.00906448f $X=0.7 $Y=1.41 $X2=0 $Y2=0
cc_27 N_A_c_23_n N_Y_c_56_n 0.00871655f $X=0.725 $Y=0.995 $X2=0 $Y2=0
cc_28 N_A_c_22_n Y 8.79174e-19 $X=0.7 $Y=1.41 $X2=0 $Y2=0
cc_29 N_A_c_23_n Y 0.0151236f $X=0.725 $Y=0.995 $X2=0 $Y2=0
cc_30 N_A_c_24_n Y 0.0114518f $X=0.485 $Y=1.16 $X2=0 $Y2=0
cc_31 N_A_c_22_n Y 0.00398335f $X=0.7 $Y=1.41 $X2=0 $Y2=0
cc_32 N_A_c_22_n N_VGND_c_75_n 0.00585411f $X=0.7 $Y=1.41 $X2=0 $Y2=0
cc_33 N_A_c_23_n N_VGND_c_75_n 0.00736901f $X=0.725 $Y=0.995 $X2=0 $Y2=0
cc_34 N_A_c_24_n N_VGND_c_75_n 0.0188164f $X=0.485 $Y=1.16 $X2=0 $Y2=0
cc_35 N_A_c_23_n N_VGND_c_78_n 0.00541359f $X=0.725 $Y=0.995 $X2=0 $Y2=0
cc_36 N_A_c_23_n N_VGND_c_79_n 0.0118398f $X=0.725 $Y=0.995 $X2=0 $Y2=0
cc_37 N_VPWR_c_42_n N_Y_M1001_d 0.00217517f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_38 N_VPWR_c_46_n N_Y_c_58_n 0.0343232f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_39 N_VPWR_c_42_n N_Y_c_58_n 0.0195972f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_40 N_VPWR_c_43_n Y 0.0617158f $X=0.465 $Y=1.66 $X2=0 $Y2=0
cc_41 N_Y_c_56_n N_VGND_c_75_n 0.0403728f $X=0.935 $Y=0.4 $X2=0 $Y2=0
cc_42 N_Y_c_56_n N_VGND_c_78_n 0.034237f $X=0.935 $Y=0.4 $X2=0 $Y2=0
cc_43 N_Y_M1000_d N_VGND_c_79_n 0.00209319f $X=0.8 $Y=0.235 $X2=0 $Y2=0
cc_44 N_Y_c_56_n N_VGND_c_79_n 0.0195344f $X=0.935 $Y=0.4 $X2=0 $Y2=0
