* File: sky130_fd_sc_hdll__a32o_1.spice
* Created: Thu Aug 27 18:56:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a32o_1.pex.spice"
.subckt sky130_fd_sc_hdll__a32o_1  VNB VPB A3 A2 A1 B1 B2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_93_21#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.199875 AS=0.2145 PD=1.265 PS=1.96 NRD=10.152 NRS=11.988 M=1 R=4.33333
+ SA=75000.3 SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1000 A_276_47# N_A3_M1000_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65 AD=0.0975
+ AS=0.199875 PD=0.95 PS=1.265 NRD=17.532 NRS=51.684 M=1 R=4.33333 SA=75001
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1004 A_366_47# N_A2_M1004_g A_276_47# VNB NSHORT L=0.15 W=0.65 AD=0.17875
+ AS=0.0975 PD=1.2 PS=0.95 NRD=40.608 NRS=17.532 M=1 R=4.33333 SA=75001.5
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1003 N_A_93_21#_M1003_d N_A1_M1003_g A_366_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.15925 AS=0.17875 PD=1.14 PS=1.2 NRD=13.836 NRS=40.608 M=1 R=4.33333
+ SA=75002.2 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1006 A_634_47# N_B1_M1006_g N_A_93_21#_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.15925 PD=0.86 PS=1.14 NRD=9.228 NRS=24.912 M=1 R=4.33333
+ SA=75002.8 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_B2_M1011_g A_634_47# VNB NSHORT L=0.15 W=0.65 AD=0.20475
+ AS=0.06825 PD=1.93 PS=0.86 NRD=9.228 NRS=9.228 M=1 R=4.33333 SA=75003.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_A_93_21#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.2525 AS=0.34 PD=1.505 PS=2.68 NRD=18.715 NRS=14.775 M=1 R=5.55556
+ SA=90000.2 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1009 N_A_268_297#_M1009_d N_A3_M1009_g N_VPWR_M1001_d VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.2525 PD=1.35 PS=1.505 NRD=6.8753 NRS=25.5903 M=1 R=5.55556
+ SA=90000.9 SB=90002.4 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_A2_M1007_g N_A_268_297#_M1009_d VPB PHIGHVT L=0.18 W=1
+ AD=0.235 AS=0.175 PD=1.47 PS=1.35 NRD=18.715 NRS=6.8753 M=1 R=5.55556
+ SA=90001.5 SB=90001.9 A=0.18 P=2.36 MULT=1
MM1008 N_A_268_297#_M1008_d N_A1_M1008_g N_VPWR_M1007_d VPB PHIGHVT L=0.18 W=1
+ AD=0.195 AS=0.235 PD=1.39 PS=1.47 NRD=9.8303 NRS=18.715 M=1 R=5.55556
+ SA=90002.1 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1002 N_A_93_21#_M1002_d N_B1_M1002_g N_A_268_297#_M1008_d VPB PHIGHVT L=0.18
+ W=1 AD=0.15 AS=0.195 PD=1.3 PS=1.39 NRD=1.9503 NRS=11.8003 M=1 R=5.55556
+ SA=90002.7 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1010 N_A_268_297#_M1010_d N_B2_M1010_g N_A_93_21#_M1002_d VPB PHIGHVT L=0.18
+ W=1 AD=0.275 AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556
+ SA=90003.2 SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hdll__a32o_1.pxi.spice"
*
.ends
*
*
