* File: sky130_fd_sc_hdll__and4bb_4.pxi.spice
* Created: Wed Sep  2 08:23:48 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND4BB_4%B_N N_B_N_c_101_n N_B_N_c_102_n N_B_N_M1002_g
+ N_B_N_M1014_g B_N B_N B_N N_B_N_c_100_n PM_SKY130_FD_SC_HDLL__AND4BB_4%B_N
x_PM_SKY130_FD_SC_HDLL__AND4BB_4%A_184_21# N_A_184_21#_M1003_d
+ N_A_184_21#_M1011_d N_A_184_21#_M1004_d N_A_184_21#_M1005_g
+ N_A_184_21#_c_147_n N_A_184_21#_M1008_g N_A_184_21#_M1007_g
+ N_A_184_21#_c_148_n N_A_184_21#_M1010_g N_A_184_21#_M1015_g
+ N_A_184_21#_c_149_n N_A_184_21#_M1013_g N_A_184_21#_M1016_g
+ N_A_184_21#_c_150_n N_A_184_21#_M1019_g N_A_184_21#_c_141_n
+ N_A_184_21#_c_142_n N_A_184_21#_c_143_n N_A_184_21#_c_162_p
+ N_A_184_21#_c_248_p N_A_184_21#_c_196_p N_A_184_21#_c_168_p
+ N_A_184_21#_c_163_p N_A_184_21#_c_169_p N_A_184_21#_c_164_p
+ N_A_184_21#_c_144_n N_A_184_21#_c_145_n N_A_184_21#_c_146_n
+ PM_SKY130_FD_SC_HDLL__AND4BB_4%A_184_21#
x_PM_SKY130_FD_SC_HDLL__AND4BB_4%D N_D_c_286_n N_D_M1000_g N_D_c_287_n
+ N_D_M1011_g D PM_SKY130_FD_SC_HDLL__AND4BB_4%D
x_PM_SKY130_FD_SC_HDLL__AND4BB_4%C N_C_c_321_n N_C_M1017_g N_C_c_322_n
+ N_C_M1006_g C C C PM_SKY130_FD_SC_HDLL__AND4BB_4%C
x_PM_SKY130_FD_SC_HDLL__AND4BB_4%A_27_47# N_A_27_47#_M1014_s N_A_27_47#_M1002_s
+ N_A_27_47#_c_354_n N_A_27_47#_M1009_g N_A_27_47#_c_355_n N_A_27_47#_M1004_g
+ N_A_27_47#_c_356_n N_A_27_47#_c_362_n N_A_27_47#_c_363_n N_A_27_47#_c_357_n
+ N_A_27_47#_c_365_n N_A_27_47#_c_358_n N_A_27_47#_c_366_n N_A_27_47#_c_359_n
+ PM_SKY130_FD_SC_HDLL__AND4BB_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__AND4BB_4%A_912_21# N_A_912_21#_M1012_d
+ N_A_912_21#_M1001_d N_A_912_21#_M1003_g N_A_912_21#_c_452_n
+ N_A_912_21#_M1018_g N_A_912_21#_c_447_n N_A_912_21#_c_448_n
+ N_A_912_21#_c_449_n N_A_912_21#_c_450_n N_A_912_21#_c_451_n
+ N_A_912_21#_c_456_n N_A_912_21#_c_457_n N_A_912_21#_c_476_p
+ N_A_912_21#_c_479_p PM_SKY130_FD_SC_HDLL__AND4BB_4%A_912_21#
x_PM_SKY130_FD_SC_HDLL__AND4BB_4%A_N N_A_N_M1012_g N_A_N_c_519_n N_A_N_c_520_n
+ N_A_N_M1001_g A_N A_N N_A_N_c_518_n PM_SKY130_FD_SC_HDLL__AND4BB_4%A_N
x_PM_SKY130_FD_SC_HDLL__AND4BB_4%VPWR N_VPWR_M1002_d N_VPWR_M1010_d
+ N_VPWR_M1019_d N_VPWR_M1006_d N_VPWR_M1018_d N_VPWR_c_544_n N_VPWR_c_545_n
+ N_VPWR_c_546_n N_VPWR_c_547_n VPWR N_VPWR_c_548_n N_VPWR_c_549_n
+ N_VPWR_c_550_n N_VPWR_c_551_n N_VPWR_c_552_n N_VPWR_c_543_n N_VPWR_c_554_n
+ N_VPWR_c_555_n N_VPWR_c_556_n N_VPWR_c_557_n N_VPWR_c_558_n
+ PM_SKY130_FD_SC_HDLL__AND4BB_4%VPWR
x_PM_SKY130_FD_SC_HDLL__AND4BB_4%X N_X_M1005_s N_X_M1015_s N_X_M1008_s
+ N_X_M1013_s N_X_c_641_n N_X_c_642_n N_X_c_646_n N_X_c_651_n X X X N_X_c_637_n
+ X X PM_SKY130_FD_SC_HDLL__AND4BB_4%X
x_PM_SKY130_FD_SC_HDLL__AND4BB_4%VGND N_VGND_M1014_d N_VGND_M1007_d
+ N_VGND_M1016_d N_VGND_M1012_s N_VGND_c_682_n N_VGND_c_683_n N_VGND_c_684_n
+ N_VGND_c_685_n N_VGND_c_686_n N_VGND_c_687_n N_VGND_c_688_n VGND
+ N_VGND_c_689_n N_VGND_c_690_n N_VGND_c_691_n N_VGND_c_692_n N_VGND_c_693_n
+ N_VGND_c_694_n VGND PM_SKY130_FD_SC_HDLL__AND4BB_4%VGND
cc_1 VNB N_B_N_M1014_g 0.0337551f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB B_N 0.00596462f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=0.765
cc_3 VNB N_B_N_c_100_n 0.0272715f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_4 VNB N_A_184_21#_M1005_g 0.0178615f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.445
cc_5 VNB N_A_184_21#_M1007_g 0.0183071f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_6 VNB N_A_184_21#_M1015_g 0.0183515f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_184_21#_M1016_g 0.0193318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_184_21#_c_141_n 0.00132792f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_184_21#_c_142_n 0.00362687f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_184_21#_c_143_n 9.97074e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_184_21#_c_144_n 0.00136342f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_184_21#_c_145_n 0.0123871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_184_21#_c_146_n 0.0687494f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_D_c_286_n 0.0187399f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_15 VNB N_D_c_287_n 0.0300175f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_16 VNB D 0.00163636f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_17 VNB N_C_c_321_n 0.0177525f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_18 VNB N_C_c_322_n 0.0250738f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_19 VNB C 0.00644538f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_20 VNB N_A_27_47#_c_354_n 0.0187555f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_21 VNB N_A_27_47#_c_355_n 0.0251891f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=0.765
cc_22 VNB N_A_27_47#_c_356_n 0.0332169f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_357_n 0.00721425f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=0.85
cc_24 VNB N_A_27_47#_c_358_n 0.0128993f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_359_n 0.00179704f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_912_21#_M1003_g 0.0233479f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_912_21#_c_447_n 0.0113258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_912_21#_c_448_n 0.0051116f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_29 VNB N_A_912_21#_c_449_n 0.0608773f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.325
cc_30 VNB N_A_912_21#_c_450_n 0.023054f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=0.85
cc_31 VNB N_A_912_21#_c_451_n 0.00315239f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_N_M1012_g 0.0431418f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.99
cc_33 VNB A_N 0.0175776f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=0.765
cc_34 VNB N_A_N_c_518_n 0.0322479f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VPWR_c_543_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB X 0.00136782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_682_n 0.00271958f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_38 VNB N_VGND_c_683_n 3.22956e-19 $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=0.85
cc_39 VNB N_VGND_c_684_n 0.0137618f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_685_n 0.00283014f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.53
cc_41 VNB N_VGND_c_686_n 0.00564356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_687_n 0.0633558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_688_n 0.00631443f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_689_n 0.0126369f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_690_n 0.0220027f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_691_n 0.328789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_692_n 0.0245177f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_693_n 0.00502664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_694_n 0.00518879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VPB N_B_N_c_101_n 0.0348063f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_51 VPB N_B_N_c_102_n 0.0263351f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_52 VPB B_N 0.00193771f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=0.765
cc_53 VPB N_B_N_c_100_n 0.00485173f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_54 VPB N_A_184_21#_c_147_n 0.0164656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_184_21#_c_148_n 0.0157879f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=0.85
cc_56 VPB N_A_184_21#_c_149_n 0.016086f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_184_21#_c_150_n 0.0164917f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_184_21#_c_143_n 0.00382282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_184_21#_c_146_n 0.045789f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_D_c_287_n 0.0297536f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_61 VPB D 0.0011597f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_62 VPB N_C_c_322_n 0.0304949f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_63 VPB C 0.00307174f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_64 VPB N_A_27_47#_c_355_n 0.0282712f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=0.765
cc_65 VPB N_A_27_47#_c_356_n 0.0290594f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_27_47#_c_362_n 0.0147617f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_67 VPB N_A_27_47#_c_363_n 0.00204048f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_68 VPB N_A_27_47#_c_357_n 0.00252093f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=0.85
cc_69 VPB N_A_27_47#_c_365_n 0.00242581f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.16
cc_70 VPB N_A_27_47#_c_366_n 0.0110158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_47#_c_359_n 7.40731e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_912_21#_c_452_n 0.0197653f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_73 VPB N_A_912_21#_c_447_n 0.00532644f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_912_21#_c_448_n 0.0132433f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_75 VPB N_A_912_21#_c_449_n 0.0423328f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.325
cc_76 VPB N_A_912_21#_c_456_n 0.0179016f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_912_21#_c_457_n 0.00255295f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.16
cc_78 VPB N_A_N_c_519_n 0.0472542f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_79 VPB N_A_N_c_520_n 0.0317967f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_80 VPB A_N 0.0182963f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=0.765
cc_81 VPB N_A_N_c_518_n 0.00624817f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_544_n 0.0132269f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.16
cc_83 VPB N_VPWR_c_545_n 0.00561645f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.325
cc_84 VPB N_VPWR_c_546_n 0.0113234f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.19
cc_85 VPB N_VPWR_c_547_n 0.00872728f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_548_n 0.0143107f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_549_n 0.0157854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_550_n 0.0232448f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_551_n 0.00874105f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_552_n 0.0190623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_543_n 0.0456593f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_554_n 0.00810608f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_555_n 0.00538861f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_556_n 0.00862719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_557_n 0.00631443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_558_n 0.0218481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB X 0.00108433f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 N_B_N_M1014_g N_A_184_21#_M1005_g 0.019485f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_99 B_N N_A_184_21#_M1005_g 0.00509309f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_100 N_B_N_c_100_n N_A_184_21#_M1005_g 0.0201607f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_101 N_B_N_c_101_n N_A_184_21#_c_147_n 0.0208356f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_102 N_B_N_c_102_n N_A_184_21#_c_147_n 0.015366f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_103 B_N N_A_184_21#_c_147_n 0.00177729f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_104 N_B_N_c_101_n N_A_184_21#_c_146_n 0.00297917f $X=0.495 $Y=1.89 $X2=0
+ $Y2=0
cc_105 N_B_N_c_101_n N_A_27_47#_c_356_n 0.0168126f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_106 N_B_N_M1014_g N_A_27_47#_c_356_n 0.00714298f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_107 B_N N_A_27_47#_c_356_n 0.0674358f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_108 N_B_N_c_100_n N_A_27_47#_c_356_n 0.00780387f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_109 N_B_N_c_102_n N_A_27_47#_c_362_n 0.00467732f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_110 N_B_N_c_102_n N_A_27_47#_c_363_n 0.0169508f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_111 B_N N_A_27_47#_c_363_n 0.0217857f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_112 N_B_N_c_100_n N_A_27_47#_c_363_n 7.40595e-19 $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_113 B_N N_VPWR_M1002_d 0.00388739f $X=0.66 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_114 N_B_N_c_102_n N_VPWR_c_548_n 0.00315013f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_115 N_B_N_c_102_n N_VPWR_c_543_n 0.0046225f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_116 N_B_N_c_102_n N_VPWR_c_554_n 0.0109875f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_117 N_B_N_M1014_g X 6.24427e-19 $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_118 B_N X 0.0043968f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_119 N_B_N_c_101_n N_X_c_637_n 4.9522e-19 $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_120 B_N N_X_c_637_n 0.00719478f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_121 B_N X 0.0554706f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_122 N_B_N_c_100_n X 2.83674e-19 $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_123 B_N N_VGND_M1014_d 0.00337877f $X=0.66 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_124 N_B_N_M1014_g N_VGND_c_682_n 0.00310635f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_125 B_N N_VGND_c_682_n 0.0101817f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_126 N_B_N_c_100_n N_VGND_c_682_n 2.92234e-19 $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_127 N_B_N_M1014_g N_VGND_c_691_n 0.00707553f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_128 B_N N_VGND_c_691_n 0.00780194f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_129 N_B_N_M1014_g N_VGND_c_692_n 0.00585385f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_130 N_A_184_21#_M1016_g N_D_c_286_n 0.0127239f $X=2.405 $Y=0.56 $X2=-0.19
+ $Y2=-0.24
cc_131 N_A_184_21#_c_142_n N_D_c_286_n 0.00302527f $X=2.615 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_132 N_A_184_21#_c_162_p N_D_c_286_n 0.0115936f $X=2.975 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_133 N_A_184_21#_c_163_p N_D_c_286_n 0.00458463f $X=3.085 $Y=0.615 $X2=-0.19
+ $Y2=-0.24
cc_134 N_A_184_21#_c_164_p N_D_c_286_n 0.0056695f $X=3.195 $Y=0.385 $X2=-0.19
+ $Y2=-0.24
cc_135 N_A_184_21#_c_150_n N_D_c_287_n 0.0331972f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A_184_21#_c_143_n N_D_c_287_n 0.00529983f $X=2.615 $Y=1.545 $X2=0 $Y2=0
cc_137 N_A_184_21#_c_162_p N_D_c_287_n 0.00103495f $X=2.975 $Y=0.7 $X2=0 $Y2=0
cc_138 N_A_184_21#_c_168_p N_D_c_287_n 0.0156375f $X=4.385 $Y=1.63 $X2=0 $Y2=0
cc_139 N_A_184_21#_c_169_p N_D_c_287_n 0.00102461f $X=4.71 $Y=0.385 $X2=0 $Y2=0
cc_140 N_A_184_21#_c_144_n N_D_c_287_n 0.00153128f $X=2.615 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A_184_21#_c_146_n N_D_c_287_n 0.0159255f $X=2.405 $Y=1.217 $X2=0 $Y2=0
cc_142 N_A_184_21#_c_142_n D 0.00514029f $X=2.615 $Y=1.075 $X2=0 $Y2=0
cc_143 N_A_184_21#_c_143_n D 0.00514029f $X=2.615 $Y=1.545 $X2=0 $Y2=0
cc_144 N_A_184_21#_c_162_p D 0.0169298f $X=2.975 $Y=0.7 $X2=0 $Y2=0
cc_145 N_A_184_21#_c_168_p D 0.0153904f $X=4.385 $Y=1.63 $X2=0 $Y2=0
cc_146 N_A_184_21#_c_144_n D 0.0123502f $X=2.615 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_184_21#_c_162_p N_C_c_321_n 0.00116634f $X=2.975 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_148 N_A_184_21#_c_163_p N_C_c_321_n 0.00300221f $X=3.085 $Y=0.615 $X2=-0.19
+ $Y2=-0.24
cc_149 N_A_184_21#_c_169_p N_C_c_321_n 0.0113637f $X=4.71 $Y=0.385 $X2=-0.19
+ $Y2=-0.24
cc_150 N_A_184_21#_c_168_p N_C_c_322_n 0.0119485f $X=4.385 $Y=1.63 $X2=0 $Y2=0
cc_151 N_A_184_21#_c_169_p N_C_c_322_n 6.80209e-19 $X=4.71 $Y=0.385 $X2=0 $Y2=0
cc_152 N_A_184_21#_c_142_n C 0.00621169f $X=2.615 $Y=1.075 $X2=0 $Y2=0
cc_153 N_A_184_21#_c_162_p C 0.012653f $X=2.975 $Y=0.7 $X2=0 $Y2=0
cc_154 N_A_184_21#_c_168_p C 0.0270167f $X=4.385 $Y=1.63 $X2=0 $Y2=0
cc_155 N_A_184_21#_c_169_p C 0.0268867f $X=4.71 $Y=0.385 $X2=0 $Y2=0
cc_156 N_A_184_21#_c_169_p N_A_27_47#_c_354_n 0.0139343f $X=4.71 $Y=0.385 $X2=0
+ $Y2=0
cc_157 N_A_184_21#_c_168_p N_A_27_47#_c_355_n 0.0124336f $X=4.385 $Y=1.63 $X2=0
+ $Y2=0
cc_158 N_A_184_21#_c_169_p N_A_27_47#_c_355_n 0.00177565f $X=4.71 $Y=0.385 $X2=0
+ $Y2=0
cc_159 N_A_184_21#_M1011_d N_A_27_47#_c_363_n 0.00794166f $X=3.07 $Y=1.485 $X2=0
+ $Y2=0
cc_160 N_A_184_21#_M1004_d N_A_27_47#_c_363_n 0.00672518f $X=4.22 $Y=1.485 $X2=0
+ $Y2=0
cc_161 N_A_184_21#_c_147_n N_A_27_47#_c_363_n 0.016342f $X=1.02 $Y=1.41 $X2=0
+ $Y2=0
cc_162 N_A_184_21#_c_148_n N_A_27_47#_c_363_n 0.0131122f $X=1.49 $Y=1.41 $X2=0
+ $Y2=0
cc_163 N_A_184_21#_c_149_n N_A_27_47#_c_363_n 0.0135818f $X=1.96 $Y=1.41 $X2=0
+ $Y2=0
cc_164 N_A_184_21#_c_150_n N_A_27_47#_c_363_n 0.0156415f $X=2.43 $Y=1.41 $X2=0
+ $Y2=0
cc_165 N_A_184_21#_c_141_n N_A_27_47#_c_363_n 0.00371062f $X=2.53 $Y=1.16 $X2=0
+ $Y2=0
cc_166 N_A_184_21#_c_196_p N_A_27_47#_c_363_n 0.00882574f $X=2.7 $Y=1.63 $X2=0
+ $Y2=0
cc_167 N_A_184_21#_c_168_p N_A_27_47#_c_363_n 0.0919942f $X=4.385 $Y=1.63 $X2=0
+ $Y2=0
cc_168 N_A_184_21#_c_146_n N_A_27_47#_c_363_n 7.06015e-19 $X=2.405 $Y=1.217
+ $X2=0 $Y2=0
cc_169 N_A_184_21#_c_168_p N_A_27_47#_c_357_n 0.017148f $X=4.385 $Y=1.63 $X2=0
+ $Y2=0
cc_170 N_A_184_21#_c_145_n N_A_27_47#_c_357_n 0.0086059f $X=4.895 $Y=0.385 $X2=0
+ $Y2=0
cc_171 N_A_184_21#_c_168_p N_A_27_47#_c_359_n 0.0141955f $X=4.385 $Y=1.63 $X2=0
+ $Y2=0
cc_172 N_A_184_21#_c_169_p N_A_27_47#_c_359_n 0.00564306f $X=4.71 $Y=0.385 $X2=0
+ $Y2=0
cc_173 N_A_184_21#_c_169_p N_A_912_21#_M1003_g 0.0130123f $X=4.71 $Y=0.385 $X2=0
+ $Y2=0
cc_174 N_A_184_21#_c_145_n N_A_912_21#_c_447_n 0.0104098f $X=4.895 $Y=0.385
+ $X2=0 $Y2=0
cc_175 N_A_184_21#_c_145_n N_A_912_21#_c_451_n 0.00926983f $X=4.895 $Y=0.385
+ $X2=0 $Y2=0
cc_176 N_A_184_21#_c_143_n N_VPWR_M1019_d 0.00109221f $X=2.615 $Y=1.545 $X2=0
+ $Y2=0
cc_177 N_A_184_21#_c_196_p N_VPWR_M1019_d 0.00260913f $X=2.7 $Y=1.63 $X2=0 $Y2=0
cc_178 N_A_184_21#_c_168_p N_VPWR_M1019_d 0.00658236f $X=4.385 $Y=1.63 $X2=0
+ $Y2=0
cc_179 N_A_184_21#_c_168_p N_VPWR_M1006_d 0.0106675f $X=4.385 $Y=1.63 $X2=0
+ $Y2=0
cc_180 N_A_184_21#_c_149_n N_VPWR_c_544_n 0.00453434f $X=1.96 $Y=1.41 $X2=0
+ $Y2=0
cc_181 N_A_184_21#_c_150_n N_VPWR_c_544_n 0.00311736f $X=2.43 $Y=1.41 $X2=0
+ $Y2=0
cc_182 N_A_184_21#_c_147_n N_VPWR_c_549_n 0.00510113f $X=1.02 $Y=1.41 $X2=0
+ $Y2=0
cc_183 N_A_184_21#_c_148_n N_VPWR_c_549_n 0.00311736f $X=1.49 $Y=1.41 $X2=0
+ $Y2=0
cc_184 N_A_184_21#_M1011_d N_VPWR_c_543_n 0.00449607f $X=3.07 $Y=1.485 $X2=0
+ $Y2=0
cc_185 N_A_184_21#_M1004_d N_VPWR_c_543_n 0.00408734f $X=4.22 $Y=1.485 $X2=0
+ $Y2=0
cc_186 N_A_184_21#_c_147_n N_VPWR_c_543_n 0.00683693f $X=1.02 $Y=1.41 $X2=0
+ $Y2=0
cc_187 N_A_184_21#_c_148_n N_VPWR_c_543_n 0.00375605f $X=1.49 $Y=1.41 $X2=0
+ $Y2=0
cc_188 N_A_184_21#_c_149_n N_VPWR_c_543_n 0.00518254f $X=1.96 $Y=1.41 $X2=0
+ $Y2=0
cc_189 N_A_184_21#_c_150_n N_VPWR_c_543_n 0.00375605f $X=2.43 $Y=1.41 $X2=0
+ $Y2=0
cc_190 N_A_184_21#_c_147_n N_VPWR_c_554_n 0.00294646f $X=1.02 $Y=1.41 $X2=0
+ $Y2=0
cc_191 N_A_184_21#_c_147_n N_VPWR_c_555_n 0.00122179f $X=1.02 $Y=1.41 $X2=0
+ $Y2=0
cc_192 N_A_184_21#_c_148_n N_VPWR_c_555_n 0.0113834f $X=1.49 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A_184_21#_c_149_n N_VPWR_c_555_n 0.00820729f $X=1.96 $Y=1.41 $X2=0
+ $Y2=0
cc_194 N_A_184_21#_c_150_n N_VPWR_c_555_n 0.00106505f $X=2.43 $Y=1.41 $X2=0
+ $Y2=0
cc_195 N_A_184_21#_c_149_n N_VPWR_c_556_n 0.00118604f $X=1.96 $Y=1.41 $X2=0
+ $Y2=0
cc_196 N_A_184_21#_c_150_n N_VPWR_c_556_n 0.0111044f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A_184_21#_M1005_g N_X_c_641_n 0.00418768f $X=0.995 $Y=0.56 $X2=0 $Y2=0
cc_198 N_A_184_21#_M1007_g N_X_c_642_n 0.0158372f $X=1.465 $Y=0.56 $X2=0 $Y2=0
cc_199 N_A_184_21#_M1015_g N_X_c_642_n 0.0121812f $X=1.935 $Y=0.56 $X2=0 $Y2=0
cc_200 N_A_184_21#_c_141_n N_X_c_642_n 0.035252f $X=2.53 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A_184_21#_c_146_n N_X_c_642_n 0.00647965f $X=2.405 $Y=1.217 $X2=0 $Y2=0
cc_202 N_A_184_21#_c_148_n N_X_c_646_n 0.0136903f $X=1.49 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A_184_21#_c_149_n N_X_c_646_n 0.0108985f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A_184_21#_c_150_n N_X_c_646_n 0.00242896f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A_184_21#_c_141_n N_X_c_646_n 0.0324737f $X=2.53 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A_184_21#_c_146_n N_X_c_646_n 0.0133137f $X=2.405 $Y=1.217 $X2=0 $Y2=0
cc_207 N_A_184_21#_M1015_g N_X_c_651_n 0.00418768f $X=1.935 $Y=0.56 $X2=0 $Y2=0
cc_208 N_A_184_21#_M1005_g X 0.00703379f $X=0.995 $Y=0.56 $X2=0 $Y2=0
cc_209 N_A_184_21#_c_147_n N_X_c_637_n 0.0051553f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A_184_21#_M1005_g X 0.00479821f $X=0.995 $Y=0.56 $X2=0 $Y2=0
cc_211 N_A_184_21#_c_147_n X 0.00285709f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A_184_21#_M1007_g X 0.00417507f $X=1.465 $Y=0.56 $X2=0 $Y2=0
cc_213 N_A_184_21#_c_148_n X 0.00338287f $X=1.49 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A_184_21#_c_141_n X 0.0134106f $X=2.53 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A_184_21#_c_146_n X 0.0344015f $X=2.405 $Y=1.217 $X2=0 $Y2=0
cc_216 N_A_184_21#_c_142_n N_VGND_M1016_d 0.00235205f $X=2.615 $Y=1.075 $X2=0
+ $Y2=0
cc_217 N_A_184_21#_c_162_p N_VGND_M1016_d 0.00604511f $X=2.975 $Y=0.7 $X2=0
+ $Y2=0
cc_218 N_A_184_21#_c_248_p N_VGND_M1016_d 0.00319468f $X=2.7 $Y=0.7 $X2=0 $Y2=0
cc_219 N_A_184_21#_M1005_g N_VGND_c_682_n 0.00808243f $X=0.995 $Y=0.56 $X2=0
+ $Y2=0
cc_220 N_A_184_21#_M1007_g N_VGND_c_682_n 5.11974e-19 $X=1.465 $Y=0.56 $X2=0
+ $Y2=0
cc_221 N_A_184_21#_M1005_g N_VGND_c_683_n 4.99752e-19 $X=0.995 $Y=0.56 $X2=0
+ $Y2=0
cc_222 N_A_184_21#_M1007_g N_VGND_c_683_n 0.00707579f $X=1.465 $Y=0.56 $X2=0
+ $Y2=0
cc_223 N_A_184_21#_M1015_g N_VGND_c_683_n 0.00737164f $X=1.935 $Y=0.56 $X2=0
+ $Y2=0
cc_224 N_A_184_21#_M1016_g N_VGND_c_683_n 5.22065e-19 $X=2.405 $Y=0.56 $X2=0
+ $Y2=0
cc_225 N_A_184_21#_M1015_g N_VGND_c_684_n 0.00341112f $X=1.935 $Y=0.56 $X2=0
+ $Y2=0
cc_226 N_A_184_21#_M1016_g N_VGND_c_684_n 0.00544582f $X=2.405 $Y=0.56 $X2=0
+ $Y2=0
cc_227 N_A_184_21#_M1015_g N_VGND_c_685_n 4.79042e-19 $X=1.935 $Y=0.56 $X2=0
+ $Y2=0
cc_228 N_A_184_21#_M1016_g N_VGND_c_685_n 0.00591224f $X=2.405 $Y=0.56 $X2=0
+ $Y2=0
cc_229 N_A_184_21#_c_141_n N_VGND_c_685_n 9.53459e-19 $X=2.53 $Y=1.16 $X2=0
+ $Y2=0
cc_230 N_A_184_21#_c_162_p N_VGND_c_685_n 0.00747245f $X=2.975 $Y=0.7 $X2=0
+ $Y2=0
cc_231 N_A_184_21#_c_248_p N_VGND_c_685_n 0.0136474f $X=2.7 $Y=0.7 $X2=0 $Y2=0
cc_232 N_A_184_21#_c_164_p N_VGND_c_685_n 0.0116817f $X=3.195 $Y=0.385 $X2=0
+ $Y2=0
cc_233 N_A_184_21#_c_145_n N_VGND_c_686_n 0.0085358f $X=4.895 $Y=0.385 $X2=0
+ $Y2=0
cc_234 N_A_184_21#_c_162_p N_VGND_c_687_n 0.00262114f $X=2.975 $Y=0.7 $X2=0
+ $Y2=0
cc_235 N_A_184_21#_c_169_p N_VGND_c_687_n 0.0678215f $X=4.71 $Y=0.385 $X2=0
+ $Y2=0
cc_236 N_A_184_21#_c_164_p N_VGND_c_687_n 0.0101706f $X=3.195 $Y=0.385 $X2=0
+ $Y2=0
cc_237 N_A_184_21#_c_145_n N_VGND_c_687_n 0.0172128f $X=4.895 $Y=0.385 $X2=0
+ $Y2=0
cc_238 N_A_184_21#_M1005_g N_VGND_c_689_n 0.00403236f $X=0.995 $Y=0.56 $X2=0
+ $Y2=0
cc_239 N_A_184_21#_M1007_g N_VGND_c_689_n 0.00341112f $X=1.465 $Y=0.56 $X2=0
+ $Y2=0
cc_240 N_A_184_21#_M1003_d N_VGND_c_691_n 0.00253533f $X=4.71 $Y=0.235 $X2=0
+ $Y2=0
cc_241 N_A_184_21#_M1005_g N_VGND_c_691_n 0.00609114f $X=0.995 $Y=0.56 $X2=0
+ $Y2=0
cc_242 N_A_184_21#_M1007_g N_VGND_c_691_n 0.00410013f $X=1.465 $Y=0.56 $X2=0
+ $Y2=0
cc_243 N_A_184_21#_M1015_g N_VGND_c_691_n 0.00410013f $X=1.935 $Y=0.56 $X2=0
+ $Y2=0
cc_244 N_A_184_21#_M1016_g N_VGND_c_691_n 0.00924731f $X=2.405 $Y=0.56 $X2=0
+ $Y2=0
cc_245 N_A_184_21#_c_162_p N_VGND_c_691_n 0.00505267f $X=2.975 $Y=0.7 $X2=0
+ $Y2=0
cc_246 N_A_184_21#_c_248_p N_VGND_c_691_n 8.89004e-19 $X=2.7 $Y=0.7 $X2=0 $Y2=0
cc_247 N_A_184_21#_c_169_p N_VGND_c_691_n 0.0527448f $X=4.71 $Y=0.385 $X2=0
+ $Y2=0
cc_248 N_A_184_21#_c_164_p N_VGND_c_691_n 0.00794239f $X=3.195 $Y=0.385 $X2=0
+ $Y2=0
cc_249 N_A_184_21#_c_145_n N_VGND_c_691_n 0.0129906f $X=4.895 $Y=0.385 $X2=0
+ $Y2=0
cc_250 N_A_184_21#_c_162_p A_606_47# 0.00267788f $X=2.975 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_251 N_A_184_21#_c_163_p A_606_47# 0.00181752f $X=3.085 $Y=0.615 $X2=-0.19
+ $Y2=-0.24
cc_252 N_A_184_21#_c_169_p A_606_47# 0.00834202f $X=4.71 $Y=0.385 $X2=-0.19
+ $Y2=-0.24
cc_253 N_A_184_21#_c_164_p A_606_47# 0.00115112f $X=3.195 $Y=0.385 $X2=-0.19
+ $Y2=-0.24
cc_254 N_A_184_21#_c_169_p A_719_47# 0.0109295f $X=4.71 $Y=0.385 $X2=-0.19
+ $Y2=-0.24
cc_255 N_A_184_21#_c_169_p A_836_47# 0.0105502f $X=4.71 $Y=0.385 $X2=-0.19
+ $Y2=-0.24
cc_256 N_D_c_286_n N_C_c_321_n 0.0235322f $X=2.955 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_257 N_D_c_287_n N_C_c_322_n 0.059645f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_258 D N_C_c_322_n 3.29137e-19 $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_259 N_D_c_286_n C 0.00253751f $X=2.955 $Y=0.995 $X2=0 $Y2=0
cc_260 N_D_c_287_n C 0.00211299f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_261 D C 0.0266489f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_262 N_D_c_287_n N_A_27_47#_c_363_n 0.0146023f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_263 N_D_c_287_n N_VPWR_c_550_n 0.00510113f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_264 N_D_c_287_n N_VPWR_c_543_n 0.00719739f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_265 N_D_c_287_n N_VPWR_c_556_n 0.00963324f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_266 N_D_c_286_n N_VGND_c_685_n 0.00587062f $X=2.955 $Y=0.995 $X2=0 $Y2=0
cc_267 N_D_c_286_n N_VGND_c_687_n 0.00401874f $X=2.955 $Y=0.995 $X2=0 $Y2=0
cc_268 N_D_c_286_n N_VGND_c_691_n 0.00626181f $X=2.955 $Y=0.995 $X2=0 $Y2=0
cc_269 N_C_c_321_n N_A_27_47#_c_354_n 0.0237144f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_270 C N_A_27_47#_c_354_n 0.0114751f $X=3.365 $Y=0.705 $X2=0 $Y2=0
cc_271 N_C_c_322_n N_A_27_47#_c_355_n 0.0565301f $X=3.545 $Y=1.41 $X2=0 $Y2=0
cc_272 N_C_c_322_n N_A_27_47#_c_363_n 0.0147595f $X=3.545 $Y=1.41 $X2=0 $Y2=0
cc_273 N_C_c_322_n N_A_27_47#_c_359_n 6.48745e-19 $X=3.545 $Y=1.41 $X2=0 $Y2=0
cc_274 C N_A_27_47#_c_359_n 0.0202367f $X=3.365 $Y=0.705 $X2=0 $Y2=0
cc_275 N_C_c_322_n N_VPWR_c_545_n 0.00452422f $X=3.545 $Y=1.41 $X2=0 $Y2=0
cc_276 N_C_c_322_n N_VPWR_c_550_n 0.00510113f $X=3.545 $Y=1.41 $X2=0 $Y2=0
cc_277 N_C_c_322_n N_VPWR_c_543_n 0.00723252f $X=3.545 $Y=1.41 $X2=0 $Y2=0
cc_278 N_C_c_321_n N_VGND_c_687_n 0.00367119f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_279 N_C_c_321_n N_VGND_c_691_n 0.00603216f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_280 C A_606_47# 0.00322241f $X=3.365 $Y=0.705 $X2=-0.19 $Y2=-0.24
cc_281 C A_719_47# 0.00587888f $X=3.365 $Y=0.705 $X2=-0.19 $Y2=-0.24
cc_282 N_A_27_47#_c_354_n N_A_912_21#_M1003_g 0.0307237f $X=4.105 $Y=0.995 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_355_n N_A_912_21#_M1003_g 0.0226707f $X=4.13 $Y=1.41 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_359_n N_A_912_21#_M1003_g 0.00141943f $X=4.165 $Y=1.16 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_355_n N_A_912_21#_c_452_n 0.0320852f $X=4.13 $Y=1.41 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_363_n N_A_912_21#_c_452_n 0.0168854f $X=4.77 $Y=2 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_365_n N_A_912_21#_c_452_n 0.0119723f $X=4.855 $Y=1.915 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_355_n N_A_912_21#_c_447_n 0.00327934f $X=4.13 $Y=1.41 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_357_n N_A_912_21#_c_447_n 0.0170008f $X=4.77 $Y=1.29 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_365_n N_A_912_21#_c_447_n 0.00145475f $X=4.855 $Y=1.915
+ $X2=0 $Y2=0
cc_291 N_A_27_47#_c_357_n N_A_912_21#_c_448_n 0.00619071f $X=4.77 $Y=1.29 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_365_n N_A_912_21#_c_448_n 0.0210622f $X=4.855 $Y=1.915 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_357_n N_A_912_21#_c_449_n 0.0137205f $X=4.77 $Y=1.29 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_363_n N_A_912_21#_c_457_n 0.00811893f $X=4.77 $Y=2 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_363_n N_VPWR_M1002_d 0.00612294f $X=4.77 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_296 N_A_27_47#_c_363_n N_VPWR_M1010_d 0.00360071f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_297 N_A_27_47#_c_363_n N_VPWR_M1019_d 0.00557992f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_298 N_A_27_47#_c_363_n N_VPWR_M1006_d 0.00658468f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_299 N_A_27_47#_c_363_n N_VPWR_M1018_d 0.00439432f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_300 N_A_27_47#_c_365_n N_VPWR_M1018_d 0.00847327f $X=4.855 $Y=1.915 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_363_n N_VPWR_c_544_n 0.00861424f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_302 N_A_27_47#_c_355_n N_VPWR_c_545_n 0.00320899f $X=4.13 $Y=1.41 $X2=0 $Y2=0
cc_303 N_A_27_47#_c_363_n N_VPWR_c_545_n 0.0222024f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_304 N_A_27_47#_c_362_n N_VPWR_c_548_n 0.0181194f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_305 N_A_27_47#_c_363_n N_VPWR_c_548_n 0.00238709f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_306 N_A_27_47#_c_363_n N_VPWR_c_549_n 0.00928399f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_307 N_A_27_47#_c_363_n N_VPWR_c_550_n 0.0127906f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_308 N_A_27_47#_c_363_n N_VPWR_c_551_n 0.0108559f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_309 N_A_27_47#_M1002_s N_VPWR_c_543_n 0.00238238f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_355_n N_VPWR_c_543_n 0.00706411f $X=4.13 $Y=1.41 $X2=0 $Y2=0
cc_311 N_A_27_47#_c_362_n N_VPWR_c_543_n 0.00991829f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_312 N_A_27_47#_c_363_n N_VPWR_c_543_n 0.0850937f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_313 N_A_27_47#_c_362_n N_VPWR_c_554_n 0.0161786f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_314 N_A_27_47#_c_363_n N_VPWR_c_554_n 0.0225111f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_315 N_A_27_47#_c_363_n N_VPWR_c_555_n 0.0196308f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_316 N_A_27_47#_c_363_n N_VPWR_c_556_n 0.0241133f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_317 N_A_27_47#_c_355_n N_VPWR_c_558_n 0.00510113f $X=4.13 $Y=1.41 $X2=0 $Y2=0
cc_318 N_A_27_47#_c_363_n N_VPWR_c_558_n 0.0120278f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_319 N_A_27_47#_c_363_n N_X_M1008_s 0.00475608f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_320 N_A_27_47#_c_363_n N_X_M1013_s 0.0048704f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_321 N_A_27_47#_c_363_n N_X_c_646_n 0.0452881f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_322 N_A_27_47#_c_363_n N_X_c_637_n 0.0190391f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_323 N_A_27_47#_c_354_n N_VGND_c_687_n 0.00367119f $X=4.105 $Y=0.995 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_M1014_s N_VGND_c_691_n 0.00559556f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_354_n N_VGND_c_691_n 0.00596085f $X=4.105 $Y=0.995 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_358_n N_VGND_c_691_n 0.00987844f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_327 N_A_27_47#_c_358_n N_VGND_c_692_n 0.0179125f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_328 N_A_912_21#_c_448_n N_A_N_M1012_g 0.00559584f $X=5.445 $Y=1.16 $X2=0
+ $Y2=0
cc_329 N_A_912_21#_c_450_n N_A_N_M1012_g 0.0177832f $X=6.095 $Y=0.74 $X2=0 $Y2=0
cc_330 N_A_912_21#_c_476_p N_A_N_M1012_g 0.00534863f $X=6.18 $Y=0.42 $X2=0 $Y2=0
cc_331 N_A_912_21#_c_448_n N_A_N_c_519_n 0.0135882f $X=5.445 $Y=1.16 $X2=0 $Y2=0
cc_332 N_A_912_21#_c_456_n N_A_N_c_520_n 0.0203397f $X=6.095 $Y=2 $X2=0 $Y2=0
cc_333 N_A_912_21#_c_479_p N_A_N_c_520_n 0.00460257f $X=6.18 $Y=2.3 $X2=0 $Y2=0
cc_334 N_A_912_21#_c_448_n A_N 0.0235853f $X=5.445 $Y=1.16 $X2=0 $Y2=0
cc_335 N_A_912_21#_c_449_n A_N 0.00130291f $X=5.445 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A_912_21#_c_450_n A_N 0.0274908f $X=6.095 $Y=0.74 $X2=0 $Y2=0
cc_337 N_A_912_21#_c_456_n A_N 0.0187174f $X=6.095 $Y=2 $X2=0 $Y2=0
cc_338 N_A_912_21#_c_448_n N_A_N_c_518_n 0.00111951f $X=5.445 $Y=1.16 $X2=0
+ $Y2=0
cc_339 N_A_912_21#_c_449_n N_A_N_c_518_n 0.0228023f $X=5.445 $Y=1.16 $X2=0 $Y2=0
cc_340 N_A_912_21#_c_450_n N_A_N_c_518_n 0.00155154f $X=6.095 $Y=0.74 $X2=0
+ $Y2=0
cc_341 N_A_912_21#_c_456_n N_A_N_c_518_n 6.43001e-19 $X=6.095 $Y=2 $X2=0 $Y2=0
cc_342 N_A_912_21#_c_456_n N_VPWR_M1018_d 0.00287786f $X=6.095 $Y=2 $X2=0 $Y2=0
cc_343 N_A_912_21#_c_457_n N_VPWR_M1018_d 0.00229205f $X=5.53 $Y=2 $X2=0 $Y2=0
cc_344 N_A_912_21#_c_456_n N_VPWR_c_546_n 0.0202626f $X=6.095 $Y=2 $X2=0 $Y2=0
cc_345 N_A_912_21#_c_457_n N_VPWR_c_546_n 0.014249f $X=5.53 $Y=2 $X2=0 $Y2=0
cc_346 N_A_912_21#_c_452_n N_VPWR_c_551_n 0.0155007f $X=4.66 $Y=1.41 $X2=0 $Y2=0
cc_347 N_A_912_21#_c_456_n N_VPWR_c_552_n 0.00386522f $X=6.095 $Y=2 $X2=0 $Y2=0
cc_348 N_A_912_21#_c_479_p N_VPWR_c_552_n 0.0116326f $X=6.18 $Y=2.3 $X2=0 $Y2=0
cc_349 N_A_912_21#_M1001_d N_VPWR_c_543_n 0.00380573f $X=6.035 $Y=2.065 $X2=0
+ $Y2=0
cc_350 N_A_912_21#_c_452_n N_VPWR_c_543_n 0.00824f $X=4.66 $Y=1.41 $X2=0 $Y2=0
cc_351 N_A_912_21#_c_456_n N_VPWR_c_543_n 0.00809766f $X=6.095 $Y=2 $X2=0 $Y2=0
cc_352 N_A_912_21#_c_457_n N_VPWR_c_543_n 8.59428e-19 $X=5.53 $Y=2 $X2=0 $Y2=0
cc_353 N_A_912_21#_c_479_p N_VPWR_c_543_n 0.00643448f $X=6.18 $Y=2.3 $X2=0 $Y2=0
cc_354 N_A_912_21#_c_452_n N_VPWR_c_558_n 0.00510113f $X=4.66 $Y=1.41 $X2=0
+ $Y2=0
cc_355 N_A_912_21#_c_451_n N_VGND_M1012_s 0.0016104f $X=5.53 $Y=0.74 $X2=0 $Y2=0
cc_356 N_A_912_21#_M1003_g N_VGND_c_686_n 0.00226228f $X=4.635 $Y=0.56 $X2=0
+ $Y2=0
cc_357 N_A_912_21#_c_449_n N_VGND_c_686_n 6.88104e-19 $X=5.445 $Y=1.16 $X2=0
+ $Y2=0
cc_358 N_A_912_21#_c_450_n N_VGND_c_686_n 0.0129893f $X=6.095 $Y=0.74 $X2=0
+ $Y2=0
cc_359 N_A_912_21#_c_451_n N_VGND_c_686_n 0.011044f $X=5.53 $Y=0.74 $X2=0 $Y2=0
cc_360 N_A_912_21#_c_476_p N_VGND_c_686_n 0.00886884f $X=6.18 $Y=0.42 $X2=0
+ $Y2=0
cc_361 N_A_912_21#_M1003_g N_VGND_c_687_n 0.00367119f $X=4.635 $Y=0.56 $X2=0
+ $Y2=0
cc_362 N_A_912_21#_c_451_n N_VGND_c_687_n 4.7797e-19 $X=5.53 $Y=0.74 $X2=0 $Y2=0
cc_363 N_A_912_21#_c_450_n N_VGND_c_690_n 0.00635723f $X=6.095 $Y=0.74 $X2=0
+ $Y2=0
cc_364 N_A_912_21#_c_476_p N_VGND_c_690_n 0.0116627f $X=6.18 $Y=0.42 $X2=0 $Y2=0
cc_365 N_A_912_21#_M1012_d N_VGND_c_691_n 0.00430827f $X=5.995 $Y=0.235 $X2=0
+ $Y2=0
cc_366 N_A_912_21#_M1003_g N_VGND_c_691_n 0.0068535f $X=4.635 $Y=0.56 $X2=0
+ $Y2=0
cc_367 N_A_912_21#_c_450_n N_VGND_c_691_n 0.0106696f $X=6.095 $Y=0.74 $X2=0
+ $Y2=0
cc_368 N_A_912_21#_c_451_n N_VGND_c_691_n 0.00148077f $X=5.53 $Y=0.74 $X2=0
+ $Y2=0
cc_369 N_A_912_21#_c_476_p N_VGND_c_691_n 0.00644035f $X=6.18 $Y=0.42 $X2=0
+ $Y2=0
cc_370 N_A_N_c_520_n N_VPWR_c_547_n 0.00967552f $X=5.945 $Y=1.99 $X2=0 $Y2=0
cc_371 N_A_N_c_520_n N_VPWR_c_552_n 0.00516667f $X=5.945 $Y=1.99 $X2=0 $Y2=0
cc_372 N_A_N_c_520_n N_VPWR_c_543_n 0.00887641f $X=5.945 $Y=1.99 $X2=0 $Y2=0
cc_373 N_A_N_M1012_g N_VGND_c_686_n 0.00957124f $X=5.92 $Y=0.445 $X2=0 $Y2=0
cc_374 N_A_N_M1012_g N_VGND_c_690_n 0.00428022f $X=5.92 $Y=0.445 $X2=0 $Y2=0
cc_375 N_A_N_M1012_g N_VGND_c_691_n 0.00825815f $X=5.92 $Y=0.445 $X2=0 $Y2=0
cc_376 N_VPWR_c_543_n N_X_M1008_s 0.00338665f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_377 N_VPWR_c_543_n N_X_M1013_s 0.00338665f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_378 N_VPWR_M1010_d N_X_c_646_n 0.00386574f $X=1.58 $Y=1.485 $X2=0 $Y2=0
cc_379 N_X_c_642_n N_VGND_M1007_d 0.00440003f $X=2.11 $Y=0.735 $X2=0 $Y2=0
cc_380 N_X_c_641_n N_VGND_c_682_n 0.0130167f $X=1.255 $Y=0.42 $X2=0 $Y2=0
cc_381 N_X_c_642_n N_VGND_c_683_n 0.0188758f $X=2.11 $Y=0.735 $X2=0 $Y2=0
cc_382 N_X_c_651_n N_VGND_c_683_n 0.01316f $X=2.195 $Y=0.42 $X2=0 $Y2=0
cc_383 N_X_c_642_n N_VGND_c_684_n 0.00314446f $X=2.11 $Y=0.735 $X2=0 $Y2=0
cc_384 N_X_c_651_n N_VGND_c_684_n 0.0114519f $X=2.195 $Y=0.42 $X2=0 $Y2=0
cc_385 N_X_c_641_n N_VGND_c_689_n 0.0116048f $X=1.255 $Y=0.42 $X2=0 $Y2=0
cc_386 N_X_c_642_n N_VGND_c_689_n 0.00235782f $X=2.11 $Y=0.735 $X2=0 $Y2=0
cc_387 X N_VGND_c_689_n 0.00238407f $X=1.085 $Y=0.765 $X2=0 $Y2=0
cc_388 N_X_M1005_s N_VGND_c_691_n 0.00310807f $X=1.07 $Y=0.235 $X2=0 $Y2=0
cc_389 N_X_M1015_s N_VGND_c_691_n 0.00466393f $X=2.01 $Y=0.235 $X2=0 $Y2=0
cc_390 N_X_c_641_n N_VGND_c_691_n 0.00646998f $X=1.255 $Y=0.42 $X2=0 $Y2=0
cc_391 N_X_c_642_n N_VGND_c_691_n 0.0113475f $X=2.11 $Y=0.735 $X2=0 $Y2=0
cc_392 N_X_c_651_n N_VGND_c_691_n 0.0064389f $X=2.195 $Y=0.42 $X2=0 $Y2=0
cc_393 X N_VGND_c_691_n 0.0044122f $X=1.085 $Y=0.765 $X2=0 $Y2=0
cc_394 N_VGND_c_691_n A_606_47# 0.00338587f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_395 N_VGND_c_691_n A_719_47# 0.0035526f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_396 N_VGND_c_691_n A_836_47# 0.00309241f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
