# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nor4_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor4_6 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.42000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.505000 1.075000 2.875000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.325000 1.075000 5.695000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.665000 1.075000 9.035000 1.285000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  1.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.395000 1.075000 11.085000 1.285000 ;
    END
  END D
  PIN VGND
    ANTENNADIFFAREA  3.419000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.420000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  0.870000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.420000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  2.976000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.585000 0.255000  0.915000 0.725000 ;
        RECT  0.585000 0.725000 11.835000 0.905000 ;
        RECT  1.525000 0.255000  1.855000 0.725000 ;
        RECT  2.465000 0.255000  2.795000 0.725000 ;
        RECT  3.405000 0.255000  3.735000 0.725000 ;
        RECT  4.345000 0.255000  4.675000 0.725000 ;
        RECT  5.285000 0.255000  5.615000 0.725000 ;
        RECT  6.745000 0.255000  7.075000 0.725000 ;
        RECT  7.685000 0.255000  8.015000 0.725000 ;
        RECT  8.625000 0.255000  8.955000 0.725000 ;
        RECT  9.565000 0.255000  9.895000 0.725000 ;
        RECT  9.605000 1.455000 11.835000 1.625000 ;
        RECT  9.605000 1.625000  9.855000 2.125000 ;
        RECT 10.505000 0.255000 10.835000 0.725000 ;
        RECT 10.545000 1.625000 10.795000 2.125000 ;
        RECT 11.445000 0.255000 11.835000 0.725000 ;
        RECT 11.445000 0.905000 11.835000 1.455000 ;
        RECT 11.445000 1.625000 11.835000 2.125000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.420000 0.085000 ;
      RECT  0.000000  2.635000 12.420000 2.805000 ;
      RECT  0.115000  0.085000  0.415000 0.905000 ;
      RECT  0.115000  1.455000  3.225000 1.625000 ;
      RECT  0.115000  1.625000  0.405000 2.465000 ;
      RECT  0.625000  1.795000  0.875000 2.635000 ;
      RECT  1.085000  0.085000  1.355000 0.555000 ;
      RECT  1.095000  1.625000  1.345000 2.465000 ;
      RECT  1.565000  1.795000  1.815000 2.635000 ;
      RECT  2.025000  0.085000  2.295000 0.555000 ;
      RECT  2.035000  1.625000  2.285000 2.465000 ;
      RECT  2.505000  1.795000  2.755000 2.635000 ;
      RECT  2.965000  0.085000  3.235000 0.555000 ;
      RECT  2.975000  1.625000  3.225000 2.295000 ;
      RECT  2.975000  2.295000  6.085000 2.465000 ;
      RECT  3.445000  1.455000  8.915000 1.625000 ;
      RECT  3.445000  1.625000  3.695000 2.125000 ;
      RECT  3.905000  0.085000  4.175000 0.555000 ;
      RECT  3.915000  1.795000  4.165000 2.295000 ;
      RECT  4.385000  1.625000  4.635000 2.125000 ;
      RECT  4.845000  0.085000  5.115000 0.555000 ;
      RECT  4.855000  1.795000  5.105000 2.295000 ;
      RECT  5.325000  1.625000  5.575000 2.125000 ;
      RECT  5.785000  0.085000  6.575000 0.555000 ;
      RECT  5.795000  1.795000  6.085000 2.295000 ;
      RECT  6.275000  1.795000  6.565000 2.295000 ;
      RECT  6.275000  2.295000 12.255000 2.465000 ;
      RECT  6.785000  1.625000  7.035000 2.125000 ;
      RECT  7.245000  0.085000  7.515000 0.555000 ;
      RECT  7.255000  1.795000  7.505000 2.295000 ;
      RECT  7.725000  1.625000  7.975000 2.125000 ;
      RECT  8.185000  0.085000  8.455000 0.555000 ;
      RECT  8.195000  1.795000  8.445000 2.295000 ;
      RECT  8.665000  1.625000  8.915000 2.125000 ;
      RECT  9.125000  0.085000  9.395000 0.555000 ;
      RECT  9.135000  1.455000  9.385000 2.295000 ;
      RECT 10.065000  0.085000 10.335000 0.555000 ;
      RECT 10.075000  1.795000 10.325000 2.295000 ;
      RECT 11.005000  0.085000 11.275000 0.555000 ;
      RECT 11.015000  1.795000 11.265000 2.295000 ;
      RECT 12.005000  0.085000 12.255000 0.905000 ;
      RECT 12.005000  1.455000 12.255000 2.295000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4_6
END LIBRARY
