# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a21oi_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.815000 1.065000 4.400000 1.310000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.250000 1.065000 2.645000 1.480000 ;
        RECT 2.250000 1.480000 6.070000 1.705000 ;
        RECT 4.675000 1.075000 6.070000 1.480000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.400000 1.035000 ;
        RECT 0.090000 1.035000 1.580000 1.415000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.523000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.630000 1.585000 2.080000 1.705000 ;
        RECT 0.630000 1.705000 1.895000 2.035000 ;
        RECT 0.645000 0.370000 0.835000 0.615000 ;
        RECT 0.645000 0.615000 1.795000 0.695000 ;
        RECT 0.645000 0.695000 4.305000 0.865000 ;
        RECT 1.605000 0.255000 1.795000 0.615000 ;
        RECT 1.750000 0.865000 4.305000 0.895000 ;
        RECT 1.750000 0.895000 2.080000 1.585000 ;
        RECT 2.475000 0.675000 4.305000 0.695000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.805000 ;
      RECT 0.180000  1.795000 0.375000 2.215000 ;
      RECT 0.180000  2.215000 2.315000 2.465000 ;
      RECT 1.005000  0.085000 1.385000 0.445000 ;
      RECT 1.005000  2.205000 2.315000 2.215000 ;
      RECT 1.985000  0.085000 2.315000 0.525000 ;
      RECT 2.115000  1.875000 6.225000 2.105000 ;
      RECT 2.115000  2.105000 2.315000 2.205000 ;
      RECT 2.485000  0.255000 4.785000 0.505000 ;
      RECT 2.485000  2.275000 2.865000 2.635000 ;
      RECT 3.085000  2.105000 3.275000 2.465000 ;
      RECT 3.445000  2.275000 3.825000 2.635000 ;
      RECT 4.045000  2.105000 4.235000 2.465000 ;
      RECT 4.405000  2.275000 4.785000 2.635000 ;
      RECT 4.525000  0.505000 4.785000 0.735000 ;
      RECT 4.525000  0.735000 5.745000 0.905000 ;
      RECT 5.005000  0.085000 5.195000 0.565000 ;
      RECT 5.005000  2.105000 5.185000 2.465000 ;
      RECT 5.365000  0.255000 5.745000 0.735000 ;
      RECT 5.365000  2.275000 5.745000 2.635000 ;
      RECT 5.965000  0.085000 6.225000 0.885000 ;
      RECT 5.965000  2.105000 6.225000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21oi_4
