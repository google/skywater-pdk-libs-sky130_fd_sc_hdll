* NGSPICE file created from sky130_fd_sc_hdll__sdlclkp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__sdlclkp_4 CLK GATE SCE VGND VNB VPB VPWR GCLK
M1000 a_425_47# a_277_243# a_310_47# VNB nshort w=360000u l=150000u
+  ad=2.196e+11p pd=1.96e+06u as=1.53e+11p ps=1.57e+06u
M1001 a_27_47# GATE VGND VNB nshort w=420000u l=150000u
+  ad=2.664e+11p pd=2.97e+06u as=1.3078e+12p ps=1.141e+07u
M1002 a_27_47# GATE a_117_369# VPB phighvt w=640000u l=180000u
+  ad=2.373e+11p pd=2.08e+06u as=1.472e+11p ps=1.74e+06u
M1003 GCLK a_1125_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=7.15e+11p pd=5.43e+06u as=2.2235e+12p ps=1.837e+07u
M1004 GCLK a_1125_47# VGND VNB nshort w=650000u l=150000u
+  ad=5.3625e+11p pd=4.25e+06u as=0p ps=0u
M1005 a_421_413# a_280_21# a_310_47# VPB phighvt w=420000u l=180000u
+  ad=1.806e+11p pd=1.7e+06u as=1.47e+11p ps=1.54e+06u
M1006 a_280_21# CLK VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1007 a_117_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_280_21# a_277_243# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1009 VPWR CLK a_1125_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1010 VPWR a_505_315# a_421_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1125_47# a_505_315# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_310_47# a_277_243# a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_280_21# a_277_243# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1014 VGND a_1125_47# GCLK VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_505_315# a_425_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND SCE a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 GCLK a_1125_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1217_47# a_505_315# a_1125_47# VNB nshort w=650000u l=150000u
+  ad=1.365e+11p pd=1.72e+06u as=2.015e+11p ps=1.92e+06u
M1019 a_505_315# a_310_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1020 VPWR a_1125_47# GCLK VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND CLK a_1217_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 GCLK a_1125_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_280_21# CLK VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1024 VGND a_1125_47# GCLK VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_1125_47# GCLK VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_310_47# a_280_21# a_27_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_505_315# a_310_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
.ends

