* File: sky130_fd_sc_hdll__o32ai_1.spice
* Created: Thu Aug 27 19:22:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o32ai_1.pex.spice"
.subckt sky130_fd_sc_hdll__o32ai_1  VNB VPB B1 B2 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1006 N_Y_M1006_d N_B1_M1006_g N_A_27_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.121875 AS=0.2015 PD=1.025 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1005 N_A_27_47#_M1005_d N_B2_M1005_g N_Y_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.09425 AS=0.121875 PD=0.94 PS=1.025 NRD=0 NRS=18.456 M=1 R=4.33333
+ SA=75000.8 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_A3_M1001_g N_A_27_47#_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.203125 AS=0.09425 PD=1.275 PS=0.94 NRD=20.304 NRS=2.76 M=1 R=4.33333
+ SA=75001.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1008 N_A_27_47#_M1008_d N_A2_M1008_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.203125 PD=0.92 PS=1.275 NRD=0 NRS=43.38 M=1 R=4.33333 SA=75002
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A1_M1007_g N_A_27_47#_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.195 AS=0.08775 PD=1.9 PS=0.92 NRD=2.76 NRS=0 M=1 R=4.33333 SA=75002.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 A_117_297# N_B1_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.115
+ AS=0.27 PD=1.23 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90002.4 A=0.18 P=2.36 MULT=1
MM1002 N_Y_M1002_d N_B2_M1002_g A_117_297# VPB PHIGHVT L=0.18 W=1 AD=0.2575
+ AS=0.115 PD=1.515 PS=1.23 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90000.6
+ SB=90002 A=0.18 P=2.36 MULT=1
MM1009 A_338_297# N_A3_M1009_g N_Y_M1002_d VPB PHIGHVT L=0.18 W=1 AD=0.2275
+ AS=0.2575 PD=1.455 PS=1.515 NRD=33.9628 NRS=45.2903 M=1 R=5.55556 SA=90001.3
+ SB=90001.3 A=0.18 P=2.36 MULT=1
MM1004 A_465_297# N_A2_M1004_g A_338_297# VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.2275 PD=1.29 PS=1.455 NRD=17.7103 NRS=33.9628 M=1 R=5.55556 SA=90001.9
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g A_465_297# VPB PHIGHVT L=0.18 W=1 AD=0.29
+ AS=0.145 PD=2.58 PS=1.29 NRD=0.9653 NRS=17.7103 M=1 R=5.55556 SA=90002.4
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hdll__o32ai_1.pxi.spice"
*
.ends
*
*
