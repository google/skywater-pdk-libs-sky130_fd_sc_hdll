* File: sky130_fd_sc_hdll__nand2_2.pex.spice
* Created: Wed Sep  2 08:36:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND2_2%B 1 3 4 6 7 9 10 12 13 14 22
c45 14 0 1.58116e-19 $X=0.695 $Y=1.19
c46 10 0 9.09144e-20 $X=0.99 $Y=0.995
r47 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r48 20 22 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=0.73 $Y=1.202
+ $X2=0.965 $Y2=1.202
r49 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.73 $Y2=1.202
r50 17 18 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r51 14 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.73
+ $Y=1.16 $X2=0.73 $Y2=1.16
r52 13 14 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=1.2
+ $X2=0.695 $Y2=1.2
r53 10 23 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r54 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r55 7 22 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r56 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r57 4 18 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r58 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r59 1 17 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.202
r60 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_2%A 1 3 4 6 7 9 10 12 13 14 22 27
c46 22 0 1.58116e-19 $X=1.905 $Y=1.202
r47 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=1.93 $Y2=1.202
r48 20 22 46.9316 $w=3.8e-07 $l=3.7e-07 $layer=POLY_cond $X=1.535 $Y=1.202
+ $X2=1.905 $Y2=1.202
r49 20 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.535
+ $Y=1.16 $X2=1.535 $Y2=1.16
r50 18 20 12.6842 $w=3.8e-07 $l=1e-07 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.535 $Y2=1.202
r51 17 18 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.202
+ $X2=1.435 $Y2=1.202
r52 14 27 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=1.63 $Y=1.2
+ $X2=1.535 $Y2=1.2
r53 13 27 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=1.255 $Y=1.2
+ $X2=1.535 $Y2=1.2
r54 10 23 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r55 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r56 7 22 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r57 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r58 4 18 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r59 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r60 1 17 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.202
r61 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995 $X2=1.41
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_2%VPWR 1 2 3 10 12 16 20 22 26 28 32 33 39
+ 42
r40 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r41 40 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r42 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r43 33 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r44 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r45 30 42 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=2.31 $Y=2.72
+ $X2=2.182 $Y2=2.72
r46 30 32 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.31 $Y=2.72
+ $X2=2.53 $Y2=2.72
r47 28 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r48 28 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r49 24 42 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.182 $Y=2.635
+ $X2=2.182 $Y2=2.72
r50 24 26 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=2.182 $Y=2.635
+ $X2=2.182 $Y2=2
r51 23 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.72 $X2=1.2
+ $Y2=2.72
r52 22 42 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=2.182 $Y2=2.72
r53 22 23 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=1.285 $Y2=2.72
r54 18 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.72
r55 18 20 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r56 17 36 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r57 16 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.72 $X2=1.2
+ $Y2=2.72
r58 16 17 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=0.345 $Y2=2.72
r59 12 15 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=0.215 $Y=1.66
+ $X2=0.215 $Y2=2.34
r60 10 36 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r61 10 15 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2.34
r62 3 26 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r63 2 20 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r64 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r65 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_2%Y 1 2 3 10 12 14 16 22 26 27 28 34 46
c54 16 0 9.09144e-20 $X=1.95 $Y=0.78
r55 28 46 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.09 $Y=1.58
+ $X2=2.095 $Y2=1.58
r56 27 28 11.5244 $w=2.78e-07 $l=2.8e-07 $layer=LI1_cond $X=2.09 $Y=1.19
+ $X2=2.09 $Y2=1.47
r57 26 34 3.22874 $w=2.8e-07 $l=1.25e-07 $layer=LI1_cond $X=2.09 $Y=0.78
+ $X2=2.09 $Y2=0.905
r58 26 27 11.1128 $w=2.78e-07 $l=2.7e-07 $layer=LI1_cond $X=2.09 $Y=0.92
+ $X2=2.09 $Y2=1.19
r59 26 34 0.61738 $w=2.78e-07 $l=1.5e-08 $layer=LI1_cond $X=2.09 $Y=0.92
+ $X2=2.09 $Y2=0.905
r60 20 28 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.645 $Y=1.58
+ $X2=2.09 $Y2=1.58
r61 20 22 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.645 $Y2=2.34
r62 16 26 3.61619 $w=2.5e-07 $l=1.4e-07 $layer=LI1_cond $X=1.95 $Y=0.78 $X2=2.09
+ $Y2=0.78
r63 16 18 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=1.95 $Y=0.78
+ $X2=1.67 $Y2=0.78
r64 15 25 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.705 $Y2=1.58
r65 14 20 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=1.58
+ $X2=1.645 $Y2=1.58
r66 14 15 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.455 $Y=1.58
+ $X2=0.895 $Y2=1.58
r67 10 25 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=1.58
r68 10 12 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=2.34
r69 3 20 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r70 3 22 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
r71 2 25 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r72 2 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r73 1 18 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_2%A_27_47# 1 2 3 12 14 15 16 17 20
r42 18 23 3.94658 $w=2.3e-07 $l=1.5e-07 $layer=LI1_cond $X=1.285 $Y=0.37
+ $X2=1.135 $Y2=0.37
r43 18 20 42.8408 $w=2.28e-07 $l=8.55e-07 $layer=LI1_cond $X=1.285 $Y=0.37
+ $X2=2.14 $Y2=0.37
r44 17 25 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0.715
+ $X2=1.135 $Y2=0.8
r45 16 23 3.02571 $w=3e-07 $l=1.15e-07 $layer=LI1_cond $X=1.135 $Y=0.485
+ $X2=1.135 $Y2=0.37
r46 16 17 8.8354 $w=2.98e-07 $l=2.3e-07 $layer=LI1_cond $X=1.135 $Y=0.485
+ $X2=1.135 $Y2=0.715
r47 14 25 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.985 $Y=0.8
+ $X2=1.135 $Y2=0.8
r48 14 15 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.985 $Y=0.8
+ $X2=0.425 $Y2=0.8
r49 10 15 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.255 $Y=0.715
+ $X2=0.425 $Y2=0.8
r50 10 12 11.355 $w=3.38e-07 $l=3.35e-07 $layer=LI1_cond $X=0.255 $Y=0.715
+ $X2=0.255 $Y2=0.38
r51 3 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.38
r52 2 25 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.72
r53 2 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.38
r54 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_2%VGND 1 8 10 17 18 21 24
r32 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r33 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r34 15 18 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r35 15 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r36 14 17 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r37 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r38 12 21 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.73
+ $Y2=0
r39 12 14 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=1.15
+ $Y2=0
r40 10 22 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r41 10 24 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r42 6 21 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085 $X2=0.73
+ $Y2=0
r43 6 8 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=0.085 $X2=0.73
+ $Y2=0.38
r44 1 8 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

