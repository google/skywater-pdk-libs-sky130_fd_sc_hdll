* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__clkbuf_1 A VGND VNB VPB VPWR X
X0 X a_75_212# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=180000u
X1 VPWR A a_75_212# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=180000u
X2 X a_75_212# VGND SUBS sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X3 VGND A a_75_212# SUBS sky130_fd_pr__nfet_01v8 w=520000u l=150000u
.ends
