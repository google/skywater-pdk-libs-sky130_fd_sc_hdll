# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__o32ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o32ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.200000 1.075000 6.295000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.720000 1.075000 4.930000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.655000 1.075000 3.365000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.075000 1.815000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.895000 1.325000 ;
    END
  END B2
  PIN VGND
    ANTENNADIFFAREA  1.059500 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  0.850000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  1.061000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.655000 2.245000 0.905000 ;
        RECT 0.515000 1.495000 3.405000 1.665000 ;
        RECT 0.515000 1.665000 0.895000 2.095000 ;
        RECT 1.985000 0.905000 2.245000 1.105000 ;
        RECT 1.985000 1.105000 2.370000 1.495000 ;
        RECT 3.025000 1.665000 3.405000 2.085000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.090000  0.255000 2.655000 0.485000 ;
      RECT 0.090000  0.485000 0.345000 0.905000 ;
      RECT 0.090000  1.495000 0.345000 2.295000 ;
      RECT 0.090000  2.295000 1.365000 2.465000 ;
      RECT 1.115000  1.835000 2.305000 2.005000 ;
      RECT 1.115000  2.005000 1.365000 2.295000 ;
      RECT 1.585000  2.175000 1.755000 2.635000 ;
      RECT 1.925000  2.005000 2.305000 2.455000 ;
      RECT 2.485000  0.485000 2.655000 0.715000 ;
      RECT 2.485000  0.715000 6.305000 0.905000 ;
      RECT 2.585000  1.835000 2.835000 2.255000 ;
      RECT 2.585000  2.255000 4.835000 2.445000 ;
      RECT 2.870000  0.085000 3.250000 0.545000 ;
      RECT 3.435000  0.255000 3.815000 0.715000 ;
      RECT 3.625000  1.495000 3.795000 2.255000 ;
      RECT 4.015000  1.495000 5.825000 1.665000 ;
      RECT 4.015000  1.665000 4.345000 2.085000 ;
      RECT 4.035000  0.085000 4.205000 0.545000 ;
      RECT 4.505000  0.255000 5.175000 0.715000 ;
      RECT 4.585000  1.835000 4.835000 2.255000 ;
      RECT 5.070000  1.835000 5.275000 2.635000 ;
      RECT 5.355000  0.085000 5.735000 0.545000 ;
      RECT 5.495000  1.665000 5.825000 2.460000 ;
      RECT 5.975000  0.255000 6.305000 0.715000 ;
      RECT 6.045000  1.495000 6.265000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o32ai_2
END LIBRARY
