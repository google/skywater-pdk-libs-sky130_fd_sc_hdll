* File: sky130_fd_sc_hdll__or2b_4.pex.spice
* Created: Thu Aug 27 19:23:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR2B_4%B_N 2 3 5 8 10 11 12 21
c26 10 0 1.70525e-19 $X=0.23 $Y=1.19
r27 20 21 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r28 17 20 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.495 $Y2=1.16
r29 11 12 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=0.257 $Y=1.53
+ $X2=0.257 $Y2=1.87
r30 10 11 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.257 $Y=1.16
+ $X2=0.257 $Y2=1.53
r31 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r32 6 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.16
r33 6 8 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.475
r34 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r35 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.89 $X2=0.495
+ $Y2=1.99
r36 1 20 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r37 1 2 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_4%A_27_53# 1 2 7 9 10 12 13 14 17 19 20 21 23
c61 13 0 1.70525e-19 $X=1.395 $Y=1.16
r62 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.055
+ $Y=1.16 $X2=1.055 $Y2=1.16
r63 21 27 9.1679 $w=4.03e-07 $l=2.46037e-07 $layer=LI1_cond $X=0.73 $Y=1.325
+ $X2=0.907 $Y2=1.16
r64 21 23 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=0.73 $Y=1.325
+ $X2=0.73 $Y2=2.2
r65 19 27 10.2928 $w=4.03e-07 $l=4.52416e-07 $layer=LI1_cond $X=0.645 $Y=0.82
+ $X2=0.907 $Y2=1.16
r66 19 20 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.645 $Y=0.82
+ $X2=0.42 $Y2=0.82
r67 15 20 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=0.265 $Y=0.735
+ $X2=0.42 $Y2=0.82
r68 15 17 10.7809 $w=3.08e-07 $l=2.9e-07 $layer=LI1_cond $X=0.265 $Y=0.735
+ $X2=0.265 $Y2=0.445
r69 13 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.395 $Y=1.16
+ $X2=1.055 $Y2=1.16
r70 13 14 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=1.16
+ $X2=1.395 $Y2=0.995
r71 10 14 34.7346 $w=1.65e-07 $l=4.66771e-07 $layer=POLY_cond $X=1.505 $Y=1.41
+ $X2=1.395 $Y2=0.995
r72 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.505 $Y=1.41
+ $X2=1.505 $Y2=1.985
r73 7 14 34.7346 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.47 $Y=0.995
+ $X2=1.395 $Y2=0.995
r74 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.47 $Y=0.995 $X2=1.47
+ $Y2=0.56
r75 2 23 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.065 $X2=0.73 $Y2=2.2
r76 1 17 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_4%A 1 3 4 6 7 15
c31 4 0 8.22775e-20 $X=1.915 $Y=1.41
r32 11 15 6.65455 $w=1.98e-07 $l=1.2e-07 $layer=LI1_cond $X=1.95 $Y=1.175
+ $X2=2.07 $Y2=1.175
r33 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.95
+ $Y=1.16 $X2=1.95 $Y2=1.16
r34 7 15 8.31818 $w=1.98e-07 $l=1.5e-07 $layer=LI1_cond $X=2.22 $Y=1.175
+ $X2=2.07 $Y2=1.175
r35 4 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=1.915 $Y=1.41
+ $X2=1.975 $Y2=1.16
r36 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.915 $Y=1.41
+ $X2=1.915 $Y2=1.985
r37 1 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.89 $Y=0.995
+ $X2=1.975 $Y2=1.16
r38 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.89 $Y=0.995 $X2=1.89
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_4%A_229_297# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 33 38 41 43 45 46 49 52 54 66
c126 45 0 8.22775e-20 $X=2.775 $Y=1.245
r127 66 67 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.865 $Y=1.202
+ $X2=3.89 $Y2=1.202
r128 63 64 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.37 $Y=1.202
+ $X2=3.395 $Y2=1.202
r129 62 63 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=2.925 $Y=1.202
+ $X2=3.37 $Y2=1.202
r130 61 62 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.9 $Y=1.202
+ $X2=2.925 $Y2=1.202
r131 58 59 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.43 $Y=1.202
+ $X2=2.455 $Y2=1.202
r132 57 61 5.83065 $w=3.72e-07 $l=4.5e-08 $layer=POLY_cond $X=2.855 $Y=1.202
+ $X2=2.9 $Y2=1.202
r133 57 59 51.828 $w=3.72e-07 $l=4e-07 $layer=POLY_cond $X=2.855 $Y=1.202
+ $X2=2.455 $Y2=1.202
r134 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.855
+ $Y=1.16 $X2=2.855 $Y2=1.16
r135 53 54 7.18162 $w=3.78e-07 $l=1.7e-07 $layer=LI1_cond $X=1.592 $Y=0.735
+ $X2=1.592 $Y2=0.905
r136 50 66 29.8011 $w=3.72e-07 $l=2.3e-07 $layer=POLY_cond $X=3.635 $Y=1.202
+ $X2=3.865 $Y2=1.202
r137 50 64 31.0968 $w=3.72e-07 $l=2.4e-07 $layer=POLY_cond $X=3.635 $Y=1.202
+ $X2=3.395 $Y2=1.202
r138 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.635
+ $Y=1.16 $X2=3.635 $Y2=1.16
r139 47 56 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=1.16
+ $X2=2.775 $Y2=1.16
r140 47 49 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.86 $Y=1.16
+ $X2=3.635 $Y2=1.16
r141 45 56 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=1.245
+ $X2=2.775 $Y2=1.16
r142 45 46 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.775 $Y=1.245
+ $X2=2.775 $Y2=1.445
r143 44 52 4.24538 $w=1.7e-07 $l=5.37215e-07 $layer=LI1_cond $X=1.56 $Y=1.53
+ $X2=1.04 $Y2=1.495
r144 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.69 $Y=1.53
+ $X2=2.775 $Y2=1.445
r145 43 44 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=2.69 $Y=1.53
+ $X2=1.56 $Y2=1.53
r146 41 53 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.655 $Y=0.4
+ $X2=1.655 $Y2=0.735
r147 38 52 2.59952 $w=3.7e-07 $l=4.34281e-07 $layer=LI1_cond $X=1.45 $Y=1.445
+ $X2=1.04 $Y2=1.495
r148 38 54 28.2872 $w=2.18e-07 $l=5.4e-07 $layer=LI1_cond $X=1.45 $Y=1.445
+ $X2=1.45 $Y2=0.905
r149 33 35 15.641 $w=5.18e-07 $l=6.8e-07 $layer=LI1_cond $X=1.3 $Y=1.63 $X2=1.3
+ $Y2=2.31
r150 31 52 2.59952 $w=3.7e-07 $l=3.14325e-07 $layer=LI1_cond $X=1.3 $Y=1.615
+ $X2=1.04 $Y2=1.495
r151 31 33 0.345023 $w=5.18e-07 $l=1.5e-08 $layer=LI1_cond $X=1.3 $Y=1.615
+ $X2=1.3 $Y2=1.63
r152 28 67 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.89 $Y=0.995
+ $X2=3.89 $Y2=1.202
r153 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.89 $Y=0.995
+ $X2=3.89 $Y2=0.56
r154 25 66 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.865 $Y=1.41
+ $X2=3.865 $Y2=1.202
r155 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.865 $Y=1.41
+ $X2=3.865 $Y2=1.985
r156 22 64 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.395 $Y=1.41
+ $X2=3.395 $Y2=1.202
r157 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.395 $Y=1.41
+ $X2=3.395 $Y2=1.985
r158 19 63 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.37 $Y=0.995
+ $X2=3.37 $Y2=1.202
r159 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.37 $Y=0.995
+ $X2=3.37 $Y2=0.56
r160 16 62 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.925 $Y=1.41
+ $X2=2.925 $Y2=1.202
r161 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.925 $Y=1.41
+ $X2=2.925 $Y2=1.985
r162 13 61 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.9 $Y=0.995
+ $X2=2.9 $Y2=1.202
r163 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.9 $Y=0.995
+ $X2=2.9 $Y2=0.56
r164 10 59 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.455 $Y=1.41
+ $X2=2.455 $Y2=1.202
r165 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.455 $Y=1.41
+ $X2=2.455 $Y2=1.985
r166 7 58 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.43 $Y=0.995
+ $X2=2.43 $Y2=1.202
r167 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.43 $Y=0.995
+ $X2=2.43 $Y2=0.56
r168 2 35 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.485 $X2=1.27 $Y2=2.31
r169 2 33 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.485 $X2=1.27 $Y2=1.63
r170 1 41 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=1.545
+ $Y=0.235 $X2=1.68 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_4%VPWR 1 2 3 4 13 15 19 23 27 30 31 33 34 35
+ 37 50 51 57
c59 3 0 1.83248e-19 $X=3.015 $Y=1.485
r60 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r61 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r62 48 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r63 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r64 45 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r65 45 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r66 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r67 42 57 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.345 $Y=2.72
+ $X2=2.205 $Y2=2.72
r68 42 44 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=2.345 $Y=2.72
+ $X2=2.99 $Y2=2.72
r69 41 58 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r70 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r71 38 54 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r72 38 40 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r73 37 57 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=2.205 $Y2=2.72
r74 37 40 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=0.69 $Y2=2.72
r75 35 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r76 35 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r77 33 47 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.975 $Y=2.72
+ $X2=3.91 $Y2=2.72
r78 33 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.975 $Y=2.72
+ $X2=4.1 $Y2=2.72
r79 32 50 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=4.37 $Y2=2.72
r80 32 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=4.1 $Y2=2.72
r81 30 44 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.035 $Y=2.72
+ $X2=2.99 $Y2=2.72
r82 30 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.035 $Y=2.72
+ $X2=3.16 $Y2=2.72
r83 29 47 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.285 $Y=2.72
+ $X2=3.91 $Y2=2.72
r84 29 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.285 $Y=2.72
+ $X2=3.16 $Y2=2.72
r85 25 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.1 $Y=2.635
+ $X2=4.1 $Y2=2.72
r86 25 27 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.1 $Y=2.635 $X2=4.1
+ $Y2=1.96
r87 21 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.16 $Y=2.635
+ $X2=3.16 $Y2=2.72
r88 21 23 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.16 $Y=2.635
+ $X2=3.16 $Y2=2.3
r89 17 57 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.205 $Y=2.635
+ $X2=2.205 $Y2=2.72
r90 17 19 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.205 $Y=2.635
+ $X2=2.205 $Y2=2
r91 13 54 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r92 13 15 15.5919 $w=2.53e-07 $l=3.45e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.29
r93 4 27 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.955
+ $Y=1.485 $X2=4.1 $Y2=1.96
r94 3 23 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.015
+ $Y=1.485 $X2=3.16 $Y2=2.3
r95 2 19 300 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=2 $X=2.005
+ $Y=1.485 $X2=2.215 $Y2=2
r96 1 15 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_4%X 1 2 3 4 15 19 22 23 24 27 31 33 35 39 40
+ 41 44 47
c75 39 0 1.83248e-19 $X=3.08 $Y=1.7
r76 44 47 0.449004 $w=3.83e-07 $l=1.5e-08 $layer=LI1_cond $X=4.297 $Y=1.2
+ $X2=4.297 $Y2=1.185
r77 43 44 7.33373 $w=3.83e-07 $l=2.45e-07 $layer=LI1_cond $X=4.297 $Y=1.445
+ $X2=4.297 $Y2=1.2
r78 42 47 8.3814 $w=3.83e-07 $l=2.8e-07 $layer=LI1_cond $X=4.297 $Y=0.905
+ $X2=4.297 $Y2=1.185
r79 38 40 8.64074 $w=5.08e-07 $l=1.25e-07 $layer=LI1_cond $X=3.63 $Y=1.7
+ $X2=3.755 $Y2=1.7
r80 38 39 18.6081 $w=5.08e-07 $l=5.5e-07 $layer=LI1_cond $X=3.63 $Y=1.7 $X2=3.08
+ $Y2=1.7
r81 36 41 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.795 $Y=0.82
+ $X2=3.605 $Y2=0.82
r82 35 42 8.24022 $w=1.7e-07 $l=2.30617e-07 $layer=LI1_cond $X=4.105 $Y=0.82
+ $X2=4.297 $Y2=0.905
r83 35 36 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.105 $Y=0.82
+ $X2=3.795 $Y2=0.82
r84 33 43 8.24022 $w=1.7e-07 $l=2.30617e-07 $layer=LI1_cond $X=4.105 $Y=1.53
+ $X2=4.297 $Y2=1.445
r85 33 40 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.105 $Y=1.53
+ $X2=3.755 $Y2=1.53
r86 29 38 4.91917 $w=2.5e-07 $l=2.55e-07 $layer=LI1_cond $X=3.63 $Y=1.955
+ $X2=3.63 $Y2=1.7
r87 29 31 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=3.63 $Y=1.955
+ $X2=3.63 $Y2=1.96
r88 25 41 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.605 $Y=0.735
+ $X2=3.605 $Y2=0.82
r89 25 27 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.605 $Y=0.735
+ $X2=3.605 $Y2=0.4
r90 23 41 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.415 $Y=0.82
+ $X2=3.605 $Y2=0.82
r91 23 24 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.415 $Y=0.82
+ $X2=2.855 $Y2=0.82
r92 22 39 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.815 $Y=1.87
+ $X2=3.08 $Y2=1.87
r93 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.69 $Y=1.955
+ $X2=2.815 $Y2=1.87
r94 17 19 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=2.69 $Y=1.955
+ $X2=2.69 $Y2=1.96
r95 13 24 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=2.665 $Y=0.735
+ $X2=2.855 $Y2=0.82
r96 13 15 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.665 $Y=0.735
+ $X2=2.665 $Y2=0.4
r97 4 38 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.485
+ $Y=1.485 $X2=3.63 $Y2=1.62
r98 4 31 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.485
+ $Y=1.485 $X2=3.63 $Y2=1.96
r99 3 19 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.545
+ $Y=1.485 $X2=2.69 $Y2=1.96
r100 2 27 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=3.445
+ $Y=0.235 $X2=3.63 $Y2=0.4
r101 1 15 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=2.505
+ $Y=0.235 $X2=2.69 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_4%VGND 1 2 3 4 17 21 25 28 29 31 32 34 35 36
+ 49 50 53 63
r67 62 63 9.00983 $w=6.48e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.24
+ $X2=1.295 $Y2=0.24
r68 59 62 1.10407 $w=6.48e-07 $l=6e-08 $layer=LI1_cond $X=1.15 $Y=0.24 $X2=1.21
+ $Y2=0.24
r69 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r70 57 59 7.72851 $w=6.48e-07 $l=4.2e-07 $layer=LI1_cond $X=0.73 $Y=0.24
+ $X2=1.15 $Y2=0.24
r71 54 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r72 53 57 0.736048 $w=6.48e-07 $l=4e-08 $layer=LI1_cond $X=0.69 $Y=0.24 $X2=0.73
+ $Y2=0.24
r73 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r74 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r75 47 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r76 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r77 44 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r78 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r79 41 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r80 41 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r81 40 63 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.295
+ $Y2=0
r82 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r83 36 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r84 34 46 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.015 $Y=0 $X2=3.91
+ $Y2=0
r85 34 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.015 $Y=0 $X2=4.1
+ $Y2=0
r86 33 49 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.185 $Y=0 $X2=4.37
+ $Y2=0
r87 33 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.185 $Y=0 $X2=4.1
+ $Y2=0
r88 31 43 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=0 $X2=2.99
+ $Y2=0
r89 31 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=0 $X2=3.16
+ $Y2=0
r90 30 46 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.245 $Y=0 $X2=3.91
+ $Y2=0
r91 30 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.245 $Y=0 $X2=3.16
+ $Y2=0
r92 28 40 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.13 $Y=0 $X2=2.07
+ $Y2=0
r93 28 29 5.29182 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=2.13 $Y=0 $X2=2.217
+ $Y2=0
r94 27 43 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.99
+ $Y2=0
r95 27 29 5.29182 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.217
+ $Y2=0
r96 23 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.1 $Y=0.085 $X2=4.1
+ $Y2=0
r97 23 25 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.1 $Y=0.085 $X2=4.1
+ $Y2=0.385
r98 19 32 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.16 $Y=0.085
+ $X2=3.16 $Y2=0
r99 19 21 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.16 $Y=0.085 $X2=3.16
+ $Y2=0.385
r100 15 29 1.23839 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.217 $Y=0.085
+ $X2=2.217 $Y2=0
r101 15 17 19.9636 $w=1.73e-07 $l=3.15e-07 $layer=LI1_cond $X=2.217 $Y=0.085
+ $X2=2.217 $Y2=0.4
r102 4 25 182 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=1 $X=3.965
+ $Y=0.235 $X2=4.1 $Y2=0.385
r103 3 21 182 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_NDIFF $count=1 $X=2.975
+ $Y=0.235 $X2=3.16 $Y2=0.385
r104 2 17 91 $w=1.7e-07 $l=3.27261e-07 $layer=licon1_NDIFF $count=2 $X=1.965
+ $Y=0.235 $X2=2.22 $Y2=0.4
r105 1 62 182 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.265 $X2=1.21 $Y2=0.4
r106 1 57 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.265 $X2=0.73 $Y2=0.4
.ends

