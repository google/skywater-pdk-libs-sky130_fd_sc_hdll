* File: sky130_fd_sc_hdll__xnor2_1.pxi.spice
* Created: Wed Sep  2 08:53:36 2020
* 
x_PM_SKY130_FD_SC_HDLL__XNOR2_1%B N_B_c_54_n N_B_M1008_g N_B_c_55_n N_B_M1002_g
+ N_B_c_56_n N_B_M1000_g N_B_c_57_n N_B_M1006_g N_B_c_64_n N_B_c_58_n N_B_c_59_n
+ N_B_c_60_n B N_B_c_61_n PM_SKY130_FD_SC_HDLL__XNOR2_1%B
x_PM_SKY130_FD_SC_HDLL__XNOR2_1%A N_A_c_137_n N_A_M1007_g N_A_c_140_n
+ N_A_M1003_g N_A_c_138_n N_A_M1004_g N_A_c_141_n N_A_M1001_g A N_A_c_139_n
+ N_A_c_156_n A PM_SKY130_FD_SC_HDLL__XNOR2_1%A
x_PM_SKY130_FD_SC_HDLL__XNOR2_1%A_47_47# N_A_47_47#_M1002_s N_A_47_47#_M1008_d
+ N_A_47_47#_c_186_n N_A_47_47#_M1009_g N_A_47_47#_c_187_n N_A_47_47#_M1005_g
+ N_A_47_47#_c_188_n N_A_47_47#_c_206_n N_A_47_47#_c_193_n N_A_47_47#_c_208_n
+ N_A_47_47#_c_209_n N_A_47_47#_c_212_n N_A_47_47#_c_194_n N_A_47_47#_c_195_n
+ N_A_47_47#_c_189_n N_A_47_47#_c_190_n N_A_47_47#_c_225_n
+ PM_SKY130_FD_SC_HDLL__XNOR2_1%A_47_47#
x_PM_SKY130_FD_SC_HDLL__XNOR2_1%VPWR N_VPWR_M1008_s N_VPWR_M1003_d
+ N_VPWR_M1009_d N_VPWR_c_283_n N_VPWR_c_284_n N_VPWR_c_285_n N_VPWR_c_286_n
+ VPWR N_VPWR_c_287_n N_VPWR_c_288_n N_VPWR_c_289_n N_VPWR_c_282_n
+ PM_SKY130_FD_SC_HDLL__XNOR2_1%VPWR
x_PM_SKY130_FD_SC_HDLL__XNOR2_1%Y N_Y_M1005_d N_Y_M1000_d N_Y_c_340_n
+ N_Y_c_337_n N_Y_c_350_n N_Y_c_341_n N_Y_c_338_n Y N_Y_c_358_n Y
+ PM_SKY130_FD_SC_HDLL__XNOR2_1%Y
x_PM_SKY130_FD_SC_HDLL__XNOR2_1%VGND N_VGND_M1007_d N_VGND_M1006_s
+ N_VGND_c_375_n N_VGND_c_376_n N_VGND_c_377_n N_VGND_c_378_n N_VGND_c_379_n
+ VGND N_VGND_c_380_n N_VGND_c_381_n PM_SKY130_FD_SC_HDLL__XNOR2_1%VGND
x_PM_SKY130_FD_SC_HDLL__XNOR2_1%A_315_47# N_A_315_47#_M1004_d
+ N_A_315_47#_M1006_d N_A_315_47#_c_421_n N_A_315_47#_c_422_n
+ N_A_315_47#_c_423_n N_A_315_47#_c_451_n
+ PM_SKY130_FD_SC_HDLL__XNOR2_1%A_315_47#
cc_1 VNB N_B_c_54_n 0.0255925f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.41
cc_2 VNB N_B_c_55_n 0.0191259f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=0.995
cc_3 VNB N_B_c_56_n 0.0230879f $X=-0.19 $Y=-0.24 $X2=2.395 $Y2=1.41
cc_4 VNB N_B_c_57_n 0.0217877f $X=-0.19 $Y=-0.24 $X2=2.54 $Y2=0.995
cc_5 VNB N_B_c_58_n 5.70308e-19 $X=-0.19 $Y=-0.24 $X2=2.055 $Y2=1.445
cc_6 VNB N_B_c_59_n 8.63483e-19 $X=-0.19 $Y=-0.24 $X2=2.165 $Y2=1.16
cc_7 VNB N_B_c_60_n 0.00504383f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=1.16
cc_8 VNB N_B_c_61_n 0.00801549f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_9 VNB N_A_c_137_n 0.0165656f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.41
cc_10 VNB N_A_c_138_n 0.0228986f $X=-0.19 $Y=-0.24 $X2=2.395 $Y2=1.41
cc_11 VNB N_A_c_139_n 0.0654623f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=1.16
cc_12 VNB N_A_47_47#_c_186_n 0.029185f $X=-0.19 $Y=-0.24 $X2=2.395 $Y2=1.41
cc_13 VNB N_A_47_47#_c_187_n 0.0201451f $X=-0.19 $Y=-0.24 $X2=2.54 $Y2=0.995
cc_14 VNB N_A_47_47#_c_188_n 0.022254f $X=-0.19 $Y=-0.24 $X2=0.81 $Y2=1.53
cc_15 VNB N_A_47_47#_c_189_n 0.00213909f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_47_47#_c_190_n 0.0253194f $X=-0.19 $Y=-0.24 $X2=0.617 $Y2=1.53
cc_17 VNB N_VPWR_c_282_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Y_c_337_n 0.0253256f $X=-0.19 $Y=-0.24 $X2=2.54 $Y2=0.995
cc_19 VNB N_Y_c_338_n 0.024449f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=1.16
cc_20 VNB N_VGND_c_375_n 0.00613291f $X=-0.19 $Y=-0.24 $X2=2.395 $Y2=1.985
cc_21 VNB N_VGND_c_376_n 0.0347342f $X=-0.19 $Y=-0.24 $X2=2.54 $Y2=0.56
cc_22 VNB N_VGND_c_377_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=1.945 $Y2=1.53
cc_23 VNB N_VGND_c_378_n 0.0128031f $X=-0.19 $Y=-0.24 $X2=0.81 $Y2=1.53
cc_24 VNB N_VGND_c_379_n 0.0198204f $X=-0.19 $Y=-0.24 $X2=2.055 $Y2=1.245
cc_25 VNB N_VGND_c_380_n 0.0326411f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_381_n 0.204723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_315_47#_c_421_n 0.00541433f $X=-0.19 $Y=-0.24 $X2=2.395 $Y2=1.985
cc_28 VNB N_A_315_47#_c_422_n 0.00747803f $X=-0.19 $Y=-0.24 $X2=2.54 $Y2=0.56
cc_29 VNB N_A_315_47#_c_423_n 6.36702e-19 $X=-0.19 $Y=-0.24 $X2=2.54 $Y2=0.56
cc_30 VPB N_B_c_54_n 0.0300443f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=1.41
cc_31 VPB N_B_c_56_n 0.0259166f $X=-0.19 $Y=1.305 $X2=2.395 $Y2=1.41
cc_32 VPB N_B_c_64_n 0.00919532f $X=-0.19 $Y=1.305 $X2=1.945 $Y2=1.53
cc_33 VPB N_B_c_58_n 0.00123012f $X=-0.19 $Y=1.305 $X2=2.055 $Y2=1.445
cc_34 VPB B 3.66229e-19 $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.445
cc_35 VPB N_B_c_61_n 0.00252492f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_36 VPB N_A_c_140_n 0.0201924f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=0.995
cc_37 VPB N_A_c_141_n 0.0194477f $X=-0.19 $Y=1.305 $X2=2.54 $Y2=0.995
cc_38 VPB N_A_c_139_n 0.0372919f $X=-0.19 $Y=1.305 $X2=2.43 $Y2=1.16
cc_39 VPB N_A_47_47#_c_186_n 0.0312229f $X=-0.19 $Y=1.305 $X2=2.395 $Y2=1.41
cc_40 VPB N_A_47_47#_c_188_n 0.0191416f $X=-0.19 $Y=1.305 $X2=0.81 $Y2=1.53
cc_41 VPB N_A_47_47#_c_193_n 0.00766781f $X=-0.19 $Y=1.305 $X2=2.055 $Y2=1.445
cc_42 VPB N_A_47_47#_c_194_n 0.00431297f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=1.16
cc_43 VPB N_A_47_47#_c_195_n 4.15035e-19 $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_44 VPB N_A_47_47#_c_189_n 9.61643e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_283_n 0.0106536f $X=-0.19 $Y=1.305 $X2=2.54 $Y2=0.995
cc_46 VPB N_VPWR_c_284_n 0.019684f $X=-0.19 $Y=1.305 $X2=2.54 $Y2=0.56
cc_47 VPB N_VPWR_c_285_n 0.0157698f $X=-0.19 $Y=1.305 $X2=0.81 $Y2=1.53
cc_48 VPB N_VPWR_c_286_n 0.0192743f $X=-0.19 $Y=1.305 $X2=2.055 $Y2=1.445
cc_49 VPB N_VPWR_c_287_n 0.0381054f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=1.16
cc_50 VPB N_VPWR_c_288_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_289_n 0.020711f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_282_n 0.044649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_Y_c_337_n 0.0338203f $X=-0.19 $Y=1.305 $X2=2.54 $Y2=0.995
cc_54 N_B_c_55_n N_A_c_137_n 0.0378292f $X=0.62 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_55 N_B_c_54_n N_A_c_140_n 0.0220848f $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_56 N_B_c_64_n N_A_c_140_n 0.0158512f $X=1.945 $Y=1.53 $X2=0 $Y2=0
cc_57 N_B_c_61_n N_A_c_140_n 9.02456e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_58 N_B_c_56_n N_A_c_141_n 0.0689351f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_59 N_B_c_64_n N_A_c_141_n 0.0114263f $X=1.945 $Y=1.53 $X2=0 $Y2=0
cc_60 N_B_c_58_n N_A_c_141_n 0.00179613f $X=2.055 $Y=1.445 $X2=0 $Y2=0
cc_61 N_B_c_54_n N_A_c_139_n 0.0414856f $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_62 N_B_c_56_n N_A_c_139_n 0.0274605f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_63 N_B_c_64_n N_A_c_139_n 0.0213795f $X=1.945 $Y=1.53 $X2=0 $Y2=0
cc_64 N_B_c_58_n N_A_c_139_n 0.00891934f $X=2.055 $Y=1.445 $X2=0 $Y2=0
cc_65 N_B_c_59_n N_A_c_139_n 0.00751709f $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_66 N_B_c_61_n N_A_c_139_n 0.00728712f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_67 N_B_c_64_n N_A_c_156_n 0.0571101f $X=1.945 $Y=1.53 $X2=0 $Y2=0
cc_68 N_B_c_58_n N_A_c_156_n 0.00221359f $X=2.055 $Y=1.445 $X2=0 $Y2=0
cc_69 N_B_c_59_n N_A_c_156_n 0.0143374f $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_70 N_B_c_61_n N_A_c_156_n 0.0168087f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_71 N_B_c_64_n N_A_47_47#_M1008_d 4.99619e-19 $X=1.945 $Y=1.53 $X2=0 $Y2=0
cc_72 B N_A_47_47#_M1008_d 0.00140146f $X=0.62 $Y=1.445 $X2=0 $Y2=0
cc_73 N_B_c_56_n N_A_47_47#_c_186_n 0.0578847f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_74 N_B_c_60_n N_A_47_47#_c_186_n 0.00116306f $X=2.43 $Y=1.16 $X2=0 $Y2=0
cc_75 N_B_c_57_n N_A_47_47#_c_187_n 0.0195811f $X=2.54 $Y=0.995 $X2=0 $Y2=0
cc_76 N_B_c_54_n N_A_47_47#_c_188_n 0.0155717f $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_77 N_B_c_55_n N_A_47_47#_c_188_n 0.00419745f $X=0.62 $Y=0.995 $X2=0 $Y2=0
cc_78 B N_A_47_47#_c_188_n 0.008073f $X=0.62 $Y=1.445 $X2=0 $Y2=0
cc_79 N_B_c_61_n N_A_47_47#_c_188_n 0.0346833f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_80 N_B_c_54_n N_A_47_47#_c_206_n 0.0100529f $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_81 B N_A_47_47#_c_206_n 0.00828055f $X=0.62 $Y=1.445 $X2=0 $Y2=0
cc_82 N_B_c_54_n N_A_47_47#_c_208_n 0.0136353f $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_83 N_B_c_56_n N_A_47_47#_c_209_n 0.0107681f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_84 N_B_c_64_n N_A_47_47#_c_209_n 0.0763009f $X=1.945 $Y=1.53 $X2=0 $Y2=0
cc_85 N_B_c_60_n N_A_47_47#_c_209_n 0.00436385f $X=2.43 $Y=1.16 $X2=0 $Y2=0
cc_86 N_B_c_56_n N_A_47_47#_c_212_n 0.00646571f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_87 N_B_c_64_n N_A_47_47#_c_212_n 0.0023738f $X=1.945 $Y=1.53 $X2=0 $Y2=0
cc_88 N_B_c_56_n N_A_47_47#_c_194_n 0.00173414f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_89 N_B_c_60_n N_A_47_47#_c_194_n 0.00651241f $X=2.43 $Y=1.16 $X2=0 $Y2=0
cc_90 N_B_c_56_n N_A_47_47#_c_195_n 0.00991543f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_91 N_B_c_64_n N_A_47_47#_c_195_n 0.0123064f $X=1.945 $Y=1.53 $X2=0 $Y2=0
cc_92 N_B_c_58_n N_A_47_47#_c_195_n 0.00240338f $X=2.055 $Y=1.445 $X2=0 $Y2=0
cc_93 N_B_c_60_n N_A_47_47#_c_195_n 0.0167445f $X=2.43 $Y=1.16 $X2=0 $Y2=0
cc_94 N_B_c_56_n N_A_47_47#_c_189_n 0.00171718f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_95 N_B_c_60_n N_A_47_47#_c_189_n 0.0110294f $X=2.43 $Y=1.16 $X2=0 $Y2=0
cc_96 N_B_c_54_n N_A_47_47#_c_190_n 0.00293839f $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_97 N_B_c_55_n N_A_47_47#_c_190_n 0.00917823f $X=0.62 $Y=0.995 $X2=0 $Y2=0
cc_98 N_B_c_61_n N_A_47_47#_c_190_n 0.00796078f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_99 N_B_c_54_n N_A_47_47#_c_225_n 0.00225422f $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_100 N_B_c_64_n N_A_47_47#_c_225_n 0.00535012f $X=1.945 $Y=1.53 $X2=0 $Y2=0
cc_101 B N_A_47_47#_c_225_n 0.0173047f $X=0.62 $Y=1.445 $X2=0 $Y2=0
cc_102 N_B_c_64_n N_VPWR_M1003_d 0.0103878f $X=1.945 $Y=1.53 $X2=0 $Y2=0
cc_103 N_B_c_54_n N_VPWR_c_284_n 0.0063674f $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_104 N_B_c_56_n N_VPWR_c_287_n 0.00702461f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_105 N_B_c_54_n N_VPWR_c_288_n 0.00597712f $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_106 N_B_c_54_n N_VPWR_c_282_n 0.0075679f $X=0.535 $Y=1.41 $X2=0 $Y2=0
cc_107 N_B_c_56_n N_VPWR_c_282_n 0.0072605f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_108 N_B_c_64_n A_415_297# 0.00147486f $X=1.945 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_109 N_B_c_56_n N_Y_c_340_n 0.00334902f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_110 N_B_c_56_n N_Y_c_341_n 7.14003e-19 $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_111 N_B_c_55_n N_VGND_c_376_n 0.0057945f $X=0.62 $Y=0.995 $X2=0 $Y2=0
cc_112 N_B_c_57_n N_VGND_c_378_n 0.00923235f $X=2.54 $Y=0.995 $X2=0 $Y2=0
cc_113 N_B_c_57_n N_VGND_c_380_n 0.00342417f $X=2.54 $Y=0.995 $X2=0 $Y2=0
cc_114 N_B_c_55_n N_VGND_c_381_n 0.0115332f $X=0.62 $Y=0.995 $X2=0 $Y2=0
cc_115 N_B_c_57_n N_VGND_c_381_n 0.00417726f $X=2.54 $Y=0.995 $X2=0 $Y2=0
cc_116 N_B_c_57_n N_A_315_47#_c_421_n 0.00317826f $X=2.54 $Y=0.995 $X2=0 $Y2=0
cc_117 N_B_c_56_n N_A_315_47#_c_422_n 0.00443205f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_118 N_B_c_57_n N_A_315_47#_c_422_n 0.0129248f $X=2.54 $Y=0.995 $X2=0 $Y2=0
cc_119 N_B_c_64_n N_A_315_47#_c_422_n 0.0019096f $X=1.945 $Y=1.53 $X2=0 $Y2=0
cc_120 N_B_c_59_n N_A_315_47#_c_422_n 0.0132597f $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_121 N_B_c_60_n N_A_315_47#_c_422_n 0.0229216f $X=2.43 $Y=1.16 $X2=0 $Y2=0
cc_122 N_B_c_64_n N_A_315_47#_c_423_n 0.00321907f $X=1.945 $Y=1.53 $X2=0 $Y2=0
cc_123 N_A_c_140_n N_A_47_47#_c_208_n 0.0118097f $X=1.005 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A_c_140_n N_A_47_47#_c_209_n 0.0122434f $X=1.005 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A_c_141_n N_A_47_47#_c_209_n 0.0149524f $X=1.985 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A_c_141_n N_A_47_47#_c_212_n 0.00108532f $X=1.985 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A_c_137_n N_A_47_47#_c_190_n 0.00152741f $X=0.98 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A_c_140_n N_A_47_47#_c_225_n 5.65079e-19 $X=1.005 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_c_141_n N_VPWR_c_287_n 0.00702461f $X=1.985 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_c_140_n N_VPWR_c_288_n 0.00673617f $X=1.005 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A_c_140_n N_VPWR_c_289_n 0.00685571f $X=1.005 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A_c_141_n N_VPWR_c_289_n 0.0118832f $X=1.985 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A_c_140_n N_VPWR_c_282_n 0.00821261f $X=1.005 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_c_141_n N_VPWR_c_282_n 0.00823077f $X=1.985 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_c_137_n N_VGND_c_375_n 0.00904649f $X=0.98 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_c_138_n N_VGND_c_375_n 0.00592912f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_c_139_n N_VGND_c_375_n 0.00431355f $X=1.535 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_c_156_n N_VGND_c_375_n 0.0136981f $X=1.535 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A_c_137_n N_VGND_c_376_n 0.00585385f $X=0.98 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_c_138_n N_VGND_c_378_n 0.00226905f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_c_138_n N_VGND_c_379_n 0.00465454f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_c_137_n N_VGND_c_381_n 0.0108435f $X=0.98 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A_c_138_n N_VGND_c_381_n 0.00934344f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_c_138_n N_A_315_47#_c_421_n 0.00622515f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A_c_139_n N_A_315_47#_c_422_n 0.00587625f $X=1.535 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A_c_138_n N_A_315_47#_c_423_n 0.0037554f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_c_139_n N_A_315_47#_c_423_n 0.00755011f $X=1.535 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_c_156_n N_A_315_47#_c_423_n 0.0142478f $X=1.535 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_47_47#_c_188_n N_VPWR_M1008_s 0.00503262f $X=0.17 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_150 N_A_47_47#_c_206_n N_VPWR_M1008_s 0.0061513f $X=0.555 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_151 N_A_47_47#_c_193_n N_VPWR_M1008_s 0.00242f $X=0.255 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_152 N_A_47_47#_c_209_n N_VPWR_M1003_d 0.0176062f $X=2.335 $Y=1.87 $X2=0 $Y2=0
cc_153 N_A_47_47#_c_194_n N_VPWR_M1009_d 0.00158813f $X=2.875 $Y=1.5 $X2=0 $Y2=0
cc_154 N_A_47_47#_c_206_n N_VPWR_c_284_n 0.0101619f $X=0.555 $Y=1.87 $X2=0 $Y2=0
cc_155 N_A_47_47#_c_193_n N_VPWR_c_284_n 0.0148845f $X=0.255 $Y=1.87 $X2=0 $Y2=0
cc_156 N_A_47_47#_c_208_n N_VPWR_c_284_n 0.0264782f $X=0.77 $Y=1.96 $X2=0 $Y2=0
cc_157 N_A_47_47#_c_186_n N_VPWR_c_286_n 0.00885685f $X=2.925 $Y=1.41 $X2=0
+ $Y2=0
cc_158 N_A_47_47#_c_186_n N_VPWR_c_287_n 0.00624655f $X=2.925 $Y=1.41 $X2=0
+ $Y2=0
cc_159 N_A_47_47#_c_208_n N_VPWR_c_288_n 0.0223557f $X=0.77 $Y=1.96 $X2=0 $Y2=0
cc_160 N_A_47_47#_c_208_n N_VPWR_c_289_n 0.0231743f $X=0.77 $Y=1.96 $X2=0 $Y2=0
cc_161 N_A_47_47#_c_209_n N_VPWR_c_289_n 0.0534723f $X=2.335 $Y=1.87 $X2=0 $Y2=0
cc_162 N_A_47_47#_M1008_d N_VPWR_c_282_n 0.00231261f $X=0.625 $Y=1.485 $X2=0
+ $Y2=0
cc_163 N_A_47_47#_c_186_n N_VPWR_c_282_n 0.00810898f $X=2.925 $Y=1.41 $X2=0
+ $Y2=0
cc_164 N_A_47_47#_c_206_n N_VPWR_c_282_n 0.0058815f $X=0.555 $Y=1.87 $X2=0 $Y2=0
cc_165 N_A_47_47#_c_193_n N_VPWR_c_282_n 6.8277e-19 $X=0.255 $Y=1.87 $X2=0 $Y2=0
cc_166 N_A_47_47#_c_208_n N_VPWR_c_282_n 0.0140101f $X=0.77 $Y=1.96 $X2=0 $Y2=0
cc_167 N_A_47_47#_c_209_n N_VPWR_c_282_n 0.0323404f $X=2.335 $Y=1.87 $X2=0 $Y2=0
cc_168 N_A_47_47#_c_209_n A_415_297# 0.00410382f $X=2.335 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_169 N_A_47_47#_c_209_n N_Y_M1000_d 0.00168082f $X=2.335 $Y=1.87 $X2=0 $Y2=0
cc_170 N_A_47_47#_c_212_n N_Y_M1000_d 0.00245781f $X=2.445 $Y=1.785 $X2=0 $Y2=0
cc_171 N_A_47_47#_c_194_n N_Y_M1000_d 0.00374406f $X=2.875 $Y=1.5 $X2=0 $Y2=0
cc_172 N_A_47_47#_c_186_n N_Y_c_340_n 0.00816929f $X=2.925 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_47_47#_c_186_n N_Y_c_337_n 0.014057f $X=2.925 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_47_47#_c_187_n N_Y_c_337_n 0.00543279f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A_47_47#_c_194_n N_Y_c_337_n 0.0105787f $X=2.875 $Y=1.5 $X2=0 $Y2=0
cc_176 N_A_47_47#_c_189_n N_Y_c_337_n 0.0232673f $X=2.96 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_47_47#_c_186_n N_Y_c_350_n 0.00365702f $X=2.925 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A_47_47#_c_209_n N_Y_c_350_n 0.00100206f $X=2.335 $Y=1.87 $X2=0 $Y2=0
cc_179 N_A_47_47#_c_194_n N_Y_c_350_n 0.0052308f $X=2.875 $Y=1.5 $X2=0 $Y2=0
cc_180 N_A_47_47#_c_186_n N_Y_c_341_n 0.00352866f $X=2.925 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_47_47#_c_209_n N_Y_c_341_n 0.0153272f $X=2.335 $Y=1.87 $X2=0 $Y2=0
cc_182 N_A_47_47#_c_212_n N_Y_c_341_n 0.00244591f $X=2.445 $Y=1.785 $X2=0 $Y2=0
cc_183 N_A_47_47#_c_194_n N_Y_c_341_n 0.00853686f $X=2.875 $Y=1.5 $X2=0 $Y2=0
cc_184 N_A_47_47#_c_187_n N_Y_c_338_n 0.0040016f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_47_47#_c_186_n N_Y_c_358_n 0.0127661f $X=2.925 $Y=1.41 $X2=0 $Y2=0
cc_186 N_A_47_47#_c_194_n N_Y_c_358_n 0.0109729f $X=2.875 $Y=1.5 $X2=0 $Y2=0
cc_187 N_A_47_47#_c_190_n N_VGND_c_375_n 0.0151223f $X=0.36 $Y=0.39 $X2=0 $Y2=0
cc_188 N_A_47_47#_c_190_n N_VGND_c_376_n 0.026295f $X=0.36 $Y=0.39 $X2=0 $Y2=0
cc_189 N_A_47_47#_c_187_n N_VGND_c_378_n 0.0011396f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_47_47#_c_187_n N_VGND_c_380_n 0.00585385f $X=3.01 $Y=0.995 $X2=0
+ $Y2=0
cc_191 N_A_47_47#_M1002_s N_VGND_c_381_n 0.00251629f $X=0.235 $Y=0.235 $X2=0
+ $Y2=0
cc_192 N_A_47_47#_c_187_n N_VGND_c_381_n 0.0121034f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_47_47#_c_190_n N_VGND_c_381_n 0.0174561f $X=0.36 $Y=0.39 $X2=0 $Y2=0
cc_194 N_A_47_47#_c_186_n N_A_315_47#_c_422_n 0.00175161f $X=2.925 $Y=1.41 $X2=0
+ $Y2=0
cc_195 N_A_47_47#_c_194_n N_A_315_47#_c_422_n 0.0066596f $X=2.875 $Y=1.5 $X2=0
+ $Y2=0
cc_196 N_A_47_47#_c_189_n N_A_315_47#_c_422_n 8.74825e-19 $X=2.96 $Y=1.16 $X2=0
+ $Y2=0
cc_197 N_VPWR_c_282_n A_415_297# 0.00312774f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_198 N_VPWR_c_282_n N_Y_M1000_d 0.00329321f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_199 N_VPWR_M1009_d N_Y_c_337_n 0.00449987f $X=3.015 $Y=1.485 $X2=0 $Y2=0
cc_200 N_VPWR_c_285_n N_Y_c_337_n 0.00284759f $X=3.265 $Y=2.635 $X2=0 $Y2=0
cc_201 N_VPWR_c_286_n N_Y_c_337_n 0.00520959f $X=3.2 $Y=2.29 $X2=0 $Y2=0
cc_202 N_VPWR_c_282_n N_Y_c_337_n 0.00519022f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_203 N_VPWR_c_286_n N_Y_c_350_n 0.0107722f $X=3.2 $Y=2.29 $X2=0 $Y2=0
cc_204 N_VPWR_c_287_n N_Y_c_350_n 0.0103369f $X=3.115 $Y=2.72 $X2=0 $Y2=0
cc_205 N_VPWR_c_282_n N_Y_c_350_n 0.0123216f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_206 N_VPWR_M1009_d N_Y_c_358_n 0.0141575f $X=3.015 $Y=1.485 $X2=0 $Y2=0
cc_207 N_VPWR_c_286_n N_Y_c_358_n 0.0190567f $X=3.2 $Y=2.29 $X2=0 $Y2=0
cc_208 N_VPWR_c_282_n N_Y_c_358_n 0.00815801f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_209 N_Y_c_338_n N_VGND_c_380_n 0.0183504f $X=3.475 $Y=0.585 $X2=0 $Y2=0
cc_210 N_Y_M1005_d N_VGND_c_381_n 0.00562368f $X=3.085 $Y=0.235 $X2=0 $Y2=0
cc_211 N_Y_c_338_n N_VGND_c_381_n 0.0152277f $X=3.475 $Y=0.585 $X2=0 $Y2=0
cc_212 A_139_47# N_VGND_c_381_n 0.00897657f $X=0.695 $Y=0.235 $X2=3.45 $Y2=0
cc_213 N_VGND_c_381_n N_A_315_47#_M1004_d 0.00209319f $X=3.45 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_214 N_VGND_c_381_n N_A_315_47#_M1006_d 0.00418178f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_215 N_VGND_c_375_n N_A_315_47#_c_421_n 0.0298239f $X=1.24 $Y=0.39 $X2=0 $Y2=0
cc_216 N_VGND_c_378_n N_A_315_47#_c_421_n 0.0156864f $X=2.295 $Y=0 $X2=0 $Y2=0
cc_217 N_VGND_c_379_n N_A_315_47#_c_421_n 0.0241599f $X=2.095 $Y=0 $X2=0 $Y2=0
cc_218 N_VGND_c_381_n N_A_315_47#_c_421_n 0.0140576f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_219 N_VGND_M1006_s N_A_315_47#_c_422_n 0.00674008f $X=2.155 $Y=0.235 $X2=0
+ $Y2=0
cc_220 N_VGND_c_378_n N_A_315_47#_c_422_n 0.0248804f $X=2.295 $Y=0 $X2=0 $Y2=0
cc_221 N_VGND_c_379_n N_A_315_47#_c_422_n 0.00384718f $X=2.095 $Y=0 $X2=0 $Y2=0
cc_222 N_VGND_c_380_n N_A_315_47#_c_422_n 0.00233324f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_223 N_VGND_c_381_n N_A_315_47#_c_422_n 0.0120675f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_224 N_VGND_c_375_n N_A_315_47#_c_423_n 0.0133617f $X=1.24 $Y=0.39 $X2=0 $Y2=0
cc_225 N_VGND_c_380_n N_A_315_47#_c_451_n 0.0150812f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_226 N_VGND_c_381_n N_A_315_47#_c_451_n 0.00874048f $X=3.45 $Y=0 $X2=0 $Y2=0
