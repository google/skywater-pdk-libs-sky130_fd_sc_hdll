* File: sky130_fd_sc_hdll__o221a_1.pex.spice
* Created: Thu Aug 27 19:20:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O221A_1%C1 1 3 4 6 7 12
c29 4 0 1.69639e-19 $X=0.545 $Y=0.995
r30 12 13 3.31956 $w=3.63e-07 $l=2.5e-08 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.545 $Y2=1.202
r31 10 12 35.8512 $w=3.63e-07 $l=2.7e-07 $layer=POLY_cond $X=0.25 $Y=1.202
+ $X2=0.52 $Y2=1.202
r32 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r33 4 13 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.545 $Y=0.995
+ $X2=0.545 $Y2=1.202
r34 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.545 $Y=0.995
+ $X2=0.545 $Y2=0.56
r35 1 12 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.52 $Y=1.41
+ $X2=0.52 $Y2=1.202
r36 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.52 $Y=1.41 $X2=0.52
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_1%B1 1 3 4 6 7 15
c36 15 0 2.7937e-20 $X=1.09 $Y=1.19
r37 7 15 2.54215 $w=3.38e-07 $l=7.5e-08 $layer=LI1_cond $X=1.015 $Y=1.155
+ $X2=1.09 $Y2=1.155
r38 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.015
+ $Y=1.16 $X2=1.015 $Y2=1.16
r39 4 10 41.1443 $w=2.56e-07 $l=2.02793e-07 $layer=POLY_cond $X=1.075 $Y=0.985
+ $X2=1.015 $Y2=1.16
r40 4 6 136.567 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=1.075 $Y=0.985
+ $X2=1.075 $Y2=0.56
r41 1 10 51.3767 $w=2.56e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.05 $Y=1.41
+ $X2=1.015 $Y2=1.16
r42 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.05 $Y=1.41 $X2=1.05
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_1%B2 1 3 4 6 7 8 18
c34 7 0 2.58934e-20 $X=1.575 $Y=1.19
c35 4 0 7.5851e-20 $X=1.52 $Y=0.995
r36 8 18 0.598672 $w=3.83e-07 $l=2e-08 $layer=LI1_cond $X=1.597 $Y=1.55
+ $X2=1.597 $Y2=1.53
r37 7 18 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=1.597 $Y=1.16
+ $X2=1.597 $Y2=1.53
r38 7 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.495
+ $Y=1.16 $X2=1.495 $Y2=1.16
r39 4 12 39.2931 $w=2.55e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.52 $Y=0.995
+ $X2=1.495 $Y2=1.16
r40 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.52 $Y=0.995 $X2=1.52
+ $Y2=0.56
r41 1 12 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.46 $Y=1.41
+ $X2=1.495 $Y2=1.16
r42 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.46 $Y=1.41 $X2=1.46
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_1%A2 1 3 4 6 9 12 13 18
c38 18 0 4.7914e-20 $X=2.147 $Y=1.255
c39 4 0 2.58934e-20 $X=2.51 $Y=0.995
r40 12 18 3.08287 $w=3.35e-07 $l=1.35e-07 $layer=LI1_cond $X=2.147 $Y=1.12
+ $X2=2.147 $Y2=1.255
r41 12 13 9.11634 $w=3.33e-07 $l=2.65e-07 $layer=LI1_cond $X=2.147 $Y=1.265
+ $X2=2.147 $Y2=1.53
r42 12 18 0.344013 $w=3.33e-07 $l=1e-08 $layer=LI1_cond $X=2.147 $Y=1.265
+ $X2=2.147 $Y2=1.255
r43 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.45
+ $Y=1.16 $X2=2.45 $Y2=1.16
r44 7 12 3.83646 $w=2.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.315 $Y=1.12
+ $X2=2.147 $Y2=1.12
r45 7 9 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.315 $Y=1.12
+ $X2=2.45 $Y2=1.12
r46 4 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.51 $Y=0.995
+ $X2=2.45 $Y2=1.16
r47 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.51 $Y=0.995 $X2=2.51
+ $Y2=0.56
r48 1 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.485 $Y=1.41
+ $X2=2.45 $Y2=1.16
r49 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.485 $Y=1.41
+ $X2=2.485 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_1%A1 1 3 4 6 7 13
c32 1 0 1.64731e-19 $X=2.895 $Y=1.41
r33 7 13 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=2.935 $Y=1.18 $X2=2.93
+ $Y2=1.18
r34 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.98
+ $Y=1.16 $X2=2.98 $Y2=1.16
r35 4 10 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=2.98 $Y=0.995
+ $X2=2.955 $Y2=1.16
r36 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.98 $Y=0.995 $X2=2.98
+ $Y2=0.56
r37 1 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.955 $Y2=1.16
r38 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_1%A_27_297# 1 2 3 10 12 13 15 18 22 25 26 29
+ 31 32 35 36 37 40 48 51 55 56
c116 10 0 1.22937e-19 $X=3.4 $Y=0.995
r117 54 56 8.87457 $w=5.88e-07 $l=1.05e-07 $layer=LI1_cond $X=2.25 $Y=2.17
+ $X2=2.355 $Y2=2.17
r118 54 55 21.9503 $w=5.88e-07 $l=7.5e-07 $layer=LI1_cond $X=2.25 $Y=2.17
+ $X2=1.5 $Y2=2.17
r119 43 46 2.39186 $w=2.63e-07 $l=5.5e-08 $layer=LI1_cond $X=0.225 $Y=1.587
+ $X2=0.28 $Y2=1.587
r120 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.46
+ $Y=1.16 $X2=3.46 $Y2=1.16
r121 38 40 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.46 $Y=1.455
+ $X2=3.46 $Y2=1.16
r122 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.375 $Y=1.54
+ $X2=3.46 $Y2=1.455
r123 36 37 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.375 $Y=1.54
+ $X2=2.745 $Y2=1.54
r124 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.66 $Y=1.625
+ $X2=2.745 $Y2=1.54
r125 34 35 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.66 $Y=1.625
+ $X2=2.66 $Y2=1.875
r126 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.575 $Y=1.96
+ $X2=2.66 $Y2=1.875
r127 32 56 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.575 $Y=1.96
+ $X2=2.355 $Y2=1.96
r128 31 55 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.235 $Y=1.96
+ $X2=1.5 $Y2=1.96
r129 29 31 6.89401 $w=1.7e-07 $l=1.39155e-07 $layer=LI1_cond $X=1.132 $Y=1.875
+ $X2=1.235 $Y2=1.96
r130 28 29 8.38581 $w=2.03e-07 $l=1.55e-07 $layer=LI1_cond $X=1.132 $Y=1.72
+ $X2=1.132 $Y2=1.875
r131 26 28 6.83569 $w=2.25e-07 $l=1.55869e-07 $layer=LI1_cond $X=1.03 $Y=1.607
+ $X2=1.132 $Y2=1.72
r132 26 48 14.0854 $w=2.23e-07 $l=2.75e-07 $layer=LI1_cond $X=1.03 $Y=1.607
+ $X2=0.755 $Y2=1.607
r133 25 48 3.99221 $w=2.63e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=1.587
+ $X2=0.755 $Y2=1.587
r134 25 46 16.9605 $w=2.63e-07 $l=3.9e-07 $layer=LI1_cond $X=0.67 $Y=1.587
+ $X2=0.28 $Y2=1.587
r135 24 51 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=0.67 $Y=0.825 $X2=0.67
+ $Y2=0.735
r136 24 25 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=0.67 $Y=0.825
+ $X2=0.67 $Y2=1.455
r137 20 51 20.6414 $w=1.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.335 $Y=0.735
+ $X2=0.67 $Y2=0.735
r138 20 22 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=0.335 $Y=0.645
+ $X2=0.335 $Y2=0.39
r139 16 43 0.377927 $w=2.8e-07 $l=1.33e-07 $layer=LI1_cond $X=0.225 $Y=1.72
+ $X2=0.225 $Y2=1.587
r140 16 18 9.87808 $w=2.78e-07 $l=2.4e-07 $layer=LI1_cond $X=0.225 $Y=1.72
+ $X2=0.225 $Y2=1.96
r141 13 41 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.425 $Y=1.41
+ $X2=3.46 $Y2=1.16
r142 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.425 $Y=1.41
+ $X2=3.425 $Y2=1.985
r143 10 41 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.4 $Y=0.995
+ $X2=3.46 $Y2=1.16
r144 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.4 $Y=0.995
+ $X2=3.4 $Y2=0.56
r145 3 54 150 $w=1.7e-07 $l=9.06918e-07 $layer=licon1_PDIFF $count=4 $X=1.55
+ $Y=1.485 $X2=2.25 $Y2=1.96
r146 2 46 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r147 2 18 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.96
r148 1 22 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.21
+ $Y=0.235 $X2=0.335 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_1%VPWR 1 2 9 13 15 17 22 29 30 33 36
r52 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r54 30 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=2.99 $Y2=2.72
r55 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r56 27 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.295 $Y=2.72
+ $X2=3.105 $Y2=2.72
r57 27 29 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.295 $Y=2.72
+ $X2=3.91 $Y2=2.72
r58 26 37 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r59 26 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r60 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r61 23 33 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.86 $Y=2.72 $X2=0.71
+ $Y2=2.72
r62 23 25 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.86 $Y=2.72
+ $X2=1.15 $Y2=2.72
r63 22 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=3.105 $Y2=2.72
r64 22 25 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=1.15 $Y2=2.72
r65 17 33 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.56 $Y=2.72 $X2=0.71
+ $Y2=2.72
r66 17 19 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.56 $Y=2.72
+ $X2=0.23 $Y2=2.72
r67 15 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r68 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r69 11 36 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=2.635
+ $X2=3.105 $Y2=2.72
r70 11 13 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=3.105 $Y=2.635
+ $X2=3.105 $Y2=1.96
r71 7 33 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=2.635 $X2=0.71
+ $Y2=2.72
r72 7 9 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=0.71 $Y=2.635
+ $X2=0.71 $Y2=2.3
r73 2 13 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.985
+ $Y=1.485 $X2=3.13 $Y2=1.96
r74 1 9 600 $w=1.7e-07 $l=8.937e-07 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.485 $X2=0.775 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_1%X 1 2 9 12 18
c18 9 0 1.4466e-19 $X=3.66 $Y=0.39
r19 18 20 0.182927 $w=3.13e-07 $l=5e-09 $layer=LI1_cond $X=3.872 $Y=1.87
+ $X2=3.872 $Y2=1.875
r20 12 22 0.952629 $w=5.63e-07 $l=4.5e-08 $layer=LI1_cond $X=3.747 $Y=1.915
+ $X2=3.747 $Y2=1.96
r21 12 20 3.17011 $w=5.63e-07 $l=4e-08 $layer=LI1_cond $X=3.747 $Y=1.915
+ $X2=3.747 $Y2=1.875
r22 12 18 1.46342 $w=3.13e-07 $l=4e-08 $layer=LI1_cond $X=3.872 $Y=1.83
+ $X2=3.872 $Y2=1.87
r23 11 12 36.7684 $w=3.13e-07 $l=1.005e-06 $layer=LI1_cond $X=3.872 $Y=0.825
+ $X2=3.872 $Y2=1.83
r24 9 11 11.4254 $w=5.83e-07 $l=4.35e-07 $layer=LI1_cond $X=3.737 $Y=0.39
+ $X2=3.737 $Y2=0.825
r25 2 22 300 $w=1.7e-07 $l=5.51362e-07 $layer=licon1_PDIFF $count=2 $X=3.515
+ $Y=1.485 $X2=3.68 $Y2=1.96
r26 1 9 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.475
+ $Y=0.235 $X2=3.66 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_1%A_124_47# 1 2 11
r18 8 11 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=0.865 $Y=0.39
+ $X2=1.73 $Y2=0.39
r19 2 11 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.73 $Y2=0.39
r20 1 8 182 $w=1.7e-07 $l=3.1305e-07 $layer=licon1_NDIFF $count=1 $X=0.62
+ $Y=0.235 $X2=0.865 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_1%A_230_47# 1 2 7 11 13
c31 13 0 2.67597e-19 $X=2.77 $Y=0.39
c32 7 0 1.69639e-19 $X=2.605 $Y=0.73
r33 11 16 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.77 $Y=0.645 $X2=2.77
+ $Y2=0.73
r34 11 13 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.77 $Y=0.645
+ $X2=2.77 $Y2=0.39
r35 7 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.605 $Y=0.73
+ $X2=2.77 $Y2=0.73
r36 7 9 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=2.605 $Y=0.73
+ $X2=1.285 $Y2=0.73
r37 2 16 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=2.585
+ $Y=0.235 $X2=2.77 $Y2=0.73
r38 2 13 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.585
+ $Y=0.235 $X2=2.77 $Y2=0.39
r39 1 9 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.15
+ $Y=0.235 $X2=1.285 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221A_1%VGND 1 2 9 13 16 17 19 20 21 34 35
c47 13 0 1.64731e-19 $X=3.19 $Y=0.39
r48 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r49 32 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r50 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r51 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r52 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r53 24 28 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r54 21 29 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r55 21 24 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r56 19 31 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=2.99
+ $Y2=0
r57 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=0 $X2=3.19
+ $Y2=0
r58 18 34 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.275 $Y=0 $X2=3.91
+ $Y2=0
r59 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=0 $X2=3.19
+ $Y2=0
r60 16 28 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.085 $Y=0 $X2=2.07
+ $Y2=0
r61 16 17 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.085 $Y=0 $X2=2.255
+ $Y2=0
r62 15 31 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.99
+ $Y2=0
r63 15 17 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.255
+ $Y2=0
r64 11 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.19 $Y=0.085
+ $X2=3.19 $Y2=0
r65 11 13 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.19 $Y=0.085
+ $X2=3.19 $Y2=0.39
r66 7 17 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=0.085
+ $X2=2.255 $Y2=0
r67 7 9 10.3381 $w=3.38e-07 $l=3.05e-07 $layer=LI1_cond $X=2.255 $Y=0.085
+ $X2=2.255 $Y2=0.39
r68 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.055
+ $Y=0.235 $X2=3.19 $Y2=0.39
r69 1 9 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.125
+ $Y=0.235 $X2=2.25 $Y2=0.39
.ends

