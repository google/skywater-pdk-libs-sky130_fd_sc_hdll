* File: sky130_fd_sc_hdll__or4b_4.pex.spice
* Created: Thu Aug 27 19:25:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR4B_4%D_N 2 3 5 8 9 10 11 16 17 18
c25 17 0 1.9892e-19 $X=0.36 $Y=1.16
r26 16 19 36.6898 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.42 $Y=1.16
+ $X2=0.42 $Y2=1.325
r27 16 18 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.42 $Y=1.16
+ $X2=0.42 $Y2=0.995
r28 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.36
+ $Y=1.16 $X2=0.36 $Y2=1.16
r29 10 11 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.275 $Y=1.53
+ $X2=0.275 $Y2=1.87
r30 9 10 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.275 $Y=1.19
+ $X2=0.275 $Y2=1.53
r31 9 17 1.01686 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=0.275 $Y=1.19 $X2=0.275
+ $Y2=1.16
r32 8 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.52 $Y=0.675
+ $X2=0.52 $Y2=0.995
r33 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r34 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.89 $X2=0.495
+ $Y2=1.99
r35 2 19 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.495 $Y=1.89
+ $X2=0.495 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_4%A_117_413# 1 2 7 9 10 12 13 14 17 21 26
c49 13 0 1.9892e-19 $X=1.385 $Y=1.16
r50 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.18
+ $Y=1.16 $X2=1.18 $Y2=1.16
r51 23 26 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.74 $Y=1.16
+ $X2=1.18 $Y2=1.16
r52 19 23 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.74 $Y=1.325
+ $X2=0.74 $Y2=1.16
r53 19 21 55.4545 $w=1.88e-07 $l=9.5e-07 $layer=LI1_cond $X=0.74 $Y=1.325
+ $X2=0.74 $Y2=2.275
r54 15 23 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.74 $Y=0.995
+ $X2=0.74 $Y2=1.16
r55 15 17 14.8852 $w=1.88e-07 $l=2.55e-07 $layer=LI1_cond $X=0.74 $Y=0.995
+ $X2=0.74 $Y2=0.74
r56 13 27 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.385 $Y=1.16
+ $X2=1.18 $Y2=1.16
r57 13 14 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.385 $Y=1.16
+ $X2=1.485 $Y2=1.202
r58 10 14 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.485 $Y2=1.202
r59 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=0.56
r60 7 14 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.202
r61 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.985
r62 2 21 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.065 $X2=0.73 $Y2=2.275
r63 1 17 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.465 $X2=0.73 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_4%C 1 3 4 6 7 8 13
r33 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.98
+ $Y=1.16 $X2=1.98 $Y2=1.16
r34 7 8 13.5114 $w=2.88e-07 $l=3.4e-07 $layer=LI1_cond $X=2.04 $Y=1.87 $X2=2.04
+ $Y2=2.21
r35 7 13 28.215 $w=2.88e-07 $l=7.1e-07 $layer=LI1_cond $X=2.04 $Y=1.87 $X2=2.04
+ $Y2=1.16
r36 4 12 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.09 $Y=0.995
+ $X2=2.005 $Y2=1.16
r37 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.09 $Y=0.995 $X2=2.09
+ $Y2=0.56
r38 1 12 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.065 $Y=1.41
+ $X2=2.005 $Y2=1.16
r39 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.065 $Y=1.41
+ $X2=2.065 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_4%B 1 3 4 6 7 8 13
c31 1 0 5.72837e-20 $X=2.535 $Y=1.41
r32 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.54
+ $Y=1.16 $X2=2.54 $Y2=1.16
r33 7 8 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.54 $Y=1.87 $X2=2.54
+ $Y2=2.21
r34 7 13 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.54 $Y=1.87 $X2=2.54
+ $Y2=1.16
r35 4 12 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=2.56 $Y=0.995
+ $X2=2.535 $Y2=1.16
r36 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.56 $Y=0.995 $X2=2.56
+ $Y2=0.56
r37 1 12 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=2.535 $Y=1.41
+ $X2=2.535 $Y2=1.16
r38 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.535 $Y=1.41
+ $X2=2.535 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_4%A 1 3 4 6 7 12 18
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.04
+ $Y=1.16 $X2=3.04 $Y2=1.16
r39 7 18 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.025 $Y=1.53
+ $X2=2.99 $Y2=1.53
r40 7 12 10.3241 $w=3.18e-07 $l=2.85e-07 $layer=LI1_cond $X=3.025 $Y=1.445
+ $X2=3.025 $Y2=1.16
r41 4 11 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=3.005 $Y=1.41
+ $X2=3.065 $Y2=1.16
r42 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.005 $Y=1.41
+ $X2=3.005 $Y2=1.985
r43 1 11 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.98 $Y=0.995
+ $X2=3.065 $Y2=1.16
r44 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.98 $Y=0.995 $X2=2.98
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_4%A_225_297# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 36 39 42 44 45 48 50 53 54 59 70 79
c141 70 0 5.72837e-20 $X=2.77 $Y=0.74
c142 50 0 1.60701e-19 $X=3.345 $Y=0.74
r143 79 80 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.995 $Y=1.202
+ $X2=5.02 $Y2=1.202
r144 76 77 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.5 $Y=1.202
+ $X2=4.525 $Y2=1.202
r145 75 76 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=4.055 $Y=1.202
+ $X2=4.5 $Y2=1.202
r146 74 75 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.03 $Y=1.202
+ $X2=4.055 $Y2=1.202
r147 71 72 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.56 $Y=1.202
+ $X2=3.585 $Y2=1.202
r148 60 79 26.5618 $w=3.72e-07 $l=2.05e-07 $layer=POLY_cond $X=4.79 $Y=1.202
+ $X2=4.995 $Y2=1.202
r149 60 77 34.336 $w=3.72e-07 $l=2.65e-07 $layer=POLY_cond $X=4.79 $Y=1.202
+ $X2=4.525 $Y2=1.202
r150 59 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.79
+ $Y=1.16 $X2=4.79 $Y2=1.16
r151 57 74 53.1237 $w=3.72e-07 $l=4.1e-07 $layer=POLY_cond $X=3.62 $Y=1.202
+ $X2=4.03 $Y2=1.202
r152 57 72 4.53495 $w=3.72e-07 $l=3.5e-08 $layer=POLY_cond $X=3.62 $Y=1.202
+ $X2=3.585 $Y2=1.202
r153 56 59 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=3.62 $Y=1.16
+ $X2=4.79 $Y2=1.16
r154 56 57 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.62
+ $Y=1.16 $X2=3.62 $Y2=1.16
r155 54 56 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.515 $Y=1.16
+ $X2=3.62 $Y2=1.16
r156 53 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.43 $Y=1.075
+ $X2=3.515 $Y2=1.16
r157 52 53 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.43 $Y=0.825
+ $X2=3.43 $Y2=1.075
r158 51 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=0.74
+ $X2=2.77 $Y2=0.74
r159 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.345 $Y=0.74
+ $X2=3.43 $Y2=0.825
r160 50 51 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.345 $Y=0.74
+ $X2=2.855 $Y2=0.74
r161 46 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.77 $Y=0.655
+ $X2=2.77 $Y2=0.74
r162 46 48 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.77 $Y=0.655
+ $X2=2.77 $Y2=0.49
r163 45 69 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.885 $Y=0.74
+ $X2=1.8 $Y2=0.74
r164 44 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.685 $Y=0.74
+ $X2=2.77 $Y2=0.74
r165 44 45 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=2.685 $Y=0.74
+ $X2=1.885 $Y2=0.74
r166 40 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.8 $Y=0.655
+ $X2=1.8 $Y2=0.74
r167 40 42 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.8 $Y=0.655
+ $X2=1.8 $Y2=0.49
r168 39 63 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.615 $Y=1.66
+ $X2=1.25 $Y2=1.66
r169 38 69 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.615 $Y=0.74
+ $X2=1.8 $Y2=0.74
r170 38 39 39.2878 $w=2.18e-07 $l=7.5e-07 $layer=LI1_cond $X=1.615 $Y=0.825
+ $X2=1.615 $Y2=1.575
r171 36 63 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=1.25 $Y=2.34
+ $X2=1.25 $Y2=1.745
r172 31 80 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.02 $Y=0.995
+ $X2=5.02 $Y2=1.202
r173 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.02 $Y=0.995
+ $X2=5.02 $Y2=0.56
r174 28 79 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.995 $Y=1.41
+ $X2=4.995 $Y2=1.202
r175 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.995 $Y=1.41
+ $X2=4.995 $Y2=1.985
r176 25 77 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.525 $Y=1.41
+ $X2=4.525 $Y2=1.202
r177 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.525 $Y=1.41
+ $X2=4.525 $Y2=1.985
r178 22 76 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.5 $Y=0.995
+ $X2=4.5 $Y2=1.202
r179 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.5 $Y=0.995
+ $X2=4.5 $Y2=0.56
r180 19 75 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.055 $Y=1.41
+ $X2=4.055 $Y2=1.202
r181 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.055 $Y=1.41
+ $X2=4.055 $Y2=1.985
r182 16 74 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.03 $Y=0.995
+ $X2=4.03 $Y2=1.202
r183 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.03 $Y=0.995
+ $X2=4.03 $Y2=0.56
r184 13 72 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.585 $Y=1.41
+ $X2=3.585 $Y2=1.202
r185 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.585 $Y=1.41
+ $X2=3.585 $Y2=1.985
r186 10 71 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.56 $Y=0.995
+ $X2=3.56 $Y2=1.202
r187 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.56 $Y=0.995
+ $X2=3.56 $Y2=0.56
r188 3 63 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.25 $Y2=1.66
r189 3 36 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.25 $Y2=2.34
r190 2 48 182 $w=1.7e-07 $l=3.15357e-07 $layer=licon1_NDIFF $count=1 $X=2.635
+ $Y=0.235 $X2=2.77 $Y2=0.49
r191 1 42 182 $w=1.7e-07 $l=3.46194e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.235 $X2=1.8 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_4%VPWR 1 2 3 4 13 15 19 23 25 27 30 31 33 34
+ 35 47 56
r65 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r66 50 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r67 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r68 47 55 3.95357 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=5.105 $Y=2.72
+ $X2=5.312 $Y2=2.72
r69 47 49 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.105 $Y=2.72
+ $X2=4.83 $Y2=2.72
r70 46 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r71 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r72 43 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r73 42 43 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r74 40 43 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.99 $Y2=2.72
r75 39 42 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.99 $Y2=2.72
r76 39 40 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r77 37 52 4.33083 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=2.72
+ $X2=0.182 $Y2=2.72
r78 37 39 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=2.72
+ $X2=0.69 $Y2=2.72
r79 35 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r80 35 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r81 33 45 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.165 $Y=2.72
+ $X2=3.91 $Y2=2.72
r82 33 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.165 $Y=2.72
+ $X2=4.29 $Y2=2.72
r83 32 49 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.415 $Y=2.72
+ $X2=4.83 $Y2=2.72
r84 32 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.415 $Y=2.72
+ $X2=4.29 $Y2=2.72
r85 30 42 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.17 $Y=2.72
+ $X2=2.99 $Y2=2.72
r86 30 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.17 $Y=2.72
+ $X2=3.295 $Y2=2.72
r87 29 45 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.42 $Y=2.72
+ $X2=3.91 $Y2=2.72
r88 29 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.42 $Y=2.72
+ $X2=3.295 $Y2=2.72
r89 25 55 3.18959 $w=2.5e-07 $l=1.19143e-07 $layer=LI1_cond $X=5.23 $Y=2.635
+ $X2=5.312 $Y2=2.72
r90 25 27 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.23 $Y=2.635
+ $X2=5.23 $Y2=1.96
r91 21 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.29 $Y=2.635
+ $X2=4.29 $Y2=2.72
r92 21 23 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.29 $Y=2.635
+ $X2=4.29 $Y2=1.96
r93 17 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.295 $Y=2.635
+ $X2=3.295 $Y2=2.72
r94 17 19 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.295 $Y=2.635
+ $X2=3.295 $Y2=1.96
r95 13 52 3.02922 $w=2.8e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.225 $Y=2.635
+ $X2=0.182 $Y2=2.72
r96 13 15 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.225 $Y=2.635
+ $X2=0.225 $Y2=2.3
r97 4 27 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.085
+ $Y=1.485 $X2=5.23 $Y2=1.96
r98 3 23 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.145
+ $Y=1.485 $X2=4.29 $Y2=1.96
r99 2 19 300 $w=1.7e-07 $l=5.66238e-07 $layer=licon1_PDIFF $count=2 $X=3.095
+ $Y=1.485 $X2=3.295 $Y2=1.96
r100 1 15 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_4%X 1 2 3 4 13 15 19 21 23 24 27 31 33 35 39
+ 41 43 46
r79 43 46 2.99957 $w=2.4e-07 $l=9e-08 $layer=LI1_cond $X=5.295 $Y=0.815
+ $X2=5.295 $Y2=0.905
r80 43 46 0.720277 $w=2.38e-07 $l=1.5e-08 $layer=LI1_cond $X=5.295 $Y=0.92
+ $X2=5.295 $Y2=0.905
r81 42 43 25.6899 $w=2.38e-07 $l=5.35e-07 $layer=LI1_cond $X=5.295 $Y=1.455
+ $X2=5.295 $Y2=0.92
r82 36 39 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.925 $Y=0.815
+ $X2=4.735 $Y2=0.815
r83 35 43 3.99943 $w=1.8e-07 $l=1.2e-07 $layer=LI1_cond $X=5.175 $Y=0.815
+ $X2=5.295 $Y2=0.815
r84 35 36 15.404 $w=1.78e-07 $l=2.5e-07 $layer=LI1_cond $X=5.175 $Y=0.815
+ $X2=4.925 $Y2=0.815
r85 34 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.885 $Y=1.54
+ $X2=4.76 $Y2=1.54
r86 33 42 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=5.175 $Y=1.54
+ $X2=5.295 $Y2=1.455
r87 33 34 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.175 $Y=1.54
+ $X2=4.885 $Y2=1.54
r88 29 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.76 $Y=1.625
+ $X2=4.76 $Y2=1.54
r89 29 31 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.76 $Y=1.625
+ $X2=4.76 $Y2=2.3
r90 25 39 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=4.735 $Y=0.725
+ $X2=4.735 $Y2=0.815
r91 25 27 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.735 $Y=0.725
+ $X2=4.735 $Y2=0.39
r92 23 39 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.545 $Y=0.815
+ $X2=4.735 $Y2=0.815
r93 23 24 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.545 $Y=0.815
+ $X2=3.985 $Y2=0.815
r94 22 38 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.945 $Y=1.54
+ $X2=3.82 $Y2=1.54
r95 21 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.635 $Y=1.54
+ $X2=4.76 $Y2=1.54
r96 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.635 $Y=1.54
+ $X2=3.945 $Y2=1.54
r97 17 24 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=3.86 $Y=0.725
+ $X2=3.985 $Y2=0.815
r98 17 19 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=3.86 $Y=0.725
+ $X2=3.86 $Y2=0.485
r99 13 38 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.82 $Y=1.625
+ $X2=3.82 $Y2=1.54
r100 13 15 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.82 $Y=1.625
+ $X2=3.82 $Y2=2.3
r101 4 41 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.615
+ $Y=1.485 $X2=4.76 $Y2=1.62
r102 4 31 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.615
+ $Y=1.485 $X2=4.76 $Y2=2.3
r103 3 38 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.675
+ $Y=1.485 $X2=3.82 $Y2=1.62
r104 3 15 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.675
+ $Y=1.485 $X2=3.82 $Y2=2.3
r105 2 27 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.575
+ $Y=0.235 $X2=4.76 $Y2=0.39
r106 1 19 182 $w=1.7e-07 $l=3.29773e-07 $layer=licon1_NDIFF $count=1 $X=3.635
+ $Y=0.235 $X2=3.82 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_4%VGND 1 2 3 4 5 6 19 21 23 27 31 35 39 41 43
+ 46 47 49 50 52 53 54 66 74 78
c96 52 0 1.60701e-19 $X=4.205 $Y=0
r97 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r98 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r99 69 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r100 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r101 66 77 3.40825 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=5.145 $Y=0
+ $X2=5.332 $Y2=0
r102 66 68 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.145 $Y=0
+ $X2=4.83 $Y2=0
r103 65 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r104 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r105 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r106 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r107 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r108 59 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r109 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r110 56 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.21
+ $Y2=0
r111 56 58 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.335 $Y=0
+ $X2=2.07 $Y2=0
r112 54 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r113 54 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r114 52 64 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.205 $Y=0 $X2=3.91
+ $Y2=0
r115 52 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.205 $Y=0 $X2=4.29
+ $Y2=0
r116 51 68 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=4.375 $Y=0
+ $X2=4.83 $Y2=0
r117 51 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.375 $Y=0 $X2=4.29
+ $Y2=0
r118 49 61 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.125 $Y=0
+ $X2=2.99 $Y2=0
r119 49 50 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.315
+ $Y2=0
r120 48 64 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.505 $Y=0
+ $X2=3.91 $Y2=0
r121 48 50 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.505 $Y=0 $X2=3.315
+ $Y2=0
r122 46 58 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.085 $Y=0 $X2=2.07
+ $Y2=0
r123 46 47 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.085 $Y=0 $X2=2.275
+ $Y2=0
r124 45 61 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.465 $Y=0
+ $X2=2.99 $Y2=0
r125 45 47 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.275
+ $Y2=0
r126 41 77 3.40825 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=5.23 $Y=0.085
+ $X2=5.332 $Y2=0
r127 41 43 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.23 $Y=0.085
+ $X2=5.23 $Y2=0.39
r128 37 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.29 $Y=0.085
+ $X2=4.29 $Y2=0
r129 37 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.29 $Y=0.085
+ $X2=4.29 $Y2=0.39
r130 33 50 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.315 $Y=0.085
+ $X2=3.315 $Y2=0
r131 33 35 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=3.315 $Y=0.085
+ $X2=3.315 $Y2=0.4
r132 29 47 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=0.085
+ $X2=2.275 $Y2=0
r133 29 31 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.275 $Y=0.085
+ $X2=2.275 $Y2=0.4
r134 25 74 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0
r135 25 27 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0.38
r136 24 71 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r137 23 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.085 $Y=0 $X2=1.21
+ $Y2=0
r138 23 24 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.085 $Y=0
+ $X2=0.345 $Y2=0
r139 19 71 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.172 $Y2=0
r140 19 21 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.215 $Y2=0.66
r141 6 43 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.095
+ $Y=0.235 $X2=5.23 $Y2=0.39
r142 5 39 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.105
+ $Y=0.235 $X2=4.29 $Y2=0.39
r143 4 35 182 $w=1.7e-07 $l=3.5812e-07 $layer=licon1_NDIFF $count=1 $X=3.055
+ $Y=0.235 $X2=3.34 $Y2=0.4
r144 3 31 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.165
+ $Y=0.235 $X2=2.3 $Y2=0.4
r145 2 27 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.25 $Y2=0.38
r146 1 21 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.66
.ends

