# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a21boi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21boi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.865000 1.065000 5.440000 1.310000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.300000 1.065000 3.695000 1.480000 ;
        RECT 3.300000 1.480000 7.120000 1.705000 ;
        RECT 5.725000 1.075000 7.120000 1.480000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 1.075000 0.670000 1.615000 ;
        RECT 0.450000 0.995000 0.670000 1.075000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.490500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.375000 0.370000 1.565000 0.615000 ;
        RECT 1.375000 0.615000 2.525000 0.695000 ;
        RECT 1.375000 0.695000 5.385000 0.865000 ;
        RECT 1.680000 1.585000 3.130000 1.705000 ;
        RECT 1.680000 1.705000 2.945000 2.035000 ;
        RECT 2.335000 0.255000 2.525000 0.615000 ;
        RECT 2.820000 0.865000 5.385000 0.895000 ;
        RECT 2.820000 0.895000 3.130000 1.585000 ;
        RECT 3.555000 0.675000 5.385000 0.695000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.360000 0.085000 ;
        RECT 0.770000  0.085000 1.155000 0.445000 ;
        RECT 1.785000  0.085000 2.165000 0.445000 ;
        RECT 2.745000  0.085000 3.385000 0.525000 ;
        RECT 6.085000  0.085000 6.275000 0.565000 ;
        RECT 7.000000  0.085000 7.240000 0.885000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 7.360000 2.805000 ;
        RECT 0.645000 2.175000 0.905000 2.635000 ;
        RECT 3.535000 2.275000 3.915000 2.635000 ;
        RECT 4.495000 2.275000 4.875000 2.635000 ;
        RECT 5.455000 2.275000 5.835000 2.635000 ;
        RECT 6.415000 2.275000 6.795000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 0.255000 0.445000 0.615000 ;
      RECT 0.090000 0.615000 1.155000 0.795000 ;
      RECT 0.095000 1.785000 1.010000 2.005000 ;
      RECT 0.095000 2.005000 0.425000 2.465000 ;
      RECT 0.840000 0.795000 1.155000 1.035000 ;
      RECT 0.840000 1.035000 2.620000 1.345000 ;
      RECT 0.840000 1.345000 1.010000 1.785000 ;
      RECT 1.180000 1.795000 1.425000 2.215000 ;
      RECT 1.180000 2.215000 3.365000 2.465000 ;
      RECT 2.055000 2.205000 3.365000 2.215000 ;
      RECT 3.165000 1.875000 7.240000 2.105000 ;
      RECT 3.165000 2.105000 3.365000 2.205000 ;
      RECT 3.565000 0.255000 5.865000 0.505000 ;
      RECT 5.095000 2.105000 5.285000 2.465000 ;
      RECT 5.605000 0.505000 5.865000 0.735000 ;
      RECT 5.605000 0.735000 6.825000 0.905000 ;
      RECT 6.050000 2.105000 6.235000 2.465000 ;
      RECT 6.445000 0.255000 6.825000 0.735000 ;
      RECT 6.990000 2.105000 7.240000 2.465000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21boi_4
