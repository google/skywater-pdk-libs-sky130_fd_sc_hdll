* File: sky130_fd_sc_hdll__nor3b_1.pxi.spice
* Created: Thu Aug 27 19:16:32 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR3B_1%A_91_199# N_A_91_199#_M1000_d
+ N_A_91_199#_M1003_d N_A_91_199#_c_46_n N_A_91_199#_M1002_g N_A_91_199#_c_47_n
+ N_A_91_199#_M1005_g N_A_91_199#_c_48_n N_A_91_199#_c_49_n N_A_91_199#_c_54_n
+ N_A_91_199#_c_87_p N_A_91_199#_c_50_n N_A_91_199#_c_51_n
+ PM_SKY130_FD_SC_HDLL__NOR3B_1%A_91_199#
x_PM_SKY130_FD_SC_HDLL__NOR3B_1%B N_B_c_102_n N_B_M1001_g N_B_c_103_n
+ N_B_M1004_g B PM_SKY130_FD_SC_HDLL__NOR3B_1%B
x_PM_SKY130_FD_SC_HDLL__NOR3B_1%A N_A_c_132_n N_A_M1006_g N_A_c_133_n
+ N_A_M1007_g A A PM_SKY130_FD_SC_HDLL__NOR3B_1%A
x_PM_SKY130_FD_SC_HDLL__NOR3B_1%C_N N_C_N_c_165_n N_C_N_c_166_n N_C_N_M1003_g
+ N_C_N_M1000_g C_N N_C_N_c_163_n N_C_N_c_164_n
+ PM_SKY130_FD_SC_HDLL__NOR3B_1%C_N
x_PM_SKY130_FD_SC_HDLL__NOR3B_1%Y N_Y_M1005_s N_Y_M1004_d N_Y_M1002_s
+ N_Y_c_199_n N_Y_c_223_p N_Y_c_195_n Y Y PM_SKY130_FD_SC_HDLL__NOR3B_1%Y
x_PM_SKY130_FD_SC_HDLL__NOR3B_1%VPWR N_VPWR_M1007_d N_VPWR_c_236_n
+ N_VPWR_c_237_n N_VPWR_c_238_n VPWR N_VPWR_c_239_n N_VPWR_c_235_n
+ PM_SKY130_FD_SC_HDLL__NOR3B_1%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR3B_1%VGND N_VGND_M1005_d N_VGND_M1006_d
+ N_VGND_c_262_n N_VGND_c_263_n N_VGND_c_264_n N_VGND_c_265_n N_VGND_c_266_n
+ N_VGND_c_267_n VGND N_VGND_c_268_n N_VGND_c_269_n
+ PM_SKY130_FD_SC_HDLL__NOR3B_1%VGND
cc_1 VNB N_A_91_199#_c_46_n 0.0312726f $X=-0.19 $Y=-0.24 $X2=0.755 $Y2=1.41
cc_2 VNB N_A_91_199#_c_47_n 0.0199704f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.995
cc_3 VNB N_A_91_199#_c_48_n 0.0035278f $X=-0.19 $Y=-0.24 $X2=0.715 $Y2=1.16
cc_4 VNB N_A_91_199#_c_49_n 3.55466e-19 $X=-0.19 $Y=-0.24 $X2=0.8 $Y2=1.785
cc_5 VNB N_A_91_199#_c_50_n 0.0219551f $X=-0.19 $Y=-0.24 $X2=2.59 $Y2=1.785
cc_6 VNB N_A_91_199#_c_51_n 0.0123834f $X=-0.19 $Y=-0.24 $X2=2.465 $Y2=0.66
cc_7 VNB N_B_c_102_n 0.0229715f $X=-0.19 $Y=-0.24 $X2=2.33 $Y2=0.465
cc_8 VNB N_B_c_103_n 0.01695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB B 0.00231247f $X=-0.19 $Y=-0.24 $X2=0.755 $Y2=1.41
cc_10 VNB N_A_c_132_n 0.0188734f $X=-0.19 $Y=-0.24 $X2=2.33 $Y2=0.465
cc_11 VNB N_A_c_133_n 0.0223932f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB A 0.00448676f $X=-0.19 $Y=-0.24 $X2=0.755 $Y2=1.41
cc_13 VNB C_N 0.0036812f $X=-0.19 $Y=-0.24 $X2=0.755 $Y2=1.985
cc_14 VNB N_C_N_c_163_n 0.0287963f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.56
cc_15 VNB N_C_N_c_164_n 0.0207066f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_16 VNB N_Y_c_195_n 0.0298186f $X=-0.19 $Y=-0.24 $X2=0.8 $Y2=1.245
cc_17 VNB Y 0.0235522f $X=-0.19 $Y=-0.24 $X2=2.465 $Y2=1.87
cc_18 VNB N_VPWR_c_235_n 0.117919f $X=-0.19 $Y=-0.24 $X2=2.465 $Y2=1.87
cc_19 VNB N_VGND_c_262_n 0.00214417f $X=-0.19 $Y=-0.24 $X2=0.755 $Y2=1.985
cc_20 VNB N_VGND_c_263_n 0.00813837f $X=-0.19 $Y=-0.24 $X2=0.715 $Y2=1.16
cc_21 VNB N_VGND_c_264_n 0.020151f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_22 VNB N_VGND_c_265_n 0.00573782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_266_n 0.0143427f $X=-0.19 $Y=-0.24 $X2=0.8 $Y2=1.785
cc_24 VNB N_VGND_c_267_n 0.00606646f $X=-0.19 $Y=-0.24 $X2=2.505 $Y2=1.87
cc_25 VNB N_VGND_c_268_n 0.021578f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_269_n 0.173768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VPB N_A_91_199#_c_46_n 0.035419f $X=-0.19 $Y=1.305 $X2=0.755 $Y2=1.41
cc_28 VPB N_A_91_199#_c_49_n 0.00111031f $X=-0.19 $Y=1.305 $X2=0.8 $Y2=1.785
cc_29 VPB N_A_91_199#_c_54_n 0.00906618f $X=-0.19 $Y=1.305 $X2=2.505 $Y2=1.87
cc_30 VPB N_A_91_199#_c_50_n 0.0211305f $X=-0.19 $Y=1.305 $X2=2.59 $Y2=1.785
cc_31 VPB N_B_c_102_n 0.0259285f $X=-0.19 $Y=1.305 $X2=2.33 $Y2=0.465
cc_32 VPB B 0.00110414f $X=-0.19 $Y=1.305 $X2=0.755 $Y2=1.41
cc_33 VPB N_A_c_133_n 0.0265102f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB A 0.00211969f $X=-0.19 $Y=1.305 $X2=0.755 $Y2=1.41
cc_35 VPB N_C_N_c_165_n 0.00968692f $X=-0.19 $Y=1.305 $X2=2.32 $Y2=1.65
cc_36 VPB N_C_N_c_166_n 0.0291017f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB C_N 0.00472078f $X=-0.19 $Y=1.305 $X2=0.755 $Y2=1.985
cc_38 VPB N_C_N_c_163_n 0.00520898f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=0.56
cc_39 VPB Y 0.0217083f $X=-0.19 $Y=1.305 $X2=2.465 $Y2=1.87
cc_40 VPB Y 0.0392564f $X=-0.19 $Y=1.305 $X2=2.465 $Y2=1.87
cc_41 VPB N_VPWR_c_236_n 0.0151799f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_237_n 0.0514459f $X=-0.19 $Y=1.305 $X2=0.755 $Y2=1.985
cc_43 VPB N_VPWR_c_238_n 0.00580385f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=0.995
cc_44 VPB N_VPWR_c_239_n 0.0233049f $X=-0.19 $Y=1.305 $X2=0.885 $Y2=1.87
cc_45 VPB N_VPWR_c_235_n 0.0522888f $X=-0.19 $Y=1.305 $X2=2.465 $Y2=1.87
cc_46 N_A_91_199#_c_46_n N_B_c_102_n 0.0795081f $X=0.755 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_47 N_A_91_199#_c_48_n N_B_c_102_n 5.77871e-19 $X=0.715 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_48 N_A_91_199#_c_49_n N_B_c_102_n 7.37579e-19 $X=0.8 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_49 N_A_91_199#_c_54_n N_B_c_102_n 0.0148341f $X=2.505 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_50 N_A_91_199#_c_47_n N_B_c_103_n 0.0218768f $X=0.78 $Y=0.995 $X2=0 $Y2=0
cc_51 N_A_91_199#_c_46_n B 0.0033106f $X=0.755 $Y=1.41 $X2=0 $Y2=0
cc_52 N_A_91_199#_c_48_n B 0.0143616f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_53 N_A_91_199#_c_49_n B 0.0236161f $X=0.8 $Y=1.785 $X2=0 $Y2=0
cc_54 N_A_91_199#_c_54_n B 0.0146342f $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_55 N_A_91_199#_c_54_n N_A_c_133_n 0.0152226f $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_56 N_A_91_199#_c_54_n A 0.019405f $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_57 N_A_91_199#_c_50_n N_C_N_c_165_n 0.0017419f $X=2.59 $Y=1.785 $X2=0 $Y2=0
cc_58 N_A_91_199#_c_54_n N_C_N_c_166_n 0.0112684f $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_59 N_A_91_199#_c_50_n N_C_N_c_166_n 0.0042189f $X=2.59 $Y=1.785 $X2=0 $Y2=0
cc_60 N_A_91_199#_c_54_n C_N 0.0247264f $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_61 N_A_91_199#_c_50_n C_N 0.0480802f $X=2.59 $Y=1.785 $X2=0 $Y2=0
cc_62 N_A_91_199#_c_54_n N_C_N_c_163_n 0.00250852f $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_63 N_A_91_199#_c_50_n N_C_N_c_163_n 0.00844447f $X=2.59 $Y=1.785 $X2=0 $Y2=0
cc_64 N_A_91_199#_c_51_n N_C_N_c_163_n 0.00255699f $X=2.465 $Y=0.66 $X2=0 $Y2=0
cc_65 N_A_91_199#_c_50_n N_C_N_c_164_n 0.00525065f $X=2.59 $Y=1.785 $X2=0 $Y2=0
cc_66 N_A_91_199#_c_51_n N_C_N_c_164_n 0.00142049f $X=2.465 $Y=0.66 $X2=0 $Y2=0
cc_67 N_A_91_199#_c_46_n N_Y_c_199_n 0.00232517f $X=0.755 $Y=1.41 $X2=0 $Y2=0
cc_68 N_A_91_199#_c_47_n N_Y_c_199_n 0.0125139f $X=0.78 $Y=0.995 $X2=0 $Y2=0
cc_69 N_A_91_199#_c_48_n N_Y_c_199_n 0.0130315f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A_91_199#_c_46_n N_Y_c_195_n 0.00362982f $X=0.755 $Y=1.41 $X2=0 $Y2=0
cc_71 N_A_91_199#_c_47_n N_Y_c_195_n 0.0133191f $X=0.78 $Y=0.995 $X2=0 $Y2=0
cc_72 N_A_91_199#_c_48_n N_Y_c_195_n 0.0104687f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_91_199#_c_46_n Y 0.041499f $X=0.755 $Y=1.41 $X2=0 $Y2=0
cc_74 N_A_91_199#_c_47_n Y 0.00304618f $X=0.78 $Y=0.995 $X2=0 $Y2=0
cc_75 N_A_91_199#_c_48_n Y 0.0223568f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_91_199#_c_49_n Y 0.0309189f $X=0.8 $Y=1.785 $X2=0 $Y2=0
cc_77 N_A_91_199#_c_87_p Y 0.0143562f $X=0.885 $Y=1.87 $X2=0 $Y2=0
cc_78 N_A_91_199#_c_54_n A_169_297# 0.00939003f $X=2.505 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_79 N_A_91_199#_c_54_n A_263_297# 0.00772933f $X=2.505 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_80 N_A_91_199#_c_54_n N_VPWR_M1007_d 0.00754471f $X=2.505 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_81 N_A_91_199#_c_54_n N_VPWR_c_236_n 0.0246758f $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_82 N_A_91_199#_c_46_n N_VPWR_c_237_n 0.00702461f $X=0.755 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A_91_199#_c_46_n N_VPWR_c_235_n 0.00990948f $X=0.755 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_91_199#_c_54_n N_VPWR_c_235_n 0.0511636f $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_85 N_A_91_199#_c_87_p N_VPWR_c_235_n 0.00606489f $X=0.885 $Y=1.87 $X2=0 $Y2=0
cc_86 N_A_91_199#_c_47_n N_VGND_c_262_n 0.0115037f $X=0.78 $Y=0.995 $X2=0 $Y2=0
cc_87 N_A_91_199#_c_51_n N_VGND_c_263_n 0.0134413f $X=2.465 $Y=0.66 $X2=0 $Y2=0
cc_88 N_A_91_199#_c_47_n N_VGND_c_264_n 0.00199015f $X=0.78 $Y=0.995 $X2=0 $Y2=0
cc_89 N_A_91_199#_c_51_n N_VGND_c_268_n 0.00846211f $X=2.465 $Y=0.66 $X2=0 $Y2=0
cc_90 N_A_91_199#_c_47_n N_VGND_c_269_n 0.00384791f $X=0.78 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A_91_199#_c_51_n N_VGND_c_269_n 0.00964063f $X=2.465 $Y=0.66 $X2=0 $Y2=0
cc_92 N_B_c_103_n N_A_c_132_n 0.0241646f $X=1.25 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_93 N_B_c_102_n N_A_c_133_n 0.0791974f $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_94 B N_A_c_133_n 5.79914e-19 $X=1.115 $Y=1.105 $X2=0 $Y2=0
cc_95 N_B_c_102_n A 0.00398212f $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_96 B A 0.0483033f $X=1.115 $Y=1.105 $X2=0 $Y2=0
cc_97 N_B_c_102_n N_Y_c_199_n 0.00277939f $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_98 N_B_c_103_n N_Y_c_199_n 0.0118666f $X=1.25 $Y=0.995 $X2=0 $Y2=0
cc_99 B N_Y_c_199_n 0.0170682f $X=1.115 $Y=1.105 $X2=0 $Y2=0
cc_100 B A_169_297# 0.00136066f $X=1.115 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_101 N_B_c_102_n N_VPWR_c_236_n 0.00287642f $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_102 N_B_c_102_n N_VPWR_c_237_n 0.00702461f $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_103 N_B_c_102_n N_VPWR_c_235_n 0.00727922f $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_104 N_B_c_103_n N_VGND_c_262_n 0.00162962f $X=1.25 $Y=0.995 $X2=0 $Y2=0
cc_105 N_B_c_103_n N_VGND_c_263_n 8.65906e-19 $X=1.25 $Y=0.995 $X2=0 $Y2=0
cc_106 N_B_c_103_n N_VGND_c_266_n 0.00428022f $X=1.25 $Y=0.995 $X2=0 $Y2=0
cc_107 N_B_c_103_n N_VGND_c_269_n 0.00585784f $X=1.25 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A_c_133_n N_C_N_c_165_n 0.00864271f $X=1.695 $Y=1.41 $X2=0 $Y2=0
cc_109 A N_C_N_c_165_n 4.80258e-19 $X=1.645 $Y=1.105 $X2=0 $Y2=0
cc_110 N_A_c_133_n N_C_N_c_166_n 0.0198867f $X=1.695 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A_c_133_n C_N 0.00322412f $X=1.695 $Y=1.41 $X2=0 $Y2=0
cc_112 A C_N 0.0452322f $X=1.645 $Y=1.105 $X2=0 $Y2=0
cc_113 N_A_c_133_n N_C_N_c_163_n 0.0203255f $X=1.695 $Y=1.41 $X2=0 $Y2=0
cc_114 A N_C_N_c_163_n 2.77811e-19 $X=1.645 $Y=1.105 $X2=0 $Y2=0
cc_115 N_A_c_132_n N_C_N_c_164_n 0.00917075f $X=1.67 $Y=0.995 $X2=0 $Y2=0
cc_116 A N_Y_c_199_n 0.00593246f $X=1.645 $Y=1.105 $X2=0 $Y2=0
cc_117 A A_263_297# 0.00190371f $X=1.645 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_118 N_A_c_133_n N_VPWR_c_236_n 0.0179797f $X=1.695 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_c_133_n N_VPWR_c_237_n 0.00427505f $X=1.695 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_c_133_n N_VPWR_c_235_n 0.00401989f $X=1.695 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_c_132_n N_VGND_c_263_n 0.0121247f $X=1.67 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A_c_133_n N_VGND_c_263_n 0.00562536f $X=1.695 $Y=1.41 $X2=0 $Y2=0
cc_123 A N_VGND_c_263_n 0.00587298f $X=1.645 $Y=1.105 $X2=0 $Y2=0
cc_124 N_A_c_132_n N_VGND_c_266_n 0.0046653f $X=1.67 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_c_132_n N_VGND_c_269_n 0.00799591f $X=1.67 $Y=0.995 $X2=0 $Y2=0
cc_126 C_N N_VPWR_M1007_d 0.00188663f $X=2.165 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_127 N_C_N_c_166_n N_VPWR_c_236_n 0.002206f $X=2.23 $Y=1.575 $X2=0 $Y2=0
cc_128 N_C_N_c_166_n N_VPWR_c_239_n 0.00482866f $X=2.23 $Y=1.575 $X2=0 $Y2=0
cc_129 N_C_N_c_166_n N_VPWR_c_235_n 0.00551811f $X=2.23 $Y=1.575 $X2=0 $Y2=0
cc_130 C_N N_VGND_c_263_n 0.0099047f $X=2.165 $Y=1.105 $X2=0 $Y2=0
cc_131 N_C_N_c_164_n N_VGND_c_263_n 0.00652097f $X=2.28 $Y=0.995 $X2=0 $Y2=0
cc_132 N_C_N_c_164_n N_VGND_c_268_n 0.00510437f $X=2.28 $Y=0.995 $X2=0 $Y2=0
cc_133 N_C_N_c_164_n N_VGND_c_269_n 0.00512902f $X=2.28 $Y=0.995 $X2=0 $Y2=0
cc_134 Y N_VPWR_c_237_n 0.0306029f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_135 N_Y_M1002_s N_VPWR_c_235_n 0.00687828f $X=0.335 $Y=1.485 $X2=0 $Y2=0
cc_136 Y N_VPWR_c_235_n 0.017555f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_137 N_Y_c_199_n N_VGND_M1005_d 0.00812071f $X=1.375 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_138 N_Y_c_199_n N_VGND_c_262_n 0.0214497f $X=1.375 $Y=0.74 $X2=0 $Y2=0
cc_139 N_Y_c_195_n N_VGND_c_262_n 0.0186889f $X=0.44 $Y=0.39 $X2=0 $Y2=0
cc_140 N_Y_c_199_n N_VGND_c_264_n 0.00233441f $X=1.375 $Y=0.74 $X2=0 $Y2=0
cc_141 N_Y_c_195_n N_VGND_c_264_n 0.0364239f $X=0.44 $Y=0.39 $X2=0 $Y2=0
cc_142 N_Y_c_199_n N_VGND_c_266_n 0.0029785f $X=1.375 $Y=0.74 $X2=0 $Y2=0
cc_143 N_Y_c_223_p N_VGND_c_266_n 0.00825814f $X=1.46 $Y=0.495 $X2=0 $Y2=0
cc_144 N_Y_M1005_s N_VGND_c_269_n 0.00357812f $X=0.315 $Y=0.235 $X2=0 $Y2=0
cc_145 N_Y_M1004_d N_VGND_c_269_n 0.00415164f $X=1.325 $Y=0.235 $X2=0 $Y2=0
cc_146 N_Y_c_199_n N_VGND_c_269_n 0.011344f $X=1.375 $Y=0.74 $X2=0 $Y2=0
cc_147 N_Y_c_223_p N_VGND_c_269_n 0.00623764f $X=1.46 $Y=0.495 $X2=0 $Y2=0
cc_148 N_Y_c_195_n N_VGND_c_269_n 0.0198876f $X=0.44 $Y=0.39 $X2=0 $Y2=0
cc_149 A_169_297# N_VPWR_c_235_n 0.00394308f $X=0.845 $Y=1.485 $X2=2.465
+ $Y2=1.87
cc_150 A_263_297# N_VPWR_c_235_n 0.00394367f $X=1.315 $Y=1.485 $X2=2.465
+ $Y2=1.87
