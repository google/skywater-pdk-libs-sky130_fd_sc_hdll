* File: sky130_fd_sc_hdll__nor4_2.pxi.spice
* Created: Wed Sep  2 08:41:05 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR4_2%A N_A_c_71_n N_A_M1006_g N_A_c_75_n N_A_M1001_g
+ N_A_c_76_n N_A_M1011_g N_A_c_72_n N_A_M1013_g A N_A_c_74_n A
+ PM_SKY130_FD_SC_HDLL__NOR4_2%A
x_PM_SKY130_FD_SC_HDLL__NOR4_2%B N_B_c_108_n N_B_M1007_g N_B_c_112_n N_B_M1003_g
+ N_B_c_113_n N_B_M1005_g N_B_c_109_n N_B_M1012_g B N_B_c_111_n B
+ PM_SKY130_FD_SC_HDLL__NOR4_2%B
x_PM_SKY130_FD_SC_HDLL__NOR4_2%C N_C_c_149_n N_C_M1002_g N_C_c_153_n N_C_M1000_g
+ N_C_c_154_n N_C_M1015_g N_C_c_150_n N_C_M1009_g C N_C_c_151_n N_C_c_152_n C
+ PM_SKY130_FD_SC_HDLL__NOR4_2%C
x_PM_SKY130_FD_SC_HDLL__NOR4_2%D N_D_c_187_n N_D_M1004_g N_D_c_191_n N_D_M1008_g
+ N_D_c_192_n N_D_M1010_g N_D_c_188_n N_D_M1014_g D N_D_c_189_n N_D_c_190_n D
+ PM_SKY130_FD_SC_HDLL__NOR4_2%D
x_PM_SKY130_FD_SC_HDLL__NOR4_2%A_27_297# N_A_27_297#_M1001_s N_A_27_297#_M1011_s
+ N_A_27_297#_M1005_d N_A_27_297#_c_230_n N_A_27_297#_c_253_p
+ N_A_27_297#_c_231_n N_A_27_297#_c_249_p N_A_27_297#_c_232_n
+ N_A_27_297#_c_233_n N_A_27_297#_c_234_n PM_SKY130_FD_SC_HDLL__NOR4_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__NOR4_2%VPWR N_VPWR_M1001_d N_VPWR_c_267_n VPWR
+ N_VPWR_c_268_n N_VPWR_c_266_n N_VPWR_c_270_n VPWR
+ PM_SKY130_FD_SC_HDLL__NOR4_2%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR4_2%A_309_297# N_A_309_297#_M1003_s
+ N_A_309_297#_M1000_d N_A_309_297#_c_316_n N_A_309_297#_c_312_n
+ N_A_309_297#_c_324_n N_A_309_297#_c_329_p
+ PM_SKY130_FD_SC_HDLL__NOR4_2%A_309_297#
x_PM_SKY130_FD_SC_HDLL__NOR4_2%A_515_297# N_A_515_297#_M1000_s
+ N_A_515_297#_M1015_s N_A_515_297#_M1010_d N_A_515_297#_c_331_n
+ N_A_515_297#_c_332_n N_A_515_297#_c_349_n N_A_515_297#_c_333_n
+ N_A_515_297#_c_363_p N_A_515_297#_c_334_n
+ PM_SKY130_FD_SC_HDLL__NOR4_2%A_515_297#
x_PM_SKY130_FD_SC_HDLL__NOR4_2%Y N_Y_M1006_d N_Y_M1007_s N_Y_M1002_s N_Y_M1004_d
+ N_Y_M1008_s N_Y_c_380_n N_Y_c_367_n N_Y_c_368_n N_Y_c_390_n N_Y_c_369_n
+ N_Y_c_398_n N_Y_c_370_n N_Y_c_406_n N_Y_c_377_n N_Y_c_371_n N_Y_c_372_n
+ N_Y_c_373_n N_Y_c_374_n N_Y_c_378_n Y N_Y_c_376_n
+ PM_SKY130_FD_SC_HDLL__NOR4_2%Y
x_PM_SKY130_FD_SC_HDLL__NOR4_2%VGND N_VGND_M1006_s N_VGND_M1013_s N_VGND_M1012_d
+ N_VGND_M1002_d N_VGND_M1009_d N_VGND_M1014_s N_VGND_c_470_n N_VGND_c_471_n
+ N_VGND_c_472_n N_VGND_c_473_n N_VGND_c_474_n N_VGND_c_475_n N_VGND_c_476_n
+ N_VGND_c_477_n N_VGND_c_478_n VGND N_VGND_c_479_n N_VGND_c_480_n
+ N_VGND_c_481_n N_VGND_c_482_n N_VGND_c_483_n PM_SKY130_FD_SC_HDLL__NOR4_2%VGND
cc_1 VNB N_A_c_71_n 0.0223809f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_72_n 0.0169338f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_3 VNB A 0.0140266f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_4 VNB N_A_c_74_n 0.0440201f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_5 VNB N_B_c_108_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_6 VNB N_B_c_109_n 0.0224106f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_7 VNB B 0.0080257f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_8 VNB N_B_c_111_n 0.0426802f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_9 VNB N_C_c_149_n 0.0224149f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_10 VNB N_C_c_150_n 0.0169338f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_11 VNB N_C_c_151_n 0.0167322f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_12 VNB N_C_c_152_n 0.0440143f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_13 VNB N_D_c_187_n 0.0169148f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_14 VNB N_D_c_188_n 0.0201356f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_15 VNB N_D_c_189_n 0.00459812f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_16 VNB N_D_c_190_n 0.0391131f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_17 VNB N_VPWR_c_266_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_18 VNB N_Y_c_367_n 0.00338427f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_19 VNB N_Y_c_368_n 0.00295675f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.202
cc_20 VNB N_Y_c_369_n 0.0158955f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_370_n 0.00317397f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_Y_c_371_n 0.00199628f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_Y_c_372_n 0.00276479f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_Y_c_373_n 0.00289004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_Y_c_374_n 0.00292451f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB Y 0.0231557f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_Y_c_376_n 0.0117119f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_470_n 0.0103614f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_29 VNB N_VGND_c_471_n 0.0356812f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.202
cc_30 VNB N_VGND_c_472_n 0.020063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_473_n 0.00471543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_474_n 0.00471543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_475_n 0.0153448f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_476_n 0.0187002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_477_n 0.0192928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_478_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_479_n 0.0192928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_480_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_481_n 0.0192928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_482_n 0.0276407f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_483_n 0.258393f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VPB N_A_c_75_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_43 VPB N_A_c_76_n 0.0161064f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_44 VPB N_A_c_74_n 0.022695f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_45 VPB N_B_c_112_n 0.0161064f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_46 VPB N_B_c_113_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_47 VPB N_B_c_111_n 0.022695f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_48 VPB N_C_c_153_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_49 VPB N_C_c_154_n 0.0161064f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_50 VPB N_C_c_152_n 0.022695f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_51 VPB N_D_c_191_n 0.0164226f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_52 VPB N_D_c_192_n 0.0191753f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_53 VPB N_D_c_190_n 0.021846f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_54 VPB N_A_27_297#_c_230_n 0.00403131f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_55 VPB N_A_27_297#_c_231_n 0.0020765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_297#_c_232_n 0.00199216f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_57 VPB N_A_27_297#_c_233_n 0.00322557f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_297#_c_234_n 0.00360002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_267_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.985
cc_60 VPB N_VPWR_c_268_n 0.104745f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.202
cc_61 VPB N_VPWR_c_266_n 0.0579497f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_62 VPB N_VPWR_c_270_n 0.0244347f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.202
cc_63 VPB N_A_309_297#_c_312_n 0.0128761f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.56
cc_64 VPB N_A_515_297#_c_331_n 0.0020765f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.56
cc_65 VPB N_A_515_297#_c_332_n 0.00326945f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_515_297#_c_333_n 0.00692367f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_67 VPB N_A_515_297#_c_334_n 0.00269738f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_Y_c_377_n 0.0196351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_Y_c_378_n 0.00164325f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB Y 0.0088309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 N_A_c_72_n N_B_c_108_n 0.0242642f $X=1.01 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_72 N_A_c_76_n N_B_c_112_n 0.00985632f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_73 A B 0.0152605f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A_c_74_n B 0.0018186f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_75 N_A_c_74_n N_B_c_111_n 0.0242642f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_76 A N_A_27_297#_c_230_n 0.0175673f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_77 N_A_c_75_n N_A_27_297#_c_231_n 0.0158351f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A_c_76_n N_A_27_297#_c_231_n 0.016363f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_79 A N_A_27_297#_c_231_n 0.0431894f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_80 N_A_c_74_n N_A_27_297#_c_231_n 0.00794509f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_81 N_A_c_75_n N_VPWR_c_267_n 0.00300743f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A_c_76_n N_VPWR_c_267_n 0.00300743f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A_c_76_n N_VPWR_c_268_n 0.00702461f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_c_75_n N_VPWR_c_266_n 0.0133387f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A_c_76_n N_VPWR_c_266_n 0.0124344f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A_c_75_n N_VPWR_c_270_n 0.00702461f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_c_72_n N_Y_c_380_n 0.00594127f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_88 N_A_c_72_n N_Y_c_367_n 0.010339f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_89 A N_Y_c_367_n 0.00446377f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_90 N_A_c_71_n N_Y_c_368_n 2.15763e-19 $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A_c_72_n N_Y_c_368_n 6.9417e-19 $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_92 A N_Y_c_368_n 0.0309026f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_93 N_A_c_74_n N_Y_c_368_n 0.00486271f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_94 N_A_c_71_n N_VGND_c_471_n 0.00497868f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_95 A N_VGND_c_471_n 0.0140538f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_96 N_A_c_71_n N_VGND_c_472_n 0.00585385f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_c_72_n N_VGND_c_472_n 0.00431352f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_98 N_A_c_72_n N_VGND_c_473_n 0.00268723f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A_c_71_n N_VGND_c_483_n 0.0117523f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_100 N_A_c_72_n N_VGND_c_483_n 0.00606926f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_101 B N_C_c_151_n 0.0140819f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_102 N_B_c_111_n N_C_c_151_n 0.0012237f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_103 N_B_c_112_n N_A_27_297#_c_232_n 0.0156202f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_104 N_B_c_113_n N_A_27_297#_c_232_n 0.013085f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_105 B N_A_27_297#_c_232_n 0.0487774f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_106 N_B_c_111_n N_A_27_297#_c_232_n 0.00789593f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_107 B N_A_27_297#_c_233_n 0.00942636f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_108 B N_A_27_297#_c_234_n 0.0089871f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_109 N_B_c_112_n N_VPWR_c_268_n 0.00702461f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_110 N_B_c_113_n N_VPWR_c_268_n 0.00429453f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_111 N_B_c_112_n N_VPWR_c_266_n 0.0126324f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_112 N_B_c_113_n N_VPWR_c_266_n 0.00739666f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_113 N_B_c_113_n N_A_309_297#_c_312_n 0.0136098f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_114 N_B_c_113_n N_A_515_297#_c_334_n 4.82843e-19 $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_115 N_B_c_108_n N_Y_c_380_n 5.22185e-19 $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_116 N_B_c_108_n N_Y_c_367_n 0.0106151f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_117 B N_Y_c_367_n 0.0199299f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_118 N_B_c_109_n N_Y_c_390_n 0.0105452f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_119 N_B_c_109_n N_Y_c_369_n 0.0117693f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_120 B N_Y_c_369_n 0.0181464f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_121 N_B_c_109_n N_Y_c_372_n 7.24382e-19 $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_122 B N_Y_c_372_n 0.0309026f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_123 N_B_c_111_n N_Y_c_372_n 0.00486271f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_124 N_B_c_108_n N_VGND_c_473_n 0.00268723f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_125 N_B_c_108_n N_VGND_c_481_n 0.00437852f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_126 N_B_c_109_n N_VGND_c_481_n 0.00431352f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_127 N_B_c_109_n N_VGND_c_482_n 0.00483063f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_128 N_B_c_108_n N_VGND_c_483_n 0.00615622f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_129 N_B_c_109_n N_VGND_c_483_n 0.00736566f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_130 N_C_c_150_n N_D_c_187_n 0.0242362f $X=3.45 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_131 N_C_c_154_n N_D_c_191_n 0.00971598f $X=3.425 $Y=1.41 $X2=0 $Y2=0
cc_132 N_C_c_151_n N_D_c_189_n 0.0125035f $X=3.19 $Y=1.16 $X2=0 $Y2=0
cc_133 N_C_c_152_n N_D_c_189_n 0.00215304f $X=3.425 $Y=1.202 $X2=0 $Y2=0
cc_134 N_C_c_152_n N_D_c_190_n 0.0242362f $X=3.425 $Y=1.202 $X2=0 $Y2=0
cc_135 N_C_c_153_n N_A_27_297#_c_234_n 4.82843e-19 $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_136 N_C_c_153_n N_VPWR_c_268_n 0.00429453f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_137 N_C_c_154_n N_VPWR_c_268_n 0.00702461f $X=3.425 $Y=1.41 $X2=0 $Y2=0
cc_138 N_C_c_153_n N_VPWR_c_266_n 0.00739666f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_139 N_C_c_154_n N_VPWR_c_266_n 0.0126324f $X=3.425 $Y=1.41 $X2=0 $Y2=0
cc_140 N_C_c_153_n N_A_309_297#_c_312_n 0.0136098f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_141 N_C_c_153_n N_A_515_297#_c_331_n 0.013085f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_142 N_C_c_154_n N_A_515_297#_c_331_n 0.0175467f $X=3.425 $Y=1.41 $X2=0 $Y2=0
cc_143 N_C_c_151_n N_A_515_297#_c_331_n 0.0362994f $X=3.19 $Y=1.16 $X2=0 $Y2=0
cc_144 N_C_c_152_n N_A_515_297#_c_331_n 0.00794509f $X=3.425 $Y=1.202 $X2=0
+ $Y2=0
cc_145 N_C_c_151_n N_A_515_297#_c_334_n 0.0213978f $X=3.19 $Y=1.16 $X2=0 $Y2=0
cc_146 N_C_c_149_n N_Y_c_369_n 0.01289f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_147 N_C_c_151_n N_Y_c_369_n 0.0449088f $X=3.19 $Y=1.16 $X2=0 $Y2=0
cc_148 N_C_c_150_n N_Y_c_398_n 0.00594127f $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_149 N_C_c_150_n N_Y_c_370_n 0.0111336f $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_150 N_C_c_150_n N_Y_c_373_n 9.09687e-19 $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_151 N_C_c_151_n N_Y_c_373_n 0.0281168f $X=3.19 $Y=1.16 $X2=0 $Y2=0
cc_152 N_C_c_152_n N_Y_c_373_n 0.00486271f $X=3.425 $Y=1.202 $X2=0 $Y2=0
cc_153 N_C_c_150_n N_VGND_c_474_n 0.00268723f $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_154 N_C_c_149_n N_VGND_c_477_n 0.00437852f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_155 N_C_c_150_n N_VGND_c_477_n 0.00431352f $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_156 N_C_c_149_n N_VGND_c_482_n 0.00483063f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_157 N_C_c_149_n N_VGND_c_483_n 0.00745263f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_158 N_C_c_150_n N_VGND_c_483_n 0.00606926f $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_159 N_D_c_191_n N_VPWR_c_268_n 0.00429453f $X=3.895 $Y=1.41 $X2=0 $Y2=0
cc_160 N_D_c_192_n N_VPWR_c_268_n 0.00429453f $X=4.365 $Y=1.41 $X2=0 $Y2=0
cc_161 N_D_c_191_n N_VPWR_c_266_n 0.00609021f $X=3.895 $Y=1.41 $X2=0 $Y2=0
cc_162 N_D_c_192_n N_VPWR_c_266_n 0.00711643f $X=4.365 $Y=1.41 $X2=0 $Y2=0
cc_163 N_D_c_191_n N_A_515_297#_c_332_n 3.19638e-19 $X=3.895 $Y=1.41 $X2=0 $Y2=0
cc_164 N_D_c_189_n N_A_515_297#_c_332_n 0.0124257f $X=4.11 $Y=1.16 $X2=0 $Y2=0
cc_165 N_D_c_191_n N_A_515_297#_c_333_n 0.0143578f $X=3.895 $Y=1.41 $X2=0 $Y2=0
cc_166 N_D_c_192_n N_A_515_297#_c_333_n 0.0113679f $X=4.365 $Y=1.41 $X2=0 $Y2=0
cc_167 N_D_c_187_n N_Y_c_398_n 5.22185e-19 $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_168 N_D_c_187_n N_Y_c_370_n 0.0106151f $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_169 N_D_c_189_n N_Y_c_370_n 0.0226199f $X=4.11 $Y=1.16 $X2=0 $Y2=0
cc_170 N_D_c_188_n N_Y_c_406_n 0.0105201f $X=4.39 $Y=0.995 $X2=0 $Y2=0
cc_171 N_D_c_192_n N_Y_c_377_n 0.0152669f $X=4.365 $Y=1.41 $X2=0 $Y2=0
cc_172 N_D_c_190_n N_Y_c_377_n 3.54534e-19 $X=4.365 $Y=1.202 $X2=0 $Y2=0
cc_173 N_D_c_188_n N_Y_c_371_n 0.0130105f $X=4.39 $Y=0.995 $X2=0 $Y2=0
cc_174 N_D_c_188_n N_Y_c_374_n 8.76687e-19 $X=4.39 $Y=0.995 $X2=0 $Y2=0
cc_175 N_D_c_189_n N_Y_c_374_n 0.0264866f $X=4.11 $Y=1.16 $X2=0 $Y2=0
cc_176 N_D_c_190_n N_Y_c_374_n 0.00486271f $X=4.365 $Y=1.202 $X2=0 $Y2=0
cc_177 N_D_c_191_n N_Y_c_378_n 2.97034e-19 $X=3.895 $Y=1.41 $X2=0 $Y2=0
cc_178 N_D_c_192_n N_Y_c_378_n 0.0117238f $X=4.365 $Y=1.41 $X2=0 $Y2=0
cc_179 N_D_c_189_n N_Y_c_378_n 0.0191995f $X=4.11 $Y=1.16 $X2=0 $Y2=0
cc_180 N_D_c_190_n N_Y_c_378_n 0.00596982f $X=4.365 $Y=1.202 $X2=0 $Y2=0
cc_181 N_D_c_192_n Y 0.00168498f $X=4.365 $Y=1.41 $X2=0 $Y2=0
cc_182 N_D_c_188_n Y 0.0182825f $X=4.39 $Y=0.995 $X2=0 $Y2=0
cc_183 N_D_c_189_n Y 0.0103327f $X=4.11 $Y=1.16 $X2=0 $Y2=0
cc_184 N_D_c_187_n N_VGND_c_474_n 0.00268723f $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_185 N_D_c_188_n N_VGND_c_476_n 0.0045387f $X=4.39 $Y=0.995 $X2=0 $Y2=0
cc_186 N_D_c_187_n N_VGND_c_479_n 0.00437852f $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_187 N_D_c_188_n N_VGND_c_479_n 0.00431352f $X=4.39 $Y=0.995 $X2=0 $Y2=0
cc_188 N_D_c_187_n N_VGND_c_483_n 0.00615622f $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_189 N_D_c_188_n N_VGND_c_483_n 0.00714059f $X=4.39 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_27_297#_c_231_n N_VPWR_M1001_d 0.00187091f $X=1.095 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_191 N_A_27_297#_c_231_n N_VPWR_c_267_n 0.0143191f $X=1.095 $Y=1.54 $X2=0
+ $Y2=0
cc_192 N_A_27_297#_c_249_p N_VPWR_c_268_n 0.0149311f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_193 N_A_27_297#_M1001_s N_VPWR_c_266_n 0.00358889f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_194 N_A_27_297#_M1011_s N_VPWR_c_266_n 0.00370124f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_195 N_A_27_297#_M1005_d N_VPWR_c_266_n 0.00234744f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_196 N_A_27_297#_c_253_p N_VPWR_c_266_n 0.00974347f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_197 N_A_27_297#_c_249_p N_VPWR_c_266_n 0.00955092f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_198 N_A_27_297#_c_253_p N_VPWR_c_270_n 0.0165369f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_199 N_A_27_297#_c_232_n N_A_309_297#_M1003_s 0.00187091f $X=2.035 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_200 N_A_27_297#_c_232_n N_A_309_297#_c_316_n 0.0143018f $X=2.035 $Y=1.54
+ $X2=0 $Y2=0
cc_201 N_A_27_297#_M1005_d N_A_309_297#_c_312_n 0.00622794f $X=2.015 $Y=1.485
+ $X2=0 $Y2=0
cc_202 N_A_27_297#_c_232_n N_A_309_297#_c_312_n 0.00385532f $X=2.035 $Y=1.54
+ $X2=0 $Y2=0
cc_203 N_A_27_297#_c_234_n N_A_309_297#_c_312_n 0.0161349f $X=2.16 $Y=1.62 $X2=0
+ $Y2=0
cc_204 N_A_27_297#_c_234_n N_A_515_297#_c_334_n 0.0346205f $X=2.16 $Y=1.62 $X2=0
+ $Y2=0
cc_205 N_A_27_297#_c_231_n N_Y_c_367_n 0.00217122f $X=1.095 $Y=1.54 $X2=0 $Y2=0
cc_206 N_A_27_297#_c_233_n N_Y_c_367_n 0.00524452f $X=1.22 $Y=1.62 $X2=0 $Y2=0
cc_207 N_A_27_297#_c_234_n N_Y_c_369_n 0.00542522f $X=2.16 $Y=1.62 $X2=0 $Y2=0
cc_208 N_A_27_297#_c_230_n N_VGND_c_471_n 0.00206382f $X=0.277 $Y=1.625 $X2=0
+ $Y2=0
cc_209 N_VPWR_c_266_n N_A_309_297#_M1003_s 0.00297222f $X=4.83 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_210 N_VPWR_c_266_n N_A_309_297#_M1000_d 0.00297222f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_211 N_VPWR_c_268_n N_A_309_297#_c_312_n 0.089449f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_212 N_VPWR_c_266_n N_A_309_297#_c_312_n 0.0543961f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_213 N_VPWR_c_268_n N_A_309_297#_c_324_n 0.0149886f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_214 N_VPWR_c_266_n N_A_309_297#_c_324_n 0.00962421f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_215 N_VPWR_c_266_n N_A_515_297#_M1000_s 0.00234744f $X=4.83 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_216 N_VPWR_c_266_n N_A_515_297#_M1015_s 0.00297222f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_217 N_VPWR_c_266_n N_A_515_297#_M1010_d 0.00217519f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_218 N_VPWR_c_268_n N_A_515_297#_c_349_n 0.015002f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_219 N_VPWR_c_266_n N_A_515_297#_c_349_n 0.00962794f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_220 N_VPWR_c_268_n N_A_515_297#_c_333_n 0.0549564f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_221 N_VPWR_c_266_n N_A_515_297#_c_333_n 0.0335386f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_222 N_VPWR_c_266_n N_Y_M1008_s 0.00232895f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_223 N_A_309_297#_c_312_n N_A_515_297#_M1000_s 0.00622794f $X=3.065 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_224 N_A_309_297#_M1000_d N_A_515_297#_c_331_n 0.00187091f $X=3.045 $Y=1.485
+ $X2=0 $Y2=0
cc_225 N_A_309_297#_c_312_n N_A_515_297#_c_331_n 0.00385532f $X=3.065 $Y=2.38
+ $X2=0 $Y2=0
cc_226 N_A_309_297#_c_329_p N_A_515_297#_c_331_n 0.0143018f $X=3.19 $Y=1.96
+ $X2=0 $Y2=0
cc_227 N_A_309_297#_c_312_n N_A_515_297#_c_334_n 0.0161349f $X=3.065 $Y=2.38
+ $X2=0 $Y2=0
cc_228 N_A_515_297#_c_333_n N_Y_M1008_s 0.00352392f $X=4.475 $Y=2.38 $X2=0 $Y2=0
cc_229 N_A_515_297#_c_331_n N_Y_c_370_n 0.00384583f $X=3.535 $Y=1.54 $X2=0 $Y2=0
cc_230 N_A_515_297#_c_332_n N_Y_c_370_n 0.00393339f $X=3.66 $Y=1.625 $X2=0 $Y2=0
cc_231 N_A_515_297#_M1010_d N_Y_c_377_n 0.00298791f $X=4.455 $Y=1.485 $X2=0
+ $Y2=0
cc_232 N_A_515_297#_c_333_n N_Y_c_377_n 0.00353225f $X=4.475 $Y=2.38 $X2=0 $Y2=0
cc_233 N_A_515_297#_c_363_p N_Y_c_377_n 0.0181502f $X=4.6 $Y=1.96 $X2=0 $Y2=0
cc_234 N_A_515_297#_c_331_n N_Y_c_373_n 0.00110124f $X=3.535 $Y=1.54 $X2=0 $Y2=0
cc_235 N_A_515_297#_c_332_n N_Y_c_378_n 0.00203916f $X=3.66 $Y=1.625 $X2=0 $Y2=0
cc_236 N_A_515_297#_c_333_n N_Y_c_378_n 0.0143553f $X=4.475 $Y=2.38 $X2=0 $Y2=0
cc_237 N_Y_c_367_n N_VGND_M1013_s 0.00162089f $X=1.51 $Y=0.815 $X2=0 $Y2=0
cc_238 N_Y_c_369_n N_VGND_M1012_d 0.00320259f $X=3.01 $Y=0.815 $X2=0 $Y2=0
cc_239 N_Y_c_369_n N_VGND_M1002_d 0.00320259f $X=3.01 $Y=0.815 $X2=0 $Y2=0
cc_240 N_Y_c_370_n N_VGND_M1009_d 0.00162089f $X=3.95 $Y=0.815 $X2=0 $Y2=0
cc_241 N_Y_c_371_n N_VGND_M1014_s 9.55912e-19 $X=4.615 $Y=0.815 $X2=0 $Y2=0
cc_242 N_Y_c_376_n N_VGND_M1014_s 0.00189615f $X=4.782 $Y=0.905 $X2=0 $Y2=0
cc_243 N_Y_c_368_n N_VGND_c_471_n 0.0014523f $X=0.95 $Y=0.815 $X2=0 $Y2=0
cc_244 N_Y_c_380_n N_VGND_c_472_n 0.0226935f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_245 N_Y_c_367_n N_VGND_c_472_n 0.00218853f $X=1.51 $Y=0.815 $X2=0 $Y2=0
cc_246 N_Y_c_367_n N_VGND_c_473_n 0.0122559f $X=1.51 $Y=0.815 $X2=0 $Y2=0
cc_247 N_Y_c_370_n N_VGND_c_474_n 0.0122559f $X=3.95 $Y=0.815 $X2=0 $Y2=0
cc_248 N_Y_c_376_n N_VGND_c_475_n 0.00247473f $X=4.782 $Y=0.905 $X2=0 $Y2=0
cc_249 N_Y_c_371_n N_VGND_c_476_n 0.00727234f $X=4.615 $Y=0.815 $X2=0 $Y2=0
cc_250 N_Y_c_376_n N_VGND_c_476_n 0.0166121f $X=4.782 $Y=0.905 $X2=0 $Y2=0
cc_251 N_Y_c_369_n N_VGND_c_477_n 0.00242888f $X=3.01 $Y=0.815 $X2=0 $Y2=0
cc_252 N_Y_c_398_n N_VGND_c_477_n 0.0226935f $X=3.19 $Y=0.39 $X2=0 $Y2=0
cc_253 N_Y_c_370_n N_VGND_c_477_n 0.00218853f $X=3.95 $Y=0.815 $X2=0 $Y2=0
cc_254 N_Y_c_370_n N_VGND_c_479_n 0.00242888f $X=3.95 $Y=0.815 $X2=0 $Y2=0
cc_255 N_Y_c_406_n N_VGND_c_479_n 0.0226935f $X=4.13 $Y=0.39 $X2=0 $Y2=0
cc_256 N_Y_c_371_n N_VGND_c_479_n 0.00218853f $X=4.615 $Y=0.815 $X2=0 $Y2=0
cc_257 N_Y_c_367_n N_VGND_c_481_n 0.00242888f $X=1.51 $Y=0.815 $X2=0 $Y2=0
cc_258 N_Y_c_390_n N_VGND_c_481_n 0.0226935f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_259 N_Y_c_369_n N_VGND_c_481_n 0.00218853f $X=3.01 $Y=0.815 $X2=0 $Y2=0
cc_260 N_Y_c_369_n N_VGND_c_482_n 0.0567707f $X=3.01 $Y=0.815 $X2=0 $Y2=0
cc_261 N_Y_M1006_d N_VGND_c_483_n 0.00312858f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_262 N_Y_M1007_s N_VGND_c_483_n 0.00291485f $X=1.505 $Y=0.235 $X2=0 $Y2=0
cc_263 N_Y_M1002_s N_VGND_c_483_n 0.00291485f $X=3.005 $Y=0.235 $X2=0 $Y2=0
cc_264 N_Y_M1004_d N_VGND_c_483_n 0.00291485f $X=3.945 $Y=0.235 $X2=0 $Y2=0
cc_265 N_Y_c_380_n N_VGND_c_483_n 0.0144038f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_266 N_Y_c_367_n N_VGND_c_483_n 0.0094091f $X=1.51 $Y=0.815 $X2=0 $Y2=0
cc_267 N_Y_c_390_n N_VGND_c_483_n 0.0144038f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_268 N_Y_c_369_n N_VGND_c_483_n 0.0115297f $X=3.01 $Y=0.815 $X2=0 $Y2=0
cc_269 N_Y_c_398_n N_VGND_c_483_n 0.0144038f $X=3.19 $Y=0.39 $X2=0 $Y2=0
cc_270 N_Y_c_370_n N_VGND_c_483_n 0.0094091f $X=3.95 $Y=0.815 $X2=0 $Y2=0
cc_271 N_Y_c_406_n N_VGND_c_483_n 0.0144038f $X=4.13 $Y=0.39 $X2=0 $Y2=0
cc_272 N_Y_c_371_n N_VGND_c_483_n 0.0045573f $X=4.615 $Y=0.815 $X2=0 $Y2=0
cc_273 N_Y_c_376_n N_VGND_c_483_n 0.00494103f $X=4.782 $Y=0.905 $X2=0 $Y2=0
