* File: sky130_fd_sc_hdll__a32oi_4.pxi.spice
* Created: Thu Aug 27 18:56:38 2020
* 
x_PM_SKY130_FD_SC_HDLL__A32OI_4%B2 N_B2_c_109_n N_B2_M1001_g N_B2_c_102_n
+ N_B2_M1002_g N_B2_c_110_n N_B2_M1012_g N_B2_c_103_n N_B2_M1024_g N_B2_c_111_n
+ N_B2_M1021_g N_B2_c_104_n N_B2_M1025_g N_B2_c_112_n N_B2_M1035_g N_B2_c_105_n
+ N_B2_M1039_g B2 B2 B2 B2 B2 B2 N_B2_c_106_n N_B2_c_107_n N_B2_c_108_n B2 B2
+ PM_SKY130_FD_SC_HDLL__A32OI_4%B2
x_PM_SKY130_FD_SC_HDLL__A32OI_4%B1 N_B1_c_186_n N_B1_M1010_g N_B1_c_192_n
+ N_B1_M1000_g N_B1_c_187_n N_B1_M1017_g N_B1_c_193_n N_B1_M1004_g N_B1_c_188_n
+ N_B1_M1030_g N_B1_c_194_n N_B1_M1009_g N_B1_c_195_n N_B1_M1016_g N_B1_c_189_n
+ N_B1_M1033_g B1 B1 N_B1_c_190_n N_B1_c_191_n B1 B1
+ PM_SKY130_FD_SC_HDLL__A32OI_4%B1
x_PM_SKY130_FD_SC_HDLL__A32OI_4%A1 N_A1_c_270_n N_A1_M1005_g N_A1_c_271_n
+ N_A1_M1011_g N_A1_c_264_n N_A1_M1007_g N_A1_c_272_n N_A1_M1026_g N_A1_c_265_n
+ N_A1_M1013_g N_A1_c_266_n N_A1_M1031_g N_A1_c_273_n N_A1_M1029_g N_A1_c_267_n
+ N_A1_M1034_g A1 A1 A1 A1 N_A1_c_269_n A1 A1 A1
+ PM_SKY130_FD_SC_HDLL__A32OI_4%A1
x_PM_SKY130_FD_SC_HDLL__A32OI_4%A2 N_A2_c_333_n N_A2_M1003_g N_A2_c_339_n
+ N_A2_M1008_g N_A2_c_334_n N_A2_M1018_g N_A2_c_340_n N_A2_M1014_g N_A2_c_335_n
+ N_A2_M1020_g N_A2_c_341_n N_A2_M1019_g N_A2_c_342_n N_A2_M1027_g N_A2_c_336_n
+ N_A2_M1036_g A2 A2 A2 A2 N_A2_c_337_n A2 A2 PM_SKY130_FD_SC_HDLL__A32OI_4%A2
x_PM_SKY130_FD_SC_HDLL__A32OI_4%A3 N_A3_c_400_n N_A3_M1015_g N_A3_c_408_n
+ N_A3_M1006_g N_A3_c_401_n N_A3_M1022_g N_A3_c_409_n N_A3_M1023_g N_A3_c_402_n
+ N_A3_M1037_g N_A3_c_410_n N_A3_M1028_g N_A3_c_411_n N_A3_M1032_g N_A3_c_403_n
+ N_A3_M1038_g A3 A3 A3 A3 A3 N_A3_c_405_n N_A3_c_406_n A3 A3 N_A3_c_407_n
+ PM_SKY130_FD_SC_HDLL__A32OI_4%A3
x_PM_SKY130_FD_SC_HDLL__A32OI_4%A_27_297# N_A_27_297#_M1001_d
+ N_A_27_297#_M1012_d N_A_27_297#_M1035_d N_A_27_297#_M1004_d
+ N_A_27_297#_M1016_d N_A_27_297#_M1011_d N_A_27_297#_M1029_d
+ N_A_27_297#_M1014_d N_A_27_297#_M1027_d N_A_27_297#_M1023_s
+ N_A_27_297#_M1032_s N_A_27_297#_c_478_n N_A_27_297#_c_489_n
+ N_A_27_297#_c_493_n N_A_27_297#_c_490_n N_A_27_297#_c_497_n
+ N_A_27_297#_c_499_n N_A_27_297#_c_503_n N_A_27_297#_c_508_n
+ N_A_27_297#_c_512_n N_A_27_297#_c_514_n N_A_27_297#_c_518_n
+ N_A_27_297#_c_523_n N_A_27_297#_c_527_n N_A_27_297#_c_529_n
+ N_A_27_297#_c_534_n N_A_27_297#_c_504_n N_A_27_297#_c_506_n
+ N_A_27_297#_c_519_n N_A_27_297#_c_521_n N_A_27_297#_c_535_n
+ PM_SKY130_FD_SC_HDLL__A32OI_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A32OI_4%Y N_Y_M1010_s N_Y_M1030_s N_Y_M1007_s
+ N_Y_M1031_s N_Y_M1001_s N_Y_M1021_s N_Y_M1000_s N_Y_M1009_s N_Y_c_607_n
+ N_Y_c_611_n N_Y_c_631_n N_Y_c_603_n N_Y_c_637_n N_Y_c_613_n N_Y_c_619_n
+ N_Y_c_642_n Y Y Y Y N_Y_c_605_n Y PM_SKY130_FD_SC_HDLL__A32OI_4%Y
x_PM_SKY130_FD_SC_HDLL__A32OI_4%VPWR N_VPWR_M1005_s N_VPWR_M1026_s
+ N_VPWR_M1008_s N_VPWR_M1019_s N_VPWR_M1006_d N_VPWR_M1028_d N_VPWR_c_706_n
+ N_VPWR_c_707_n N_VPWR_c_708_n N_VPWR_c_709_n N_VPWR_c_710_n VPWR
+ N_VPWR_c_711_n N_VPWR_c_712_n N_VPWR_c_713_n N_VPWR_c_714_n N_VPWR_c_715_n
+ N_VPWR_c_716_n N_VPWR_c_717_n N_VPWR_c_705_n N_VPWR_c_719_n N_VPWR_c_720_n
+ N_VPWR_c_721_n N_VPWR_c_722_n N_VPWR_c_723_n N_VPWR_c_724_n
+ PM_SKY130_FD_SC_HDLL__A32OI_4%VPWR
x_PM_SKY130_FD_SC_HDLL__A32OI_4%A_27_47# N_A_27_47#_M1002_d N_A_27_47#_M1024_d
+ N_A_27_47#_M1039_d N_A_27_47#_M1017_d N_A_27_47#_M1033_d N_A_27_47#_c_837_n
+ N_A_27_47#_c_838_n N_A_27_47#_c_843_n N_A_27_47#_c_846_n N_A_27_47#_c_847_n
+ N_A_27_47#_c_874_p N_A_27_47#_c_836_n N_A_27_47#_c_851_n
+ PM_SKY130_FD_SC_HDLL__A32OI_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__A32OI_4%VGND N_VGND_M1002_s N_VGND_M1025_s
+ N_VGND_M1015_s N_VGND_M1022_s N_VGND_M1038_s N_VGND_c_892_n VGND
+ N_VGND_c_893_n N_VGND_c_894_n N_VGND_c_895_n N_VGND_c_896_n N_VGND_c_897_n
+ N_VGND_c_898_n N_VGND_c_899_n N_VGND_c_900_n N_VGND_c_901_n N_VGND_c_902_n
+ N_VGND_c_903_n PM_SKY130_FD_SC_HDLL__A32OI_4%VGND
x_PM_SKY130_FD_SC_HDLL__A32OI_4%A_893_47# N_A_893_47#_M1007_d
+ N_A_893_47#_M1013_d N_A_893_47#_M1034_d N_A_893_47#_M1018_d
+ N_A_893_47#_M1036_d N_A_893_47#_c_1023_n
+ PM_SKY130_FD_SC_HDLL__A32OI_4%A_893_47#
x_PM_SKY130_FD_SC_HDLL__A32OI_4%A_1379_47# N_A_1379_47#_M1003_s
+ N_A_1379_47#_M1020_s N_A_1379_47#_M1015_d N_A_1379_47#_M1037_d
+ N_A_1379_47#_c_1052_n N_A_1379_47#_c_1063_n N_A_1379_47#_c_1064_n
+ N_A_1379_47#_c_1069_n N_A_1379_47#_c_1071_n
+ PM_SKY130_FD_SC_HDLL__A32OI_4%A_1379_47#
cc_1 VNB N_B2_c_102_n 0.0219558f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB N_B2_c_103_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB N_B2_c_104_n 0.0163871f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_4 VNB N_B2_c_105_n 0.0166494f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_5 VNB N_B2_c_106_n 0.0263946f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.165
cc_6 VNB N_B2_c_107_n 0.0720805f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_7 VNB N_B2_c_108_n 0.00936732f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.305
cc_8 VNB N_B1_c_186_n 0.0161073f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_9 VNB N_B1_c_187_n 0.0169334f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_10 VNB N_B1_c_188_n 0.0174137f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_11 VNB N_B1_c_189_n 0.0229091f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_12 VNB N_B1_c_190_n 0.00328581f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_13 VNB N_B1_c_191_n 0.0730516f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A1_c_264_n 0.022465f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_15 VNB N_A1_c_265_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_16 VNB N_A1_c_266_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_17 VNB N_A1_c_267_n 0.0188029f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_18 VNB A1 0.00147415f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.105
cc_19 VNB N_A1_c_269_n 0.108629f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.202
cc_20 VNB N_A2_c_333_n 0.0179218f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_21 VNB N_A2_c_334_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_22 VNB N_A2_c_335_n 0.0174167f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_23 VNB N_A2_c_336_n 0.0241689f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_24 VNB N_A2_c_337_n 0.0805231f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.202
cc_25 VNB A2 0.00982743f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A3_c_400_n 0.0215708f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_27 VNB N_A3_c_401_n 0.0167427f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_28 VNB N_A3_c_402_n 0.0171787f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_29 VNB N_A3_c_403_n 0.0189425f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_30 VNB A3 0.00598505f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_31 VNB N_A3_c_405_n 0.103647f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.202
cc_32 VNB N_A3_c_406_n 0.00332226f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.305
cc_33 VNB N_A3_c_407_n 0.00834913f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=1.19
cc_34 VNB N_Y_c_603_n 0.00881835f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.165
cc_35 VNB Y 0.00384158f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_Y_c_605_n 0.00100529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_705_n 0.478484f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_27_47#_c_836_n 0.00234081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_892_n 0.00551967f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_40 VNB N_VGND_c_893_n 0.0151574f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_41 VNB N_VGND_c_894_n 0.0134288f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_42 VNB N_VGND_c_895_n 0.164929f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_896_n 0.0123546f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_44 VNB N_VGND_c_897_n 0.0134624f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=1.16
cc_45 VNB N_VGND_c_898_n 0.00792095f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.53
cc_46 VNB N_VGND_c_899_n 0.00849831f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_47 VNB N_VGND_c_900_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=1.19
cc_48 VNB N_VGND_c_901_n 0.00537227f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_902_n 0.0350712f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_903_n 0.545272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_893_47#_c_1023_n 0.00444027f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_52 VNB N_A_1379_47#_c_1052_n 0.0140526f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_53 VPB N_B2_c_109_n 0.01915f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_54 VPB N_B2_c_110_n 0.0162612f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_55 VPB N_B2_c_111_n 0.0162625f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_56 VPB N_B2_c_112_n 0.0164246f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_57 VPB B2 0.0257344f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_58 VPB N_B2_c_106_n 0.00944663f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.165
cc_59 VPB N_B2_c_107_n 0.0474397f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_60 VPB N_B1_c_192_n 0.0156532f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_61 VPB N_B1_c_193_n 0.0162424f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_62 VPB N_B1_c_194_n 0.0162621f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.995
cc_63 VPB N_B1_c_195_n 0.0166003f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_64 VPB N_B1_c_190_n 0.00230149f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_65 VPB N_B1_c_191_n 0.0463185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A1_c_270_n 0.0161497f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_67 VPB N_A1_c_271_n 0.0160921f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_68 VPB N_A1_c_272_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_69 VPB N_A1_c_273_n 0.0227977f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_70 VPB N_A1_c_269_n 0.0679469f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.202
cc_71 VPB N_A2_c_339_n 0.0175227f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_72 VPB N_A2_c_340_n 0.0160921f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_73 VPB N_A2_c_341_n 0.0158129f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.995
cc_74 VPB N_A2_c_342_n 0.0209165f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_75 VPB N_A2_c_337_n 0.050339f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.202
cc_76 VPB N_A3_c_408_n 0.0206372f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_77 VPB N_A3_c_409_n 0.0160921f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_78 VPB N_A3_c_410_n 0.0158129f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.995
cc_79 VPB N_A3_c_411_n 0.0209165f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_80 VPB N_A3_c_405_n 0.0618209f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.202
cc_81 VPB N_A_27_297#_c_478_n 0.00821562f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB Y 0.00363513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_706_n 4.17955e-19 $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_84 VPB N_VPWR_c_707_n 4.04661e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_85 VPB N_VPWR_c_708_n 4.04661e-19 $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_86 VPB N_VPWR_c_709_n 4.04661e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_710_n 4.04661e-19 $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.165
cc_88 VPB N_VPWR_c_711_n 0.10295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_712_n 0.0178661f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=1.202
cc_90 VPB N_VPWR_c_713_n 0.0235941f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_91 VPB N_VPWR_c_714_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.87
cc_92 VPB N_VPWR_c_715_n 0.03063f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.19
cc_93 VPB N_VPWR_c_716_n 0.0140826f $X=-0.19 $Y=1.305 $X2=1.61 $Y2=1.19
cc_94 VPB N_VPWR_c_717_n 0.0286331f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_705_n 0.0619708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_719_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_720_n 0.0210912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_721_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_722_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_723_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_724_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 N_B2_c_105_n N_B1_c_186_n 0.0215202f $X=1.93 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_103 N_B2_c_112_n N_B1_c_192_n 0.03651f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_104 N_B2_c_107_n N_B1_c_191_n 0.0215202f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_105 B2 N_B1_c_191_n 2.14426e-19 $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_106 B2 N_A_27_297#_M1001_d 0.0121575f $X=0.15 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_107 N_B2_c_109_n N_A_27_297#_c_478_n 0.0125689f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_108 N_B2_c_110_n N_A_27_297#_c_478_n 0.0110013f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_109 N_B2_c_111_n N_A_27_297#_c_478_n 0.0104321f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_110 N_B2_c_112_n N_A_27_297#_c_478_n 0.0110013f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_111 B2 N_A_27_297#_c_478_n 0.0106869f $X=0.15 $Y=1.445 $X2=0 $Y2=0
cc_112 N_B2_c_110_n N_Y_c_607_n 0.0123803f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_113 N_B2_c_111_n N_Y_c_607_n 0.00899481f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_114 N_B2_c_107_n N_Y_c_607_n 0.005986f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_115 B2 N_Y_c_607_n 0.0246069f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_116 N_B2_c_112_n N_Y_c_611_n 0.0137815f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_117 B2 N_Y_c_611_n 0.00311671f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_118 N_B2_c_109_n N_Y_c_613_n 0.0137867f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_119 N_B2_c_110_n N_Y_c_613_n 0.00766271f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_120 N_B2_c_111_n N_Y_c_613_n 0.00105163f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_121 B2 N_Y_c_613_n 0.0277972f $X=0.15 $Y=1.445 $X2=0 $Y2=0
cc_122 N_B2_c_107_n N_Y_c_613_n 0.00613621f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_123 B2 N_Y_c_613_n 0.0170672f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_124 N_B2_c_110_n N_Y_c_619_n 0.00116208f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_125 N_B2_c_111_n N_Y_c_619_n 0.0112429f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_126 N_B2_c_112_n N_Y_c_619_n 0.00627445f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_127 N_B2_c_107_n N_Y_c_619_n 0.00613621f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_128 B2 N_Y_c_619_n 0.0170672f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_129 N_B2_c_112_n Y 0.00408716f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_130 N_B2_c_105_n Y 0.0034652f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_131 N_B2_c_107_n Y 0.0034652f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_132 B2 Y 0.0136023f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_133 N_B2_c_112_n Y 0.00319402f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_134 N_B2_c_105_n N_Y_c_605_n 9.14188e-19 $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_135 N_B2_c_109_n N_VPWR_c_711_n 0.00439333f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_136 N_B2_c_110_n N_VPWR_c_711_n 0.00439333f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_137 N_B2_c_111_n N_VPWR_c_711_n 0.00439333f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_138 N_B2_c_112_n N_VPWR_c_711_n 0.00439333f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_139 N_B2_c_109_n N_VPWR_c_705_n 0.00699435f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_140 N_B2_c_110_n N_VPWR_c_705_n 0.00608292f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_141 N_B2_c_111_n N_VPWR_c_705_n 0.00608292f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_142 N_B2_c_112_n N_VPWR_c_705_n 0.00610813f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_143 N_B2_c_102_n N_A_27_47#_c_837_n 0.00405771f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_144 N_B2_c_102_n N_A_27_47#_c_838_n 0.0132138f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_145 N_B2_c_103_n N_A_27_47#_c_838_n 0.0129187f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_146 N_B2_c_106_n N_A_27_47#_c_838_n 0.00214654f $X=0.395 $Y=1.165 $X2=0 $Y2=0
cc_147 N_B2_c_107_n N_A_27_47#_c_838_n 0.00322095f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_148 B2 N_A_27_47#_c_838_n 0.0322963f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_149 N_B2_c_106_n N_A_27_47#_c_843_n 0.00381493f $X=0.395 $Y=1.165 $X2=0 $Y2=0
cc_150 N_B2_c_108_n N_A_27_47#_c_843_n 0.00931784f $X=0.22 $Y=1.305 $X2=0 $Y2=0
cc_151 B2 N_A_27_47#_c_843_n 8.08679e-19 $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_152 N_B2_c_104_n N_A_27_47#_c_846_n 0.00377939f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_153 N_B2_c_104_n N_A_27_47#_c_847_n 0.0120987f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_154 N_B2_c_105_n N_A_27_47#_c_847_n 0.0147393f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_155 N_B2_c_107_n N_A_27_47#_c_847_n 0.00344781f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_156 B2 N_A_27_47#_c_847_n 0.0260597f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_157 N_B2_c_107_n N_A_27_47#_c_851_n 0.00312289f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_158 B2 N_A_27_47#_c_851_n 0.0092175f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_159 N_B2_c_102_n N_VGND_c_893_n 0.00198377f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_160 N_B2_c_103_n N_VGND_c_894_n 0.00425094f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_161 N_B2_c_104_n N_VGND_c_894_n 0.00198377f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_162 N_B2_c_105_n N_VGND_c_895_n 0.00425094f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_163 N_B2_c_102_n N_VGND_c_898_n 0.0112154f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_164 N_B2_c_103_n N_VGND_c_898_n 0.00162962f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_165 N_B2_c_103_n N_VGND_c_899_n 5.64511e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_166 N_B2_c_104_n N_VGND_c_899_n 0.00960147f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_167 N_B2_c_105_n N_VGND_c_899_n 0.00317372f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_168 N_B2_c_102_n N_VGND_c_903_n 0.00358947f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_169 N_B2_c_103_n N_VGND_c_903_n 0.00584696f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_170 N_B2_c_104_n N_VGND_c_903_n 0.00271758f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_171 N_B2_c_105_n N_VGND_c_903_n 0.00579121f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B1_c_195_n N_A1_c_270_n 0.0309206f $X=3.785 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_173 N_B1_c_190_n A1 0.015263f $X=3.7 $Y=1.16 $X2=0 $Y2=0
cc_174 N_B1_c_191_n A1 2.33231e-19 $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_175 N_B1_c_190_n N_A1_c_269_n 0.0041816f $X=3.7 $Y=1.16 $X2=0 $Y2=0
cc_176 N_B1_c_191_n N_A1_c_269_n 0.0190036f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_177 N_B1_c_192_n N_A_27_297#_c_478_n 0.00920483f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_178 N_B1_c_193_n N_A_27_297#_c_478_n 0.0110013f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_179 N_B1_c_194_n N_A_27_297#_c_478_n 0.010389f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_180 N_B1_c_195_n N_A_27_297#_c_478_n 0.014098f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_181 N_B1_c_195_n N_A_27_297#_c_489_n 0.00600033f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_182 N_B1_c_195_n N_A_27_297#_c_490_n 0.00163f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_183 N_B1_c_190_n N_A_27_297#_c_490_n 0.00131284f $X=3.7 $Y=1.16 $X2=0 $Y2=0
cc_184 N_B1_c_192_n N_Y_c_611_n 2.31742e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_185 N_B1_c_186_n N_Y_c_631_n 0.00217694f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_186 N_B1_c_187_n N_Y_c_603_n 0.0114045f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_187 N_B1_c_188_n N_Y_c_603_n 0.0087742f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_188 N_B1_c_189_n N_Y_c_603_n 0.010581f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_189 N_B1_c_190_n N_Y_c_603_n 0.0657163f $X=3.7 $Y=1.16 $X2=0 $Y2=0
cc_190 N_B1_c_191_n N_Y_c_603_n 0.00875686f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_191 N_B1_c_193_n N_Y_c_637_n 0.0134376f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_192 N_B1_c_194_n N_Y_c_637_n 0.00938864f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_193 N_B1_c_190_n N_Y_c_637_n 0.0238259f $X=3.7 $Y=1.16 $X2=0 $Y2=0
cc_194 N_B1_c_191_n N_Y_c_637_n 0.00595224f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_195 N_B1_c_192_n N_Y_c_619_n 3.03958e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_196 N_B1_c_193_n N_Y_c_642_n 0.00116208f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_197 N_B1_c_194_n N_Y_c_642_n 0.0111902f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_198 N_B1_c_195_n N_Y_c_642_n 0.00652611f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_199 N_B1_c_190_n N_Y_c_642_n 0.0186876f $X=3.7 $Y=1.16 $X2=0 $Y2=0
cc_200 N_B1_c_191_n N_Y_c_642_n 0.00591164f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_201 N_B1_c_186_n Y 0.00330483f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_202 N_B1_c_192_n Y 0.00438448f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_203 N_B1_c_193_n Y 0.00393734f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_204 N_B1_c_190_n Y 0.021702f $X=3.7 $Y=1.16 $X2=0 $Y2=0
cc_205 N_B1_c_191_n Y 0.0286604f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_206 N_B1_c_192_n Y 0.0145125f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_207 N_B1_c_193_n Y 0.00823589f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_208 N_B1_c_194_n Y 0.00104879f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_209 N_B1_c_191_n Y 0.00444485f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_210 N_B1_c_186_n N_Y_c_605_n 0.00421096f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_211 N_B1_c_187_n N_Y_c_605_n 0.00407254f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_212 N_B1_c_195_n N_VPWR_c_706_n 0.00125028f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_213 N_B1_c_192_n N_VPWR_c_711_n 0.00439333f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_214 N_B1_c_193_n N_VPWR_c_711_n 0.00439333f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_215 N_B1_c_194_n N_VPWR_c_711_n 0.00439333f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_216 N_B1_c_195_n N_VPWR_c_711_n 0.00439333f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_217 N_B1_c_192_n N_VPWR_c_705_n 0.00610813f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_218 N_B1_c_193_n N_VPWR_c_705_n 0.00608292f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_219 N_B1_c_194_n N_VPWR_c_705_n 0.00608292f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_220 N_B1_c_195_n N_VPWR_c_705_n 0.00619886f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_221 N_B1_c_186_n N_A_27_47#_c_836_n 0.00958023f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_222 N_B1_c_187_n N_A_27_47#_c_836_n 0.00813248f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_223 N_B1_c_188_n N_A_27_47#_c_836_n 0.00844662f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_224 N_B1_c_189_n N_A_27_47#_c_836_n 0.00844662f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_225 N_B1_c_191_n N_A_27_47#_c_836_n 3.86154e-19 $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_226 N_B1_c_186_n N_VGND_c_895_n 0.00366111f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_227 N_B1_c_187_n N_VGND_c_895_n 0.00366111f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_228 N_B1_c_188_n N_VGND_c_895_n 0.00366111f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_229 N_B1_c_189_n N_VGND_c_895_n 0.00366111f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_230 N_B1_c_186_n N_VGND_c_903_n 0.00543917f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_231 N_B1_c_187_n N_VGND_c_903_n 0.00549891f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_232 N_B1_c_188_n N_VGND_c_903_n 0.00561869f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_233 N_B1_c_189_n N_VGND_c_903_n 0.00681779f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A1_c_267_n N_A2_c_333_n 0.0170727f $X=6.26 $Y=1.01 $X2=-0.19 $Y2=-0.24
cc_235 N_A1_c_273_n N_A2_c_339_n 0.0169064f $X=6.14 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A1_c_269_n N_A2_c_337_n 0.0198396f $X=6.14 $Y=1.202 $X2=0 $Y2=0
cc_237 A1 A2 0.00547493f $X=5.69 $Y=1.105 $X2=0 $Y2=0
cc_238 N_A1_c_269_n A2 0.0011957f $X=6.14 $Y=1.202 $X2=0 $Y2=0
cc_239 N_A1_c_270_n N_A_27_297#_c_489_n 0.00567952f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_240 N_A1_c_270_n N_A_27_297#_c_493_n 0.0157734f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_241 N_A1_c_271_n N_A_27_297#_c_493_n 0.0176505f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_242 A1 N_A_27_297#_c_493_n 0.0287231f $X=5.69 $Y=1.105 $X2=0 $Y2=0
cc_243 N_A1_c_269_n N_A_27_297#_c_493_n 0.00574723f $X=6.14 $Y=1.202 $X2=0 $Y2=0
cc_244 N_A1_c_271_n N_A_27_297#_c_497_n 0.00530373f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_245 N_A1_c_272_n N_A_27_297#_c_497_n 0.00557226f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_246 N_A1_c_272_n N_A_27_297#_c_499_n 0.0202314f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_247 N_A1_c_273_n N_A_27_297#_c_499_n 0.0254294f $X=6.14 $Y=1.41 $X2=0 $Y2=0
cc_248 A1 N_A_27_297#_c_499_n 0.0426246f $X=5.69 $Y=1.105 $X2=0 $Y2=0
cc_249 N_A1_c_269_n N_A_27_297#_c_499_n 0.0176371f $X=6.14 $Y=1.202 $X2=0 $Y2=0
cc_250 N_A1_c_273_n N_A_27_297#_c_503_n 0.00559194f $X=6.14 $Y=1.41 $X2=0 $Y2=0
cc_251 A1 N_A_27_297#_c_504_n 0.00903496f $X=5.69 $Y=1.105 $X2=0 $Y2=0
cc_252 N_A1_c_269_n N_A_27_297#_c_504_n 0.00443401f $X=6.14 $Y=1.202 $X2=0 $Y2=0
cc_253 N_A1_c_269_n N_A_27_297#_c_506_n 0.00199819f $X=6.14 $Y=1.202 $X2=0 $Y2=0
cc_254 N_A1_c_264_n N_Y_c_603_n 0.0110355f $X=4.85 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A1_c_265_n N_Y_c_603_n 0.00922871f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_256 N_A1_c_266_n N_Y_c_603_n 0.00922871f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_257 A1 N_Y_c_603_n 0.0849667f $X=5.69 $Y=1.105 $X2=0 $Y2=0
cc_258 N_A1_c_269_n N_Y_c_603_n 0.0252705f $X=6.14 $Y=1.202 $X2=0 $Y2=0
cc_259 N_A1_c_270_n N_Y_c_642_n 2.26437e-19 $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A1_c_270_n N_VPWR_c_706_n 0.0158902f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A1_c_271_n N_VPWR_c_706_n 0.0109404f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A1_c_272_n N_VPWR_c_706_n 6.26289e-19 $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A1_c_273_n N_VPWR_c_707_n 9.90794e-19 $X=6.14 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A1_c_270_n N_VPWR_c_711_n 0.00427505f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A1_c_271_n N_VPWR_c_712_n 0.00622633f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A1_c_272_n N_VPWR_c_712_n 0.00702461f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_267 N_A1_c_273_n N_VPWR_c_713_n 0.00702461f $X=6.14 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A1_c_270_n N_VPWR_c_705_n 0.00748259f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A1_c_271_n N_VPWR_c_705_n 0.0104011f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_270 N_A1_c_272_n N_VPWR_c_705_n 0.013679f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_271 N_A1_c_273_n N_VPWR_c_705_n 0.014276f $X=6.14 $Y=1.41 $X2=0 $Y2=0
cc_272 N_A1_c_272_n N_VPWR_c_720_n 0.00362675f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_273 N_A1_c_273_n N_VPWR_c_720_n 0.0171741f $X=6.14 $Y=1.41 $X2=0 $Y2=0
cc_274 N_A1_c_264_n N_VGND_c_895_n 0.00366111f $X=4.85 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A1_c_265_n N_VGND_c_895_n 0.00366111f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_276 N_A1_c_266_n N_VGND_c_895_n 0.00366111f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_277 N_A1_c_267_n N_VGND_c_895_n 0.00366111f $X=6.26 $Y=1.01 $X2=0 $Y2=0
cc_278 N_A1_c_264_n N_VGND_c_903_n 0.00669801f $X=4.85 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A1_c_265_n N_VGND_c_903_n 0.00549891f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_280 N_A1_c_266_n N_VGND_c_903_n 0.00549891f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_281 N_A1_c_267_n N_VGND_c_903_n 0.00570488f $X=6.26 $Y=1.01 $X2=0 $Y2=0
cc_282 N_A1_c_264_n N_A_893_47#_c_1023_n 0.00818766f $X=4.85 $Y=0.995 $X2=0
+ $Y2=0
cc_283 N_A1_c_265_n N_A_893_47#_c_1023_n 0.00818766f $X=5.32 $Y=0.995 $X2=0
+ $Y2=0
cc_284 N_A1_c_266_n N_A_893_47#_c_1023_n 0.00818766f $X=5.79 $Y=0.995 $X2=0
+ $Y2=0
cc_285 N_A1_c_267_n N_A_893_47#_c_1023_n 0.0127383f $X=6.26 $Y=1.01 $X2=0 $Y2=0
cc_286 N_A1_c_267_n N_A_1379_47#_c_1052_n 7.71295e-19 $X=6.26 $Y=1.01 $X2=0
+ $Y2=0
cc_287 A2 N_A3_c_405_n 0.00189259f $X=8.455 $Y=1.19 $X2=0 $Y2=0
cc_288 A2 N_A3_c_406_n 0.00693886f $X=8.455 $Y=1.19 $X2=0 $Y2=0
cc_289 N_A2_c_339_n N_A_27_297#_c_503_n 0.00805067f $X=6.845 $Y=1.41 $X2=0 $Y2=0
cc_290 N_A2_c_339_n N_A_27_297#_c_508_n 0.0169991f $X=6.845 $Y=1.41 $X2=0 $Y2=0
cc_291 N_A2_c_340_n N_A_27_297#_c_508_n 0.0175543f $X=7.315 $Y=1.41 $X2=0 $Y2=0
cc_292 N_A2_c_337_n N_A_27_297#_c_508_n 0.0061683f $X=8.255 $Y=1.202 $X2=0 $Y2=0
cc_293 A2 N_A_27_297#_c_508_n 0.0301395f $X=8.455 $Y=1.19 $X2=0 $Y2=0
cc_294 N_A2_c_340_n N_A_27_297#_c_512_n 0.00530373f $X=7.315 $Y=1.41 $X2=0 $Y2=0
cc_295 N_A2_c_341_n N_A_27_297#_c_512_n 0.00490547f $X=7.785 $Y=1.41 $X2=0 $Y2=0
cc_296 N_A2_c_341_n N_A_27_297#_c_514_n 0.0160251f $X=7.785 $Y=1.41 $X2=0 $Y2=0
cc_297 N_A2_c_342_n N_A_27_297#_c_514_n 0.0195541f $X=8.255 $Y=1.41 $X2=0 $Y2=0
cc_298 N_A2_c_337_n N_A_27_297#_c_514_n 0.00596011f $X=8.255 $Y=1.202 $X2=0
+ $Y2=0
cc_299 A2 N_A_27_297#_c_514_n 0.0315459f $X=8.455 $Y=1.19 $X2=0 $Y2=0
cc_300 N_A2_c_342_n N_A_27_297#_c_518_n 0.00561135f $X=8.255 $Y=1.41 $X2=0 $Y2=0
cc_301 N_A2_c_337_n N_A_27_297#_c_519_n 0.00412388f $X=8.255 $Y=1.202 $X2=0
+ $Y2=0
cc_302 A2 N_A_27_297#_c_519_n 0.00945295f $X=8.455 $Y=1.19 $X2=0 $Y2=0
cc_303 A2 N_A_27_297#_c_521_n 0.00835061f $X=8.455 $Y=1.19 $X2=0 $Y2=0
cc_304 N_A2_c_339_n N_VPWR_c_707_n 0.018551f $X=6.845 $Y=1.41 $X2=0 $Y2=0
cc_305 N_A2_c_340_n N_VPWR_c_707_n 0.0107665f $X=7.315 $Y=1.41 $X2=0 $Y2=0
cc_306 N_A2_c_341_n N_VPWR_c_707_n 5.96427e-19 $X=7.785 $Y=1.41 $X2=0 $Y2=0
cc_307 N_A2_c_340_n N_VPWR_c_708_n 6.33692e-19 $X=7.315 $Y=1.41 $X2=0 $Y2=0
cc_308 N_A2_c_341_n N_VPWR_c_708_n 0.0170578f $X=7.785 $Y=1.41 $X2=0 $Y2=0
cc_309 N_A2_c_342_n N_VPWR_c_708_n 0.0154308f $X=8.255 $Y=1.41 $X2=0 $Y2=0
cc_310 N_A2_c_339_n N_VPWR_c_713_n 0.00427505f $X=6.845 $Y=1.41 $X2=0 $Y2=0
cc_311 N_A2_c_340_n N_VPWR_c_714_n 0.00622633f $X=7.315 $Y=1.41 $X2=0 $Y2=0
cc_312 N_A2_c_341_n N_VPWR_c_714_n 0.00427505f $X=7.785 $Y=1.41 $X2=0 $Y2=0
cc_313 N_A2_c_342_n N_VPWR_c_715_n 0.00622633f $X=8.255 $Y=1.41 $X2=0 $Y2=0
cc_314 N_A2_c_339_n N_VPWR_c_705_n 0.00790874f $X=6.845 $Y=1.41 $X2=0 $Y2=0
cc_315 N_A2_c_340_n N_VPWR_c_705_n 0.0104011f $X=7.315 $Y=1.41 $X2=0 $Y2=0
cc_316 N_A2_c_341_n N_VPWR_c_705_n 0.00732977f $X=7.785 $Y=1.41 $X2=0 $Y2=0
cc_317 N_A2_c_342_n N_VPWR_c_705_n 0.0116835f $X=8.255 $Y=1.41 $X2=0 $Y2=0
cc_318 N_A2_c_336_n N_VGND_c_892_n 0.00294182f $X=8.28 $Y=1.01 $X2=0 $Y2=0
cc_319 N_A2_c_333_n N_VGND_c_895_n 0.00366111f $X=6.82 $Y=0.995 $X2=0 $Y2=0
cc_320 N_A2_c_334_n N_VGND_c_895_n 0.00366111f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_321 N_A2_c_335_n N_VGND_c_895_n 0.00366111f $X=7.76 $Y=0.995 $X2=0 $Y2=0
cc_322 N_A2_c_336_n N_VGND_c_895_n 0.00366111f $X=8.28 $Y=1.01 $X2=0 $Y2=0
cc_323 N_A2_c_333_n N_VGND_c_903_n 0.00575667f $X=6.82 $Y=0.995 $X2=0 $Y2=0
cc_324 N_A2_c_334_n N_VGND_c_903_n 0.00549891f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_325 N_A2_c_335_n N_VGND_c_903_n 0.00561869f $X=7.76 $Y=0.995 $X2=0 $Y2=0
cc_326 N_A2_c_336_n N_VGND_c_903_n 0.00681779f $X=8.28 $Y=1.01 $X2=0 $Y2=0
cc_327 N_A2_c_333_n N_A_893_47#_c_1023_n 0.0125017f $X=6.82 $Y=0.995 $X2=0 $Y2=0
cc_328 N_A2_c_334_n N_A_893_47#_c_1023_n 0.00818766f $X=7.29 $Y=0.995 $X2=0
+ $Y2=0
cc_329 N_A2_c_335_n N_A_893_47#_c_1023_n 0.00844662f $X=7.76 $Y=0.995 $X2=0
+ $Y2=0
cc_330 N_A2_c_336_n N_A_893_47#_c_1023_n 0.00844662f $X=8.28 $Y=1.01 $X2=0 $Y2=0
cc_331 A2 N_A_893_47#_c_1023_n 0.00288497f $X=8.455 $Y=1.19 $X2=0 $Y2=0
cc_332 N_A2_c_333_n N_A_1379_47#_c_1052_n 0.00463711f $X=6.82 $Y=0.995 $X2=0
+ $Y2=0
cc_333 N_A2_c_334_n N_A_1379_47#_c_1052_n 0.00922871f $X=7.29 $Y=0.995 $X2=0
+ $Y2=0
cc_334 N_A2_c_335_n N_A_1379_47#_c_1052_n 0.00922871f $X=7.76 $Y=0.995 $X2=0
+ $Y2=0
cc_335 N_A2_c_336_n N_A_1379_47#_c_1052_n 0.0110355f $X=8.28 $Y=1.01 $X2=0 $Y2=0
cc_336 N_A2_c_337_n N_A_1379_47#_c_1052_n 0.0108232f $X=8.255 $Y=1.202 $X2=0
+ $Y2=0
cc_337 A2 N_A_1379_47#_c_1052_n 0.0736794f $X=8.455 $Y=1.19 $X2=0 $Y2=0
cc_338 N_A3_c_408_n N_A_27_297#_c_518_n 0.016418f $X=9.245 $Y=1.41 $X2=0 $Y2=0
cc_339 N_A3_c_408_n N_A_27_297#_c_523_n 0.0181528f $X=9.245 $Y=1.41 $X2=0 $Y2=0
cc_340 N_A3_c_409_n N_A_27_297#_c_523_n 0.0176821f $X=9.715 $Y=1.41 $X2=0 $Y2=0
cc_341 N_A3_c_405_n N_A_27_297#_c_523_n 0.0060275f $X=10.68 $Y=1.202 $X2=0 $Y2=0
cc_342 N_A3_c_406_n N_A_27_297#_c_523_n 0.0282764f $X=10.755 $Y=1.177 $X2=0
+ $Y2=0
cc_343 N_A3_c_409_n N_A_27_297#_c_527_n 0.00530373f $X=9.715 $Y=1.41 $X2=0 $Y2=0
cc_344 N_A3_c_410_n N_A_27_297#_c_527_n 0.00490547f $X=10.185 $Y=1.41 $X2=0
+ $Y2=0
cc_345 N_A3_c_410_n N_A_27_297#_c_529_n 0.0161099f $X=10.185 $Y=1.41 $X2=0 $Y2=0
cc_346 N_A3_c_411_n N_A_27_297#_c_529_n 0.018798f $X=10.655 $Y=1.41 $X2=0 $Y2=0
cc_347 N_A3_c_405_n N_A_27_297#_c_529_n 0.00955388f $X=10.68 $Y=1.202 $X2=0
+ $Y2=0
cc_348 N_A3_c_406_n N_A_27_297#_c_529_n 0.028254f $X=10.755 $Y=1.177 $X2=0 $Y2=0
cc_349 N_A3_c_407_n N_A_27_297#_c_529_n 0.00952377f $X=10.895 $Y=1.075 $X2=0
+ $Y2=0
cc_350 N_A3_c_411_n N_A_27_297#_c_534_n 0.00561135f $X=10.655 $Y=1.41 $X2=0
+ $Y2=0
cc_351 N_A3_c_405_n N_A_27_297#_c_535_n 0.00403737f $X=10.68 $Y=1.202 $X2=0
+ $Y2=0
cc_352 N_A3_c_406_n N_A_27_297#_c_535_n 0.00890343f $X=10.755 $Y=1.177 $X2=0
+ $Y2=0
cc_353 N_A3_c_408_n N_VPWR_c_709_n 0.0344287f $X=9.245 $Y=1.41 $X2=0 $Y2=0
cc_354 N_A3_c_409_n N_VPWR_c_709_n 0.0107665f $X=9.715 $Y=1.41 $X2=0 $Y2=0
cc_355 N_A3_c_410_n N_VPWR_c_709_n 5.96427e-19 $X=10.185 $Y=1.41 $X2=0 $Y2=0
cc_356 N_A3_c_409_n N_VPWR_c_710_n 6.33692e-19 $X=9.715 $Y=1.41 $X2=0 $Y2=0
cc_357 N_A3_c_410_n N_VPWR_c_710_n 0.0141913f $X=10.185 $Y=1.41 $X2=0 $Y2=0
cc_358 N_A3_c_411_n N_VPWR_c_710_n 0.0125643f $X=10.655 $Y=1.41 $X2=0 $Y2=0
cc_359 N_A3_c_408_n N_VPWR_c_715_n 0.00427505f $X=9.245 $Y=1.41 $X2=0 $Y2=0
cc_360 N_A3_c_409_n N_VPWR_c_716_n 0.00622633f $X=9.715 $Y=1.41 $X2=0 $Y2=0
cc_361 N_A3_c_410_n N_VPWR_c_716_n 0.00427505f $X=10.185 $Y=1.41 $X2=0 $Y2=0
cc_362 N_A3_c_411_n N_VPWR_c_717_n 0.00622633f $X=10.655 $Y=1.41 $X2=0 $Y2=0
cc_363 N_A3_c_408_n N_VPWR_c_705_n 0.00873932f $X=9.245 $Y=1.41 $X2=0 $Y2=0
cc_364 N_A3_c_409_n N_VPWR_c_705_n 0.0104011f $X=9.715 $Y=1.41 $X2=0 $Y2=0
cc_365 N_A3_c_410_n N_VPWR_c_705_n 0.00732977f $X=10.185 $Y=1.41 $X2=0 $Y2=0
cc_366 N_A3_c_411_n N_VPWR_c_705_n 0.0116835f $X=10.655 $Y=1.41 $X2=0 $Y2=0
cc_367 A3 N_VGND_M1038_s 0.0092806f $X=10.765 $Y=0.765 $X2=0 $Y2=0
cc_368 N_A3_c_400_n N_VGND_c_892_n 0.00812954f $X=9.22 $Y=0.995 $X2=0 $Y2=0
cc_369 N_A3_c_401_n N_VGND_c_892_n 5.10336e-19 $X=9.69 $Y=0.995 $X2=0 $Y2=0
cc_370 N_A3_c_400_n N_VGND_c_896_n 0.00339367f $X=9.22 $Y=0.995 $X2=0 $Y2=0
cc_371 N_A3_c_401_n N_VGND_c_896_n 0.00340075f $X=9.69 $Y=0.995 $X2=0 $Y2=0
cc_372 N_A3_c_402_n N_VGND_c_897_n 0.00340075f $X=10.16 $Y=0.995 $X2=0 $Y2=0
cc_373 N_A3_c_403_n N_VGND_c_897_n 0.00312205f $X=10.68 $Y=0.995 $X2=0 $Y2=0
cc_374 N_A3_c_400_n N_VGND_c_901_n 4.98468e-19 $X=9.22 $Y=0.995 $X2=0 $Y2=0
cc_375 N_A3_c_401_n N_VGND_c_901_n 0.00701096f $X=9.69 $Y=0.995 $X2=0 $Y2=0
cc_376 N_A3_c_402_n N_VGND_c_901_n 0.00730174f $X=10.16 $Y=0.995 $X2=0 $Y2=0
cc_377 N_A3_c_403_n N_VGND_c_901_n 4.81687e-19 $X=10.68 $Y=0.995 $X2=0 $Y2=0
cc_378 N_A3_c_402_n N_VGND_c_902_n 5.20018e-19 $X=10.16 $Y=0.995 $X2=0 $Y2=0
cc_379 N_A3_c_403_n N_VGND_c_902_n 0.0113014f $X=10.68 $Y=0.995 $X2=0 $Y2=0
cc_380 A3 N_VGND_c_902_n 0.0116947f $X=10.765 $Y=0.765 $X2=0 $Y2=0
cc_381 N_A3_c_405_n N_VGND_c_902_n 0.0011054f $X=10.68 $Y=1.202 $X2=0 $Y2=0
cc_382 N_A3_c_406_n N_VGND_c_902_n 0.00178385f $X=10.755 $Y=1.177 $X2=0 $Y2=0
cc_383 N_A3_c_400_n N_VGND_c_903_n 0.00407103f $X=9.22 $Y=0.995 $X2=0 $Y2=0
cc_384 N_A3_c_401_n N_VGND_c_903_n 0.00407108f $X=9.69 $Y=0.995 $X2=0 $Y2=0
cc_385 N_A3_c_402_n N_VGND_c_903_n 0.00418642f $X=10.16 $Y=0.995 $X2=0 $Y2=0
cc_386 N_A3_c_403_n N_VGND_c_903_n 0.00572495f $X=10.68 $Y=0.995 $X2=0 $Y2=0
cc_387 A3 N_VGND_c_903_n 0.00147231f $X=10.765 $Y=0.765 $X2=0 $Y2=0
cc_388 N_A3_c_400_n N_A_1379_47#_c_1052_n 0.0144302f $X=9.22 $Y=0.995 $X2=0
+ $Y2=0
cc_389 N_A3_c_405_n N_A_1379_47#_c_1052_n 2.26856e-19 $X=10.68 $Y=1.202 $X2=0
+ $Y2=0
cc_390 N_A3_c_406_n N_A_1379_47#_c_1052_n 0.0106232f $X=10.755 $Y=1.177 $X2=0
+ $Y2=0
cc_391 N_A3_c_400_n N_A_1379_47#_c_1063_n 0.00391984f $X=9.22 $Y=0.995 $X2=0
+ $Y2=0
cc_392 N_A3_c_401_n N_A_1379_47#_c_1064_n 0.0126234f $X=9.69 $Y=0.995 $X2=0
+ $Y2=0
cc_393 N_A3_c_402_n N_A_1379_47#_c_1064_n 0.0123716f $X=10.16 $Y=0.995 $X2=0
+ $Y2=0
cc_394 N_A3_c_403_n N_A_1379_47#_c_1064_n 0.00421533f $X=10.68 $Y=0.995 $X2=0
+ $Y2=0
cc_395 N_A3_c_405_n N_A_1379_47#_c_1064_n 0.00753178f $X=10.68 $Y=1.202 $X2=0
+ $Y2=0
cc_396 N_A3_c_406_n N_A_1379_47#_c_1064_n 0.0413512f $X=10.755 $Y=1.177 $X2=0
+ $Y2=0
cc_397 N_A3_c_402_n N_A_1379_47#_c_1069_n 0.00393134f $X=10.16 $Y=0.995 $X2=0
+ $Y2=0
cc_398 N_A3_c_403_n N_A_1379_47#_c_1069_n 0.00381946f $X=10.68 $Y=0.995 $X2=0
+ $Y2=0
cc_399 N_A3_c_405_n N_A_1379_47#_c_1071_n 0.00312289f $X=10.68 $Y=1.202 $X2=0
+ $Y2=0
cc_400 N_A3_c_406_n N_A_1379_47#_c_1071_n 0.00914423f $X=10.755 $Y=1.177 $X2=0
+ $Y2=0
cc_401 N_A_27_297#_c_478_n N_Y_M1001_s 0.00367145f $X=3.935 $Y=2.34 $X2=0 $Y2=0
cc_402 N_A_27_297#_c_478_n N_Y_M1021_s 0.00367145f $X=3.935 $Y=2.34 $X2=0 $Y2=0
cc_403 N_A_27_297#_c_478_n N_Y_M1000_s 0.00367145f $X=3.935 $Y=2.34 $X2=0 $Y2=0
cc_404 N_A_27_297#_c_478_n N_Y_M1009_s 0.00367145f $X=3.935 $Y=2.34 $X2=0 $Y2=0
cc_405 N_A_27_297#_M1012_d N_Y_c_607_n 0.00504278f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_406 N_A_27_297#_c_478_n N_Y_c_607_n 0.0130979f $X=3.935 $Y=2.34 $X2=0 $Y2=0
cc_407 N_A_27_297#_M1035_d N_Y_c_611_n 0.00733799f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_408 N_A_27_297#_c_478_n N_Y_c_611_n 0.008366f $X=3.935 $Y=2.34 $X2=0 $Y2=0
cc_409 N_A_27_297#_M1004_d N_Y_c_637_n 0.00498385f $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_410 N_A_27_297#_c_478_n N_Y_c_637_n 0.0130979f $X=3.935 $Y=2.34 $X2=0 $Y2=0
cc_411 N_A_27_297#_c_478_n N_Y_c_613_n 0.0193386f $X=3.935 $Y=2.34 $X2=0 $Y2=0
cc_412 N_A_27_297#_c_478_n N_Y_c_619_n 0.0193386f $X=3.935 $Y=2.34 $X2=0 $Y2=0
cc_413 N_A_27_297#_c_478_n N_Y_c_642_n 0.0193386f $X=3.935 $Y=2.34 $X2=0 $Y2=0
cc_414 N_A_27_297#_c_489_n N_Y_c_642_n 0.0207808f $X=4.02 $Y=2.255 $X2=0 $Y2=0
cc_415 N_A_27_297#_c_490_n N_Y_c_642_n 0.0116213f $X=4.105 $Y=1.66 $X2=0 $Y2=0
cc_416 N_A_27_297#_M1035_d Y 0.00116564f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_417 N_A_27_297#_M1035_d Y 0.00430665f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_418 N_A_27_297#_c_478_n Y 0.0315499f $X=3.935 $Y=2.34 $X2=0 $Y2=0
cc_419 N_A_27_297#_c_493_n N_VPWR_M1005_s 0.00374243f $X=4.895 $Y=1.66 $X2=-0.19
+ $Y2=1.305
cc_420 N_A_27_297#_c_499_n N_VPWR_M1026_s 0.0169975f $X=6.29 $Y=1.66 $X2=0 $Y2=0
cc_421 N_A_27_297#_c_508_n N_VPWR_M1008_s 0.00370015f $X=7.465 $Y=1.66 $X2=0
+ $Y2=0
cc_422 N_A_27_297#_c_514_n N_VPWR_M1019_s 0.00370015f $X=8.405 $Y=1.66 $X2=0
+ $Y2=0
cc_423 N_A_27_297#_c_523_n N_VPWR_M1006_d 0.00377217f $X=9.865 $Y=1.66 $X2=0
+ $Y2=0
cc_424 N_A_27_297#_c_529_n N_VPWR_M1028_d 0.00377217f $X=10.805 $Y=1.66 $X2=0
+ $Y2=0
cc_425 N_A_27_297#_c_489_n N_VPWR_c_706_n 0.0362681f $X=4.02 $Y=2.255 $X2=0
+ $Y2=0
cc_426 N_A_27_297#_c_493_n N_VPWR_c_706_n 0.0209383f $X=4.895 $Y=1.66 $X2=0
+ $Y2=0
cc_427 N_A_27_297#_c_497_n N_VPWR_c_706_n 0.0336646f $X=4.98 $Y=1.96 $X2=0 $Y2=0
cc_428 N_A_27_297#_c_503_n N_VPWR_c_707_n 0.0210095f $X=6.375 $Y=1.96 $X2=0
+ $Y2=0
cc_429 N_A_27_297#_c_508_n N_VPWR_c_707_n 0.0209383f $X=7.465 $Y=1.66 $X2=0
+ $Y2=0
cc_430 N_A_27_297#_c_512_n N_VPWR_c_707_n 0.0336646f $X=7.55 $Y=1.96 $X2=0 $Y2=0
cc_431 N_A_27_297#_c_512_n N_VPWR_c_708_n 0.0410603f $X=7.55 $Y=1.96 $X2=0 $Y2=0
cc_432 N_A_27_297#_c_514_n N_VPWR_c_708_n 0.0210225f $X=8.405 $Y=1.66 $X2=0
+ $Y2=0
cc_433 N_A_27_297#_c_518_n N_VPWR_c_708_n 0.0336646f $X=8.49 $Y=1.96 $X2=0 $Y2=0
cc_434 N_A_27_297#_c_523_n N_VPWR_c_709_n 0.0209383f $X=9.865 $Y=1.66 $X2=0
+ $Y2=0
cc_435 N_A_27_297#_c_527_n N_VPWR_c_709_n 0.0336646f $X=9.95 $Y=1.96 $X2=0 $Y2=0
cc_436 N_A_27_297#_c_527_n N_VPWR_c_710_n 0.0410603f $X=9.95 $Y=1.96 $X2=0 $Y2=0
cc_437 N_A_27_297#_c_529_n N_VPWR_c_710_n 0.0209383f $X=10.805 $Y=1.66 $X2=0
+ $Y2=0
cc_438 N_A_27_297#_c_534_n N_VPWR_c_710_n 0.0336646f $X=10.89 $Y=1.96 $X2=0
+ $Y2=0
cc_439 N_A_27_297#_c_478_n N_VPWR_c_711_n 0.171502f $X=3.935 $Y=2.34 $X2=0 $Y2=0
cc_440 N_A_27_297#_c_489_n N_VPWR_c_711_n 0.00950266f $X=4.02 $Y=2.255 $X2=0
+ $Y2=0
cc_441 N_A_27_297#_c_497_n N_VPWR_c_712_n 0.0118139f $X=4.98 $Y=1.96 $X2=0 $Y2=0
cc_442 N_A_27_297#_c_503_n N_VPWR_c_713_n 0.0118139f $X=6.375 $Y=1.96 $X2=0
+ $Y2=0
cc_443 N_A_27_297#_c_512_n N_VPWR_c_714_n 0.0118139f $X=7.55 $Y=1.96 $X2=0 $Y2=0
cc_444 N_A_27_297#_c_518_n N_VPWR_c_715_n 0.0118139f $X=8.49 $Y=1.96 $X2=0 $Y2=0
cc_445 N_A_27_297#_c_527_n N_VPWR_c_716_n 0.0118139f $X=9.95 $Y=1.96 $X2=0 $Y2=0
cc_446 N_A_27_297#_c_534_n N_VPWR_c_717_n 0.0118139f $X=10.89 $Y=1.96 $X2=0
+ $Y2=0
cc_447 N_A_27_297#_M1001_d N_VPWR_c_705_n 0.0021994f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_448 N_A_27_297#_M1012_d N_VPWR_c_705_n 0.00233855f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_449 N_A_27_297#_M1035_d N_VPWR_c_705_n 0.00233855f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_450 N_A_27_297#_M1004_d N_VPWR_c_705_n 0.00233855f $X=2.935 $Y=1.485 $X2=0
+ $Y2=0
cc_451 N_A_27_297#_M1016_d N_VPWR_c_705_n 0.00528666f $X=3.875 $Y=1.485 $X2=0
+ $Y2=0
cc_452 N_A_27_297#_M1011_d N_VPWR_c_705_n 0.00647849f $X=4.835 $Y=1.485 $X2=0
+ $Y2=0
cc_453 N_A_27_297#_M1029_d N_VPWR_c_705_n 0.0165942f $X=6.23 $Y=1.485 $X2=0
+ $Y2=0
cc_454 N_A_27_297#_M1014_d N_VPWR_c_705_n 0.00647849f $X=7.405 $Y=1.485 $X2=0
+ $Y2=0
cc_455 N_A_27_297#_M1027_d N_VPWR_c_705_n 0.0288246f $X=8.345 $Y=1.485 $X2=0
+ $Y2=0
cc_456 N_A_27_297#_M1023_s N_VPWR_c_705_n 0.00647849f $X=9.805 $Y=1.485 $X2=0
+ $Y2=0
cc_457 N_A_27_297#_M1032_s N_VPWR_c_705_n 0.00568146f $X=10.745 $Y=1.485 $X2=0
+ $Y2=0
cc_458 N_A_27_297#_c_478_n N_VPWR_c_705_n 0.132351f $X=3.935 $Y=2.34 $X2=0 $Y2=0
cc_459 N_A_27_297#_c_489_n N_VPWR_c_705_n 0.00641762f $X=4.02 $Y=2.255 $X2=0
+ $Y2=0
cc_460 N_A_27_297#_c_497_n N_VPWR_c_705_n 0.00646998f $X=4.98 $Y=1.96 $X2=0
+ $Y2=0
cc_461 N_A_27_297#_c_503_n N_VPWR_c_705_n 0.00646998f $X=6.375 $Y=1.96 $X2=0
+ $Y2=0
cc_462 N_A_27_297#_c_512_n N_VPWR_c_705_n 0.00646998f $X=7.55 $Y=1.96 $X2=0
+ $Y2=0
cc_463 N_A_27_297#_c_518_n N_VPWR_c_705_n 0.00646998f $X=8.49 $Y=1.96 $X2=0
+ $Y2=0
cc_464 N_A_27_297#_c_527_n N_VPWR_c_705_n 0.00646998f $X=9.95 $Y=1.96 $X2=0
+ $Y2=0
cc_465 N_A_27_297#_c_534_n N_VPWR_c_705_n 0.00646998f $X=10.89 $Y=1.96 $X2=0
+ $Y2=0
cc_466 N_A_27_297#_c_499_n N_VPWR_c_720_n 0.0513372f $X=6.29 $Y=1.66 $X2=0 $Y2=0
cc_467 N_Y_M1001_s N_VPWR_c_705_n 0.00235479f $X=0.585 $Y=1.485 $X2=0 $Y2=0
cc_468 N_Y_M1021_s N_VPWR_c_705_n 0.00235479f $X=1.525 $Y=1.485 $X2=0 $Y2=0
cc_469 N_Y_M1000_s N_VPWR_c_705_n 0.00235479f $X=2.465 $Y=1.485 $X2=0 $Y2=0
cc_470 N_Y_M1009_s N_VPWR_c_705_n 0.00235479f $X=3.405 $Y=1.485 $X2=0 $Y2=0
cc_471 N_Y_c_603_n N_A_27_47#_M1017_d 0.00407984f $X=6 $Y=0.72 $X2=0 $Y2=0
cc_472 N_Y_c_603_n N_A_27_47#_M1033_d 0.0102196f $X=6 $Y=0.72 $X2=0 $Y2=0
cc_473 Y N_A_27_47#_c_847_n 0.00386389f $X=2.41 $Y=1.105 $X2=0 $Y2=0
cc_474 N_Y_M1010_s N_A_27_47#_c_836_n 0.00413629f $X=2.425 $Y=0.235 $X2=0 $Y2=0
cc_475 N_Y_M1030_s N_A_27_47#_c_836_n 0.00523126f $X=3.365 $Y=0.235 $X2=0 $Y2=0
cc_476 N_Y_c_631_n N_A_27_47#_c_836_n 0.0123377f $X=2.505 $Y=0.805 $X2=0 $Y2=0
cc_477 N_Y_c_603_n N_A_27_47#_c_836_n 0.0824481f $X=6 $Y=0.72 $X2=0 $Y2=0
cc_478 Y N_A_27_47#_c_836_n 0.00467444f $X=2.41 $Y=1.105 $X2=0 $Y2=0
cc_479 N_Y_c_603_n N_VGND_c_895_n 0.00438623f $X=6 $Y=0.72 $X2=0 $Y2=0
cc_480 N_Y_M1010_s N_VGND_c_903_n 0.00259839f $X=2.425 $Y=0.235 $X2=0 $Y2=0
cc_481 N_Y_M1030_s N_VGND_c_903_n 0.00300439f $X=3.365 $Y=0.235 $X2=0 $Y2=0
cc_482 N_Y_M1007_s N_VGND_c_903_n 0.00259839f $X=4.925 $Y=0.235 $X2=0 $Y2=0
cc_483 N_Y_M1031_s N_VGND_c_903_n 0.00259839f $X=5.865 $Y=0.235 $X2=0 $Y2=0
cc_484 N_Y_c_603_n N_VGND_c_903_n 0.0128891f $X=6 $Y=0.72 $X2=0 $Y2=0
cc_485 N_Y_c_603_n N_A_893_47#_M1007_d 0.0063705f $X=6 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_486 N_Y_c_603_n N_A_893_47#_M1013_d 0.00439968f $X=6 $Y=0.72 $X2=0 $Y2=0
cc_487 N_Y_M1007_s N_A_893_47#_c_1023_n 0.00414886f $X=4.925 $Y=0.235 $X2=0
+ $Y2=0
cc_488 N_Y_M1031_s N_A_893_47#_c_1023_n 0.00415474f $X=5.865 $Y=0.235 $X2=0
+ $Y2=0
cc_489 N_Y_c_603_n N_A_893_47#_c_1023_n 0.0916483f $X=6 $Y=0.72 $X2=0 $Y2=0
cc_490 N_A_27_47#_c_838_n N_VGND_M1002_s 0.00439476f $X=1.115 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_491 N_A_27_47#_c_847_n N_VGND_M1025_s 0.00439476f $X=2.055 $Y=0.72 $X2=0
+ $Y2=0
cc_492 N_A_27_47#_c_837_n N_VGND_c_893_n 0.0116326f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_493 N_A_27_47#_c_838_n N_VGND_c_893_n 0.00244812f $X=1.115 $Y=0.72 $X2=0
+ $Y2=0
cc_494 N_A_27_47#_c_838_n N_VGND_c_894_n 0.00313948f $X=1.115 $Y=0.72 $X2=0
+ $Y2=0
cc_495 N_A_27_47#_c_846_n N_VGND_c_894_n 0.01143f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_496 N_A_27_47#_c_847_n N_VGND_c_894_n 0.00244812f $X=2.055 $Y=0.72 $X2=0
+ $Y2=0
cc_497 N_A_27_47#_c_847_n N_VGND_c_895_n 0.0031329f $X=2.055 $Y=0.72 $X2=0 $Y2=0
cc_498 N_A_27_47#_c_874_p N_VGND_c_895_n 0.00894629f $X=2.14 $Y=0.465 $X2=0
+ $Y2=0
cc_499 N_A_27_47#_c_836_n N_VGND_c_895_n 0.0881863f $X=4.02 $Y=0.38 $X2=0 $Y2=0
cc_500 N_A_27_47#_c_837_n N_VGND_c_898_n 0.0156777f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_501 N_A_27_47#_c_838_n N_VGND_c_898_n 0.0213178f $X=1.115 $Y=0.72 $X2=0 $Y2=0
cc_502 N_A_27_47#_c_846_n N_VGND_c_899_n 0.0156777f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_503 N_A_27_47#_c_847_n N_VGND_c_899_n 0.0213178f $X=2.055 $Y=0.72 $X2=0 $Y2=0
cc_504 N_A_27_47#_M1002_d N_VGND_c_903_n 0.00430496f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_505 N_A_27_47#_M1024_d N_VGND_c_903_n 0.00309604f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_506 N_A_27_47#_M1039_d N_VGND_c_903_n 0.00236972f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_507 N_A_27_47#_M1017_d N_VGND_c_903_n 0.00258215f $X=2.895 $Y=0.235 $X2=0
+ $Y2=0
cc_508 N_A_27_47#_M1033_d N_VGND_c_903_n 0.00211652f $X=3.885 $Y=0.235 $X2=0
+ $Y2=0
cc_509 N_A_27_47#_c_837_n N_VGND_c_903_n 0.00643448f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_510 N_A_27_47#_c_838_n N_VGND_c_903_n 0.0114934f $X=1.115 $Y=0.72 $X2=0 $Y2=0
cc_511 N_A_27_47#_c_846_n N_VGND_c_903_n 0.00643448f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_512 N_A_27_47#_c_847_n N_VGND_c_903_n 0.0115249f $X=2.055 $Y=0.72 $X2=0 $Y2=0
cc_513 N_A_27_47#_c_874_p N_VGND_c_903_n 0.00636368f $X=2.14 $Y=0.465 $X2=0
+ $Y2=0
cc_514 N_A_27_47#_c_836_n N_VGND_c_903_n 0.068219f $X=4.02 $Y=0.38 $X2=0 $Y2=0
cc_515 N_A_27_47#_c_836_n N_A_893_47#_c_1023_n 0.0123435f $X=4.02 $Y=0.38 $X2=0
+ $Y2=0
cc_516 N_VGND_c_903_n N_A_893_47#_M1007_d 0.00253093f $X=10.81 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_517 N_VGND_c_903_n N_A_893_47#_M1013_d 0.00258215f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_518 N_VGND_c_903_n N_A_893_47#_M1034_d 0.00332948f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_519 N_VGND_c_903_n N_A_893_47#_M1018_d 0.00258215f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_520 N_VGND_c_903_n N_A_893_47#_M1036_d 0.00211652f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_521 N_VGND_c_892_n N_A_893_47#_c_1023_n 0.0137364f $X=9.01 $Y=0.38 $X2=0
+ $Y2=0
cc_522 N_VGND_c_895_n N_A_893_47#_c_1023_n 0.19176f $X=8.845 $Y=0 $X2=0 $Y2=0
cc_523 N_VGND_c_903_n N_A_893_47#_c_1023_n 0.147661f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_524 N_VGND_c_903_n N_A_1379_47#_M1003_s 0.00259839f $X=10.81 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_525 N_VGND_c_903_n N_A_1379_47#_M1020_s 0.00300439f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_526 N_VGND_c_903_n N_A_1379_47#_M1015_d 0.00307738f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_527 N_VGND_c_903_n N_A_1379_47#_M1037_d 0.00680846f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_528 N_VGND_M1015_s N_A_1379_47#_c_1052_n 0.0105655f $X=8.885 $Y=0.235 $X2=0
+ $Y2=0
cc_529 N_VGND_c_892_n N_A_1379_47#_c_1052_n 0.0206068f $X=9.01 $Y=0.38 $X2=0
+ $Y2=0
cc_530 N_VGND_c_895_n N_A_1379_47#_c_1052_n 0.00346265f $X=8.845 $Y=0 $X2=0
+ $Y2=0
cc_531 N_VGND_c_896_n N_A_1379_47#_c_1052_n 0.00325651f $X=9.735 $Y=0 $X2=0
+ $Y2=0
cc_532 N_VGND_c_903_n N_A_1379_47#_c_1052_n 0.0157842f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_533 N_VGND_c_892_n N_A_1379_47#_c_1063_n 0.012714f $X=9.01 $Y=0.38 $X2=0
+ $Y2=0
cc_534 N_VGND_c_896_n N_A_1379_47#_c_1063_n 0.01143f $X=9.735 $Y=0 $X2=0 $Y2=0
cc_535 N_VGND_c_903_n N_A_1379_47#_c_1063_n 0.00643448f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_536 N_VGND_M1022_s N_A_1379_47#_c_1064_n 0.00439476f $X=9.765 $Y=0.235 $X2=0
+ $Y2=0
cc_537 N_VGND_c_896_n N_A_1379_47#_c_1064_n 0.00245287f $X=9.735 $Y=0 $X2=0
+ $Y2=0
cc_538 N_VGND_c_897_n N_A_1379_47#_c_1064_n 0.0032663f $X=10.685 $Y=0 $X2=0
+ $Y2=0
cc_539 N_VGND_c_901_n N_A_1379_47#_c_1064_n 0.0197774f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_540 N_VGND_c_903_n N_A_1379_47#_c_1064_n 0.011481f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_541 N_VGND_c_897_n N_A_1379_47#_c_1069_n 0.0116326f $X=10.685 $Y=0 $X2=0
+ $Y2=0
cc_542 N_VGND_c_901_n N_A_1379_47#_c_1069_n 0.0128539f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_543 N_VGND_c_902_n N_A_1379_47#_c_1069_n 0.0150302f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_544 N_VGND_c_903_n N_A_1379_47#_c_1069_n 0.00643448f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_545 N_A_893_47#_c_1023_n N_A_1379_47#_M1003_s 0.00414886f $X=8.49 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_546 N_A_893_47#_c_1023_n N_A_1379_47#_M1020_s 0.00523924f $X=8.49 $Y=0.38
+ $X2=0 $Y2=0
cc_547 N_A_893_47#_M1018_d N_A_1379_47#_c_1052_n 0.00439968f $X=7.365 $Y=0.235
+ $X2=0 $Y2=0
cc_548 N_A_893_47#_M1036_d N_A_1379_47#_c_1052_n 0.00724259f $X=8.355 $Y=0.235
+ $X2=0 $Y2=0
cc_549 N_A_893_47#_c_1023_n N_A_1379_47#_c_1052_n 0.0935475f $X=8.49 $Y=0.38
+ $X2=0 $Y2=0
