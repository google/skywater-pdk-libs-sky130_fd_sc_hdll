* File: sky130_fd_sc_hdll__a22o_2.pxi.spice
* Created: Wed Sep  2 08:18:37 2020
* 
x_PM_SKY130_FD_SC_HDLL__A22O_2%B2 N_B2_c_58_n N_B2_M1005_g N_B2_c_59_n
+ N_B2_M1009_g B2 N_B2_c_60_n PM_SKY130_FD_SC_HDLL__A22O_2%B2
x_PM_SKY130_FD_SC_HDLL__A22O_2%B1 N_B1_c_82_n N_B1_M1010_g N_B1_c_83_n
+ N_B1_M1000_g B1 B1 N_B1_c_85_n B1 PM_SKY130_FD_SC_HDLL__A22O_2%B1
x_PM_SKY130_FD_SC_HDLL__A22O_2%A1 N_A1_c_118_n N_A1_M1008_g N_A1_c_119_n
+ N_A1_M1006_g A1 A1 N_A1_c_121_n PM_SKY130_FD_SC_HDLL__A22O_2%A1
x_PM_SKY130_FD_SC_HDLL__A22O_2%A2 N_A2_c_154_n N_A2_M1003_g N_A2_c_155_n
+ N_A2_M1007_g A2 PM_SKY130_FD_SC_HDLL__A22O_2%A2
x_PM_SKY130_FD_SC_HDLL__A22O_2%A_27_297# N_A_27_297#_M1010_d N_A_27_297#_M1006_s
+ N_A_27_297#_M1005_s N_A_27_297#_M1000_d N_A_27_297#_c_194_n
+ N_A_27_297#_M1001_g N_A_27_297#_c_187_n N_A_27_297#_M1002_g
+ N_A_27_297#_c_195_n N_A_27_297#_M1011_g N_A_27_297#_c_188_n
+ N_A_27_297#_M1004_g N_A_27_297#_c_196_n N_A_27_297#_c_197_n
+ N_A_27_297#_c_198_n N_A_27_297#_c_199_n N_A_27_297#_c_189_n
+ N_A_27_297#_c_228_n N_A_27_297#_c_190_n N_A_27_297#_c_191_n
+ N_A_27_297#_c_192_n N_A_27_297#_c_201_n N_A_27_297#_c_210_n
+ N_A_27_297#_c_193_n PM_SKY130_FD_SC_HDLL__A22O_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A22O_2%A_117_297# N_A_117_297#_M1005_d
+ N_A_117_297#_M1008_d N_A_117_297#_c_312_n N_A_117_297#_c_321_n
+ N_A_117_297#_c_327_p N_A_117_297#_c_322_n
+ PM_SKY130_FD_SC_HDLL__A22O_2%A_117_297#
x_PM_SKY130_FD_SC_HDLL__A22O_2%VPWR N_VPWR_M1008_s N_VPWR_M1003_d N_VPWR_M1011_s
+ N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n
+ N_VPWR_c_341_n VPWR N_VPWR_c_342_n N_VPWR_c_343_n N_VPWR_c_344_n
+ N_VPWR_c_335_n PM_SKY130_FD_SC_HDLL__A22O_2%VPWR
x_PM_SKY130_FD_SC_HDLL__A22O_2%X N_X_M1002_s N_X_M1001_d X X X X X X N_X_c_405_n
+ X PM_SKY130_FD_SC_HDLL__A22O_2%X
x_PM_SKY130_FD_SC_HDLL__A22O_2%VGND N_VGND_M1009_s N_VGND_M1007_d N_VGND_M1004_d
+ N_VGND_c_416_n N_VGND_c_417_n N_VGND_c_418_n N_VGND_c_419_n N_VGND_c_420_n
+ VGND N_VGND_c_421_n N_VGND_c_422_n N_VGND_c_423_n N_VGND_c_424_n
+ PM_SKY130_FD_SC_HDLL__A22O_2%VGND
cc_1 VNB N_B2_c_58_n 0.030174f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_B2_c_59_n 0.0202522f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_3 VNB N_B2_c_60_n 0.0143633f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_4 VNB N_B1_c_82_n 0.0190413f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_B1_c_83_n 0.0272683f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB B1 0.00528653f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_B1_c_85_n 0.00534702f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A1_c_118_n 0.0328269f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_9 VNB N_A1_c_119_n 0.0203751f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_10 VNB A1 0.00494419f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_11 VNB N_A1_c_121_n 0.00250827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A2_c_154_n 0.0223122f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_13 VNB N_A2_c_155_n 0.01741f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_14 VNB A2 0.00512384f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_15 VNB N_A_27_297#_c_187_n 0.0168637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_297#_c_188_n 0.0195177f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_297#_c_189_n 0.0129014f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_297#_c_190_n 0.00388218f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_297#_c_191_n 0.00182992f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_297#_c_192_n 9.16142e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_297#_c_193_n 0.0560156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_335_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB X 7.1422e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_24 VNB N_VGND_c_416_n 0.0128958f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_25 VNB N_VGND_c_417_n 0.0283775f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.175
cc_26 VNB N_VGND_c_418_n 0.0028208f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_419_n 0.0123291f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_420_n 0.0118305f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_421_n 0.0442162f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_422_n 0.023147f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_423_n 0.00574292f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_424_n 0.224509f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VPB N_B2_c_58_n 0.0333642f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_34 VPB N_B1_c_83_n 0.0334904f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_35 VPB N_A1_c_118_n 0.0349922f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_36 VPB N_A2_c_154_n 0.0270079f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_37 VPB N_A_27_297#_c_194_n 0.0160769f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_27_297#_c_195_n 0.0197262f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_297#_c_196_n 0.00746643f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_297#_c_197_n 0.025859f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_297#_c_198_n 0.0303613f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_297#_c_199_n 0.00978665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_297#_c_192_n 0.00133183f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_27_297#_c_201_n 0.00257199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_297#_c_193_n 0.0282458f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_117_297#_c_312_n 0.00819467f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_47 VPB N_VPWR_c_336_n 0.00606222f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.175
cc_48 VPB N_VPWR_c_337_n 0.00285945f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_338_n 0.0123032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_339_n 0.00901916f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_340_n 0.01762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_341_n 0.00513801f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_342_n 0.0386236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_343_n 0.0211125f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_344_n 0.00546578f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_335_n 0.0496942f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB X 0.00104381f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_58 N_B2_c_59_n N_B1_c_82_n 0.0339429f $X=0.52 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_59 N_B2_c_58_n N_B1_c_83_n 0.0754187f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_60 N_B2_c_60_n N_B1_c_83_n 7.27588e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_61 N_B2_c_58_n B1 3.46207e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_62 N_B2_c_58_n N_B1_c_85_n 9.36086e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_63 N_B2_c_60_n N_B1_c_85_n 0.0165024f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_64 N_B2_c_58_n N_A_27_297#_c_196_n 4.66918e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_65 N_B2_c_58_n N_A_27_297#_c_197_n 0.010181f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_66 N_B2_c_58_n N_A_27_297#_c_198_n 0.0116083f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_67 N_B2_c_60_n N_A_27_297#_c_198_n 0.013348f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_68 N_B2_c_58_n N_A_27_297#_c_199_n 0.00443521f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_69 N_B2_c_60_n N_A_27_297#_c_199_n 0.0263882f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_70 N_B2_c_59_n N_A_27_297#_c_189_n 7.24737e-19 $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_71 N_B2_c_58_n N_A_27_297#_c_210_n 0.0104293f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_72 N_B2_c_58_n N_VPWR_c_342_n 0.00429425f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_73 N_B2_c_58_n N_VPWR_c_335_n 0.00700259f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_74 N_B2_c_58_n N_VGND_c_417_n 0.00417825f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_75 N_B2_c_59_n N_VGND_c_417_n 0.0265784f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_76 N_B2_c_60_n N_VGND_c_417_n 0.0302791f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_77 N_B2_c_59_n N_VGND_c_424_n 7.20442e-19 $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_78 N_B1_c_83_n N_A1_c_118_n 0.00760856f $X=0.965 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_79 B1 N_A1_c_118_n 2.45417e-19 $X=1.085 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_80 N_B1_c_85_n N_A1_c_118_n 6.95005e-19 $X=1.202 $Y=1.075 $X2=-0.19 $Y2=-0.24
cc_81 N_B1_c_83_n A1 2.12489e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_82 B1 A1 0.0306521f $X=1.085 $Y=0.765 $X2=0 $Y2=0
cc_83 N_B1_c_83_n N_A1_c_121_n 5.87023e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_84 N_B1_c_85_n N_A1_c_121_n 0.0172678f $X=1.202 $Y=1.075 $X2=0 $Y2=0
cc_85 B1 N_A_27_297#_M1010_d 0.00660077f $X=1.085 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_86 N_B1_c_83_n N_A_27_297#_c_197_n 0.00138485f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_87 N_B1_c_83_n N_A_27_297#_c_198_n 0.0178995f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_88 N_B1_c_85_n N_A_27_297#_c_198_n 0.0381822f $X=1.202 $Y=1.075 $X2=0 $Y2=0
cc_89 N_B1_c_82_n N_A_27_297#_c_189_n 0.00810253f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_90 N_B1_c_83_n N_A_27_297#_c_189_n 0.00204237f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_91 B1 N_A_27_297#_c_189_n 0.0210337f $X=1.085 $Y=0.765 $X2=0 $Y2=0
cc_92 N_B1_c_85_n N_A_27_297#_c_189_n 0.00447978f $X=1.202 $Y=1.075 $X2=0 $Y2=0
cc_93 N_B1_c_83_n N_A_27_297#_c_201_n 0.00151714f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_94 N_B1_c_83_n N_A_27_297#_c_210_n 0.00864172f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_95 N_B1_c_83_n N_A_117_297#_c_312_n 0.0153152f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_96 N_B1_c_83_n N_VPWR_c_336_n 0.00236094f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_97 N_B1_c_83_n N_VPWR_c_342_n 0.00429453f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_98 N_B1_c_83_n N_VPWR_c_335_n 0.00737353f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_99 N_B1_c_82_n N_VGND_c_417_n 0.00413342f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_100 B1 N_VGND_c_417_n 0.00627099f $X=1.085 $Y=0.765 $X2=0 $Y2=0
cc_101 N_B1_c_82_n N_VGND_c_421_n 0.0042613f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_102 N_B1_c_82_n N_VGND_c_424_n 0.0081372f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A1_c_118_n N_A2_c_154_n 0.0442241f $X=1.955 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_104 A1 N_A2_c_154_n 3.46144e-19 $X=1.565 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_105 N_A1_c_121_n N_A2_c_154_n 2.33401e-19 $X=1.775 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_106 N_A1_c_119_n N_A2_c_155_n 0.0245323f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_107 N_A1_c_118_n A2 0.0015187f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A1_c_121_n A2 0.0135294f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_109 A1 N_A_27_297#_M1006_s 0.0062896f $X=1.565 $Y=0.765 $X2=0 $Y2=0
cc_110 N_A1_c_118_n N_A_27_297#_c_198_n 0.0232209f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A1_c_121_n N_A_27_297#_c_198_n 0.032215f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A1_c_118_n N_A_27_297#_c_189_n 0.00213831f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A1_c_119_n N_A_27_297#_c_189_n 0.0138667f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_114 A1 N_A_27_297#_c_189_n 0.0233314f $X=1.565 $Y=0.765 $X2=0 $Y2=0
cc_115 N_A1_c_121_n N_A_27_297#_c_189_n 0.00241976f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A1_c_119_n N_A_27_297#_c_228_n 0.0047574f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_117 A1 N_A_27_297#_c_228_n 0.002932f $X=1.565 $Y=0.765 $X2=0 $Y2=0
cc_118 N_A1_c_119_n N_A_27_297#_c_191_n 0.00197969f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_119 A1 N_A_27_297#_c_191_n 0.00939017f $X=1.565 $Y=0.765 $X2=0 $Y2=0
cc_120 N_A1_c_118_n N_A_117_297#_c_312_n 0.0161386f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A1_c_118_n N_VPWR_c_336_n 0.0109451f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A1_c_118_n N_VPWR_c_340_n 0.00388325f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A1_c_118_n N_VPWR_c_335_n 0.00469535f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A1_c_119_n N_VGND_c_418_n 0.00132905f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A1_c_119_n N_VGND_c_421_n 0.00357877f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A1_c_119_n N_VGND_c_424_n 0.00683557f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A2_c_154_n N_A_27_297#_c_194_n 0.0182273f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A2_c_155_n N_A_27_297#_c_187_n 0.0213207f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A2_c_154_n N_A_27_297#_c_198_n 0.0213791f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_130 A2 N_A_27_297#_c_198_n 0.0313942f $X=2.42 $Y=1.105 $X2=0 $Y2=0
cc_131 N_A2_c_155_n N_A_27_297#_c_189_n 0.00214141f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A2_c_155_n N_A_27_297#_c_228_n 0.00425788f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A2_c_154_n N_A_27_297#_c_190_n 0.00363179f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A2_c_155_n N_A_27_297#_c_190_n 0.0118333f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_135 A2 N_A_27_297#_c_190_n 0.0226779f $X=2.42 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A2_c_154_n N_A_27_297#_c_191_n 7.67796e-19 $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_137 A2 N_A_27_297#_c_191_n 0.0113712f $X=2.42 $Y=1.105 $X2=0 $Y2=0
cc_138 N_A2_c_154_n N_A_27_297#_c_192_n 0.00351724f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A2_c_155_n N_A_27_297#_c_192_n 0.00171795f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_140 A2 N_A_27_297#_c_192_n 0.0123149f $X=2.42 $Y=1.105 $X2=0 $Y2=0
cc_141 N_A2_c_154_n N_A_27_297#_c_193_n 0.0258002f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_142 A2 N_A_27_297#_c_193_n 0.00141899f $X=2.42 $Y=1.105 $X2=0 $Y2=0
cc_143 N_A2_c_154_n N_VPWR_c_336_n 0.00103987f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A2_c_154_n N_VPWR_c_337_n 0.00313517f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A2_c_154_n N_VPWR_c_340_n 0.00702461f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A2_c_154_n N_VPWR_c_335_n 0.0127114f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A2_c_155_n N_VGND_c_418_n 0.0125614f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A2_c_155_n N_VGND_c_421_n 0.0020416f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A2_c_155_n N_VGND_c_424_n 0.00303429f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A_27_297#_c_198_n N_A_117_297#_M1005_d 0.00184351f $X=2.845 $Y=1.54
+ $X2=-0.19 $Y2=-0.24
cc_151 N_A_27_297#_c_210_n N_A_117_297#_M1005_d 0.00349652f $X=1.035 $Y=2.36
+ $X2=-0.19 $Y2=-0.24
cc_152 N_A_27_297#_c_198_n N_A_117_297#_M1008_d 0.00250945f $X=2.845 $Y=1.54
+ $X2=0 $Y2=0
cc_153 N_A_27_297#_M1000_d N_A_117_297#_c_312_n 0.00589053f $X=1.055 $Y=1.485
+ $X2=0 $Y2=0
cc_154 N_A_27_297#_c_201_n N_A_117_297#_c_312_n 0.0157862f $X=1.2 $Y=2.34 $X2=0
+ $Y2=0
cc_155 N_A_27_297#_c_210_n N_A_117_297#_c_312_n 0.00707535f $X=1.035 $Y=2.36
+ $X2=0 $Y2=0
cc_156 N_A_27_297#_c_198_n N_A_117_297#_c_321_n 0.0169022f $X=2.845 $Y=1.54
+ $X2=0 $Y2=0
cc_157 N_A_27_297#_c_197_n N_A_117_297#_c_322_n 0.0217133f $X=0.26 $Y=1.66 $X2=0
+ $Y2=0
cc_158 N_A_27_297#_c_198_n N_A_117_297#_c_322_n 0.0929038f $X=2.845 $Y=1.54
+ $X2=0 $Y2=0
cc_159 N_A_27_297#_c_210_n N_A_117_297#_c_322_n 0.0124153f $X=1.035 $Y=2.36
+ $X2=0 $Y2=0
cc_160 N_A_27_297#_c_198_n N_VPWR_M1008_s 0.00296218f $X=2.845 $Y=1.54 $X2=-0.19
+ $Y2=-0.24
cc_161 N_A_27_297#_c_198_n N_VPWR_M1003_d 0.00278342f $X=2.845 $Y=1.54 $X2=0
+ $Y2=0
cc_162 N_A_27_297#_c_201_n N_VPWR_c_336_n 0.0169231f $X=1.2 $Y=2.34 $X2=0 $Y2=0
cc_163 N_A_27_297#_c_194_n N_VPWR_c_337_n 0.0122777f $X=3 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_27_297#_c_195_n N_VPWR_c_337_n 9.95344e-19 $X=3.47 $Y=1.41 $X2=0
+ $Y2=0
cc_165 N_A_27_297#_c_198_n N_VPWR_c_337_n 0.0146838f $X=2.845 $Y=1.54 $X2=0
+ $Y2=0
cc_166 N_A_27_297#_c_193_n N_VPWR_c_337_n 2.53351e-19 $X=3.47 $Y=1.202 $X2=0
+ $Y2=0
cc_167 N_A_27_297#_c_195_n N_VPWR_c_339_n 0.0239562f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A_27_297#_c_196_n N_VPWR_c_342_n 0.0211994f $X=0.26 $Y=2.295 $X2=0
+ $Y2=0
cc_169 N_A_27_297#_c_210_n N_VPWR_c_342_n 0.0543516f $X=1.035 $Y=2.36 $X2=0
+ $Y2=0
cc_170 N_A_27_297#_c_194_n N_VPWR_c_343_n 0.00622633f $X=3 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_27_297#_c_195_n N_VPWR_c_343_n 0.00430719f $X=3.47 $Y=1.41 $X2=0
+ $Y2=0
cc_172 N_A_27_297#_M1005_s N_VPWR_c_335_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_173 N_A_27_297#_M1000_d N_VPWR_c_335_n 0.00217543f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_174 N_A_27_297#_c_194_n N_VPWR_c_335_n 0.0104011f $X=3 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_27_297#_c_195_n N_VPWR_c_335_n 0.00713389f $X=3.47 $Y=1.41 $X2=0
+ $Y2=0
cc_176 N_A_27_297#_c_196_n N_VPWR_c_335_n 0.012545f $X=0.26 $Y=2.295 $X2=0 $Y2=0
cc_177 N_A_27_297#_c_210_n N_VPWR_c_335_n 0.0334433f $X=1.035 $Y=2.36 $X2=0
+ $Y2=0
cc_178 N_A_27_297#_c_194_n X 0.00531251f $X=3 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_27_297#_c_187_n X 0.00550066f $X=3.025 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_27_297#_c_195_n X 0.0120688f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_27_297#_c_188_n X 0.011401f $X=3.495 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_27_297#_c_198_n X 0.011299f $X=2.845 $Y=1.54 $X2=0 $Y2=0
cc_183 N_A_27_297#_c_190_n X 0.0112831f $X=2.845 $Y=0.82 $X2=0 $Y2=0
cc_184 N_A_27_297#_c_192_n X 0.0321275f $X=2.93 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_27_297#_c_193_n X 0.039785f $X=3.47 $Y=1.202 $X2=0 $Y2=0
cc_186 N_A_27_297#_c_195_n X 0.00454654f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_187 N_A_27_297#_c_193_n X 0.00300738f $X=3.47 $Y=1.202 $X2=0 $Y2=0
cc_188 N_A_27_297#_c_195_n X 0.0120374f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A_27_297#_c_188_n N_X_c_405_n 0.00736996f $X=3.495 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_27_297#_c_193_n N_X_c_405_n 0.00157084f $X=3.47 $Y=1.202 $X2=0 $Y2=0
cc_191 N_A_27_297#_c_190_n N_VGND_M1007_d 0.00270407f $X=2.845 $Y=0.82 $X2=0
+ $Y2=0
cc_192 N_A_27_297#_c_189_n N_VGND_c_417_n 0.0138716f $X=2.125 $Y=0.38 $X2=0
+ $Y2=0
cc_193 N_A_27_297#_c_187_n N_VGND_c_418_n 0.00659659f $X=3.025 $Y=0.995 $X2=0
+ $Y2=0
cc_194 N_A_27_297#_c_189_n N_VGND_c_418_n 0.0177122f $X=2.125 $Y=0.38 $X2=0
+ $Y2=0
cc_195 N_A_27_297#_c_228_n N_VGND_c_418_n 0.00377501f $X=2.21 $Y=0.735 $X2=0
+ $Y2=0
cc_196 N_A_27_297#_c_190_n N_VGND_c_418_n 0.0250392f $X=2.845 $Y=0.82 $X2=0
+ $Y2=0
cc_197 N_A_27_297#_c_193_n N_VGND_c_418_n 2.76193e-19 $X=3.47 $Y=1.202 $X2=0
+ $Y2=0
cc_198 N_A_27_297#_c_188_n N_VGND_c_420_n 0.017969f $X=3.495 $Y=0.995 $X2=0
+ $Y2=0
cc_199 N_A_27_297#_c_189_n N_VGND_c_421_n 0.0882414f $X=2.125 $Y=0.38 $X2=0
+ $Y2=0
cc_200 N_A_27_297#_c_190_n N_VGND_c_421_n 0.00251212f $X=2.845 $Y=0.82 $X2=0
+ $Y2=0
cc_201 N_A_27_297#_c_187_n N_VGND_c_422_n 0.00521982f $X=3.025 $Y=0.995 $X2=0
+ $Y2=0
cc_202 N_A_27_297#_c_188_n N_VGND_c_422_n 0.00374367f $X=3.495 $Y=0.995 $X2=0
+ $Y2=0
cc_203 N_A_27_297#_c_190_n N_VGND_c_422_n 0.00148976f $X=2.845 $Y=0.82 $X2=0
+ $Y2=0
cc_204 N_A_27_297#_M1010_d N_VGND_c_424_n 0.00250339f $X=0.975 $Y=0.235 $X2=0
+ $Y2=0
cc_205 N_A_27_297#_M1006_s N_VGND_c_424_n 0.00250339f $X=1.595 $Y=0.235 $X2=0
+ $Y2=0
cc_206 N_A_27_297#_c_187_n N_VGND_c_424_n 0.00899703f $X=3.025 $Y=0.995 $X2=0
+ $Y2=0
cc_207 N_A_27_297#_c_188_n N_VGND_c_424_n 0.00688545f $X=3.495 $Y=0.995 $X2=0
+ $Y2=0
cc_208 N_A_27_297#_c_189_n N_VGND_c_424_n 0.052369f $X=2.125 $Y=0.38 $X2=0 $Y2=0
cc_209 N_A_27_297#_c_190_n N_VGND_c_424_n 0.00993099f $X=2.845 $Y=0.82 $X2=0
+ $Y2=0
cc_210 N_A_27_297#_c_189_n A_411_47# 0.00542732f $X=2.125 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_211 N_A_27_297#_c_228_n A_411_47# 0.00559046f $X=2.21 $Y=0.735 $X2=-0.19
+ $Y2=-0.24
cc_212 N_A_27_297#_c_190_n A_411_47# 0.00158968f $X=2.845 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_213 N_A_27_297#_c_191_n A_411_47# 0.00269653f $X=2.295 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_214 N_A_117_297#_c_312_n N_VPWR_M1008_s 0.00553503f $X=2.13 $Y=1.915
+ $X2=-0.19 $Y2=1.305
cc_215 N_A_117_297#_c_312_n N_VPWR_c_336_n 0.0221579f $X=2.13 $Y=1.915 $X2=0
+ $Y2=0
cc_216 N_A_117_297#_c_327_p N_VPWR_c_336_n 0.0156675f $X=2.215 $Y=2.3 $X2=0
+ $Y2=0
cc_217 N_A_117_297#_c_312_n N_VPWR_c_340_n 0.00293436f $X=2.13 $Y=1.915 $X2=0
+ $Y2=0
cc_218 N_A_117_297#_c_327_p N_VPWR_c_340_n 0.0159953f $X=2.215 $Y=2.3 $X2=0
+ $Y2=0
cc_219 N_A_117_297#_c_312_n N_VPWR_c_342_n 0.00320421f $X=2.13 $Y=1.915 $X2=0
+ $Y2=0
cc_220 N_A_117_297#_M1005_d N_VPWR_c_335_n 0.00232895f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_221 N_A_117_297#_M1008_d N_VPWR_c_335_n 0.00367486f $X=2.045 $Y=1.485 $X2=0
+ $Y2=0
cc_222 N_A_117_297#_c_312_n N_VPWR_c_335_n 0.0133318f $X=2.13 $Y=1.915 $X2=0
+ $Y2=0
cc_223 N_A_117_297#_c_327_p N_VPWR_c_335_n 0.00954719f $X=2.215 $Y=2.3 $X2=0
+ $Y2=0
cc_224 N_VPWR_c_335_n N_X_M1001_d 0.00439555f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_225 N_VPWR_c_339_n X 0.0684531f $X=3.84 $Y=1.63 $X2=0 $Y2=0
cc_226 N_VPWR_c_337_n X 0.0381758f $X=2.765 $Y=1.96 $X2=0 $Y2=0
cc_227 N_VPWR_c_343_n X 0.0262891f $X=3.755 $Y=2.72 $X2=0 $Y2=0
cc_228 N_VPWR_c_335_n X 0.0148218f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_229 N_VPWR_c_339_n N_VGND_c_420_n 0.00786978f $X=3.84 $Y=1.63 $X2=0 $Y2=0
cc_230 N_X_c_405_n N_VGND_c_420_n 0.0489013f $X=3.235 $Y=0.42 $X2=0 $Y2=0
cc_231 N_X_c_405_n N_VGND_c_422_n 0.0258717f $X=3.235 $Y=0.42 $X2=0 $Y2=0
cc_232 N_X_M1002_s N_VGND_c_424_n 0.00428929f $X=3.1 $Y=0.235 $X2=0 $Y2=0
cc_233 N_X_c_405_n N_VGND_c_424_n 0.0149437f $X=3.235 $Y=0.42 $X2=0 $Y2=0
cc_234 N_VGND_c_424_n A_119_47# 0.00978874f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_235 N_VGND_c_424_n A_411_47# 0.00379705f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
