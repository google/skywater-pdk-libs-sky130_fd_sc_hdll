* File: sky130_fd_sc_hdll__o21bai_2.pxi.spice
* Created: Thu Aug 27 19:20:03 2020
* 
x_PM_SKY130_FD_SC_HDLL__O21BAI_2%B1_N N_B1_N_c_70_n N_B1_N_M1004_g N_B1_N_c_71_n
+ N_B1_N_M1003_g B1_N B1_N PM_SKY130_FD_SC_HDLL__O21BAI_2%B1_N
x_PM_SKY130_FD_SC_HDLL__O21BAI_2%A_28_297# N_A_28_297#_M1003_d
+ N_A_28_297#_M1004_s N_A_28_297#_c_103_n N_A_28_297#_M1005_g
+ N_A_28_297#_c_104_n N_A_28_297#_M1009_g N_A_28_297#_c_96_n N_A_28_297#_M1001_g
+ N_A_28_297#_c_97_n N_A_28_297#_M1002_g N_A_28_297#_c_109_n N_A_28_297#_c_98_n
+ N_A_28_297#_c_99_n N_A_28_297#_c_100_n N_A_28_297#_c_106_n N_A_28_297#_c_101_n
+ N_A_28_297#_c_102_n PM_SKY130_FD_SC_HDLL__O21BAI_2%A_28_297#
x_PM_SKY130_FD_SC_HDLL__O21BAI_2%A2 N_A2_c_163_n N_A2_M1006_g N_A2_c_167_n
+ N_A2_M1011_g N_A2_c_168_n N_A2_M1013_g N_A2_c_164_n N_A2_M1012_g A2
+ N_A2_c_166_n PM_SKY130_FD_SC_HDLL__O21BAI_2%A2
x_PM_SKY130_FD_SC_HDLL__O21BAI_2%A1 N_A1_c_214_n N_A1_M1000_g N_A1_c_218_n
+ N_A1_M1007_g N_A1_c_219_n N_A1_M1010_g N_A1_c_215_n N_A1_M1008_g A1
+ N_A1_c_216_n A1 PM_SKY130_FD_SC_HDLL__O21BAI_2%A1
x_PM_SKY130_FD_SC_HDLL__O21BAI_2%VPWR N_VPWR_M1004_d N_VPWR_M1009_d
+ N_VPWR_M1007_s N_VPWR_c_253_n N_VPWR_c_254_n N_VPWR_c_255_n N_VPWR_c_256_n
+ N_VPWR_c_257_n N_VPWR_c_258_n N_VPWR_c_259_n VPWR N_VPWR_c_260_n
+ N_VPWR_c_252_n N_VPWR_c_262_n PM_SKY130_FD_SC_HDLL__O21BAI_2%VPWR
x_PM_SKY130_FD_SC_HDLL__O21BAI_2%Y N_Y_M1001_s N_Y_M1005_s N_Y_M1011_s
+ N_Y_c_340_n N_Y_c_316_n N_Y_c_348_p N_Y_c_317_n Y N_Y_c_315_n Y
+ PM_SKY130_FD_SC_HDLL__O21BAI_2%Y
x_PM_SKY130_FD_SC_HDLL__O21BAI_2%A_437_297# N_A_437_297#_M1011_d
+ N_A_437_297#_M1013_d N_A_437_297#_M1010_d N_A_437_297#_c_355_n
+ N_A_437_297#_c_361_n N_A_437_297#_c_356_n N_A_437_297#_c_357_n
+ N_A_437_297#_c_380_n N_A_437_297#_c_358_n N_A_437_297#_c_359_n
+ N_A_437_297#_c_360_n PM_SKY130_FD_SC_HDLL__O21BAI_2%A_437_297#
x_PM_SKY130_FD_SC_HDLL__O21BAI_2%VGND N_VGND_M1003_s N_VGND_M1006_s
+ N_VGND_M1000_s N_VGND_c_395_n N_VGND_c_396_n N_VGND_c_397_n N_VGND_c_398_n
+ N_VGND_c_399_n N_VGND_c_400_n N_VGND_c_401_n N_VGND_c_402_n VGND
+ N_VGND_c_403_n N_VGND_c_404_n PM_SKY130_FD_SC_HDLL__O21BAI_2%VGND
x_PM_SKY130_FD_SC_HDLL__O21BAI_2%A_226_47# N_A_226_47#_M1001_d
+ N_A_226_47#_M1002_d N_A_226_47#_M1012_d N_A_226_47#_M1008_d
+ N_A_226_47#_c_459_n N_A_226_47#_c_460_n N_A_226_47#_c_472_n
+ N_A_226_47#_c_475_n N_A_226_47#_c_461_n N_A_226_47#_c_462_n
+ N_A_226_47#_c_483_n N_A_226_47#_c_463_n N_A_226_47#_c_464_n
+ N_A_226_47#_c_465_n PM_SKY130_FD_SC_HDLL__O21BAI_2%A_226_47#
cc_1 VNB N_B1_N_c_70_n 0.0391278f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_2 VNB N_B1_N_c_71_n 0.0216313f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_3 VNB B1_N 0.0151337f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.19
cc_4 VNB N_A_28_297#_c_96_n 0.0199367f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_28_297#_c_97_n 0.0166801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_28_297#_c_98_n 0.0083295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_28_297#_c_99_n 0.00108972f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_28_297#_c_100_n 9.61753e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_28_297#_c_101_n 0.0053919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_28_297#_c_102_n 0.0755054f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A2_c_163_n 0.0169271f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_12 VNB N_A2_c_164_n 0.0169324f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_13 VNB A2 0.0121984f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A2_c_166_n 0.0359564f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A1_c_214_n 0.0169324f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_16 VNB N_A1_c_215_n 0.0223965f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_17 VNB N_A1_c_216_n 0.0430121f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB A1 0.020968f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_252_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_315_n 0.00474942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_395_n 0.0112126f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_22 VNB N_VGND_c_396_n 0.018448f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_23 VNB N_VGND_c_397_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_398_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_399_n 0.058968f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_400_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_401_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_402_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_403_n 0.0230835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_404_n 0.267585f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_226_47#_c_459_n 0.00618298f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_226_47#_c_460_n 0.00633933f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.19
cc_33 VNB N_A_226_47#_c_461_n 0.00221554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_226_47#_c_462_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_226_47#_c_463_n 0.0139603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_226_47#_c_464_n 0.0186133f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_226_47#_c_465_n 0.00253348f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VPB N_B1_N_c_70_n 0.0398113f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_39 VPB B1_N 0.00407848f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.19
cc_40 VPB N_A_28_297#_c_103_n 0.0182655f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_41 VPB N_A_28_297#_c_104_n 0.0193978f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.16
cc_42 VPB N_A_28_297#_c_99_n 0.00356026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_28_297#_c_106_n 0.00362304f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_28_297#_c_102_n 0.0389537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A2_c_167_n 0.0193736f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=0.995
cc_46 VPB N_A2_c_168_n 0.01642f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_47 VPB N_A2_c_166_n 0.0212542f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A1_c_218_n 0.0156552f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=0.995
cc_49 VPB N_A1_c_219_n 0.0201729f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_50 VPB N_A1_c_216_n 0.022695f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_253_n 0.0215305f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.16
cc_52 VPB N_VPWR_c_254_n 0.0106018f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_255_n 4.89699e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_256_n 0.0181525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_257_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_258_n 0.0390623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_259_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_260_n 0.0212809f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_252_n 0.0730686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_262_n 0.0274883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_Y_c_316_n 0.0111041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_Y_c_317_n 0.0081557f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_Y_c_315_n 0.00165176f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_437_297#_c_355_n 0.00610594f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.16
cc_65 VPB N_A_437_297#_c_356_n 0.00247174f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.19
cc_66 VPB N_A_437_297#_c_357_n 0.00188871f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_437_297#_c_358_n 0.00290609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_437_297#_c_359_n 0.0116576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_437_297#_c_360_n 0.0307403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 N_B1_N_c_70_n N_A_28_297#_c_103_n 0.0142472f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_71 N_B1_N_c_70_n N_A_28_297#_c_109_n 0.0195698f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_72 B1_N N_A_28_297#_c_109_n 0.00735917f $X=0.36 $Y=1.19 $X2=0 $Y2=0
cc_73 N_B1_N_c_71_n N_A_28_297#_c_98_n 0.00604734f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_74 B1_N N_A_28_297#_c_98_n 0.00601073f $X=0.36 $Y=1.19 $X2=0 $Y2=0
cc_75 N_B1_N_c_70_n N_A_28_297#_c_99_n 0.00534646f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_76 B1_N N_A_28_297#_c_99_n 0.00621616f $X=0.36 $Y=1.19 $X2=0 $Y2=0
cc_77 N_B1_N_c_70_n N_A_28_297#_c_106_n 0.00864563f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_78 B1_N N_A_28_297#_c_106_n 0.0133535f $X=0.36 $Y=1.19 $X2=0 $Y2=0
cc_79 N_B1_N_c_70_n N_A_28_297#_c_101_n 0.00172703f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_80 B1_N N_A_28_297#_c_101_n 0.0146005f $X=0.36 $Y=1.19 $X2=0 $Y2=0
cc_81 N_B1_N_c_70_n N_A_28_297#_c_102_n 0.0133915f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_82 N_B1_N_c_70_n N_VPWR_c_253_n 0.00370547f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_83 N_B1_N_c_70_n N_VPWR_c_252_n 0.00500987f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_84 N_B1_N_c_70_n N_VPWR_c_262_n 0.00393512f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_85 N_B1_N_c_70_n N_VGND_c_396_n 0.00391367f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_86 N_B1_N_c_71_n N_VGND_c_396_n 0.00602843f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_87 B1_N N_VGND_c_396_n 0.0138735f $X=0.36 $Y=1.19 $X2=0 $Y2=0
cc_88 N_B1_N_c_71_n N_VGND_c_399_n 0.00510437f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_89 N_B1_N_c_71_n N_VGND_c_404_n 0.00512902f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_90 N_B1_N_c_71_n N_A_226_47#_c_459_n 0.00340559f $X=0.525 $Y=0.995 $X2=0
+ $Y2=0
cc_91 N_A_28_297#_c_97_n N_A2_c_163_n 0.0146683f $X=2.1 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_92 N_A_28_297#_c_102_n A2 0.00215915f $X=1.63 $Y=1.202 $X2=0 $Y2=0
cc_93 N_A_28_297#_c_102_n N_A2_c_166_n 0.0146683f $X=1.63 $Y=1.202 $X2=0 $Y2=0
cc_94 N_A_28_297#_c_109_n N_VPWR_M1004_d 0.0039833f $X=0.65 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_95 N_A_28_297#_c_103_n N_VPWR_c_253_n 0.0127297f $X=1.035 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A_28_297#_c_104_n N_VPWR_c_253_n 6.39761e-19 $X=1.505 $Y=1.41 $X2=0
+ $Y2=0
cc_97 N_A_28_297#_c_109_n N_VPWR_c_253_n 0.0182266f $X=0.65 $Y=1.58 $X2=0 $Y2=0
cc_98 N_A_28_297#_c_100_n N_VPWR_c_253_n 8.7362e-19 $X=1.175 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_28_297#_c_106_n N_VPWR_c_253_n 0.00126814f $X=0.265 $Y=1.58 $X2=0
+ $Y2=0
cc_100 N_A_28_297#_c_104_n N_VPWR_c_254_n 0.00341296f $X=1.505 $Y=1.41 $X2=0
+ $Y2=0
cc_101 N_A_28_297#_c_102_n N_VPWR_c_254_n 9.86422e-19 $X=1.63 $Y=1.202 $X2=0
+ $Y2=0
cc_102 N_A_28_297#_c_103_n N_VPWR_c_256_n 0.00622633f $X=1.035 $Y=1.41 $X2=0
+ $Y2=0
cc_103 N_A_28_297#_c_104_n N_VPWR_c_256_n 0.00702461f $X=1.505 $Y=1.41 $X2=0
+ $Y2=0
cc_104 N_A_28_297#_c_103_n N_VPWR_c_252_n 0.0104011f $X=1.035 $Y=1.41 $X2=0
+ $Y2=0
cc_105 N_A_28_297#_c_104_n N_VPWR_c_252_n 0.0137041f $X=1.505 $Y=1.41 $X2=0
+ $Y2=0
cc_106 N_A_28_297#_c_106_n N_VPWR_c_252_n 0.00647432f $X=0.265 $Y=1.58 $X2=0
+ $Y2=0
cc_107 N_A_28_297#_c_102_n N_Y_c_316_n 0.00743111f $X=1.63 $Y=1.202 $X2=0 $Y2=0
cc_108 N_A_28_297#_c_103_n N_Y_c_317_n 0.00116321f $X=1.035 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A_28_297#_c_104_n N_Y_c_317_n 0.0198117f $X=1.505 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A_28_297#_c_99_n N_Y_c_317_n 0.0028058f $X=0.782 $Y=1.495 $X2=0 $Y2=0
cc_111 N_A_28_297#_c_100_n N_Y_c_317_n 0.0110727f $X=1.175 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_28_297#_c_102_n N_Y_c_317_n 0.00706074f $X=1.63 $Y=1.202 $X2=0 $Y2=0
cc_113 N_A_28_297#_c_104_n N_Y_c_315_n 0.00148689f $X=1.505 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_28_297#_c_96_n N_Y_c_315_n 0.0134547f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A_28_297#_c_97_n N_Y_c_315_n 0.00299628f $X=2.1 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A_28_297#_c_99_n N_Y_c_315_n 0.00610543f $X=0.782 $Y=1.495 $X2=0 $Y2=0
cc_117 N_A_28_297#_c_100_n N_Y_c_315_n 0.0138315f $X=1.175 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_28_297#_c_102_n N_Y_c_315_n 0.0447722f $X=1.63 $Y=1.202 $X2=0 $Y2=0
cc_119 N_A_28_297#_c_98_n N_VGND_c_396_n 0.00959344f $X=0.735 $Y=0.66 $X2=0
+ $Y2=0
cc_120 N_A_28_297#_c_96_n N_VGND_c_399_n 0.00357877f $X=1.63 $Y=0.995 $X2=0
+ $Y2=0
cc_121 N_A_28_297#_c_97_n N_VGND_c_399_n 0.00357877f $X=2.1 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A_28_297#_c_98_n N_VGND_c_399_n 0.00542302f $X=0.735 $Y=0.66 $X2=0
+ $Y2=0
cc_123 N_A_28_297#_c_96_n N_VGND_c_404_n 0.00677297f $X=1.63 $Y=0.995 $X2=0
+ $Y2=0
cc_124 N_A_28_297#_c_97_n N_VGND_c_404_n 0.00538422f $X=2.1 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_28_297#_c_98_n N_VGND_c_404_n 0.00578545f $X=0.735 $Y=0.66 $X2=0
+ $Y2=0
cc_126 N_A_28_297#_c_98_n N_A_226_47#_c_459_n 0.00197505f $X=0.735 $Y=0.66 $X2=0
+ $Y2=0
cc_127 N_A_28_297#_c_96_n N_A_226_47#_c_460_n 0.00757452f $X=1.63 $Y=0.995 $X2=0
+ $Y2=0
cc_128 N_A_28_297#_c_98_n N_A_226_47#_c_460_n 0.0258345f $X=0.735 $Y=0.66 $X2=0
+ $Y2=0
cc_129 N_A_28_297#_c_100_n N_A_226_47#_c_460_n 0.0223399f $X=1.175 $Y=1.16 $X2=0
+ $Y2=0
cc_130 N_A_28_297#_c_102_n N_A_226_47#_c_460_n 0.00740214f $X=1.63 $Y=1.202
+ $X2=0 $Y2=0
cc_131 N_A_28_297#_c_96_n N_A_226_47#_c_472_n 0.0142483f $X=1.63 $Y=0.995 $X2=0
+ $Y2=0
cc_132 N_A_28_297#_c_97_n N_A_226_47#_c_472_n 0.0140389f $X=2.1 $Y=0.995 $X2=0
+ $Y2=0
cc_133 N_A_28_297#_c_102_n N_A_226_47#_c_472_n 0.00514929f $X=1.63 $Y=1.202
+ $X2=0 $Y2=0
cc_134 N_A2_c_164_n N_A1_c_214_n 0.0176256f $X=3.04 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_135 N_A2_c_168_n N_A1_c_218_n 0.00966756f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_136 A2 N_A1_c_216_n 0.00578274f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_137 N_A2_c_166_n N_A1_c_216_n 0.0176256f $X=3.015 $Y=1.202 $X2=0 $Y2=0
cc_138 A2 A1 0.0136085f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_139 N_A2_c_167_n N_VPWR_c_254_n 0.0019773f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A2_c_168_n N_VPWR_c_255_n 0.00110692f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A2_c_167_n N_VPWR_c_258_n 0.00429453f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A2_c_168_n N_VPWR_c_258_n 0.00429453f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A2_c_167_n N_VPWR_c_252_n 0.00734734f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A2_c_168_n N_VPWR_c_252_n 0.00609021f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A2_c_167_n N_Y_c_316_n 0.0176655f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A2_c_168_n N_Y_c_316_n 6.53978e-19 $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_147 A2 N_Y_c_316_n 0.0550513f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_148 N_A2_c_166_n N_Y_c_316_n 0.00717692f $X=3.015 $Y=1.202 $X2=0 $Y2=0
cc_149 N_A2_c_167_n N_Y_c_315_n 0.00100699f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_150 A2 N_Y_c_315_n 0.0162828f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_151 N_A2_c_166_n N_Y_c_315_n 0.00339447f $X=3.015 $Y=1.202 $X2=0 $Y2=0
cc_152 N_A2_c_167_n N_A_437_297#_c_361_n 0.0143148f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A2_c_168_n N_A_437_297#_c_361_n 0.0143578f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A2_c_168_n N_A_437_297#_c_357_n 0.00132962f $X=3.015 $Y=1.41 $X2=0
+ $Y2=0
cc_155 A2 N_A_437_297#_c_357_n 0.0139423f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_156 A2 N_A_437_297#_c_358_n 0.0040358f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_157 N_A2_c_163_n N_VGND_c_397_n 0.00385178f $X=2.52 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A2_c_164_n N_VGND_c_397_n 0.00365402f $X=3.04 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A2_c_163_n N_VGND_c_399_n 0.00421816f $X=2.52 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A2_c_164_n N_VGND_c_401_n 0.00396605f $X=3.04 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A2_c_163_n N_VGND_c_404_n 0.00611766f $X=2.52 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A2_c_164_n N_VGND_c_404_n 0.00583042f $X=3.04 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A2_c_163_n N_A_226_47#_c_475_n 0.00284788f $X=2.52 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A2_c_163_n N_A_226_47#_c_461_n 0.00518775f $X=2.52 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A2_c_164_n N_A_226_47#_c_461_n 4.72003e-19 $X=3.04 $Y=0.995 $X2=0 $Y2=0
cc_166 A2 N_A_226_47#_c_461_n 0.0210224f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_167 N_A2_c_163_n N_A_226_47#_c_462_n 0.00929182f $X=2.52 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A2_c_164_n N_A_226_47#_c_462_n 0.00650032f $X=3.04 $Y=0.995 $X2=0 $Y2=0
cc_169 A2 N_A_226_47#_c_462_n 0.0399344f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_170 N_A2_c_166_n N_A_226_47#_c_462_n 0.00468948f $X=3.015 $Y=1.202 $X2=0
+ $Y2=0
cc_171 N_A2_c_163_n N_A_226_47#_c_483_n 5.69266e-19 $X=2.52 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A2_c_164_n N_A_226_47#_c_483_n 0.00857123f $X=3.04 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A2_c_164_n N_A_226_47#_c_465_n 0.00269873f $X=3.04 $Y=0.995 $X2=0 $Y2=0
cc_174 A2 N_A_226_47#_c_465_n 0.0294984f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_175 N_A1_c_218_n N_VPWR_c_255_n 0.0163934f $X=3.485 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A1_c_219_n N_VPWR_c_255_n 0.0135516f $X=3.955 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A1_c_218_n N_VPWR_c_258_n 0.00427505f $X=3.485 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A1_c_219_n N_VPWR_c_260_n 0.00622633f $X=3.955 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A1_c_218_n N_VPWR_c_252_n 0.00735499f $X=3.485 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A1_c_219_n N_VPWR_c_252_n 0.0114251f $X=3.955 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A1_c_218_n N_A_437_297#_c_358_n 0.0170057f $X=3.485 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A1_c_219_n N_A_437_297#_c_358_n 0.0166678f $X=3.955 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A1_c_216_n N_A_437_297#_c_358_n 0.00815835f $X=3.955 $Y=1.202 $X2=0
+ $Y2=0
cc_184 A1 N_A_437_297#_c_358_n 0.0343628f $X=3.815 $Y=1.19 $X2=0 $Y2=0
cc_185 A1 N_A_437_297#_c_359_n 0.0225537f $X=3.815 $Y=1.19 $X2=0 $Y2=0
cc_186 N_A1_c_214_n N_VGND_c_398_n 0.00385467f $X=3.46 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A1_c_215_n N_VGND_c_398_n 0.00381583f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A1_c_214_n N_VGND_c_401_n 0.00423334f $X=3.46 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A1_c_215_n N_VGND_c_403_n 0.00397706f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A1_c_214_n N_VGND_c_404_n 0.00610858f $X=3.46 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A1_c_215_n N_VGND_c_404_n 0.00687453f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A1_c_214_n N_A_226_47#_c_483_n 0.00693563f $X=3.46 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A1_c_215_n N_A_226_47#_c_483_n 5.34196e-19 $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A1_c_214_n N_A_226_47#_c_463_n 0.0107693f $X=3.46 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A1_c_215_n N_A_226_47#_c_463_n 0.00937294f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A1_c_216_n N_A_226_47#_c_463_n 0.00468948f $X=3.955 $Y=1.202 $X2=0
+ $Y2=0
cc_197 A1 N_A_226_47#_c_463_n 0.0599937f $X=3.815 $Y=1.19 $X2=0 $Y2=0
cc_198 N_A1_c_214_n N_A_226_47#_c_464_n 5.66376e-19 $X=3.46 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A1_c_215_n N_A_226_47#_c_464_n 0.0084675f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A1_c_214_n N_A_226_47#_c_465_n 0.00142536f $X=3.46 $Y=0.995 $X2=0 $Y2=0
cc_201 N_VPWR_c_252_n N_Y_M1005_s 0.00647849f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_202 N_VPWR_c_252_n N_Y_M1011_s 0.00232895f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_203 N_VPWR_c_253_n N_Y_c_340_n 0.0357198f $X=0.8 $Y=1.96 $X2=0 $Y2=0
cc_204 N_VPWR_c_256_n N_Y_c_340_n 0.0118139f $X=1.62 $Y=2.72 $X2=0 $Y2=0
cc_205 N_VPWR_c_252_n N_Y_c_340_n 0.00646998f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_206 N_VPWR_M1009_d N_Y_c_317_n 0.00291581f $X=1.595 $Y=1.485 $X2=0 $Y2=0
cc_207 N_VPWR_c_254_n N_Y_c_317_n 0.0187556f $X=1.74 $Y=1.96 $X2=0 $Y2=0
cc_208 N_VPWR_c_252_n N_A_437_297#_M1011_d 0.00217519f $X=4.37 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_209 N_VPWR_c_252_n N_A_437_297#_M1013_d 0.00436089f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_210 N_VPWR_c_252_n N_A_437_297#_M1010_d 0.00442207f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_211 N_VPWR_c_254_n N_A_437_297#_c_355_n 0.0324951f $X=1.74 $Y=1.96 $X2=0
+ $Y2=0
cc_212 N_VPWR_c_258_n N_A_437_297#_c_361_n 0.0400924f $X=3.505 $Y=2.72 $X2=0
+ $Y2=0
cc_213 N_VPWR_c_252_n N_A_437_297#_c_361_n 0.0253962f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_214 N_VPWR_c_254_n N_A_437_297#_c_356_n 0.0117483f $X=1.74 $Y=1.96 $X2=0
+ $Y2=0
cc_215 N_VPWR_c_258_n N_A_437_297#_c_356_n 0.0220041f $X=3.505 $Y=2.72 $X2=0
+ $Y2=0
cc_216 N_VPWR_c_252_n N_A_437_297#_c_356_n 0.0127039f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_217 N_VPWR_c_255_n N_A_437_297#_c_380_n 0.0484833f $X=3.72 $Y=2 $X2=0 $Y2=0
cc_218 N_VPWR_c_258_n N_A_437_297#_c_380_n 0.0119545f $X=3.505 $Y=2.72 $X2=0
+ $Y2=0
cc_219 N_VPWR_c_252_n N_A_437_297#_c_380_n 0.006547f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_220 N_VPWR_M1007_s N_A_437_297#_c_358_n 0.00188315f $X=3.575 $Y=1.485 $X2=0
+ $Y2=0
cc_221 N_VPWR_c_255_n N_A_437_297#_c_358_n 0.0212439f $X=3.72 $Y=2 $X2=0 $Y2=0
cc_222 N_VPWR_c_255_n N_A_437_297#_c_360_n 0.0399729f $X=3.72 $Y=2 $X2=0 $Y2=0
cc_223 N_VPWR_c_260_n N_A_437_297#_c_360_n 0.019258f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_224 N_VPWR_c_252_n N_A_437_297#_c_360_n 0.0105137f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_225 N_Y_c_316_n N_A_437_297#_M1011_d 0.00296183f $X=2.655 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_226 N_Y_c_316_n N_A_437_297#_c_355_n 0.0229833f $X=2.655 $Y=1.53 $X2=0 $Y2=0
cc_227 N_Y_M1011_s N_A_437_297#_c_361_n 0.00352392f $X=2.635 $Y=1.485 $X2=0
+ $Y2=0
cc_228 N_Y_c_348_p N_A_437_297#_c_361_n 0.0134104f $X=2.78 $Y=1.62 $X2=0 $Y2=0
cc_229 N_Y_c_316_n N_A_437_297#_c_357_n 0.00623033f $X=2.655 $Y=1.53 $X2=0 $Y2=0
cc_230 N_Y_M1001_s N_VGND_c_404_n 0.00256987f $X=1.705 $Y=0.235 $X2=0 $Y2=0
cc_231 N_Y_c_315_n N_A_226_47#_c_460_n 0.0110448f $X=1.84 $Y=0.73 $X2=0 $Y2=0
cc_232 N_Y_M1001_s N_A_226_47#_c_472_n 0.00399909f $X=1.705 $Y=0.235 $X2=0 $Y2=0
cc_233 N_Y_c_315_n N_A_226_47#_c_472_n 0.0271308f $X=1.84 $Y=0.73 $X2=0 $Y2=0
cc_234 N_Y_c_315_n N_A_226_47#_c_461_n 0.00144197f $X=1.84 $Y=0.73 $X2=0 $Y2=0
cc_235 N_A_437_297#_c_358_n N_A_226_47#_c_463_n 0.00554576f $X=4.105 $Y=1.56
+ $X2=0 $Y2=0
cc_236 N_A_437_297#_c_358_n N_A_226_47#_c_465_n 7.50318e-19 $X=4.105 $Y=1.56
+ $X2=0 $Y2=0
cc_237 N_VGND_c_404_n N_A_226_47#_M1001_d 0.00345409f $X=4.37 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_238 N_VGND_c_404_n N_A_226_47#_M1002_d 0.00215206f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_239 N_VGND_c_404_n N_A_226_47#_M1012_d 0.00215201f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_240 N_VGND_c_404_n N_A_226_47#_M1008_d 0.00226063f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_241 N_VGND_c_399_n N_A_226_47#_c_459_n 0.0197205f $X=2.695 $Y=0 $X2=0 $Y2=0
cc_242 N_VGND_c_404_n N_A_226_47#_c_459_n 0.0107706f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_243 N_VGND_c_399_n N_A_226_47#_c_472_n 0.0499893f $X=2.695 $Y=0 $X2=0 $Y2=0
cc_244 N_VGND_c_404_n N_A_226_47#_c_472_n 0.0317007f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_245 N_VGND_c_397_n N_A_226_47#_c_475_n 0.0141571f $X=2.78 $Y=0.39 $X2=0 $Y2=0
cc_246 N_VGND_c_399_n N_A_226_47#_c_475_n 0.0152108f $X=2.695 $Y=0 $X2=0 $Y2=0
cc_247 N_VGND_c_404_n N_A_226_47#_c_475_n 0.00940698f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_248 N_VGND_c_397_n N_A_226_47#_c_461_n 0.00471242f $X=2.78 $Y=0.39 $X2=0
+ $Y2=0
cc_249 N_VGND_M1006_s N_A_226_47#_c_462_n 0.00348805f $X=2.595 $Y=0.235 $X2=0
+ $Y2=0
cc_250 N_VGND_c_397_n N_A_226_47#_c_462_n 0.0131987f $X=2.78 $Y=0.39 $X2=0 $Y2=0
cc_251 N_VGND_c_399_n N_A_226_47#_c_462_n 0.00266636f $X=2.695 $Y=0 $X2=0 $Y2=0
cc_252 N_VGND_c_401_n N_A_226_47#_c_462_n 0.00199443f $X=3.635 $Y=0 $X2=0 $Y2=0
cc_253 N_VGND_c_404_n N_A_226_47#_c_462_n 0.0100158f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_254 N_VGND_c_397_n N_A_226_47#_c_483_n 0.0223967f $X=2.78 $Y=0.39 $X2=0 $Y2=0
cc_255 N_VGND_c_398_n N_A_226_47#_c_483_n 0.0183628f $X=3.72 $Y=0.39 $X2=0 $Y2=0
cc_256 N_VGND_c_401_n N_A_226_47#_c_483_n 0.0222529f $X=3.635 $Y=0 $X2=0 $Y2=0
cc_257 N_VGND_c_404_n N_A_226_47#_c_483_n 0.0139016f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_258 N_VGND_M1000_s N_A_226_47#_c_463_n 0.00348805f $X=3.535 $Y=0.235 $X2=0
+ $Y2=0
cc_259 N_VGND_c_398_n N_A_226_47#_c_463_n 0.0131987f $X=3.72 $Y=0.39 $X2=0 $Y2=0
cc_260 N_VGND_c_401_n N_A_226_47#_c_463_n 0.00266636f $X=3.635 $Y=0 $X2=0 $Y2=0
cc_261 N_VGND_c_403_n N_A_226_47#_c_463_n 0.00199443f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_262 N_VGND_c_404_n N_A_226_47#_c_463_n 0.0100158f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_263 N_VGND_c_398_n N_A_226_47#_c_464_n 0.021759f $X=3.72 $Y=0.39 $X2=0 $Y2=0
cc_264 N_VGND_c_403_n N_A_226_47#_c_464_n 0.0245357f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_265 N_VGND_c_404_n N_A_226_47#_c_464_n 0.0149859f $X=4.37 $Y=0 $X2=0 $Y2=0
