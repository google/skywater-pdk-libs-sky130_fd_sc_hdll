* File: sky130_fd_sc_hdll__nand4b_2.pex.spice
* Created: Wed Sep  2 08:38:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND4B_2%A_N 2 3 5 8 10 11 19
c31 10 0 1.09696e-19 $X=0.235 $Y=1.19
r32 18 19 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r33 15 18 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.495 $Y2=1.16
r34 10 11 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.16
+ $X2=0.21 $Y2=1.53
r35 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r36 6 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.16
r37 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r38 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r39 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.89 $X2=0.495
+ $Y2=1.99
r40 1 18 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r41 1 2 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_2%A_27_47# 1 2 7 9 10 12 13 15 16 18 19 22
+ 26 30 32 33 35 38 49
c89 19 0 1.09696e-19 $X=1.385 $Y=1.16
c90 16 0 1.05021e-19 $X=1.98 $Y=0.995
r91 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.16 $X2=1.17 $Y2=1.16
r92 36 49 2.28545 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.16 $X2=0.61
+ $Y2=1.16
r93 36 38 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.72 $Y=1.16
+ $X2=1.17 $Y2=1.16
r94 34 49 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=1.245
+ $X2=0.61 $Y2=1.16
r95 34 35 35.0971 $w=2.18e-07 $l=6.7e-07 $layer=LI1_cond $X=0.61 $Y=1.245
+ $X2=0.61 $Y2=1.915
r96 33 49 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=1.075
+ $X2=0.61 $Y2=1.16
r97 32 33 14.1436 $w=2.18e-07 $l=2.7e-07 $layer=LI1_cond $X=0.61 $Y=0.805
+ $X2=0.61 $Y2=1.075
r98 28 35 25.6396 $w=1.68e-07 $l=3.93e-07 $layer=LI1_cond $X=0.217 $Y=2 $X2=0.61
+ $Y2=2
r99 28 30 9.26474 $w=2.53e-07 $l=2.05e-07 $layer=LI1_cond $X=0.217 $Y=2.085
+ $X2=0.217 $Y2=2.29
r100 24 32 25.6396 $w=1.68e-07 $l=3.93e-07 $layer=LI1_cond $X=0.217 $Y=0.72
+ $X2=0.61 $Y2=0.72
r101 24 26 9.26474 $w=2.53e-07 $l=2.05e-07 $layer=LI1_cond $X=0.217 $Y=0.635
+ $X2=0.217 $Y2=0.43
r102 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.955 $Y=1.202
+ $X2=1.98 $Y2=1.202
r103 21 22 56.4447 $w=3.8e-07 $l=4.45e-07 $layer=POLY_cond $X=1.51 $Y=1.202
+ $X2=1.955 $Y2=1.202
r104 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.485 $Y=1.202
+ $X2=1.51 $Y2=1.202
r105 19 39 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.385 $Y=1.16
+ $X2=1.17 $Y2=1.16
r106 19 20 13.6483 $w=3.8e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.385 $Y=1.16
+ $X2=1.485 $Y2=1.202
r107 16 23 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.98 $Y=0.995
+ $X2=1.98 $Y2=1.202
r108 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.98 $Y=0.995
+ $X2=1.98 $Y2=0.56
r109 13 22 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.202
r110 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.985
r111 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=1.202
r112 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=0.56
r113 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.202
r114 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.985
r115 2 30 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.29
r116 1 26 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_2%B 1 3 4 6 7 9 10 12 13 14 20 23 27 29
c49 4 0 1.55098e-19 $X=2.425 $Y=1.41
r50 27 29 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=2.555 $Y=1.175
+ $X2=3.015 $Y2=1.175
r51 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.115
+ $Y=1.16 $X2=3.115 $Y2=1.16
r52 20 22 29.0521 $w=3.65e-07 $l=2.2e-07 $layer=POLY_cond $X=2.895 $Y=1.202
+ $X2=3.115 $Y2=1.202
r53 19 20 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=2.87 $Y=1.202
+ $X2=2.895 $Y2=1.202
r54 18 19 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=2.425 $Y=1.202
+ $X2=2.87 $Y2=1.202
r55 17 18 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=2.4 $Y=1.202
+ $X2=2.425 $Y2=1.202
r56 14 23 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=3.02 $Y=1.175
+ $X2=3.115 $Y2=1.175
r57 14 29 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=3.02 $Y=1.175
+ $X2=3.015 $Y2=1.175
r58 13 27 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=2.54 $Y=1.175
+ $X2=2.555 $Y2=1.175
r59 10 20 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.202
r60 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.985
r61 7 19 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.87 $Y=0.995
+ $X2=2.87 $Y2=1.202
r62 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.87 $Y=0.995 $X2=2.87
+ $Y2=0.56
r63 4 18 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.202
r64 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.985
r65 1 17 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.4 $Y=0.995 $X2=2.4
+ $Y2=1.202
r66 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.4 $Y=0.995 $X2=2.4
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_2%C 1 3 4 6 7 9 10 12 13 14 21 27 30
c47 21 0 1.44136e-19 $X=4.32 $Y=1.16
r48 21 23 7.79515 $w=3.71e-07 $l=6e-08 $layer=POLY_cond $X=4.32 $Y=1.202
+ $X2=4.38 $Y2=1.202
r49 19 21 1.94879 $w=3.71e-07 $l=1.5e-08 $layer=POLY_cond $X=4.305 $Y=1.202
+ $X2=4.32 $Y2=1.202
r50 18 19 51.3181 $w=3.71e-07 $l=3.95e-07 $layer=POLY_cond $X=3.91 $Y=1.202
+ $X2=4.305 $Y2=1.202
r51 17 18 9.74394 $w=3.71e-07 $l=7.5e-08 $layer=POLY_cond $X=3.835 $Y=1.202
+ $X2=3.91 $Y2=1.202
r52 14 30 2.49545 $w=1.98e-07 $l=4.5e-08 $layer=LI1_cond $X=4.32 $Y=1.175
+ $X2=4.365 $Y2=1.175
r53 14 27 23.0136 $w=1.98e-07 $l=4.15e-07 $layer=LI1_cond $X=4.32 $Y=1.175
+ $X2=3.905 $Y2=1.175
r54 14 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.32
+ $Y=1.16 $X2=4.32 $Y2=1.16
r55 13 27 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=3.9 $Y=1.175
+ $X2=3.905 $Y2=1.175
r56 10 23 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.38 $Y=0.995
+ $X2=4.38 $Y2=1.202
r57 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.38 $Y=0.995
+ $X2=4.38 $Y2=0.56
r58 7 19 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.202
r59 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.985
r60 4 18 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.91 $Y=0.995
+ $X2=3.91 $Y2=1.202
r61 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.91 $Y=0.995 $X2=3.91
+ $Y2=0.56
r62 1 17 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.202
r63 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_2%D 1 3 4 6 7 9 10 12 13 18 19 23 29 31
c45 19 0 1.44136e-19 $X=5.65 $Y=1.105
r46 29 31 22.7364 $w=1.98e-07 $l=4.1e-07 $layer=LI1_cond $X=5.285 $Y=1.175
+ $X2=5.695 $Y2=1.175
r47 23 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.695
+ $Y=1.16 $X2=5.695 $Y2=1.16
r48 19 31 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=5.735 $Y=1.175
+ $X2=5.695 $Y2=1.175
r49 18 29 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=5.265 $Y=1.175
+ $X2=5.285 $Y2=1.175
r50 16 17 9.58886 $w=3.77e-07 $l=7.5e-08 $layer=POLY_cond $X=5.335 $Y=1.202
+ $X2=5.41 $Y2=1.202
r51 15 16 50.5013 $w=3.77e-07 $l=3.95e-07 $layer=POLY_cond $X=4.94 $Y=1.202
+ $X2=5.335 $Y2=1.202
r52 14 15 9.58886 $w=3.77e-07 $l=7.5e-08 $layer=POLY_cond $X=4.865 $Y=1.202
+ $X2=4.94 $Y2=1.202
r53 13 23 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.485 $Y=1.16
+ $X2=5.695 $Y2=1.16
r54 13 17 10.4633 $w=3.77e-07 $l=9.3675e-08 $layer=POLY_cond $X=5.485 $Y=1.16
+ $X2=5.41 $Y2=1.202
r55 10 17 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.41 $Y=0.995
+ $X2=5.41 $Y2=1.202
r56 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.41 $Y=0.995
+ $X2=5.41 $Y2=0.56
r57 7 16 20.0566 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.335 $Y=1.41
+ $X2=5.335 $Y2=1.202
r58 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.335 $Y=1.41
+ $X2=5.335 $Y2=1.985
r59 4 15 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.94 $Y=0.995
+ $X2=4.94 $Y2=1.202
r60 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.94 $Y=0.995 $X2=4.94
+ $Y2=0.56
r61 1 14 20.0566 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.865 $Y=1.41
+ $X2=4.865 $Y2=1.202
r62 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.865 $Y=1.41
+ $X2=4.865 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_2%VPWR 1 2 3 4 5 6 19 20 23 27 31 35 37 39
+ 46 48 49 51 52 53 63 71 76 80 84
r91 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r92 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r93 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r94 74 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r95 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r96 71 83 5.38443 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=5.485 $Y=2.72
+ $X2=5.732 $Y2=2.72
r97 71 73 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.485 $Y=2.72
+ $X2=5.29 $Y2=2.72
r98 70 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r99 70 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.45 $Y2=2.72
r100 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r101 67 80 13.0174 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=3.365 $Y2=2.72
r102 67 69 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=4.37 $Y2=2.72
r103 66 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r104 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r105 63 80 13.0174 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=3.045 $Y=2.72
+ $X2=3.365 $Y2=2.72
r106 63 65 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.045 $Y=2.72
+ $X2=2.99 $Y2=2.72
r107 62 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r108 62 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r109 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r110 59 76 3.7769 $w=3.6e-07 $l=2.44643e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.21 $Y2=2.53
r111 59 61 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=2.07 $Y2=2.72
r112 53 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r113 53 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r114 51 69 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=2.72
+ $X2=4.37 $Y2=2.72
r115 51 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.455 $Y=2.72
+ $X2=4.585 $Y2=2.72
r116 50 73 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=4.715 $Y=2.72
+ $X2=5.29 $Y2=2.72
r117 50 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.715 $Y=2.72
+ $X2=4.585 $Y2=2.72
r118 48 61 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.07 $Y2=2.72
r119 48 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.19 $Y2=2.72
r120 47 65 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.99 $Y2=2.72
r121 47 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.19 $Y2=2.72
r122 46 56 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r123 45 46 10.9193 $w=5.48e-07 $l=2.15e-07 $layer=LI1_cond $X=0.73 $Y=2.53
+ $X2=0.515 $Y2=2.53
r124 39 42 19.8395 $w=3.93e-07 $l=6.8e-07 $layer=LI1_cond $X=5.682 $Y=1.66
+ $X2=5.682 $Y2=2.34
r125 37 83 2.94291 $w=3.95e-07 $l=1.07121e-07 $layer=LI1_cond $X=5.682 $Y=2.635
+ $X2=5.732 $Y2=2.72
r126 37 42 8.60685 $w=3.93e-07 $l=2.95e-07 $layer=LI1_cond $X=5.682 $Y=2.635
+ $X2=5.682 $Y2=2.34
r127 33 52 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.585 $Y=2.635
+ $X2=4.585 $Y2=2.72
r128 33 35 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=4.585 $Y=2.635
+ $X2=4.585 $Y2=2
r129 29 80 2.66764 $w=6.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.365 $Y=2.635
+ $X2=3.365 $Y2=2.72
r130 29 31 11.8673 $w=6.38e-07 $l=6.35e-07 $layer=LI1_cond $X=3.365 $Y=2.635
+ $X2=3.365 $Y2=2
r131 25 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2.72
r132 25 27 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2
r133 21 76 2.68304 $w=2.5e-07 $l=2.75e-07 $layer=LI1_cond $X=1.21 $Y=2.255
+ $X2=1.21 $Y2=2.53
r134 21 23 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=1.21 $Y=2.255
+ $X2=1.21 $Y2=1.66
r135 20 45 1.30481 $w=5.48e-07 $l=6e-08 $layer=LI1_cond $X=0.79 $Y=2.53 $X2=0.73
+ $Y2=2.53
r136 19 76 3.7769 $w=3.6e-07 $l=1.25e-07 $layer=LI1_cond $X=1.085 $Y=2.53
+ $X2=1.21 $Y2=2.53
r137 19 20 6.41533 $w=5.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.085 $Y=2.53
+ $X2=0.79 $Y2=2.53
r138 6 42 400 $w=1.7e-07 $l=9.60937e-07 $layer=licon1_PDIFF $count=1 $X=5.425
+ $Y=1.485 $X2=5.65 $Y2=2.34
r139 6 39 400 $w=1.7e-07 $l=3e-07 $layer=licon1_PDIFF $count=1 $X=5.425 $Y=1.485
+ $X2=5.65 $Y2=1.66
r140 5 35 300 $w=1.7e-07 $l=5.98268e-07 $layer=licon1_PDIFF $count=2 $X=4.395
+ $Y=1.485 $X2=4.575 $Y2=2
r141 4 31 150 $w=1.7e-07 $l=7.495e-07 $layer=licon1_PDIFF $count=4 $X=2.985
+ $Y=1.485 $X2=3.52 $Y2=2
r142 3 27 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=1.485 $X2=2.19 $Y2=2
r143 2 76 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.25 $Y2=2.34
r144 2 23 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.25 $Y2=1.66
r145 1 45 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.065 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_2%Y 1 2 3 4 5 18 20 24 26 30 32 36 39 41 42
+ 43 44 51
c92 51 0 1.55098e-19 $X=1.72 $Y=0.72
r93 43 44 6.69888 $w=5.48e-07 $l=2.55e-07 $layer=LI1_cond $X=1.695 $Y=1.19
+ $X2=1.695 $Y2=1.445
r94 42 43 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=1.695 $Y=0.85
+ $X2=1.695 $Y2=1.19
r95 42 51 3.94257 $w=3.78e-07 $l=1.3e-07 $layer=LI1_cond $X=1.695 $Y=0.85
+ $X2=1.695 $Y2=0.72
r96 34 36 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.075 $Y=1.665
+ $X2=5.075 $Y2=2
r97 33 41 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=4.235 $Y=1.555
+ $X2=4.045 $Y2=1.555
r98 32 34 7.46666 $w=2.2e-07 $l=2.38747e-07 $layer=LI1_cond $X=4.885 $Y=1.555
+ $X2=5.075 $Y2=1.665
r99 32 33 34.0495 $w=2.18e-07 $l=6.5e-07 $layer=LI1_cond $X=4.885 $Y=1.555
+ $X2=4.235 $Y2=1.555
r100 28 41 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=4.045 $Y=1.665
+ $X2=4.045 $Y2=1.555
r101 28 30 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=4.045 $Y=1.665
+ $X2=4.045 $Y2=2.34
r102 27 39 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.825 $Y=1.555
+ $X2=2.635 $Y2=1.555
r103 26 41 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=3.855 $Y=1.555
+ $X2=4.045 $Y2=1.555
r104 26 27 53.9553 $w=2.18e-07 $l=1.03e-06 $layer=LI1_cond $X=3.855 $Y=1.555
+ $X2=2.825 $Y2=1.555
r105 22 39 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=2.635 $Y=1.665
+ $X2=2.635 $Y2=1.555
r106 22 24 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=2.635 $Y=1.665
+ $X2=2.635 $Y2=2.34
r107 21 44 3.36699 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.885 $Y=1.555
+ $X2=1.695 $Y2=1.555
r108 20 39 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.445 $Y=1.555
+ $X2=2.635 $Y2=1.555
r109 20 21 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=2.445 $Y=1.555
+ $X2=1.885 $Y2=1.555
r110 16 44 3.21057 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=1.555
r111 16 18 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=2.34
r112 5 36 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.955
+ $Y=1.485 $X2=5.1 $Y2=2
r113 4 41 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=1.66
r114 4 30 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=2.34
r115 3 39 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=1.485 $X2=2.66 $Y2=1.66
r116 3 24 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=1.485 $X2=2.66 $Y2=2.34
r117 2 44 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=1.485 $X2=1.72 $Y2=1.66
r118 2 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=1.485 $X2=1.72 $Y2=2.34
r119 1 51 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.235 $X2=1.72 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_2%VGND 1 2 9 12 13 14 16 29 30 34
r70 34 37 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0 $X2=0.705
+ $Y2=0.38
r71 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r72 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r73 27 30 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r74 26 27 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r75 24 27 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=4.83
+ $Y2=0
r76 24 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r77 23 26 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=4.83
+ $Y2=0
r78 23 24 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r79 21 34 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r80 21 23 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.15
+ $Y2=0
r81 16 34 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r82 16 18 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r83 14 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r84 14 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r85 12 26 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.065 $Y=0 $X2=4.83
+ $Y2=0
r86 12 13 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=0 $X2=5.15
+ $Y2=0
r87 11 29 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=5.235 $Y=0 $X2=5.75
+ $Y2=0
r88 11 13 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.235 $Y=0 $X2=5.15
+ $Y2=0
r89 7 13 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.15 $Y=0.085 $X2=5.15
+ $Y2=0
r90 7 9 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.15 $Y=0.085 $X2=5.15
+ $Y2=0.38
r91 2 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.015
+ $Y=0.235 $X2=5.15 $Y2=0.38
r92 1 37 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_2%A_225_47# 1 2 3 10 12 14 20 22
r40 20 22 36.494 $w=2.68e-07 $l=8.55e-07 $layer=LI1_cond $X=2.275 $Y=0.77
+ $X2=3.13 $Y2=0.77
r41 17 20 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.19 $Y=0.635
+ $X2=2.275 $Y2=0.77
r42 17 19 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=0.635
+ $X2=2.19 $Y2=0.55
r43 16 19 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=0.465
+ $X2=2.19 $Y2=0.55
r44 15 25 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.335 $Y=0.36
+ $X2=1.21 $Y2=0.36
r45 14 16 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.105 $Y=0.36
+ $X2=2.19 $Y2=0.465
r46 14 15 40.6667 $w=2.08e-07 $l=7.7e-07 $layer=LI1_cond $X=2.105 $Y=0.36
+ $X2=1.335 $Y2=0.36
r47 10 25 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.21 $Y=0.465
+ $X2=1.21 $Y2=0.36
r48 10 12 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=1.21 $Y=0.465
+ $X2=1.21 $Y2=0.72
r49 3 22 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=2.945
+ $Y=0.235 $X2=3.13 $Y2=0.72
r50 2 19 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=2.055
+ $Y=0.235 $X2=2.19 $Y2=0.55
r51 1 25 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.25 $Y2=0.38
r52 1 12 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.25 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_2%A_495_47# 1 2 11
c15 11 0 1.05021e-19 $X=4.12 $Y=0.38
r16 8 11 77.1082 $w=2.08e-07 $l=1.46e-06 $layer=LI1_cond $X=2.66 $Y=0.36
+ $X2=4.12 $Y2=0.36
r17 2 11 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.985
+ $Y=0.235 $X2=4.12 $Y2=0.38
r18 1 8 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=2.66 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_2%A_705_47# 1 2 3 10 16 18 22 25
r45 20 22 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=5.622 $Y=0.715
+ $X2=5.622 $Y2=0.38
r46 19 25 5.71385 $w=2.3e-07 $l=1.73205e-07 $layer=LI1_cond $X=4.805 $Y=0.81
+ $X2=4.655 $Y2=0.76
r47 18 20 7.51555 $w=1.9e-07 $l=2.09175e-07 $layer=LI1_cond $X=5.455 $Y=0.81
+ $X2=5.622 $Y2=0.715
r48 18 19 37.9426 $w=1.88e-07 $l=6.5e-07 $layer=LI1_cond $X=5.455 $Y=0.81
+ $X2=4.805 $Y2=0.81
r49 14 25 0.905018 $w=2.6e-07 $l=1.54677e-07 $layer=LI1_cond $X=4.635 $Y=0.615
+ $X2=4.655 $Y2=0.76
r50 14 16 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=4.635 $Y=0.615
+ $X2=4.635 $Y2=0.42
r51 10 25 5.71385 $w=2.3e-07 $l=1.54919e-07 $layer=LI1_cond $X=4.505 $Y=0.77
+ $X2=4.655 $Y2=0.76
r52 10 12 36.494 $w=2.68e-07 $l=8.55e-07 $layer=LI1_cond $X=4.505 $Y=0.77
+ $X2=3.65 $Y2=0.77
r53 3 22 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.485
+ $Y=0.235 $X2=5.62 $Y2=0.38
r54 2 25 182 $w=1.7e-07 $l=6.08379e-07 $layer=licon1_NDIFF $count=1 $X=4.455
+ $Y=0.235 $X2=4.635 $Y2=0.76
r55 2 16 182 $w=1.7e-07 $l=2.59856e-07 $layer=licon1_NDIFF $count=1 $X=4.455
+ $Y=0.235 $X2=4.635 $Y2=0.42
r56 1 12 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=3.525
+ $Y=0.235 $X2=3.65 $Y2=0.72
.ends

