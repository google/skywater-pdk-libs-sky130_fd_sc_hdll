* File: sky130_fd_sc_hdll__a21boi_2.pxi.spice
* Created: Wed Sep  2 08:16:52 2020
* 
x_PM_SKY130_FD_SC_HDLL__A21BOI_2%B1_N N_B1_N_c_74_n N_B1_N_c_75_n N_B1_N_M1007_g
+ N_B1_N_M1010_g N_B1_N_c_69_n N_B1_N_c_70_n N_B1_N_c_71_n B1_N N_B1_N_c_73_n
+ PM_SKY130_FD_SC_HDLL__A21BOI_2%B1_N
x_PM_SKY130_FD_SC_HDLL__A21BOI_2%A_61_47# N_A_61_47#_M1010_s N_A_61_47#_M1007_d
+ N_A_61_47#_c_113_n N_A_61_47#_M1003_g N_A_61_47#_c_104_n N_A_61_47#_M1006_g
+ N_A_61_47#_c_114_n N_A_61_47#_M1005_g N_A_61_47#_M1012_g N_A_61_47#_c_106_n
+ N_A_61_47#_c_107_n N_A_61_47#_c_108_n N_A_61_47#_c_109_n N_A_61_47#_c_110_n
+ N_A_61_47#_c_111_n N_A_61_47#_c_112_n PM_SKY130_FD_SC_HDLL__A21BOI_2%A_61_47#
x_PM_SKY130_FD_SC_HDLL__A21BOI_2%A2 N_A2_c_176_n N_A2_M1001_g N_A2_c_177_n
+ N_A2_M1009_g N_A2_c_178_n N_A2_M1013_g N_A2_c_179_n N_A2_M1002_g N_A2_c_180_n
+ N_A2_c_198_p N_A2_c_193_n N_A2_c_181_n A2 N_A2_c_182_n N_A2_c_217_p
+ PM_SKY130_FD_SC_HDLL__A21BOI_2%A2
x_PM_SKY130_FD_SC_HDLL__A21BOI_2%A1 N_A1_c_257_n N_A1_M1004_g N_A1_c_261_n
+ N_A1_M1000_g N_A1_c_258_n N_A1_M1011_g N_A1_c_262_n N_A1_M1008_g A1
+ N_A1_c_260_n A1 PM_SKY130_FD_SC_HDLL__A21BOI_2%A1
x_PM_SKY130_FD_SC_HDLL__A21BOI_2%VPWR N_VPWR_M1007_s N_VPWR_M1001_d
+ N_VPWR_M1008_s N_VPWR_c_305_n N_VPWR_c_306_n N_VPWR_c_307_n N_VPWR_c_308_n
+ N_VPWR_c_309_n N_VPWR_c_310_n N_VPWR_c_311_n VPWR N_VPWR_c_312_n
+ N_VPWR_c_304_n PM_SKY130_FD_SC_HDLL__A21BOI_2%VPWR
x_PM_SKY130_FD_SC_HDLL__A21BOI_2%A_228_297# N_A_228_297#_M1003_d
+ N_A_228_297#_M1005_d N_A_228_297#_M1000_d N_A_228_297#_M1002_s
+ N_A_228_297#_c_371_n N_A_228_297#_c_379_n N_A_228_297#_c_372_n
+ N_A_228_297#_c_381_n N_A_228_297#_c_382_n N_A_228_297#_c_392_n
+ N_A_228_297#_c_420_n N_A_228_297#_c_395_n N_A_228_297#_c_373_n
+ N_A_228_297#_c_374_n N_A_228_297#_c_399_n
+ PM_SKY130_FD_SC_HDLL__A21BOI_2%A_228_297#
x_PM_SKY130_FD_SC_HDLL__A21BOI_2%Y N_Y_M1006_s N_Y_M1004_s N_Y_M1003_s
+ N_Y_c_436_n N_Y_c_444_n N_Y_c_445_n N_Y_c_455_n Y N_Y_c_447_n
+ PM_SKY130_FD_SC_HDLL__A21BOI_2%Y
x_PM_SKY130_FD_SC_HDLL__A21BOI_2%VGND N_VGND_M1010_d N_VGND_M1012_d
+ N_VGND_M1013_d N_VGND_c_484_n N_VGND_c_485_n N_VGND_c_486_n N_VGND_c_487_n
+ N_VGND_c_488_n N_VGND_c_489_n VGND N_VGND_c_490_n N_VGND_c_491_n
+ N_VGND_c_492_n N_VGND_c_493_n PM_SKY130_FD_SC_HDLL__A21BOI_2%VGND
cc_1 VNB N_B1_N_c_69_n 0.019806f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.73
cc_2 VNB N_B1_N_c_70_n 0.0389355f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.88
cc_3 VNB N_B1_N_c_71_n 0.00809188f $X=-0.19 $Y=-0.24 $X2=0.387 $Y2=1.435
cc_4 VNB B1_N 0.0209655f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_5 VNB N_B1_N_c_73_n 0.0333977f $X=-0.19 $Y=-0.24 $X2=0.34 $Y2=0.93
cc_6 VNB N_A_61_47#_c_104_n 0.019148f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.73
cc_7 VNB N_A_61_47#_M1012_g 0.0186736f $X=-0.19 $Y=-0.24 $X2=0.34 $Y2=0.93
cc_8 VNB N_A_61_47#_c_106_n 0.0325873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_61_47#_c_107_n 0.032938f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_61_47#_c_108_n 0.00754218f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_61_47#_c_109_n 0.0082377f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_61_47#_c_110_n 4.363e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_61_47#_c_111_n 0.0165811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_61_47#_c_112_n 0.00279787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A2_c_176_n 0.0222553f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.435
cc_16 VNB N_A2_c_177_n 0.0168453f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=2.1
cc_17 VNB N_A2_c_178_n 0.0227688f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=0.445
cc_18 VNB N_A2_c_179_n 0.0315085f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.73
cc_19 VNB N_A2_c_180_n 8.72475e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_20 VNB N_A2_c_181_n 0.00312578f $X=-0.19 $Y=-0.24 $X2=0.34 $Y2=0.93
cc_21 VNB N_A2_c_182_n 0.00709264f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A1_c_257_n 0.0162246f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.435
cc_23 VNB N_A1_c_258_n 0.0173683f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=0.445
cc_24 VNB A1 0.00437149f $X=-0.19 $Y=-0.24 $X2=0.387 $Y2=1.435
cc_25 VNB N_A1_c_260_n 0.0381875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_304_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_Y_c_436_n 0.0013059f $X=-0.19 $Y=-0.24 $X2=0.387 $Y2=1.223
cc_28 VNB N_VGND_c_484_n 0.00660273f $X=-0.19 $Y=-0.24 $X2=0.387 $Y2=1.223
cc_29 VNB N_VGND_c_485_n 0.00561552f $X=-0.19 $Y=-0.24 $X2=0.387 $Y2=0.93
cc_30 VNB N_VGND_c_486_n 0.0173534f $X=-0.19 $Y=-0.24 $X2=0.34 $Y2=0.93
cc_31 VNB N_VGND_c_487_n 0.0279067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_488_n 0.0212289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_489_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_490_n 0.032381f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_491_n 0.0421381f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_492_n 0.00461634f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_493_n 0.247963f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VPB N_B1_N_c_74_n 0.019936f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.715
cc_39 VPB N_B1_N_c_75_n 0.0294891f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.815
cc_40 VPB N_B1_N_c_71_n 0.0190975f $X=-0.19 $Y=1.305 $X2=0.387 $Y2=1.435
cc_41 VPB B1_N 0.0222924f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_42 VPB N_A_61_47#_c_113_n 0.0195217f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=0.445
cc_43 VPB N_A_61_47#_c_114_n 0.0164008f $X=-0.19 $Y=1.305 $X2=0.387 $Y2=1.435
cc_44 VPB N_A_61_47#_c_106_n 0.0159576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_61_47#_c_107_n 0.0228611f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_61_47#_c_110_n 0.0155902f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A2_c_176_n 0.0247855f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.435
cc_48 VPB N_A2_c_179_n 0.0289514f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=0.73
cc_49 VPB N_A2_c_180_n 0.00337424f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_50 VPB N_A2_c_182_n 0.00784196f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A1_c_261_n 0.016507f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=2.1
cc_52 VPB N_A1_c_262_n 0.0161202f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=0.73
cc_53 VPB A1 2.42596e-19 $X=-0.19 $Y=1.305 $X2=0.387 $Y2=1.435
cc_54 VPB N_A1_c_260_n 0.0204622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_305_n 0.0115529f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=0.73
cc_56 VPB N_VPWR_c_306_n 0.0230729f $X=-0.19 $Y=1.305 $X2=0.387 $Y2=1.223
cc_57 VPB N_VPWR_c_307_n 0.00420232f $X=-0.19 $Y=1.305 $X2=0.387 $Y2=0.93
cc_58 VPB N_VPWR_c_308_n 0.0554921f $X=-0.19 $Y=1.305 $X2=0.272 $Y2=0.85
cc_59 VPB N_VPWR_c_309_n 0.00324214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_310_n 0.00547845f $X=-0.19 $Y=1.305 $X2=0.272 $Y2=0.93
cc_61 VPB N_VPWR_c_311_n 0.0161222f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_312_n 0.0218501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_304_n 0.0699824f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_228_297#_c_371_n 0.00537941f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_228_297#_c_372_n 0.00293587f $X=-0.19 $Y=1.305 $X2=0.34 $Y2=0.93
cc_66 VPB N_A_228_297#_c_373_n 0.0111305f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_228_297#_c_374_n 0.0133845f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_Y_c_436_n 0.00146972f $X=-0.19 $Y=1.305 $X2=0.387 $Y2=1.223
cc_69 N_B1_N_c_69_n N_A_61_47#_c_104_n 0.00801723f $X=0.49 $Y=0.73 $X2=0 $Y2=0
cc_70 N_B1_N_c_73_n N_A_61_47#_c_106_n 0.00699351f $X=0.34 $Y=0.93 $X2=0 $Y2=0
cc_71 N_B1_N_c_69_n N_A_61_47#_c_108_n 0.00969164f $X=0.49 $Y=0.73 $X2=0 $Y2=0
cc_72 N_B1_N_c_70_n N_A_61_47#_c_108_n 0.0119208f $X=0.49 $Y=0.88 $X2=0 $Y2=0
cc_73 B1_N N_A_61_47#_c_108_n 0.00907806f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_74 N_B1_N_c_69_n N_A_61_47#_c_109_n 0.00756969f $X=0.49 $Y=0.73 $X2=0 $Y2=0
cc_75 N_B1_N_c_70_n N_A_61_47#_c_109_n 0.0112161f $X=0.49 $Y=0.88 $X2=0 $Y2=0
cc_76 B1_N N_A_61_47#_c_109_n 0.0183558f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_77 N_B1_N_c_73_n N_A_61_47#_c_109_n 0.00410312f $X=0.34 $Y=0.93 $X2=0 $Y2=0
cc_78 N_B1_N_c_75_n N_A_61_47#_c_110_n 0.00325111f $X=0.5 $Y=1.815 $X2=0 $Y2=0
cc_79 N_B1_N_c_71_n N_A_61_47#_c_110_n 0.0129344f $X=0.387 $Y=1.435 $X2=0 $Y2=0
cc_80 B1_N N_A_61_47#_c_110_n 0.0320633f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_81 B1_N N_A_61_47#_c_112_n 0.0148889f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_82 N_B1_N_c_73_n N_A_61_47#_c_112_n 0.00283179f $X=0.34 $Y=0.93 $X2=0 $Y2=0
cc_83 N_B1_N_c_75_n N_VPWR_c_306_n 0.00930811f $X=0.5 $Y=1.815 $X2=0 $Y2=0
cc_84 N_B1_N_c_71_n N_VPWR_c_306_n 7.59231e-19 $X=0.387 $Y=1.435 $X2=0 $Y2=0
cc_85 B1_N N_VPWR_c_306_n 0.0177312f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_86 N_B1_N_c_75_n N_VPWR_c_308_n 0.00602273f $X=0.5 $Y=1.815 $X2=0 $Y2=0
cc_87 N_B1_N_c_75_n N_VPWR_c_304_n 0.00586437f $X=0.5 $Y=1.815 $X2=0 $Y2=0
cc_88 N_B1_N_c_75_n N_A_228_297#_c_372_n 0.00265527f $X=0.5 $Y=1.815 $X2=0 $Y2=0
cc_89 N_B1_N_c_69_n N_VGND_c_484_n 0.00706259f $X=0.49 $Y=0.73 $X2=0 $Y2=0
cc_90 N_B1_N_c_69_n N_VGND_c_490_n 0.0037867f $X=0.49 $Y=0.73 $X2=0 $Y2=0
cc_91 N_B1_N_c_70_n N_VGND_c_490_n 0.00220222f $X=0.49 $Y=0.88 $X2=0 $Y2=0
cc_92 N_B1_N_c_69_n N_VGND_c_493_n 0.00728882f $X=0.49 $Y=0.73 $X2=0 $Y2=0
cc_93 N_B1_N_c_70_n N_VGND_c_493_n 0.00244058f $X=0.49 $Y=0.88 $X2=0 $Y2=0
cc_94 B1_N N_VGND_c_493_n 0.00603494f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_95 N_A_61_47#_c_114_n N_A2_c_176_n 0.023682f $X=2.015 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_96 N_A_61_47#_M1012_g N_A2_c_176_n 0.0222633f $X=2.04 $Y=0.56 $X2=-0.19
+ $Y2=-0.24
cc_97 N_A_61_47#_c_107_n N_A2_c_176_n 0.00370749f $X=2.015 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_98 N_A_61_47#_M1012_g N_A2_c_177_n 0.0189598f $X=2.04 $Y=0.56 $X2=0 $Y2=0
cc_99 N_A_61_47#_c_114_n N_A2_c_180_n 7.72205e-19 $X=2.015 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A_61_47#_c_107_n N_A2_c_180_n 0.00151698f $X=2.015 $Y=1.202 $X2=0 $Y2=0
cc_101 N_A_61_47#_c_114_n N_A2_c_193_n 0.00182399f $X=2.015 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_61_47#_c_107_n N_A2_c_181_n 0.0016157f $X=2.015 $Y=1.202 $X2=0 $Y2=0
cc_103 N_A_61_47#_c_113_n N_VPWR_c_308_n 0.00429453f $X=1.545 $Y=1.41 $X2=0
+ $Y2=0
cc_104 N_A_61_47#_c_114_n N_VPWR_c_308_n 0.00429355f $X=2.015 $Y=1.41 $X2=0
+ $Y2=0
cc_105 N_A_61_47#_c_110_n N_VPWR_c_308_n 0.00537589f $X=0.74 $Y=2.1 $X2=0 $Y2=0
cc_106 N_A_61_47#_c_113_n N_VPWR_c_304_n 0.00734734f $X=1.545 $Y=1.41 $X2=0
+ $Y2=0
cc_107 N_A_61_47#_c_114_n N_VPWR_c_304_n 0.00609013f $X=2.015 $Y=1.41 $X2=0
+ $Y2=0
cc_108 N_A_61_47#_c_110_n N_VPWR_c_304_n 0.00608145f $X=0.74 $Y=2.1 $X2=0 $Y2=0
cc_109 N_A_61_47#_c_106_n N_A_228_297#_c_371_n 0.00481342f $X=1.445 $Y=1.16
+ $X2=0 $Y2=0
cc_110 N_A_61_47#_c_110_n N_A_228_297#_c_371_n 0.0256566f $X=0.74 $Y=2.1 $X2=0
+ $Y2=0
cc_111 N_A_61_47#_c_111_n N_A_228_297#_c_371_n 0.00853716f $X=1.19 $Y=1.16 $X2=0
+ $Y2=0
cc_112 N_A_61_47#_c_113_n N_A_228_297#_c_379_n 0.0113402f $X=1.545 $Y=1.41 $X2=0
+ $Y2=0
cc_113 N_A_61_47#_c_114_n N_A_228_297#_c_379_n 0.0115699f $X=2.015 $Y=1.41 $X2=0
+ $Y2=0
cc_114 N_A_61_47#_c_114_n N_A_228_297#_c_381_n 0.00592015f $X=2.015 $Y=1.41
+ $X2=0 $Y2=0
cc_115 N_A_61_47#_c_113_n N_A_228_297#_c_382_n 7.90282e-19 $X=1.545 $Y=1.41
+ $X2=0 $Y2=0
cc_116 N_A_61_47#_c_114_n N_A_228_297#_c_382_n 0.00506665f $X=2.015 $Y=1.41
+ $X2=0 $Y2=0
cc_117 N_A_61_47#_c_113_n N_Y_c_436_n 0.0272528f $X=1.545 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A_61_47#_c_104_n N_Y_c_436_n 0.00839378f $X=1.57 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A_61_47#_c_114_n N_Y_c_436_n 0.00723354f $X=2.015 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_61_47#_M1012_g N_Y_c_436_n 0.00558221f $X=2.04 $Y=0.56 $X2=0 $Y2=0
cc_121 N_A_61_47#_c_107_n N_Y_c_436_n 0.0383087f $X=2.015 $Y=1.202 $X2=0 $Y2=0
cc_122 N_A_61_47#_c_111_n N_Y_c_436_n 0.0170986f $X=1.19 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A_61_47#_M1012_g N_Y_c_444_n 0.0147337f $X=2.04 $Y=0.56 $X2=0 $Y2=0
cc_124 N_A_61_47#_c_104_n N_Y_c_445_n 0.0030072f $X=1.57 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_61_47#_c_107_n N_Y_c_445_n 2.05567e-19 $X=2.015 $Y=1.202 $X2=0 $Y2=0
cc_126 N_A_61_47#_c_104_n N_Y_c_447_n 0.00734847f $X=1.57 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_61_47#_c_104_n N_VGND_c_484_n 0.00931367f $X=1.57 $Y=0.995 $X2=0
+ $Y2=0
cc_128 N_A_61_47#_c_106_n N_VGND_c_484_n 0.00602899f $X=1.445 $Y=1.16 $X2=0
+ $Y2=0
cc_129 N_A_61_47#_c_109_n N_VGND_c_484_n 0.0163983f $X=0.735 $Y=1.07 $X2=0 $Y2=0
cc_130 N_A_61_47#_c_111_n N_VGND_c_484_n 0.0178755f $X=1.19 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_61_47#_M1012_g N_VGND_c_485_n 0.00318876f $X=2.04 $Y=0.56 $X2=0 $Y2=0
cc_132 N_A_61_47#_c_104_n N_VGND_c_488_n 0.00404729f $X=1.57 $Y=0.995 $X2=0
+ $Y2=0
cc_133 N_A_61_47#_M1012_g N_VGND_c_488_n 0.00422112f $X=2.04 $Y=0.56 $X2=0 $Y2=0
cc_134 N_A_61_47#_c_108_n N_VGND_c_490_n 0.0203667f $X=0.645 $Y=0.445 $X2=0
+ $Y2=0
cc_135 N_A_61_47#_M1010_s N_VGND_c_493_n 0.00299073f $X=0.305 $Y=0.235 $X2=0
+ $Y2=0
cc_136 N_A_61_47#_c_104_n N_VGND_c_493_n 0.00728096f $X=1.57 $Y=0.995 $X2=0
+ $Y2=0
cc_137 N_A_61_47#_M1012_g N_VGND_c_493_n 0.00595896f $X=2.04 $Y=0.56 $X2=0 $Y2=0
cc_138 N_A_61_47#_c_108_n N_VGND_c_493_n 0.0190389f $X=0.645 $Y=0.445 $X2=0
+ $Y2=0
cc_139 N_A2_c_177_n N_A1_c_257_n 0.0388034f $X=2.57 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_140 N_A2_c_176_n N_A1_c_261_n 0.0396504f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A2_c_180_n N_A1_c_261_n 0.00200016f $X=2.487 $Y=1.495 $X2=0 $Y2=0
cc_142 N_A2_c_198_p N_A1_c_261_n 0.0124289f $X=3.735 $Y=1.585 $X2=0 $Y2=0
cc_143 N_A2_c_178_n N_A1_c_258_n 0.0332704f $X=3.89 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A2_c_179_n N_A1_c_262_n 0.0375814f $X=3.915 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A2_c_198_p N_A1_c_262_n 0.0124894f $X=3.735 $Y=1.585 $X2=0 $Y2=0
cc_146 N_A2_c_182_n N_A1_c_262_n 0.00193514f $X=3.95 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A2_c_176_n A1 8.51484e-19 $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A2_c_179_n A1 3.56938e-19 $X=3.915 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A2_c_198_p A1 0.045762f $X=3.735 $Y=1.585 $X2=0 $Y2=0
cc_150 N_A2_c_181_n A1 0.0202426f $X=2.46 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A2_c_182_n A1 0.0277378f $X=3.95 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A2_c_176_n N_A1_c_260_n 0.0425075f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A2_c_179_n N_A1_c_260_n 0.0208702f $X=3.915 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A2_c_180_n N_A1_c_260_n 0.00206091f $X=2.487 $Y=1.495 $X2=0 $Y2=0
cc_155 N_A2_c_198_p N_A1_c_260_n 0.00658914f $X=3.735 $Y=1.585 $X2=0 $Y2=0
cc_156 N_A2_c_181_n N_A1_c_260_n 8.45859e-19 $X=2.46 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A2_c_182_n N_A1_c_260_n 0.00309543f $X=3.95 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A2_c_198_p N_VPWR_M1001_d 0.006471f $X=3.735 $Y=1.585 $X2=0 $Y2=0
cc_159 N_A2_c_193_n N_VPWR_M1001_d 4.30199e-19 $X=2.675 $Y=1.585 $X2=0 $Y2=0
cc_160 N_A2_c_198_p N_VPWR_M1008_s 0.00750181f $X=3.735 $Y=1.585 $X2=0 $Y2=0
cc_161 N_A2_c_217_p N_VPWR_M1008_s 3.63664e-19 $X=3.91 $Y=1.495 $X2=0 $Y2=0
cc_162 N_A2_c_176_n N_VPWR_c_307_n 0.0039542f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A2_c_176_n N_VPWR_c_308_n 0.0051032f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A2_c_179_n N_VPWR_c_310_n 0.0078402f $X=3.915 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A2_c_179_n N_VPWR_c_312_n 0.00464324f $X=3.915 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A2_c_176_n N_VPWR_c_304_n 0.00678224f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A2_c_179_n N_VPWR_c_304_n 0.00627369f $X=3.915 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A2_c_193_n N_A_228_297#_M1005_d 0.00277296f $X=2.675 $Y=1.585 $X2=0
+ $Y2=0
cc_169 N_A2_c_198_p N_A_228_297#_M1000_d 0.00358863f $X=3.735 $Y=1.585 $X2=0
+ $Y2=0
cc_170 N_A2_c_182_n N_A_228_297#_M1002_s 3.74695e-19 $X=3.95 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A2_c_217_p N_A_228_297#_M1002_s 0.00836932f $X=3.91 $Y=1.495 $X2=0
+ $Y2=0
cc_172 N_A2_c_176_n N_A_228_297#_c_379_n 0.00227366f $X=2.485 $Y=1.41 $X2=0
+ $Y2=0
cc_173 N_A2_c_176_n N_A_228_297#_c_381_n 7.36455e-19 $X=2.485 $Y=1.41 $X2=0
+ $Y2=0
cc_174 N_A2_c_193_n N_A_228_297#_c_381_n 0.00473113f $X=2.675 $Y=1.585 $X2=0
+ $Y2=0
cc_175 N_A2_c_176_n N_A_228_297#_c_382_n 0.00423695f $X=2.485 $Y=1.41 $X2=0
+ $Y2=0
cc_176 N_A2_c_176_n N_A_228_297#_c_392_n 0.010823f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A2_c_198_p N_A_228_297#_c_392_n 0.0214606f $X=3.735 $Y=1.585 $X2=0
+ $Y2=0
cc_178 N_A2_c_193_n N_A_228_297#_c_392_n 0.0147606f $X=2.675 $Y=1.585 $X2=0
+ $Y2=0
cc_179 N_A2_c_179_n N_A_228_297#_c_395_n 0.0136586f $X=3.915 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A2_c_198_p N_A_228_297#_c_395_n 0.0235438f $X=3.735 $Y=1.585 $X2=0
+ $Y2=0
cc_181 N_A2_c_217_p N_A_228_297#_c_395_n 0.0160146f $X=3.91 $Y=1.495 $X2=0 $Y2=0
cc_182 N_A2_c_217_p N_A_228_297#_c_373_n 0.00192735f $X=3.91 $Y=1.495 $X2=0
+ $Y2=0
cc_183 N_A2_c_198_p N_A_228_297#_c_399_n 0.0131878f $X=3.735 $Y=1.585 $X2=0
+ $Y2=0
cc_184 N_A2_c_176_n N_Y_c_436_n 4.54742e-19 $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A2_c_180_n N_Y_c_436_n 0.0106235f $X=2.487 $Y=1.495 $X2=0 $Y2=0
cc_186 N_A2_c_193_n N_Y_c_436_n 0.00764665f $X=2.675 $Y=1.585 $X2=0 $Y2=0
cc_187 N_A2_c_181_n N_Y_c_436_n 0.00681678f $X=2.46 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A2_c_176_n N_Y_c_444_n 0.00405236f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A2_c_177_n N_Y_c_444_n 0.0124372f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A2_c_181_n N_Y_c_444_n 0.0172611f $X=2.46 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A2_c_177_n N_Y_c_455_n 0.00145841f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A2_c_178_n N_Y_c_455_n 0.00163897f $X=3.89 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A2_c_177_n N_VGND_c_485_n 0.00318876f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A2_c_178_n N_VGND_c_487_n 0.00479247f $X=3.89 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A2_c_179_n N_VGND_c_487_n 6.09842e-19 $X=3.915 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A2_c_182_n N_VGND_c_487_n 0.00570392f $X=3.95 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A2_c_177_n N_VGND_c_491_n 0.00422112f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A2_c_178_n N_VGND_c_491_n 0.00585385f $X=3.89 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A2_c_177_n N_VGND_c_493_n 0.00574008f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A2_c_178_n N_VGND_c_493_n 0.0118428f $X=3.89 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A1_c_261_n N_VPWR_c_307_n 0.00285238f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A1_c_261_n N_VPWR_c_310_n 5.56307e-19 $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A1_c_262_n N_VPWR_c_310_n 0.00913948f $X=3.435 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A1_c_261_n N_VPWR_c_311_n 0.0052046f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A1_c_262_n N_VPWR_c_311_n 0.0032362f $X=3.435 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A1_c_261_n N_VPWR_c_304_n 0.00687867f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A1_c_262_n N_VPWR_c_304_n 0.00384231f $X=3.435 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A1_c_261_n N_A_228_297#_c_382_n 7.49249e-19 $X=2.955 $Y=1.41 $X2=0
+ $Y2=0
cc_209 N_A1_c_261_n N_A_228_297#_c_392_n 0.0117763f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A1_c_262_n N_A_228_297#_c_395_n 0.0132365f $X=3.435 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A1_c_257_n N_Y_c_444_n 0.00916468f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_212 A1 N_Y_c_444_n 0.00753835f $X=3.23 $Y=1.105 $X2=0 $Y2=0
cc_213 N_A1_c_257_n N_Y_c_455_n 0.00761699f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A1_c_258_n N_Y_c_455_n 0.0107845f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_215 A1 N_Y_c_455_n 0.0215803f $X=3.23 $Y=1.105 $X2=0 $Y2=0
cc_216 N_A1_c_260_n N_Y_c_455_n 0.00338805f $X=3.41 $Y=1.202 $X2=0 $Y2=0
cc_217 N_A1_c_257_n N_VGND_c_491_n 0.0041289f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A1_c_258_n N_VGND_c_491_n 0.0054895f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A1_c_257_n N_VGND_c_493_n 0.00570321f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A1_c_258_n N_VGND_c_493_n 0.0102103f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_221 N_VPWR_c_304_n N_A_228_297#_M1003_d 0.00254418f $X=4.37 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_222 N_VPWR_c_304_n N_A_228_297#_M1005_d 0.00231261f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_223 N_VPWR_c_304_n N_A_228_297#_M1000_d 0.00288166f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_224 N_VPWR_c_304_n N_A_228_297#_M1002_s 0.00255363f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_225 N_VPWR_c_306_n N_A_228_297#_c_371_n 5.25358e-19 $X=0.26 $Y=2.165 $X2=0
+ $Y2=0
cc_226 N_VPWR_c_307_n N_A_228_297#_c_379_n 0.0115829f $X=2.72 $Y=2.36 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_308_n N_A_228_297#_c_379_n 0.0604576f $X=2.635 $Y=2.72 $X2=0
+ $Y2=0
cc_228 N_VPWR_c_304_n N_A_228_297#_c_379_n 0.0381843f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_229 N_VPWR_c_306_n N_A_228_297#_c_372_n 0.00542158f $X=0.26 $Y=2.165 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_308_n N_A_228_297#_c_372_n 0.017616f $X=2.635 $Y=2.72 $X2=0
+ $Y2=0
cc_231 N_VPWR_c_304_n N_A_228_297#_c_372_n 0.00962421f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_232 N_VPWR_c_307_n N_A_228_297#_c_382_n 0.00547755f $X=2.72 $Y=2.36 $X2=0
+ $Y2=0
cc_233 N_VPWR_M1001_d N_A_228_297#_c_392_n 0.00362947f $X=2.575 $Y=1.485 $X2=0
+ $Y2=0
cc_234 N_VPWR_c_307_n N_A_228_297#_c_392_n 0.0130459f $X=2.72 $Y=2.36 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_308_n N_A_228_297#_c_392_n 0.0027955f $X=2.635 $Y=2.72 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_311_n N_A_228_297#_c_392_n 0.00367471f $X=3.46 $Y=2.72 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_304_n N_A_228_297#_c_392_n 0.0131151f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_307_n N_A_228_297#_c_420_n 0.0127516f $X=2.72 $Y=2.36 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_310_n N_A_228_297#_c_420_n 0.0135709f $X=3.675 $Y=2.36 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_311_n N_A_228_297#_c_420_n 0.0117203f $X=3.46 $Y=2.72 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_304_n N_A_228_297#_c_420_n 0.00645162f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_242 N_VPWR_M1008_s N_A_228_297#_c_395_n 0.00395992f $X=3.525 $Y=1.485 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_310_n N_A_228_297#_c_395_n 0.0200578f $X=3.675 $Y=2.36 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_311_n N_A_228_297#_c_395_n 0.00274283f $X=3.46 $Y=2.72 $X2=0
+ $Y2=0
cc_245 N_VPWR_c_312_n N_A_228_297#_c_395_n 0.00345885f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_304_n N_A_228_297#_c_395_n 0.0119994f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_247 N_VPWR_c_312_n N_A_228_297#_c_374_n 0.0179903f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_248 N_VPWR_c_304_n N_A_228_297#_c_374_n 0.00990273f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_249 N_VPWR_c_304_n N_Y_M1003_s 0.00232895f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_250 N_A_228_297#_c_379_n N_Y_M1003_s 0.00344991f $X=2.035 $Y=2.375 $X2=0
+ $Y2=0
cc_251 N_A_228_297#_c_371_n N_Y_c_436_n 0.0238336f $X=1.265 $Y=1.96 $X2=0 $Y2=0
cc_252 N_A_228_297#_c_379_n N_Y_c_436_n 0.0209745f $X=2.035 $Y=2.375 $X2=0 $Y2=0
cc_253 N_A_228_297#_c_381_n N_Y_c_436_n 0.0140391f $X=2.225 $Y=2.025 $X2=0 $Y2=0
cc_254 N_A_228_297#_c_382_n N_Y_c_436_n 0.00703767f $X=2.225 $Y=2.285 $X2=0
+ $Y2=0
cc_255 N_Y_c_444_n N_VGND_M1012_d 0.009211f $X=2.98 $Y=0.7 $X2=0 $Y2=0
cc_256 N_Y_c_436_n N_VGND_c_484_n 0.00666656f $X=1.78 $Y=1.61 $X2=0 $Y2=0
cc_257 N_Y_c_445_n N_VGND_c_484_n 0.0120674f $X=1.78 $Y=0.76 $X2=0 $Y2=0
cc_258 N_Y_c_447_n N_VGND_c_484_n 0.0241122f $X=1.78 $Y=0.42 $X2=0 $Y2=0
cc_259 N_Y_c_444_n N_VGND_c_485_n 0.020165f $X=2.98 $Y=0.7 $X2=0 $Y2=0
cc_260 N_Y_c_444_n N_VGND_c_488_n 0.00408888f $X=2.98 $Y=0.7 $X2=0 $Y2=0
cc_261 N_Y_c_447_n N_VGND_c_488_n 0.0218467f $X=1.78 $Y=0.42 $X2=0 $Y2=0
cc_262 N_Y_c_444_n N_VGND_c_491_n 0.00789715f $X=2.98 $Y=0.7 $X2=0 $Y2=0
cc_263 N_Y_c_455_n N_VGND_c_491_n 0.0221123f $X=3.195 $Y=0.36 $X2=0 $Y2=0
cc_264 N_Y_M1006_s N_VGND_c_493_n 0.00286149f $X=1.645 $Y=0.235 $X2=0 $Y2=0
cc_265 N_Y_M1004_s N_VGND_c_493_n 0.0026338f $X=3.005 $Y=0.235 $X2=0 $Y2=0
cc_266 N_Y_c_444_n N_VGND_c_493_n 0.0216805f $X=2.98 $Y=0.7 $X2=0 $Y2=0
cc_267 N_Y_c_455_n N_VGND_c_493_n 0.0141007f $X=3.195 $Y=0.36 $X2=0 $Y2=0
cc_268 N_Y_c_447_n N_VGND_c_493_n 0.0125929f $X=1.78 $Y=0.42 $X2=0 $Y2=0
cc_269 N_Y_c_444_n A_529_47# 0.00529826f $X=2.98 $Y=0.7 $X2=-0.19 $Y2=-0.24
cc_270 N_VGND_c_493_n A_529_47# 0.00239227f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
cc_271 N_VGND_c_493_n A_697_47# 0.014106f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
