* File: sky130_fd_sc_hdll__nor4bb_1.pex.spice
* Created: Thu Aug 27 19:17:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_1%C_N 2 3 5 8 9 10 14 15 16
r34 14 17 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.16
+ $X2=0.53 $Y2=1.325
r35 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.16
+ $X2=0.53 $Y2=0.995
r36 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.16 $X2=0.53 $Y2=1.16
r37 9 10 9.79577 $w=3.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.63 $Y=1.19 $X2=0.63
+ $Y2=1.53
r38 9 15 0.864332 $w=3.98e-07 $l=3e-08 $layer=LI1_cond $X=0.63 $Y=1.19 $X2=0.63
+ $Y2=1.16
r39 8 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.56 $Y=0.675
+ $X2=0.56 $Y2=0.995
r40 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.975
+ $X2=0.495 $Y2=2.26
r41 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.875 $X2=0.495
+ $Y2=1.975
r42 2 17 182.367 $w=2e-07 $l=5.5e-07 $layer=POLY_cond $X=0.495 $Y=1.875
+ $X2=0.495 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_1%D_N 1 3 4 6 7 14
r30 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.085
+ $Y=1.16 $X2=1.085 $Y2=1.16
r31 7 14 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.255 $Y=1.16
+ $X2=1.085 $Y2=1.16
r32 4 10 49.9093 $w=2.71e-07 $l=2.7157e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.075 $Y2=1.16
r33 4 6 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.03 $Y=1.41 $X2=1.03
+ $Y2=1.695
r34 1 10 38.8824 $w=2.71e-07 $l=1.96914e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.075 $Y2=1.16
r35 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_1%A_216_93# 1 2 7 9 10 12 13 14 15 19 24 27
r60 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.705
+ $Y=1.16 $X2=1.705 $Y2=1.16
r61 22 24 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=1.525
+ $X2=1.705 $Y2=1.16
r62 21 24 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.705 $Y=0.825
+ $X2=1.705 $Y2=1.16
r63 20 27 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.345 $Y=0.74
+ $X2=1.26 $Y2=0.66
r64 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.62 $Y=0.74
+ $X2=1.705 $Y2=0.825
r65 19 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.62 $Y=0.74
+ $X2=1.345 $Y2=0.74
r66 15 22 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.62 $Y=1.62
+ $X2=1.705 $Y2=1.525
r67 15 17 20.7225 $w=1.88e-07 $l=3.55e-07 $layer=LI1_cond $X=1.62 $Y=1.62
+ $X2=1.265 $Y2=1.62
r68 13 25 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.92 $Y=1.16
+ $X2=1.705 $Y2=1.16
r69 13 14 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.92 $Y=1.16
+ $X2=2.02 $Y2=1.202
r70 10 14 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=2.045 $Y=0.995
+ $X2=2.02 $Y2=1.202
r71 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.045 $Y=0.995
+ $X2=2.045 $Y2=0.56
r72 7 14 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=2.02 $Y=1.41
+ $X2=2.02 $Y2=1.202
r73 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.02 $Y=1.41 $X2=2.02
+ $Y2=1.985
r74 2 17 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.485 $X2=1.265 $Y2=1.63
r75 1 27 182 $w=1.7e-07 $l=2.70416e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.465 $X2=1.26 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_1%A_27_410# 1 2 7 9 10 12 14 17 19 22 23 24
+ 27 33 35
r77 30 33 3.93367 $w=3.73e-07 $l=1.28e-07 $layer=LI1_cond $X=0.172 $Y=0.637
+ $X2=0.3 $Y2=0.637
r78 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.465
+ $Y=1.16 $X2=2.465 $Y2=1.16
r79 25 27 55.6605 $w=2.33e-07 $l=1.135e-06 $layer=LI1_cond $X=2.497 $Y=2.295
+ $X2=2.497 $Y2=1.16
r80 23 25 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=2.38 $Y=2.38
+ $X2=2.497 $Y2=2.295
r81 23 24 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=2.38 $Y=2.38
+ $X2=1.305 $Y2=2.38
r82 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.22 $Y=2.295
+ $X2=1.305 $Y2=2.38
r83 21 22 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.22 $Y=2.07
+ $X2=1.22 $Y2=2.295
r84 20 35 1.93133 $w=1.85e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.977
+ $X2=0.215 $Y2=1.977
r85 19 21 6.83233 $w=1.85e-07 $l=1.28662e-07 $layer=LI1_cond $X=1.135 $Y=1.977
+ $X2=1.22 $Y2=2.07
r86 19 20 47.3612 $w=1.83e-07 $l=7.9e-07 $layer=LI1_cond $X=1.135 $Y=1.977
+ $X2=0.345 $Y2=1.977
r87 15 35 4.5059 $w=2.17e-07 $l=9.3e-08 $layer=LI1_cond $X=0.215 $Y=2.07
+ $X2=0.215 $Y2=1.977
r88 15 17 9.75144 $w=2.58e-07 $l=2.2e-07 $layer=LI1_cond $X=0.215 $Y=2.07
+ $X2=0.215 $Y2=2.29
r89 14 35 4.5059 $w=2.17e-07 $l=1.11445e-07 $layer=LI1_cond $X=0.172 $Y=1.885
+ $X2=0.215 $Y2=1.977
r90 13 30 5.2298 $w=1.75e-07 $l=1.88e-07 $layer=LI1_cond $X=0.172 $Y=0.825
+ $X2=0.172 $Y2=0.637
r91 13 14 67.1792 $w=1.73e-07 $l=1.06e-06 $layer=LI1_cond $X=0.172 $Y=0.825
+ $X2=0.172 $Y2=1.885
r92 10 28 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.525 $Y=0.995
+ $X2=2.465 $Y2=1.16
r93 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.525 $Y=0.995
+ $X2=2.525 $Y2=0.56
r94 7 28 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.5 $Y=1.41
+ $X2=2.465 $Y2=1.16
r95 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.5 $Y=1.41 $X2=2.5
+ $Y2=1.985
r96 2 17 600 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.05 $X2=0.26 $Y2=2.29
r97 1 33 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.465 $X2=0.3 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_1%B 1 3 4 6 7 11
r28 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.985
+ $Y=1.16 $X2=2.985 $Y2=1.16
r29 7 11 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.975 $Y=1.53
+ $X2=2.975 $Y2=1.16
r30 4 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.045 $Y=0.995
+ $X2=2.985 $Y2=1.16
r31 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.045 $Y=0.995
+ $X2=3.045 $Y2=0.56
r32 1 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.02 $Y=1.41
+ $X2=2.985 $Y2=1.16
r33 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.02 $Y=1.41 $X2=3.02
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_1%A 1 3 4 6 7
r20 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.525
+ $Y=1.16 $X2=3.525 $Y2=1.16
r21 4 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.49 $Y=1.41
+ $X2=3.525 $Y2=1.16
r22 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.49 $Y=1.41 $X2=3.49
+ $Y2=1.985
r23 1 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.465 $Y=0.995
+ $X2=3.525 $Y2=1.16
r24 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.465 $Y=0.995
+ $X2=3.465 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_1%VPWR 1 2 9 11 13 15 17 22 31 35
r45 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r46 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r47 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r48 28 29 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r49 26 29 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r50 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r51 25 28 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r52 25 26 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r53 23 31 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r54 23 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r55 22 34 6.00926 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=3.51 $Y=2.72
+ $X2=3.825 $Y2=2.72
r56 22 28 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.51 $Y=2.72 $X2=3.45
+ $Y2=2.72
r57 17 31 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r58 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r59 15 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r60 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r61 11 34 3.05232 $w=4.8e-07 $l=1.16619e-07 $layer=LI1_cond $X=3.75 $Y=2.635
+ $X2=3.825 $Y2=2.72
r62 11 13 15.8231 $w=4.78e-07 $l=6.35e-07 $layer=LI1_cond $X=3.75 $Y=2.635
+ $X2=3.75 $Y2=2
r63 7 31 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r64 7 9 9.40151 $w=3.78e-07 $l=3.1e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.325
r65 2 13 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.58
+ $Y=1.485 $X2=3.725 $Y2=2
r66 1 9 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.05 $X2=0.73 $Y2=2.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_1%Y 1 2 3 10 15 18 20 22 24
r48 23 24 8.87273 $w=1.98e-07 $l=1.6e-07 $layer=LI1_cond $X=3.24 $Y=0.655
+ $X2=3.24 $Y2=0.495
r49 21 22 2.36881 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.37 $Y=0.74
+ $X2=2.165 $Y2=0.74
r50 20 23 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.14 $Y=0.74
+ $X2=3.24 $Y2=0.655
r51 20 21 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.14 $Y=0.74
+ $X2=2.37 $Y2=0.74
r52 16 22 4.06715 $w=2.25e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.27 $Y=0.655
+ $X2=2.165 $Y2=0.74
r53 16 18 8.87273 $w=1.98e-07 $l=1.6e-07 $layer=LI1_cond $X=2.27 $Y=0.655
+ $X2=2.27 $Y2=0.495
r54 14 22 4.06715 $w=2.25e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.085 $Y=0.825
+ $X2=2.165 $Y2=0.74
r55 14 15 52.0904 $w=2.48e-07 $l=1.13e-06 $layer=LI1_cond $X=2.085 $Y=0.825
+ $X2=2.085 $Y2=1.955
r56 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.96 $Y=2.04
+ $X2=2.085 $Y2=1.955
r57 10 12 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.96 $Y=2.04
+ $X2=1.785 $Y2=2.04
r58 3 12 600 $w=1.7e-07 $l=6.14329e-07 $layer=licon1_PDIFF $count=1 $X=1.66
+ $Y=1.485 $X2=1.785 $Y2=2.04
r59 2 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=3.12
+ $Y=0.235 $X2=3.255 $Y2=0.495
r60 1 18 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=2.12
+ $Y=0.235 $X2=2.255 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_1%VGND 1 2 3 4 15 19 23 25 27 30 31 33 34
+ 36 37 38 50 56 58
r64 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r65 53 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r66 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r67 50 55 6.00926 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=3.51 $Y=0 $X2=3.825
+ $Y2=0
r68 50 52 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.51 $Y=0 $X2=3.45
+ $Y2=0
r69 49 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r70 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r71 46 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r72 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r73 42 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r74 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r75 38 42 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r76 38 58 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r77 36 48 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.59 $Y=0 $X2=2.53
+ $Y2=0
r78 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=0 $X2=2.755
+ $Y2=0
r79 35 52 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.92 $Y=0 $X2=3.45
+ $Y2=0
r80 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.92 $Y=0 $X2=2.755
+ $Y2=0
r81 33 45 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.62 $Y=0 $X2=1.61
+ $Y2=0
r82 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.62 $Y=0 $X2=1.785
+ $Y2=0
r83 32 48 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=1.95 $Y=0 $X2=2.53
+ $Y2=0
r84 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.95 $Y=0 $X2=1.785
+ $Y2=0
r85 30 41 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.705 $Y=0 $X2=0.69
+ $Y2=0
r86 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0 $X2=0.79
+ $Y2=0
r87 29 45 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.61
+ $Y2=0
r88 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.79
+ $Y2=0
r89 25 55 3.05232 $w=4.8e-07 $l=1.16619e-07 $layer=LI1_cond $X=3.75 $Y=0.085
+ $X2=3.825 $Y2=0
r90 25 27 7.60008 $w=4.78e-07 $l=3.05e-07 $layer=LI1_cond $X=3.75 $Y=0.085
+ $X2=3.75 $Y2=0.39
r91 21 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=0.085
+ $X2=2.755 $Y2=0
r92 21 23 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.755 $Y=0.085
+ $X2=2.755 $Y2=0.39
r93 17 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=0.085
+ $X2=1.785 $Y2=0
r94 17 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.785 $Y=0.085
+ $X2=1.785 $Y2=0.38
r95 13 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r96 13 15 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.66
r97 4 27 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.54
+ $Y=0.235 $X2=3.725 $Y2=0.39
r98 3 23 182 $w=1.7e-07 $l=2.19203e-07 $layer=licon1_NDIFF $count=1 $X=2.6
+ $Y=0.235 $X2=2.755 $Y2=0.39
r99 2 19 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.66
+ $Y=0.235 $X2=1.785 $Y2=0.38
r100 1 15 182 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_NDIFF $count=1 $X=0.635
+ $Y=0.465 $X2=0.79 $Y2=0.66
.ends

