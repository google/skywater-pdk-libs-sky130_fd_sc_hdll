# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__and3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.745000 0.410000 1.325000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.915000 2.125000 2.490000 2.465000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.305000 2.370000 0.765000 ;
        RECT 1.985000 0.765000 2.620000 1.245000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.125000 1.795000 3.590000 2.465000 ;
        RECT 3.165000 0.255000 3.570000 0.715000 ;
        RECT 3.240000 0.715000 3.570000 0.925000 ;
        RECT 3.240000 0.925000 4.040000 1.445000 ;
        RECT 3.240000 1.445000 3.590000 1.795000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.085000 0.355000 0.575000 ;
      RECT 0.085000  1.575000 0.400000 2.635000 ;
      RECT 0.630000  0.305000 0.905000 1.015000 ;
      RECT 0.630000  1.015000 1.465000 1.245000 ;
      RECT 0.630000  1.245000 0.905000 1.905000 ;
      RECT 1.080000  2.130000 1.745000 2.635000 ;
      RECT 1.100000  1.425000 3.020000 1.595000 ;
      RECT 1.100000  1.595000 1.335000 1.960000 ;
      RECT 1.105000  0.305000 1.815000 0.570000 ;
      RECT 1.505000  1.765000 1.885000 1.955000 ;
      RECT 1.505000  1.955000 1.745000 2.130000 ;
      RECT 1.645000  0.570000 1.815000 1.425000 ;
      RECT 2.160000  1.595000 2.350000 1.890000 ;
      RECT 2.610000  0.085000 2.940000 0.580000 ;
      RECT 2.660000  1.790000 2.875000 2.635000 ;
      RECT 2.790000  0.995000 3.020000 1.425000 ;
      RECT 3.760000  0.085000 4.025000 0.745000 ;
      RECT 3.760000  1.625000 4.025000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and3b_2
END LIBRARY
