* File: sky130_fd_sc_hdll__o21bai_4.pex.spice
* Created: Wed Sep  2 08:44:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O21BAI_4%B1_N 1 3 4 6 7 15
c26 15 0 1.46056e-19 $X=0.375 $Y=1.19
c27 1 0 1.30421e-19 $X=0.545 $Y=1.41
r28 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.345
+ $Y=1.16 $X2=0.345 $Y2=1.16
r29 7 15 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=0.23 $Y=1.18
+ $X2=0.345 $Y2=1.18
r30 4 10 39.3227 $w=3.86e-07 $l=2.25433e-07 $layer=POLY_cond $X=0.57 $Y=0.995
+ $X2=0.427 $Y2=1.16
r31 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.57 $Y=0.995 $X2=0.57
+ $Y2=0.56
r32 1 10 45.0491 $w=3.86e-07 $l=3.03315e-07 $layer=POLY_cond $X=0.545 $Y=1.41
+ $X2=0.427 $Y2=1.16
r33 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.545 $Y=1.41
+ $X2=0.545 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_4%A_33_297# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 31 33 35 39 42 44 50 55 56 65
c98 65 0 1.46056e-19 $X=2.55 $Y=1.202
c99 28 0 1.76278e-19 $X=3.02 $Y=0.995
r100 65 66 62.7535 $w=3.61e-07 $l=4.7e-07 $layer=POLY_cond $X=2.55 $Y=1.202
+ $X2=3.02 $Y2=1.202
r101 64 65 16.6898 $w=3.61e-07 $l=1.25e-07 $layer=POLY_cond $X=2.425 $Y=1.202
+ $X2=2.55 $Y2=1.202
r102 61 62 16.6898 $w=3.61e-07 $l=1.25e-07 $layer=POLY_cond $X=1.955 $Y=1.202
+ $X2=2.08 $Y2=1.202
r103 60 61 46.0637 $w=3.61e-07 $l=3.45e-07 $layer=POLY_cond $X=1.61 $Y=1.202
+ $X2=1.955 $Y2=1.202
r104 59 60 16.6898 $w=3.61e-07 $l=1.25e-07 $layer=POLY_cond $X=1.485 $Y=1.202
+ $X2=1.61 $Y2=1.202
r105 51 64 23.3657 $w=3.61e-07 $l=1.75e-07 $layer=POLY_cond $X=2.25 $Y=1.202
+ $X2=2.425 $Y2=1.202
r106 51 62 22.6981 $w=3.61e-07 $l=1.7e-07 $layer=POLY_cond $X=2.25 $Y=1.202
+ $X2=2.08 $Y2=1.202
r107 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.25
+ $Y=1.16 $X2=2.25 $Y2=1.16
r108 48 59 54.0748 $w=3.61e-07 $l=4.05e-07 $layer=POLY_cond $X=1.08 $Y=1.202
+ $X2=1.485 $Y2=1.202
r109 48 57 8.67867 $w=3.61e-07 $l=6.5e-08 $layer=POLY_cond $X=1.08 $Y=1.202
+ $X2=1.015 $Y2=1.202
r110 47 50 61.7922 $w=2.08e-07 $l=1.17e-06 $layer=LI1_cond $X=1.08 $Y=1.18
+ $X2=2.25 $Y2=1.18
r111 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.08
+ $Y=1.16 $X2=1.08 $Y2=1.16
r112 45 56 1.46923 $w=2.1e-07 $l=1.33e-07 $layer=LI1_cond $X=0.945 $Y=1.18
+ $X2=0.812 $Y2=1.18
r113 45 47 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=0.945 $Y=1.18
+ $X2=1.08 $Y2=1.18
r114 43 56 5.01685 $w=2.17e-07 $l=1.26333e-07 $layer=LI1_cond $X=0.765 $Y=1.285
+ $X2=0.812 $Y2=1.18
r115 43 44 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.765 $Y=1.285
+ $X2=0.765 $Y2=1.455
r116 42 56 5.01685 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=0.812 $Y=1.075
+ $X2=0.812 $Y2=1.18
r117 42 55 7.82791 $w=2.63e-07 $l=1.8e-07 $layer=LI1_cond $X=0.812 $Y=1.075
+ $X2=0.812 $Y2=0.895
r118 37 55 6.82995 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=0.755 $Y=0.705
+ $X2=0.755 $Y2=0.895
r119 37 39 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.755 $Y=0.705
+ $X2=0.755 $Y2=0.39
r120 36 54 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.475 $Y=1.54
+ $X2=0.31 $Y2=1.54
r121 35 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.68 $Y=1.54
+ $X2=0.765 $Y2=1.455
r122 35 36 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.68 $Y=1.54
+ $X2=0.475 $Y2=1.54
r123 31 54 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.31 $Y=1.625
+ $X2=0.31 $Y2=1.54
r124 31 33 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.31 $Y=1.625
+ $X2=0.31 $Y2=2.3
r125 28 66 23.3725 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.02 $Y=0.995
+ $X2=3.02 $Y2=1.202
r126 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.02 $Y=0.995
+ $X2=3.02 $Y2=0.56
r127 25 65 23.3725 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.55 $Y=0.995
+ $X2=2.55 $Y2=1.202
r128 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.55 $Y=0.995
+ $X2=2.55 $Y2=0.56
r129 22 64 19.0337 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.202
r130 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.985
r131 19 62 23.3725 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.08 $Y=0.995
+ $X2=2.08 $Y2=1.202
r132 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.08 $Y=0.995
+ $X2=2.08 $Y2=0.56
r133 16 61 19.0337 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.202
r134 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.985
r135 13 60 23.3725 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.61 $Y=0.995
+ $X2=1.61 $Y2=1.202
r136 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.61 $Y=0.995
+ $X2=1.61 $Y2=0.56
r137 10 59 19.0337 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.202
r138 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.985
r139 7 57 19.0337 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.015 $Y=1.41
+ $X2=1.015 $Y2=1.202
r140 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.015 $Y=1.41
+ $X2=1.015 $Y2=1.985
r141 2 54 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.485 $X2=0.31 $Y2=1.62
r142 2 33 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.485 $X2=0.31 $Y2=2.3
r143 1 39 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.645
+ $Y=0.235 $X2=0.78 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_4%A2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39 44
r86 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.875 $Y=1.202
+ $X2=4.9 $Y2=1.202
r87 37 39 22.6747 $w=3.72e-07 $l=1.75e-07 $layer=POLY_cond $X=4.7 $Y=1.202
+ $X2=4.875 $Y2=1.202
r88 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.7 $Y=1.16
+ $X2=4.7 $Y2=1.16
r89 35 37 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=4.405 $Y=1.202
+ $X2=4.7 $Y2=1.202
r90 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.38 $Y=1.202
+ $X2=4.405 $Y2=1.202
r91 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=3.935 $Y=1.202
+ $X2=4.38 $Y2=1.202
r92 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.91 $Y=1.202
+ $X2=3.935 $Y2=1.202
r93 31 44 21.0727 $w=1.98e-07 $l=3.8e-07 $layer=LI1_cond $X=3.53 $Y=1.175
+ $X2=3.91 $Y2=1.175
r94 30 32 49.2366 $w=3.72e-07 $l=3.8e-07 $layer=POLY_cond $X=3.53 $Y=1.202
+ $X2=3.91 $Y2=1.202
r95 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.53
+ $Y=1.16 $X2=3.53 $Y2=1.16
r96 28 30 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=3.465 $Y=1.202
+ $X2=3.53 $Y2=1.202
r97 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.44 $Y=1.202
+ $X2=3.465 $Y2=1.202
r98 25 38 21.6273 $w=1.98e-07 $l=3.9e-07 $layer=LI1_cond $X=4.31 $Y=1.175
+ $X2=4.7 $Y2=1.175
r99 25 44 22.1818 $w=1.98e-07 $l=4e-07 $layer=LI1_cond $X=4.31 $Y=1.175 $X2=3.91
+ $Y2=1.175
r100 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.9 $Y=0.995
+ $X2=4.9 $Y2=1.202
r101 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.9 $Y=0.995
+ $X2=4.9 $Y2=0.56
r102 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.875 $Y=1.41
+ $X2=4.875 $Y2=1.202
r103 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.875 $Y=1.41
+ $X2=4.875 $Y2=1.985
r104 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.405 $Y=1.41
+ $X2=4.405 $Y2=1.202
r105 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.405 $Y=1.41
+ $X2=4.405 $Y2=1.985
r106 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.38 $Y=0.995
+ $X2=4.38 $Y2=1.202
r107 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.38 $Y=0.995
+ $X2=4.38 $Y2=0.56
r108 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.935 $Y=1.41
+ $X2=3.935 $Y2=1.202
r109 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.935 $Y=1.41
+ $X2=3.935 $Y2=1.985
r110 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.91 $Y=0.995
+ $X2=3.91 $Y2=1.202
r111 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.91 $Y=0.995
+ $X2=3.91 $Y2=0.56
r112 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.465 $Y=1.41
+ $X2=3.465 $Y2=1.202
r113 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.465 $Y=1.41
+ $X2=3.465 $Y2=1.985
r114 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.44 $Y=0.995
+ $X2=3.44 $Y2=1.202
r115 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.44 $Y=0.995
+ $X2=3.44 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_4%A1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 41 44
r75 41 42 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.755 $Y=1.202
+ $X2=6.78 $Y2=1.202
r76 39 41 26.5618 $w=3.72e-07 $l=2.05e-07 $layer=POLY_cond $X=6.55 $Y=1.202
+ $X2=6.755 $Y2=1.202
r77 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.55
+ $Y=1.16 $X2=6.55 $Y2=1.16
r78 37 39 34.336 $w=3.72e-07 $l=2.65e-07 $layer=POLY_cond $X=6.285 $Y=1.202
+ $X2=6.55 $Y2=1.202
r79 36 37 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.26 $Y=1.202
+ $X2=6.285 $Y2=1.202
r80 35 36 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=5.815 $Y=1.202
+ $X2=6.26 $Y2=1.202
r81 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.79 $Y=1.202
+ $X2=5.815 $Y2=1.202
r82 33 44 4.75325 $w=2.08e-07 $l=9e-08 $layer=LI1_cond $X=5.38 $Y=1.18 $X2=5.29
+ $Y2=1.18
r83 32 34 53.1237 $w=3.72e-07 $l=4.1e-07 $layer=POLY_cond $X=5.38 $Y=1.202
+ $X2=5.79 $Y2=1.202
r84 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.38
+ $Y=1.16 $X2=5.38 $Y2=1.16
r85 30 32 4.53495 $w=3.72e-07 $l=3.5e-08 $layer=POLY_cond $X=5.345 $Y=1.202
+ $X2=5.38 $Y2=1.202
r86 29 30 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.32 $Y=1.202
+ $X2=5.345 $Y2=1.202
r87 26 40 16.3723 $w=2.08e-07 $l=3.1e-07 $layer=LI1_cond $X=6.86 $Y=1.18
+ $X2=6.55 $Y2=1.18
r88 25 40 37.4978 $w=2.08e-07 $l=7.1e-07 $layer=LI1_cond $X=5.84 $Y=1.18
+ $X2=6.55 $Y2=1.18
r89 25 33 24.2944 $w=2.08e-07 $l=4.6e-07 $layer=LI1_cond $X=5.84 $Y=1.18
+ $X2=5.38 $Y2=1.18
r90 22 42 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.78 $Y=0.995
+ $X2=6.78 $Y2=1.202
r91 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.78 $Y=0.995
+ $X2=6.78 $Y2=0.56
r92 19 41 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.755 $Y=1.41
+ $X2=6.755 $Y2=1.202
r93 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.755 $Y=1.41
+ $X2=6.755 $Y2=1.985
r94 16 37 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.285 $Y=1.41
+ $X2=6.285 $Y2=1.202
r95 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.285 $Y=1.41
+ $X2=6.285 $Y2=1.985
r96 13 36 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.26 $Y=0.995
+ $X2=6.26 $Y2=1.202
r97 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.26 $Y=0.995
+ $X2=6.26 $Y2=0.56
r98 10 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.815 $Y=1.41
+ $X2=5.815 $Y2=1.202
r99 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.815 $Y=1.41
+ $X2=5.815 $Y2=1.985
r100 7 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.79 $Y=0.995
+ $X2=5.79 $Y2=1.202
r101 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.79 $Y=0.995
+ $X2=5.79 $Y2=0.56
r102 4 30 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.345 $Y=1.41
+ $X2=5.345 $Y2=1.202
r103 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.345 $Y=1.41
+ $X2=5.345 $Y2=1.985
r104 1 29 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.32 $Y=0.995
+ $X2=5.32 $Y2=1.202
r105 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.32 $Y=0.995
+ $X2=5.32 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_4%VPWR 1 2 3 4 5 18 20 24 28 32 36 38 39 41
+ 42 44 45 47 48 49 69 70 73
r100 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r101 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r102 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r103 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r104 64 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r105 63 64 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r106 61 64 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=5.29 $Y2=2.72
r107 60 63 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=5.29 $Y2=2.72
r108 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r109 58 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r110 58 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r111 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r112 55 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.845 $Y=2.72
+ $X2=1.72 $Y2=2.72
r113 55 57 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.845 $Y=2.72
+ $X2=2.53 $Y2=2.72
r114 53 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r115 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r116 49 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r117 47 66 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.395 $Y=2.72
+ $X2=6.21 $Y2=2.72
r118 47 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.395 $Y=2.72
+ $X2=6.52 $Y2=2.72
r119 46 69 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=6.645 $Y=2.72
+ $X2=7.13 $Y2=2.72
r120 46 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.645 $Y=2.72
+ $X2=6.52 $Y2=2.72
r121 44 63 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.455 $Y=2.72
+ $X2=5.29 $Y2=2.72
r122 44 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.455 $Y=2.72
+ $X2=5.58 $Y2=2.72
r123 43 66 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=5.705 $Y=2.72
+ $X2=6.21 $Y2=2.72
r124 43 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.705 $Y=2.72
+ $X2=5.58 $Y2=2.72
r125 41 57 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.535 $Y=2.72
+ $X2=2.53 $Y2=2.72
r126 41 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.535 $Y=2.72
+ $X2=2.66 $Y2=2.72
r127 40 60 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.785 $Y=2.72
+ $X2=2.99 $Y2=2.72
r128 40 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.785 $Y=2.72
+ $X2=2.66 $Y2=2.72
r129 38 52 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.695 $Y=2.72
+ $X2=0.69 $Y2=2.72
r130 38 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=2.72
+ $X2=0.78 $Y2=2.72
r131 34 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=2.635
+ $X2=6.52 $Y2=2.72
r132 34 36 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=6.52 $Y=2.635
+ $X2=6.52 $Y2=1.96
r133 30 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.58 $Y=2.635
+ $X2=5.58 $Y2=2.72
r134 30 32 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.58 $Y=2.635
+ $X2=5.58 $Y2=1.96
r135 26 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=2.635
+ $X2=2.66 $Y2=2.72
r136 26 28 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.66 $Y=2.635
+ $X2=2.66 $Y2=1.96
r137 22 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=2.635
+ $X2=1.72 $Y2=2.72
r138 22 24 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.72 $Y=2.635
+ $X2=1.72 $Y2=1.96
r139 21 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.865 $Y=2.72
+ $X2=0.78 $Y2=2.72
r140 20 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.595 $Y=2.72
+ $X2=1.72 $Y2=2.72
r141 20 21 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.595 $Y=2.72
+ $X2=0.865 $Y2=2.72
r142 16 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=2.635
+ $X2=0.78 $Y2=2.72
r143 16 18 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.78 $Y=2.635
+ $X2=0.78 $Y2=1.96
r144 5 36 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.375
+ $Y=1.485 $X2=6.52 $Y2=1.96
r145 4 32 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.435
+ $Y=1.485 $X2=5.58 $Y2=1.96
r146 3 28 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.515
+ $Y=1.485 $X2=2.66 $Y2=1.96
r147 2 24 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.575
+ $Y=1.485 $X2=1.72 $Y2=1.96
r148 1 18 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.635
+ $Y=1.485 $X2=0.78 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_4%Y 1 2 3 4 5 6 19 21 23 25 31 33 35 39 47
+ 51 53 54 61
c88 19 0 1.30421e-19 $X=1.205 $Y=1.625
r89 62 63 0.119608 $w=4.98e-07 $l=5e-09 $layer=LI1_cond $X=2.945 $Y=1.535
+ $X2=2.945 $Y2=1.54
r90 54 63 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=2.695 $Y=1.54
+ $X2=2.945 $Y2=1.54
r91 54 62 0.119608 $w=4.98e-07 $l=5e-09 $layer=LI1_cond $X=2.945 $Y=1.53
+ $X2=2.945 $Y2=1.535
r92 54 61 14.4049 $w=4.98e-07 $l=4.55e-07 $layer=LI1_cond $X=2.945 $Y=1.53
+ $X2=2.945 $Y2=1.075
r93 45 54 14.6641 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=2.315 $Y=1.54
+ $X2=2.695 $Y2=1.54
r94 45 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.315 $Y=1.54
+ $X2=2.19 $Y2=1.54
r95 40 51 6.72674 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.825 $Y=1.535
+ $X2=3.7 $Y2=1.535
r96 39 53 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.515 $Y=1.535
+ $X2=4.64 $Y2=1.535
r97 39 40 42.5152 $w=1.78e-07 $l=6.9e-07 $layer=LI1_cond $X=4.515 $Y=1.535
+ $X2=3.825 $Y2=1.535
r98 36 62 6.79934 $w=1.8e-07 $l=2.5e-07 $layer=LI1_cond $X=3.195 $Y=1.535
+ $X2=2.945 $Y2=1.535
r99 35 51 6.72674 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.575 $Y=1.535
+ $X2=3.7 $Y2=1.535
r100 35 36 23.4141 $w=1.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.575 $Y=1.535
+ $X2=3.195 $Y2=1.535
r101 33 49 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=0.815
+ $X2=2.81 $Y2=0.73
r102 33 61 13.0276 $w=2.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.81 $Y=0.815
+ $X2=2.81 $Y2=1.075
r103 29 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=1.625
+ $X2=2.19 $Y2=1.54
r104 29 31 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.19 $Y=1.625
+ $X2=2.19 $Y2=2.3
r105 25 49 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.695 $Y=0.73
+ $X2=2.81 $Y2=0.73
r106 25 27 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.695 $Y=0.73
+ $X2=1.82 $Y2=0.73
r107 24 44 5.2341 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.375 $Y=1.54
+ $X2=1.205 $Y2=1.54
r108 23 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.065 $Y=1.54
+ $X2=2.19 $Y2=1.54
r109 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.065 $Y=1.54
+ $X2=1.375 $Y2=1.54
r110 19 44 2.61705 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=1.625
+ $X2=1.205 $Y2=1.54
r111 19 21 22.8794 $w=3.38e-07 $l=6.75e-07 $layer=LI1_cond $X=1.205 $Y=1.625
+ $X2=1.205 $Y2=2.3
r112 6 53 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=4.495
+ $Y=1.485 $X2=4.64 $Y2=1.62
r113 5 51 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.555
+ $Y=1.485 $X2=3.7 $Y2=1.62
r114 4 47 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.485 $X2=2.19 $Y2=1.62
r115 4 31 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.485 $X2=2.19 $Y2=2.3
r116 3 44 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.105
+ $Y=1.485 $X2=1.25 $Y2=1.62
r117 3 21 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.105
+ $Y=1.485 $X2=1.25 $Y2=2.3
r118 2 49 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.625
+ $Y=0.235 $X2=2.76 $Y2=0.73
r119 1 27 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.685
+ $Y=0.235 $X2=1.82 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_4%A_621_297# 1 2 3 4 5 18 20 21 24 26 28 29
+ 30 34 36 38 40 42 48
r65 38 50 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.99 $Y=1.625
+ $X2=6.99 $Y2=1.54
r66 38 40 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=6.99 $Y=1.625
+ $X2=6.99 $Y2=2.3
r67 37 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.175 $Y=1.54
+ $X2=6.05 $Y2=1.54
r68 36 50 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.865 $Y=1.54
+ $X2=6.99 $Y2=1.54
r69 36 37 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.865 $Y=1.54
+ $X2=6.175 $Y2=1.54
r70 32 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.05 $Y=1.625
+ $X2=6.05 $Y2=1.54
r71 32 34 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=6.05 $Y=1.625
+ $X2=6.05 $Y2=2.3
r72 31 44 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.235 $Y=1.54
+ $X2=5.11 $Y2=1.54
r73 30 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.925 $Y=1.54
+ $X2=6.05 $Y2=1.54
r74 30 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.925 $Y=1.54
+ $X2=5.235 $Y2=1.54
r75 29 46 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.11 $Y=2.295
+ $X2=5.11 $Y2=2.38
r76 28 44 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.11 $Y=1.625
+ $X2=5.11 $Y2=1.54
r77 28 29 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=5.11 $Y=1.625
+ $X2=5.11 $Y2=2.295
r78 27 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.295 $Y=2.38
+ $X2=4.17 $Y2=2.38
r79 26 46 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.985 $Y=2.38
+ $X2=5.11 $Y2=2.38
r80 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.985 $Y=2.38
+ $X2=4.295 $Y2=2.38
r81 22 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.17 $Y=2.295
+ $X2=4.17 $Y2=2.38
r82 22 24 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.17 $Y=2.295
+ $X2=4.17 $Y2=1.96
r83 20 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.045 $Y=2.38
+ $X2=4.17 $Y2=2.38
r84 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.045 $Y=2.38
+ $X2=3.355 $Y2=2.38
r85 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.19 $Y=2.295
+ $X2=3.355 $Y2=2.38
r86 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.19 $Y=2.295
+ $X2=3.19 $Y2=1.96
r87 5 50 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.845
+ $Y=1.485 $X2=6.99 $Y2=1.62
r88 5 40 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=6.845
+ $Y=1.485 $X2=6.99 $Y2=2.3
r89 4 48 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.905
+ $Y=1.485 $X2=6.05 $Y2=1.62
r90 4 34 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.905
+ $Y=1.485 $X2=6.05 $Y2=2.3
r91 3 46 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=1.485 $X2=5.11 $Y2=2.3
r92 3 44 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=1.485 $X2=5.11 $Y2=1.62
r93 2 24 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.025
+ $Y=1.485 $X2=4.17 $Y2=1.96
r94 1 18 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=3.105
+ $Y=1.485 $X2=3.23 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_4%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 40
+ 41 43 44 46 47 48 67 68
r105 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r106 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r107 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r108 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r109 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r110 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r111 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r112 56 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r113 55 56 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r114 53 56 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=3.45 $Y2=0
r115 52 55 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=3.45
+ $Y2=0
r116 52 53 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r117 50 71 3.40825 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.197 $Y2=0
r118 50 52 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.69
+ $Y2=0
r119 48 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r120 48 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r121 46 64 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.435 $Y=0
+ $X2=6.21 $Y2=0
r122 46 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=0 $X2=6.52
+ $Y2=0
r123 45 67 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=6.605 $Y=0
+ $X2=7.13 $Y2=0
r124 45 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.605 $Y=0 $X2=6.52
+ $Y2=0
r125 43 61 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.495 $Y=0
+ $X2=5.29 $Y2=0
r126 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.495 $Y=0 $X2=5.58
+ $Y2=0
r127 42 64 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=5.665 $Y=0
+ $X2=6.21 $Y2=0
r128 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.665 $Y=0 $X2=5.58
+ $Y2=0
r129 40 58 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.555 $Y=0
+ $X2=4.37 $Y2=0
r130 40 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.555 $Y=0 $X2=4.64
+ $Y2=0
r131 39 61 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=4.725 $Y=0 $X2=5.29
+ $Y2=0
r132 39 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.725 $Y=0 $X2=4.64
+ $Y2=0
r133 37 55 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=0
+ $X2=3.45 $Y2=0
r134 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=0 $X2=3.7
+ $Y2=0
r135 36 58 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.785 $Y=0
+ $X2=4.37 $Y2=0
r136 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.785 $Y=0 $X2=3.7
+ $Y2=0
r137 32 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=0.085
+ $X2=6.52 $Y2=0
r138 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.52 $Y=0.085
+ $X2=6.52 $Y2=0.39
r139 28 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.58 $Y=0.085
+ $X2=5.58 $Y2=0
r140 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.58 $Y=0.085
+ $X2=5.58 $Y2=0.39
r141 24 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0
r142 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0.39
r143 20 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.085 $X2=3.7
+ $Y2=0
r144 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0.39
r145 16 71 3.40825 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=0.31 $Y=0.085
+ $X2=0.197 $Y2=0
r146 16 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.31 $Y=0.085
+ $X2=0.31 $Y2=0.39
r147 5 34 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=6.335
+ $Y=0.235 $X2=6.52 $Y2=0.39
r148 4 30 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=5.395
+ $Y=0.235 $X2=5.58 $Y2=0.39
r149 3 26 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.455
+ $Y=0.235 $X2=4.64 $Y2=0.39
r150 2 22 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=3.515
+ $Y=0.235 $X2=3.7 $Y2=0.39
r151 1 18 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.235 $X2=0.31 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_4%A_245_47# 1 2 3 4 5 6 7 22 28 29 30 34 36
+ 40 42 46 48 52 58 59 60
c119 29 0 1.76278e-19 $X=3.27 $Y=0.725
r120 50 52 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.965 $Y=0.725
+ $X2=6.965 $Y2=0.39
r121 49 60 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.215 $Y=0.815
+ $X2=6.025 $Y2=0.815
r122 48 50 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=6.775 $Y=0.815
+ $X2=6.965 $Y2=0.725
r123 48 49 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=6.775 $Y=0.815
+ $X2=6.215 $Y2=0.815
r124 44 60 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=6.025 $Y=0.725
+ $X2=6.025 $Y2=0.815
r125 44 46 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.025 $Y=0.725
+ $X2=6.025 $Y2=0.39
r126 43 59 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.275 $Y=0.815
+ $X2=5.085 $Y2=0.815
r127 42 60 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.835 $Y=0.815
+ $X2=6.025 $Y2=0.815
r128 42 43 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=5.835 $Y=0.815
+ $X2=5.275 $Y2=0.815
r129 38 59 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=5.085 $Y=0.725
+ $X2=5.085 $Y2=0.815
r130 38 40 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.085 $Y=0.725
+ $X2=5.085 $Y2=0.39
r131 37 58 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.335 $Y=0.815
+ $X2=4.145 $Y2=0.815
r132 36 59 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.895 $Y=0.815
+ $X2=5.085 $Y2=0.815
r133 36 37 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.895 $Y=0.815
+ $X2=4.335 $Y2=0.815
r134 32 58 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=4.145 $Y=0.725
+ $X2=4.145 $Y2=0.815
r135 32 34 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.145 $Y=0.725
+ $X2=4.145 $Y2=0.39
r136 31 57 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.395 $Y=0.815
+ $X2=3.27 $Y2=0.815
r137 30 58 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.955 $Y=0.815
+ $X2=4.145 $Y2=0.815
r138 30 31 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.955 $Y=0.815
+ $X2=3.395 $Y2=0.815
r139 29 57 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=3.27 $Y=0.725 $X2=3.27
+ $Y2=0.815
r140 28 55 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=0.475
+ $X2=3.27 $Y2=0.39
r141 28 29 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=3.27 $Y=0.475
+ $X2=3.27 $Y2=0.725
r142 24 27 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.35 $Y=0.39
+ $X2=2.29 $Y2=0.39
r143 22 55 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.145 $Y=0.39
+ $X2=3.27 $Y2=0.39
r144 22 27 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=3.145 $Y=0.39
+ $X2=2.29 $Y2=0.39
r145 7 52 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.855
+ $Y=0.235 $X2=6.99 $Y2=0.39
r146 6 46 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=5.865
+ $Y=0.235 $X2=6.05 $Y2=0.39
r147 5 40 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.975
+ $Y=0.235 $X2=5.11 $Y2=0.39
r148 4 34 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.985
+ $Y=0.235 $X2=4.17 $Y2=0.39
r149 3 57 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.095
+ $Y=0.235 $X2=3.23 $Y2=0.73
r150 3 55 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.095
+ $Y=0.235 $X2=3.23 $Y2=0.39
r151 2 27 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.155
+ $Y=0.235 $X2=2.29 $Y2=0.39
r152 1 24 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.225
+ $Y=0.235 $X2=1.35 $Y2=0.39
.ends

