* File: sky130_fd_sc_hdll__clkbuf_6.pex.spice
* Created: Wed Sep  2 08:25:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_6%A 1 3 6 10 12 14 15 16 24
r41 24 25 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.202
+ $X2=0.965 $Y2=1.202
r42 23 24 55.463 $w=3.65e-07 $l=4.2e-07 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.94 $Y2=1.202
r43 22 23 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r44 20 22 29.7123 $w=3.65e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.202
+ $X2=0.495 $Y2=1.202
r45 16 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r46 15 16 11.5244 $w=3.08e-07 $l=3.1e-07 $layer=LI1_cond $X=0.24 $Y=0.85
+ $X2=0.24 $Y2=1.16
r47 12 25 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r48 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r49 8 24 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=1.202
r50 8 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=0.445
r51 4 23 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r52 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r53 1 22 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r54 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_6%A_117_297# 1 2 7 9 12 16 18 20 21 23 26
+ 30 32 34 35 37 40 44 46 48 51 55 64 67 80
r139 80 81 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=3.76 $Y=1.202
+ $X2=3.785 $Y2=1.202
r140 79 80 54.7135 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.34 $Y=1.202
+ $X2=3.76 $Y2=1.202
r141 78 79 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=3.315 $Y=1.202
+ $X2=3.34 $Y2=1.202
r142 75 76 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.845 $Y2=1.202
r143 74 75 55.3649 $w=3.7e-07 $l=4.25e-07 $layer=POLY_cond $X=2.395 $Y=1.202
+ $X2=2.82 $Y2=1.202
r144 73 74 2.60541 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.395 $Y2=1.202
r145 72 73 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=2.375 $Y2=1.202
r146 71 72 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.88 $Y=1.202
+ $X2=1.905 $Y2=1.202
r147 68 69 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.46 $Y2=1.202
r148 65 78 11.7243 $w=3.7e-07 $l=9e-08 $layer=POLY_cond $X=3.225 $Y=1.202
+ $X2=3.315 $Y2=1.202
r149 65 76 49.5027 $w=3.7e-07 $l=3.8e-07 $layer=POLY_cond $X=3.225 $Y=1.202
+ $X2=2.845 $Y2=1.202
r150 64 65 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3.225
+ $Y=1.16 $X2=3.225 $Y2=1.16
r151 62 71 46.2459 $w=3.7e-07 $l=3.55e-07 $layer=POLY_cond $X=1.525 $Y=1.202
+ $X2=1.88 $Y2=1.202
r152 62 69 8.46757 $w=3.7e-07 $l=6.5e-08 $layer=POLY_cond $X=1.525 $Y=1.202
+ $X2=1.46 $Y2=1.202
r153 61 64 78.3661 $w=2.48e-07 $l=1.7e-06 $layer=LI1_cond $X=1.525 $Y=1.2
+ $X2=3.225 $Y2=1.2
r154 61 62 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=1.525
+ $Y=1.16 $X2=1.525 $Y2=1.16
r155 59 67 2.3589 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.2
+ $X2=0.73 $Y2=1.2
r156 59 61 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=0.895 $Y=1.2
+ $X2=1.525 $Y2=1.2
r157 55 57 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.73 $Y=1.66
+ $X2=0.73 $Y2=2.34
r158 53 67 4.07664 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.73 $Y=1.325
+ $X2=0.73 $Y2=1.2
r159 53 55 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.73 $Y=1.325
+ $X2=0.73 $Y2=1.66
r160 49 67 4.07664 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.73 $Y=1.075
+ $X2=0.73 $Y2=1.2
r161 49 51 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=0.73 $Y=1.075
+ $X2=0.73 $Y2=0.445
r162 46 81 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.202
r163 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r164 42 80 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.76 $Y=0.995
+ $X2=3.76 $Y2=1.202
r165 42 44 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.76 $Y=0.995
+ $X2=3.76 $Y2=0.445
r166 38 79 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.34 $Y=0.995
+ $X2=3.34 $Y2=1.202
r167 38 40 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.34 $Y=0.995
+ $X2=3.34 $Y2=0.445
r168 35 78 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.202
r169 35 37 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r170 32 76 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r171 32 34 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r172 28 75 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=1.202
r173 28 30 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=0.445
r174 24 74 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.395 $Y=0.995
+ $X2=2.395 $Y2=1.202
r175 24 26 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.395 $Y=0.995
+ $X2=2.395 $Y2=0.445
r176 21 73 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r177 21 23 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r178 18 72 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r179 18 20 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r180 14 71 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.88 $Y=0.995
+ $X2=1.88 $Y2=1.202
r181 14 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.88 $Y=0.995
+ $X2=1.88 $Y2=0.445
r182 10 69 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=1.202
r183 10 12 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=0.445
r184 7 68 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r185 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r186 2 57 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r187 2 55 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r188 1 51 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_6%VPWR 1 2 3 4 5 16 18 24 28 32 34 38 40 44
+ 46 48 55 56 62 65 68 71
r63 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r64 69 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r65 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r66 66 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r67 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r68 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r69 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r70 56 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r71 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r72 53 71 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.155 $Y=2.72
+ $X2=4.02 $Y2=2.72
r73 53 55 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.155 $Y=2.72
+ $X2=4.37 $Y2=2.72
r74 52 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r75 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r76 49 59 4.49698 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r77 49 51 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.69 $Y2=2.72
r78 48 62 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=1.2 $Y2=2.72
r79 48 51 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=0.69 $Y2=2.72
r80 46 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r81 46 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r82 42 71 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=2.72
r83 42 44 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=2
r84 41 68 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=3.08 $Y2=2.72
r85 40 71 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=4.02 $Y2=2.72
r86 40 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=3.215 $Y2=2.72
r87 36 68 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2.72
r88 36 38 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2
r89 35 65 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.14 $Y2=2.72
r90 34 68 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=3.08 $Y2=2.72
r91 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=2.275 $Y2=2.72
r92 30 65 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.72
r93 30 32 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2
r94 29 62 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.2 $Y2=2.72
r95 28 65 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=2.14 $Y2=2.72
r96 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=1.335 $Y2=2.72
r97 24 27 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.2 $Y=1.66 $X2=1.2
+ $Y2=2.34
r98 22 62 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.72
r99 22 27 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.34
r100 18 21 26.122 $w=2.98e-07 $l=6.8e-07 $layer=LI1_cond $X=0.245 $Y=1.66
+ $X2=0.245 $Y2=2.34
r101 16 59 3.0207 $w=3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.197 $Y2=2.72
r102 16 21 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.245 $Y2=2.34
r103 5 44 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=2
r104 4 38 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2
r105 3 32 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r106 2 27 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.34
r107 2 24 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.66
r108 1 21 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r109 1 18 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_6%X 1 2 3 4 5 6 21 23 25 27 28 29 33 37 39
+ 41 45 49 53 55 58 63 65
r111 63 65 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=3.91 $Y=1.495
+ $X2=3.91 $Y2=1.19
r112 61 63 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.55 $Y=1.58
+ $X2=3.91 $Y2=1.58
r113 58 65 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.91 $Y=0.905
+ $X2=3.91 $Y2=1.19
r114 49 61 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.55 $Y=2.34
+ $X2=3.55 $Y2=1.665
r115 43 58 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.55 $Y=0.82
+ $X2=3.91 $Y2=0.82
r116 43 45 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=3.55 $Y=0.735
+ $X2=3.55 $Y2=0.445
r117 42 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=1.58
+ $X2=2.61 $Y2=1.58
r118 41 61 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=1.58
+ $X2=3.55 $Y2=1.58
r119 41 42 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.385 $Y=1.58
+ $X2=2.775 $Y2=1.58
r120 40 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=0.82
+ $X2=2.61 $Y2=0.82
r121 39 43 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=0.82
+ $X2=3.55 $Y2=0.82
r122 39 40 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.385 $Y=0.82
+ $X2=2.775 $Y2=0.82
r123 35 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=1.58
r124 35 37 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=2.34
r125 31 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.735
+ $X2=2.61 $Y2=0.82
r126 31 33 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=2.61 $Y=0.735
+ $X2=2.61 $Y2=0.445
r127 30 52 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=1.58
+ $X2=1.67 $Y2=1.58
r128 29 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=1.58
+ $X2=2.61 $Y2=1.58
r129 29 30 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.445 $Y=1.58
+ $X2=1.835 $Y2=1.58
r130 27 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=0.82
+ $X2=2.61 $Y2=0.82
r131 27 28 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.445 $Y=0.82
+ $X2=1.835 $Y2=0.82
r132 23 52 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=1.58
r133 23 25 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=2.34
r134 19 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.67 $Y=0.735
+ $X2=1.835 $Y2=0.82
r135 19 21 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.67 $Y=0.735
+ $X2=1.67 $Y2=0.445
r136 6 61 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.66
r137 6 49 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2.34
r138 5 55 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.66
r139 5 37 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.34
r140 4 52 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r141 4 25 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
r142 3 45 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.235 $X2=3.55 $Y2=0.445
r143 2 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.47
+ $Y=0.235 $X2=2.61 $Y2=0.445
r144 1 21 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_6%VGND 1 2 3 4 5 16 18 22 24 28 30 34 36 40
+ 42 44 51 52 58 61 64 67
r67 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r68 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r69 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r70 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r71 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r72 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r73 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r74 52 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r75 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r76 49 67 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.155 $Y=0 $X2=4.02
+ $Y2=0
r77 49 51 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.155 $Y=0 $X2=4.37
+ $Y2=0
r78 48 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r79 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r80 45 55 3.97288 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.197
+ $Y2=0
r81 45 47 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.69
+ $Y2=0
r82 44 58 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.2
+ $Y2=0
r83 44 47 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.69
+ $Y2=0
r84 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r85 42 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r86 38 67 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0
r87 38 40 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0.4
r88 37 64 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.08
+ $Y2=0
r89 36 67 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.885 $Y=0 $X2=4.02
+ $Y2=0
r90 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.885 $Y=0 $X2=3.215
+ $Y2=0
r91 32 64 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0
r92 32 34 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.4
r93 31 61 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.14
+ $Y2=0
r94 30 64 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=3.08
+ $Y2=0
r95 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=2.275
+ $Y2=0
r96 26 61 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0
r97 26 28 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0.4
r98 25 58 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.2
+ $Y2=0
r99 24 61 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=2.14
+ $Y2=0
r100 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=0
+ $X2=1.335 $Y2=0
r101 20 58 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0
r102 20 22 15.3659 $w=2.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0.445
r103 16 55 3.17028 $w=2.5e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.197 $Y2=0
r104 16 18 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.38
r105 5 40 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.835
+ $Y=0.235 $X2=4.02 $Y2=0.4
r106 4 34 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.4
r107 3 28 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.235 $X2=2.14 $Y2=0.4
r108 2 22 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.445
r109 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

