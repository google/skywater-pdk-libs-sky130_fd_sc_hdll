* File: sky130_fd_sc_hdll__nor4_1.spice
* Created: Thu Aug 27 19:16:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nor4_1.pex.spice"
.subckt sky130_fd_sc_hdll__nor4_1  VNB VPB D C B A Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1006 N_Y_M1006_d N_D_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.2015 PD=0.97 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2 SB=75001.7
+ A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_C_M1001_g N_Y_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.104 PD=0.98 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1003 N_Y_M1003_d N_B_M1003_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65 AD=0.1105
+ AS=0.10725 PD=0.99 PS=0.98 NRD=0 NRS=10.152 M=1 R=4.33333 SA=75001.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.65 AD=0.1885
+ AS=0.1105 PD=1.88 PS=0.99 NRD=0 NRS=11.988 M=1 R=4.33333 SA=75001.7 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1004 A_117_297# N_D_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.18 W=1 AD=0.17 AS=0.27
+ PD=1.34 PS=2.54 NRD=22.6353 NRS=0.9653 M=1 R=5.55556 SA=90000.2 SB=90001.7
+ A=0.18 P=2.36 MULT=1
MM1000 A_221_297# N_C_M1000_g A_117_297# VPB PHIGHVT L=0.18 W=1 AD=0.15 AS=0.17
+ PD=1.3 PS=1.34 NRD=18.6953 NRS=22.6353 M=1 R=5.55556 SA=90000.7 SB=90001.1
+ A=0.18 P=2.36 MULT=1
MM1005 A_317_297# N_B_M1005_g A_221_297# VPB PHIGHVT L=0.18 W=1 AD=0.155 AS=0.15
+ PD=1.31 PS=1.3 NRD=19.6803 NRS=18.6953 M=1 R=5.55556 SA=90001.2 SB=90000.7
+ A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g A_317_297# VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.155 PD=2.54 PS=1.31 NRD=0.9653 NRS=19.6803 M=1 R=5.55556 SA=90001.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hdll__nor4_1.pxi.spice"
*
.ends
*
*
