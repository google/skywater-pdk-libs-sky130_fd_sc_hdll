* File: sky130_fd_sc_hdll__clkinvlp_4.pex.spice
* Created: Wed Sep  2 08:26:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKINVLP_4%A 3 7 11 15 19 23 27 31 33 34 48
c65 33 0 1.46135e-19 $X=0.23 $Y=0.85
r66 47 48 79.5619 $w=3.3e-07 $l=4.55e-07 $layer=POLY_cond $X=1.625 $Y=1.16
+ $X2=2.08 $Y2=1.16
r67 46 47 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=1.56 $Y=1.16
+ $X2=1.625 $Y2=1.16
r68 45 46 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=1.265 $Y=1.16
+ $X2=1.56 $Y2=1.16
r69 44 45 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.04 $Y=1.16
+ $X2=1.265 $Y2=1.16
r70 43 44 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.835 $Y=1.16
+ $X2=1.04 $Y2=1.16
r71 42 43 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=0.52 $Y=1.16
+ $X2=0.835 $Y2=1.16
r72 41 42 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=0.475 $Y=1.16
+ $X2=0.52 $Y2=1.16
r73 38 41 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.315 $Y=1.16
+ $X2=0.475 $Y2=1.16
r74 34 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.315
+ $Y=1.16 $X2=0.315 $Y2=1.16
r75 33 34 10.5076 $w=3.38e-07 $l=3.1e-07 $layer=LI1_cond $X=0.255 $Y=0.85
+ $X2=0.255 $Y2=1.16
r76 29 48 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.08 $Y=1.325
+ $X2=2.08 $Y2=1.16
r77 29 31 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.08 $Y=1.325
+ $X2=2.08 $Y2=1.985
r78 25 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.625 $Y=0.995
+ $X2=1.625 $Y2=1.16
r79 25 27 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.625 $Y=0.995
+ $X2=1.625 $Y2=0.51
r80 21 46 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.56 $Y=1.325
+ $X2=1.56 $Y2=1.16
r81 21 23 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.56 $Y=1.325
+ $X2=1.56 $Y2=1.985
r82 17 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.265 $Y=0.995
+ $X2=1.265 $Y2=1.16
r83 17 19 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.265 $Y=0.995
+ $X2=1.265 $Y2=0.51
r84 13 44 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.04 $Y=1.325
+ $X2=1.04 $Y2=1.16
r85 13 15 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.04 $Y=1.325
+ $X2=1.04 $Y2=1.985
r86 9 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.835 $Y=0.995
+ $X2=0.835 $Y2=1.16
r87 9 11 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.835 $Y=0.995
+ $X2=0.835 $Y2=0.51
r88 5 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=1.16
r89 5 7 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=0.51
r90 1 42 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.325
+ $X2=0.52 $Y2=1.16
r91 1 3 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.52 $Y=1.325 $X2=0.52
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINVLP_4%VPWR 1 2 3 10 12 18 22 24 29 30 31 37
+ 46
r38 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r39 40 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r40 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r41 37 45 4.10258 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.492 $Y2=2.72
r42 37 39 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.07 $Y2=2.72
r43 36 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r44 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r45 33 42 4.74282 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=0.42 $Y=2.72 $X2=0.21
+ $Y2=2.72
r46 33 35 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=0.42 $Y=2.72
+ $X2=1.15 $Y2=2.72
r47 31 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r48 31 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r49 29 35 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.15 $Y2=2.72
r50 29 30 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.322 $Y2=2.72
r51 28 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.46 $Y=2.72
+ $X2=2.07 $Y2=2.72
r52 28 30 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=1.46 $Y=2.72
+ $X2=1.322 $Y2=2.72
r53 24 27 29.2227 $w=2.78e-07 $l=7.1e-07 $layer=LI1_cond $X=2.365 $Y=1.63
+ $X2=2.365 $Y2=2.34
r54 22 45 3.25748 $w=2.8e-07 $l=1.64085e-07 $layer=LI1_cond $X=2.365 $Y=2.635
+ $X2=2.492 $Y2=2.72
r55 22 27 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=2.365 $Y=2.635
+ $X2=2.365 $Y2=2.34
r56 18 21 29.754 $w=2.73e-07 $l=7.1e-07 $layer=LI1_cond $X=1.322 $Y=1.63
+ $X2=1.322 $Y2=2.34
r57 16 30 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.322 $Y=2.635
+ $X2=1.322 $Y2=2.72
r58 16 21 12.3626 $w=2.73e-07 $l=2.95e-07 $layer=LI1_cond $X=1.322 $Y=2.635
+ $X2=1.322 $Y2=2.34
r59 12 15 24.1127 $w=3.23e-07 $l=6.8e-07 $layer=LI1_cond $X=0.257 $Y=1.66
+ $X2=0.257 $Y2=2.34
r60 10 42 2.9812 $w=3.25e-07 $l=1.05924e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.21 $Y2=2.72
r61 10 15 10.4606 $w=3.23e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.257 $Y2=2.34
r62 3 27 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.205
+ $Y=1.485 $X2=2.34 $Y2=2.34
r63 3 24 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.205
+ $Y=1.485 $X2=2.34 $Y2=1.63
r64 2 21 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.165
+ $Y=1.485 $X2=1.3 $Y2=2.34
r65 2 18 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.165
+ $Y=1.485 $X2=1.3 $Y2=1.63
r66 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r67 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINVLP_4%Y 1 2 3 10 14 18 19 20 21 22 23 47 52
r37 50 52 7.3214 $w=4.23e-07 $l=2.7e-07 $layer=LI1_cond $X=0.78 $Y=0.467
+ $X2=1.05 $Y2=0.467
r38 42 50 1.87632 $w=3.5e-07 $l=2.13e-07 $layer=LI1_cond $X=0.78 $Y=0.68
+ $X2=0.78 $Y2=0.467
r39 23 43 4.32773 $w=3.45e-07 $l=1.4e-07 $layer=LI1_cond $X=0.78 $Y=1.155
+ $X2=0.78 $Y2=1.015
r40 23 30 4.32773 $w=3.45e-07 $l=1.42478e-07 $layer=LI1_cond $X=0.78 $Y=1.155
+ $X2=0.775 $Y2=1.295
r41 22 43 5.43295 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.78 $Y=0.85
+ $X2=0.78 $Y2=1.015
r42 22 42 5.59758 $w=3.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.78 $Y=0.85
+ $X2=0.78 $Y2=0.68
r43 21 50 1.03042 $w=4.23e-07 $l=3.8e-08 $layer=LI1_cond $X=0.742 $Y=0.467
+ $X2=0.78 $Y2=0.467
r44 21 47 1.41005 $w=4.23e-07 $l=5.2e-08 $layer=LI1_cond $X=0.742 $Y=0.467
+ $X2=0.69 $Y2=0.467
r45 20 40 4.4064 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=0.775 $Y=2.21
+ $X2=0.775 $Y2=2.34
r46 19 20 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.775 $Y=1.87
+ $X2=0.775 $Y2=2.21
r47 19 34 8.13489 $w=3.38e-07 $l=2.4e-07 $layer=LI1_cond $X=0.775 $Y=1.87
+ $X2=0.775 $Y2=1.63
r48 18 34 3.38954 $w=3.38e-07 $l=1e-07 $layer=LI1_cond $X=0.775 $Y=1.53
+ $X2=0.775 $Y2=1.63
r49 18 30 7.96542 $w=3.38e-07 $l=2.35e-07 $layer=LI1_cond $X=0.775 $Y=1.53
+ $X2=0.775 $Y2=1.295
r50 14 16 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.82 $Y=1.63 $X2=1.82
+ $Y2=2.34
r51 12 14 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.82 $Y=1.295
+ $X2=1.82 $Y2=1.63
r52 11 23 2.10399 $w=2.8e-07 $l=1.75e-07 $layer=LI1_cond $X=0.955 $Y=1.155
+ $X2=0.78 $Y2=1.155
r53 10 12 6.87623 $w=2.8e-07 $l=2.24332e-07 $layer=LI1_cond $X=1.655 $Y=1.155
+ $X2=1.82 $Y2=1.295
r54 10 11 28.8111 $w=2.78e-07 $l=7e-07 $layer=LI1_cond $X=1.655 $Y=1.155
+ $X2=0.955 $Y2=1.155
r55 3 16 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.685
+ $Y=1.485 $X2=1.82 $Y2=2.34
r56 3 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.685
+ $Y=1.485 $X2=1.82 $Y2=1.63
r57 2 40 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.645
+ $Y=1.485 $X2=0.78 $Y2=2.34
r58 2 34 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.645
+ $Y=1.485 $X2=0.78 $Y2=1.63
r59 1 52 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.235 $X2=1.05 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINVLP_4%VGND 1 2 7 9 13 16 17 18 28 29
c30 7 0 1.46135e-19 $X=0.26 $Y=0.085
r31 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r32 26 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r33 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r34 23 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r35 22 25 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r36 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r37 20 32 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r38 20 22 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r39 18 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r40 18 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r41 16 25 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=1.675 $Y=0 $X2=1.61
+ $Y2=0
r42 16 17 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=1.675 $Y=0 $X2=1.837
+ $Y2=0
r43 15 28 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2 $Y=0 $X2=2.53
+ $Y2=0
r44 15 17 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=2 $Y=0 $X2=1.837
+ $Y2=0
r45 11 17 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.837 $Y=0.085
+ $X2=1.837 $Y2=0
r46 11 13 15.0704 $w=3.23e-07 $l=4.25e-07 $layer=LI1_cond $X=1.837 $Y=0.085
+ $X2=1.837 $Y2=0.51
r47 7 32 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r48 7 9 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.43
r49 2 13 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.7
+ $Y=0.235 $X2=1.835 $Y2=0.51
r50 1 9 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends

