# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nand2_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand2_12 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  3.330000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.625000 1.055000 10.695000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  3.330000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.335000 1.055000 5.765000 1.325000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  4.858000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.565000 1.495000 11.235000 1.665000 ;
        RECT  0.565000 1.665000  0.895000 2.465000 ;
        RECT  1.505000 1.665000  1.835000 2.465000 ;
        RECT  2.445000 1.665000  2.775000 2.465000 ;
        RECT  3.385000 1.665000  3.715000 2.465000 ;
        RECT  4.325000 1.665000  4.655000 2.465000 ;
        RECT  5.265000 1.665000  5.595000 2.465000 ;
        RECT  6.045000 1.055000  6.455000 1.495000 ;
        RECT  6.155000 0.635000 11.235000 0.885000 ;
        RECT  6.155000 0.885000  6.455000 1.055000 ;
        RECT  6.205000 1.665000  6.535000 2.465000 ;
        RECT  7.145000 1.665000  7.475000 2.465000 ;
        RECT  8.085000 1.665000  8.415000 2.465000 ;
        RECT  9.025000 1.665000  9.355000 2.465000 ;
        RECT  9.965000 1.665000 10.295000 2.465000 ;
        RECT 10.905000 1.665000 11.235000 2.465000 ;
        RECT 10.965000 0.885000 11.235000 1.055000 ;
        RECT 10.965000 1.055000 11.435000 1.325000 ;
        RECT 10.965000 1.325000 11.235000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.150000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.090000  0.255000  0.425000 0.715000 ;
      RECT  0.090000  0.715000  5.985000 0.885000 ;
      RECT  0.125000  1.495000  0.395000 2.635000 ;
      RECT  0.595000  0.085000  0.865000 0.545000 ;
      RECT  1.035000  0.255000  1.365000 0.715000 ;
      RECT  1.065000  1.835000  1.335000 2.635000 ;
      RECT  1.535000  0.085000  1.805000 0.545000 ;
      RECT  1.975000  0.255000  2.305000 0.715000 ;
      RECT  2.005000  1.835000  2.275000 2.635000 ;
      RECT  2.475000  0.085000  2.745000 0.545000 ;
      RECT  2.915000  0.255000  3.245000 0.715000 ;
      RECT  2.945000  1.835000  3.215000 2.635000 ;
      RECT  3.415000  0.085000  3.685000 0.545000 ;
      RECT  3.855000  0.255000  4.185000 0.715000 ;
      RECT  3.885000  1.835000  4.155000 2.635000 ;
      RECT  4.355000  0.085000  4.625000 0.545000 ;
      RECT  4.795000  0.255000  5.125000 0.715000 ;
      RECT  4.825000  1.835000  5.095000 2.635000 ;
      RECT  5.295000  0.085000  5.565000 0.545000 ;
      RECT  5.735000  0.255000 11.705000 0.465000 ;
      RECT  5.735000  0.465000  5.985000 0.715000 ;
      RECT  5.765000  1.835000  6.035000 2.635000 ;
      RECT  6.705000  1.835000  6.975000 2.635000 ;
      RECT  7.645000  1.835000  7.915000 2.635000 ;
      RECT  8.585000  1.835000  8.855000 2.635000 ;
      RECT  9.525000  1.835000  9.795000 2.635000 ;
      RECT 10.465000  1.835000 10.735000 2.635000 ;
      RECT 11.405000  1.495000 11.675000 2.635000 ;
      RECT 11.455000  0.465000 11.705000 0.885000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2_12
END LIBRARY
