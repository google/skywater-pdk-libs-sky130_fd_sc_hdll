# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__or2_6
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.415000 1.075000 1.085000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.075000 2.025000 1.275000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.396500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985000 0.255000 3.285000 0.725000 ;
        RECT 2.985000 0.725000 5.415000 0.905000 ;
        RECT 2.985000 1.495000 5.415000 1.665000 ;
        RECT 2.985000 1.665000 3.315000 2.465000 ;
        RECT 3.925000 1.665000 4.255000 2.465000 ;
        RECT 3.955000 0.255000 4.225000 0.725000 ;
        RECT 4.865000 1.665000 5.195000 2.465000 ;
        RECT 4.895000 0.255000 5.165000 0.725000 ;
        RECT 5.015000 0.905000 5.415000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.090000  1.455000 1.355000 1.665000 ;
      RECT 0.090000  1.665000 0.415000 2.465000 ;
      RECT 0.145000  0.085000 0.415000 0.905000 ;
      RECT 0.585000  0.255000 0.915000 0.725000 ;
      RECT 0.585000  0.725000 1.855000 0.735000 ;
      RECT 0.585000  0.735000 2.375000 0.905000 ;
      RECT 0.585000  1.835000 0.915000 2.635000 ;
      RECT 1.085000  0.085000 1.355000 0.555000 ;
      RECT 1.085000  1.665000 1.355000 2.295000 ;
      RECT 1.085000  2.295000 2.325000 2.465000 ;
      RECT 1.525000  0.255000 1.855000 0.725000 ;
      RECT 1.525000  1.445000 2.375000 1.665000 ;
      RECT 1.525000  1.665000 1.855000 2.125000 ;
      RECT 2.025000  0.085000 2.815000 0.555000 ;
      RECT 2.025000  1.835000 2.325000 2.295000 ;
      RECT 2.195000  0.905000 2.375000 1.075000 ;
      RECT 2.195000  1.075000 4.845000 1.275000 ;
      RECT 2.195000  1.275000 2.375000 1.445000 ;
      RECT 2.545000  0.555000 2.815000 0.905000 ;
      RECT 2.545000  1.495000 2.815000 2.635000 ;
      RECT 3.455000  0.085000 3.785000 0.555000 ;
      RECT 3.485000  1.835000 3.755000 2.635000 ;
      RECT 4.395000  0.085000 4.725000 0.555000 ;
      RECT 4.425000  1.835000 4.695000 2.635000 ;
      RECT 5.335000  0.085000 5.665000 0.555000 ;
      RECT 5.365000  1.835000 5.635000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2_6
