* File: sky130_fd_sc_hdll__sdlclkp_1.pex.spice
* Created: Wed Sep  2 08:52:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_1%SCE 2 3 5 8 10 11 19
c29 8 0 1.15416e-19 $X=0.52 $Y=0.445
c30 3 0 1.81037e-19 $X=0.495 $Y=1.77
r31 18 19 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r32 15 18 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.495 $Y2=1.16
r33 10 11 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.207 $Y=1.16
+ $X2=0.207 $Y2=1.53
r34 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r35 6 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.16
r36 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r37 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.77
+ $X2=0.495 $Y2=2.165
r38 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.67 $X2=0.495
+ $Y2=1.77
r39 1 18 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r40 1 2 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_1%GATE 2 3 5 8 10 11 15 16
c40 16 0 3.25666e-19 $X=0.94 $Y=1.16
c41 15 0 9.19878e-20 $X=0.94 $Y=1.16
c42 2 0 1.70274e-19 $X=0.905 $Y=1.67
r43 15 18 39.5599 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=0.957 $Y=1.16
+ $X2=0.957 $Y2=1.325
r44 15 17 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=0.957 $Y=1.16
+ $X2=0.957 $Y2=0.995
r45 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r46 10 11 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=1.045 $Y=1.53
+ $X2=1.045 $Y2=1.87
r47 10 16 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.045 $Y=1.53
+ $X2=1.045 $Y2=1.16
r48 8 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.945 $Y=0.445
+ $X2=0.945 $Y2=0.995
r49 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.905 $Y=1.77
+ $X2=0.905 $Y2=2.165
r50 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.905 $Y=1.67 $X2=0.905
+ $Y2=1.77
r51 2 18 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=0.905 $Y=1.67
+ $X2=0.905 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_269_21# 1 2 9 11 13 16 18 21 25 26 28
+ 34 36 37 38 41 45 47 49 50 51 54 57
c174 50 0 1.44161e-19 $X=4.305 $Y=1.53
c175 47 0 3.87639e-19 $X=1.712 $Y=1.452
c176 34 0 1.48075e-19 $X=4.457 $Y=1.495
c177 25 0 2.99785e-20 $X=1.55 $Y=0.87
c178 9 0 2.2455e-20 $X=1.42 $Y=0.415
r179 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.875
+ $Y=1.74 $X2=1.875 $Y2=1.74
r180 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.45 $Y=1.53
+ $X2=4.45 $Y2=1.53
r181 54 66 5.07427 $w=4.93e-07 $l=2.1e-07 $layer=LI1_cond $X=1.712 $Y=1.53
+ $X2=1.712 $Y2=1.74
r182 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.71 $Y=1.53
+ $X2=1.71 $Y2=1.53
r183 51 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.855 $Y=1.53
+ $X2=1.71 $Y2=1.53
r184 50 57 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.305 $Y=1.53
+ $X2=4.45 $Y2=1.53
r185 50 51 3.03217 $w=1.4e-07 $l=2.45e-06 $layer=MET1_cond $X=4.305 $Y=1.53
+ $X2=1.855 $Y2=1.53
r186 47 54 1.88473 $w=4.93e-07 $l=7.8e-08 $layer=LI1_cond $X=1.712 $Y=1.452
+ $X2=1.712 $Y2=1.53
r187 47 48 7.22426 $w=4.93e-07 $l=2.47e-07 $layer=LI1_cond $X=1.712 $Y=1.452
+ $X2=1.712 $Y2=1.205
r188 43 45 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=5.09 $Y=0.615
+ $X2=5.09 $Y2=0.465
r189 39 58 2.99321 $w=2.5e-07 $l=9.3e-08 $layer=LI1_cond $X=4.55 $Y=1.62
+ $X2=4.457 $Y2=1.62
r190 39 41 23.0489 $w=2.48e-07 $l=5e-07 $layer=LI1_cond $X=4.55 $Y=1.62 $X2=5.05
+ $Y2=1.62
r191 37 43 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.965 $Y=0.7
+ $X2=5.09 $Y2=0.615
r192 37 38 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.965 $Y=0.7
+ $X2=4.55 $Y2=0.7
r193 36 49 4.98297 $w=1.77e-07 $l=8.89101e-08 $layer=LI1_cond $X=4.465 $Y=1.105
+ $X2=4.457 $Y2=1.19
r194 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.465 $Y=0.785
+ $X2=4.55 $Y2=0.7
r195 35 36 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.465 $Y=0.785
+ $X2=4.465 $Y2=1.105
r196 34 58 4.02313 $w=1.85e-07 $l=1.25e-07 $layer=LI1_cond $X=4.457 $Y=1.495
+ $X2=4.457 $Y2=1.62
r197 33 49 4.98297 $w=1.77e-07 $l=8.5e-08 $layer=LI1_cond $X=4.457 $Y=1.275
+ $X2=4.457 $Y2=1.19
r198 33 34 13.1892 $w=1.83e-07 $l=2.2e-07 $layer=LI1_cond $X=4.457 $Y=1.275
+ $X2=4.457 $Y2=1.495
r199 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.28
+ $Y=1.19 $X2=4.28 $Y2=1.19
r200 28 49 1.49848 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=4.365 $Y=1.19
+ $X2=4.457 $Y2=1.19
r201 28 30 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.365 $Y=1.19
+ $X2=4.28 $Y2=1.19
r202 26 60 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=1.55 $Y=0.87
+ $X2=1.42 $Y2=0.87
r203 25 48 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=1.632 $Y=0.87
+ $X2=1.632 $Y2=1.205
r204 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.55
+ $Y=0.87 $X2=1.55 $Y2=0.87
r205 18 31 48.0587 $w=2.96e-07 $l=2.80624e-07 $layer=POLY_cond $X=4.215 $Y=1.44
+ $X2=4.28 $Y2=1.19
r206 18 21 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=4.215 $Y=1.44
+ $X2=4.215 $Y2=1.835
r207 14 31 43.457 $w=2.96e-07 $l=2.35743e-07 $layer=POLY_cond $X=4.19 $Y=0.995
+ $X2=4.28 $Y2=1.19
r208 14 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.19 $Y=0.995
+ $X2=4.19 $Y2=0.445
r209 11 65 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=1.96 $Y=1.99
+ $X2=1.9 $Y2=1.74
r210 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.96 $Y=1.99
+ $X2=1.96 $Y2=2.275
r211 7 60 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.42 $Y=0.735
+ $X2=1.42 $Y2=0.87
r212 7 9 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.42 $Y=0.735
+ $X2=1.42 $Y2=0.415
r213 2 41 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.905
+ $Y=1.515 $X2=5.05 $Y2=1.66
r214 1 45 182 $w=1.7e-07 $l=3.0895e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.235 $X2=5.05 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_266_243# 1 2 8 9 11 12 13 16 18 21 24
+ 28 30 31 37 38 41 42 43
c116 42 0 2.2455e-20 $X=2.06 $Y=0.87
c117 41 0 2.73089e-19 $X=2.06 $Y=0.87
c118 28 0 1.17835e-19 $X=3.98 $Y=1.66
c119 18 0 2.92127e-20 $X=2.022 $Y=1.215
c120 8 0 3.15944e-20 $X=1.43 $Y=1.89
r121 41 44 41.3874 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.06 $Y=0.87
+ $X2=2.06 $Y2=1.035
r122 41 43 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.06 $Y=0.87
+ $X2=2.06 $Y2=0.705
r123 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.06
+ $Y=0.87 $X2=2.06 $Y2=0.87
r124 38 49 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.9 $Y=0.85 $X2=3.9
+ $Y2=0.935
r125 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.885 $Y=0.85
+ $X2=3.885 $Y2=0.85
r126 33 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.22 $Y=0.85
+ $X2=2.22 $Y2=0.85
r127 31 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.365 $Y=0.85
+ $X2=2.22 $Y2=0.85
r128 30 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.74 $Y=0.85
+ $X2=3.885 $Y2=0.85
r129 30 31 1.70173 $w=1.4e-07 $l=1.375e-06 $layer=MET1_cond $X=3.74 $Y=0.85
+ $X2=2.365 $Y2=0.85
r130 25 28 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.82 $Y=1.66
+ $X2=3.98 $Y2=1.66
r131 24 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.82 $Y=1.575
+ $X2=3.82 $Y2=1.66
r132 24 49 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.82 $Y=1.575
+ $X2=3.82 $Y2=0.935
r133 19 38 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.9 $Y=0.77 $X2=3.9
+ $Y2=0.85
r134 19 21 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=3.9 $Y=0.77
+ $X2=3.9 $Y2=0.465
r135 18 44 61.2142 $w=1.95e-07 $l=1.8e-07 $layer=POLY_cond $X=2.022 $Y=1.215
+ $X2=2.022 $Y2=1.035
r136 16 43 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2 $Y=0.415 $X2=2
+ $Y2=0.705
r137 12 18 27.531 $w=1.5e-07 $l=1.29167e-07 $layer=POLY_cond $X=1.925 $Y=1.29
+ $X2=2.022 $Y2=1.215
r138 12 13 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.925 $Y=1.29
+ $X2=1.53 $Y2=1.29
r139 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.43 $Y=1.99
+ $X2=1.43 $Y2=2.275
r140 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.43 $Y=1.89 $X2=1.43
+ $Y2=1.99
r141 7 13 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=1.43 $Y=1.365
+ $X2=1.53 $Y2=1.29
r142 7 8 174.078 $w=2e-07 $l=5.25e-07 $layer=POLY_cond $X=1.43 $Y=1.365 $X2=1.43
+ $Y2=1.89
r143 2 28 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.855
+ $Y=1.515 $X2=3.98 $Y2=1.66
r144 1 21 182 $w=1.7e-07 $l=2.85745e-07 $layer=licon1_NDIFF $count=1 $X=3.855
+ $Y=0.235 $X2=3.98 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_484_315# 1 2 7 9 12 15 16 18 21 23 27
+ 31 33 37 44 45 50
c130 37 0 1.04371e-19 $X=5.61 $Y=1.16
c131 33 0 5.75693e-20 $X=5.385 $Y=2
c132 12 0 1.25378e-19 $X=2.655 $Y=0.445
r133 49 50 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=5.805 $Y=1.16
+ $X2=5.83 $Y2=1.16
r134 41 44 4.25649 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=2.555 $Y=1.74
+ $X2=2.665 $Y2=1.74
r135 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.555
+ $Y=1.74 $X2=2.555 $Y2=1.74
r136 38 49 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=5.61 $Y=1.16
+ $X2=5.805 $Y2=1.16
r137 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.61
+ $Y=1.16 $X2=5.61 $Y2=1.16
r138 35 37 24.8598 $w=3.48e-07 $l=7.55e-07 $layer=LI1_cond $X=5.56 $Y=1.915
+ $X2=5.56 $Y2=1.16
r139 34 45 2.69039 $w=1.7e-07 $l=1.87083e-07 $layer=LI1_cond $X=3.545 $Y=2
+ $X2=3.435 $Y2=1.86
r140 33 35 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=5.385 $Y=2
+ $X2=5.56 $Y2=1.915
r141 33 34 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=5.385 $Y=2
+ $X2=3.545 $Y2=2
r142 29 45 3.42573 $w=1.7e-07 $l=2.37171e-07 $layer=LI1_cond $X=3.46 $Y=1.635
+ $X2=3.435 $Y2=1.86
r143 29 31 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=3.46 $Y=1.635
+ $X2=3.46 $Y2=0.42
r144 25 45 3.42573 $w=2.2e-07 $l=2.25e-07 $layer=LI1_cond $X=3.435 $Y=2.085
+ $X2=3.435 $Y2=1.86
r145 25 27 6.28605 $w=2.18e-07 $l=1.2e-07 $layer=LI1_cond $X=3.435 $Y=2.085
+ $X2=3.435 $Y2=2.205
r146 23 45 2.69039 $w=2.7e-07 $l=1.48324e-07 $layer=LI1_cond $X=3.325 $Y=1.77
+ $X2=3.435 $Y2=1.86
r147 23 44 28.1708 $w=2.68e-07 $l=6.6e-07 $layer=LI1_cond $X=3.325 $Y=1.77
+ $X2=2.665 $Y2=1.77
r148 19 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.83 $Y=0.995
+ $X2=5.83 $Y2=1.16
r149 19 21 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.83 $Y=0.995
+ $X2=5.83 $Y2=0.445
r150 16 18 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=5.805 $Y=1.77
+ $X2=5.805 $Y2=2.165
r151 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=5.805 $Y=1.67 $X2=5.805
+ $Y2=1.77
r152 14 49 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=5.805 $Y=1.325
+ $X2=5.805 $Y2=1.16
r153 14 15 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=5.805 $Y=1.325
+ $X2=5.805 $Y2=1.67
r154 10 42 38.6443 $w=2.87e-07 $l=2.0106e-07 $layer=POLY_cond $X=2.655 $Y=1.575
+ $X2=2.575 $Y2=1.74
r155 10 12 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=2.655 $Y=1.575
+ $X2=2.655 $Y2=0.445
r156 7 42 48.651 $w=2.87e-07 $l=2.76134e-07 $layer=POLY_cond $X=2.52 $Y=1.99
+ $X2=2.575 $Y2=1.74
r157 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.52 $Y=1.99
+ $X2=2.52 $Y2=2.275
r158 2 27 600 $w=1.7e-07 $l=7.89177e-07 $layer=licon1_PDIFF $count=1 $X=3.315
+ $Y=1.485 $X2=3.46 $Y2=2.205
r159 1 31 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.325
+ $Y=0.235 $X2=3.46 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_299_47# 1 2 7 9 10 12 13 17 22 23 24
+ 26 29 32
c102 32 0 1.28928e-19 $X=2.56 $Y=1.185
c103 26 0 2.99785e-20 $X=2.56 $Y=0.995
c104 24 0 3.15944e-20 $X=2.3 $Y=1.29
r105 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.12
+ $Y=1.16 $X2=3.12 $Y2=1.16
r106 27 32 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=1.185
+ $X2=2.56 $Y2=1.185
r107 27 29 14.4055 $w=3.78e-07 $l=4.75e-07 $layer=LI1_cond $X=2.645 $Y=1.185
+ $X2=3.12 $Y2=1.185
r108 26 32 3.11956 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.56 $Y=0.995
+ $X2=2.56 $Y2=1.185
r109 25 26 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.56 $Y=0.535
+ $X2=2.56 $Y2=0.995
r110 23 32 3.40559 $w=2.75e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.475 $Y=1.29
+ $X2=2.56 $Y2=1.185
r111 23 24 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.475 $Y=1.29
+ $X2=2.3 $Y2=1.29
r112 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.215 $Y=1.375
+ $X2=2.3 $Y2=1.29
r113 21 22 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.215 $Y=1.375
+ $X2=2.215 $Y2=2.125
r114 17 22 7.85115 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.13 $Y=2.295
+ $X2=2.215 $Y2=2.125
r115 17 19 14.7445 $w=3.38e-07 $l=4.35e-07 $layer=LI1_cond $X=2.13 $Y=2.295
+ $X2=1.695 $Y2=2.295
r116 13 25 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.475 $Y=0.395
+ $X2=2.56 $Y2=0.535
r117 13 15 30.6632 $w=2.78e-07 $l=7.45e-07 $layer=LI1_cond $X=2.475 $Y=0.395
+ $X2=1.73 $Y2=0.395
r118 10 30 38.532 $w=3.11e-07 $l=2.07123e-07 $layer=POLY_cond $X=3.25 $Y=0.995
+ $X2=3.155 $Y2=1.16
r119 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.25 $Y=0.995
+ $X2=3.25 $Y2=0.56
r120 7 30 47.2262 $w=3.11e-07 $l=2.82843e-07 $layer=POLY_cond $X=3.225 $Y=1.41
+ $X2=3.155 $Y2=1.16
r121 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.225 $Y=1.41
+ $X2=3.225 $Y2=1.985
r122 2 19 600 $w=1.7e-07 $l=3e-07 $layer=licon1_PDIFF $count=1 $X=1.52 $Y=2.065
+ $X2=1.695 $Y2=2.29
r123 1 15 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.73 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_1%CLK 3 5 8 10 11 13 16 19 20 22 23 25 31
+ 36 44
c95 36 0 1.64862e-19 $X=4.89 $Y=1.19
c96 11 0 1.6194e-19 $X=6.285 $Y=1.77
c97 8 0 1.17835e-19 $X=4.815 $Y=1.835
r98 31 34 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.25 $Y=1.16
+ $X2=6.25 $Y2=1.325
r99 31 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.25 $Y=1.16
+ $X2=6.25 $Y2=0.995
r100 28 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.925
+ $Y=1.16 $X2=4.925 $Y2=1.16
r101 25 44 0.00320802 $w=2.3e-07 $l=5e-09 $layer=MET1_cond $X=4.83 $Y=1.19
+ $X2=4.825 $Y2=1.19
r102 25 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.89 $Y=1.19
+ $X2=4.89 $Y2=1.19
r103 23 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.25
+ $Y=1.16 $X2=6.25 $Y2=1.16
r104 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.085 $Y=1.19
+ $X2=6.085 $Y2=1.19
r105 20 25 0.153963 $w=2.3e-07 $l=2.05e-07 $layer=MET1_cond $X=5.035 $Y=1.19
+ $X2=4.83 $Y2=1.19
r106 19 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.94 $Y=1.19
+ $X2=6.085 $Y2=1.19
r107 19 20 1.12005 $w=1.4e-07 $l=9.05e-07 $layer=MET1_cond $X=5.94 $Y=1.19
+ $X2=5.035 $Y2=1.19
r108 16 33 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.31 $Y=0.445
+ $X2=6.31 $Y2=0.995
r109 11 13 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=6.285 $Y=1.77
+ $X2=6.285 $Y2=2.165
r110 10 11 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=6.285 $Y=1.67 $X2=6.285
+ $Y2=1.77
r111 10 34 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=6.285 $Y=1.67
+ $X2=6.285 $Y2=1.325
r112 5 28 52.1409 $w=3.07e-07 $l=3.13943e-07 $layer=POLY_cond $X=4.815 $Y=1.44
+ $X2=4.887 $Y2=1.16
r113 5 8 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=4.815 $Y=1.44
+ $X2=4.815 $Y2=1.835
r114 1 28 38.5336 $w=3.07e-07 $l=2.07918e-07 $layer=POLY_cond $X=4.79 $Y=0.995
+ $X2=4.887 $Y2=1.16
r115 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.79 $Y=0.995
+ $X2=4.79 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_1089_47# 1 2 7 9 10 12 15 17 18 19 25
+ 29
c74 25 0 1.74496e-19 $X=6.73 $Y=1.16
r75 27 29 13.988 $w=5.88e-07 $l=6.9e-07 $layer=LI1_cond $X=6.04 $Y=1.79 $X2=6.73
+ $Y2=1.79
r76 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.73
+ $Y=1.16 $X2=6.73 $Y2=1.16
r77 23 29 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=6.73 $Y=1.495
+ $X2=6.73 $Y2=1.79
r78 23 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.73 $Y=1.495
+ $X2=6.73 $Y2=1.16
r79 22 25 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.73 $Y=0.785
+ $X2=6.73 $Y2=1.16
r80 19 27 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=6.04 $Y=2.085
+ $X2=6.04 $Y2=1.79
r81 19 21 2.87059 $w=1.7e-07 $l=4e-08 $layer=LI1_cond $X=6.04 $Y=2.085 $X2=6.04
+ $Y2=2.125
r82 17 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.645 $Y=0.7
+ $X2=6.73 $Y2=0.785
r83 17 18 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=6.645 $Y=0.7
+ $X2=5.705 $Y2=0.7
r84 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.62 $Y=0.615
+ $X2=5.705 $Y2=0.7
r85 13 15 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.62 $Y=0.615
+ $X2=5.62 $Y2=0.46
r86 10 26 38.6072 $w=2.91e-07 $l=2.02287e-07 $layer=POLY_cond $X=6.835 $Y=0.995
+ $X2=6.752 $Y2=1.16
r87 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.835 $Y=0.995
+ $X2=6.835 $Y2=0.56
r88 7 26 48.3784 $w=2.91e-07 $l=2.77489e-07 $layer=POLY_cond $X=6.81 $Y=1.41
+ $X2=6.752 $Y2=1.16
r89 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.81 $Y=1.41 $X2=6.81
+ $Y2=1.985
r90 2 21 600 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_PDIFF $count=1 $X=5.895
+ $Y=1.845 $X2=6.04 $Y2=2.125
r91 1 15 182 $w=1.7e-07 $l=3e-07 $layer=licon1_NDIFF $count=1 $X=5.445 $Y=0.235
+ $X2=5.62 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_1%VPWR 1 2 3 4 5 16 18 24 27 30 32 33 34
+ 41 54 55 63 69 73
c93 5 0 1.74496e-19 $X=6.375 $Y=1.845
r94 71 73 6.78742 $w=5.48e-07 $l=2.5e-08 $layer=LI1_cond $X=3.91 $Y=2.53
+ $X2=3.885 $Y2=2.53
r95 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r96 69 73 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.105 $Y=2.72
+ $X2=3.885 $Y2=2.72
r97 68 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r98 67 69 10.1774 $w=7.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.99 $Y=2.44
+ $X2=3.105 $Y2=2.44
r99 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r100 65 67 1.72039 $w=7.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.885 $Y=2.44
+ $X2=2.99 $Y2=2.44
r101 62 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r102 61 65 5.81655 $w=7.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.53 $Y=2.44
+ $X2=2.885 $Y2=2.44
r103 61 63 8.45698 $w=7.28e-07 $l=1e-08 $layer=LI1_cond $X=2.53 $Y=2.44 $X2=2.52
+ $Y2=2.44
r104 61 62 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r105 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r106 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r107 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r108 49 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r109 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r110 46 48 16.8538 $w=5.48e-07 $l=7.75e-07 $layer=LI1_cond $X=4.515 $Y=2.53
+ $X2=5.29 $Y2=2.53
r111 44 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r112 44 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r113 43 46 3.1533 $w=5.48e-07 $l=1.45e-07 $layer=LI1_cond $X=4.37 $Y=2.53
+ $X2=4.515 $Y2=2.53
r114 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r115 41 71 5.43672 $w=5.48e-07 $l=2.5e-07 $layer=LI1_cond $X=4.16 $Y=2.53
+ $X2=3.91 $Y2=2.53
r116 41 43 4.56684 $w=5.48e-07 $l=2.1e-07 $layer=LI1_cond $X=4.16 $Y=2.53
+ $X2=4.37 $Y2=2.53
r117 40 62 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r118 39 63 119.39 $w=1.68e-07 $l=1.83e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.52 $Y2=2.72
r119 39 40 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r120 37 58 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r121 37 39 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r122 34 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r123 34 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r124 32 51 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.385 $Y=2.72
+ $X2=6.21 $Y2=2.72
r125 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.385 $Y=2.72
+ $X2=6.55 $Y2=2.72
r126 31 54 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.715 $Y=2.72
+ $X2=7.13 $Y2=2.72
r127 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.715 $Y=2.72
+ $X2=6.55 $Y2=2.72
r128 30 51 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=5.735 $Y=2.72
+ $X2=6.21 $Y2=2.72
r129 29 30 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.57 $Y=2.53
+ $X2=5.735 $Y2=2.53
r130 27 48 3.69697 $w=5.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.46 $Y=2.53
+ $X2=5.29 $Y2=2.53
r131 27 29 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=5.46 $Y=2.53
+ $X2=5.57 $Y2=2.53
r132 22 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.55 $Y=2.635
+ $X2=6.55 $Y2=2.72
r133 22 24 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.55 $Y=2.635
+ $X2=6.55 $Y2=2.36
r134 16 58 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r135 16 18 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2
r136 5 24 600 $w=1.7e-07 $l=5.96112e-07 $layer=licon1_PDIFF $count=1 $X=6.375
+ $Y=1.845 $X2=6.55 $Y2=2.36
r137 4 29 600 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_PDIFF $count=1 $X=5.445
+ $Y=1.845 $X2=5.57 $Y2=2.34
r138 3 46 600 $w=1.7e-07 $l=9.24054e-07 $layer=licon1_PDIFF $count=1 $X=4.305
+ $Y=1.515 $X2=4.515 $Y2=2.34
r139 2 65 600 $w=1.7e-07 $l=4.10061e-07 $layer=licon1_PDIFF $count=1 $X=2.61
+ $Y=2.065 $X2=2.885 $Y2=2.36
r140 1 18 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_27_47# 1 2 3 12 15 16 17 18 20 24
c53 24 0 1.74968e-19 $X=1.2 $Y=0.42
r54 22 24 12.0152 $w=1.78e-07 $l=1.95e-07 $layer=LI1_cond $X=1.205 $Y=0.615
+ $X2=1.205 $Y2=0.42
r55 18 20 17.2866 $w=3.38e-07 $l=5.1e-07 $layer=LI1_cond $X=0.685 $Y=2.295
+ $X2=1.195 $Y2=2.295
r56 17 28 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=0.7 $X2=0.6
+ $Y2=0.7
r57 16 22 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.115 $Y=0.7
+ $X2=1.205 $Y2=0.615
r58 16 17 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.115 $Y=0.7
+ $X2=0.685 $Y2=0.7
r59 15 18 7.85115 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.6 $Y=2.125
+ $X2=0.685 $Y2=2.295
r60 14 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.6 $Y=0.785 $X2=0.6
+ $Y2=0.7
r61 14 15 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=0.6 $Y=0.785
+ $X2=0.6 $Y2=2.125
r62 10 28 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.215 $Y=0.7
+ $X2=0.6 $Y2=0.7
r63 10 12 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=0.215 $Y=0.615
+ $X2=0.215 $Y2=0.43
r64 3 20 600 $w=1.7e-07 $l=5.35747e-07 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.845 $X2=1.195 $Y2=2.29
r65 2 24 182 $w=1.7e-07 $l=2.59856e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.235 $X2=1.2 $Y2=0.42
r66 1 12 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_1%GCLK 1 2 7 8 9 10
r14 9 10 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=7.11 $Y=1.815
+ $X2=7.11 $Y2=2.21
r15 8 9 28.8111 $w=2.48e-07 $l=6.25e-07 $layer=LI1_cond $X=7.11 $Y=1.19 $X2=7.11
+ $Y2=1.815
r16 8 19 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=7.11 $Y=1.19 $X2=7.11
+ $Y2=0.64
r17 7 19 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=7.11 $Y=0.51 $X2=7.11
+ $Y2=0.64
r18 2 9 300 $w=1.7e-07 $l=4.06202e-07 $layer=licon1_PDIFF $count=2 $X=6.9
+ $Y=1.485 $X2=7.07 $Y2=1.815
r19 1 19 182 $w=1.7e-07 $l=4.78357e-07 $layer=licon1_NDIFF $count=1 $X=6.91
+ $Y=0.235 $X2=7.07 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_1%VGND 1 2 3 4 15 19 21 22 28 30 35 40 53
+ 54 58 64 67
r108 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r109 64 65 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r110 58 61 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.36
r111 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r112 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r113 51 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r114 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r115 48 51 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=6.21 $Y2=0
r116 48 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=4.37
+ $Y2=0
r117 47 50 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.83 $Y=0 $X2=6.21
+ $Y2=0
r118 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r119 45 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.615 $Y=0 $X2=4.45
+ $Y2=0
r120 45 47 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.615 $Y=0
+ $X2=4.83 $Y2=0
r121 44 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r122 44 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=2.99
+ $Y2=0
r123 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r124 41 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0 $X2=2.995
+ $Y2=0
r125 41 43 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.08 $Y=0 $X2=3.91
+ $Y2=0
r126 40 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.285 $Y=0 $X2=4.45
+ $Y2=0
r127 40 43 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.285 $Y=0
+ $X2=3.91 $Y2=0
r128 39 65 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.99 $Y2=0
r129 39 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r130 38 39 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r131 36 58 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r132 36 38 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r133 35 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.91 $Y=0 $X2=2.995
+ $Y2=0
r134 35 38 114.824 $w=1.68e-07 $l=1.76e-06 $layer=LI1_cond $X=2.91 $Y=0 $X2=1.15
+ $Y2=0
r135 30 58 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r136 30 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r137 28 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r138 28 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r139 24 53 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=6.685 $Y=0
+ $X2=7.13 $Y2=0
r140 22 50 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.325 $Y=0
+ $X2=6.21 $Y2=0
r141 21 26 11.5244 $w=3.58e-07 $l=3.6e-07 $layer=LI1_cond $X=6.505 $Y=0
+ $X2=6.505 $Y2=0.36
r142 21 24 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=6.505 $Y=0 $X2=6.685
+ $Y2=0
r143 21 22 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=6.505 $Y=0 $X2=6.325
+ $Y2=0
r144 17 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.45 $Y=0.085
+ $X2=4.45 $Y2=0
r145 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.45 $Y=0.085
+ $X2=4.45 $Y2=0.36
r146 13 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=0.085
+ $X2=2.995 $Y2=0
r147 13 15 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.995 $Y=0.085
+ $X2=2.995 $Y2=0.51
r148 4 26 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=6.385
+ $Y=0.235 $X2=6.52 $Y2=0.36
r149 3 19 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=4.265
+ $Y=0.235 $X2=4.45 $Y2=0.36
r150 2 15 182 $w=1.7e-07 $l=3.85357e-07 $layer=licon1_NDIFF $count=1 $X=2.73
+ $Y=0.235 $X2=2.995 $Y2=0.51
r151 1 61 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.36
.ends

