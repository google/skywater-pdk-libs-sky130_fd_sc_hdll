* File: sky130_fd_sc_hdll__a32oi_1.pex.spice
* Created: Thu Aug 27 18:56:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A32OI_1%B2 1 3 4 6 7 12
c26 1 0 1.7339e-19 $X=0.495 $Y=1.41
r27 12 13 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r28 10 12 33.7665 $w=3.64e-07 $l=2.55e-07 $layer=POLY_cond $X=0.24 $Y=1.202
+ $X2=0.495 $Y2=1.202
r29 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r30 4 13 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r31 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r32 1 12 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r33 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_1%B1 1 3 4 6 7 11
c32 11 0 1.7339e-19 $X=1.03 $Y=1.16
r33 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.03
+ $Y=1.16 $X2=1.03 $Y2=1.16
r34 7 11 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.09 $Y=1.53 $X2=1.09
+ $Y2=1.16
r35 4 10 49.2447 $w=2.79e-07 $l=2.73861e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=1.015 $Y2=1.16
r36 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r37 1 10 38.7444 $w=2.79e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=1.015 $Y2=1.16
r38 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995 $X2=0.94
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_1%A1 1 3 4 6 7
r32 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.56
+ $Y=1.16 $X2=1.56 $Y2=1.16
r33 7 11 34.0495 $w=2.18e-07 $l=6.5e-07 $layer=LI1_cond $X=1.585 $Y=0.51
+ $X2=1.585 $Y2=1.16
r34 4 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.62 $Y=0.995
+ $X2=1.56 $Y2=1.16
r35 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.62 $Y=0.995 $X2=1.62
+ $Y2=0.56
r36 1 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.595 $Y=1.41
+ $X2=1.56 $Y2=1.16
r37 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.595 $Y=1.41
+ $X2=1.595 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_1%A2 1 3 4 6 7 8 9
r31 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.1 $Y=1.16
+ $X2=2.1 $Y2=1.16
r32 8 9 17.1909 $w=1.98e-07 $l=3.1e-07 $layer=LI1_cond $X=2.085 $Y=0.85
+ $X2=2.085 $Y2=1.16
r33 7 8 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=2.085 $Y=0.51
+ $X2=2.085 $Y2=0.85
r34 4 14 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.065 $Y=1.41
+ $X2=2.1 $Y2=1.16
r35 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.065 $Y=1.41
+ $X2=2.065 $Y2=1.985
r36 1 14 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.04 $Y=0.995
+ $X2=2.1 $Y2=1.16
r37 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.04 $Y=0.995 $X2=2.04
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_1%A3 3 6 7 8 10 11 14
r23 11 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.58
+ $Y=1.16 $X2=2.58 $Y2=1.16
r24 9 14 25.55 $w=2.7e-07 $l=1.15e-07 $layer=POLY_cond $X=2.58 $Y=1.275 $X2=2.58
+ $Y2=1.16
r25 9 10 35.4596 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.58 $Y=1.275
+ $X2=2.58 $Y2=1.41
r26 7 14 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=2.58 $Y=1.095
+ $X2=2.58 $Y2=1.16
r27 7 8 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.58 $Y=1.095
+ $X2=2.58 $Y2=0.96
r28 6 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.545 $Y=1.985
+ $X2=2.545 $Y2=1.41
r29 3 8 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.52 $Y=0.56 $X2=2.52
+ $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_1%A_27_297# 1 2 3 10 12 14 16 17 18 29
r38 19 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.445 $Y=1.87
+ $X2=1.32 $Y2=1.87
r39 18 29 3.40825 $w=1.7e-07 $l=9.44722e-08 $layer=LI1_cond $X=2.215 $Y=1.87
+ $X2=2.3 $Y2=1.85
r40 18 19 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.215 $Y=1.87
+ $X2=1.445 $Y2=1.87
r41 17 27 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.32 $Y=2.255
+ $X2=1.32 $Y2=2.36
r42 16 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.32 $Y=1.955
+ $X2=1.32 $Y2=1.87
r43 16 17 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=1.32 $Y=1.955 $X2=1.32
+ $Y2=2.255
r44 15 23 3.8266 $w=2.1e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=2.36
+ $X2=0.215 $Y2=2.36
r45 14 27 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.195 $Y=2.36
+ $X2=1.32 $Y2=2.36
r46 14 15 44.8918 $w=2.08e-07 $l=8.5e-07 $layer=LI1_cond $X=1.195 $Y=2.36
+ $X2=0.345 $Y2=2.36
r47 10 23 3.09071 $w=2.6e-07 $l=1.05e-07 $layer=LI1_cond $X=0.215 $Y=2.255
+ $X2=0.215 $Y2=2.36
r48 10 12 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.215 $Y=2.255
+ $X2=0.215 $Y2=2
r49 3 29 300 $w=1.7e-07 $l=4.92189e-07 $layer=licon1_PDIFF $count=2 $X=2.155
+ $Y=1.485 $X2=2.3 $Y2=1.91
r50 2 27 600 $w=1.7e-07 $l=9.55406e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.36 $Y2=2.3
r51 2 25 600 $w=1.7e-07 $l=5.15412e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.36 $Y2=1.87
r52 1 23 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r53 1 12 600 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_1%Y 1 2 7 8 11 14 22
r36 19 22 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=0.645 $Y=1.935
+ $X2=0.68 $Y2=1.935
r37 14 22 1.92074 $w=2.98e-07 $l=5e-08 $layer=LI1_cond $X=0.73 $Y=1.935 $X2=0.68
+ $Y2=1.935
r38 14 19 1.57516 $w=2.6e-07 $l=1.5e-07 $layer=LI1_cond $X=0.645 $Y=1.785
+ $X2=0.645 $Y2=1.935
r39 13 14 30.2423 $w=3.88e-07 $l=9.8e-07 $layer=LI1_cond $X=0.645 $Y=0.805
+ $X2=0.645 $Y2=1.785
r40 9 11 4.03355 $w=2.98e-07 $l=1.05e-07 $layer=LI1_cond $X=1.115 $Y=0.635
+ $X2=1.115 $Y2=0.53
r41 8 13 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.775 $Y=0.72
+ $X2=0.645 $Y2=0.805
r42 7 9 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=0.965 $Y=0.72
+ $X2=1.115 $Y2=0.635
r43 7 8 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.965 $Y=0.72
+ $X2=0.775 $Y2=0.72
r44 2 14 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2
r45 1 11 182 $w=1.7e-07 $l=3.68375e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.18 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_1%VPWR 1 2 9 13 18 19 20 21 22 23 37
r40 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r41 34 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r42 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r43 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r44 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r45 26 30 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r46 23 31 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r47 23 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r48 21 33 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.555 $Y=2.72
+ $X2=2.53 $Y2=2.72
r49 21 22 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.555 $Y=2.72
+ $X2=2.75 $Y2=2.72
r50 20 36 3.22941 $w=1.7e-07 $l=4.5e-08 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=2.99 $Y2=2.72
r51 20 22 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=2.75 $Y2=2.72
r52 18 30 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.705 $Y=2.72
+ $X2=1.61 $Y2=2.72
r53 18 19 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.705 $Y=2.72
+ $X2=1.83 $Y2=2.72
r54 17 33 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.53 $Y2=2.72
r55 17 19 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.83 $Y2=2.72
r56 13 16 20.0939 $w=3.88e-07 $l=6.8e-07 $layer=LI1_cond $X=2.75 $Y=1.66
+ $X2=2.75 $Y2=2.34
r57 11 22 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.75 $Y=2.635
+ $X2=2.75 $Y2=2.72
r58 11 16 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=2.75 $Y=2.635
+ $X2=2.75 $Y2=2.34
r59 7 19 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.83 $Y=2.635
+ $X2=1.83 $Y2=2.72
r60 7 9 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.83 $Y=2.635
+ $X2=1.83 $Y2=2.3
r61 2 16 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=1.485 $X2=2.78 $Y2=2.34
r62 2 13 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=1.485 $X2=2.78 $Y2=1.66
r63 1 9 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.685
+ $Y=1.485 $X2=1.83 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_1%VGND 1 2 7 9 13 15 16 17 18 29
r39 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r40 26 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r41 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r42 23 26 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r43 22 25 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r44 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r45 20 31 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.22
+ $Y2=0
r46 20 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.69
+ $Y2=0
r47 18 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r48 18 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r49 16 25 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.57 $Y=0 $X2=2.53
+ $Y2=0
r50 16 17 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.57 $Y=0 $X2=2.765
+ $Y2=0
r51 15 28 2.15294 $w=1.7e-07 $l=3e-08 $layer=LI1_cond $X=2.96 $Y=0 $X2=2.99
+ $Y2=0
r52 15 17 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.96 $Y=0 $X2=2.765
+ $Y2=0
r53 11 17 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.765 $Y=0.085
+ $X2=2.765 $Y2=0
r54 11 13 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=2.765 $Y=0.085
+ $X2=2.765 $Y2=0.38
r55 7 31 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.22 $Y2=0
r56 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.38
r57 2 13 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=2.595
+ $Y=0.235 $X2=2.78 $Y2=0.38
r58 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.275 $Y2=0.38
.ends

