* File: sky130_fd_sc_hdll__or2_4.pxi.spice
* Created: Thu Aug 27 19:23:22 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR2_4%B N_B_c_57_n N_B_M1009_g N_B_c_60_n N_B_M1003_g B
+ B N_B_c_59_n PM_SKY130_FD_SC_HDLL__OR2_4%B
x_PM_SKY130_FD_SC_HDLL__OR2_4%A N_A_c_86_n N_A_M1004_g N_A_c_87_n N_A_M1001_g A
+ A PM_SKY130_FD_SC_HDLL__OR2_4%A
x_PM_SKY130_FD_SC_HDLL__OR2_4%A_35_297# N_A_35_297#_M1009_d N_A_35_297#_M1003_s
+ N_A_35_297#_c_117_n N_A_35_297#_M1000_g N_A_35_297#_c_123_n
+ N_A_35_297#_M1002_g N_A_35_297#_c_118_n N_A_35_297#_M1005_g
+ N_A_35_297#_c_124_n N_A_35_297#_M1006_g N_A_35_297#_c_119_n
+ N_A_35_297#_M1007_g N_A_35_297#_c_125_n N_A_35_297#_M1010_g
+ N_A_35_297#_c_126_n N_A_35_297#_M1011_g N_A_35_297#_c_120_n
+ N_A_35_297#_M1008_g N_A_35_297#_c_127_n N_A_35_297#_c_121_n
+ N_A_35_297#_c_147_n N_A_35_297#_c_149_n N_A_35_297#_c_129_n
+ N_A_35_297#_c_180_p N_A_35_297#_c_130_n N_A_35_297#_c_139_n
+ N_A_35_297#_c_122_n PM_SKY130_FD_SC_HDLL__OR2_4%A_35_297#
x_PM_SKY130_FD_SC_HDLL__OR2_4%VPWR N_VPWR_M1001_d N_VPWR_M1006_s N_VPWR_M1011_s
+ N_VPWR_c_236_n N_VPWR_c_237_n N_VPWR_c_238_n N_VPWR_c_239_n N_VPWR_c_240_n
+ N_VPWR_c_241_n N_VPWR_c_242_n N_VPWR_c_243_n N_VPWR_c_244_n VPWR
+ N_VPWR_c_245_n N_VPWR_c_235_n PM_SKY130_FD_SC_HDLL__OR2_4%VPWR
x_PM_SKY130_FD_SC_HDLL__OR2_4%X N_X_M1000_s N_X_M1007_s N_X_M1002_d N_X_M1010_d
+ N_X_c_295_n N_X_c_289_n N_X_c_290_n N_X_c_306_n N_X_c_310_n N_X_c_311_n
+ N_X_c_314_n N_X_c_291_n X X PM_SKY130_FD_SC_HDLL__OR2_4%X
x_PM_SKY130_FD_SC_HDLL__OR2_4%VGND N_VGND_M1009_s N_VGND_M1004_d N_VGND_M1005_d
+ N_VGND_M1008_d N_VGND_c_366_n N_VGND_c_367_n N_VGND_c_368_n N_VGND_c_369_n
+ N_VGND_c_370_n N_VGND_c_371_n N_VGND_c_372_n N_VGND_c_373_n N_VGND_c_374_n
+ N_VGND_c_375_n N_VGND_c_376_n VGND N_VGND_c_377_n N_VGND_c_378_n
+ PM_SKY130_FD_SC_HDLL__OR2_4%VGND
cc_1 VNB N_B_c_57_n 0.0187851f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB B 0.0206963f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_B_c_59_n 0.0425581f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_4 VNB N_A_c_86_n 0.0176117f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_5 VNB N_A_c_87_n 0.0273798f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.41
cc_6 VNB A 0.00390991f $X=-0.19 $Y=-0.24 $X2=0.217 $Y2=0.85
cc_7 VNB N_A_35_297#_c_117_n 0.0178713f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_8 VNB N_A_35_297#_c_118_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_9 VNB N_A_35_297#_c_119_n 0.0171643f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_35_297#_c_120_n 0.0203186f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_35_297#_c_121_n 0.00289902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_35_297#_c_122_n 0.0783018f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VPWR_c_235_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_X_c_289_n 0.00264486f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_X_c_290_n 0.00256943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_X_c_291_n 0.0039559f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB X 0.016601f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_366_n 0.0100926f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_19 VNB N_VGND_c_367_n 0.0185223f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.202
cc_20 VNB N_VGND_c_368_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_369_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_370_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_371_n 0.0225503f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_372_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_373_n 0.021597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_374_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_375_n 0.0195326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_376_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_377_n 0.0158267f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_378_n 0.211191f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VPB N_B_c_60_n 0.0202918f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.41
cc_32 VPB B 0.00503328f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_33 VPB N_B_c_59_n 0.0181807f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_34 VPB N_A_c_87_n 0.0264022f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.41
cc_35 VPB A 0.00155242f $X=-0.19 $Y=1.305 $X2=0.217 $Y2=0.85
cc_36 VPB N_A_35_297#_c_123_n 0.0167342f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_35_297#_c_124_n 0.0162421f $X=-0.19 $Y=1.305 $X2=0.217 $Y2=0.85
cc_38 VPB N_A_35_297#_c_125_n 0.0162497f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_35_297#_c_126_n 0.0192858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_35_297#_c_127_n 0.0307964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_35_297#_c_121_n 0.00167261f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_35_297#_c_129_n 0.00157469f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_35_297#_c_130_n 0.00716461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_35_297#_c_122_n 0.0495328f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_236_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_46 VPB N_VPWR_c_237_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.217 $Y2=0.85
cc_47 VPB N_VPWR_c_238_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_239_n 0.035553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_240_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_241_n 0.0212608f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_242_n 0.00323937f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_243_n 0.0197985f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_244_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_245_n 0.0158267f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_235_n 0.0574578f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB X 0.00854525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 N_B_c_57_n N_A_c_86_n 0.0114141f $X=0.52 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_58 N_B_c_60_n N_A_c_87_n 0.0673708f $X=0.555 $Y=1.41 $X2=0 $Y2=0
cc_59 N_B_c_59_n N_A_c_87_n 0.025578f $X=0.52 $Y=1.202 $X2=0 $Y2=0
cc_60 N_B_c_59_n A 3.13535e-19 $X=0.52 $Y=1.202 $X2=0 $Y2=0
cc_61 N_B_c_60_n N_A_35_297#_c_127_n 0.0172825f $X=0.555 $Y=1.41 $X2=0 $Y2=0
cc_62 N_B_c_57_n N_A_35_297#_c_121_n 0.00319101f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_63 N_B_c_60_n N_A_35_297#_c_121_n 0.00460399f $X=0.555 $Y=1.41 $X2=0 $Y2=0
cc_64 N_B_c_59_n N_A_35_297#_c_121_n 0.0165783f $X=0.52 $Y=1.202 $X2=0 $Y2=0
cc_65 N_B_c_60_n N_A_35_297#_c_130_n 0.0137741f $X=0.555 $Y=1.41 $X2=0 $Y2=0
cc_66 B N_A_35_297#_c_130_n 0.0163216f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_67 N_B_c_59_n N_A_35_297#_c_130_n 0.00533125f $X=0.52 $Y=1.202 $X2=0 $Y2=0
cc_68 N_B_c_57_n N_A_35_297#_c_139_n 0.0142588f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_69 B N_A_35_297#_c_139_n 0.0409157f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_70 N_B_c_60_n N_VPWR_c_239_n 0.00628074f $X=0.555 $Y=1.41 $X2=0 $Y2=0
cc_71 N_B_c_60_n N_VPWR_c_235_n 0.0117413f $X=0.555 $Y=1.41 $X2=0 $Y2=0
cc_72 B N_VGND_M1009_s 0.00380678f $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_73 B N_VGND_c_366_n 2.18612e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_74 N_B_c_57_n N_VGND_c_367_n 0.00600179f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_75 B N_VGND_c_367_n 0.0205967f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_76 N_B_c_59_n N_VGND_c_367_n 0.00102593f $X=0.52 $Y=1.202 $X2=0 $Y2=0
cc_77 N_B_c_57_n N_VGND_c_371_n 0.0046926f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_78 N_B_c_57_n N_VGND_c_378_n 0.00880731f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_79 B N_VGND_c_378_n 0.0013663f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_80 N_A_c_86_n N_A_35_297#_c_117_n 0.0175599f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A_c_87_n N_A_35_297#_c_123_n 0.0184999f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A_c_87_n N_A_35_297#_c_127_n 0.00278317f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A_c_86_n N_A_35_297#_c_121_n 0.00763597f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_84 N_A_c_87_n N_A_35_297#_c_121_n 0.00189596f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_85 A N_A_35_297#_c_121_n 0.0258394f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_86 N_A_c_87_n N_A_35_297#_c_147_n 0.020895f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_87 A N_A_35_297#_c_147_n 0.0296092f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_88 A N_A_35_297#_c_149_n 0.0146115f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_89 N_A_c_87_n N_A_35_297#_c_129_n 9.39515e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_90 A N_A_35_297#_c_129_n 0.0062586f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_91 N_A_c_86_n N_A_35_297#_c_139_n 0.00796059f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_92 N_A_c_87_n N_A_35_297#_c_122_n 0.0215331f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_93 A N_A_35_297#_c_122_n 0.00428159f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_94 N_A_c_87_n N_VPWR_c_236_n 0.00780108f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A_c_87_n N_VPWR_c_239_n 0.00702461f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A_c_87_n N_VPWR_c_235_n 0.0127674f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A_c_86_n N_VGND_c_368_n 0.00801937f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_98 N_A_c_87_n N_VGND_c_368_n 5.59096e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_99 A N_VGND_c_368_n 0.0144654f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_100 N_A_c_86_n N_VGND_c_371_n 0.00542757f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A_c_86_n N_VGND_c_378_n 0.0100653f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A_35_297#_c_147_n A_129_297# 0.00418862f $X=1.51 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_103 N_A_35_297#_c_130_n A_129_297# 0.00189464f $X=0.32 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_104 N_A_35_297#_c_147_n N_VPWR_M1001_d 0.00898896f $X=1.51 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_105 N_A_35_297#_c_123_n N_VPWR_c_236_n 0.00525051f $X=1.52 $Y=1.41 $X2=0
+ $Y2=0
cc_106 N_A_35_297#_c_127_n N_VPWR_c_236_n 0.0161967f $X=0.32 $Y=2.3 $X2=0 $Y2=0
cc_107 N_A_35_297#_c_147_n N_VPWR_c_236_n 0.0136682f $X=1.51 $Y=1.58 $X2=0 $Y2=0
cc_108 N_A_35_297#_c_124_n N_VPWR_c_237_n 0.00381622f $X=1.99 $Y=1.41 $X2=0
+ $Y2=0
cc_109 N_A_35_297#_c_125_n N_VPWR_c_237_n 0.00402622f $X=2.46 $Y=1.41 $X2=0
+ $Y2=0
cc_110 N_A_35_297#_c_126_n N_VPWR_c_238_n 0.0064303f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A_35_297#_c_127_n N_VPWR_c_239_n 0.0230775f $X=0.32 $Y=2.3 $X2=0 $Y2=0
cc_112 N_A_35_297#_c_123_n N_VPWR_c_241_n 0.00673617f $X=1.52 $Y=1.41 $X2=0
+ $Y2=0
cc_113 N_A_35_297#_c_124_n N_VPWR_c_241_n 0.0048852f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_35_297#_c_125_n N_VPWR_c_243_n 0.00514793f $X=2.46 $Y=1.41 $X2=0
+ $Y2=0
cc_115 N_A_35_297#_c_126_n N_VPWR_c_243_n 0.00597712f $X=2.93 $Y=1.41 $X2=0
+ $Y2=0
cc_116 N_A_35_297#_M1003_s N_VPWR_c_235_n 0.00233913f $X=0.175 $Y=1.485 $X2=0
+ $Y2=0
cc_117 N_A_35_297#_c_123_n N_VPWR_c_235_n 0.012155f $X=1.52 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A_35_297#_c_124_n N_VPWR_c_235_n 0.00650546f $X=1.99 $Y=1.41 $X2=0
+ $Y2=0
cc_119 N_A_35_297#_c_125_n N_VPWR_c_235_n 0.00677533f $X=2.46 $Y=1.41 $X2=0
+ $Y2=0
cc_120 N_A_35_297#_c_126_n N_VPWR_c_235_n 0.0110717f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_35_297#_c_127_n N_VPWR_c_235_n 0.0134907f $X=0.32 $Y=2.3 $X2=0 $Y2=0
cc_122 N_A_35_297#_c_147_n N_X_M1002_d 0.00334924f $X=1.51 $Y=1.58 $X2=0 $Y2=0
cc_123 N_A_35_297#_c_118_n N_X_c_295_n 0.00854453f $X=1.965 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A_35_297#_c_119_n N_X_c_295_n 5.82315e-19 $X=2.435 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_35_297#_c_118_n N_X_c_289_n 0.0060427f $X=1.965 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_35_297#_c_119_n N_X_c_289_n 0.0107277f $X=2.435 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_35_297#_c_180_p N_X_c_289_n 0.0455988f $X=2.455 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_35_297#_c_122_n N_X_c_289_n 0.00345061f $X=2.93 $Y=1.202 $X2=0 $Y2=0
cc_129 N_A_35_297#_c_117_n N_X_c_290_n 6.43527e-19 $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_35_297#_c_118_n N_X_c_290_n 0.00262358f $X=1.965 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_35_297#_c_149_n N_X_c_290_n 0.0153702f $X=1.637 $Y=1.245 $X2=0 $Y2=0
cc_132 N_A_35_297#_c_180_p N_X_c_290_n 0.0160635f $X=2.455 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_35_297#_c_122_n N_X_c_290_n 0.00357932f $X=2.93 $Y=1.202 $X2=0 $Y2=0
cc_134 N_A_35_297#_c_124_n N_X_c_306_n 0.00947543f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_35_297#_c_125_n N_X_c_306_n 0.0128736f $X=2.46 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A_35_297#_c_180_p N_X_c_306_n 0.0125645f $X=2.455 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_35_297#_c_122_n N_X_c_306_n 0.00481395f $X=2.93 $Y=1.202 $X2=0 $Y2=0
cc_138 N_A_35_297#_c_120_n N_X_c_310_n 0.0111926f $X=2.955 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_35_297#_c_124_n N_X_c_311_n 5.16456e-19 $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_35_297#_c_125_n N_X_c_311_n 0.00665381f $X=2.46 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_35_297#_c_126_n N_X_c_311_n 0.00723796f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_35_297#_c_123_n N_X_c_314_n 0.00846409f $X=1.52 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_35_297#_c_124_n N_X_c_314_n 0.011379f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_35_297#_c_125_n N_X_c_314_n 5.5123e-19 $X=2.46 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_35_297#_c_147_n N_X_c_314_n 0.0102737f $X=1.51 $Y=1.58 $X2=0 $Y2=0
cc_146 N_A_35_297#_c_180_p N_X_c_314_n 0.00486487f $X=2.455 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_35_297#_c_122_n N_X_c_314_n 0.00288832f $X=2.93 $Y=1.202 $X2=0 $Y2=0
cc_148 N_A_35_297#_c_120_n N_X_c_291_n 0.00924052f $X=2.955 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_35_297#_c_122_n N_X_c_291_n 0.00551758f $X=2.93 $Y=1.202 $X2=0 $Y2=0
cc_150 N_A_35_297#_c_119_n X 0.00186312f $X=2.435 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_35_297#_c_125_n X 0.00156711f $X=2.46 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_35_297#_c_126_n X 0.00310484f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_35_297#_c_120_n X 0.00384363f $X=2.955 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_35_297#_c_180_p X 0.0115725f $X=2.455 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_35_297#_c_122_n X 0.0279195f $X=2.93 $Y=1.202 $X2=0 $Y2=0
cc_156 N_A_35_297#_c_124_n X 0.00157305f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_35_297#_c_125_n X 0.00728727f $X=2.46 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_35_297#_c_126_n X 0.0221888f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_35_297#_c_180_p X 0.00327411f $X=2.455 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_35_297#_c_122_n X 0.00718514f $X=2.93 $Y=1.202 $X2=0 $Y2=0
cc_161 N_A_35_297#_c_139_n N_VGND_c_367_n 0.0233571f $X=0.73 $Y=0.4 $X2=0 $Y2=0
cc_162 N_A_35_297#_c_117_n N_VGND_c_368_n 0.00637569f $X=1.495 $Y=0.995 $X2=0
+ $Y2=0
cc_163 N_A_35_297#_c_139_n N_VGND_c_368_n 0.0283955f $X=0.73 $Y=0.4 $X2=0 $Y2=0
cc_164 N_A_35_297#_c_118_n N_VGND_c_369_n 0.00377869f $X=1.965 $Y=0.995 $X2=0
+ $Y2=0
cc_165 N_A_35_297#_c_119_n N_VGND_c_369_n 0.00276126f $X=2.435 $Y=0.995 $X2=0
+ $Y2=0
cc_166 N_A_35_297#_c_120_n N_VGND_c_370_n 0.00438629f $X=2.955 $Y=0.995 $X2=0
+ $Y2=0
cc_167 N_A_35_297#_c_139_n N_VGND_c_371_n 0.0181506f $X=0.73 $Y=0.4 $X2=0 $Y2=0
cc_168 N_A_35_297#_c_117_n N_VGND_c_373_n 0.00585385f $X=1.495 $Y=0.995 $X2=0
+ $Y2=0
cc_169 N_A_35_297#_c_118_n N_VGND_c_373_n 0.00398337f $X=1.965 $Y=0.995 $X2=0
+ $Y2=0
cc_170 N_A_35_297#_c_119_n N_VGND_c_375_n 0.00439206f $X=2.435 $Y=0.995 $X2=0
+ $Y2=0
cc_171 N_A_35_297#_c_120_n N_VGND_c_375_n 0.00423846f $X=2.955 $Y=0.995 $X2=0
+ $Y2=0
cc_172 N_A_35_297#_M1009_d N_VGND_c_378_n 0.00217091f $X=0.595 $Y=0.235 $X2=0
+ $Y2=0
cc_173 N_A_35_297#_c_117_n N_VGND_c_378_n 0.0111758f $X=1.495 $Y=0.995 $X2=0
+ $Y2=0
cc_174 N_A_35_297#_c_118_n N_VGND_c_378_n 0.0058274f $X=1.965 $Y=0.995 $X2=0
+ $Y2=0
cc_175 N_A_35_297#_c_119_n N_VGND_c_378_n 0.00628058f $X=2.435 $Y=0.995 $X2=0
+ $Y2=0
cc_176 N_A_35_297#_c_120_n N_VGND_c_378_n 0.00711863f $X=2.955 $Y=0.995 $X2=0
+ $Y2=0
cc_177 N_A_35_297#_c_139_n N_VGND_c_378_n 0.0136221f $X=0.73 $Y=0.4 $X2=0 $Y2=0
cc_178 A_129_297# N_VPWR_c_235_n 0.00983149f $X=0.645 $Y=1.485 $X2=0.705 $Y2=0.4
cc_179 N_VPWR_c_235_n N_X_M1002_d 0.00231261f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_180 N_VPWR_c_235_n N_X_M1010_d 0.00231261f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_181 N_VPWR_M1006_s N_X_c_306_n 0.00463882f $X=2.08 $Y=1.485 $X2=0 $Y2=0
cc_182 N_VPWR_c_237_n N_X_c_306_n 0.0131159f $X=2.225 $Y=2.34 $X2=0 $Y2=0
cc_183 N_VPWR_c_241_n N_X_c_306_n 0.00198891f $X=2.14 $Y=2.72 $X2=0 $Y2=0
cc_184 N_VPWR_c_243_n N_X_c_306_n 0.00267292f $X=3.08 $Y=2.72 $X2=0 $Y2=0
cc_185 N_VPWR_c_235_n N_X_c_306_n 0.00968081f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_186 N_VPWR_c_237_n N_X_c_311_n 0.0177504f $X=2.225 $Y=2.34 $X2=0 $Y2=0
cc_187 N_VPWR_c_238_n N_X_c_311_n 0.034303f $X=3.165 $Y=2 $X2=0 $Y2=0
cc_188 N_VPWR_c_243_n N_X_c_311_n 0.0223557f $X=3.08 $Y=2.72 $X2=0 $Y2=0
cc_189 N_VPWR_c_235_n N_X_c_311_n 0.0139997f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_190 N_VPWR_c_236_n N_X_c_314_n 0.0343633f $X=1.245 $Y=2.01 $X2=0 $Y2=0
cc_191 N_VPWR_c_237_n N_X_c_314_n 0.02165f $X=2.225 $Y=2.34 $X2=0 $Y2=0
cc_192 N_VPWR_c_241_n N_X_c_314_n 0.0222542f $X=2.14 $Y=2.72 $X2=0 $Y2=0
cc_193 N_VPWR_c_235_n N_X_c_314_n 0.0139813f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_194 N_VPWR_M1011_s X 3.74046e-19 $X=3.02 $Y=1.485 $X2=0 $Y2=0
cc_195 N_VPWR_M1011_s X 0.00858714f $X=3.02 $Y=1.485 $X2=0 $Y2=0
cc_196 N_VPWR_c_238_n X 0.021341f $X=3.165 $Y=2 $X2=0 $Y2=0
cc_197 N_X_c_289_n N_VGND_M1005_d 0.00251598f $X=2.53 $Y=0.82 $X2=0 $Y2=0
cc_198 N_X_c_291_n N_VGND_M1008_d 0.00758342f $X=2.997 $Y=0.905 $X2=0 $Y2=0
cc_199 N_X_c_295_n N_VGND_c_369_n 0.0223967f $X=1.755 $Y=0.4 $X2=0 $Y2=0
cc_200 N_X_c_289_n N_VGND_c_369_n 0.0127122f $X=2.53 $Y=0.82 $X2=0 $Y2=0
cc_201 N_X_c_291_n N_VGND_c_370_n 0.00651305f $X=2.997 $Y=0.905 $X2=0 $Y2=0
cc_202 N_X_c_295_n N_VGND_c_373_n 0.0216696f $X=1.755 $Y=0.4 $X2=0 $Y2=0
cc_203 N_X_c_289_n N_VGND_c_373_n 0.00194552f $X=2.53 $Y=0.82 $X2=0 $Y2=0
cc_204 N_X_c_289_n N_VGND_c_375_n 0.00444586f $X=2.53 $Y=0.82 $X2=0 $Y2=0
cc_205 N_X_c_310_n N_VGND_c_375_n 0.0213655f $X=2.695 $Y=0.4 $X2=0 $Y2=0
cc_206 N_X_M1000_s N_VGND_c_378_n 0.00325153f $X=1.57 $Y=0.235 $X2=0 $Y2=0
cc_207 N_X_M1007_s N_VGND_c_378_n 0.00306175f $X=2.51 $Y=0.235 $X2=0 $Y2=0
cc_208 N_X_c_295_n N_VGND_c_378_n 0.0140292f $X=1.755 $Y=0.4 $X2=0 $Y2=0
cc_209 N_X_c_289_n N_VGND_c_378_n 0.0135311f $X=2.53 $Y=0.82 $X2=0 $Y2=0
cc_210 N_X_c_310_n N_VGND_c_378_n 0.0141427f $X=2.695 $Y=0.4 $X2=0 $Y2=0
cc_211 N_X_c_291_n N_VGND_c_378_n 3.33075e-19 $X=2.997 $Y=0.905 $X2=0 $Y2=0
