* File: sky130_fd_sc_hdll__sdfstp_1.pex.spice
* Created: Thu Aug 27 19:27:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%SCD 1 2 3 5 6 8 13 14
c33 3 0 3.49297e-20 $X=0.495 $Y=1.77
r34 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.255
+ $Y=1.16 $X2=0.255 $Y2=1.16
r35 14 19 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.212 $Y=1.53
+ $X2=0.212 $Y2=1.16
r36 13 19 14.0101 $w=2.53e-07 $l=3.1e-07 $layer=LI1_cond $X=0.212 $Y=0.85
+ $X2=0.212 $Y2=1.16
r37 6 18 85.0704 $w=2.76e-07 $l=5.07937e-07 $layer=POLY_cond $X=0.52 $Y=0.73
+ $X2=0.35 $Y2=1.16
r38 6 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.445
r39 3 9 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.495 $Y=1.695
+ $X2=0.315 $Y2=1.695
r40 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.77
+ $X2=0.495 $Y2=2.165
r41 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.315 $Y=1.62
+ $X2=0.315 $Y2=1.695
r42 1 18 38.7914 $w=2.76e-07 $l=1.81659e-07 $layer=POLY_cond $X=0.315 $Y=1.325
+ $X2=0.35 $Y2=1.16
r43 1 2 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.315 $Y=1.325
+ $X2=0.315 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%SCE 3 6 7 9 11 12 14 17 19 20 22 25 30 33
+ 34 38 46
c110 30 0 4.39648e-20 $X=0.93 $Y=1.25
c111 22 0 1.07953e-19 $X=2.73 $Y=1.19
c112 7 0 1.40323e-19 $X=0.965 $Y=1.77
r113 33 36 37.7919 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.782 $Y=1.16
+ $X2=2.782 $Y2=1.325
r114 33 35 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.782 $Y=1.16
+ $X2=2.782 $Y2=0.995
r115 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.735
+ $Y=1.16 $X2=2.735 $Y2=1.16
r116 30 31 5.56766 $w=3.03e-07 $l=3.5e-08 $layer=POLY_cond $X=0.93 $Y=1.25
+ $X2=0.965 $Y2=1.25
r117 28 30 23.066 $w=3.03e-07 $l=1.45e-07 $layer=POLY_cond $X=0.785 $Y=1.25
+ $X2=0.93 $Y2=1.25
r118 28 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.785
+ $Y=1.25 $X2=0.785 $Y2=1.25
r119 25 46 0.0320802 $w=2.3e-07 $l=5e-08 $layer=MET1_cond $X=0.69 $Y=1.19
+ $X2=0.64 $Y2=1.19
r120 25 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.725 $Y=1.19
+ $X2=0.725 $Y2=1.19
r121 22 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.73 $Y=1.19
+ $X2=2.73 $Y2=1.19
r122 20 25 0.137923 $w=2.3e-07 $l=1.8e-07 $layer=MET1_cond $X=0.87 $Y=1.19
+ $X2=0.69 $Y2=1.19
r123 19 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.585 $Y=1.19
+ $X2=2.73 $Y2=1.19
r124 19 20 2.12252 $w=1.4e-07 $l=1.715e-06 $layer=MET1_cond $X=2.585 $Y=1.19
+ $X2=0.87 $Y2=1.19
r125 17 35 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.89 $Y=0.445
+ $X2=2.89 $Y2=0.995
r126 12 14 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.835 $Y=1.77
+ $X2=2.835 $Y2=2.165
r127 11 12 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.835 $Y=1.67 $X2=2.835
+ $Y2=1.77
r128 11 36 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=2.835 $Y=1.67
+ $X2=2.835 $Y2=1.325
r129 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.965 $Y=1.77
+ $X2=0.965 $Y2=2.165
r130 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.67 $X2=0.965
+ $Y2=1.77
r131 5 31 12.5184 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.415
+ $X2=0.965 $Y2=1.25
r132 5 6 84.5522 $w=2e-07 $l=2.55e-07 $layer=POLY_cond $X=0.965 $Y=1.415
+ $X2=0.965 $Y2=1.67
r133 1 30 19.2026 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.085
+ $X2=0.93 $Y2=1.25
r134 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.93 $Y=1.085 $X2=0.93
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%D 2 3 5 8 9 10 14 16
c49 9 0 3.49297e-20 $X=1.15 $Y=0.85
r50 14 16 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=0.93
+ $X2=1.375 $Y2=0.765
r51 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.35
+ $Y=0.93 $X2=1.35 $Y2=0.93
r52 10 15 15.5386 $w=4.43e-07 $l=6e-07 $layer=LI1_cond $X=1.262 $Y=1.53
+ $X2=1.262 $Y2=0.93
r53 9 15 2.07181 $w=4.43e-07 $l=8e-08 $layer=LI1_cond $X=1.262 $Y=0.85 $X2=1.262
+ $Y2=0.93
r54 8 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.4 $Y=0.445 $X2=1.4
+ $Y2=0.765
r55 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.375 $Y=1.77
+ $X2=1.375 $Y2=2.165
r56 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.375 $Y=1.67 $X2=1.375
+ $Y2=1.77
r57 1 14 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.095
+ $X2=1.375 $Y2=0.93
r58 1 2 190.657 $w=2e-07 $l=5.75e-07 $layer=POLY_cond $X=1.375 $Y=1.095
+ $X2=1.375 $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_349_21# 1 2 9 12 13 15 17 21 22 23 25
+ 35 37
c79 22 0 1.4475e-19 $X=2.15 $Y=1.16
r80 35 37 0.182927 $w=3.13e-07 $l=5e-09 $layer=LI1_cond $X=2.595 $Y=1.927
+ $X2=2.6 $Y2=1.927
r81 23 25 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=2.59 $Y=0.715
+ $X2=2.59 $Y2=0.44
r82 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=1.16 $X2=2.15 $Y2=1.16
r83 19 35 13.2805 $w=3.13e-07 $l=3.63e-07 $layer=LI1_cond $X=2.232 $Y=1.927
+ $X2=2.595 $Y2=1.927
r84 19 21 20.9848 $w=3.33e-07 $l=6.1e-07 $layer=LI1_cond $X=2.232 $Y=1.77
+ $X2=2.232 $Y2=1.16
r85 18 23 20.8976 $w=1.88e-07 $l=3.58e-07 $layer=LI1_cond $X=2.232 $Y=0.81
+ $X2=2.59 $Y2=0.81
r86 18 21 8.77233 $w=3.33e-07 $l=2.55e-07 $layer=LI1_cond $X=2.232 $Y=0.905
+ $X2=2.232 $Y2=1.16
r87 16 22 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.945 $Y=1.16
+ $X2=2.15 $Y2=1.16
r88 16 17 3.18546 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=1.945 $Y=1.16
+ $X2=1.845 $Y2=1.16
r89 13 15 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.845 $Y=1.77
+ $X2=1.845 $Y2=2.165
r90 12 13 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.845 $Y=1.67 $X2=1.845
+ $Y2=1.77
r91 11 17 33.332 $w=1.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.325
+ $X2=1.845 $Y2=1.16
r92 11 12 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=1.845 $Y=1.325
+ $X2=1.845 $Y2=1.67
r93 7 17 33.332 $w=1.75e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.82 $Y=0.995
+ $X2=1.845 $Y2=1.16
r94 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.82 $Y=0.995 $X2=1.82
+ $Y2=0.445
r95 2 37 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.475
+ $Y=1.845 $X2=2.6 $Y2=1.99
r96 1 25 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=2.505
+ $Y=0.235 $X2=2.63 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%CLK 7 8 10 13 15 16 17 20 21 22
c58 21 0 3.28604e-20 $X=3.68 $Y=1.255
c59 13 0 1.06712e-19 $X=3.88 $Y=0.805
r60 20 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.68 $Y=1.255
+ $X2=3.68 $Y2=1.42
r61 20 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.68 $Y=1.255
+ $X2=3.68 $Y2=1.09
r62 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.68
+ $Y=1.255 $X2=3.68 $Y2=1.255
r63 17 21 4.6235 $w=5.93e-07 $l=2.3e-07 $layer=LI1_cond $X=3.45 $Y=1.352
+ $X2=3.68 $Y2=1.352
r64 15 16 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.795 $Y=1.62
+ $X2=3.795 $Y2=1.77
r65 15 23 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.74 $Y=1.62 $X2=3.74
+ $Y2=1.42
r66 11 13 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=3.74 $Y=0.805
+ $X2=3.88 $Y2=0.805
r67 8 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.88 $Y=0.73 $X2=3.88
+ $Y2=0.805
r68 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.88 $Y=0.73 $X2=3.88
+ $Y2=0.445
r69 7 16 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.825 $Y=2.165
+ $X2=3.825 $Y2=1.77
r70 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.74 $Y=0.88 $X2=3.74
+ $Y2=0.805
r71 1 22 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.74 $Y=0.88 $X2=3.74
+ $Y2=1.09
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_693_369# 1 2 8 9 11 14 16 17 19 21 22
+ 24 26 27 29 32 34 37 41 43 44 45 46 48 50 51 55 56 57 58 61 62 64 65 66 67 68
+ 77 81 85
c289 85 0 1.8066e-19 $X=5.73 $Y=1.74
c290 81 0 3.28604e-20 $X=4.235 $Y=1.09
c291 77 0 3.33234e-19 $X=8.295 $Y=1.87
c292 62 0 5.96508e-20 $X=9.64 $Y=1.09
c293 34 0 6.74919e-20 $X=4.317 $Y=0.805
r294 84 85 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.73
+ $Y=1.74 $X2=5.73 $Y2=1.74
r295 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.295 $Y=1.87
+ $X2=8.295 $Y2=1.87
r296 74 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.69 $Y=1.87
+ $X2=5.69 $Y2=1.87
r297 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.21 $Y=1.87
+ $X2=4.21 $Y2=1.87
r298 68 74 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=5.885 $Y=1.87
+ $X2=5.69 $Y2=1.87
r299 67 77 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.15 $Y=1.87
+ $X2=8.295 $Y2=1.87
r300 67 68 2.80321 $w=1.4e-07 $l=2.265e-06 $layer=MET1_cond $X=8.15 $Y=1.87
+ $X2=5.885 $Y2=1.87
r301 66 70 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=4.405 $Y=1.87
+ $X2=4.21 $Y2=1.87
r302 65 74 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.545 $Y=1.87
+ $X2=5.69 $Y2=1.87
r303 65 66 1.41089 $w=1.4e-07 $l=1.14e-06 $layer=MET1_cond $X=5.545 $Y=1.87
+ $X2=4.405 $Y2=1.87
r304 64 78 8.13333 $w=2.85e-07 $l=1.9e-07 $layer=LI1_cond $X=8.485 $Y=1.812
+ $X2=8.295 $Y2=1.812
r305 62 90 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.64 $Y=1.09
+ $X2=9.64 $Y2=0.925
r306 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.64
+ $Y=1.09 $X2=9.64 $Y2=1.09
r307 59 61 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=9.685 $Y=0.905
+ $X2=9.685 $Y2=1.09
r308 57 59 7.54394 $w=1.85e-07 $l=2.06325e-07 $layer=LI1_cond $X=9.52 $Y=0.812
+ $X2=9.685 $Y2=0.905
r309 57 58 44.0639 $w=1.83e-07 $l=7.35e-07 $layer=LI1_cond $X=9.52 $Y=0.812
+ $X2=8.785 $Y2=0.812
r310 56 88 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.57 $Y=1.16
+ $X2=8.57 $Y2=1.325
r311 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.57
+ $Y=1.16 $X2=8.57 $Y2=1.16
r312 53 64 6.82232 $w=2.85e-07 $l=2.09285e-07 $layer=LI1_cond $X=8.635 $Y=1.67
+ $X2=8.485 $Y2=1.812
r313 53 55 19.5915 $w=2.98e-07 $l=5.1e-07 $layer=LI1_cond $X=8.635 $Y=1.67
+ $X2=8.635 $Y2=1.16
r314 52 58 7.32714 $w=1.85e-07 $l=1.90919e-07 $layer=LI1_cond $X=8.635 $Y=0.905
+ $X2=8.785 $Y2=0.812
r315 52 55 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=8.635 $Y=0.905
+ $X2=8.635 $Y2=1.16
r316 51 82 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.235 $Y=1.255
+ $X2=4.235 $Y2=1.42
r317 51 81 39.9376 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.235 $Y=1.255
+ $X2=4.235 $Y2=1.09
r318 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.21
+ $Y=1.255 $X2=4.21 $Y2=1.255
r319 48 71 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.165 $Y=1.83
+ $X2=4.165 $Y2=1.915
r320 48 50 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=4.165 $Y=1.83
+ $X2=4.165 $Y2=1.255
r321 47 50 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=4.165 $Y=0.885
+ $X2=4.165 $Y2=1.255
r322 45 47 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.035 $Y=0.8
+ $X2=4.165 $Y2=0.885
r323 45 46 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.035 $Y=0.8
+ $X2=3.705 $Y2=0.8
r324 43 71 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.035 $Y=1.915
+ $X2=4.165 $Y2=1.915
r325 43 44 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.035 $Y=1.915
+ $X2=3.675 $Y2=1.915
r326 39 46 6.83233 $w=1.7e-07 $l=1.28662e-07 $layer=LI1_cond $X=3.612 $Y=0.715
+ $X2=3.705 $Y2=0.8
r327 39 41 16.4865 $w=1.83e-07 $l=2.75e-07 $layer=LI1_cond $X=3.612 $Y=0.715
+ $X2=3.612 $Y2=0.44
r328 35 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.59 $Y=2
+ $X2=3.675 $Y2=1.915
r329 35 37 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.59 $Y=2 $X2=3.59
+ $Y2=2.16
r330 32 90 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.7 $Y=0.445
+ $X2=9.7 $Y2=0.925
r331 27 29 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=8.535 $Y=1.57
+ $X2=8.535 $Y2=2.065
r332 26 27 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=8.535 $Y=1.47 $X2=8.535
+ $Y2=1.57
r333 26 88 48.0787 $w=2e-07 $l=1.45e-07 $layer=POLY_cond $X=8.535 $Y=1.47
+ $X2=8.535 $Y2=1.325
r334 22 84 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=5.755 $Y=1.99
+ $X2=5.755 $Y2=1.74
r335 22 24 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.755 $Y=1.99
+ $X2=5.755 $Y2=2.275
r336 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.34 $Y=0.73
+ $X2=5.34 $Y2=0.445
r337 18 34 6.88539 $w=1.5e-07 $l=1.08e-07 $layer=POLY_cond $X=4.425 $Y=0.805
+ $X2=4.317 $Y2=0.805
r338 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.265 $Y=0.805
+ $X2=5.34 $Y2=0.73
r339 17 18 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=5.265 $Y=0.805
+ $X2=4.425 $Y2=0.805
r340 14 34 18.6014 $w=1.67e-07 $l=9e-08 $layer=POLY_cond $X=4.35 $Y=0.73
+ $X2=4.317 $Y2=0.805
r341 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.35 $Y=0.73
+ $X2=4.35 $Y2=0.445
r342 12 34 18.6014 $w=1.67e-07 $l=8.21584e-08 $layer=POLY_cond $X=4.302 $Y=0.88
+ $X2=4.317 $Y2=0.805
r343 12 81 77.5789 $w=1.85e-07 $l=2.1e-07 $layer=POLY_cond $X=4.302 $Y=0.88
+ $X2=4.302 $Y2=1.09
r344 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=4.295 $Y=1.77
+ $X2=4.295 $Y2=2.165
r345 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.295 $Y=1.67 $X2=4.295
+ $Y2=1.77
r346 8 82 82.8943 $w=2e-07 $l=2.5e-07 $layer=POLY_cond $X=4.295 $Y=1.67
+ $X2=4.295 $Y2=1.42
r347 2 37 600 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_PDIFF $count=1 $X=3.465
+ $Y=1.845 $X2=3.59 $Y2=2.16
r348 1 41 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=3.495
+ $Y=0.235 $X2=3.62 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_877_369# 1 2 8 9 11 12 13 15 18 22 24
+ 26 29 34 35 37 39 41 42 46 48 54
c184 46 0 1.33492e-19 $X=4.72 $Y=1.185
c185 42 0 1.03798e-20 $X=9.135 $Y=1.19
c186 39 0 1.24362e-19 $X=9.055 $Y=1.19
c187 29 0 7.95993e-20 $X=4.56 $Y=0.42
c188 24 0 1.39178e-19 $X=9.115 $Y=1.99
c189 18 0 1.00357e-19 $X=5.81 $Y=0.445
c190 11 0 2.89743e-19 $X=5.195 $Y=1.915
c191 9 0 1.70908e-19 $X=5.735 $Y=1.165
c192 8 0 1.8066e-19 $X=4.965 $Y=1.84
r193 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.205
+ $Y=1.74 $X2=9.205 $Y2=1.74
r194 53 54 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.965 $Y=1.255
+ $X2=5.04 $Y2=1.255
r195 50 53 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.755 $Y=1.255
+ $X2=4.965 $Y2=1.255
r196 46 64 7.6678 $w=3.63e-07 $l=2.35e-07 $layer=LI1_cond $X=4.657 $Y=1.185
+ $X2=4.657 $Y2=1.42
r197 46 63 5.21818 $w=3.63e-07 $l=1e-07 $layer=LI1_cond $X=4.657 $Y=1.185
+ $X2=4.657 $Y2=1.085
r198 46 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.755
+ $Y=1.255 $X2=4.755 $Y2=1.255
r199 45 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.72 $Y=1.185
+ $X2=4.865 $Y2=1.185
r200 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.72 $Y=1.185
+ $X2=4.72 $Y2=1.185
r201 42 57 18.9207 $w=3.33e-07 $l=5.5e-07 $layer=LI1_cond $X=9.122 $Y=1.19
+ $X2=9.122 $Y2=1.74
r202 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.135 $Y=1.19
+ $X2=9.135 $Y2=1.19
r203 39 41 0.0513283 $w=2.3e-07 $l=8e-08 $layer=MET1_cond $X=9.055 $Y=1.19
+ $X2=9.135 $Y2=1.19
r204 37 39 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=8.94 $Y=1.19
+ $X2=9.055 $Y2=1.19
r205 37 48 5.04331 $w=1.4e-07 $l=4.075e-06 $layer=MET1_cond $X=8.94 $Y=1.19
+ $X2=4.865 $Y2=1.19
r206 35 64 26.1586 $w=3.13e-07 $l=7.15e-07 $layer=LI1_cond $X=4.632 $Y=2.135
+ $X2=4.632 $Y2=1.42
r207 34 35 5.62076 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=4.617 $Y=2.3
+ $X2=4.617 $Y2=2.135
r208 29 63 35.1212 $w=2.08e-07 $l=6.65e-07 $layer=LI1_cond $X=4.58 $Y=0.42
+ $X2=4.58 $Y2=1.085
r209 24 56 47.8775 $w=2.99e-07 $l=2.79285e-07 $layer=POLY_cond $X=9.115 $Y=1.99
+ $X2=9.177 $Y2=1.74
r210 24 26 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=9.115 $Y=1.99
+ $X2=9.115 $Y2=2.275
r211 20 56 38.5562 $w=2.99e-07 $l=2.03912e-07 $layer=POLY_cond $X=9.09 $Y=1.575
+ $X2=9.177 $Y2=1.74
r212 20 22 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=9.09 $Y=1.575
+ $X2=9.09 $Y2=0.555
r213 16 18 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=5.81 $Y=1.09
+ $X2=5.81 $Y2=0.445
r214 13 15 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.285 $Y=1.99
+ $X2=5.285 $Y2=2.275
r215 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.195 $Y=1.915
+ $X2=5.285 $Y2=1.99
r216 11 12 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=5.195 $Y=1.915
+ $X2=5.04 $Y2=1.915
r217 9 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.735 $Y=1.165
+ $X2=5.81 $Y2=1.09
r218 9 54 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=5.735 $Y=1.165
+ $X2=5.04 $Y2=1.165
r219 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.965 $Y=1.84
+ $X2=5.04 $Y2=1.915
r220 7 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.965 $Y=1.42
+ $X2=4.965 $Y2=1.255
r221 7 8 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=4.965 $Y=1.42
+ $X2=4.965 $Y2=1.84
r222 2 34 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=4.385
+ $Y=1.845 $X2=4.53 $Y2=2.3
r223 1 29 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_1229_21# 1 2 9 12 13 15 18 21 23 24 27
+ 31 33 37
c95 33 0 4.30126e-20 $X=6.285 $Y=0.72
c96 23 0 3.13156e-20 $X=7.155 $Y=2.02
c97 21 0 3.97233e-20 $X=6.785 $Y=0.72
r98 37 41 32.4954 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.31 $Y=0.93
+ $X2=6.31 $Y2=1.065
r99 37 40 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.31 $Y=0.93
+ $X2=6.31 $Y2=0.795
r100 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.31
+ $Y=0.93 $X2=6.31 $Y2=0.93
r101 33 36 6.36876 $w=3.78e-07 $l=2.1e-07 $layer=LI1_cond $X=6.285 $Y=0.72
+ $X2=6.285 $Y2=0.93
r102 29 31 7.82791 $w=2.63e-07 $l=1.8e-07 $layer=LI1_cond $X=7.287 $Y=2.105
+ $X2=7.287 $Y2=2.285
r103 25 27 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.91 $Y=0.635
+ $X2=6.91 $Y2=0.51
r104 23 29 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=7.155 $Y=2.02
+ $X2=7.287 $Y2=2.105
r105 23 24 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.155 $Y=2.02
+ $X2=6.595 $Y2=2.02
r106 22 33 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.475 $Y=0.72
+ $X2=6.285 $Y2=0.72
r107 21 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.785 $Y=0.72
+ $X2=6.91 $Y2=0.635
r108 21 22 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.785 $Y=0.72
+ $X2=6.475 $Y2=0.72
r109 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.51
+ $Y=1.74 $X2=6.51 $Y2=1.74
r110 16 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.51 $Y=1.935
+ $X2=6.595 $Y2=2.02
r111 16 18 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.51 $Y=1.935
+ $X2=6.51 $Y2=1.74
r112 13 19 45.1054 $w=3.82e-07 $l=3.02076e-07 $layer=POLY_cond $X=6.315 $Y=1.99
+ $X2=6.43 $Y2=1.74
r113 13 15 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.315 $Y=1.99
+ $X2=6.315 $Y2=2.275
r114 12 19 31.7097 $w=3.82e-07 $l=2.14942e-07 $layer=POLY_cond $X=6.315 $Y=1.575
+ $X2=6.43 $Y2=1.74
r115 12 41 169.104 $w=2e-07 $l=5.1e-07 $layer=POLY_cond $X=6.315 $Y=1.575
+ $X2=6.315 $Y2=1.065
r116 9 40 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.22 $Y=0.445
+ $X2=6.22 $Y2=0.795
r117 2 31 600 $w=1.7e-07 $l=2.92916e-07 $layer=licon1_PDIFF $count=1 $X=7.095
+ $Y=2.065 $X2=7.265 $Y2=2.285
r118 1 27 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=6.825
+ $Y=0.235 $X2=6.95 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_1075_413# 1 2 8 10 11 13 14 16 18 19 21
+ 24 27 29 35 38 40 49 50 52 53 54 58 61
c155 8 0 4.30126e-20 $X=7.005 $Y=1.095
r156 53 62 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.09 $Y=1.16
+ $X2=8.09 $Y2=1.325
r157 53 61 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.09 $Y=1.16
+ $X2=8.09 $Y2=0.995
r158 52 54 6.35905 $w=3.48e-07 $l=1.85e-07 $layer=LI1_cond $X=8.09 $Y=1.15
+ $X2=7.905 $Y2=1.15
r159 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.09
+ $Y=1.16 $X2=8.09 $Y2=1.16
r160 50 54 35.7257 $w=2.98e-07 $l=9.3e-07 $layer=LI1_cond $X=6.975 $Y=1.125
+ $X2=7.905 $Y2=1.125
r161 48 58 25.55 $w=2.7e-07 $l=1.15e-07 $layer=POLY_cond $X=6.89 $Y=1.23
+ $X2=7.005 $Y2=1.23
r162 47 50 3.29018 $w=4.18e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=1.185
+ $X2=6.975 $Y2=1.185
r163 47 49 6.54147 $w=4.18e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=1.185
+ $X2=6.805 $Y2=1.185
r164 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.89
+ $Y=1.23 $X2=6.89 $Y2=1.23
r165 40 45 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.205 $Y=1.31
+ $X2=6.12 $Y2=1.31
r166 40 49 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.205 $Y=1.31
+ $X2=6.805 $Y2=1.31
r167 37 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.12 $Y=1.395
+ $X2=6.12 $Y2=1.31
r168 37 38 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=6.12 $Y=1.395
+ $X2=6.12 $Y2=2.135
r169 33 45 28.9016 $w=1.68e-07 $l=4.43e-07 $layer=LI1_cond $X=5.677 $Y=1.31
+ $X2=6.12 $Y2=1.31
r170 33 35 21.8286 $w=4.23e-07 $l=8.05e-07 $layer=LI1_cond $X=5.677 $Y=1.225
+ $X2=5.677 $Y2=0.42
r171 29 38 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.035 $Y=2.3
+ $X2=6.12 $Y2=2.135
r172 29 31 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=6.035 $Y=2.3
+ $X2=5.52 $Y2=2.3
r173 24 61 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.15 $Y=0.555
+ $X2=8.15 $Y2=0.995
r174 19 21 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=8.125 $Y=1.57
+ $X2=8.125 $Y2=2.065
r175 18 19 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=8.125 $Y=1.47 $X2=8.125
+ $Y2=1.57
r176 18 62 48.0787 $w=2e-07 $l=1.45e-07 $layer=POLY_cond $X=8.125 $Y=1.47
+ $X2=8.125 $Y2=1.325
r177 14 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.26 $Y=0.73
+ $X2=7.26 $Y2=0.805
r178 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.26 $Y=0.73
+ $X2=7.26 $Y2=0.445
r179 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.005 $Y=1.99
+ $X2=7.005 $Y2=2.275
r180 10 11 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.005 $Y=1.89 $X2=7.005
+ $Y2=1.99
r181 9 58 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=7.005 $Y=1.365
+ $X2=7.005 $Y2=1.23
r182 9 10 174.078 $w=2e-07 $l=5.25e-07 $layer=POLY_cond $X=7.005 $Y=1.365
+ $X2=7.005 $Y2=1.89
r183 8 58 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=7.005 $Y=1.095
+ $X2=7.005 $Y2=1.23
r184 7 27 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=7.005 $Y=0.805
+ $X2=7.26 $Y2=0.805
r185 7 8 71.2891 $w=2e-07 $l=2.15e-07 $layer=POLY_cond $X=7.005 $Y=0.88
+ $X2=7.005 $Y2=1.095
r186 2 31 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=5.375
+ $Y=2.065 $X2=5.52 $Y2=2.3
r187 1 35 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=5.415
+ $Y=0.235 $X2=5.55 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%SET_B 1 3 6 8 10 13 18 22 23 25 26 28 29
+ 31 38
c133 38 0 4.64199e-20 $X=7.52 $Y=1.53
c134 26 0 3.13156e-20 $X=7.715 $Y=1.53
c135 8 0 3.88079e-19 $X=10.26 $Y=1.99
c136 6 0 3.97233e-20 $X=7.62 $Y=0.445
c137 1 0 1.47636e-19 $X=7.595 $Y=1.99
r138 35 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.45
+ $Y=1.68 $X2=7.45 $Y2=1.68
r139 31 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.52 $Y=1.53
+ $X2=7.52 $Y2=1.53
r140 29 44 4.32166 $w=2.78e-07 $l=1.05e-07 $layer=LI1_cond $X=9.72 $Y=1.53
+ $X2=9.72 $Y2=1.635
r141 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.71 $Y=1.53
+ $X2=9.71 $Y2=1.53
r142 26 31 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=7.715 $Y=1.53
+ $X2=7.52 $Y2=1.53
r143 25 28 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.565 $Y=1.53
+ $X2=9.71 $Y2=1.53
r144 25 26 2.2896 $w=1.4e-07 $l=1.85e-06 $layer=MET1_cond $X=9.565 $Y=1.53
+ $X2=7.715 $Y2=1.53
r145 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.53
+ $Y=1.63 $X2=10.53 $Y2=1.63
r146 20 44 3.32261 $w=1.8e-07 $l=1.4e-07 $layer=LI1_cond $X=9.86 $Y=1.635
+ $X2=9.72 $Y2=1.635
r147 20 22 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=9.86 $Y=1.635
+ $X2=10.53 $Y2=1.635
r148 18 23 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=10.53 $Y=1.6
+ $X2=10.53 $Y2=1.63
r149 18 19 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=10.53 $Y=1.6
+ $X2=10.53 $Y2=1.465
r150 17 23 45.5456 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=10.53 $Y=1.835
+ $X2=10.53 $Y2=1.63
r151 13 19 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=10.59 $Y=0.445
+ $X2=10.59 $Y2=1.465
r152 8 17 86.1854 $w=1.51e-07 $l=2.7e-07 $layer=POLY_cond $X=10.26 $Y=1.912
+ $X2=10.53 $Y2=1.912
r153 8 10 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=10.26 $Y=1.99
+ $X2=10.26 $Y2=2.275
r154 4 35 38.571 $w=3.25e-07 $l=2.14942e-07 $layer=POLY_cond $X=7.62 $Y=1.515
+ $X2=7.505 $Y2=1.68
r155 4 6 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=7.62 $Y=1.515
+ $X2=7.62 $Y2=0.445
r156 1 35 55.4962 $w=3.25e-07 $l=3.52136e-07 $layer=POLY_cond $X=7.595 $Y=1.99
+ $X2=7.505 $Y2=1.68
r157 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.595 $Y=1.99
+ $X2=7.595 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_1921_295# 1 2 8 9 11 12 13 16 19 22 23
+ 25 26 29 32 34 37
c104 37 0 1.50109e-19 $X=11.555 $Y=1.28
c105 26 0 5.96508e-20 $X=10.28 $Y=1.28
c106 9 0 1.03798e-20 $X=9.705 $Y=1.99
r107 34 36 6.80499 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=11.515 $Y=0.42
+ $X2=11.515 $Y2=0.585
r108 32 37 3.77418 $w=2.45e-07 $l=9.21954e-08 $layer=LI1_cond $X=11.57 $Y=1.195
+ $X2=11.555 $Y2=1.28
r109 32 36 30.5648 $w=2.28e-07 $l=6.1e-07 $layer=LI1_cond $X=11.57 $Y=1.195
+ $X2=11.57 $Y2=0.585
r110 27 37 3.77418 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=11.555 $Y=1.365
+ $X2=11.555 $Y2=1.28
r111 27 29 40.7788 $w=2.58e-07 $l=9.2e-07 $layer=LI1_cond $X=11.555 $Y=1.365
+ $X2=11.555 $Y2=2.285
r112 25 37 2.68609 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.425 $Y=1.28
+ $X2=11.555 $Y2=1.28
r113 25 26 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=11.425 $Y=1.28
+ $X2=10.28 $Y2=1.28
r114 23 40 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=10.145 $Y=1.02
+ $X2=10.145 $Y2=1.185
r115 23 39 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=10.145 $Y=1.02
+ $X2=10.145 $Y2=0.855
r116 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.12
+ $Y=1.02 $X2=10.12 $Y2=1.02
r117 20 26 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=10.157 $Y=1.195
+ $X2=10.28 $Y2=1.28
r118 20 22 8.23174 $w=2.43e-07 $l=1.75e-07 $layer=LI1_cond $X=10.157 $Y=1.195
+ $X2=10.157 $Y2=1.02
r119 19 40 96.1574 $w=2e-07 $l=2.9e-07 $layer=POLY_cond $X=10.085 $Y=1.475
+ $X2=10.085 $Y2=1.185
r120 16 39 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=10.06 $Y=0.445
+ $X2=10.06 $Y2=0.855
r121 12 19 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=9.985 $Y=1.55
+ $X2=10.085 $Y2=1.475
r122 12 13 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=9.985 $Y=1.55
+ $X2=9.805 $Y2=1.55
r123 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=9.705 $Y=1.99
+ $X2=9.705 $Y2=2.275
r124 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=9.705 $Y=1.89 $X2=9.705
+ $Y2=1.99
r125 7 13 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=9.705 $Y=1.625
+ $X2=9.805 $Y2=1.55
r126 7 8 87.868 $w=2e-07 $l=2.65e-07 $layer=POLY_cond $X=9.705 $Y=1.625
+ $X2=9.705 $Y2=1.89
r127 2 29 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=11.365
+ $Y=2.065 $X2=11.51 $Y2=2.285
r128 1 34 182 $w=1.7e-07 $l=3.34963e-07 $layer=licon1_NDIFF $count=1 $X=11.255
+ $Y=0.235 $X2=11.51 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_1725_329# 1 2 3 12 13 15 16 20 24 26 27
+ 28 29 30 31 35 39 43 46 47 49 51 52 54 58 60
c155 60 0 2.95922e-19 $X=11.04 $Y=1.69
c156 54 0 4.36044e-20 $X=9.605 $Y=1.98
c157 30 0 3.88523e-20 $X=12.265 $Y=1.535
c158 20 0 3.87572e-20 $X=12.24 $Y=0.445
r159 65 67 11.2698 $w=4.1e-07 $l=8.87412e-08 $layer=POLY_cond $X=11.095 $Y=1.205
+ $X2=11.125 $Y2=1.28
r160 61 67 48.2 $w=4.1e-07 $l=4.1e-07 $layer=POLY_cond $X=11.125 $Y=1.69
+ $X2=11.125 $Y2=1.28
r161 60 63 8.79496 $w=3.78e-07 $l=2.9e-07 $layer=LI1_cond $X=11.065 $Y=1.69
+ $X2=11.065 $Y2=1.98
r162 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.04
+ $Y=1.69 $X2=11.04 $Y2=1.69
r163 52 65 49.5896 $w=3.2e-07 $l=2.75e-07 $layer=POLY_cond $X=11.095 $Y=0.93
+ $X2=11.095 $Y2=1.205
r164 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.07
+ $Y=0.93 $X2=11.07 $Y2=0.93
r165 49 51 21.0446 $w=2.28e-07 $l=4.2e-07 $layer=LI1_cond $X=10.65 $Y=0.9
+ $X2=11.07 $Y2=0.9
r166 48 58 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=10.595 $Y=1.98
+ $X2=10.495 $Y2=1.98
r167 47 63 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.875 $Y=1.98
+ $X2=11.065 $Y2=1.98
r168 47 48 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.875 $Y=1.98
+ $X2=10.595 $Y2=1.98
r169 46 49 6.85974 $w=2.3e-07 $l=1.57242e-07 $layer=LI1_cond $X=10.55 $Y=0.785
+ $X2=10.65 $Y2=0.9
r170 45 46 13.3091 $w=1.98e-07 $l=2.4e-07 $layer=LI1_cond $X=10.55 $Y=0.545
+ $X2=10.55 $Y2=0.785
r171 41 58 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=10.495 $Y=2.065
+ $X2=10.495 $Y2=1.98
r172 41 43 12.2 $w=1.98e-07 $l=2.2e-07 $layer=LI1_cond $X=10.495 $Y=2.065
+ $X2=10.495 $Y2=2.285
r173 40 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.69 $Y=1.98
+ $X2=9.605 $Y2=1.98
r174 39 58 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=10.395 $Y=1.98
+ $X2=10.495 $Y2=1.98
r175 39 40 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=10.395 $Y=1.98
+ $X2=9.69 $Y2=1.98
r176 35 45 7.01501 $w=2.7e-07 $l=1.78115e-07 $layer=LI1_cond $X=10.45 $Y=0.41
+ $X2=10.55 $Y2=0.545
r177 35 37 49.0855 $w=2.68e-07 $l=1.15e-06 $layer=LI1_cond $X=10.45 $Y=0.41
+ $X2=9.3 $Y2=0.41
r178 31 54 20.3551 $w=1.68e-07 $l=3.12e-07 $layer=LI1_cond $X=9.605 $Y=2.292
+ $X2=9.605 $Y2=1.98
r179 31 33 22.0168 $w=3.33e-07 $l=6.4e-07 $layer=LI1_cond $X=9.52 $Y=2.292
+ $X2=8.88 $Y2=2.292
r180 27 52 0.901628 $w=3.2e-07 $l=5e-09 $layer=POLY_cond $X=11.095 $Y=0.925
+ $X2=11.095 $Y2=0.93
r181 27 28 45.2492 $w=3.2e-07 $l=1.6e-07 $layer=POLY_cond $X=11.095 $Y=0.925
+ $X2=11.095 $Y2=0.765
r182 24 30 93.4966 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=12.265 $Y=1.77
+ $X2=12.265 $Y2=1.535
r183 24 26 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=12.265 $Y=1.77
+ $X2=12.265 $Y2=2.165
r184 22 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.24 $Y=1.355
+ $X2=12.24 $Y2=1.28
r185 22 30 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=12.24 $Y=1.355
+ $X2=12.24 $Y2=1.535
r186 18 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.24 $Y=1.205
+ $X2=12.24 $Y2=1.28
r187 18 20 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=12.24 $Y=1.205
+ $X2=12.24 $Y2=0.445
r188 17 67 26.4667 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=11.375 $Y=1.28
+ $X2=11.125 $Y2=1.28
r189 16 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.165 $Y=1.28
+ $X2=12.24 $Y2=1.28
r190 16 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=12.165 $Y=1.28
+ $X2=11.375 $Y2=1.28
r191 13 61 50.6865 $w=4.1e-07 $l=3.67423e-07 $layer=POLY_cond $X=11.275 $Y=1.99
+ $X2=11.125 $Y2=1.69
r192 13 15 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=11.275 $Y=1.99
+ $X2=11.275 $Y2=2.275
r193 12 28 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.18 $Y=0.445
+ $X2=11.18 $Y2=0.765
r194 3 43 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=10.35
+ $Y=2.065 $X2=10.495 $Y2=2.285
r195 2 33 600 $w=1.7e-07 $l=7.61906e-07 $layer=licon1_PDIFF $count=1 $X=8.625
+ $Y=1.645 $X2=8.88 $Y2=2.29
r196 1 37 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=9.165
+ $Y=0.235 $X2=9.3 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_2381_47# 1 2 7 9 10 12 15 19 23 26
r50 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.66
+ $Y=1.16 $X2=12.66 $Y2=1.16
r51 21 26 1.0017 $w=3.3e-07 $l=1.7e-07 $layer=LI1_cond $X=12.195 $Y=1.16
+ $X2=12.025 $Y2=1.16
r52 21 23 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=12.195 $Y=1.16
+ $X2=12.66 $Y2=1.16
r53 17 26 5.58832 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=12.025 $Y=1.325
+ $X2=12.025 $Y2=1.16
r54 17 19 22.5404 $w=3.38e-07 $l=6.65e-07 $layer=LI1_cond $X=12.025 $Y=1.325
+ $X2=12.025 $Y2=1.99
r55 13 26 5.58832 $w=3e-07 $l=1.83916e-07 $layer=LI1_cond $X=11.985 $Y=0.995
+ $X2=12.025 $Y2=1.16
r56 13 15 25.2651 $w=2.58e-07 $l=5.7e-07 $layer=LI1_cond $X=11.985 $Y=0.995
+ $X2=11.985 $Y2=0.425
r57 10 24 38.6069 $w=3.31e-07 $l=2.12238e-07 $layer=POLY_cond $X=12.815 $Y=0.995
+ $X2=12.707 $Y2=1.16
r58 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.815 $Y=0.995
+ $X2=12.815 $Y2=0.56
r59 7 24 46.3664 $w=3.31e-07 $l=2.88531e-07 $layer=POLY_cond $X=12.79 $Y=1.41
+ $X2=12.707 $Y2=1.16
r60 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.79 $Y=1.41
+ $X2=12.79 $Y2=1.985
r61 2 19 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=11.905
+ $Y=1.845 $X2=12.03 $Y2=1.99
r62 1 15 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=11.905
+ $Y=0.235 $X2=12.03 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_27_369# 1 2 7 10 11 13 14 16
r46 14 16 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=1.225 $Y=2.36
+ $X2=2.08 $Y2=2.36
r47 13 14 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.14 $Y=2.255
+ $X2=1.225 $Y2=2.36
r48 12 13 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.14 $Y=2.025
+ $X2=1.14 $Y2=2.255
r49 10 12 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.055 $Y=1.935
+ $X2=1.14 $Y2=2.025
r50 10 11 43.7475 $w=1.78e-07 $l=7.1e-07 $layer=LI1_cond $X=1.055 $Y=1.935
+ $X2=0.345 $Y2=1.935
r51 7 11 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=0.215 $Y=2.025
+ $X2=0.345 $Y2=1.935
r52 7 9 2.11154 $w=2.6e-07 $l=4.5e-08 $layer=LI1_cond $X=0.215 $Y=2.025
+ $X2=0.215 $Y2=2.07
r53 2 16 600 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.845 $X2=2.08 $Y2=2.34
r54 1 9 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.07
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%VPWR 1 2 3 4 5 6 7 8 27 31 33 37 41 45 48
+ 49 51 52 53 55 60 65 78 94 95 98 101 104 111 119 123 125
c188 95 0 1.68923e-19 $X=13.11 $Y=2.72
r189 125 126 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r190 121 123 9.7969 $w=6.78e-07 $l=1.15e-07 $layer=LI1_cond $X=8.51 $Y=2.465
+ $X2=8.625 $Y2=2.465
r191 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r192 118 121 11.1693 $w=6.78e-07 $l=6.35e-07 $layer=LI1_cond $X=7.875 $Y=2.465
+ $X2=8.51 $Y2=2.465
r193 118 119 10.6764 $w=6.78e-07 $l=1.65e-07 $layer=LI1_cond $X=7.875 $Y=2.465
+ $X2=7.71 $Y2=2.465
r194 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r195 104 107 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=4.035 $Y=2.36
+ $X2=4.035 $Y2=2.72
r196 102 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r197 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r198 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r199 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r200 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.19 $Y=2.72
+ $X2=13.11 $Y2=2.72
r201 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r202 89 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=12.19 $Y2=2.72
r203 88 91 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=11.27 $Y=2.72
+ $X2=12.19 $Y2=2.72
r204 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r205 86 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.27 $Y2=2.72
r206 86 126 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=9.89 $Y2=2.72
r207 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r208 83 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.19 $Y=2.72
+ $X2=10.025 $Y2=2.72
r209 83 85 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=10.19 $Y=2.72
+ $X2=10.81 $Y2=2.72
r210 82 126 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r211 82 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=8.51 $Y2=2.72
r212 81 123 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.97 $Y=2.72
+ $X2=8.625 $Y2=2.72
r213 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r214 78 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.86 $Y=2.72
+ $X2=10.025 $Y2=2.72
r215 78 81 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=9.86 $Y=2.72
+ $X2=8.97 $Y2=2.72
r216 77 122 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r217 77 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=6.67 $Y2=2.72
r218 76 119 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=7.59 $Y=2.72
+ $X2=7.71 $Y2=2.72
r219 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r220 74 76 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=6.83 $Y=2.72
+ $X2=7.59 $Y2=2.72
r221 72 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r222 71 72 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r223 69 72 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=6.21 $Y2=2.72
r224 69 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r225 68 71 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=6.21 $Y2=2.72
r226 68 69 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r227 66 107 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=4.035 $Y2=2.72
r228 66 68 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=4.37 $Y2=2.72
r229 65 74 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=6.637 $Y=2.72
+ $X2=6.83 $Y2=2.72
r230 65 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r231 65 111 10.7761 $w=3.83e-07 $l=3.6e-07 $layer=LI1_cond $X=6.637 $Y=2.72
+ $X2=6.637 $Y2=2.36
r232 65 71 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.445 $Y=2.72
+ $X2=6.21 $Y2=2.72
r233 64 102 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r234 64 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r235 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r236 61 98 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.835 $Y=2.72
+ $X2=0.675 $Y2=2.72
r237 61 63 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.835 $Y=2.72
+ $X2=1.15 $Y2=2.72
r238 60 101 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=2.94 $Y=2.72
+ $X2=3.087 $Y2=2.72
r239 60 63 116.781 $w=1.68e-07 $l=1.79e-06 $layer=LI1_cond $X=2.94 $Y=2.72
+ $X2=1.15 $Y2=2.72
r240 55 98 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.675 $Y2=2.72
r241 55 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r242 53 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r243 53 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r244 51 91 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=12.435 $Y=2.72
+ $X2=12.19 $Y2=2.72
r245 51 52 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=12.435 $Y=2.72
+ $X2=12.562 $Y2=2.72
r246 50 94 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=12.69 $Y=2.72
+ $X2=13.11 $Y2=2.72
r247 50 52 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=12.69 $Y=2.72
+ $X2=12.562 $Y2=2.72
r248 48 85 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=10.875 $Y=2.72
+ $X2=10.81 $Y2=2.72
r249 48 49 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.875 $Y=2.72
+ $X2=11.065 $Y2=2.72
r250 47 88 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=11.255 $Y=2.72
+ $X2=11.27 $Y2=2.72
r251 47 49 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.255 $Y=2.72
+ $X2=11.065 $Y2=2.72
r252 43 52 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=12.562 $Y=2.635
+ $X2=12.562 $Y2=2.72
r253 43 45 27.7942 $w=2.53e-07 $l=6.15e-07 $layer=LI1_cond $X=12.562 $Y=2.635
+ $X2=12.562 $Y2=2.02
r254 39 49 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=11.065 $Y=2.635
+ $X2=11.065 $Y2=2.72
r255 39 41 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=11.065 $Y=2.635
+ $X2=11.065 $Y2=2.34
r256 35 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.025 $Y=2.635
+ $X2=10.025 $Y2=2.72
r257 35 37 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=10.025 $Y=2.635
+ $X2=10.025 $Y2=2.36
r258 34 101 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=3.235 $Y=2.72
+ $X2=3.087 $Y2=2.72
r259 33 107 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.845 $Y=2.72
+ $X2=4.035 $Y2=2.72
r260 33 34 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.845 $Y=2.72
+ $X2=3.235 $Y2=2.72
r261 29 101 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.087 $Y=2.635
+ $X2=3.087 $Y2=2.72
r262 29 31 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=3.087 $Y=2.635
+ $X2=3.087 $Y2=2.34
r263 25 98 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.675 $Y=2.635
+ $X2=0.675 $Y2=2.72
r264 25 27 9.90381 $w=3.18e-07 $l=2.75e-07 $layer=LI1_cond $X=0.675 $Y=2.635
+ $X2=0.675 $Y2=2.36
r265 8 45 300 $w=1.7e-07 $l=2.45713e-07 $layer=licon1_PDIFF $count=2 $X=12.355
+ $Y=1.845 $X2=12.525 $Y2=2.02
r266 7 41 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=10.915
+ $Y=2.065 $X2=11.04 $Y2=2.34
r267 6 37 600 $w=1.7e-07 $l=3.93542e-07 $layer=licon1_PDIFF $count=1 $X=9.795
+ $Y=2.065 $X2=10.025 $Y2=2.36
r268 5 118 600 $w=1.7e-07 $l=3.78253e-07 $layer=licon1_PDIFF $count=1 $X=7.685
+ $Y=2.065 $X2=7.875 $Y2=2.36
r269 4 111 600 $w=1.7e-07 $l=3.84057e-07 $layer=licon1_PDIFF $count=1 $X=6.405
+ $Y=2.065 $X2=6.61 $Y2=2.36
r270 3 104 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=3.915
+ $Y=1.845 $X2=4.06 $Y2=2.36
r271 2 31 600 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.845 $X2=3.07 $Y2=2.34
r272 1 27 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.845 $X2=0.73 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_201_47# 1 2 3 4 13 19 21 23 28 33 36 37
+ 40 43 44
c126 43 0 4.73773e-19 $X=5.095 $Y=1.53
c127 37 0 1.4475e-19 $X=1.955 $Y=1.53
c128 33 0 1.00357e-19 $X=5.017 $Y=0.78
c129 28 0 1.40323e-19 $X=1.75 $Y=1.965
c130 13 0 4.39648e-20 $X=1.655 $Y=0.425
r131 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.095 $Y=1.53
+ $X2=5.095 $Y2=1.53
r132 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.76 $Y=1.53
+ $X2=1.76 $Y2=1.53
r133 37 39 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=1.955 $Y=1.53
+ $X2=1.76 $Y2=1.53
r134 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.95 $Y=1.53
+ $X2=5.095 $Y2=1.53
r135 36 37 3.70668 $w=1.4e-07 $l=2.995e-06 $layer=MET1_cond $X=4.95 $Y=1.53
+ $X2=1.955 $Y2=1.53
r136 35 44 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=5.095 $Y=1.59
+ $X2=5.095 $Y2=1.53
r137 33 44 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.095 $Y=0.78
+ $X2=5.095 $Y2=1.53
r138 31 40 54.5789 $w=1.88e-07 $l=9.35e-07 $layer=LI1_cond $X=1.75 $Y=0.595
+ $X2=1.75 $Y2=1.53
r139 29 40 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=1.75 $Y=1.845
+ $X2=1.75 $Y2=1.53
r140 28 29 2.10789 $w=1.9e-07 $l=1.2e-07 $layer=LI1_cond $X=1.75 $Y=1.965
+ $X2=1.75 $Y2=1.845
r141 26 28 6.72258 $w=2.38e-07 $l=1.4e-07 $layer=LI1_cond $X=1.61 $Y=1.965
+ $X2=1.75 $Y2=1.965
r142 21 35 6.27261 $w=2.13e-07 $l=1.07e-07 $layer=LI1_cond $X=5.072 $Y=1.697
+ $X2=5.072 $Y2=1.59
r143 21 23 32.322 $w=2.13e-07 $l=6.03e-07 $layer=LI1_cond $X=5.072 $Y=1.697
+ $X2=5.072 $Y2=2.3
r144 17 33 8.35379 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=5.017 $Y=0.618
+ $X2=5.017 $Y2=0.78
r145 17 19 7.02104 $w=3.23e-07 $l=1.98e-07 $layer=LI1_cond $X=5.017 $Y=0.618
+ $X2=5.017 $Y2=0.42
r146 13 31 7.55181 $w=3.4e-07 $l=2.1225e-07 $layer=LI1_cond $X=1.655 $Y=0.425
+ $X2=1.75 $Y2=0.595
r147 13 15 17.4561 $w=3.38e-07 $l=5.15e-07 $layer=LI1_cond $X=1.655 $Y=0.425
+ $X2=1.14 $Y2=0.425
r148 4 23 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=4.925
+ $Y=2.065 $X2=5.05 $Y2=2.3
r149 3 26 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.465
+ $Y=1.845 $X2=1.61 $Y2=1.97
r150 2 19 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.235 $X2=5.08 $Y2=0.42
r151 1 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.235 $X2=1.14 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%Q 1 2 7 8 9 10 11 12 20
r11 12 35 2.65948 $w=3.23e-07 $l=7.5e-08 $layer=LI1_cond $X=13.077 $Y=2.21
+ $X2=13.077 $Y2=2.285
r12 11 12 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=13.077 $Y=1.87
+ $X2=13.077 $Y2=2.21
r13 10 11 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=13.077 $Y=1.53
+ $X2=13.077 $Y2=1.87
r14 9 10 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=13.077 $Y=1.19
+ $X2=13.077 $Y2=1.53
r15 8 9 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=13.077 $Y=0.85
+ $X2=13.077 $Y2=1.19
r16 7 8 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=13.077 $Y=0.51
+ $X2=13.077 $Y2=0.85
r17 7 20 2.48218 $w=3.23e-07 $l=7e-08 $layer=LI1_cond $X=13.077 $Y=0.51
+ $X2=13.077 $Y2=0.44
r18 2 35 600 $w=1.7e-07 $l=8.69483e-07 $layer=licon1_PDIFF $count=1 $X=12.88
+ $Y=1.485 $X2=13.025 $Y2=2.285
r19 1 20 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=12.89
+ $Y=0.235 $X2=13.025 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_1%VGND 1 2 3 4 5 6 7 8 25 26 29 31 35 39 43
+ 47 50 51 53 54 56 57 58 64 90 91 102 105 116 120
c172 91 0 2.71124e-20 $X=13.11 $Y=0
c173 64 0 6.74919e-20 $X=6.06 $Y=0
r174 118 120 13.5844 $w=8.88e-07 $l=2.65e-07 $layer=LI1_cond $X=8.05 $Y=0.36
+ $X2=8.315 $Y2=0.36
r175 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r176 115 118 2.19326 $w=8.88e-07 $l=1.6e-07 $layer=LI1_cond $X=7.89 $Y=0.36
+ $X2=8.05 $Y2=0.36
r177 115 116 18.6563 $w=8.88e-07 $l=6.35e-07 $layer=LI1_cond $X=7.89 $Y=0.36
+ $X2=7.255 $Y2=0.36
r178 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r179 103 106 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=2.99 $Y2=0
r180 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r181 100 103 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=2.07 $Y2=0
r182 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r183 97 99 8.43408 $w=6.22e-07 $l=4.3e-07 $layer=LI1_cond $X=0.26 $Y=0.255
+ $X2=0.69 $Y2=0.255
r184 94 97 0.588424 $w=6.22e-07 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=0.255
+ $X2=0.26 $Y2=0.255
r185 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r186 88 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.19 $Y=0
+ $X2=13.11 $Y2=0
r187 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r188 85 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=12.19 $Y2=0
r189 84 87 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=11.27 $Y=0
+ $X2=12.19 $Y2=0
r190 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r191 82 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.27 $Y2=0
r192 81 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r193 79 82 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=10.81 $Y2=0
r194 79 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.05 $Y2=0
r195 78 81 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=8.51 $Y=0 $X2=10.81
+ $Y2=0
r196 78 120 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=8.51 $Y=0
+ $X2=8.315 $Y2=0
r197 78 79 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r198 75 119 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r199 75 110 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=6.21 $Y2=0
r200 74 116 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.13 $Y=0
+ $X2=7.255 $Y2=0
r201 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r202 72 74 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=6.595 $Y=0
+ $X2=7.13 $Y2=0
r203 70 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.21 $Y2=0
r204 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r205 67 70 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.75 $Y2=0
r206 66 69 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.37 $Y=0 $X2=5.75
+ $Y2=0
r207 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r208 64 112 8.49551 $w=5.33e-07 $l=3.8e-07 $layer=LI1_cond $X=6.327 $Y=0
+ $X2=6.327 $Y2=0.38
r209 64 72 7.58357 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=6.327 $Y=0
+ $X2=6.595 $Y2=0
r210 64 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r211 64 69 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.06 $Y=0 $X2=5.75
+ $Y2=0
r212 63 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r213 63 106 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=2.99 $Y2=0
r214 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r215 60 105 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.35 $Y=0
+ $X2=3.145 $Y2=0
r216 60 62 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.35 $Y=0 $X2=3.91
+ $Y2=0
r217 58 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r218 58 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r219 56 87 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=12.285 $Y=0
+ $X2=12.19 $Y2=0
r220 56 57 9.89127 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=12.285 $Y=0
+ $X2=12.487 $Y2=0
r221 55 90 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=12.69 $Y=0
+ $X2=13.11 $Y2=0
r222 55 57 9.89127 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=12.69 $Y=0
+ $X2=12.487 $Y2=0
r223 53 81 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=10.835 $Y=0
+ $X2=10.81 $Y2=0
r224 53 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.835 $Y=0
+ $X2=10.96 $Y2=0
r225 52 84 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=11.085 $Y=0
+ $X2=11.27 $Y2=0
r226 52 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.085 $Y=0
+ $X2=10.96 $Y2=0
r227 50 62 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.925 $Y=0 $X2=3.91
+ $Y2=0
r228 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.925 $Y=0 $X2=4.09
+ $Y2=0
r229 49 66 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.255 $Y=0
+ $X2=4.37 $Y2=0
r230 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.255 $Y=0 $X2=4.09
+ $Y2=0
r231 45 57 1.50354 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=12.487 $Y=0.085
+ $X2=12.487 $Y2=0
r232 45 47 7.82523 $w=4.03e-07 $l=2.75e-07 $layer=LI1_cond $X=12.487 $Y=0.085
+ $X2=12.487 $Y2=0.36
r233 41 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.96 $Y=0.085
+ $X2=10.96 $Y2=0
r234 41 43 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=10.96 $Y=0.085
+ $X2=10.96 $Y2=0.36
r235 37 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.09 $Y=0.085
+ $X2=4.09 $Y2=0
r236 37 39 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.09 $Y=0.085
+ $X2=4.09 $Y2=0.36
r237 33 105 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.145 $Y=0.085
+ $X2=3.145 $Y2=0
r238 33 35 8.29197 $w=4.08e-07 $l=2.95e-07 $layer=LI1_cond $X=3.145 $Y=0.085
+ $X2=3.145 $Y2=0.38
r239 32 102 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.29 $Y=0
+ $X2=2.157 $Y2=0
r240 31 105 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.94 $Y=0
+ $X2=3.145 $Y2=0
r241 31 32 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.94 $Y=0 $X2=2.29
+ $Y2=0
r242 27 102 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.157 $Y=0.085
+ $X2=2.157 $Y2=0
r243 27 29 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=2.157 $Y=0.085
+ $X2=2.157 $Y2=0.38
r244 26 99 8.44605 $w=6.22e-07 $l=2.83417e-07 $layer=LI1_cond $X=0.75 $Y=0
+ $X2=0.69 $Y2=0.255
r245 25 102 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=2.157 $Y2=0
r246 25 26 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=0.75 $Y2=0
r247 8 47 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=12.315
+ $Y=0.235 $X2=12.525 $Y2=0.36
r248 7 43 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=10.665
+ $Y=0.235 $X2=10.92 $Y2=0.36
r249 6 115 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=7.695
+ $Y=0.235 $X2=7.89 $Y2=0.36
r250 5 112 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.295
+ $Y=0.235 $X2=6.43 $Y2=0.38
r251 4 39 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.955
+ $Y=0.235 $X2=4.09 $Y2=0.36
r252 3 35 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.965
+ $Y=0.235 $X2=3.1 $Y2=0.38
r253 2 29 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.235 $X2=2.11 $Y2=0.38
r254 1 97 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends

