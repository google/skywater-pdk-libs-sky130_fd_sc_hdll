* NGSPICE file created from sky130_fd_sc_hdll__and4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__and4b_1 A_N B C D VGND VNB VPB VPWR X
M1000 a_379_47# B a_307_47# VNB nshort w=420000u l=150000u
+  ad=2.1e+11p pd=1.84e+06u as=8.82e+10p ps=1.26e+06u
M1001 VPWR A_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=7.115e+11p pd=6.35e+06u as=1.134e+11p ps=1.38e+06u
M1002 a_509_47# C a_379_47# VNB nshort w=420000u l=150000u
+  ad=1.491e+11p pd=1.55e+06u as=0p ps=0u
M1003 X a_213_413# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=3.422e+11p ps=3.43e+06u
M1004 VPWR B a_213_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=3.171e+11p ps=3.19e+06u
M1005 VGND D a_509_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_213_413# a_27_47# VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_213_413# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1008 VGND A_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1009 a_213_413# C VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR D a_213_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_307_47# a_27_47# a_213_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
.ends

