* File: sky130_fd_sc_hdll__nand4bb_4.spice
* Created: Thu Aug 27 19:15:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nand4bb_4.pex.spice"
.subckt sky130_fd_sc_hdll__nand4bb_4  VNB VPB A_N B_N C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B_N	B_N
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1021 N_VGND_M1021_d N_A_N_M1021_g N_A_27_47#_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.092625 AS=0.2015 PD=0.935 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1013 N_A_206_47#_M1013_d N_B_N_M1013_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.65
+ AD=0.312 AS=0.092625 PD=2.26 PS=0.935 NRD=20.304 NRS=1.836 M=1 R=4.33333
+ SA=75000.7 SB=75000.4 A=0.0975 P=1.6 MULT=1
MM1007 N_Y_M1007_d N_A_27_47#_M1007_g N_A_395_47#_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.2015 PD=0.97 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1032 N_Y_M1007_d N_A_27_47#_M1032_g N_A_395_47#_M1032_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75003 A=0.0975 P=1.6 MULT=1
MM1033 N_Y_M1033_d N_A_27_47#_M1033_g N_A_395_47#_M1032_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.2 SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1035 N_Y_M1033_d N_A_27_47#_M1035_g N_A_395_47#_M1035_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1002 N_A_395_47#_M1035_s N_A_206_47#_M1002_g N_A_853_47#_M1002_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1
+ R=4.33333 SA=75002.1 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1008 N_A_395_47#_M1008_d N_A_206_47#_M1008_g N_A_853_47#_M1002_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75002.5 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1025 N_A_395_47#_M1008_d N_A_206_47#_M1025_g N_A_853_47#_M1025_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1
+ R=4.33333 SA=75003 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1028 N_A_395_47#_M1028_d N_A_206_47#_M1028_g N_A_853_47#_M1025_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1
+ R=4.33333 SA=75003.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_A_1251_47#_M1000_d N_C_M1000_g N_A_853_47#_M1000_s VNB NSHORT L=0.15
+ W=0.65 AD=0.221 AS=0.104 PD=1.98 PS=0.97 NRD=4.608 NRS=3.684 M=1 R=4.33333
+ SA=75000.3 SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1009 N_A_1251_47#_M1009_d N_C_M1009_g N_A_853_47#_M1000_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=2.76 NRS=3.684 M=1 R=4.33333
+ SA=75000.7 SB=75003 A=0.0975 P=1.6 MULT=1
MM1011 N_A_1251_47#_M1009_d N_C_M1011_g N_A_853_47#_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=4.608 NRS=3.684 M=1 R=4.33333
+ SA=75001.2 SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1020 N_A_1251_47#_M1020_d N_C_M1020_g N_A_853_47#_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75001.7 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1016 N_A_1251_47#_M1020_d N_D_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.1
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1018 N_A_1251_47#_M1018_d N_D_M1018_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=5.532 NRS=0 M=1 R=4.33333 SA=75002.6
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1026 N_A_1251_47#_M1018_d N_D_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=1.836 NRS=8.304 M=1 R=4.33333 SA=75003
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1030 N_A_1251_47#_M1030_d N_D_M1030_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.21125 AS=0.104 PD=1.95 PS=0.97 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1014 N_VPWR_M1014_d N_A_N_M1014_g N_A_27_47#_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1001 N_A_206_47#_M1001_d N_B_N_M1001_g N_VPWR_M1014_d VPB PHIGHVT L=0.18 W=1
+ AD=0.455 AS=0.145 PD=2.91 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.4 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A_27_47#_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90007.8 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1010_d N_A_27_47#_M1010_g N_Y_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90007.3 A=0.18 P=2.36 MULT=1
MM1022 N_VPWR_M1010_d N_A_27_47#_M1022_g N_Y_M1022_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90006.9 A=0.18 P=2.36 MULT=1
MM1034 N_VPWR_M1034_d N_A_27_47#_M1034_g N_Y_M1022_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90006.4 A=0.18 P=2.36 MULT=1
MM1003 N_Y_M1003_d N_A_206_47#_M1003_g N_VPWR_M1034_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90005.9 A=0.18 P=2.36 MULT=1
MM1015 N_Y_M1003_d N_A_206_47#_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90005.4 A=0.18 P=2.36 MULT=1
MM1019 N_Y_M1019_d N_A_206_47#_M1019_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90005 A=0.18 P=2.36 MULT=1
MM1031 N_Y_M1019_d N_A_206_47#_M1031_g N_VPWR_M1031_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.42 PD=1.29 PS=1.84 NRD=0.9653 NRS=10.8153 M=1 R=5.55556
+ SA=90003.5 SB=90004.5 A=0.18 P=2.36 MULT=1
MM1005 N_Y_M1005_d N_C_M1005_g N_VPWR_M1031_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.42 PD=1.29 PS=1.84 NRD=0.9653 NRS=31.5003 M=1 R=5.55556 SA=90004.5
+ SB=90003.5 A=0.18 P=2.36 MULT=1
MM1023 N_Y_M1005_d N_C_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90005 SB=90003
+ A=0.18 P=2.36 MULT=1
MM1027 N_Y_M1027_d N_C_M1027_g N_VPWR_M1023_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90005.4
+ SB=90002.5 A=0.18 P=2.36 MULT=1
MM1029 N_Y_M1027_d N_C_M1029_g N_VPWR_M1029_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90005.9
+ SB=90002.1 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1029_s N_D_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90006.4
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_D_M1012_g N_Y_M1006_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90006.8
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1017 N_VPWR_M1012_d N_D_M1017_g N_Y_M1017_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90007.3
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1024 N_VPWR_M1024_d N_D_M1024_g N_Y_M1017_s VPB PHIGHVT L=0.18 W=1 AD=0.285
+ AS=0.145 PD=2.57 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90007.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX36_noxref VNB VPB NWDIODE A=17.5908 P=25.13
c_54 VNB 0 2.7314e-19 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hdll__nand4bb_4.pxi.spice"
*
.ends
*
*
