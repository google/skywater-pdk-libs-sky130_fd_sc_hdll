# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__mux2i_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__mux2i_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.590000 0.995000 1.235000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.355000 0.995000 4.050000 1.325000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  1.387500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.245000 1.075000 6.530000 1.290000 ;
        RECT 6.360000 1.290000 6.530000 1.425000 ;
        RECT 6.360000 1.425000 8.650000 1.595000 ;
        RECT 8.480000 0.995000 8.650000 1.425000 ;
    END
  END S
  PIN VGND
    ANTENNADIFFAREA  1.030250 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.475000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  2.339500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.315000 4.185000 0.485000 ;
        RECT 0.095000 0.485000 0.320000 2.255000 ;
        RECT 0.095000 2.255000 4.185000 2.425000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.515000  0.655000 1.850000 0.825000 ;
      RECT 0.515000  1.575000 6.130000 1.745000 ;
      RECT 1.455000  0.825000 1.850000 0.935000 ;
      RECT 2.395000  0.655000 6.035000 0.825000 ;
      RECT 2.395000  1.915000 7.915000 2.085000 ;
      RECT 4.375000  0.085000 4.705000 0.465000 ;
      RECT 4.375000  2.255000 4.705000 2.635000 ;
      RECT 4.925000  0.255000 5.095000 0.655000 ;
      RECT 5.265000  0.085000 5.645000 0.465000 ;
      RECT 5.265000  2.255000 5.645000 2.635000 ;
      RECT 5.865000  0.255000 6.035000 0.655000 ;
      RECT 6.205000  0.085000 6.580000 0.590000 ;
      RECT 6.205000  2.255000 6.585000 2.635000 ;
      RECT 6.800000  0.255000 6.975000 0.715000 ;
      RECT 6.800000  0.715000 7.915000 0.905000 ;
      RECT 6.800000  0.905000 7.100000 0.935000 ;
      RECT 6.805000  1.795000 6.975000 1.915000 ;
      RECT 6.805000  2.085000 6.975000 2.465000 ;
      RECT 7.145000  2.255000 7.525000 2.635000 ;
      RECT 7.245000  0.085000 7.495000 0.545000 ;
      RECT 7.430000  1.075000 8.310000 1.245000 ;
      RECT 7.745000  0.510000 7.915000 0.715000 ;
      RECT 7.745000  1.795000 7.915000 1.915000 ;
      RECT 7.745000  2.085000 7.915000 2.465000 ;
      RECT 8.090000  0.655000 9.045000 0.825000 ;
      RECT 8.090000  0.825000 8.310000 1.075000 ;
      RECT 8.235000  0.085000 8.565000 0.465000 ;
      RECT 8.235000  2.255000 8.565000 2.635000 ;
      RECT 8.785000  0.255000 9.045000 0.655000 ;
      RECT 8.785000  1.795000 9.045000 2.465000 ;
      RECT 8.870000  0.825000 9.045000 1.795000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.680000  0.765000 1.850000 0.935000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.800000  0.765000 6.970000 0.935000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
    LAYER met1 ;
      RECT 1.620000 0.735000 1.910000 0.780000 ;
      RECT 1.620000 0.780000 7.030000 0.920000 ;
      RECT 1.620000 0.920000 1.910000 0.965000 ;
      RECT 6.690000 0.735000 7.030000 0.780000 ;
      RECT 6.690000 0.920000 7.030000 0.965000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2i_4
END LIBRARY
