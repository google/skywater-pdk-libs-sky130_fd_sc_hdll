* NGSPICE file created from sky130_fd_sc_hdll__and2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__and2b_1 A_N B VGND VNB VPB VPWR X
M1000 VPWR A_N a_27_413# VPB phighvt w=420000u l=180000u
+  ad=6.422e+11p pd=5.18e+06u as=1.134e+11p ps=1.38e+06u
M1001 VGND B a_327_47# VNB nshort w=420000u l=150000u
+  ad=3.653e+11p pd=3.54e+06u as=1.218e+11p ps=1.42e+06u
M1002 a_225_413# a_27_413# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1003 a_327_47# a_27_413# a_225_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1004 X a_225_413# VGND VNB nshort w=650000u l=150000u
+  ad=1.95e+11p pd=1.9e+06u as=0p ps=0u
M1005 X a_225_413# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.1e+11p pd=2.62e+06u as=0p ps=0u
M1006 a_27_413# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1007 VPWR B a_225_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

