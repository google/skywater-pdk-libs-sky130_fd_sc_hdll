* File: sky130_fd_sc_hdll__xnor3_2.pex.spice
* Created: Wed Sep  2 08:54:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__XNOR3_2%A_79_21# 1 2 7 9 10 12 13 15 16 18 22 24
+ 25 26 27 29 31 33 34 36 38 40 42 46
r108 45 46 0.654891 $w=3.68e-07 $l=5e-09 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=0.99 $Y2=1.202
r109 44 45 64.1793 $w=3.68e-07 $l=4.9e-07 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.985 $Y2=1.202
r110 43 44 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r111 38 42 11.3723 $w=1.98e-07 $l=2e-07 $layer=LI1_cond $X=2.88 $Y=0.355
+ $X2=2.68 $Y2=0.355
r112 38 40 6.65455 $w=1.98e-07 $l=1.2e-07 $layer=LI1_cond $X=2.88 $Y=0.355 $X2=3
+ $Y2=0.355
r113 34 36 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=1.83 $Y=2.32
+ $X2=2.925 $Y2=2.32
r114 33 42 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=1.715 $Y=0.34
+ $X2=2.68 $Y2=0.34
r115 31 34 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.72 $Y=2.235
+ $X2=1.83 $Y2=2.32
r116 30 31 9.95292 $w=2.18e-07 $l=1.9e-07 $layer=LI1_cond $X=1.72 $Y=2.045
+ $X2=1.72 $Y2=2.235
r117 28 33 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.605 $Y=0.425
+ $X2=1.715 $Y2=0.34
r118 28 29 14.1436 $w=2.18e-07 $l=2.7e-07 $layer=LI1_cond $X=1.605 $Y=0.425
+ $X2=1.605 $Y2=0.695
r119 26 30 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.61 $Y=1.96
+ $X2=1.72 $Y2=2.045
r120 26 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.61 $Y=1.96
+ $X2=1.265 $Y2=1.96
r121 24 29 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.495 $Y=0.78
+ $X2=1.605 $Y2=0.695
r122 24 25 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.495 $Y=0.78
+ $X2=1.265 $Y2=0.78
r123 23 46 20.3016 $w=3.68e-07 $l=1.55e-07 $layer=POLY_cond $X=1.145 $Y=1.202
+ $X2=0.99 $Y2=1.202
r124 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.145
+ $Y=1.16 $X2=1.145 $Y2=1.16
r125 20 27 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.155 $Y=1.875
+ $X2=1.265 $Y2=1.96
r126 20 22 37.4544 $w=2.18e-07 $l=7.15e-07 $layer=LI1_cond $X=1.155 $Y=1.875
+ $X2=1.155 $Y2=1.16
r127 19 25 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.155 $Y=0.865
+ $X2=1.265 $Y2=0.78
r128 19 22 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=1.155 $Y=0.865
+ $X2=1.155 $Y2=1.16
r129 16 46 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r130 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r131 13 45 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r132 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r133 10 44 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r134 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r135 7 43 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.202
r136 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r137 2 36 600 $w=1.7e-07 $l=7.64068e-07 $layer=licon1_PDIFF $count=1 $X=2.78
+ $Y=1.625 $X2=2.925 $Y2=2.32
r138 1 40 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.855
+ $Y=0.245 $X2=3 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_2%C 1 3 7 8 10 11 13 15 18 19
c60 19 0 2.74598e-20 $X=2.53 $Y=1.19
c61 1 0 1.70967e-19 $X=1.565 $Y=0.995
r62 19 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.525
+ $Y=1.16 $X2=2.525 $Y2=1.16
r63 18 22 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=2.59 $Y=1.16
+ $X2=2.525 $Y2=1.16
r64 14 22 146.009 $w=3.3e-07 $l=8.35e-07 $layer=POLY_cond $X=1.69 $Y=1.16
+ $X2=2.525 $Y2=1.16
r65 14 15 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.69 $Y=1.16
+ $X2=1.59 $Y2=1.202
r66 11 18 39.7875 $w=2.42e-07 $l=1.9182e-07 $layer=POLY_cond $X=2.78 $Y=0.995
+ $X2=2.722 $Y2=1.16
r67 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.78 $Y=0.995
+ $X2=2.78 $Y2=0.565
r68 8 18 80.9439 $w=2.42e-07 $l=4.05685e-07 $layer=POLY_cond $X=2.69 $Y=1.55
+ $X2=2.722 $Y2=1.16
r69 8 10 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=2.69 $Y=1.55 $X2=2.69
+ $Y2=2.045
r70 4 15 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=1.59 $Y=1.41
+ $X2=1.59 $Y2=1.202
r71 4 7 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.59 $Y=1.41 $X2=1.59
+ $Y2=1.805
r72 1 15 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=1.565 $Y=0.995
+ $X2=1.59 $Y2=1.202
r73 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.565 $Y=0.995
+ $X2=1.565 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_2%A_328_93# 1 2 7 9 10 12 13 18 20 23 24 28
r72 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.2
+ $Y=1.16 $X2=3.2 $Y2=1.16
r73 25 28 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.095 $Y=1.16
+ $X2=3.2 $Y2=1.16
r74 22 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=1.325
+ $X2=3.095 $Y2=1.16
r75 22 23 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.095 $Y=1.325
+ $X2=3.095 $Y2=1.535
r76 21 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=1.62
+ $X2=1.97 $Y2=1.62
r77 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.01 $Y=1.62
+ $X2=3.095 $Y2=1.535
r78 20 21 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=3.01 $Y=1.62
+ $X2=2.055 $Y2=1.62
r79 16 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.97 $Y=1.535
+ $X2=1.97 $Y2=1.62
r80 16 18 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.97 $Y=1.535
+ $X2=1.97 $Y2=0.76
r81 13 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.885 $Y=1.62
+ $X2=1.97 $Y2=1.62
r82 13 15 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=1.885 $Y=1.62 $X2=1.825
+ $Y2=1.62
r83 10 29 38.578 $w=2.95e-07 $l=1.67481e-07 $layer=POLY_cond $X=3.22 $Y=0.995
+ $X2=3.225 $Y2=1.16
r84 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.22 $Y=0.995
+ $X2=3.22 $Y2=0.565
r85 7 29 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=3.225 $Y=1.41
+ $X2=3.225 $Y2=1.16
r86 7 9 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=3.225 $Y=1.41
+ $X2=3.225 $Y2=1.905
r87 2 15 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.68
+ $Y=1.485 $X2=1.825 $Y2=1.62
r88 1 18 182 $w=1.7e-07 $l=4.54148e-07 $layer=licon1_NDIFF $count=1 $X=1.64
+ $Y=0.465 $X2=1.97 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_2%A_885_297# 1 2 7 9 12 15 16 18 21 22 23 27
+ 35 37 38 39 40 47 49 50 55 57 60
c183 55 0 1.24749e-19 $X=7.75 $Y=1.11
c184 27 0 1.36535e-19 $X=4.73 $Y=1.58
r185 55 58 37.8858 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=7.772 $Y=1.11
+ $X2=7.772 $Y2=1.275
r186 55 57 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=7.772 $Y=1.11
+ $X2=7.772 $Y2=0.945
r187 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.75
+ $Y=1.11 $X2=7.75 $Y2=1.11
r188 50 56 11.8358 $w=2.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.68 $Y=0.85
+ $X2=7.68 $Y2=1.11
r189 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.63 $Y=0.85
+ $X2=7.63 $Y2=0.85
r190 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.15 $Y=0.85
+ $X2=6.15 $Y2=0.85
r191 42 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.67 $Y=0.85
+ $X2=4.67 $Y2=0.85
r192 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.295 $Y=0.85
+ $X2=6.15 $Y2=0.85
r193 39 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.485 $Y=0.85
+ $X2=7.63 $Y2=0.85
r194 39 40 1.47277 $w=1.4e-07 $l=1.19e-06 $layer=MET1_cond $X=7.485 $Y=0.85
+ $X2=6.295 $Y2=0.85
r195 38 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.815 $Y=0.85
+ $X2=4.67 $Y2=0.85
r196 37 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.005 $Y=0.85
+ $X2=6.15 $Y2=0.85
r197 37 38 1.47277 $w=1.4e-07 $l=1.19e-06 $layer=MET1_cond $X=6.005 $Y=0.85
+ $X2=4.815 $Y2=0.85
r198 35 47 7.65801 $w=2.08e-07 $l=1.45e-07 $layer=LI1_cond $X=6.13 $Y=0.995
+ $X2=6.13 $Y2=0.85
r199 31 35 6.28605 $w=2.73e-07 $l=1.5e-07 $layer=LI1_cond $X=5.98 $Y=1.132
+ $X2=6.13 $Y2=1.132
r200 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.98
+ $Y=1.16 $X2=5.98 $Y2=1.16
r201 28 60 28.0163 $w=2.88e-07 $l=7.05e-07 $layer=LI1_cond $X=4.73 $Y=1.445
+ $X2=4.73 $Y2=0.74
r202 27 28 0.275955 $w=2.9e-07 $l=1.35e-07 $layer=LI1_cond $X=4.73 $Y=1.58
+ $X2=4.73 $Y2=1.445
r203 25 27 6.82929 $w=2.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.57 $Y=1.58
+ $X2=4.73 $Y2=1.58
r204 22 32 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=6.24 $Y=1.16
+ $X2=5.98 $Y2=1.16
r205 22 23 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=6.24 $Y=1.16
+ $X2=6.34 $Y2=1.202
r206 21 57 131.747 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=7.855 $Y=0.535
+ $X2=7.855 $Y2=0.945
r207 16 18 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=7.83 $Y=1.57
+ $X2=7.83 $Y2=2.065
r208 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.83 $Y=1.47 $X2=7.83
+ $Y2=1.57
r209 15 58 64.6575 $w=2e-07 $l=1.95e-07 $layer=POLY_cond $X=7.83 $Y=1.47
+ $X2=7.83 $Y2=1.275
r210 10 23 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=6.365 $Y=0.995
+ $X2=6.34 $Y2=1.202
r211 10 12 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=6.365 $Y=0.995
+ $X2=6.365 $Y2=0.455
r212 7 23 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=6.34 $Y=1.41
+ $X2=6.34 $Y2=1.202
r213 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=6.34 $Y=1.41
+ $X2=6.34 $Y2=1.805
r214 2 25 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.425
+ $Y=1.485 $X2=4.57 $Y2=1.63
r215 1 60 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.655
+ $Y=0.235 $X2=4.79 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_2%B 1 3 6 8 9 13 16 18 19 22 24 25 28 31 35
+ 36 38 39 42 45
c136 39 0 1.94872e-19 $X=7.5 $Y=1.445
r137 39 45 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=7.585 $Y=1.53
+ $X2=7.58 $Y2=1.53
r138 38 45 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.355 $Y=1.53
+ $X2=7.58 $Y2=1.53
r139 36 43 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.245 $Y=1.16
+ $X2=7.245 $Y2=1.325
r140 36 42 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.245 $Y=1.16
+ $X2=7.245 $Y2=0.995
r141 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.22
+ $Y=1.16 $X2=7.22 $Y2=1.16
r142 33 38 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=7.245 $Y=1.445
+ $X2=7.355 $Y2=1.53
r143 33 35 14.9294 $w=2.18e-07 $l=2.85e-07 $layer=LI1_cond $X=7.245 $Y=1.445
+ $X2=7.245 $Y2=1.16
r144 31 32 29.1618 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=5.535 $Y=1.16
+ $X2=5.535 $Y2=1.085
r145 26 28 174.919 $w=1.8e-07 $l=4.5e-07 $layer=POLY_cond $X=7.185 $Y=2.415
+ $X2=7.185 $Y2=1.965
r146 25 28 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=7.185 $Y=1.57
+ $X2=7.185 $Y2=1.965
r147 24 25 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.185 $Y=1.47 $X2=7.185
+ $Y2=1.57
r148 24 43 48.0787 $w=2e-07 $l=1.45e-07 $layer=POLY_cond $X=7.185 $Y=1.47
+ $X2=7.185 $Y2=1.325
r149 22 42 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.16 $Y=0.565
+ $X2=7.16 $Y2=0.995
r150 18 26 27.2212 $w=1.5e-07 $l=1.67705e-07 $layer=POLY_cond $X=7.085 $Y=2.54
+ $X2=7.185 $Y2=2.415
r151 18 19 743.511 $w=1.5e-07 $l=1.45e-06 $layer=POLY_cond $X=7.085 $Y=2.54
+ $X2=5.635 $Y2=2.54
r152 16 32 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.56 $Y=0.565
+ $X2=5.56 $Y2=1.085
r153 11 19 27.2212 $w=1.5e-07 $l=1.36015e-07 $layer=POLY_cond $X=5.535 $Y=2.455
+ $X2=5.635 $Y2=2.54
r154 11 13 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=5.535 $Y=2.455
+ $X2=5.535 $Y2=1.905
r155 10 31 83.702 $w=2e-07 $l=2.5e-07 $layer=POLY_cond $X=5.535 $Y=1.41
+ $X2=5.535 $Y2=1.16
r156 10 13 192.411 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=5.535 $Y=1.41
+ $X2=5.535 $Y2=1.905
r157 8 31 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=5.435 $Y=1.16
+ $X2=5.535 $Y2=1.16
r158 8 9 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=5.435 $Y=1.16
+ $X2=4.655 $Y2=1.16
r159 4 9 21.6156 $w=2.33e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.58 $Y=1.085
+ $X2=4.655 $Y2=1.16
r160 4 6 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.58 $Y=1.085
+ $X2=4.58 $Y2=0.56
r161 1 4 50.6824 $w=2.33e-07 $l=3.43642e-07 $layer=POLY_cond $X=4.335 $Y=1.322
+ $X2=4.58 $Y2=1.085
r162 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.335 $Y=1.41
+ $X2=4.335 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_2%A 1 3 4 6 7
c35 1 0 3.84251e-19 $X=8.385 $Y=1.41
r36 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.28
+ $Y=1.16 $X2=8.28 $Y2=1.16
r37 7 11 10.833 $w=2.48e-07 $l=2.35e-07 $layer=LI1_cond $X=8.515 $Y=1.2 $X2=8.28
+ $Y2=1.2
r38 4 10 38.532 $w=3.11e-07 $l=2.07123e-07 $layer=POLY_cond $X=8.41 $Y=0.995
+ $X2=8.315 $Y2=1.16
r39 4 6 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.41 $Y=0.995 $X2=8.41
+ $Y2=0.555
r40 1 10 47.2262 $w=3.11e-07 $l=2.82843e-07 $layer=POLY_cond $X=8.385 $Y=1.41
+ $X2=8.315 $Y2=1.16
r41 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.385 $Y=1.41
+ $X2=8.385 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_2%A_1003_297# 1 2 3 4 13 15 16 18 21 23 27
+ 28 29 30 36 37 40 43 44
c132 30 0 1.20335e-19 $X=8.95 $Y=1.495
c133 29 0 1.89379e-19 $X=8.95 $Y=1.325
r134 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.14 $Y=0.51
+ $X2=8.14 $Y2=0.51
r135 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.18 $Y=0.51
+ $X2=5.18 $Y2=0.51
r136 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.325 $Y=0.51
+ $X2=5.18 $Y2=0.51
r137 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.995 $Y=0.51
+ $X2=8.14 $Y2=0.51
r138 36 37 3.30445 $w=1.4e-07 $l=2.67e-06 $layer=MET1_cond $X=7.995 $Y=0.51
+ $X2=5.325 $Y2=0.51
r139 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.01
+ $Y=1.16 $X2=9.01 $Y2=1.16
r140 32 34 17.9567 $w=2.31e-07 $l=3.4e-07 $layer=LI1_cond $X=9.005 $Y=0.82
+ $X2=9.005 $Y2=1.16
r141 31 44 8.94137 $w=2.88e-07 $l=2.25e-07 $layer=LI1_cond $X=8.17 $Y=0.735
+ $X2=8.17 $Y2=0.51
r142 29 34 9.58904 $w=2.31e-07 $l=1.90526e-07 $layer=LI1_cond $X=8.95 $Y=1.325
+ $X2=9.005 $Y2=1.16
r143 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.95 $Y=1.325
+ $X2=8.95 $Y2=1.495
r144 28 31 14.5133 $w=1.17e-07 $l=1.8262e-07 $layer=LI1_cond $X=8.315 $Y=0.82
+ $X2=8.17 $Y2=0.735
r145 27 32 2.5345 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=8.865 $Y=0.82
+ $X2=9.005 $Y2=0.82
r146 27 28 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=8.865 $Y=0.82
+ $X2=8.315 $Y2=0.82
r147 23 30 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=8.865 $Y=1.6
+ $X2=8.95 $Y2=1.495
r148 23 25 37.7619 $w=2.08e-07 $l=7.15e-07 $layer=LI1_cond $X=8.865 $Y=1.6
+ $X2=8.15 $Y2=1.6
r149 19 40 3.57235 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.14 $Y=0.595
+ $X2=5.14 $Y2=0.43
r150 19 21 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=5.14 $Y=0.595
+ $X2=5.14 $Y2=1.94
r151 16 35 44.9977 $w=3.9e-07 $l=3.04138e-07 $layer=POLY_cond $X=8.855 $Y=1.41
+ $X2=8.975 $Y2=1.16
r152 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.855 $Y=1.41
+ $X2=8.855 $Y2=1.985
r153 13 35 39.3952 $w=3.9e-07 $l=2.26164e-07 $layer=POLY_cond $X=8.83 $Y=0.995
+ $X2=8.975 $Y2=1.16
r154 13 15 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.83 $Y=0.995
+ $X2=8.83 $Y2=0.555
r155 4 25 600 $w=1.7e-07 $l=2.42178e-07 $layer=licon1_PDIFF $count=1 $X=7.92
+ $Y=1.645 $X2=8.15 $Y2=1.62
r156 3 21 600 $w=1.7e-07 $l=5.13712e-07 $layer=licon1_PDIFF $count=1 $X=5.015
+ $Y=1.485 $X2=5.14 $Y2=1.94
r157 2 44 182 $w=1.7e-07 $l=4.8775e-07 $layer=licon1_NDIFF $count=1 $X=7.93
+ $Y=0.235 $X2=8.15 $Y2=0.625
r158 1 40 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=5.175
+ $Y=0.245 $X2=5.3 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_2%VPWR 1 2 3 4 13 15 21 25 29 32 33 34 36 48
+ 54 55 61 64
r97 64 65 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r98 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r99 55 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=8.51 $Y2=2.72
r100 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r101 52 64 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=8.79 $Y=2.72
+ $X2=8.622 $Y2=2.72
r102 52 54 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=8.79 $Y=2.72
+ $X2=9.43 $Y2=2.72
r103 51 65 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=8.51 $Y2=2.72
r104 50 51 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r105 48 64 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=8.455 $Y=2.72
+ $X2=8.622 $Y2=2.72
r106 48 50 266.508 $w=1.68e-07 $l=4.085e-06 $layer=LI1_cond $X=8.455 $Y=2.72
+ $X2=4.37 $Y2=2.72
r107 47 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r108 46 47 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r109 44 47 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=3.91 $Y2=2.72
r110 44 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r111 43 46 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=3.91 $Y2=2.72
r112 43 44 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r113 41 61 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.43 $Y=2.72
+ $X2=1.237 $Y2=2.72
r114 41 43 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.43 $Y=2.72
+ $X2=1.61 $Y2=2.72
r115 40 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r116 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r117 37 58 4.42505 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=2.72
+ $X2=0.187 $Y2=2.72
r118 37 39 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.375 $Y=2.72
+ $X2=0.69 $Y2=2.72
r119 36 61 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=1.045 $Y=2.72
+ $X2=1.237 $Y2=2.72
r120 36 39 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.045 $Y=2.72
+ $X2=0.69 $Y2=2.72
r121 34 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r122 34 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r123 32 46 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.935 $Y=2.72
+ $X2=3.91 $Y2=2.72
r124 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.935 $Y=2.72
+ $X2=4.1 $Y2=2.72
r125 31 50 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.265 $Y=2.72
+ $X2=4.37 $Y2=2.72
r126 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.265 $Y=2.72
+ $X2=4.1 $Y2=2.72
r127 27 64 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=8.622 $Y=2.635
+ $X2=8.622 $Y2=2.72
r128 27 29 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=8.622 $Y=2.635
+ $X2=8.622 $Y2=2.36
r129 23 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.1 $Y=2.635 $X2=4.1
+ $Y2=2.72
r130 23 25 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.1 $Y=2.635
+ $X2=4.1 $Y2=2.32
r131 19 61 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.237 $Y=2.635
+ $X2=1.237 $Y2=2.72
r132 19 21 10.0278 $w=3.83e-07 $l=3.35e-07 $layer=LI1_cond $X=1.237 $Y=2.635
+ $X2=1.237 $Y2=2.3
r133 15 18 27.0228 $w=2.88e-07 $l=6.8e-07 $layer=LI1_cond $X=0.23 $Y=1.66
+ $X2=0.23 $Y2=2.34
r134 13 58 3.0128 $w=2.9e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.23 $Y=2.635
+ $X2=0.187 $Y2=2.72
r135 13 18 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.23 $Y=2.635
+ $X2=0.23 $Y2=2.34
r136 4 29 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=8.475
+ $Y=1.485 $X2=8.62 $Y2=2.36
r137 3 25 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.975
+ $Y=2.175 $X2=4.1 $Y2=2.32
r138 2 21 600 $w=1.7e-07 $l=9.05028e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.265 $Y2=2.3
r139 1 18 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r140 1 15 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_2%X 1 2 7 10
r14 10 13 38.1747 $w=3.18e-07 $l=1.06e-06 $layer=LI1_cond $X=0.705 $Y=0.56
+ $X2=0.705 $Y2=1.62
r15 7 17 15.486 $w=3.18e-07 $l=4.3e-07 $layer=LI1_cond $X=0.705 $Y=1.87
+ $X2=0.705 $Y2=2.3
r16 7 13 9.00346 $w=3.18e-07 $l=2.5e-07 $layer=LI1_cond $X=0.705 $Y=1.87
+ $X2=0.705 $Y2=1.62
r17 2 17 400 $w=1.7e-07 $l=8.937e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.75 $Y2=2.3
r18 2 13 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.75 $Y2=1.62
r19 1 10 182 $w=1.7e-07 $l=4.1503e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.75 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_2%A_453_325# 1 2 3 4 13 17 22 24 25 28 29 30
+ 32 35 39 43 45 46 48
c155 29 0 1.36535e-19 $X=5.395 $Y=2.36
r156 46 47 17.602 $w=2.01e-07 $l=2.9e-07 $layer=LI1_cond $X=5.48 $Y=0.772
+ $X2=5.77 $Y2=0.772
r157 41 43 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.93 $Y=1.12
+ $X2=4.04 $Y2=1.12
r158 37 47 1.71937 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=5.77 $Y=0.655
+ $X2=5.77 $Y2=0.772
r159 37 39 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=5.77 $Y=0.655
+ $X2=5.77 $Y2=0.545
r160 33 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=2.36
+ $X2=5.48 $Y2=2.36
r161 33 35 131.786 $w=1.68e-07 $l=2.02e-06 $layer=LI1_cond $X=5.565 $Y=2.36
+ $X2=7.585 $Y2=2.36
r162 32 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=2.275
+ $X2=5.48 $Y2=2.36
r163 31 46 1.71937 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=5.48 $Y=0.89
+ $X2=5.48 $Y2=0.772
r164 31 32 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=5.48 $Y=0.89
+ $X2=5.48 $Y2=2.275
r165 29 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=2.36
+ $X2=5.48 $Y2=2.36
r166 29 30 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=5.395 $Y=2.36
+ $X2=4.87 $Y2=2.36
r167 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.785 $Y=2.275
+ $X2=4.87 $Y2=2.36
r168 27 28 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.785 $Y=2.065
+ $X2=4.785 $Y2=2.275
r169 26 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.125 $Y=1.98
+ $X2=4.04 $Y2=1.98
r170 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.7 $Y=1.98
+ $X2=4.785 $Y2=2.065
r171 25 26 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=4.7 $Y=1.98
+ $X2=4.125 $Y2=1.98
r172 24 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=1.895
+ $X2=4.04 $Y2=1.98
r173 23 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=1.205
+ $X2=4.04 $Y2=1.12
r174 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.04 $Y=1.205
+ $X2=4.04 $Y2=1.895
r175 22 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.93 $Y=1.035
+ $X2=3.93 $Y2=1.12
r176 21 22 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.93 $Y=0.455
+ $X2=3.93 $Y2=1.035
r177 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.845 $Y=0.37
+ $X2=3.93 $Y2=0.455
r178 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.845 $Y=0.37
+ $X2=3.55 $Y2=0.37
r179 13 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.955 $Y=1.98
+ $X2=4.04 $Y2=1.98
r180 13 15 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=3.955 $Y=1.98
+ $X2=2.455 $Y2=1.98
r181 4 35 600 $w=1.7e-07 $l=8.56081e-07 $layer=licon1_PDIFF $count=1 $X=7.275
+ $Y=1.645 $X2=7.585 $Y2=2.36
r182 3 15 600 $w=1.7e-07 $l=4.39858e-07 $layer=licon1_PDIFF $count=1 $X=2.265
+ $Y=1.625 $X2=2.455 $Y2=1.98
r183 2 39 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=5.635
+ $Y=0.245 $X2=5.77 $Y2=0.545
r184 1 19 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=3.295
+ $Y=0.245 $X2=3.55 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_2%A_477_49# 1 2 3 4 13 16 17 19 21 24 26 27
+ 29 34 35 36 37 40 43
c136 29 0 1.24749e-19 $X=7.43 $Y=0.38
c137 16 0 2.74598e-20 $X=3.59 $Y=1.375
r138 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.15 $Y=1.53
+ $X2=6.15 $Y2=1.53
r139 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.7 $Y=1.53 $X2=3.7
+ $Y2=1.53
r140 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.845 $Y=1.53
+ $X2=3.7 $Y2=1.53
r141 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.005 $Y=1.53
+ $X2=6.15 $Y2=1.53
r142 36 37 2.67326 $w=1.4e-07 $l=2.16e-06 $layer=MET1_cond $X=6.005 $Y=1.53
+ $X2=3.845 $Y2=1.53
r143 32 34 10.6148 $w=2.78e-07 $l=2.15e-07 $layer=LI1_cond $X=2.52 $Y=0.765
+ $X2=2.735 $Y2=0.765
r144 27 35 11.5258 $w=2.08e-07 $l=2.1e-07 $layer=LI1_cond $X=7.345 $Y=0.36
+ $X2=7.135 $Y2=0.36
r145 27 29 4.48918 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=7.345 $Y=0.36
+ $X2=7.43 $Y2=0.36
r146 26 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.625 $Y=0.34
+ $X2=7.135 $Y2=0.34
r147 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.54 $Y=0.425
+ $X2=6.625 $Y2=0.34
r148 23 24 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.54 $Y=0.425
+ $X2=6.54 $Y2=1.445
r149 22 44 6.03523 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=6.21 $Y=1.53
+ $X2=6.002 $Y2=1.53
r150 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.455 $Y=1.53
+ $X2=6.54 $Y2=1.445
r151 21 22 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.455 $Y=1.53
+ $X2=6.21 $Y2=1.53
r152 17 44 2.46632 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=6.002 $Y=1.615
+ $X2=6.002 $Y2=1.53
r153 17 19 0.138849 $w=4.13e-07 $l=5e-09 $layer=LI1_cond $X=6.002 $Y=1.615
+ $X2=6.002 $Y2=1.62
r154 16 40 8.59825 $w=3.35e-07 $l=1.55997e-07 $layer=LI1_cond $X=3.59 $Y=1.375
+ $X2=3.592 $Y2=1.53
r155 15 16 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.59 $Y=0.795
+ $X2=3.59 $Y2=1.375
r156 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.505 $Y=0.71
+ $X2=3.59 $Y2=0.795
r157 13 34 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.505 $Y=0.71
+ $X2=2.735 $Y2=0.71
r158 4 19 300 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_PDIFF $count=2 $X=5.625
+ $Y=1.485 $X2=5.97 $Y2=1.62
r159 3 40 600 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=3.315
+ $Y=1.485 $X2=3.565 $Y2=1.61
r160 2 29 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=7.235
+ $Y=0.245 $X2=7.43 $Y2=0.38
r161 1 32 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.385
+ $Y=0.245 $X2=2.52 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_2%A_1286_297# 1 2 3 4 15 20 23 26 29 31 36
c67 4 0 1.20335e-19 $X=8.945 $Y=1.485
r68 34 36 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=9.27 $Y=0.42 $X2=9.4
+ $Y2=0.42
r69 28 29 17.3428 $w=2.28e-07 $l=3.3e-07 $layer=LI1_cond $X=9.28 $Y=1.99
+ $X2=8.95 $Y2=1.99
r70 26 31 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.4 $Y=1.875 $X2=9.4
+ $Y2=1.99
r71 25 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.4 $Y=0.585 $X2=9.4
+ $Y2=0.42
r72 25 26 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=9.4 $Y=0.585
+ $X2=9.4 $Y2=1.875
r73 21 31 3.15669 $w=2.28e-07 $l=6.3e-08 $layer=LI1_cond $X=9.337 $Y=1.99
+ $X2=9.4 $Y2=1.99
r74 21 28 2.85605 $w=2.28e-07 $l=5.7e-08 $layer=LI1_cond $X=9.337 $Y=1.99
+ $X2=9.28 $Y2=1.99
r75 21 23 7.61784 $w=2.93e-07 $l=1.95e-07 $layer=LI1_cond $X=9.337 $Y=2.105
+ $X2=9.337 $Y2=2.3
r76 20 29 129.503 $w=1.68e-07 $l=1.985e-06 $layer=LI1_cond $X=6.965 $Y=2.02
+ $X2=8.95 $Y2=2.02
r77 15 18 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=6.88 $Y=0.76
+ $X2=6.88 $Y2=1.865
r78 13 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.88 $Y=1.935
+ $X2=6.965 $Y2=2.02
r79 13 18 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=6.88 $Y=1.935 $X2=6.88
+ $Y2=1.865
r80 4 28 600 $w=1.7e-07 $l=6.20282e-07 $layer=licon1_PDIFF $count=1 $X=8.945
+ $Y=1.485 $X2=9.28 $Y2=1.96
r81 4 23 600 $w=1.7e-07 $l=9.6601e-07 $layer=licon1_PDIFF $count=1 $X=8.945
+ $Y=1.485 $X2=9.275 $Y2=2.3
r82 3 18 600 $w=1.7e-07 $l=6.11146e-07 $layer=licon1_PDIFF $count=1 $X=6.43
+ $Y=1.485 $X2=6.88 $Y2=1.865
r83 2 34 182 $w=1.7e-07 $l=4.48051e-07 $layer=licon1_NDIFF $count=1 $X=8.905
+ $Y=0.235 $X2=9.27 $Y2=0.42
r84 1 15 182 $w=1.7e-07 $l=7.01302e-07 $layer=licon1_NDIFF $count=1 $X=6.44
+ $Y=0.245 $X2=6.88 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_2%VGND 1 2 3 4 13 15 19 23 27 30 31 33 34 35
+ 37 56 57 63
c108 57 0 1.70967e-19 $X=9.43 $Y=0
r109 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r110 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r111 54 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=9.43
+ $Y2=0
r112 53 54 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r113 51 54 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=4.37 $Y=0 $X2=8.51
+ $Y2=0
r114 50 53 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=4.37 $Y=0 $X2=8.51
+ $Y2=0
r115 50 51 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r116 48 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r117 47 48 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r118 45 48 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=3.91
+ $Y2=0
r119 45 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r120 44 47 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=3.91
+ $Y2=0
r121 44 45 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r122 42 63 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.325 $Y=0 $X2=1.18
+ $Y2=0
r123 42 44 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.325 $Y=0
+ $X2=1.61 $Y2=0
r124 41 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r125 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r126 38 60 4.42505 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=0
+ $X2=0.187 $Y2=0
r127 38 40 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.375 $Y=0
+ $X2=0.69 $Y2=0
r128 37 63 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.18
+ $Y2=0
r129 37 40 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r130 35 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r131 35 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r132 33 53 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=8.535 $Y=0 $X2=8.51
+ $Y2=0
r133 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.535 $Y=0 $X2=8.62
+ $Y2=0
r134 32 56 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=8.705 $Y=0
+ $X2=9.43 $Y2=0
r135 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.705 $Y=0 $X2=8.62
+ $Y2=0
r136 30 47 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.185 $Y=0
+ $X2=3.91 $Y2=0
r137 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.185 $Y=0 $X2=4.27
+ $Y2=0
r138 29 50 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.37
+ $Y2=0
r139 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.27
+ $Y2=0
r140 25 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.62 $Y=0.085
+ $X2=8.62 $Y2=0
r141 25 27 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.62 $Y=0.085
+ $X2=8.62 $Y2=0.4
r142 21 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=0.085
+ $X2=4.27 $Y2=0
r143 21 23 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.27 $Y=0.085
+ $X2=4.27 $Y2=0.36
r144 17 63 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0
r145 17 19 10.9283 $w=2.88e-07 $l=2.75e-07 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0.36
r146 13 60 3.0128 $w=2.9e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.23 $Y=0.085
+ $X2=0.187 $Y2=0
r147 13 15 18.8762 $w=2.88e-07 $l=4.75e-07 $layer=LI1_cond $X=0.23 $Y=0.085
+ $X2=0.23 $Y2=0.56
r148 4 27 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=8.485
+ $Y=0.235 $X2=8.62 $Y2=0.4
r149 3 23 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=4.115
+ $Y=0.235 $X2=4.27 $Y2=0.36
r150 2 19 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.24 $Y2=0.36
r151 1 15 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

