* File: sky130_fd_sc_hdll__diode_8.pex.spice
* Created: Wed Sep  2 08:29:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__DIODE_8%DIODE 1 4 10 58
r7 56 58 3.75385 $w=2.208e-06 $l=6.8e-07 $layer=LI1_cond $X=2.69 $Y=1.36
+ $X2=3.37 $Y2=1.36
r8 54 56 1.87692 $w=2.208e-06 $l=3.4e-07 $layer=LI1_cond $X=2.35 $Y=1.36
+ $X2=2.69 $Y2=1.36
r9 52 54 3.61584 $w=2.208e-06 $l=6.55e-07 $layer=LI1_cond $X=1.695 $Y=1.36
+ $X2=2.35 $Y2=1.36
r10 50 52 0.138009 $w=2.208e-06 $l=2.5e-08 $layer=LI1_cond $X=1.67 $Y=1.36
+ $X2=1.695 $Y2=1.36
r11 48 50 1.87692 $w=2.208e-06 $l=3.4e-07 $layer=LI1_cond $X=1.33 $Y=1.36
+ $X2=1.67 $Y2=1.36
r12 46 48 1.87692 $w=2.208e-06 $l=3.4e-07 $layer=LI1_cond $X=0.99 $Y=1.36
+ $X2=1.33 $Y2=1.36
r13 10 46 1.65611 $w=2.208e-06 $l=3e-07 $layer=LI1_cond $X=0.69 $Y=1.36 $X2=0.99
+ $Y2=1.36
r14 10 37 2.09774 $w=2.208e-06 $l=3.8e-07 $layer=LI1_cond $X=0.69 $Y=1.36
+ $X2=0.31 $Y2=1.36
r15 4 37 0.441629 $w=2.208e-06 $l=8e-08 $layer=LI1_cond $X=0.23 $Y=1.36 $X2=0.31
+ $Y2=1.36
r16 1 58 60.6667 $w=1.7e-07 $l=3.32135e-06 $layer=licon1_NDIFF $count=3 $X=0.135
+ $Y=0.195 $X2=3.37 $Y2=0.37
r17 1 56 60.6667 $w=1.7e-07 $l=2.64105e-06 $layer=licon1_NDIFF $count=3 $X=0.135
+ $Y=0.195 $X2=2.69 $Y2=0.37
r18 1 54 45.5 $w=1.7e-07 $l=2.45905e-06 $layer=licon1_NDIFF $count=4 $X=0.135
+ $Y=0.195 $X2=2.35 $Y2=0.71
r19 1 52 45.5 $w=1.7e-07 $l=2.07311e-06 $layer=licon1_NDIFF $count=4 $X=0.135
+ $Y=0.195 $X2=1.695 $Y2=1.39
r20 1 50 45.5 $w=1.7e-07 $l=1.62014e-06 $layer=licon1_NDIFF $count=4 $X=0.135
+ $Y=0.195 $X2=1.67 $Y2=0.37
r21 1 48 45.5 $w=1.7e-07 $l=1.42949e-06 $layer=licon1_NDIFF $count=4 $X=0.135
+ $Y=0.195 $X2=1.33 $Y2=0.71
r22 1 46 60.6667 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_NDIFF $count=3 $X=0.135
+ $Y=0.195 $X2=0.99 $Y2=0.37
r23 1 37 60.6667 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_NDIFF $count=3 $X=0.135
+ $Y=0.195 $X2=0.31 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HDLL__DIODE_8%VGND 1 8 9
r5 8 9 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r6 4 8 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=3.45
+ $Y2=0
r7 1 9 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=3.45
+ $Y2=0
r8 1 4 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HDLL__DIODE_8%VPWR 1 8 9
r5 8 9 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.45 $Y=2.72 $X2=3.45
+ $Y2=2.72
r6 4 8 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=0.23 $Y=2.72 $X2=3.45
+ $Y2=2.72
r7 1 9 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=0.23 $Y=2.72 $X2=3.45
+ $Y2=2.72
r8 1 4 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
.ends

