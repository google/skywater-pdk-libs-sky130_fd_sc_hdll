* File: sky130_fd_sc_hdll__a211o_4.spice
* Created: Wed Sep  2 08:15:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a211o_4.pex.spice"
.subckt sky130_fd_sc_hdll__a211o_4  VNB VPB B1 C1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* C1	C1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1001 N_X_M1001_d N_A_79_204#_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.20475 PD=0.98 PS=1.93 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75005.9 A=0.0975 P=1.6 MULT=1
MM1004 N_X_M1001_d N_A_79_204#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75000.7
+ SB=75005.4 A=0.0975 P=1.6 MULT=1
MM1005 N_X_M1005_d N_A_79_204#_M1005_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.128375 AS=0.10725 PD=1.045 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1011 N_X_M1005_d N_A_79_204#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.128375 AS=0.108875 PD=1.045 PS=0.985 NRD=11.988 NRS=0.912 M=1 R=4.33333
+ SA=75001.7 SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1007 N_A_79_204#_M1007_d N_B1_M1007_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.108875 PD=0.97 PS=0.985 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75002.2
+ SB=75003.9 A=0.0975 P=1.6 MULT=1
MM1012 N_A_79_204#_M1007_d N_C1_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.141375 PD=0.97 PS=1.085 NRD=7.38 NRS=11.988 M=1 R=4.33333
+ SA=75002.7 SB=75003.4 A=0.0975 P=1.6 MULT=1
MM1023 N_A_79_204#_M1023_d N_C1_M1023_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.143 AS=0.141375 PD=1.09 PS=1.085 NRD=11.076 NRS=16.608 M=1 R=4.33333
+ SA=75003.3 SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1013 N_A_79_204#_M1023_d N_B1_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.143 AS=0.156 PD=1.09 PS=1.13 NRD=18.456 NRS=7.38 M=1 R=4.33333 SA=75003.9
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1013_s N_A2_M1002_g A_1051_47# VNB NSHORT L=0.15 W=0.65 AD=0.156
+ AS=0.091 PD=1.13 PS=0.93 NRD=29.532 NRS=15.684 M=1 R=4.33333 SA=75004.5
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1016 A_1051_47# N_A1_M1016_g N_A_79_204#_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.1235 PD=0.93 PS=1.03 NRD=15.684 NRS=9.228 M=1 R=4.33333
+ SA=75004.9 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1014 A_1243_47# N_A1_M1014_g N_A_79_204#_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.1235 PD=0.93 PS=1.03 NRD=15.684 NRS=9.228 M=1 R=4.33333
+ SA=75005.5 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1019_d N_A2_M1019_g A_1243_47# VNB NSHORT L=0.15 W=0.65 AD=0.2015
+ AS=0.091 PD=1.92 PS=0.93 NRD=8.304 NRS=15.684 M=1 R=4.33333 SA=75005.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_79_204#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.15 PD=2.54 PS=1.3 NRD=0.9653 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A_79_204#_M1009_g N_X_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1009_d N_A_79_204#_M1010_g N_X_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.1
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1020 N_VPWR_M1020_d N_A_79_204#_M1020_g N_X_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.15 PD=2.54 PS=1.3 NRD=0.9653 NRS=1.9503 M=1 R=5.55556 SA=90001.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1017 N_A_523_297#_M1017_d N_B1_M1017_g A_613_297# VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.15 PD=2.54 PS=1.3 NRD=0.9653 NRS=18.6953 M=1 R=5.55556 SA=90000.2
+ SB=90003.8 A=0.18 P=2.36 MULT=1
MM1006 A_613_297# N_C1_M1006_g N_A_79_204#_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=18.6953 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90003.3 A=0.18 P=2.36 MULT=1
MM1022 A_805_297# N_C1_M1022_g N_A_79_204#_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.17 AS=0.15 PD=1.34 PS=1.3 NRD=22.6353 NRS=1.9503 M=1 R=5.55556 SA=90001.1
+ SB=90002.8 A=0.18 P=2.36 MULT=1
MM1015 N_A_523_297#_M1015_d N_B1_M1015_g A_805_297# VPB PHIGHVT L=0.18 W=1
+ AD=0.205 AS=0.17 PD=1.41 PS=1.34 NRD=9.8303 NRS=22.6353 M=1 R=5.55556
+ SA=90001.7 SB=90002.3 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_A2_M1000_g N_A_523_297#_M1015_d VPB PHIGHVT L=0.18 W=1
+ AD=0.205 AS=0.205 PD=1.41 PS=1.41 NRD=1.9503 NRS=15.7403 M=1 R=5.55556
+ SA=90002.2 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1000_d N_A1_M1008_g N_A_523_297#_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.205 AS=0.15 PD=1.41 PS=1.3 NRD=23.6203 NRS=1.9503 M=1 R=5.55556
+ SA=90002.8 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1018_d N_A1_M1018_g N_A_523_297#_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90003.3
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1021 N_VPWR_M1018_d N_A2_M1021_g N_A_523_297#_M1021_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.27 PD=1.3 PS=2.54 NRD=1.9503 NRS=0.9653 M=1 R=5.55556 SA=90003.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX24_noxref VNB VPB NWDIODE A=12.4227 P=18.69
pX25_noxref noxref_16 C1 C1 PROBETYPE=1
pX26_noxref noxref_17 B1 B1 PROBETYPE=1
pX27_noxref noxref_18 A1 A1 PROBETYPE=1
pX28_noxref noxref_19 A2 A2 PROBETYPE=1
c_92 VPB 0 2.78086e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__a211o_4.pxi.spice"
*
.ends
*
*
