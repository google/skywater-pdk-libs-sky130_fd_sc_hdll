* File: sky130_fd_sc_hdll__or3b_2.spice
* Created: Wed Sep  2 08:48:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or3b_2.pex.spice"
.subckt sky130_fd_sc_hdll__or3b_2  VNB VPB C_N A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_C_N_M1009_g N_A_27_47#_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0787009 AS=0.1302 PD=0.773271 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_186_21#_M1001_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.170625 AS=0.121799 PD=1.175 PS=1.19673 NRD=8.304 NRS=11.076 M=1 R=4.33333
+ SA=75000.5 SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1011 N_X_M1001_d N_A_186_21#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.170625 AS=0.139264 PD=1.175 PS=1.28178 NRD=36.912 NRS=10.152 M=1
+ R=4.33333 SA=75001.2 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1005 N_A_186_21#_M1005_d N_A_M1005_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.089986 PD=0.7 PS=0.828224 NRD=0 NRS=19.992 M=1 R=2.8 SA=75001.9
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_B_M1002_g N_A_186_21#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.063 AS=0.0588 PD=0.72 PS=0.7 NRD=7.14 NRS=0 M=1 R=2.8 SA=75002.3
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_A_186_21#_M1003_d N_A_27_47#_M1003_g N_VGND_M1002_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.063 PD=1.36 PS=0.72 NRD=0 NRS=0 M=1 R=2.8 SA=75002.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_C_N_M1006_g N_A_27_47#_M1006_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0904183 AS=0.1134 PD=0.801549 PS=1.38 NRD=75.1752 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1007 N_VPWR_M1006_d N_A_186_21#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.215282 AS=0.2 PD=1.90845 PS=1.4 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.4 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1010_d N_A_186_21#_M1010_g N_X_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.218803 AS=0.2 PD=1.91549 PS=1.4 NRD=1.9503 NRS=22.6353 M=1 R=5.55556
+ SA=90001 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1000 A_448_297# N_A_M1000_g N_VPWR_M1010_d VPB PHIGHVT L=0.18 W=0.42 AD=0.0651
+ AS=0.0918972 PD=0.73 PS=0.804507 NRD=46.886 NRS=76.83 M=1 R=2.33333 SA=90001.4
+ SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1004 A_546_297# N_B_M1004_g A_448_297# VPB PHIGHVT L=0.18 W=0.42 AD=0.0567
+ AS=0.0651 PD=0.69 PS=0.73 NRD=37.5088 NRS=46.886 M=1 R=2.33333 SA=90001.9
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1008 N_A_186_21#_M1008_d N_A_27_47#_M1008_g A_546_297# VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.0567 PD=1.38 PS=0.69 NRD=2.3443 NRS=37.5088 M=1
+ R=2.33333 SA=90002.4 SB=90000.2 A=0.0756 P=1.2 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
pX13_noxref noxref_13 X X PROBETYPE=1
pX14_noxref noxref_14 A A PROBETYPE=1
pX15_noxref noxref_15 B B PROBETYPE=1
c_40 VNB 0 1.58571e-19 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hdll__or3b_2.pxi.spice"
*
.ends
*
*
