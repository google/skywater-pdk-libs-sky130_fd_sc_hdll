* File: sky130_fd_sc_hdll__a211o_2.pxi.spice
* Created: Thu Aug 27 18:51:30 2020
* 
x_PM_SKY130_FD_SC_HDLL__A211O_2%A_79_21# N_A_79_21#_M1010_d N_A_79_21#_M1005_d
+ N_A_79_21#_M1009_d N_A_79_21#_c_54_n N_A_79_21#_M1008_g N_A_79_21#_c_60_n
+ N_A_79_21#_M1000_g N_A_79_21#_c_55_n N_A_79_21#_M1011_g N_A_79_21#_c_61_n
+ N_A_79_21#_M1006_g N_A_79_21#_c_56_n N_A_79_21#_c_70_p N_A_79_21#_c_130_p
+ N_A_79_21#_c_63_n N_A_79_21#_c_64_n N_A_79_21#_c_71_p N_A_79_21#_c_57_n
+ N_A_79_21#_c_58_n N_A_79_21#_c_65_n N_A_79_21#_c_82_p N_A_79_21#_c_59_n
+ PM_SKY130_FD_SC_HDLL__A211O_2%A_79_21#
x_PM_SKY130_FD_SC_HDLL__A211O_2%A2 N_A2_c_159_n N_A2_M1007_g N_A2_c_156_n
+ N_A2_M1003_g A2 N_A2_c_158_n PM_SKY130_FD_SC_HDLL__A211O_2%A2
x_PM_SKY130_FD_SC_HDLL__A211O_2%A1 N_A1_c_189_n N_A1_M1010_g N_A1_c_190_n
+ N_A1_M1004_g A1 A1 PM_SKY130_FD_SC_HDLL__A211O_2%A1
x_PM_SKY130_FD_SC_HDLL__A211O_2%B1 N_B1_c_219_n N_B1_M1002_g N_B1_c_220_n
+ N_B1_M1001_g B1 B1 PM_SKY130_FD_SC_HDLL__A211O_2%B1
x_PM_SKY130_FD_SC_HDLL__A211O_2%C1 N_C1_c_246_n N_C1_M1005_g N_C1_c_247_n
+ N_C1_M1009_g C1 PM_SKY130_FD_SC_HDLL__A211O_2%C1
x_PM_SKY130_FD_SC_HDLL__A211O_2%VPWR N_VPWR_M1000_d N_VPWR_M1006_d
+ N_VPWR_M1007_d N_VPWR_c_269_n N_VPWR_c_270_n N_VPWR_c_271_n N_VPWR_c_272_n
+ N_VPWR_c_273_n N_VPWR_c_274_n N_VPWR_c_275_n VPWR N_VPWR_c_276_n
+ N_VPWR_c_268_n N_VPWR_c_278_n PM_SKY130_FD_SC_HDLL__A211O_2%VPWR
x_PM_SKY130_FD_SC_HDLL__A211O_2%X N_X_M1008_s N_X_M1000_s X N_X_c_321_n
+ PM_SKY130_FD_SC_HDLL__A211O_2%X
x_PM_SKY130_FD_SC_HDLL__A211O_2%A_319_297# N_A_319_297#_M1007_s
+ N_A_319_297#_M1004_d N_A_319_297#_c_339_n N_A_319_297#_c_336_n
+ N_A_319_297#_c_341_n PM_SKY130_FD_SC_HDLL__A211O_2%A_319_297#
x_PM_SKY130_FD_SC_HDLL__A211O_2%VGND N_VGND_M1008_d N_VGND_M1011_d
+ N_VGND_M1002_d N_VGND_c_364_n N_VGND_c_365_n N_VGND_c_366_n N_VGND_c_367_n
+ N_VGND_c_368_n VGND N_VGND_c_369_n N_VGND_c_370_n N_VGND_c_371_n
+ N_VGND_c_372_n PM_SKY130_FD_SC_HDLL__A211O_2%VGND
cc_1 VNB N_A_79_21#_c_54_n 0.022136f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1
cc_2 VNB N_A_79_21#_c_55_n 0.0188964f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=0.995
cc_3 VNB N_A_79_21#_c_56_n 0.00468317f $X=-0.19 $Y=-0.24 $X2=1.185 $Y2=1.16
cc_4 VNB N_A_79_21#_c_57_n 0.00815748f $X=-0.19 $Y=-0.24 $X2=3.555 $Y2=0.785
cc_5 VNB N_A_79_21#_c_58_n 0.0167856f $X=-0.19 $Y=-0.24 $X2=3.77 $Y2=0.4
cc_6 VNB N_A_79_21#_c_59_n 0.0644226f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_7 VNB N_A2_c_156_n 0.0201403f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB A2 0.00305046f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A2_c_158_n 0.034931f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_10 VNB N_A1_c_189_n 0.0173247f $X=-0.19 $Y=-0.24 $X2=2.5 $Y2=0.235
cc_11 VNB N_A1_c_190_n 0.0236079f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB A1 0.00450648f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_B1_c_219_n 0.0186029f $X=-0.19 $Y=-0.24 $X2=2.5 $Y2=0.235
cc_14 VNB N_B1_c_220_n 0.0242757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB B1 0.00196466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_C1_c_246_n 0.0232607f $X=-0.19 $Y=-0.24 $X2=2.5 $Y2=0.235
cc_17 VNB N_C1_c_247_n 0.0260998f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB C1 0.0119145f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_268_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_X_c_321_n 0.0017876f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1
cc_21 VNB N_VGND_c_364_n 0.0107461f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1
cc_22 VNB N_VGND_c_365_n 0.035483f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_23 VNB N_VGND_c_366_n 0.00528059f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=0.995
cc_24 VNB N_VGND_c_367_n 0.0353556f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_25 VNB N_VGND_c_368_n 0.00526062f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_26 VNB N_VGND_c_369_n 0.02207f $X=-0.19 $Y=-0.24 $X2=2.855 $Y2=0.785
cc_27 VNB N_VGND_c_370_n 0.223067f $X=-0.19 $Y=-0.24 $X2=3.745 $Y2=0.695
cc_28 VNB N_VGND_c_371_n 0.0164684f $X=-0.19 $Y=-0.24 $X2=2.665 $Y2=0.785
cc_29 VNB N_VGND_c_372_n 0.0187377f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VPB N_A_79_21#_c_60_n 0.021062f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_31 VPB N_A_79_21#_c_61_n 0.0191132f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_32 VPB N_A_79_21#_c_56_n 0.00360556f $X=-0.19 $Y=1.305 $X2=1.185 $Y2=1.16
cc_33 VPB N_A_79_21#_c_63_n 0.019502f $X=-0.19 $Y=1.305 $X2=3.555 $Y2=1.575
cc_34 VPB N_A_79_21#_c_64_n 4.43773e-19 $X=-0.19 $Y=1.305 $X2=1.355 $Y2=1.575
cc_35 VPB N_A_79_21#_c_65_n 0.026497f $X=-0.19 $Y=1.305 $X2=3.77 $Y2=1.755
cc_36 VPB N_A_79_21#_c_59_n 0.034891f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_37 VPB N_A2_c_159_n 0.020729f $X=-0.19 $Y=1.305 $X2=2.5 $Y2=0.235
cc_38 VPB N_A2_c_158_n 0.0157302f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_39 VPB N_A1_c_190_n 0.028949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_B1_c_220_n 0.0269388f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_C1_c_247_n 0.0321792f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_269_n 0.0107202f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1
cc_43 VPB N_VPWR_c_270_n 0.0442199f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_44 VPB N_VPWR_c_271_n 0.0210262f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=0.995
cc_45 VPB N_VPWR_c_272_n 0.0114873f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_46 VPB N_VPWR_c_273_n 0.00533487f $X=-0.19 $Y=1.305 $X2=1.227 $Y2=1.16
cc_47 VPB N_VPWR_c_274_n 0.0208444f $X=-0.19 $Y=1.305 $X2=2.475 $Y2=0.785
cc_48 VPB N_VPWR_c_275_n 0.00526085f $X=-0.19 $Y=1.305 $X2=1.355 $Y2=0.785
cc_49 VPB N_VPWR_c_276_n 0.049526f $X=-0.19 $Y=1.305 $X2=3.77 $Y2=0.4
cc_50 VPB N_VPWR_c_268_n 0.0568628f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_278_n 0.00487897f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.202
cc_52 VPB N_X_c_321_n 0.00255477f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1
cc_53 VPB N_A_319_297#_c_336_n 0.00634949f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_54 N_A_79_21#_c_56_n N_A2_c_159_n 0.00192835f $X=1.185 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_55 N_A_79_21#_c_63_n N_A2_c_159_n 0.0163834f $X=3.555 $Y=1.575 $X2=-0.19
+ $Y2=-0.24
cc_56 N_A_79_21#_c_56_n N_A2_c_156_n 0.00273656f $X=1.185 $Y=1.16 $X2=0 $Y2=0
cc_57 N_A_79_21#_c_70_p N_A2_c_156_n 0.016311f $X=2.475 $Y=0.785 $X2=0 $Y2=0
cc_58 N_A_79_21#_c_71_p N_A2_c_156_n 0.00207051f $X=2.69 $Y=0.36 $X2=0 $Y2=0
cc_59 N_A_79_21#_c_56_n A2 0.0191079f $X=1.185 $Y=1.16 $X2=0 $Y2=0
cc_60 N_A_79_21#_c_70_p A2 0.0296095f $X=2.475 $Y=0.785 $X2=0 $Y2=0
cc_61 N_A_79_21#_c_63_n A2 0.0246685f $X=3.555 $Y=1.575 $X2=0 $Y2=0
cc_62 N_A_79_21#_c_59_n A2 7.7121e-19 $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_63 N_A_79_21#_c_56_n N_A2_c_158_n 0.00491009f $X=1.185 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_79_21#_c_70_p N_A2_c_158_n 0.0082533f $X=2.475 $Y=0.785 $X2=0 $Y2=0
cc_65 N_A_79_21#_c_63_n N_A2_c_158_n 0.00668061f $X=3.555 $Y=1.575 $X2=0 $Y2=0
cc_66 N_A_79_21#_c_59_n N_A2_c_158_n 0.0143728f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_67 N_A_79_21#_c_70_p N_A1_c_189_n 0.0086724f $X=2.475 $Y=0.785 $X2=-0.19
+ $Y2=-0.24
cc_68 N_A_79_21#_c_71_p N_A1_c_189_n 0.0077727f $X=2.69 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_69 N_A_79_21#_c_82_p N_A1_c_189_n 6.8073e-19 $X=2.665 $Y=0.785 $X2=-0.19
+ $Y2=-0.24
cc_70 N_A_79_21#_c_63_n N_A1_c_190_n 0.0166676f $X=3.555 $Y=1.575 $X2=0 $Y2=0
cc_71 N_A_79_21#_c_82_p N_A1_c_190_n 0.00510895f $X=2.665 $Y=0.785 $X2=0 $Y2=0
cc_72 N_A_79_21#_c_70_p A1 0.0111524f $X=2.475 $Y=0.785 $X2=0 $Y2=0
cc_73 N_A_79_21#_c_63_n A1 0.0217713f $X=3.555 $Y=1.575 $X2=0 $Y2=0
cc_74 N_A_79_21#_c_82_p A1 0.0149589f $X=2.665 $Y=0.785 $X2=0 $Y2=0
cc_75 N_A_79_21#_c_57_n N_B1_c_219_n 0.0136346f $X=3.555 $Y=0.785 $X2=-0.19
+ $Y2=-0.24
cc_76 N_A_79_21#_c_58_n N_B1_c_219_n 8.44804e-19 $X=3.77 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_77 N_A_79_21#_c_63_n N_B1_c_220_n 0.0209121f $X=3.555 $Y=1.575 $X2=0 $Y2=0
cc_78 N_A_79_21#_c_57_n N_B1_c_220_n 0.00501343f $X=3.555 $Y=0.785 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_65_n N_B1_c_220_n 0.00239548f $X=3.77 $Y=1.755 $X2=0 $Y2=0
cc_80 N_A_79_21#_c_63_n B1 0.0177736f $X=3.555 $Y=1.575 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_57_n B1 0.0203681f $X=3.555 $Y=0.785 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_57_n N_C1_c_246_n 0.0101229f $X=3.555 $Y=0.785 $X2=-0.19
+ $Y2=-0.24
cc_83 N_A_79_21#_c_58_n N_C1_c_246_n 0.00639463f $X=3.77 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_84 N_A_79_21#_c_63_n N_C1_c_247_n 0.0150745f $X=3.555 $Y=1.575 $X2=0 $Y2=0
cc_85 N_A_79_21#_c_57_n N_C1_c_247_n 0.00294707f $X=3.555 $Y=0.785 $X2=0 $Y2=0
cc_86 N_A_79_21#_c_65_n N_C1_c_247_n 0.0156516f $X=3.77 $Y=1.755 $X2=0 $Y2=0
cc_87 N_A_79_21#_c_63_n C1 0.0195108f $X=3.555 $Y=1.575 $X2=0 $Y2=0
cc_88 N_A_79_21#_c_57_n C1 0.023399f $X=3.555 $Y=0.785 $X2=0 $Y2=0
cc_89 N_A_79_21#_c_64_n N_VPWR_M1006_d 0.0041845f $X=1.355 $Y=1.575 $X2=0 $Y2=0
cc_90 N_A_79_21#_c_63_n N_VPWR_M1007_d 0.00758524f $X=3.555 $Y=1.575 $X2=0 $Y2=0
cc_91 N_A_79_21#_c_60_n N_VPWR_c_270_n 0.00484201f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A_79_21#_c_60_n N_VPWR_c_271_n 0.00702461f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_93 N_A_79_21#_c_61_n N_VPWR_c_271_n 0.00702461f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_79_21#_c_61_n N_VPWR_c_272_n 0.00459037f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A_79_21#_c_64_n N_VPWR_c_272_n 0.0219217f $X=1.355 $Y=1.575 $X2=0 $Y2=0
cc_96 N_A_79_21#_c_59_n N_VPWR_c_272_n 8.35232e-19 $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_97 N_A_79_21#_c_65_n N_VPWR_c_276_n 0.0128245f $X=3.77 $Y=1.755 $X2=0 $Y2=0
cc_98 N_A_79_21#_M1009_d N_VPWR_c_268_n 0.00237229f $X=3.625 $Y=1.485 $X2=0
+ $Y2=0
cc_99 N_A_79_21#_c_60_n N_VPWR_c_268_n 0.0133985f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A_79_21#_c_61_n N_VPWR_c_268_n 0.0138321f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_79_21#_c_65_n N_VPWR_c_268_n 0.0131136f $X=3.77 $Y=1.755 $X2=0 $Y2=0
cc_102 N_A_79_21#_c_54_n N_X_c_321_n 0.00495976f $X=0.47 $Y=1 $X2=0 $Y2=0
cc_103 N_A_79_21#_c_60_n N_X_c_321_n 0.00258957f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_79_21#_c_55_n N_X_c_321_n 0.00110025f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A_79_21#_c_61_n N_X_c_321_n 0.00126789f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_106 N_A_79_21#_c_56_n N_X_c_321_n 0.0324727f $X=1.185 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_79_21#_c_59_n N_X_c_321_n 0.0382763f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_63_n N_A_319_297#_M1007_s 0.00661259f $X=3.555 $Y=1.575
+ $X2=-0.19 $Y2=-0.24
cc_109 N_A_79_21#_c_63_n N_A_319_297#_M1004_d 0.00631695f $X=3.555 $Y=1.575
+ $X2=0 $Y2=0
cc_110 N_A_79_21#_c_63_n N_A_319_297#_c_339_n 0.0420721f $X=3.555 $Y=1.575 $X2=0
+ $Y2=0
cc_111 N_A_79_21#_c_63_n N_A_319_297#_c_336_n 0.0249887f $X=3.555 $Y=1.575 $X2=0
+ $Y2=0
cc_112 N_A_79_21#_c_63_n N_A_319_297#_c_341_n 0.0197281f $X=3.555 $Y=1.575 $X2=0
+ $Y2=0
cc_113 N_A_79_21#_c_65_n N_A_319_297#_c_341_n 0.0153157f $X=3.77 $Y=1.755 $X2=0
+ $Y2=0
cc_114 N_A_79_21#_c_63_n A_643_297# 0.00646447f $X=3.555 $Y=1.575 $X2=-0.19
+ $Y2=-0.24
cc_115 N_A_79_21#_c_56_n N_VGND_M1011_d 2.47258e-19 $X=1.185 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_70_p N_VGND_M1011_d 0.0174861f $X=2.475 $Y=0.785 $X2=0 $Y2=0
cc_117 N_A_79_21#_c_130_p N_VGND_M1011_d 0.00676892f $X=1.355 $Y=0.785 $X2=0
+ $Y2=0
cc_118 N_A_79_21#_c_57_n N_VGND_M1002_d 0.00715799f $X=3.555 $Y=0.785 $X2=0
+ $Y2=0
cc_119 N_A_79_21#_c_54_n N_VGND_c_365_n 0.00392847f $X=0.47 $Y=1 $X2=0 $Y2=0
cc_120 N_A_79_21#_c_57_n N_VGND_c_366_n 0.0208106f $X=3.555 $Y=0.785 $X2=0 $Y2=0
cc_121 N_A_79_21#_c_70_p N_VGND_c_367_n 0.0093646f $X=2.475 $Y=0.785 $X2=0 $Y2=0
cc_122 N_A_79_21#_c_71_p N_VGND_c_367_n 0.0210734f $X=2.69 $Y=0.36 $X2=0 $Y2=0
cc_123 N_A_79_21#_c_57_n N_VGND_c_367_n 0.00307876f $X=3.555 $Y=0.785 $X2=0
+ $Y2=0
cc_124 N_A_79_21#_c_57_n N_VGND_c_369_n 0.00212534f $X=3.555 $Y=0.785 $X2=0
+ $Y2=0
cc_125 N_A_79_21#_c_58_n N_VGND_c_369_n 0.0215942f $X=3.77 $Y=0.4 $X2=0 $Y2=0
cc_126 N_A_79_21#_M1010_d N_VGND_c_370_n 0.00334776f $X=2.5 $Y=0.235 $X2=0 $Y2=0
cc_127 N_A_79_21#_M1005_d N_VGND_c_370_n 0.0025127f $X=3.585 $Y=0.235 $X2=0
+ $Y2=0
cc_128 N_A_79_21#_c_54_n N_VGND_c_370_n 0.0115419f $X=0.47 $Y=1 $X2=0 $Y2=0
cc_129 N_A_79_21#_c_55_n N_VGND_c_370_n 0.00860847f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_79_21#_c_70_p N_VGND_c_370_n 0.0197196f $X=2.475 $Y=0.785 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_130_p N_VGND_c_370_n 0.00141553f $X=1.355 $Y=0.785 $X2=0
+ $Y2=0
cc_132 N_A_79_21#_c_71_p N_VGND_c_370_n 0.0141847f $X=2.69 $Y=0.36 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_57_n N_VGND_c_370_n 0.0112552f $X=3.555 $Y=0.785 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_58_n N_VGND_c_370_n 0.0141615f $X=3.77 $Y=0.4 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_54_n N_VGND_c_371_n 0.00585385f $X=0.47 $Y=1 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_55_n N_VGND_c_371_n 0.00505556f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_54_n N_VGND_c_372_n 5.1033e-19 $X=0.47 $Y=1 $X2=0 $Y2=0
cc_138 N_A_79_21#_c_55_n N_VGND_c_372_n 0.00848656f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_79_21#_c_70_p N_VGND_c_372_n 0.0227658f $X=2.475 $Y=0.785 $X2=0 $Y2=0
cc_140 N_A_79_21#_c_130_p N_VGND_c_372_n 0.0153171f $X=1.355 $Y=0.785 $X2=0
+ $Y2=0
cc_141 N_A_79_21#_c_59_n N_VGND_c_372_n 0.00229848f $X=0.965 $Y=1.202 $X2=0
+ $Y2=0
cc_142 N_A_79_21#_c_70_p A_421_47# 0.00487708f $X=2.475 $Y=0.785 $X2=-0.19
+ $Y2=-0.24
cc_143 N_A2_c_156_n N_A1_c_189_n 0.0332498f $X=2.03 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_144 N_A2_c_159_n N_A1_c_190_n 0.031436f $X=2.005 $Y=1.41 $X2=0 $Y2=0
cc_145 A2 N_A1_c_190_n 2.15878e-19 $X=1.62 $Y=1.105 $X2=0 $Y2=0
cc_146 N_A2_c_158_n N_A1_c_190_n 0.0366711f $X=2.005 $Y=1.202 $X2=0 $Y2=0
cc_147 A2 A1 0.0114795f $X=1.62 $Y=1.105 $X2=0 $Y2=0
cc_148 N_A2_c_158_n A1 0.00193773f $X=2.005 $Y=1.202 $X2=0 $Y2=0
cc_149 N_A2_c_159_n N_VPWR_c_272_n 0.00206436f $X=2.005 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A2_c_159_n N_VPWR_c_273_n 0.0061488f $X=2.005 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A2_c_159_n N_VPWR_c_274_n 0.00512582f $X=2.005 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A2_c_159_n N_VPWR_c_268_n 0.00833776f $X=2.005 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A2_c_159_n N_A_319_297#_c_339_n 0.0115703f $X=2.005 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A2_c_159_n N_A_319_297#_c_336_n 0.00749768f $X=2.005 $Y=1.41 $X2=0
+ $Y2=0
cc_155 N_A2_c_156_n N_VGND_c_367_n 0.00433717f $X=2.03 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A2_c_156_n N_VGND_c_370_n 0.0073635f $X=2.03 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A2_c_156_n N_VGND_c_372_n 0.0121728f $X=2.03 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A1_c_189_n N_B1_c_219_n 0.0163232f $X=2.425 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_159 N_A1_c_190_n N_B1_c_220_n 0.0555124f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_160 A1 N_B1_c_220_n 7.20932e-19 $X=2.435 $Y=1.105 $X2=0 $Y2=0
cc_161 N_A1_c_190_n B1 7.29446e-19 $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_162 A1 B1 0.0194549f $X=2.435 $Y=1.105 $X2=0 $Y2=0
cc_163 N_A1_c_190_n N_VPWR_c_273_n 0.00464319f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A1_c_190_n N_VPWR_c_276_n 0.00521297f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A1_c_190_n N_VPWR_c_268_n 0.00735433f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A1_c_190_n N_A_319_297#_c_339_n 0.0152751f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A1_c_190_n N_A_319_297#_c_336_n 7.48103e-19 $X=2.585 $Y=1.41 $X2=0
+ $Y2=0
cc_168 N_A1_c_189_n N_VGND_c_367_n 0.00423225f $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A1_c_189_n N_VGND_c_370_n 0.00611638f $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_170 N_B1_c_219_n N_C1_c_246_n 0.021585f $X=2.97 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_171 N_B1_c_220_n N_C1_c_247_n 0.0955909f $X=3.125 $Y=1.41 $X2=0 $Y2=0
cc_172 B1 N_C1_c_247_n 2.35867e-19 $X=2.975 $Y=1.105 $X2=0 $Y2=0
cc_173 N_B1_c_220_n C1 0.00137737f $X=3.125 $Y=1.41 $X2=0 $Y2=0
cc_174 B1 C1 0.0183874f $X=2.975 $Y=1.105 $X2=0 $Y2=0
cc_175 N_B1_c_220_n N_VPWR_c_276_n 0.00688798f $X=3.125 $Y=1.41 $X2=0 $Y2=0
cc_176 N_B1_c_220_n N_VPWR_c_268_n 0.0124404f $X=3.125 $Y=1.41 $X2=0 $Y2=0
cc_177 N_B1_c_220_n N_A_319_297#_c_341_n 0.01061f $X=3.125 $Y=1.41 $X2=0 $Y2=0
cc_178 N_B1_c_219_n N_VGND_c_366_n 0.00640381f $X=2.97 $Y=0.995 $X2=0 $Y2=0
cc_179 N_B1_c_219_n N_VGND_c_367_n 0.00433717f $X=2.97 $Y=0.995 $X2=0 $Y2=0
cc_180 N_B1_c_219_n N_VGND_c_370_n 0.00655915f $X=2.97 $Y=0.995 $X2=0 $Y2=0
cc_181 N_C1_c_247_n N_VPWR_c_276_n 0.00610391f $X=3.535 $Y=1.41 $X2=0 $Y2=0
cc_182 N_C1_c_247_n N_VPWR_c_268_n 0.0111713f $X=3.535 $Y=1.41 $X2=0 $Y2=0
cc_183 N_C1_c_247_n N_A_319_297#_c_341_n 0.00193883f $X=3.535 $Y=1.41 $X2=0
+ $Y2=0
cc_184 N_C1_c_246_n N_VGND_c_366_n 0.00299634f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_185 N_C1_c_246_n N_VGND_c_369_n 0.00420829f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_186 N_C1_c_246_n N_VGND_c_370_n 0.00702828f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_187 N_VPWR_c_268_n N_X_M1000_s 0.00462156f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_188 N_VPWR_c_271_n N_X_c_321_n 0.00774418f $X=1.1 $Y=2.72 $X2=0 $Y2=0
cc_189 N_VPWR_c_268_n N_X_c_321_n 0.00816554f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_190 N_VPWR_c_268_n N_A_319_297#_M1007_s 0.00258507f $X=3.91 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_191 N_VPWR_c_268_n N_A_319_297#_M1004_d 0.00305869f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_192 N_VPWR_M1007_d N_A_319_297#_c_339_n 0.00639376f $X=2.095 $Y=1.485 $X2=0
+ $Y2=0
cc_193 N_VPWR_c_273_n N_A_319_297#_c_339_n 0.0213073f $X=2.305 $Y=2.355 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_274_n N_A_319_297#_c_339_n 0.00277259f $X=2.155 $Y=2.72 $X2=0
+ $Y2=0
cc_195 N_VPWR_c_276_n N_A_319_297#_c_339_n 0.00346937f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_196 N_VPWR_c_268_n N_A_319_297#_c_339_n 0.0130554f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_197 N_VPWR_c_272_n N_A_319_297#_c_336_n 0.0466847f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_198 N_VPWR_c_273_n N_A_319_297#_c_336_n 0.0174485f $X=2.305 $Y=2.355 $X2=0
+ $Y2=0
cc_199 N_VPWR_c_274_n N_A_319_297#_c_336_n 0.0244364f $X=2.155 $Y=2.72 $X2=0
+ $Y2=0
cc_200 N_VPWR_c_268_n N_A_319_297#_c_336_n 0.0143661f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_201 N_VPWR_c_276_n N_A_319_297#_c_341_n 0.0203601f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_202 N_VPWR_c_268_n N_A_319_297#_c_341_n 0.0124905f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_203 N_VPWR_c_268_n A_643_297# 0.00983149f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_204 N_VPWR_c_270_n N_VGND_c_365_n 0.0104469f $X=0.26 $Y=1.655 $X2=0 $Y2=0
cc_205 N_X_c_321_n N_VGND_c_365_n 0.0210877f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_206 N_X_M1008_s N_VGND_c_370_n 0.00610537f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_207 N_X_c_321_n N_VGND_c_370_n 0.00878068f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_208 N_X_c_321_n N_VGND_c_371_n 0.0154757f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_209 N_VGND_c_370_n A_421_47# 0.00307614f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
