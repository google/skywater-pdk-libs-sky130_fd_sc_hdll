* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__probe_p_8 A VGND VNB VPB VPWR X
X0 a_399_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VGND a_27_47# a_399_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_399_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 VPWR a_27_47# a_399_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_399_297# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR a_27_47# a_399_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_399_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 a_399_297# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND a_27_47# a_399_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_399_297# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_399_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_399_297# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_399_297# X VPB short w=3.02e+06u l=5000u
X18 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 VPWR a_27_47# a_399_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 VGND a_27_47# a_399_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VPWR a_27_47# a_399_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 VGND a_27_47# a_399_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
