* File: sky130_fd_sc_hdll__dfrtp_4.pxi.spice
* Created: Wed Sep  2 08:28:14 2020
* 
x_PM_SKY130_FD_SC_HDLL__DFRTP_4%CLK N_CLK_c_218_n N_CLK_c_222_n N_CLK_c_223_n
+ N_CLK_M1004_g N_CLK_c_219_n N_CLK_M1021_g CLK CLK
+ PM_SKY130_FD_SC_HDLL__DFRTP_4%CLK
x_PM_SKY130_FD_SC_HDLL__DFRTP_4%A_27_47# N_A_27_47#_M1021_s N_A_27_47#_M1004_s
+ N_A_27_47#_c_275_n N_A_27_47#_c_276_n N_A_27_47#_M1027_g N_A_27_47#_M1002_g
+ N_A_27_47#_c_256_n N_A_27_47#_M1007_g N_A_27_47#_c_258_n N_A_27_47#_c_259_n
+ N_A_27_47#_c_279_n N_A_27_47#_c_280_n N_A_27_47#_M1000_g N_A_27_47#_c_260_n
+ N_A_27_47#_c_282_n N_A_27_47#_c_283_n N_A_27_47#_M1028_g N_A_27_47#_M1020_g
+ N_A_27_47#_c_262_n N_A_27_47#_c_263_n N_A_27_47#_c_264_n N_A_27_47#_c_284_n
+ N_A_27_47#_c_285_n N_A_27_47#_c_265_n N_A_27_47#_c_266_n N_A_27_47#_c_267_n
+ N_A_27_47#_c_268_n N_A_27_47#_c_269_n N_A_27_47#_c_270_n N_A_27_47#_c_271_n
+ N_A_27_47#_c_272_n N_A_27_47#_c_273_n N_A_27_47#_c_274_n
+ PM_SKY130_FD_SC_HDLL__DFRTP_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__DFRTP_4%D N_D_M1012_g N_D_c_503_n N_D_c_504_n
+ N_D_M1024_g N_D_c_501_n N_D_c_506_n D N_D_c_502_n
+ PM_SKY130_FD_SC_HDLL__DFRTP_4%D
x_PM_SKY130_FD_SC_HDLL__DFRTP_4%A_211_363# N_A_211_363#_M1002_d
+ N_A_211_363#_M1027_d N_A_211_363#_c_564_n N_A_211_363#_M1025_g
+ N_A_211_363#_M1014_g N_A_211_363#_c_557_n N_A_211_363#_M1005_g
+ N_A_211_363#_c_565_n N_A_211_363#_M1009_g N_A_211_363#_c_558_n
+ N_A_211_363#_c_559_n N_A_211_363#_c_560_n N_A_211_363#_c_568_n
+ N_A_211_363#_c_569_n N_A_211_363#_c_561_n N_A_211_363#_c_570_n
+ N_A_211_363#_c_571_n N_A_211_363#_c_572_n N_A_211_363#_c_573_n
+ N_A_211_363#_c_574_n N_A_211_363#_c_575_n N_A_211_363#_c_562_n
+ N_A_211_363#_c_576_n N_A_211_363#_c_563_n
+ PM_SKY130_FD_SC_HDLL__DFRTP_4%A_211_363#
x_PM_SKY130_FD_SC_HDLL__DFRTP_4%A_811_289# N_A_811_289#_M1032_d
+ N_A_811_289#_M1022_d N_A_811_289#_c_768_n N_A_811_289#_M1015_g
+ N_A_811_289#_M1001_g N_A_811_289#_c_770_n N_A_811_289#_c_791_n
+ N_A_811_289#_c_767_n N_A_811_289#_c_793_n N_A_811_289#_c_780_n
+ N_A_811_289#_c_798_n N_A_811_289#_c_783_n N_A_811_289#_c_810_p
+ N_A_811_289#_c_784_n N_A_811_289#_c_772_n
+ PM_SKY130_FD_SC_HDLL__DFRTP_4%A_811_289#
x_PM_SKY130_FD_SC_HDLL__DFRTP_4%RESET_B N_RESET_B_M1003_g N_RESET_B_c_872_n
+ N_RESET_B_c_886_n N_RESET_B_M1033_g N_RESET_B_c_873_n N_RESET_B_c_888_n
+ N_RESET_B_M1017_g N_RESET_B_M1029_g N_RESET_B_c_875_n N_RESET_B_c_876_n
+ N_RESET_B_c_877_n RESET_B N_RESET_B_c_878_n N_RESET_B_c_879_n
+ N_RESET_B_c_880_n N_RESET_B_c_881_n N_RESET_B_c_882_n N_RESET_B_c_883_n
+ RESET_B PM_SKY130_FD_SC_HDLL__DFRTP_4%RESET_B
x_PM_SKY130_FD_SC_HDLL__DFRTP_4%A_583_47# N_A_583_47#_M1007_d
+ N_A_583_47#_M1025_d N_A_583_47#_M1032_g N_A_583_47#_c_1032_n
+ N_A_583_47#_c_1033_n N_A_583_47#_M1022_g N_A_583_47#_c_1043_n
+ N_A_583_47#_c_1066_n N_A_583_47#_c_1034_n N_A_583_47#_c_1027_n
+ N_A_583_47#_c_1028_n N_A_583_47#_c_1029_n N_A_583_47#_c_1030_n
+ N_A_583_47#_c_1031_n PM_SKY130_FD_SC_HDLL__DFRTP_4%A_583_47#
x_PM_SKY130_FD_SC_HDLL__DFRTP_4%A_1403_21# N_A_1403_21#_M1013_d
+ N_A_1403_21#_M1017_d N_A_1403_21#_M1018_g N_A_1403_21#_c_1155_n
+ N_A_1403_21#_c_1171_n N_A_1403_21#_M1006_g N_A_1403_21#_c_1172_n
+ N_A_1403_21#_M1010_g N_A_1403_21#_c_1156_n N_A_1403_21#_M1008_g
+ N_A_1403_21#_c_1173_n N_A_1403_21#_M1016_g N_A_1403_21#_c_1157_n
+ N_A_1403_21#_M1023_g N_A_1403_21#_c_1174_n N_A_1403_21#_M1019_g
+ N_A_1403_21#_c_1158_n N_A_1403_21#_M1030_g N_A_1403_21#_c_1175_n
+ N_A_1403_21#_M1026_g N_A_1403_21#_c_1159_n N_A_1403_21#_M1031_g
+ N_A_1403_21#_c_1160_n N_A_1403_21#_c_1161_n N_A_1403_21#_c_1201_n
+ N_A_1403_21#_c_1206_n N_A_1403_21#_c_1255_p N_A_1403_21#_c_1176_n
+ N_A_1403_21#_c_1177_n N_A_1403_21#_c_1162_n N_A_1403_21#_c_1163_n
+ N_A_1403_21#_c_1164_n N_A_1403_21#_c_1165_n N_A_1403_21#_c_1166_n
+ N_A_1403_21#_c_1167_n N_A_1403_21#_c_1168_n N_A_1403_21#_c_1169_n
+ PM_SKY130_FD_SC_HDLL__DFRTP_4%A_1403_21#
x_PM_SKY130_FD_SC_HDLL__DFRTP_4%A_1188_47# N_A_1188_47#_M1005_d
+ N_A_1188_47#_M1028_d N_A_1188_47#_c_1355_n N_A_1188_47#_M1011_g
+ N_A_1188_47#_M1013_g N_A_1188_47#_c_1360_n N_A_1188_47#_c_1363_n
+ N_A_1188_47#_c_1354_n N_A_1188_47#_c_1357_n N_A_1188_47#_c_1358_n
+ N_A_1188_47#_c_1359_n PM_SKY130_FD_SC_HDLL__DFRTP_4%A_1188_47#
x_PM_SKY130_FD_SC_HDLL__DFRTP_4%VPWR N_VPWR_M1004_d N_VPWR_M1024_s
+ N_VPWR_M1015_d N_VPWR_M1022_s N_VPWR_M1006_d N_VPWR_M1011_d N_VPWR_M1010_d
+ N_VPWR_M1016_d N_VPWR_M1026_d N_VPWR_c_1454_n N_VPWR_c_1455_n N_VPWR_c_1456_n
+ N_VPWR_c_1457_n N_VPWR_c_1458_n N_VPWR_c_1459_n N_VPWR_c_1460_n
+ N_VPWR_c_1461_n N_VPWR_c_1462_n N_VPWR_c_1463_n N_VPWR_c_1464_n
+ N_VPWR_c_1465_n N_VPWR_c_1466_n N_VPWR_c_1467_n N_VPWR_c_1468_n
+ N_VPWR_c_1469_n N_VPWR_c_1470_n N_VPWR_c_1471_n N_VPWR_c_1472_n VPWR
+ N_VPWR_c_1473_n N_VPWR_c_1474_n N_VPWR_c_1475_n N_VPWR_c_1476_n
+ N_VPWR_c_1453_n N_VPWR_c_1478_n N_VPWR_c_1479_n N_VPWR_c_1480_n
+ N_VPWR_c_1481_n PM_SKY130_FD_SC_HDLL__DFRTP_4%VPWR
x_PM_SKY130_FD_SC_HDLL__DFRTP_4%A_468_47# N_A_468_47#_M1012_d
+ N_A_468_47#_M1024_d N_A_468_47#_c_1624_n N_A_468_47#_c_1643_n
+ N_A_468_47#_c_1632_n PM_SKY130_FD_SC_HDLL__DFRTP_4%A_468_47#
x_PM_SKY130_FD_SC_HDLL__DFRTP_4%A_699_413# N_A_699_413#_M1000_d
+ N_A_699_413#_M1033_d N_A_699_413#_c_1659_n N_A_699_413#_c_1660_n
+ N_A_699_413#_c_1661_n N_A_699_413#_c_1662_n
+ PM_SKY130_FD_SC_HDLL__DFRTP_4%A_699_413#
x_PM_SKY130_FD_SC_HDLL__DFRTP_4%Q N_Q_M1008_s N_Q_M1030_s N_Q_M1010_s
+ N_Q_M1019_s N_Q_c_1710_n N_Q_c_1704_n N_Q_c_1716_n N_Q_c_1698_n N_Q_c_1699_n
+ N_Q_c_1705_n N_Q_c_1730_n N_Q_c_1751_n N_Q_c_1706_n N_Q_c_1700_n N_Q_c_1701_n
+ N_Q_c_1707_n Q Q Q N_Q_c_1703_n N_Q_c_1709_n PM_SKY130_FD_SC_HDLL__DFRTP_4%Q
x_PM_SKY130_FD_SC_HDLL__DFRTP_4%VGND N_VGND_M1021_d N_VGND_M1012_s
+ N_VGND_M1003_d N_VGND_M1018_d N_VGND_M1008_d N_VGND_M1023_d N_VGND_M1031_d
+ N_VGND_c_1775_n N_VGND_c_1776_n N_VGND_c_1777_n N_VGND_c_1778_n
+ N_VGND_c_1779_n N_VGND_c_1780_n N_VGND_c_1781_n N_VGND_c_1782_n
+ N_VGND_c_1783_n N_VGND_c_1784_n N_VGND_c_1785_n N_VGND_c_1786_n
+ N_VGND_c_1787_n N_VGND_c_1788_n VGND N_VGND_c_1789_n N_VGND_c_1790_n
+ N_VGND_c_1791_n N_VGND_c_1792_n N_VGND_c_1793_n N_VGND_c_1794_n
+ N_VGND_c_1795_n N_VGND_c_1796_n PM_SKY130_FD_SC_HDLL__DFRTP_4%VGND
cc_1 VNB N_CLK_c_218_n 0.0612188f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.325
cc_2 VNB N_CLK_c_219_n 0.0173562f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_3 VNB CLK 0.0160726f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_A_27_47#_M1002_g 0.0398926f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_5 VNB N_A_27_47#_c_256_n 0.00994239f $X=-0.19 $Y=-0.24 $X2=0.352 $Y2=1.16
cc_6 VNB N_A_27_47#_M1007_g 0.0224944f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.16
cc_7 VNB N_A_27_47#_c_258_n 0.015931f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_259_n 0.00231033f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_9 VNB N_A_27_47#_c_260_n 0.0446574f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_M1020_g 0.0308613f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_262_n 0.0111414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_263_n 0.00233121f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_264_n 0.00783792f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_265_n 0.0267455f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_266_n 0.00242452f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_267_n 0.0332386f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_268_n 7.01061e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_269_n 0.00705679f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_270_n 0.00200162f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_271_n 0.0267704f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_272_n 0.0276305f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_273_n 0.00935418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_274_n 0.00683758f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_D_M1012_g 0.0551753f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.74
cc_25 VNB N_D_c_501_n 0.0139927f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_D_c_502_n 0.0204858f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.16
cc_27 VNB N_A_211_363#_M1014_g 0.0242964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_211_363#_c_557_n 0.0189002f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_29 VNB N_A_211_363#_c_558_n 0.00308451f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_211_363#_c_559_n 0.00571147f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_211_363#_c_560_n 0.0427899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_211_363#_c_561_n 0.0033367f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_211_363#_c_562_n 0.0315937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_211_363#_c_563_n 0.01291f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_811_289#_M1001_g 0.0484711f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_811_289#_c_767_n 0.00721918f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_RESET_B_c_872_n 0.0101914f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_38 VNB N_RESET_B_c_873_n 0.00103828f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_RESET_B_M1029_g 0.0304839f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_RESET_B_c_875_n 0.00618905f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_41 VNB N_RESET_B_c_876_n 0.0212513f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_42 VNB N_RESET_B_c_877_n 0.00104886f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_RESET_B_c_878_n 0.0295986f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_RESET_B_c_879_n 0.00913762f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_RESET_B_c_880_n 0.0180246f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_RESET_B_c_881_n 0.0288472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_RESET_B_c_882_n 0.00638876f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_RESET_B_c_883_n 0.00441814f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB RESET_B 0.00633626f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_583_47#_M1032_g 0.0198147f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_51 VNB N_A_583_47#_c_1027_n 0.0122699f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_583_47#_c_1028_n 0.0073066f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_583_47#_c_1029_n 0.00322861f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_583_47#_c_1030_n 0.00185456f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_583_47#_c_1031_n 0.0317322f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_1403_21#_M1018_g 0.0237218f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_57 VNB N_A_1403_21#_c_1155_n 0.0111493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_1403_21#_c_1156_n 0.0201651f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_59 VNB N_A_1403_21#_c_1157_n 0.0167673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_1403_21#_c_1158_n 0.0167581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_1403_21#_c_1159_n 0.0196229f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_1403_21#_c_1160_n 0.00209314f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1403_21#_c_1161_n 7.82159e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_1403_21#_c_1162_n 0.00284289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_1403_21#_c_1163_n 0.00628208f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1403_21#_c_1164_n 0.0147678f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1403_21#_c_1165_n 2.29591e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1403_21#_c_1166_n 0.016811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_1403_21#_c_1167_n 0.0081134f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_1403_21#_c_1168_n 0.0546825f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_1403_21#_c_1169_n 0.0868798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_1188_47#_M1013_g 0.0506579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1188_47#_c_1354_n 0.00743571f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_74 VNB N_VPWR_c_1453_n 0.478484f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_468_47#_c_1624_n 0.0051081f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_76 VNB N_Q_c_1698_n 0.00264486f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_Q_c_1699_n 0.00232612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_Q_c_1700_n 6.43096e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_Q_c_1701_n 0.00232612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB Q 0.0233631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_Q_c_1703_n 0.0103908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1775_n 0.00858778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1776_n 0.00564356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1777_n 0.00513781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1778_n 0.00646908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1779_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1780_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1781_n 0.0216385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1782_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1783_n 0.0381083f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1784_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1785_n 0.0199309f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1786_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1787_n 0.0193029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1788_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1789_n 0.014742f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1790_n 0.0782767f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1791_n 0.0552412f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1792_n 0.0113686f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1793_n 0.541443f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1794_n 0.0085923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1795_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1796_n 0.00458779f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VPB N_CLK_c_218_n 0.00482568f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.325
cc_105 VPB N_CLK_c_222_n 0.014844f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_106 VPB N_CLK_c_223_n 0.0466088f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.74
cc_107 VPB CLK 0.0154183f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_108 VPB N_A_27_47#_c_275_n 0.0192832f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_109 VPB N_A_27_47#_c_276_n 0.025741f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_110 VPB N_A_27_47#_c_258_n 0.0167703f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_27_47#_c_259_n 0.00701107f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.53
cc_112 VPB N_A_27_47#_c_279_n 0.0299621f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_27_47#_c_280_n 0.025222f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_27_47#_c_260_n 0.0132357f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_27_47#_c_282_n 0.0299456f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_27_47#_c_283_n 0.0240442f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_27_47#_c_284_n 0.00133165f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_27_47#_c_285_n 0.0297432f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_27_47#_c_266_n 4.26143e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_27_47#_c_269_n 0.00369171f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_27_47#_c_270_n 3.60888e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_27_47#_c_271_n 0.0125132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_27_47#_c_273_n 0.0028911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_27_47#_c_274_n 9.86971e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_D_c_503_n 0.0168054f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_126 VPB N_D_c_504_n 0.0266858f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_127 VPB N_D_c_501_n 0.0355324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_D_c_506_n 0.024376f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.665
cc_129 VPB D 0.0222332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_D_c_502_n 0.00669841f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.16
cc_131 VPB N_A_211_363#_c_564_n 0.0529433f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_132 VPB N_A_211_363#_c_565_n 0.0590351f $X=-0.19 $Y=1.305 $X2=0.352 $Y2=1.16
cc_133 VPB N_A_211_363#_c_558_n 0.00584199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_211_363#_c_559_n 0.00400344f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_211_363#_c_568_n 0.00222651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_211_363#_c_569_n 0.00167605f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_211_363#_c_570_n 0.0127037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_211_363#_c_571_n 0.00230751f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_211_363#_c_572_n 0.0161202f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_211_363#_c_573_n 0.00180228f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_211_363#_c_574_n 0.006632f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_211_363#_c_575_n 0.00254605f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_211_363#_c_576_n 0.00886602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_211_363#_c_563_n 0.0114316f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_811_289#_c_768_n 0.0629228f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_146 VPB N_A_811_289#_M1001_g 0.00836073f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_811_289#_c_770_n 0.0139674f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_148 VPB N_A_811_289#_c_767_n 0.00184276f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_811_289#_c_772_n 4.8645e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_RESET_B_c_872_n 0.0385919f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_151 VPB N_RESET_B_c_886_n 0.0266961f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_152 VPB N_RESET_B_c_873_n 0.033485f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_RESET_B_c_888_n 0.0241411f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.665
cc_154 VPB N_RESET_B_c_883_n 0.00505769f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_583_47#_c_1032_n 0.0301195f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.665
cc_156 VPB N_A_583_47#_c_1033_n 0.0188477f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_157 VPB N_A_583_47#_c_1034_n 0.0077712f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_583_47#_c_1028_n 0.00816282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_583_47#_c_1029_n 0.00346469f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_583_47#_c_1030_n 0.00113493f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_583_47#_c_1031_n 0.0256197f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_1403_21#_c_1155_n 0.0350675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_1403_21#_c_1171_n 0.0233838f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_164 VPB N_A_1403_21#_c_1172_n 0.0195138f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_1403_21#_c_1173_n 0.0159705f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_1403_21#_c_1174_n 0.0159551f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_1403_21#_c_1175_n 0.0191365f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_1403_21#_c_1176_n 0.00793653f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_1403_21#_c_1177_n 0.0031203f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_1403_21#_c_1165_n 0.0144264f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_1403_21#_c_1169_n 0.0503129f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_1188_47#_c_1355_n 0.0619838f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_173 VPB N_A_1188_47#_M1013_g 0.0114533f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_1188_47#_c_1357_n 0.00315851f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_1188_47#_c_1358_n 0.0134285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_1188_47#_c_1359_n 0.0244291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1454_n 0.00126291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1455_n 0.0093324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1456_n 0.00286019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1457_n 0.00785764f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1458_n 0.00234526f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1459_n 0.0138694f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1460_n 0.00362149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1461_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1462_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1463_n 0.0184687f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1464_n 0.0067475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_1465_n 0.0464278f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_1466_n 0.00359728f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1467_n 0.0088131f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1468_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1469_n 0.0216041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1470_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1471_n 0.0221062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1472_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1473_n 0.0146985f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1474_n 0.0281279f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1475_n 0.0529119f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1476_n 0.0121672f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1453_n 0.0714013f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1478_n 0.0054556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1479_n 0.00478085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1480_n 0.00513379f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1481_n 0.00987527f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_A_468_47#_c_1624_n 0.0079504f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_206 VPB N_A_699_413#_c_1659_n 4.96295e-19 $X=-0.19 $Y=1.305 $X2=0.305
+ $Y2=1.665
cc_207 VPB N_A_699_413#_c_1660_n 0.00909504f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.665
cc_208 VPB N_A_699_413#_c_1661_n 0.00247249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_A_699_413#_c_1662_n 7.36897e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_Q_c_1704_n 0.0019704f $X=-0.19 $Y=1.305 $X2=0.352 $Y2=1.16
cc_211 VPB N_Q_c_1705_n 0.0018222f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.53
cc_212 VPB N_Q_c_1706_n 5.77105e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_Q_c_1707_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB Q 0.00868578f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_Q_c_1709_n 0.0133798f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 N_CLK_c_222_n N_A_27_47#_c_275_n 0.00262901f $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_217 N_CLK_c_223_n N_A_27_47#_c_275_n 0.00668506f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_218 CLK N_A_27_47#_c_275_n 8.03089e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_219 N_CLK_c_223_n N_A_27_47#_c_276_n 0.0192779f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_220 N_CLK_c_218_n N_A_27_47#_M1002_g 0.00192687f $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_221 N_CLK_c_219_n N_A_27_47#_M1002_g 0.0154184f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_222 N_CLK_c_218_n N_A_27_47#_c_263_n 0.0108877f $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_223 N_CLK_c_219_n N_A_27_47#_c_263_n 0.00652815f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_224 CLK N_A_27_47#_c_263_n 0.00736322f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_225 N_CLK_c_218_n N_A_27_47#_c_264_n 0.0070116f $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_226 CLK N_A_27_47#_c_264_n 0.0220292f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_227 N_CLK_c_223_n N_A_27_47#_c_284_n 0.0171402f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_228 CLK N_A_27_47#_c_284_n 0.00731943f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_229 N_CLK_c_218_n N_A_27_47#_c_285_n 4.93713e-19 $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_230 N_CLK_c_223_n N_A_27_47#_c_285_n 0.00841026f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_231 CLK N_A_27_47#_c_285_n 0.0231715f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_232 CLK N_A_27_47#_c_266_n 0.00762548f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_233 N_CLK_c_218_n N_A_27_47#_c_269_n 0.0029245f $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_234 N_CLK_c_222_n N_A_27_47#_c_269_n 4.50807e-19 $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_235 N_CLK_c_223_n N_A_27_47#_c_269_n 0.00460739f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_236 CLK N_A_27_47#_c_269_n 0.0396442f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_237 N_CLK_c_218_n N_A_27_47#_c_271_n 0.0139997f $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_238 CLK N_A_27_47#_c_271_n 0.00161375f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_239 N_CLK_c_223_n N_VPWR_c_1454_n 0.0125197f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_240 N_CLK_c_223_n N_VPWR_c_1473_n 0.00304525f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_241 N_CLK_c_223_n N_VPWR_c_1453_n 0.00454898f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_242 N_CLK_c_218_n N_VGND_c_1789_n 6.41851e-19 $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_243 N_CLK_c_219_n N_VGND_c_1789_n 0.00198377f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_244 N_CLK_c_219_n N_VGND_c_1793_n 0.00367064f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_245 N_CLK_c_219_n N_VGND_c_1794_n 0.0142867f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_246 N_A_27_47#_c_256_n N_D_M1012_g 0.00468817f $X=2.817 $Y=1.245 $X2=0 $Y2=0
cc_247 N_A_27_47#_M1007_g N_D_M1012_g 0.0133483f $X=2.84 $Y=0.415 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_265_n N_D_M1012_g 0.00249406f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_249 N_A_27_47#_c_268_n N_D_M1012_g 0.00139106f $X=2.825 $Y=1.19 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_272_n N_D_M1012_g 0.0148947f $X=2.735 $Y=0.93 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_273_n N_D_M1012_g 0.00395248f $X=2.735 $Y=0.93 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_265_n N_D_c_501_n 0.00328759f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_253 N_A_27_47#_c_271_n N_D_c_501_n 0.00312973f $X=0.99 $Y=1.235 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_259_n N_D_c_506_n 0.00468817f $X=2.92 $Y=1.32 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_265_n N_D_c_506_n 0.00221183f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_256 N_A_27_47#_c_265_n N_D_c_502_n 0.0506264f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_257 N_A_27_47#_c_259_n N_A_211_363#_c_564_n 0.0220389f $X=2.92 $Y=1.32 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_c_279_n N_A_211_363#_c_564_n 0.0183435f $X=3.405 $Y=1.89 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_280_n N_A_211_363#_c_564_n 0.0157142f $X=3.405 $Y=1.99 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_272_n N_A_211_363#_c_564_n 6.13774e-19 $X=2.735 $Y=0.93
+ $X2=0 $Y2=0
cc_261 N_A_27_47#_c_273_n N_A_211_363#_c_564_n 0.00148383f $X=2.735 $Y=0.93
+ $X2=0 $Y2=0
cc_262 N_A_27_47#_M1007_g N_A_211_363#_M1014_g 0.0115275f $X=2.84 $Y=0.415 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_M1020_g N_A_211_363#_c_557_n 0.0138474f $X=6.51 $Y=0.415 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_260_n N_A_211_363#_c_565_n 0.00310475f $X=6.32 $Y=1.395
+ $X2=0 $Y2=0
cc_265 N_A_27_47#_c_282_n N_A_211_363#_c_565_n 0.0160483f $X=6.32 $Y=1.89 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_c_283_n N_A_211_363#_c_565_n 0.0141144f $X=6.32 $Y=1.99 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_270_n N_A_211_363#_c_565_n 0.0010284f $X=6.61 $Y=1.19 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_274_n N_A_211_363#_c_565_n 4.78088e-19 $X=6.57 $Y=1.11 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_258_n N_A_211_363#_c_558_n 0.0116146f $X=3.305 $Y=1.32 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_279_n N_A_211_363#_c_558_n 0.00442969f $X=3.405 $Y=1.89
+ $X2=0 $Y2=0
cc_271 N_A_27_47#_c_267_n N_A_211_363#_c_558_n 0.0113699f $X=6.465 $Y=1.19 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_268_n N_A_211_363#_c_558_n 4.95484e-19 $X=2.825 $Y=1.19
+ $X2=0 $Y2=0
cc_273 N_A_27_47#_c_272_n N_A_211_363#_c_558_n 0.00150125f $X=2.735 $Y=0.93
+ $X2=0 $Y2=0
cc_274 N_A_27_47#_c_273_n N_A_211_363#_c_558_n 0.0293808f $X=2.735 $Y=0.93 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_260_n N_A_211_363#_c_559_n 0.00878869f $X=6.32 $Y=1.395
+ $X2=0 $Y2=0
cc_276 N_A_27_47#_M1020_g N_A_211_363#_c_559_n 3.66012e-19 $X=6.51 $Y=0.415
+ $X2=0 $Y2=0
cc_277 N_A_27_47#_c_267_n N_A_211_363#_c_559_n 0.0148653f $X=6.465 $Y=1.19 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_270_n N_A_211_363#_c_559_n 4.59004e-19 $X=6.61 $Y=1.19 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_274_n N_A_211_363#_c_559_n 0.0462576f $X=6.57 $Y=1.11 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_M1020_g N_A_211_363#_c_560_n 0.0163952f $X=6.51 $Y=0.415 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_267_n N_A_211_363#_c_560_n 0.00222666f $X=6.465 $Y=1.19
+ $X2=0 $Y2=0
cc_282 N_A_27_47#_c_274_n N_A_211_363#_c_560_n 0.00214859f $X=6.57 $Y=1.11 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_260_n N_A_211_363#_c_568_n 0.00133124f $X=6.32 $Y=1.395
+ $X2=0 $Y2=0
cc_284 N_A_27_47#_c_282_n N_A_211_363#_c_568_n 0.0139123f $X=6.32 $Y=1.89 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_267_n N_A_211_363#_c_568_n 0.00508651f $X=6.465 $Y=1.19
+ $X2=0 $Y2=0
cc_286 N_A_27_47#_c_274_n N_A_211_363#_c_568_n 0.0117591f $X=6.57 $Y=1.11 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_258_n N_A_211_363#_c_561_n 0.00143371f $X=3.305 $Y=1.32
+ $X2=0 $Y2=0
cc_288 N_A_27_47#_c_267_n N_A_211_363#_c_561_n 0.0111717f $X=6.465 $Y=1.19 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_272_n N_A_211_363#_c_561_n 7.17844e-19 $X=2.735 $Y=0.93
+ $X2=0 $Y2=0
cc_290 N_A_27_47#_c_273_n N_A_211_363#_c_561_n 0.0187842f $X=2.735 $Y=0.93 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_265_n N_A_211_363#_c_570_n 0.0515231f $X=2.535 $Y=1.19 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_267_n N_A_211_363#_c_570_n 0.00873978f $X=6.465 $Y=1.19
+ $X2=0 $Y2=0
cc_293 N_A_27_47#_c_268_n N_A_211_363#_c_570_n 0.0133153f $X=2.825 $Y=1.19 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_273_n N_A_211_363#_c_570_n 0.00563605f $X=2.735 $Y=0.93
+ $X2=0 $Y2=0
cc_295 N_A_27_47#_c_276_n N_A_211_363#_c_571_n 0.00479165f $X=0.965 $Y=1.74
+ $X2=0 $Y2=0
cc_296 N_A_27_47#_c_284_n N_A_211_363#_c_571_n 0.00546643f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_265_n N_A_211_363#_c_571_n 0.0161767f $X=2.535 $Y=1.19 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_269_n N_A_211_363#_c_571_n 0.00111166f $X=0.745 $Y=1.19
+ $X2=0 $Y2=0
cc_299 N_A_27_47#_c_279_n N_A_211_363#_c_572_n 0.00272583f $X=3.405 $Y=1.89
+ $X2=0 $Y2=0
cc_300 N_A_27_47#_c_280_n N_A_211_363#_c_572_n 0.00153589f $X=3.405 $Y=1.99
+ $X2=0 $Y2=0
cc_301 N_A_27_47#_c_282_n N_A_211_363#_c_572_n 0.00359908f $X=6.32 $Y=1.89 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_283_n N_A_211_363#_c_572_n 0.00375592f $X=6.32 $Y=1.99 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_267_n N_A_211_363#_c_572_n 0.134385f $X=6.465 $Y=1.19 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_258_n N_A_211_363#_c_573_n 3.78985e-19 $X=3.305 $Y=1.32
+ $X2=0 $Y2=0
cc_305 N_A_27_47#_c_279_n N_A_211_363#_c_573_n 0.00162956f $X=3.405 $Y=1.89
+ $X2=0 $Y2=0
cc_306 N_A_27_47#_c_280_n N_A_211_363#_c_573_n 0.00114104f $X=3.405 $Y=1.99
+ $X2=0 $Y2=0
cc_307 N_A_27_47#_c_267_n N_A_211_363#_c_573_n 0.0129897f $X=6.465 $Y=1.19 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_258_n N_A_211_363#_c_574_n 8.09221e-19 $X=3.305 $Y=1.32
+ $X2=0 $Y2=0
cc_309 N_A_27_47#_c_259_n N_A_211_363#_c_574_n 0.00575298f $X=2.92 $Y=1.32 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_279_n N_A_211_363#_c_574_n 0.00371639f $X=3.405 $Y=1.89
+ $X2=0 $Y2=0
cc_311 N_A_27_47#_c_267_n N_A_211_363#_c_574_n 0.00544465f $X=6.465 $Y=1.19
+ $X2=0 $Y2=0
cc_312 N_A_27_47#_c_268_n N_A_211_363#_c_574_n 2.72172e-19 $X=2.825 $Y=1.19
+ $X2=0 $Y2=0
cc_313 N_A_27_47#_c_273_n N_A_211_363#_c_574_n 0.0115098f $X=2.735 $Y=0.93 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_282_n N_A_211_363#_c_575_n 7.85835e-19 $X=6.32 $Y=1.89 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_283_n N_A_211_363#_c_575_n 8.1316e-19 $X=6.32 $Y=1.99 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_270_n N_A_211_363#_c_575_n 0.0163395f $X=6.61 $Y=1.19 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_274_n N_A_211_363#_c_575_n 8.5067e-19 $X=6.57 $Y=1.11 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_258_n N_A_211_363#_c_562_n 0.0262961f $X=3.305 $Y=1.32 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_267_n N_A_211_363#_c_562_n 0.00330092f $X=6.465 $Y=1.19
+ $X2=0 $Y2=0
cc_320 N_A_27_47#_c_272_n N_A_211_363#_c_562_n 0.0175402f $X=2.735 $Y=0.93 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_273_n N_A_211_363#_c_562_n 8.5661e-19 $X=2.735 $Y=0.93 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_260_n N_A_211_363#_c_576_n 0.00487863f $X=6.32 $Y=1.395
+ $X2=0 $Y2=0
cc_323 N_A_27_47#_c_282_n N_A_211_363#_c_576_n 0.00572726f $X=6.32 $Y=1.89 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_270_n N_A_211_363#_c_576_n 0.00268408f $X=6.61 $Y=1.19 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_274_n N_A_211_363#_c_576_n 0.0184855f $X=6.57 $Y=1.11 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_276_n N_A_211_363#_c_563_n 0.0065704f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_M1002_g N_A_211_363#_c_563_n 0.0219823f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_263_n N_A_211_363#_c_563_n 0.0103201f $X=0.66 $Y=0.72 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_284_n N_A_211_363#_c_563_n 0.00841124f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_265_n N_A_211_363#_c_563_n 0.0193232f $X=2.535 $Y=1.19 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_266_n N_A_211_363#_c_563_n 0.00224499f $X=0.89 $Y=1.19 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_269_n N_A_211_363#_c_563_n 0.0568565f $X=0.745 $Y=1.19 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_c_279_n N_A_811_289#_c_768_n 0.00905857f $X=3.405 $Y=1.89
+ $X2=0 $Y2=0
cc_334 N_A_27_47#_c_280_n N_A_811_289#_c_768_n 0.00751882f $X=3.405 $Y=1.99
+ $X2=0 $Y2=0
cc_335 N_A_27_47#_c_258_n N_A_811_289#_M1001_g 0.00220848f $X=3.305 $Y=1.32
+ $X2=0 $Y2=0
cc_336 N_A_27_47#_c_267_n N_A_811_289#_M1001_g 0.0022411f $X=6.465 $Y=1.19 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_279_n N_A_811_289#_c_770_n 6.41051e-19 $X=3.405 $Y=1.89
+ $X2=0 $Y2=0
cc_338 N_A_27_47#_c_267_n N_A_811_289#_c_770_n 0.00937231f $X=6.465 $Y=1.19
+ $X2=0 $Y2=0
cc_339 N_A_27_47#_c_267_n N_A_811_289#_c_767_n 0.0135227f $X=6.465 $Y=1.19 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_c_282_n N_A_811_289#_c_780_n 0.00212864f $X=6.32 $Y=1.89 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_c_283_n N_A_811_289#_c_780_n 4.39557e-19 $X=6.32 $Y=1.99 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_267_n N_A_811_289#_c_780_n 0.00251211f $X=6.465 $Y=1.19
+ $X2=0 $Y2=0
cc_343 N_A_27_47#_c_283_n N_A_811_289#_c_783_n 0.00558596f $X=6.32 $Y=1.99 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_267_n N_A_811_289#_c_784_n 0.0015131f $X=6.465 $Y=1.19 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_267_n N_RESET_B_c_872_n 0.00187172f $X=6.465 $Y=1.19 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_267_n N_RESET_B_c_875_n 0.0676268f $X=6.465 $Y=1.19 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_260_n N_RESET_B_c_876_n 5.35574e-19 $X=6.32 $Y=1.395 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_267_n N_RESET_B_c_876_n 0.121696f $X=6.465 $Y=1.19 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_270_n N_RESET_B_c_876_n 0.0298783f $X=6.61 $Y=1.19 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_274_n N_RESET_B_c_876_n 0.0233523f $X=6.57 $Y=1.11 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_267_n N_RESET_B_c_878_n 0.00219045f $X=6.465 $Y=1.19 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_267_n N_RESET_B_c_879_n 0.004609f $X=6.465 $Y=1.19 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_282_n N_A_583_47#_c_1032_n 0.0046947f $X=6.32 $Y=1.89 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_c_267_n N_A_583_47#_c_1032_n 0.00392735f $X=6.465 $Y=1.19
+ $X2=0 $Y2=0
cc_355 N_A_27_47#_c_282_n N_A_583_47#_c_1033_n 0.0138263f $X=6.32 $Y=1.89 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_283_n N_A_583_47#_c_1033_n 0.0125159f $X=6.32 $Y=1.99 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_280_n N_A_583_47#_c_1043_n 0.0191355f $X=3.405 $Y=1.99 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_c_258_n N_A_583_47#_c_1034_n 0.00124445f $X=3.305 $Y=1.32
+ $X2=0 $Y2=0
cc_359 N_A_27_47#_c_279_n N_A_583_47#_c_1034_n 0.011704f $X=3.405 $Y=1.89 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_280_n N_A_583_47#_c_1034_n 0.00518242f $X=3.405 $Y=1.99
+ $X2=0 $Y2=0
cc_361 N_A_27_47#_c_267_n N_A_583_47#_c_1034_n 4.47512e-19 $X=6.465 $Y=1.19
+ $X2=0 $Y2=0
cc_362 N_A_27_47#_c_267_n N_A_583_47#_c_1027_n 0.0136728f $X=6.465 $Y=1.19 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_267_n N_A_583_47#_c_1028_n 0.0428999f $X=6.465 $Y=1.19 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_258_n N_A_583_47#_c_1029_n 0.00414f $X=3.305 $Y=1.32 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_267_n N_A_583_47#_c_1029_n 0.0135902f $X=6.465 $Y=1.19 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_267_n N_A_583_47#_c_1030_n 0.0103471f $X=6.465 $Y=1.19 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_267_n N_A_583_47#_c_1031_n 0.00555554f $X=6.465 $Y=1.19
+ $X2=0 $Y2=0
cc_368 N_A_27_47#_M1020_g N_A_1403_21#_M1018_g 0.0214866f $X=6.51 $Y=0.415 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_274_n N_A_1403_21#_M1018_g 7.83497e-19 $X=6.57 $Y=1.11 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_c_260_n N_A_1403_21#_c_1155_n 6.96482e-19 $X=6.32 $Y=1.395
+ $X2=0 $Y2=0
cc_371 N_A_27_47#_c_260_n N_A_1403_21#_c_1168_n 0.00673213f $X=6.32 $Y=1.395
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_c_260_n N_A_1188_47#_c_1360_n 0.00117242f $X=6.32 $Y=1.395
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_M1020_g N_A_1188_47#_c_1360_n 0.01612f $X=6.51 $Y=0.415 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_c_274_n N_A_1188_47#_c_1360_n 0.0290942f $X=6.57 $Y=1.11 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_c_283_n N_A_1188_47#_c_1363_n 0.00711535f $X=6.32 $Y=1.99
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_c_260_n N_A_1188_47#_c_1354_n 0.00263092f $X=6.32 $Y=1.395
+ $X2=0 $Y2=0
cc_377 N_A_27_47#_M1020_g N_A_1188_47#_c_1354_n 0.00177777f $X=6.51 $Y=0.415
+ $X2=0 $Y2=0
cc_378 N_A_27_47#_c_270_n N_A_1188_47#_c_1354_n 0.00756683f $X=6.61 $Y=1.19
+ $X2=0 $Y2=0
cc_379 N_A_27_47#_c_274_n N_A_1188_47#_c_1354_n 0.0344296f $X=6.57 $Y=1.11 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_c_260_n N_A_1188_47#_c_1358_n 0.00218f $X=6.32 $Y=1.395 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_c_282_n N_A_1188_47#_c_1358_n 0.0024443f $X=6.32 $Y=1.89 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_c_274_n N_A_1188_47#_c_1358_n 7.37494e-19 $X=6.57 $Y=1.11
+ $X2=0 $Y2=0
cc_383 N_A_27_47#_c_284_n N_VPWR_M1004_d 0.001889f $X=0.66 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_384 N_A_27_47#_c_276_n N_VPWR_c_1454_n 0.00960497f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_284_n N_VPWR_c_1454_n 0.0213487f $X=0.66 $Y=1.88 $X2=0 $Y2=0
cc_386 N_A_27_47#_c_285_n N_VPWR_c_1454_n 0.0254007f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_387 N_A_27_47#_c_283_n N_VPWR_c_1457_n 0.00107286f $X=6.32 $Y=1.99 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_c_283_n N_VPWR_c_1465_n 0.00632161f $X=6.32 $Y=1.99 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_c_284_n N_VPWR_c_1473_n 0.00180073f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_c_285_n N_VPWR_c_1473_n 0.0181185f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_391 N_A_27_47#_c_276_n N_VPWR_c_1474_n 0.00590576f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_280_n N_VPWR_c_1475_n 0.00431504f $X=3.405 $Y=1.99 $X2=0
+ $Y2=0
cc_393 N_A_27_47#_c_276_n N_VPWR_c_1453_n 0.00986661f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_c_280_n N_VPWR_c_1453_n 0.00680728f $X=3.405 $Y=1.99 $X2=0
+ $Y2=0
cc_395 N_A_27_47#_c_283_n N_VPWR_c_1453_n 0.00752369f $X=6.32 $Y=1.99 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_c_284_n N_VPWR_c_1453_n 0.00528325f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_c_285_n N_VPWR_c_1453_n 0.00973967f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_c_256_n N_A_468_47#_c_1624_n 3.34213e-19 $X=2.817 $Y=1.245
+ $X2=0 $Y2=0
cc_399 N_A_27_47#_M1007_g N_A_468_47#_c_1624_n 0.00157198f $X=2.84 $Y=0.415
+ $X2=0 $Y2=0
cc_400 N_A_27_47#_c_265_n N_A_468_47#_c_1624_n 0.0214246f $X=2.535 $Y=1.19 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_c_268_n N_A_468_47#_c_1624_n 0.00250208f $X=2.825 $Y=1.19
+ $X2=0 $Y2=0
cc_402 N_A_27_47#_c_272_n N_A_468_47#_c_1624_n 3.66345e-19 $X=2.735 $Y=0.93
+ $X2=0 $Y2=0
cc_403 N_A_27_47#_c_273_n N_A_468_47#_c_1624_n 0.0378917f $X=2.735 $Y=0.93 $X2=0
+ $Y2=0
cc_404 N_A_27_47#_M1007_g N_A_468_47#_c_1632_n 0.00181198f $X=2.84 $Y=0.415
+ $X2=0 $Y2=0
cc_405 N_A_27_47#_c_268_n N_A_468_47#_c_1632_n 6.44071e-19 $X=2.825 $Y=1.19
+ $X2=0 $Y2=0
cc_406 N_A_27_47#_c_272_n N_A_468_47#_c_1632_n 5.66878e-19 $X=2.735 $Y=0.93
+ $X2=0 $Y2=0
cc_407 N_A_27_47#_c_273_n N_A_468_47#_c_1632_n 0.00672775f $X=2.735 $Y=0.93
+ $X2=0 $Y2=0
cc_408 N_A_27_47#_c_280_n N_A_699_413#_c_1659_n 6.16934e-19 $X=3.405 $Y=1.99
+ $X2=0 $Y2=0
cc_409 N_A_27_47#_c_267_n N_A_699_413#_c_1660_n 3.42555e-19 $X=6.465 $Y=1.19
+ $X2=0 $Y2=0
cc_410 N_A_27_47#_c_279_n N_A_699_413#_c_1661_n 3.38294e-19 $X=3.405 $Y=1.89
+ $X2=0 $Y2=0
cc_411 N_A_27_47#_c_263_n N_VGND_M1021_d 0.00227127f $X=0.66 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_412 N_A_27_47#_M1002_g N_VGND_c_1775_n 0.00430756f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_413 N_A_27_47#_M1002_g N_VGND_c_1781_n 0.00585385f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_414 N_A_27_47#_c_262_n N_VGND_c_1789_n 0.0109767f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_415 N_A_27_47#_c_263_n N_VGND_c_1789_n 0.00244154f $X=0.66 $Y=0.72 $X2=0
+ $Y2=0
cc_416 N_A_27_47#_M1007_g N_VGND_c_1790_n 0.00585385f $X=2.84 $Y=0.415 $X2=0
+ $Y2=0
cc_417 N_A_27_47#_c_272_n N_VGND_c_1790_n 6.34045e-19 $X=2.735 $Y=0.93 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_M1020_g N_VGND_c_1791_n 0.00357877f $X=6.51 $Y=0.415 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_M1021_s N_VGND_c_1793_n 0.00296179f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_M1002_g N_VGND_c_1793_n 0.0120602f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_M1007_g N_VGND_c_1793_n 0.00679961f $X=2.84 $Y=0.415 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_M1020_g N_VGND_c_1793_n 0.00609857f $X=6.51 $Y=0.415 $X2=0
+ $Y2=0
cc_423 N_A_27_47#_c_262_n N_VGND_c_1793_n 0.00916732f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_424 N_A_27_47#_c_263_n N_VGND_c_1793_n 0.00625251f $X=0.66 $Y=0.72 $X2=0
+ $Y2=0
cc_425 N_A_27_47#_c_273_n N_VGND_c_1793_n 0.00906336f $X=2.735 $Y=0.93 $X2=0
+ $Y2=0
cc_426 N_A_27_47#_M1002_g N_VGND_c_1794_n 0.00317372f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_427 N_A_27_47#_c_262_n N_VGND_c_1794_n 0.00923148f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_c_263_n N_VGND_c_1794_n 0.0224548f $X=0.66 $Y=0.72 $X2=0 $Y2=0
cc_429 N_A_27_47#_c_266_n N_VGND_c_1794_n 9.39106e-19 $X=0.89 $Y=1.19 $X2=0
+ $Y2=0
cc_430 N_A_27_47#_c_271_n N_VGND_c_1794_n 6.78636e-19 $X=0.99 $Y=1.235 $X2=0
+ $Y2=0
cc_431 N_D_c_503_n N_A_211_363#_c_564_n 0.00444468f $X=2.35 $Y=1.89 $X2=0 $Y2=0
cc_432 N_D_c_504_n N_A_211_363#_c_564_n 0.00923409f $X=2.35 $Y=1.99 $X2=0 $Y2=0
cc_433 N_D_c_506_n N_A_211_363#_c_564_n 0.0156064f $X=2.19 $Y=1.3 $X2=0 $Y2=0
cc_434 N_D_c_506_n N_A_211_363#_c_558_n 0.00237908f $X=2.19 $Y=1.3 $X2=0 $Y2=0
cc_435 N_D_c_503_n N_A_211_363#_c_570_n 0.00196547f $X=2.35 $Y=1.89 $X2=0 $Y2=0
cc_436 N_D_c_501_n N_A_211_363#_c_570_n 0.0029768f $X=2.19 $Y=1.465 $X2=0 $Y2=0
cc_437 D N_A_211_363#_c_570_n 0.0272612f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_438 N_D_c_502_n N_A_211_363#_c_570_n 0.0072231f $X=1.89 $Y=1.465 $X2=0 $Y2=0
cc_439 D N_A_211_363#_c_571_n 0.00287144f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_440 N_D_c_506_n N_A_211_363#_c_574_n 0.00150989f $X=2.19 $Y=1.3 $X2=0 $Y2=0
cc_441 N_D_c_501_n N_A_211_363#_c_563_n 6.86957e-19 $X=2.19 $Y=1.465 $X2=0 $Y2=0
cc_442 N_D_c_502_n N_A_211_363#_c_563_n 0.143829f $X=1.89 $Y=1.465 $X2=0 $Y2=0
cc_443 N_D_c_504_n N_VPWR_c_1455_n 0.00593401f $X=2.35 $Y=1.99 $X2=0 $Y2=0
cc_444 N_D_c_501_n N_VPWR_c_1455_n 0.00539813f $X=2.19 $Y=1.465 $X2=0 $Y2=0
cc_445 D N_VPWR_c_1455_n 0.0224013f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_446 N_D_c_502_n N_VPWR_c_1455_n 4.34793e-19 $X=1.89 $Y=1.465 $X2=0 $Y2=0
cc_447 D N_VPWR_c_1474_n 0.0211539f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_448 N_D_c_504_n N_VPWR_c_1475_n 0.00518883f $X=2.35 $Y=1.99 $X2=0 $Y2=0
cc_449 N_D_c_504_n N_VPWR_c_1453_n 0.00779061f $X=2.35 $Y=1.99 $X2=0 $Y2=0
cc_450 D N_VPWR_c_1453_n 0.00588351f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_451 N_D_M1012_g N_A_468_47#_c_1624_n 0.0289233f $X=2.265 $Y=0.445 $X2=0 $Y2=0
cc_452 N_D_c_503_n N_A_468_47#_c_1624_n 0.0124776f $X=2.35 $Y=1.89 $X2=0 $Y2=0
cc_453 N_D_c_504_n N_A_468_47#_c_1624_n 0.0176479f $X=2.35 $Y=1.99 $X2=0 $Y2=0
cc_454 N_D_c_501_n N_A_468_47#_c_1624_n 0.00782245f $X=2.19 $Y=1.465 $X2=0 $Y2=0
cc_455 N_D_c_506_n N_A_468_47#_c_1624_n 0.013406f $X=2.19 $Y=1.3 $X2=0 $Y2=0
cc_456 D N_A_468_47#_c_1624_n 0.018973f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_457 N_D_c_502_n N_A_468_47#_c_1624_n 0.0803286f $X=1.89 $Y=1.465 $X2=0 $Y2=0
cc_458 N_D_M1012_g N_A_468_47#_c_1643_n 0.00588428f $X=2.265 $Y=0.445 $X2=0
+ $Y2=0
cc_459 N_D_M1012_g N_A_468_47#_c_1632_n 0.00163056f $X=2.265 $Y=0.445 $X2=0
+ $Y2=0
cc_460 N_D_c_502_n N_VGND_M1012_s 0.00431286f $X=1.89 $Y=1.465 $X2=0 $Y2=0
cc_461 N_D_M1012_g N_VGND_c_1775_n 0.00675175f $X=2.265 $Y=0.445 $X2=0 $Y2=0
cc_462 N_D_c_502_n N_VGND_c_1775_n 0.0275242f $X=1.89 $Y=1.465 $X2=0 $Y2=0
cc_463 N_D_c_502_n N_VGND_c_1781_n 0.00399177f $X=1.89 $Y=1.465 $X2=0 $Y2=0
cc_464 N_D_M1012_g N_VGND_c_1790_n 0.00367956f $X=2.265 $Y=0.445 $X2=0 $Y2=0
cc_465 N_D_M1012_g N_VGND_c_1793_n 0.00698416f $X=2.265 $Y=0.445 $X2=0 $Y2=0
cc_466 N_D_c_502_n N_VGND_c_1793_n 0.00753394f $X=1.89 $Y=1.465 $X2=0 $Y2=0
cc_467 N_A_211_363#_c_568_n N_A_811_289#_M1022_d 2.38738e-19 $X=6.47 $Y=1.58
+ $X2=0 $Y2=0
cc_468 N_A_211_363#_c_569_n N_A_811_289#_M1022_d 0.00214136f $X=6.125 $Y=1.58
+ $X2=0 $Y2=0
cc_469 N_A_211_363#_c_572_n N_A_811_289#_M1022_d 0.00268622f $X=6.465 $Y=1.87
+ $X2=0 $Y2=0
cc_470 N_A_211_363#_c_572_n N_A_811_289#_c_768_n 0.00537127f $X=6.465 $Y=1.87
+ $X2=0 $Y2=0
cc_471 N_A_211_363#_c_562_n N_A_811_289#_M1001_g 0.00294296f $X=3.37 $Y=0.9
+ $X2=0 $Y2=0
cc_472 N_A_211_363#_c_572_n N_A_811_289#_c_770_n 0.0242473f $X=6.465 $Y=1.87
+ $X2=0 $Y2=0
cc_473 N_A_211_363#_c_557_n N_A_811_289#_c_791_n 0.00372135f $X=5.865 $Y=0.705
+ $X2=0 $Y2=0
cc_474 N_A_211_363#_c_569_n N_A_811_289#_c_767_n 0.00184581f $X=6.125 $Y=1.58
+ $X2=0 $Y2=0
cc_475 N_A_211_363#_c_572_n N_A_811_289#_c_793_n 0.00749812f $X=6.465 $Y=1.87
+ $X2=0 $Y2=0
cc_476 N_A_211_363#_c_569_n N_A_811_289#_c_780_n 0.0139294f $X=6.125 $Y=1.58
+ $X2=0 $Y2=0
cc_477 N_A_211_363#_c_572_n N_A_811_289#_c_780_n 0.0205959f $X=6.465 $Y=1.87
+ $X2=0 $Y2=0
cc_478 N_A_211_363#_c_575_n N_A_811_289#_c_780_n 0.00182733f $X=6.61 $Y=1.87
+ $X2=0 $Y2=0
cc_479 N_A_211_363#_c_576_n N_A_811_289#_c_780_n 0.00405794f $X=6.815 $Y=1.74
+ $X2=0 $Y2=0
cc_480 N_A_211_363#_c_572_n N_A_811_289#_c_798_n 0.00708567f $X=6.465 $Y=1.87
+ $X2=0 $Y2=0
cc_481 N_A_211_363#_c_559_n N_A_811_289#_c_784_n 0.0432669f $X=6.04 $Y=0.87
+ $X2=0 $Y2=0
cc_482 N_A_211_363#_c_560_n N_A_811_289#_c_784_n 0.00372135f $X=6.04 $Y=0.87
+ $X2=0 $Y2=0
cc_483 N_A_211_363#_c_569_n N_A_811_289#_c_772_n 0.008521f $X=6.125 $Y=1.58
+ $X2=0 $Y2=0
cc_484 N_A_211_363#_c_572_n N_RESET_B_c_872_n 0.00331104f $X=6.465 $Y=1.87 $X2=0
+ $Y2=0
cc_485 N_A_211_363#_c_559_n N_RESET_B_c_876_n 0.0130979f $X=6.04 $Y=0.87 $X2=0
+ $Y2=0
cc_486 N_A_211_363#_c_560_n N_RESET_B_c_876_n 0.00531637f $X=6.04 $Y=0.87 $X2=0
+ $Y2=0
cc_487 N_A_211_363#_c_557_n N_A_583_47#_M1032_g 0.0104372f $X=5.865 $Y=0.705
+ $X2=0 $Y2=0
cc_488 N_A_211_363#_c_559_n N_A_583_47#_c_1032_n 8.45489e-19 $X=6.04 $Y=0.87
+ $X2=0 $Y2=0
cc_489 N_A_211_363#_c_560_n N_A_583_47#_c_1032_n 0.00332535f $X=6.04 $Y=0.87
+ $X2=0 $Y2=0
cc_490 N_A_211_363#_c_569_n N_A_583_47#_c_1032_n 9.50091e-19 $X=6.125 $Y=1.58
+ $X2=0 $Y2=0
cc_491 N_A_211_363#_c_572_n N_A_583_47#_c_1032_n 2.73565e-19 $X=6.465 $Y=1.87
+ $X2=0 $Y2=0
cc_492 N_A_211_363#_c_569_n N_A_583_47#_c_1033_n 9.06082e-19 $X=6.125 $Y=1.58
+ $X2=0 $Y2=0
cc_493 N_A_211_363#_c_572_n N_A_583_47#_c_1033_n 0.00310577f $X=6.465 $Y=1.87
+ $X2=0 $Y2=0
cc_494 N_A_211_363#_c_564_n N_A_583_47#_c_1043_n 0.00489371f $X=2.86 $Y=1.99
+ $X2=0 $Y2=0
cc_495 N_A_211_363#_c_570_n N_A_583_47#_c_1043_n 5.02408e-19 $X=3.045 $Y=1.87
+ $X2=0 $Y2=0
cc_496 N_A_211_363#_c_572_n N_A_583_47#_c_1043_n 0.00443579f $X=6.465 $Y=1.87
+ $X2=0 $Y2=0
cc_497 N_A_211_363#_c_573_n N_A_583_47#_c_1043_n 0.00467362f $X=3.335 $Y=1.87
+ $X2=0 $Y2=0
cc_498 N_A_211_363#_c_574_n N_A_583_47#_c_1043_n 0.0211562f $X=3.19 $Y=1.87
+ $X2=0 $Y2=0
cc_499 N_A_211_363#_M1014_g N_A_583_47#_c_1066_n 0.0103152f $X=3.37 $Y=0.415
+ $X2=0 $Y2=0
cc_500 N_A_211_363#_c_561_n N_A_583_47#_c_1066_n 0.0142946f $X=3.295 $Y=0.9
+ $X2=0 $Y2=0
cc_501 N_A_211_363#_c_562_n N_A_583_47#_c_1066_n 0.00423748f $X=3.37 $Y=0.9
+ $X2=0 $Y2=0
cc_502 N_A_211_363#_c_564_n N_A_583_47#_c_1034_n 4.10445e-19 $X=2.86 $Y=1.99
+ $X2=0 $Y2=0
cc_503 N_A_211_363#_c_558_n N_A_583_47#_c_1034_n 0.0127937f $X=3.19 $Y=1.575
+ $X2=0 $Y2=0
cc_504 N_A_211_363#_c_572_n N_A_583_47#_c_1034_n 0.0160321f $X=6.465 $Y=1.87
+ $X2=0 $Y2=0
cc_505 N_A_211_363#_c_573_n N_A_583_47#_c_1034_n 0.0026155f $X=3.335 $Y=1.87
+ $X2=0 $Y2=0
cc_506 N_A_211_363#_c_574_n N_A_583_47#_c_1034_n 0.0223887f $X=3.19 $Y=1.87
+ $X2=0 $Y2=0
cc_507 N_A_211_363#_M1014_g N_A_583_47#_c_1027_n 0.0092269f $X=3.37 $Y=0.415
+ $X2=0 $Y2=0
cc_508 N_A_211_363#_c_558_n N_A_583_47#_c_1027_n 0.0072769f $X=3.19 $Y=1.575
+ $X2=0 $Y2=0
cc_509 N_A_211_363#_c_561_n N_A_583_47#_c_1027_n 0.0167253f $X=3.295 $Y=0.9
+ $X2=0 $Y2=0
cc_510 N_A_211_363#_c_562_n N_A_583_47#_c_1027_n 0.00159498f $X=3.37 $Y=0.9
+ $X2=0 $Y2=0
cc_511 N_A_211_363#_c_558_n N_A_583_47#_c_1029_n 0.00987668f $X=3.19 $Y=1.575
+ $X2=0 $Y2=0
cc_512 N_A_211_363#_c_561_n N_A_583_47#_c_1029_n 7.96251e-19 $X=3.295 $Y=0.9
+ $X2=0 $Y2=0
cc_513 N_A_211_363#_c_572_n N_A_583_47#_c_1029_n 0.00764593f $X=6.465 $Y=1.87
+ $X2=0 $Y2=0
cc_514 N_A_211_363#_c_560_n N_A_583_47#_c_1031_n 0.0104372f $X=6.04 $Y=0.87
+ $X2=0 $Y2=0
cc_515 N_A_211_363#_c_565_n N_A_1403_21#_c_1155_n 0.0154755f $X=6.85 $Y=1.99
+ $X2=0 $Y2=0
cc_516 N_A_211_363#_c_576_n N_A_1403_21#_c_1155_n 0.00174759f $X=6.815 $Y=1.74
+ $X2=0 $Y2=0
cc_517 N_A_211_363#_c_565_n N_A_1403_21#_c_1171_n 0.0255792f $X=6.85 $Y=1.99
+ $X2=0 $Y2=0
cc_518 N_A_211_363#_c_557_n N_A_1188_47#_c_1360_n 0.00378498f $X=5.865 $Y=0.705
+ $X2=0 $Y2=0
cc_519 N_A_211_363#_c_559_n N_A_1188_47#_c_1360_n 0.00639761f $X=6.04 $Y=0.87
+ $X2=0 $Y2=0
cc_520 N_A_211_363#_c_560_n N_A_1188_47#_c_1360_n 0.0026746f $X=6.04 $Y=0.87
+ $X2=0 $Y2=0
cc_521 N_A_211_363#_c_565_n N_A_1188_47#_c_1363_n 0.0151193f $X=6.85 $Y=1.99
+ $X2=0 $Y2=0
cc_522 N_A_211_363#_c_568_n N_A_1188_47#_c_1363_n 0.00138883f $X=6.47 $Y=1.58
+ $X2=0 $Y2=0
cc_523 N_A_211_363#_c_572_n N_A_1188_47#_c_1363_n 0.00160054f $X=6.465 $Y=1.87
+ $X2=0 $Y2=0
cc_524 N_A_211_363#_c_575_n N_A_1188_47#_c_1363_n 0.00397729f $X=6.61 $Y=1.87
+ $X2=0 $Y2=0
cc_525 N_A_211_363#_c_576_n N_A_1188_47#_c_1363_n 0.0355415f $X=6.815 $Y=1.74
+ $X2=0 $Y2=0
cc_526 N_A_211_363#_c_565_n N_A_1188_47#_c_1357_n 0.00292771f $X=6.85 $Y=1.99
+ $X2=0 $Y2=0
cc_527 N_A_211_363#_c_575_n N_A_1188_47#_c_1357_n 0.00198562f $X=6.61 $Y=1.87
+ $X2=0 $Y2=0
cc_528 N_A_211_363#_c_576_n N_A_1188_47#_c_1357_n 0.0138125f $X=6.815 $Y=1.74
+ $X2=0 $Y2=0
cc_529 N_A_211_363#_c_565_n N_A_1188_47#_c_1358_n 0.00211311f $X=6.85 $Y=1.99
+ $X2=0 $Y2=0
cc_530 N_A_211_363#_c_576_n N_A_1188_47#_c_1358_n 0.0183661f $X=6.815 $Y=1.74
+ $X2=0 $Y2=0
cc_531 N_A_211_363#_c_572_n N_VPWR_M1022_s 0.00227884f $X=6.465 $Y=1.87 $X2=0
+ $Y2=0
cc_532 N_A_211_363#_c_563_n N_VPWR_c_1454_n 0.0202126f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_533 N_A_211_363#_c_570_n N_VPWR_c_1455_n 0.00658376f $X=3.045 $Y=1.87 $X2=0
+ $Y2=0
cc_534 N_A_211_363#_c_563_n N_VPWR_c_1455_n 4.4131e-19 $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_535 N_A_211_363#_c_572_n N_VPWR_c_1456_n 0.0013967f $X=6.465 $Y=1.87 $X2=0
+ $Y2=0
cc_536 N_A_211_363#_c_572_n N_VPWR_c_1457_n 0.0040303f $X=6.465 $Y=1.87 $X2=0
+ $Y2=0
cc_537 N_A_211_363#_c_565_n N_VPWR_c_1465_n 0.00429453f $X=6.85 $Y=1.99 $X2=0
+ $Y2=0
cc_538 N_A_211_363#_c_563_n N_VPWR_c_1474_n 0.0120448f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_539 N_A_211_363#_c_564_n N_VPWR_c_1475_n 0.00536466f $X=2.86 $Y=1.99 $X2=0
+ $Y2=0
cc_540 N_A_211_363#_c_574_n N_VPWR_c_1475_n 0.00232657f $X=3.19 $Y=1.87 $X2=0
+ $Y2=0
cc_541 N_A_211_363#_c_564_n N_VPWR_c_1453_n 0.00746423f $X=2.86 $Y=1.99 $X2=0
+ $Y2=0
cc_542 N_A_211_363#_c_565_n N_VPWR_c_1453_n 0.00634125f $X=6.85 $Y=1.99 $X2=0
+ $Y2=0
cc_543 N_A_211_363#_c_570_n N_VPWR_c_1453_n 0.0805781f $X=3.045 $Y=1.87 $X2=0
+ $Y2=0
cc_544 N_A_211_363#_c_571_n N_VPWR_c_1453_n 0.0182006f $X=1.345 $Y=1.87 $X2=0
+ $Y2=0
cc_545 N_A_211_363#_c_572_n N_VPWR_c_1453_n 0.145789f $X=6.465 $Y=1.87 $X2=0
+ $Y2=0
cc_546 N_A_211_363#_c_573_n N_VPWR_c_1453_n 0.0159704f $X=3.335 $Y=1.87 $X2=0
+ $Y2=0
cc_547 N_A_211_363#_c_574_n N_VPWR_c_1453_n 0.00188924f $X=3.19 $Y=1.87 $X2=0
+ $Y2=0
cc_548 N_A_211_363#_c_575_n N_VPWR_c_1453_n 0.0186106f $X=6.61 $Y=1.87 $X2=0
+ $Y2=0
cc_549 N_A_211_363#_c_563_n N_VPWR_c_1453_n 0.0029375f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_550 N_A_211_363#_c_564_n N_A_468_47#_c_1624_n 0.00490509f $X=2.86 $Y=1.99
+ $X2=0 $Y2=0
cc_551 N_A_211_363#_c_570_n N_A_468_47#_c_1624_n 0.0311285f $X=3.045 $Y=1.87
+ $X2=0 $Y2=0
cc_552 N_A_211_363#_c_573_n N_A_468_47#_c_1624_n 9.63027e-19 $X=3.335 $Y=1.87
+ $X2=0 $Y2=0
cc_553 N_A_211_363#_c_574_n N_A_468_47#_c_1624_n 0.01769f $X=3.19 $Y=1.87 $X2=0
+ $Y2=0
cc_554 N_A_211_363#_c_572_n N_A_699_413#_c_1660_n 0.032945f $X=6.465 $Y=1.87
+ $X2=0 $Y2=0
cc_555 N_A_211_363#_c_572_n N_A_699_413#_c_1661_n 0.00857493f $X=6.465 $Y=1.87
+ $X2=0 $Y2=0
cc_556 N_A_211_363#_c_563_n N_VGND_c_1775_n 0.00457032f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_557 N_A_211_363#_c_563_n N_VGND_c_1781_n 0.00732874f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_558 N_A_211_363#_M1014_g N_VGND_c_1790_n 0.00368123f $X=3.37 $Y=0.415 $X2=0
+ $Y2=0
cc_559 N_A_211_363#_c_557_n N_VGND_c_1791_n 0.00561318f $X=5.865 $Y=0.705 $X2=0
+ $Y2=0
cc_560 N_A_211_363#_c_559_n N_VGND_c_1791_n 0.00183172f $X=6.04 $Y=0.87 $X2=0
+ $Y2=0
cc_561 N_A_211_363#_c_560_n N_VGND_c_1791_n 3.95442e-19 $X=6.04 $Y=0.87 $X2=0
+ $Y2=0
cc_562 N_A_211_363#_M1002_d N_VGND_c_1793_n 0.00535012f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_563 N_A_211_363#_M1014_g N_VGND_c_1793_n 0.00689722f $X=3.37 $Y=0.415 $X2=0
+ $Y2=0
cc_564 N_A_211_363#_c_557_n N_VGND_c_1793_n 0.0069755f $X=5.865 $Y=0.705 $X2=0
+ $Y2=0
cc_565 N_A_211_363#_c_559_n N_VGND_c_1793_n 0.00156293f $X=6.04 $Y=0.87 $X2=0
+ $Y2=0
cc_566 N_A_211_363#_c_563_n N_VGND_c_1793_n 0.00616598f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_567 N_A_811_289#_c_768_n N_RESET_B_c_872_n 0.0307401f $X=4.155 $Y=1.99 $X2=0
+ $Y2=0
cc_568 N_A_811_289#_M1001_g N_RESET_B_c_872_n 0.0179384f $X=4.25 $Y=0.445 $X2=0
+ $Y2=0
cc_569 N_A_811_289#_c_770_n N_RESET_B_c_872_n 0.0136984f $X=5.505 $Y=1.61 $X2=0
+ $Y2=0
cc_570 N_A_811_289#_c_768_n N_RESET_B_c_886_n 0.0135184f $X=4.155 $Y=1.99 $X2=0
+ $Y2=0
cc_571 N_A_811_289#_M1001_g N_RESET_B_c_875_n 0.00261071f $X=4.25 $Y=0.445 $X2=0
+ $Y2=0
cc_572 N_A_811_289#_M1032_d N_RESET_B_c_876_n 3.28012e-19 $X=5.445 $Y=0.235
+ $X2=0 $Y2=0
cc_573 N_A_811_289#_c_770_n N_RESET_B_c_876_n 3.07379e-19 $X=5.505 $Y=1.61 $X2=0
+ $Y2=0
cc_574 N_A_811_289#_c_767_n N_RESET_B_c_876_n 0.0072536f $X=5.59 $Y=1.525 $X2=0
+ $Y2=0
cc_575 N_A_811_289#_c_810_p N_RESET_B_c_876_n 0.00227253f $X=5.6 $Y=0.36 $X2=0
+ $Y2=0
cc_576 N_A_811_289#_c_784_n N_RESET_B_c_876_n 0.0147184f $X=5.52 $Y=0.835 $X2=0
+ $Y2=0
cc_577 N_A_811_289#_c_767_n N_RESET_B_c_877_n 2.71757e-19 $X=5.59 $Y=1.525 $X2=0
+ $Y2=0
cc_578 N_A_811_289#_c_784_n N_RESET_B_c_877_n 0.00131338f $X=5.52 $Y=0.835 $X2=0
+ $Y2=0
cc_579 N_A_811_289#_M1001_g N_RESET_B_c_879_n 0.0120484f $X=4.25 $Y=0.445 $X2=0
+ $Y2=0
cc_580 N_A_811_289#_c_767_n N_RESET_B_c_879_n 0.00440619f $X=5.59 $Y=1.525 $X2=0
+ $Y2=0
cc_581 N_A_811_289#_c_784_n N_RESET_B_c_879_n 0.00188953f $X=5.52 $Y=0.835 $X2=0
+ $Y2=0
cc_582 N_A_811_289#_M1001_g N_RESET_B_c_880_n 0.0639035f $X=4.25 $Y=0.445 $X2=0
+ $Y2=0
cc_583 N_A_811_289#_c_810_p N_RESET_B_c_880_n 9.85278e-19 $X=5.6 $Y=0.36 $X2=0
+ $Y2=0
cc_584 N_A_811_289#_c_791_n N_A_583_47#_M1032_g 0.00644998f $X=5.52 $Y=0.68
+ $X2=0 $Y2=0
cc_585 N_A_811_289#_c_767_n N_A_583_47#_M1032_g 0.012632f $X=5.59 $Y=1.525 $X2=0
+ $Y2=0
cc_586 N_A_811_289#_c_810_p N_A_583_47#_M1032_g 0.00331537f $X=5.6 $Y=0.36 $X2=0
+ $Y2=0
cc_587 N_A_811_289#_c_784_n N_A_583_47#_M1032_g 0.0066202f $X=5.52 $Y=0.835
+ $X2=0 $Y2=0
cc_588 N_A_811_289#_c_770_n N_A_583_47#_c_1032_n 0.00207011f $X=5.505 $Y=1.61
+ $X2=0 $Y2=0
cc_589 N_A_811_289#_c_767_n N_A_583_47#_c_1032_n 0.0109981f $X=5.59 $Y=1.525
+ $X2=0 $Y2=0
cc_590 N_A_811_289#_c_780_n N_A_583_47#_c_1032_n 3.99612e-19 $X=5.945 $Y=1.92
+ $X2=0 $Y2=0
cc_591 N_A_811_289#_c_784_n N_A_583_47#_c_1032_n 8.88512e-19 $X=5.52 $Y=0.835
+ $X2=0 $Y2=0
cc_592 N_A_811_289#_c_772_n N_A_583_47#_c_1032_n 0.0049553f $X=5.59 $Y=1.61
+ $X2=0 $Y2=0
cc_593 N_A_811_289#_c_793_n N_A_583_47#_c_1033_n 0.00314949f $X=5.59 $Y=1.835
+ $X2=0 $Y2=0
cc_594 N_A_811_289#_c_780_n N_A_583_47#_c_1033_n 0.0158338f $X=5.945 $Y=1.92
+ $X2=0 $Y2=0
cc_595 N_A_811_289#_c_783_n N_A_583_47#_c_1033_n 0.00472286f $X=6.03 $Y=2.3
+ $X2=0 $Y2=0
cc_596 N_A_811_289#_c_772_n N_A_583_47#_c_1033_n 0.00303318f $X=5.59 $Y=1.61
+ $X2=0 $Y2=0
cc_597 N_A_811_289#_c_768_n N_A_583_47#_c_1043_n 0.00129332f $X=4.155 $Y=1.99
+ $X2=0 $Y2=0
cc_598 N_A_811_289#_M1001_g N_A_583_47#_c_1066_n 0.00592384f $X=4.25 $Y=0.445
+ $X2=0 $Y2=0
cc_599 N_A_811_289#_c_768_n N_A_583_47#_c_1034_n 0.00535568f $X=4.155 $Y=1.99
+ $X2=0 $Y2=0
cc_600 N_A_811_289#_M1001_g N_A_583_47#_c_1034_n 0.00143703f $X=4.25 $Y=0.445
+ $X2=0 $Y2=0
cc_601 N_A_811_289#_c_770_n N_A_583_47#_c_1034_n 0.00842454f $X=5.505 $Y=1.61
+ $X2=0 $Y2=0
cc_602 N_A_811_289#_M1001_g N_A_583_47#_c_1027_n 0.0135473f $X=4.25 $Y=0.445
+ $X2=0 $Y2=0
cc_603 N_A_811_289#_c_768_n N_A_583_47#_c_1028_n 0.00481281f $X=4.155 $Y=1.99
+ $X2=0 $Y2=0
cc_604 N_A_811_289#_M1001_g N_A_583_47#_c_1028_n 0.0110226f $X=4.25 $Y=0.445
+ $X2=0 $Y2=0
cc_605 N_A_811_289#_c_770_n N_A_583_47#_c_1028_n 0.0694522f $X=5.505 $Y=1.61
+ $X2=0 $Y2=0
cc_606 N_A_811_289#_c_770_n N_A_583_47#_c_1030_n 0.0116159f $X=5.505 $Y=1.61
+ $X2=0 $Y2=0
cc_607 N_A_811_289#_c_767_n N_A_583_47#_c_1030_n 0.0196285f $X=5.59 $Y=1.525
+ $X2=0 $Y2=0
cc_608 N_A_811_289#_c_770_n N_A_583_47#_c_1031_n 0.00941249f $X=5.505 $Y=1.61
+ $X2=0 $Y2=0
cc_609 N_A_811_289#_c_791_n N_A_1188_47#_c_1360_n 0.00430859f $X=5.52 $Y=0.68
+ $X2=0 $Y2=0
cc_610 N_A_811_289#_c_783_n N_A_1188_47#_c_1363_n 0.0206717f $X=6.03 $Y=2.3
+ $X2=0 $Y2=0
cc_611 N_A_811_289#_c_770_n N_VPWR_M1022_s 0.00204101f $X=5.505 $Y=1.61 $X2=0
+ $Y2=0
cc_612 N_A_811_289#_c_793_n N_VPWR_M1022_s 0.00454747f $X=5.59 $Y=1.835 $X2=0
+ $Y2=0
cc_613 N_A_811_289#_c_798_n N_VPWR_M1022_s 0.00390064f $X=5.675 $Y=1.92 $X2=0
+ $Y2=0
cc_614 N_A_811_289#_c_768_n N_VPWR_c_1456_n 0.00458065f $X=4.155 $Y=1.99 $X2=0
+ $Y2=0
cc_615 N_A_811_289#_c_770_n N_VPWR_c_1457_n 0.00346475f $X=5.505 $Y=1.61 $X2=0
+ $Y2=0
cc_616 N_A_811_289#_c_780_n N_VPWR_c_1457_n 0.00255212f $X=5.945 $Y=1.92 $X2=0
+ $Y2=0
cc_617 N_A_811_289#_c_798_n N_VPWR_c_1457_n 0.00972897f $X=5.675 $Y=1.92 $X2=0
+ $Y2=0
cc_618 N_A_811_289#_c_783_n N_VPWR_c_1457_n 0.0178901f $X=6.03 $Y=2.3 $X2=0
+ $Y2=0
cc_619 N_A_811_289#_c_780_n N_VPWR_c_1465_n 0.00269374f $X=5.945 $Y=1.92 $X2=0
+ $Y2=0
cc_620 N_A_811_289#_c_783_n N_VPWR_c_1465_n 0.0117479f $X=6.03 $Y=2.3 $X2=0
+ $Y2=0
cc_621 N_A_811_289#_c_768_n N_VPWR_c_1475_n 0.00525574f $X=4.155 $Y=1.99 $X2=0
+ $Y2=0
cc_622 N_A_811_289#_M1022_d N_VPWR_c_1453_n 0.00349593f $X=5.865 $Y=1.645 $X2=0
+ $Y2=0
cc_623 N_A_811_289#_c_768_n N_VPWR_c_1453_n 0.0072085f $X=4.155 $Y=1.99 $X2=0
+ $Y2=0
cc_624 N_A_811_289#_c_780_n N_VPWR_c_1453_n 0.00229794f $X=5.945 $Y=1.92 $X2=0
+ $Y2=0
cc_625 N_A_811_289#_c_798_n N_VPWR_c_1453_n 4.80263e-19 $X=5.675 $Y=1.92 $X2=0
+ $Y2=0
cc_626 N_A_811_289#_c_783_n N_VPWR_c_1453_n 0.00306902f $X=6.03 $Y=2.3 $X2=0
+ $Y2=0
cc_627 N_A_811_289#_c_768_n N_A_699_413#_c_1659_n 0.00428162f $X=4.155 $Y=1.99
+ $X2=0 $Y2=0
cc_628 N_A_811_289#_c_768_n N_A_699_413#_c_1660_n 0.0171824f $X=4.155 $Y=1.99
+ $X2=0 $Y2=0
cc_629 N_A_811_289#_c_770_n N_A_699_413#_c_1660_n 0.0615757f $X=5.505 $Y=1.61
+ $X2=0 $Y2=0
cc_630 N_A_811_289#_c_798_n N_A_699_413#_c_1660_n 0.004407f $X=5.675 $Y=1.92
+ $X2=0 $Y2=0
cc_631 N_A_811_289#_c_810_p N_VGND_c_1776_n 0.0179146f $X=5.6 $Y=0.36 $X2=0
+ $Y2=0
cc_632 N_A_811_289#_M1001_g N_VGND_c_1790_n 0.00585385f $X=4.25 $Y=0.445 $X2=0
+ $Y2=0
cc_633 N_A_811_289#_c_810_p N_VGND_c_1791_n 0.0215212f $X=5.6 $Y=0.36 $X2=0
+ $Y2=0
cc_634 N_A_811_289#_M1032_d N_VGND_c_1793_n 0.00246666f $X=5.445 $Y=0.235 $X2=0
+ $Y2=0
cc_635 N_A_811_289#_M1001_g N_VGND_c_1793_n 0.00693872f $X=4.25 $Y=0.445 $X2=0
+ $Y2=0
cc_636 N_A_811_289#_c_810_p N_VGND_c_1793_n 0.00688009f $X=5.6 $Y=0.36 $X2=0
+ $Y2=0
cc_637 N_RESET_B_c_876_n N_A_583_47#_M1032_g 0.00427213f $X=7.81 $Y=0.85 $X2=0
+ $Y2=0
cc_638 N_RESET_B_c_877_n N_A_583_47#_M1032_g 5.75754e-19 $X=4.925 $Y=0.85 $X2=0
+ $Y2=0
cc_639 N_RESET_B_c_878_n N_A_583_47#_M1032_g 0.00599875f $X=4.67 $Y=0.93 $X2=0
+ $Y2=0
cc_640 N_RESET_B_c_879_n N_A_583_47#_M1032_g 0.00177764f $X=4.67 $Y=0.93 $X2=0
+ $Y2=0
cc_641 N_RESET_B_c_880_n N_A_583_47#_M1032_g 0.0101386f $X=4.695 $Y=0.765 $X2=0
+ $Y2=0
cc_642 N_RESET_B_c_875_n N_A_583_47#_c_1027_n 0.00264594f $X=4.81 $Y=0.85 $X2=0
+ $Y2=0
cc_643 N_RESET_B_c_879_n N_A_583_47#_c_1027_n 0.0086523f $X=4.67 $Y=0.93 $X2=0
+ $Y2=0
cc_644 N_RESET_B_c_872_n N_A_583_47#_c_1028_n 0.0112582f $X=4.69 $Y=1.89 $X2=0
+ $Y2=0
cc_645 N_RESET_B_c_875_n N_A_583_47#_c_1028_n 0.00100061f $X=4.81 $Y=0.85 $X2=0
+ $Y2=0
cc_646 N_RESET_B_c_876_n N_A_583_47#_c_1028_n 8.33479e-19 $X=7.81 $Y=0.85 $X2=0
+ $Y2=0
cc_647 N_RESET_B_c_878_n N_A_583_47#_c_1028_n 0.00314155f $X=4.67 $Y=0.93 $X2=0
+ $Y2=0
cc_648 N_RESET_B_c_879_n N_A_583_47#_c_1028_n 0.0489652f $X=4.67 $Y=0.93 $X2=0
+ $Y2=0
cc_649 N_RESET_B_c_872_n N_A_583_47#_c_1030_n 8.14528e-19 $X=4.69 $Y=1.89 $X2=0
+ $Y2=0
cc_650 N_RESET_B_c_876_n N_A_583_47#_c_1030_n 0.00422691f $X=7.81 $Y=0.85 $X2=0
+ $Y2=0
cc_651 N_RESET_B_c_878_n N_A_583_47#_c_1030_n 5.24882e-19 $X=4.67 $Y=0.93 $X2=0
+ $Y2=0
cc_652 N_RESET_B_c_879_n N_A_583_47#_c_1030_n 7.26099e-19 $X=4.67 $Y=0.93 $X2=0
+ $Y2=0
cc_653 N_RESET_B_c_872_n N_A_583_47#_c_1031_n 0.0192408f $X=4.69 $Y=1.89 $X2=0
+ $Y2=0
cc_654 N_RESET_B_c_876_n N_A_583_47#_c_1031_n 0.00102675f $X=7.81 $Y=0.85 $X2=0
+ $Y2=0
cc_655 N_RESET_B_c_878_n N_A_583_47#_c_1031_n 0.00613982f $X=4.67 $Y=0.93 $X2=0
+ $Y2=0
cc_656 N_RESET_B_c_876_n N_A_1403_21#_M1018_g 0.00105989f $X=7.81 $Y=0.85 $X2=0
+ $Y2=0
cc_657 N_RESET_B_c_873_n N_A_1403_21#_c_1155_n 0.0103479f $X=7.96 $Y=1.89 $X2=0
+ $Y2=0
cc_658 N_RESET_B_c_881_n N_A_1403_21#_c_1155_n 0.00418864f $X=7.97 $Y=1.12 $X2=0
+ $Y2=0
cc_659 N_RESET_B_c_883_n N_A_1403_21#_c_1155_n 0.00218833f $X=8.275 $Y=1.22
+ $X2=0 $Y2=0
cc_660 N_RESET_B_c_888_n N_A_1403_21#_c_1171_n 0.0226527f $X=7.96 $Y=1.99 $X2=0
+ $Y2=0
cc_661 N_RESET_B_M1029_g N_A_1403_21#_c_1160_n 3.49437e-19 $X=7.985 $Y=0.445
+ $X2=0 $Y2=0
cc_662 N_RESET_B_c_876_n N_A_1403_21#_c_1160_n 0.0122038f $X=7.81 $Y=0.85 $X2=0
+ $Y2=0
cc_663 N_RESET_B_c_881_n N_A_1403_21#_c_1160_n 4.11328e-19 $X=7.97 $Y=1.12 $X2=0
+ $Y2=0
cc_664 N_RESET_B_c_882_n N_A_1403_21#_c_1160_n 0.00284943f $X=8.25 $Y=0.85 $X2=0
+ $Y2=0
cc_665 N_RESET_B_c_883_n N_A_1403_21#_c_1160_n 0.00782309f $X=8.275 $Y=1.22
+ $X2=0 $Y2=0
cc_666 RESET_B N_A_1403_21#_c_1160_n 0.0049647f $X=8.055 $Y=1.19 $X2=0 $Y2=0
cc_667 N_RESET_B_M1029_g N_A_1403_21#_c_1161_n 0.00778365f $X=7.985 $Y=0.445
+ $X2=0 $Y2=0
cc_668 N_RESET_B_c_876_n N_A_1403_21#_c_1161_n 4.49559e-19 $X=7.81 $Y=0.85 $X2=0
+ $Y2=0
cc_669 N_RESET_B_c_882_n N_A_1403_21#_c_1161_n 0.00361023f $X=8.25 $Y=0.85 $X2=0
+ $Y2=0
cc_670 N_RESET_B_M1029_g N_A_1403_21#_c_1201_n 0.00869977f $X=7.985 $Y=0.445
+ $X2=0 $Y2=0
cc_671 N_RESET_B_c_881_n N_A_1403_21#_c_1201_n 9.38055e-19 $X=7.97 $Y=1.12 $X2=0
+ $Y2=0
cc_672 N_RESET_B_c_882_n N_A_1403_21#_c_1201_n 0.013814f $X=8.25 $Y=0.85 $X2=0
+ $Y2=0
cc_673 N_RESET_B_c_883_n N_A_1403_21#_c_1201_n 0.00230931f $X=8.275 $Y=1.22
+ $X2=0 $Y2=0
cc_674 RESET_B N_A_1403_21#_c_1201_n 0.00367536f $X=8.055 $Y=1.19 $X2=0 $Y2=0
cc_675 N_RESET_B_M1029_g N_A_1403_21#_c_1206_n 0.00358232f $X=7.985 $Y=0.445
+ $X2=0 $Y2=0
cc_676 N_RESET_B_c_888_n N_A_1403_21#_c_1177_n 0.0026824f $X=7.96 $Y=1.99 $X2=0
+ $Y2=0
cc_677 N_RESET_B_c_882_n N_A_1403_21#_c_1163_n 0.00986473f $X=8.25 $Y=0.85 $X2=0
+ $Y2=0
cc_678 RESET_B N_A_1403_21#_c_1163_n 0.00257461f $X=8.055 $Y=1.19 $X2=0 $Y2=0
cc_679 N_RESET_B_c_882_n N_A_1403_21#_c_1164_n 0.0115715f $X=8.25 $Y=0.85 $X2=0
+ $Y2=0
cc_680 N_RESET_B_c_883_n N_A_1403_21#_c_1164_n 0.015141f $X=8.275 $Y=1.22 $X2=0
+ $Y2=0
cc_681 RESET_B N_A_1403_21#_c_1164_n 0.00895511f $X=8.055 $Y=1.19 $X2=0 $Y2=0
cc_682 N_RESET_B_c_883_n N_A_1403_21#_c_1165_n 0.00502592f $X=8.275 $Y=1.22
+ $X2=0 $Y2=0
cc_683 N_RESET_B_M1029_g N_A_1403_21#_c_1167_n 0.00524996f $X=7.985 $Y=0.445
+ $X2=0 $Y2=0
cc_684 N_RESET_B_c_876_n N_A_1403_21#_c_1167_n 0.0165891f $X=7.81 $Y=0.85 $X2=0
+ $Y2=0
cc_685 N_RESET_B_c_881_n N_A_1403_21#_c_1167_n 0.00152691f $X=7.97 $Y=1.12 $X2=0
+ $Y2=0
cc_686 N_RESET_B_c_882_n N_A_1403_21#_c_1167_n 0.00935406f $X=8.25 $Y=0.85 $X2=0
+ $Y2=0
cc_687 N_RESET_B_c_883_n N_A_1403_21#_c_1167_n 0.00885417f $X=8.275 $Y=1.22
+ $X2=0 $Y2=0
cc_688 RESET_B N_A_1403_21#_c_1167_n 0.00648772f $X=8.055 $Y=1.19 $X2=0 $Y2=0
cc_689 N_RESET_B_M1029_g N_A_1403_21#_c_1168_n 0.00673938f $X=7.985 $Y=0.445
+ $X2=0 $Y2=0
cc_690 N_RESET_B_c_876_n N_A_1403_21#_c_1168_n 0.00444753f $X=7.81 $Y=0.85 $X2=0
+ $Y2=0
cc_691 N_RESET_B_c_881_n N_A_1403_21#_c_1168_n 0.0125386f $X=7.97 $Y=1.12 $X2=0
+ $Y2=0
cc_692 N_RESET_B_c_883_n N_A_1403_21#_c_1168_n 6.63351e-19 $X=8.275 $Y=1.22
+ $X2=0 $Y2=0
cc_693 RESET_B N_A_1403_21#_c_1168_n 0.00215991f $X=8.055 $Y=1.19 $X2=0 $Y2=0
cc_694 N_RESET_B_c_873_n N_A_1188_47#_c_1355_n 0.0305666f $X=7.96 $Y=1.89 $X2=0
+ $Y2=0
cc_695 N_RESET_B_c_888_n N_A_1188_47#_c_1355_n 0.0124449f $X=7.96 $Y=1.99 $X2=0
+ $Y2=0
cc_696 N_RESET_B_c_883_n N_A_1188_47#_c_1355_n 0.00340189f $X=8.275 $Y=1.22
+ $X2=0 $Y2=0
cc_697 N_RESET_B_c_873_n N_A_1188_47#_M1013_g 0.00719773f $X=7.96 $Y=1.89 $X2=0
+ $Y2=0
cc_698 N_RESET_B_M1029_g N_A_1188_47#_M1013_g 0.0274433f $X=7.985 $Y=0.445 $X2=0
+ $Y2=0
cc_699 N_RESET_B_c_881_n N_A_1188_47#_M1013_g 0.014851f $X=7.97 $Y=1.12 $X2=0
+ $Y2=0
cc_700 N_RESET_B_c_882_n N_A_1188_47#_M1013_g 0.00346696f $X=8.25 $Y=0.85 $X2=0
+ $Y2=0
cc_701 N_RESET_B_c_883_n N_A_1188_47#_M1013_g 0.00363598f $X=8.275 $Y=1.22 $X2=0
+ $Y2=0
cc_702 RESET_B N_A_1188_47#_M1013_g 0.00629174f $X=8.055 $Y=1.19 $X2=0 $Y2=0
cc_703 N_RESET_B_c_876_n N_A_1188_47#_c_1360_n 0.0139734f $X=7.81 $Y=0.85 $X2=0
+ $Y2=0
cc_704 N_RESET_B_c_876_n N_A_1188_47#_c_1354_n 0.0197148f $X=7.81 $Y=0.85 $X2=0
+ $Y2=0
cc_705 N_RESET_B_c_883_n N_A_1188_47#_c_1354_n 0.0053446f $X=8.275 $Y=1.22 $X2=0
+ $Y2=0
cc_706 N_RESET_B_c_873_n N_A_1188_47#_c_1357_n 0.00132473f $X=7.96 $Y=1.89 $X2=0
+ $Y2=0
cc_707 N_RESET_B_c_888_n N_A_1188_47#_c_1357_n 7.88452e-19 $X=7.96 $Y=1.99 $X2=0
+ $Y2=0
cc_708 N_RESET_B_c_873_n N_A_1188_47#_c_1358_n 0.00113009f $X=7.96 $Y=1.89 $X2=0
+ $Y2=0
cc_709 N_RESET_B_c_876_n N_A_1188_47#_c_1358_n 0.00810734f $X=7.81 $Y=0.85 $X2=0
+ $Y2=0
cc_710 N_RESET_B_c_883_n N_A_1188_47#_c_1358_n 0.00462059f $X=8.275 $Y=1.22
+ $X2=0 $Y2=0
cc_711 N_RESET_B_c_873_n N_A_1188_47#_c_1359_n 0.0180181f $X=7.96 $Y=1.89 $X2=0
+ $Y2=0
cc_712 N_RESET_B_c_881_n N_A_1188_47#_c_1359_n 6.25544e-19 $X=7.97 $Y=1.12 $X2=0
+ $Y2=0
cc_713 N_RESET_B_c_883_n N_A_1188_47#_c_1359_n 0.0422493f $X=8.275 $Y=1.22 $X2=0
+ $Y2=0
cc_714 RESET_B N_A_1188_47#_c_1359_n 0.00302494f $X=8.055 $Y=1.19 $X2=0 $Y2=0
cc_715 N_RESET_B_c_886_n N_VPWR_c_1456_n 0.0117385f $X=4.69 $Y=1.99 $X2=0 $Y2=0
cc_716 N_RESET_B_c_886_n N_VPWR_c_1457_n 0.00502266f $X=4.69 $Y=1.99 $X2=0 $Y2=0
cc_717 N_RESET_B_c_888_n N_VPWR_c_1458_n 0.00848253f $X=7.96 $Y=1.99 $X2=0 $Y2=0
cc_718 N_RESET_B_c_888_n N_VPWR_c_1459_n 0.00643335f $X=7.96 $Y=1.99 $X2=0 $Y2=0
cc_719 N_RESET_B_c_886_n N_VPWR_c_1463_n 0.0046377f $X=4.69 $Y=1.99 $X2=0 $Y2=0
cc_720 N_RESET_B_c_886_n N_VPWR_c_1453_n 0.0062934f $X=4.69 $Y=1.99 $X2=0 $Y2=0
cc_721 N_RESET_B_c_888_n N_VPWR_c_1453_n 0.0107763f $X=7.96 $Y=1.99 $X2=0 $Y2=0
cc_722 N_RESET_B_c_888_n N_VPWR_c_1481_n 7.58167e-19 $X=7.96 $Y=1.99 $X2=0 $Y2=0
cc_723 N_RESET_B_c_872_n N_A_699_413#_c_1660_n 0.00268737f $X=4.69 $Y=1.89 $X2=0
+ $Y2=0
cc_724 N_RESET_B_c_886_n N_A_699_413#_c_1660_n 0.0117053f $X=4.69 $Y=1.99 $X2=0
+ $Y2=0
cc_725 N_RESET_B_c_886_n N_A_699_413#_c_1662_n 0.00449002f $X=4.69 $Y=1.99 $X2=0
+ $Y2=0
cc_726 N_RESET_B_c_876_n N_VGND_M1003_d 0.00389427f $X=7.81 $Y=0.85 $X2=0 $Y2=0
cc_727 N_RESET_B_c_876_n N_VGND_c_1776_n 0.00368623f $X=7.81 $Y=0.85 $X2=0 $Y2=0
cc_728 N_RESET_B_c_877_n N_VGND_c_1776_n 0.00121322f $X=4.925 $Y=0.85 $X2=0
+ $Y2=0
cc_729 N_RESET_B_c_878_n N_VGND_c_1776_n 4.92937e-19 $X=4.67 $Y=0.93 $X2=0 $Y2=0
cc_730 N_RESET_B_c_879_n N_VGND_c_1776_n 0.00646762f $X=4.67 $Y=0.93 $X2=0 $Y2=0
cc_731 N_RESET_B_c_880_n N_VGND_c_1776_n 0.0112955f $X=4.695 $Y=0.765 $X2=0
+ $Y2=0
cc_732 N_RESET_B_M1029_g N_VGND_c_1777_n 0.00576858f $X=7.985 $Y=0.445 $X2=0
+ $Y2=0
cc_733 N_RESET_B_c_876_n N_VGND_c_1777_n 0.00105f $X=7.81 $Y=0.85 $X2=0 $Y2=0
cc_734 N_RESET_B_M1029_g N_VGND_c_1783_n 0.00366078f $X=7.985 $Y=0.445 $X2=0
+ $Y2=0
cc_735 N_RESET_B_c_878_n N_VGND_c_1790_n 0.00168692f $X=4.67 $Y=0.93 $X2=0 $Y2=0
cc_736 N_RESET_B_c_880_n N_VGND_c_1790_n 0.00585385f $X=4.695 $Y=0.765 $X2=0
+ $Y2=0
cc_737 N_RESET_B_M1029_g N_VGND_c_1793_n 0.00682964f $X=7.985 $Y=0.445 $X2=0
+ $Y2=0
cc_738 N_RESET_B_c_875_n N_VGND_c_1793_n 0.0413081f $X=4.81 $Y=0.85 $X2=0 $Y2=0
cc_739 N_RESET_B_c_876_n N_VGND_c_1793_n 0.15099f $X=7.81 $Y=0.85 $X2=0 $Y2=0
cc_740 N_RESET_B_c_878_n N_VGND_c_1793_n 8.42898e-19 $X=4.67 $Y=0.93 $X2=0 $Y2=0
cc_741 N_RESET_B_c_879_n N_VGND_c_1793_n 0.00720014f $X=4.67 $Y=0.93 $X2=0 $Y2=0
cc_742 N_RESET_B_c_880_n N_VGND_c_1793_n 0.00624118f $X=4.695 $Y=0.765 $X2=0
+ $Y2=0
cc_743 RESET_B N_VGND_c_1793_n 0.0155345f $X=8.055 $Y=1.19 $X2=0 $Y2=0
cc_744 N_RESET_B_c_882_n A_1612_47# 0.00242692f $X=8.25 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_745 N_A_583_47#_c_1033_n N_VPWR_c_1457_n 0.0112655f $X=5.775 $Y=1.57 $X2=0
+ $Y2=0
cc_746 N_A_583_47#_c_1031_n N_VPWR_c_1457_n 0.0015757f $X=5.2 $Y=1.17 $X2=0
+ $Y2=0
cc_747 N_A_583_47#_c_1033_n N_VPWR_c_1465_n 0.00406603f $X=5.775 $Y=1.57 $X2=0
+ $Y2=0
cc_748 N_A_583_47#_c_1043_n N_VPWR_c_1475_n 0.0430883f $X=3.495 $Y=2.3 $X2=0
+ $Y2=0
cc_749 N_A_583_47#_M1025_d N_VPWR_c_1453_n 0.00234191f $X=2.95 $Y=2.065 $X2=0
+ $Y2=0
cc_750 N_A_583_47#_c_1033_n N_VPWR_c_1453_n 0.0046037f $X=5.775 $Y=1.57 $X2=0
+ $Y2=0
cc_751 N_A_583_47#_c_1043_n N_VPWR_c_1453_n 0.0122854f $X=3.495 $Y=2.3 $X2=0
+ $Y2=0
cc_752 N_A_583_47#_c_1043_n N_A_468_47#_c_1624_n 0.0188635f $X=3.495 $Y=2.3
+ $X2=0 $Y2=0
cc_753 N_A_583_47#_c_1043_n N_A_699_413#_M1000_d 0.0048981f $X=3.495 $Y=2.3
+ $X2=-0.19 $Y2=-0.24
cc_754 N_A_583_47#_c_1034_n N_A_699_413#_M1000_d 6.31229e-19 $X=3.58 $Y=2.135
+ $X2=-0.19 $Y2=-0.24
cc_755 N_A_583_47#_c_1043_n N_A_699_413#_c_1659_n 0.019526f $X=3.495 $Y=2.3
+ $X2=0 $Y2=0
cc_756 N_A_583_47#_c_1034_n N_A_699_413#_c_1659_n 0.0072692f $X=3.58 $Y=2.135
+ $X2=0 $Y2=0
cc_757 N_A_583_47#_c_1033_n N_A_699_413#_c_1660_n 0.00132889f $X=5.775 $Y=1.57
+ $X2=0 $Y2=0
cc_758 N_A_583_47#_c_1028_n N_A_699_413#_c_1660_n 4.0432e-19 $X=5.115 $Y=1.27
+ $X2=0 $Y2=0
cc_759 N_A_583_47#_c_1034_n N_A_699_413#_c_1661_n 0.0133171f $X=3.58 $Y=2.135
+ $X2=0 $Y2=0
cc_760 N_A_583_47#_c_1029_n N_A_699_413#_c_1661_n 0.0035943f $X=3.85 $Y=1.27
+ $X2=0 $Y2=0
cc_761 N_A_583_47#_c_1033_n N_A_699_413#_c_1662_n 0.00258461f $X=5.775 $Y=1.57
+ $X2=0 $Y2=0
cc_762 N_A_583_47#_M1032_g N_VGND_c_1776_n 0.00655088f $X=5.37 $Y=0.555 $X2=0
+ $Y2=0
cc_763 N_A_583_47#_c_1028_n N_VGND_c_1776_n 0.00223331f $X=5.115 $Y=1.27 $X2=0
+ $Y2=0
cc_764 N_A_583_47#_c_1030_n N_VGND_c_1776_n 6.77929e-19 $X=5.2 $Y=1.17 $X2=0
+ $Y2=0
cc_765 N_A_583_47#_c_1031_n N_VGND_c_1776_n 0.001314f $X=5.2 $Y=1.17 $X2=0 $Y2=0
cc_766 N_A_583_47#_c_1066_n N_VGND_c_1790_n 0.0411841f $X=3.68 $Y=0.39 $X2=0
+ $Y2=0
cc_767 N_A_583_47#_M1032_g N_VGND_c_1791_n 0.00467644f $X=5.37 $Y=0.555 $X2=0
+ $Y2=0
cc_768 N_A_583_47#_M1007_d N_VGND_c_1793_n 0.00350729f $X=2.915 $Y=0.235 $X2=0
+ $Y2=0
cc_769 N_A_583_47#_M1032_g N_VGND_c_1793_n 0.00663528f $X=5.37 $Y=0.555 $X2=0
+ $Y2=0
cc_770 N_A_583_47#_c_1066_n N_VGND_c_1793_n 0.0321485f $X=3.68 $Y=0.39 $X2=0
+ $Y2=0
cc_771 N_A_583_47#_c_1066_n A_689_47# 0.0149756f $X=3.68 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_772 N_A_583_47#_c_1027_n A_689_47# 0.00616231f $X=3.765 $Y=1.185 $X2=-0.19
+ $Y2=-0.24
cc_773 N_A_1403_21#_c_1176_n N_A_1188_47#_c_1355_n 0.0173951f $X=8.79 $Y=2 $X2=0
+ $Y2=0
cc_774 N_A_1403_21#_c_1177_n N_A_1188_47#_c_1355_n 2.53623e-19 $X=8.28 $Y=2
+ $X2=0 $Y2=0
cc_775 N_A_1403_21#_c_1165_n N_A_1188_47#_c_1355_n 0.00983395f $X=8.875 $Y=1.915
+ $X2=0 $Y2=0
cc_776 N_A_1403_21#_c_1161_n N_A_1188_47#_M1013_g 8.23902e-19 $X=7.85 $Y=0.695
+ $X2=0 $Y2=0
cc_777 N_A_1403_21#_c_1201_n N_A_1188_47#_M1013_g 0.0128617f $X=8.615 $Y=0.38
+ $X2=0 $Y2=0
cc_778 N_A_1403_21#_c_1163_n N_A_1188_47#_M1013_g 0.00384679f $X=8.775 $Y=0.82
+ $X2=0 $Y2=0
cc_779 N_A_1403_21#_c_1164_n N_A_1188_47#_M1013_g 0.0112999f $X=8.875 $Y=1.295
+ $X2=0 $Y2=0
cc_780 N_A_1403_21#_c_1165_n N_A_1188_47#_M1013_g 0.00510833f $X=8.875 $Y=1.915
+ $X2=0 $Y2=0
cc_781 N_A_1403_21#_M1018_g N_A_1188_47#_c_1360_n 0.0107452f $X=7.09 $Y=0.445
+ $X2=0 $Y2=0
cc_782 N_A_1403_21#_c_1161_n N_A_1188_47#_c_1360_n 2.7752e-19 $X=7.85 $Y=0.695
+ $X2=0 $Y2=0
cc_783 N_A_1403_21#_c_1171_n N_A_1188_47#_c_1363_n 0.0139423f $X=7.37 $Y=1.99
+ $X2=0 $Y2=0
cc_784 N_A_1403_21#_M1018_g N_A_1188_47#_c_1354_n 0.00857239f $X=7.09 $Y=0.445
+ $X2=0 $Y2=0
cc_785 N_A_1403_21#_c_1160_n N_A_1188_47#_c_1354_n 0.0160099f $X=7.44 $Y=0.98
+ $X2=0 $Y2=0
cc_786 N_A_1403_21#_c_1161_n N_A_1188_47#_c_1354_n 0.00405007f $X=7.85 $Y=0.695
+ $X2=0 $Y2=0
cc_787 N_A_1403_21#_c_1167_n N_A_1188_47#_c_1354_n 0.00978668f $X=7.85 $Y=0.78
+ $X2=0 $Y2=0
cc_788 N_A_1403_21#_c_1168_n N_A_1188_47#_c_1354_n 0.0114298f $X=7.37 $Y=0.98
+ $X2=0 $Y2=0
cc_789 N_A_1403_21#_c_1155_n N_A_1188_47#_c_1357_n 0.00522009f $X=7.37 $Y=1.89
+ $X2=0 $Y2=0
cc_790 N_A_1403_21#_c_1171_n N_A_1188_47#_c_1357_n 0.00784271f $X=7.37 $Y=1.99
+ $X2=0 $Y2=0
cc_791 N_A_1403_21#_c_1177_n N_A_1188_47#_c_1357_n 0.00506701f $X=8.28 $Y=2
+ $X2=0 $Y2=0
cc_792 N_A_1403_21#_c_1155_n N_A_1188_47#_c_1358_n 0.0205484f $X=7.37 $Y=1.89
+ $X2=0 $Y2=0
cc_793 N_A_1403_21#_c_1160_n N_A_1188_47#_c_1358_n 0.00856004f $X=7.44 $Y=0.98
+ $X2=0 $Y2=0
cc_794 N_A_1403_21#_c_1168_n N_A_1188_47#_c_1358_n 0.00411823f $X=7.37 $Y=0.98
+ $X2=0 $Y2=0
cc_795 N_A_1403_21#_c_1160_n N_A_1188_47#_c_1359_n 0.00570594f $X=7.44 $Y=0.98
+ $X2=0 $Y2=0
cc_796 N_A_1403_21#_c_1176_n N_A_1188_47#_c_1359_n 0.0236443f $X=8.79 $Y=2 $X2=0
+ $Y2=0
cc_797 N_A_1403_21#_c_1177_n N_A_1188_47#_c_1359_n 0.0138731f $X=8.28 $Y=2 $X2=0
+ $Y2=0
cc_798 N_A_1403_21#_c_1164_n N_A_1188_47#_c_1359_n 2.98117e-19 $X=8.875 $Y=1.295
+ $X2=0 $Y2=0
cc_799 N_A_1403_21#_c_1165_n N_A_1188_47#_c_1359_n 0.0141871f $X=8.875 $Y=1.915
+ $X2=0 $Y2=0
cc_800 N_A_1403_21#_c_1168_n N_A_1188_47#_c_1359_n 8.76062e-19 $X=7.37 $Y=0.98
+ $X2=0 $Y2=0
cc_801 N_A_1403_21#_c_1176_n N_VPWR_M1011_d 0.00235763f $X=8.79 $Y=2 $X2=0 $Y2=0
cc_802 N_A_1403_21#_c_1171_n N_VPWR_c_1458_n 0.00380702f $X=7.37 $Y=1.99 $X2=0
+ $Y2=0
cc_803 N_A_1403_21#_c_1255_p N_VPWR_c_1458_n 0.011854f $X=8.195 $Y=2.21 $X2=0
+ $Y2=0
cc_804 N_A_1403_21#_c_1255_p N_VPWR_c_1459_n 0.00725596f $X=8.195 $Y=2.21 $X2=0
+ $Y2=0
cc_805 N_A_1403_21#_c_1176_n N_VPWR_c_1459_n 0.00254414f $X=8.79 $Y=2 $X2=0
+ $Y2=0
cc_806 N_A_1403_21#_c_1172_n N_VPWR_c_1460_n 0.0128545f $X=9.455 $Y=1.41 $X2=0
+ $Y2=0
cc_807 N_A_1403_21#_c_1176_n N_VPWR_c_1460_n 0.0138368f $X=8.79 $Y=2 $X2=0 $Y2=0
cc_808 N_A_1403_21#_c_1165_n N_VPWR_c_1460_n 0.0245886f $X=8.875 $Y=1.915 $X2=0
+ $Y2=0
cc_809 N_A_1403_21#_c_1166_n N_VPWR_c_1460_n 0.00956519f $X=10.63 $Y=1.16 $X2=0
+ $Y2=0
cc_810 N_A_1403_21#_c_1169_n N_VPWR_c_1460_n 2.05489e-19 $X=10.865 $Y=1.202
+ $X2=0 $Y2=0
cc_811 N_A_1403_21#_c_1173_n N_VPWR_c_1461_n 0.00534613f $X=9.925 $Y=1.41 $X2=0
+ $Y2=0
cc_812 N_A_1403_21#_c_1174_n N_VPWR_c_1461_n 0.00571916f $X=10.395 $Y=1.41 $X2=0
+ $Y2=0
cc_813 N_A_1403_21#_c_1175_n N_VPWR_c_1462_n 0.00740098f $X=10.865 $Y=1.41 $X2=0
+ $Y2=0
cc_814 N_A_1403_21#_c_1171_n N_VPWR_c_1465_n 0.00433532f $X=7.37 $Y=1.99 $X2=0
+ $Y2=0
cc_815 N_A_1403_21#_c_1176_n N_VPWR_c_1467_n 0.00242603f $X=8.79 $Y=2 $X2=0
+ $Y2=0
cc_816 N_A_1403_21#_c_1172_n N_VPWR_c_1469_n 0.00702461f $X=9.455 $Y=1.41 $X2=0
+ $Y2=0
cc_817 N_A_1403_21#_c_1173_n N_VPWR_c_1469_n 0.00673617f $X=9.925 $Y=1.41 $X2=0
+ $Y2=0
cc_818 N_A_1403_21#_c_1174_n N_VPWR_c_1471_n 0.00702461f $X=10.395 $Y=1.41 $X2=0
+ $Y2=0
cc_819 N_A_1403_21#_c_1175_n N_VPWR_c_1471_n 0.00702461f $X=10.865 $Y=1.41 $X2=0
+ $Y2=0
cc_820 N_A_1403_21#_M1017_d N_VPWR_c_1453_n 0.00448008f $X=8.05 $Y=2.065 $X2=0
+ $Y2=0
cc_821 N_A_1403_21#_c_1171_n N_VPWR_c_1453_n 0.00654443f $X=7.37 $Y=1.99 $X2=0
+ $Y2=0
cc_822 N_A_1403_21#_c_1172_n N_VPWR_c_1453_n 0.0137919f $X=9.455 $Y=1.41 $X2=0
+ $Y2=0
cc_823 N_A_1403_21#_c_1173_n N_VPWR_c_1453_n 0.0118438f $X=9.925 $Y=1.41 $X2=0
+ $Y2=0
cc_824 N_A_1403_21#_c_1174_n N_VPWR_c_1453_n 0.0125095f $X=10.395 $Y=1.41 $X2=0
+ $Y2=0
cc_825 N_A_1403_21#_c_1175_n N_VPWR_c_1453_n 0.0135275f $X=10.865 $Y=1.41 $X2=0
+ $Y2=0
cc_826 N_A_1403_21#_c_1255_p N_VPWR_c_1453_n 0.00608739f $X=8.195 $Y=2.21 $X2=0
+ $Y2=0
cc_827 N_A_1403_21#_c_1176_n N_VPWR_c_1453_n 0.00984214f $X=8.79 $Y=2 $X2=0
+ $Y2=0
cc_828 N_A_1403_21#_c_1255_p N_VPWR_c_1481_n 0.00857111f $X=8.195 $Y=2.21 $X2=0
+ $Y2=0
cc_829 N_A_1403_21#_c_1176_n N_VPWR_c_1481_n 0.0246484f $X=8.79 $Y=2 $X2=0 $Y2=0
cc_830 N_A_1403_21#_c_1156_n N_Q_c_1710_n 0.00753207f $X=9.48 $Y=0.995 $X2=0
+ $Y2=0
cc_831 N_A_1403_21#_c_1172_n N_Q_c_1704_n 5.00384e-19 $X=9.455 $Y=1.41 $X2=0
+ $Y2=0
cc_832 N_A_1403_21#_c_1173_n N_Q_c_1704_n 8.90899e-19 $X=9.925 $Y=1.41 $X2=0
+ $Y2=0
cc_833 N_A_1403_21#_c_1165_n N_Q_c_1704_n 0.00241233f $X=8.875 $Y=1.915 $X2=0
+ $Y2=0
cc_834 N_A_1403_21#_c_1166_n N_Q_c_1704_n 0.0236329f $X=10.63 $Y=1.16 $X2=0
+ $Y2=0
cc_835 N_A_1403_21#_c_1169_n N_Q_c_1704_n 0.00716774f $X=10.865 $Y=1.202 $X2=0
+ $Y2=0
cc_836 N_A_1403_21#_c_1173_n N_Q_c_1716_n 0.0113204f $X=9.925 $Y=1.41 $X2=0
+ $Y2=0
cc_837 N_A_1403_21#_c_1174_n N_Q_c_1716_n 6.55856e-19 $X=10.395 $Y=1.41 $X2=0
+ $Y2=0
cc_838 N_A_1403_21#_c_1157_n N_Q_c_1698_n 0.0107068f $X=9.95 $Y=0.995 $X2=0
+ $Y2=0
cc_839 N_A_1403_21#_c_1158_n N_Q_c_1698_n 0.0060427f $X=10.42 $Y=0.995 $X2=0
+ $Y2=0
cc_840 N_A_1403_21#_c_1166_n N_Q_c_1698_n 0.0397876f $X=10.63 $Y=1.16 $X2=0
+ $Y2=0
cc_841 N_A_1403_21#_c_1169_n N_Q_c_1698_n 0.00345061f $X=10.865 $Y=1.202 $X2=0
+ $Y2=0
cc_842 N_A_1403_21#_c_1156_n N_Q_c_1699_n 0.00393093f $X=9.48 $Y=0.995 $X2=0
+ $Y2=0
cc_843 N_A_1403_21#_c_1164_n N_Q_c_1699_n 3.52526e-19 $X=8.875 $Y=1.295 $X2=0
+ $Y2=0
cc_844 N_A_1403_21#_c_1166_n N_Q_c_1699_n 0.0306114f $X=10.63 $Y=1.16 $X2=0
+ $Y2=0
cc_845 N_A_1403_21#_c_1169_n N_Q_c_1699_n 0.00358305f $X=10.865 $Y=1.202 $X2=0
+ $Y2=0
cc_846 N_A_1403_21#_c_1173_n N_Q_c_1705_n 0.0137916f $X=9.925 $Y=1.41 $X2=0
+ $Y2=0
cc_847 N_A_1403_21#_c_1174_n N_Q_c_1705_n 0.0156273f $X=10.395 $Y=1.41 $X2=0
+ $Y2=0
cc_848 N_A_1403_21#_c_1166_n N_Q_c_1705_n 0.0458726f $X=10.63 $Y=1.16 $X2=0
+ $Y2=0
cc_849 N_A_1403_21#_c_1169_n N_Q_c_1705_n 0.00807006f $X=10.865 $Y=1.202 $X2=0
+ $Y2=0
cc_850 N_A_1403_21#_c_1157_n N_Q_c_1730_n 6.15855e-19 $X=9.95 $Y=0.995 $X2=0
+ $Y2=0
cc_851 N_A_1403_21#_c_1158_n N_Q_c_1730_n 0.00872696f $X=10.42 $Y=0.995 $X2=0
+ $Y2=0
cc_852 N_A_1403_21#_c_1175_n N_Q_c_1706_n 0.0191333f $X=10.865 $Y=1.41 $X2=0
+ $Y2=0
cc_853 N_A_1403_21#_c_1166_n N_Q_c_1706_n 0.0027931f $X=10.63 $Y=1.16 $X2=0
+ $Y2=0
cc_854 N_A_1403_21#_c_1169_n N_Q_c_1706_n 9.33689e-19 $X=10.865 $Y=1.202 $X2=0
+ $Y2=0
cc_855 N_A_1403_21#_c_1159_n N_Q_c_1700_n 0.0138887f $X=10.89 $Y=0.995 $X2=0
+ $Y2=0
cc_856 N_A_1403_21#_c_1158_n N_Q_c_1701_n 0.00266283f $X=10.42 $Y=0.995 $X2=0
+ $Y2=0
cc_857 N_A_1403_21#_c_1166_n N_Q_c_1701_n 0.0306114f $X=10.63 $Y=1.16 $X2=0
+ $Y2=0
cc_858 N_A_1403_21#_c_1169_n N_Q_c_1701_n 0.00358305f $X=10.865 $Y=1.202 $X2=0
+ $Y2=0
cc_859 N_A_1403_21#_c_1166_n N_Q_c_1707_n 0.0204509f $X=10.63 $Y=1.16 $X2=0
+ $Y2=0
cc_860 N_A_1403_21#_c_1169_n N_Q_c_1707_n 0.00656533f $X=10.865 $Y=1.202 $X2=0
+ $Y2=0
cc_861 N_A_1403_21#_c_1175_n Q 0.00196984f $X=10.865 $Y=1.41 $X2=0 $Y2=0
cc_862 N_A_1403_21#_c_1159_n Q 0.021017f $X=10.89 $Y=0.995 $X2=0 $Y2=0
cc_863 N_A_1403_21#_c_1166_n Q 0.0156912f $X=10.63 $Y=1.16 $X2=0 $Y2=0
cc_864 N_A_1403_21#_c_1161_n N_VGND_M1018_d 0.00285522f $X=7.85 $Y=0.695 $X2=0
+ $Y2=0
cc_865 N_A_1403_21#_c_1206_n N_VGND_M1018_d 0.00263657f $X=7.935 $Y=0.38 $X2=0
+ $Y2=0
cc_866 N_A_1403_21#_M1018_g N_VGND_c_1777_n 0.00937569f $X=7.09 $Y=0.445 $X2=0
+ $Y2=0
cc_867 N_A_1403_21#_c_1161_n N_VGND_c_1777_n 0.00443718f $X=7.85 $Y=0.695 $X2=0
+ $Y2=0
cc_868 N_A_1403_21#_c_1206_n N_VGND_c_1777_n 0.0141597f $X=7.935 $Y=0.38 $X2=0
+ $Y2=0
cc_869 N_A_1403_21#_c_1167_n N_VGND_c_1777_n 0.0171519f $X=7.85 $Y=0.78 $X2=0
+ $Y2=0
cc_870 N_A_1403_21#_c_1168_n N_VGND_c_1777_n 0.00137452f $X=7.37 $Y=0.98 $X2=0
+ $Y2=0
cc_871 N_A_1403_21#_c_1156_n N_VGND_c_1778_n 0.00614193f $X=9.48 $Y=0.995 $X2=0
+ $Y2=0
cc_872 N_A_1403_21#_c_1162_n N_VGND_c_1778_n 0.0125645f $X=8.775 $Y=0.465 $X2=0
+ $Y2=0
cc_873 N_A_1403_21#_c_1163_n N_VGND_c_1778_n 0.0244808f $X=8.775 $Y=0.82 $X2=0
+ $Y2=0
cc_874 N_A_1403_21#_c_1164_n N_VGND_c_1778_n 0.00532529f $X=8.875 $Y=1.295 $X2=0
+ $Y2=0
cc_875 N_A_1403_21#_c_1166_n N_VGND_c_1778_n 0.0137893f $X=10.63 $Y=1.16 $X2=0
+ $Y2=0
cc_876 N_A_1403_21#_c_1169_n N_VGND_c_1778_n 2.29969e-19 $X=10.865 $Y=1.202
+ $X2=0 $Y2=0
cc_877 N_A_1403_21#_c_1157_n N_VGND_c_1779_n 0.00276126f $X=9.95 $Y=0.995 $X2=0
+ $Y2=0
cc_878 N_A_1403_21#_c_1158_n N_VGND_c_1779_n 0.00359159f $X=10.42 $Y=0.995 $X2=0
+ $Y2=0
cc_879 N_A_1403_21#_c_1159_n N_VGND_c_1780_n 0.00438629f $X=10.89 $Y=0.995 $X2=0
+ $Y2=0
cc_880 N_A_1403_21#_c_1201_n N_VGND_c_1783_n 0.0302738f $X=8.615 $Y=0.38 $X2=0
+ $Y2=0
cc_881 N_A_1403_21#_c_1206_n N_VGND_c_1783_n 0.00768187f $X=7.935 $Y=0.38 $X2=0
+ $Y2=0
cc_882 N_A_1403_21#_c_1162_n N_VGND_c_1783_n 0.0178412f $X=8.775 $Y=0.465 $X2=0
+ $Y2=0
cc_883 N_A_1403_21#_c_1167_n N_VGND_c_1783_n 0.00275249f $X=7.85 $Y=0.78 $X2=0
+ $Y2=0
cc_884 N_A_1403_21#_c_1156_n N_VGND_c_1785_n 0.00465454f $X=9.48 $Y=0.995 $X2=0
+ $Y2=0
cc_885 N_A_1403_21#_c_1157_n N_VGND_c_1785_n 0.00439206f $X=9.95 $Y=0.995 $X2=0
+ $Y2=0
cc_886 N_A_1403_21#_c_1158_n N_VGND_c_1787_n 0.00397237f $X=10.42 $Y=0.995 $X2=0
+ $Y2=0
cc_887 N_A_1403_21#_c_1159_n N_VGND_c_1787_n 0.00439206f $X=10.89 $Y=0.995 $X2=0
+ $Y2=0
cc_888 N_A_1403_21#_M1018_g N_VGND_c_1791_n 0.00403211f $X=7.09 $Y=0.445 $X2=0
+ $Y2=0
cc_889 N_A_1403_21#_M1013_d N_VGND_c_1793_n 0.00212393f $X=8.565 $Y=0.235 $X2=0
+ $Y2=0
cc_890 N_A_1403_21#_M1018_g N_VGND_c_1793_n 0.00721829f $X=7.09 $Y=0.445 $X2=0
+ $Y2=0
cc_891 N_A_1403_21#_c_1156_n N_VGND_c_1793_n 0.0092281f $X=9.48 $Y=0.995 $X2=0
+ $Y2=0
cc_892 N_A_1403_21#_c_1157_n N_VGND_c_1793_n 0.00616524f $X=9.95 $Y=0.995 $X2=0
+ $Y2=0
cc_893 N_A_1403_21#_c_1158_n N_VGND_c_1793_n 0.00582631f $X=10.42 $Y=0.995 $X2=0
+ $Y2=0
cc_894 N_A_1403_21#_c_1159_n N_VGND_c_1793_n 0.00710229f $X=10.89 $Y=0.995 $X2=0
+ $Y2=0
cc_895 N_A_1403_21#_c_1201_n N_VGND_c_1793_n 0.0144022f $X=8.615 $Y=0.38 $X2=0
+ $Y2=0
cc_896 N_A_1403_21#_c_1206_n N_VGND_c_1793_n 0.00290541f $X=7.935 $Y=0.38 $X2=0
+ $Y2=0
cc_897 N_A_1403_21#_c_1162_n N_VGND_c_1793_n 0.0120802f $X=8.775 $Y=0.465 $X2=0
+ $Y2=0
cc_898 N_A_1403_21#_c_1167_n N_VGND_c_1793_n 0.00257477f $X=7.85 $Y=0.78 $X2=0
+ $Y2=0
cc_899 N_A_1403_21#_c_1168_n N_VGND_c_1793_n 0.00109336f $X=7.37 $Y=0.98 $X2=0
+ $Y2=0
cc_900 N_A_1403_21#_c_1201_n A_1612_47# 0.00500514f $X=8.615 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_901 N_A_1188_47#_c_1355_n N_VPWR_c_1458_n 7.16012e-19 $X=8.43 $Y=1.99 $X2=0
+ $Y2=0
cc_902 N_A_1188_47#_c_1359_n N_VPWR_c_1458_n 0.00900963f $X=8.405 $Y=1.66 $X2=0
+ $Y2=0
cc_903 N_A_1188_47#_c_1355_n N_VPWR_c_1459_n 0.00343369f $X=8.43 $Y=1.99 $X2=0
+ $Y2=0
cc_904 N_A_1188_47#_c_1355_n N_VPWR_c_1460_n 0.00387762f $X=8.43 $Y=1.99 $X2=0
+ $Y2=0
cc_905 N_A_1188_47#_c_1363_n N_VPWR_c_1465_n 0.0667942f $X=7.25 $Y=2.295 $X2=0
+ $Y2=0
cc_906 N_A_1188_47#_M1028_d N_VPWR_c_1453_n 0.00223064f $X=6.41 $Y=2.065 $X2=0
+ $Y2=0
cc_907 N_A_1188_47#_c_1355_n N_VPWR_c_1453_n 0.00406753f $X=8.43 $Y=1.99 $X2=0
+ $Y2=0
cc_908 N_A_1188_47#_c_1363_n N_VPWR_c_1453_n 0.0313133f $X=7.25 $Y=2.295 $X2=0
+ $Y2=0
cc_909 N_A_1188_47#_c_1355_n N_VPWR_c_1481_n 0.010677f $X=8.43 $Y=1.99 $X2=0
+ $Y2=0
cc_910 N_A_1188_47#_c_1363_n A_1388_413# 0.00624991f $X=7.25 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_911 N_A_1188_47#_c_1360_n N_VGND_c_1777_n 0.0178063f $X=6.965 $Y=0.395 $X2=0
+ $Y2=0
cc_912 N_A_1188_47#_M1013_g N_VGND_c_1778_n 0.00271669f $X=8.49 $Y=0.445 $X2=0
+ $Y2=0
cc_913 N_A_1188_47#_M1013_g N_VGND_c_1783_n 0.00366111f $X=8.49 $Y=0.445 $X2=0
+ $Y2=0
cc_914 N_A_1188_47#_c_1360_n N_VGND_c_1791_n 0.0669774f $X=6.965 $Y=0.395 $X2=0
+ $Y2=0
cc_915 N_A_1188_47#_M1005_d N_VGND_c_1793_n 0.00354884f $X=5.94 $Y=0.235 $X2=0
+ $Y2=0
cc_916 N_A_1188_47#_M1013_g N_VGND_c_1793_n 0.00688669f $X=8.49 $Y=0.445 $X2=0
+ $Y2=0
cc_917 N_A_1188_47#_c_1360_n N_VGND_c_1793_n 0.0188078f $X=6.965 $Y=0.395 $X2=0
+ $Y2=0
cc_918 N_A_1188_47#_c_1360_n A_1317_47# 0.00805453f $X=6.965 $Y=0.395 $X2=-0.19
+ $Y2=-0.24
cc_919 N_VPWR_c_1453_n N_A_468_47#_M1024_d 0.00272455f $X=11.27 $Y=2.72 $X2=0
+ $Y2=0
cc_920 N_VPWR_c_1455_n N_A_468_47#_c_1624_n 0.0221376f $X=2.115 $Y=2.34 $X2=0
+ $Y2=0
cc_921 N_VPWR_c_1475_n N_A_468_47#_c_1624_n 0.0184938f $X=4.29 $Y=2.72 $X2=0
+ $Y2=0
cc_922 N_VPWR_c_1453_n N_A_468_47#_c_1624_n 0.00695694f $X=11.27 $Y=2.72 $X2=0
+ $Y2=0
cc_923 N_VPWR_c_1453_n N_A_699_413#_M1000_d 0.00531344f $X=11.27 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_924 N_VPWR_c_1453_n N_A_699_413#_M1033_d 0.00230036f $X=11.27 $Y=2.72 $X2=0
+ $Y2=0
cc_925 N_VPWR_c_1475_n N_A_699_413#_c_1659_n 0.00730735f $X=4.29 $Y=2.72 $X2=0
+ $Y2=0
cc_926 N_VPWR_c_1453_n N_A_699_413#_c_1659_n 0.00287341f $X=11.27 $Y=2.72 $X2=0
+ $Y2=0
cc_927 N_VPWR_c_1456_n N_A_699_413#_c_1660_n 0.0209399f $X=4.455 $Y=2.29 $X2=0
+ $Y2=0
cc_928 N_VPWR_c_1463_n N_A_699_413#_c_1660_n 0.00330997f $X=5.305 $Y=2.72 $X2=0
+ $Y2=0
cc_929 N_VPWR_c_1475_n N_A_699_413#_c_1660_n 0.00434397f $X=4.29 $Y=2.72 $X2=0
+ $Y2=0
cc_930 N_VPWR_c_1453_n N_A_699_413#_c_1660_n 0.00597125f $X=11.27 $Y=2.72 $X2=0
+ $Y2=0
cc_931 N_VPWR_c_1456_n N_A_699_413#_c_1662_n 0.0102921f $X=4.455 $Y=2.29 $X2=0
+ $Y2=0
cc_932 N_VPWR_c_1457_n N_A_699_413#_c_1662_n 0.010735f $X=5.54 $Y=2.34 $X2=0
+ $Y2=0
cc_933 N_VPWR_c_1463_n N_A_699_413#_c_1662_n 0.00730735f $X=5.305 $Y=2.72 $X2=0
+ $Y2=0
cc_934 N_VPWR_c_1453_n N_A_699_413#_c_1662_n 0.00287341f $X=11.27 $Y=2.72 $X2=0
+ $Y2=0
cc_935 N_VPWR_c_1453_n A_1388_413# 0.00273046f $X=11.27 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_936 N_VPWR_c_1453_n N_Q_M1010_s 0.00300692f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_937 N_VPWR_c_1453_n N_Q_M1019_s 0.00370124f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_938 N_VPWR_c_1461_n N_Q_c_1716_n 0.0401622f $X=10.16 $Y=1.96 $X2=0 $Y2=0
cc_939 N_VPWR_c_1469_n N_Q_c_1716_n 0.0169389f $X=10.075 $Y=2.72 $X2=0 $Y2=0
cc_940 N_VPWR_c_1453_n N_Q_c_1716_n 0.010932f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_941 N_VPWR_M1016_d N_Q_c_1705_n 0.00178587f $X=10.015 $Y=1.485 $X2=0 $Y2=0
cc_942 N_VPWR_c_1461_n N_Q_c_1705_n 0.0136682f $X=10.16 $Y=1.96 $X2=0 $Y2=0
cc_943 N_VPWR_c_1471_n N_Q_c_1751_n 0.0149311f $X=11.015 $Y=2.72 $X2=0 $Y2=0
cc_944 N_VPWR_c_1453_n N_Q_c_1751_n 0.00955092f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_945 N_VPWR_M1026_d N_Q_c_1709_n 0.00678475f $X=10.955 $Y=1.485 $X2=0 $Y2=0
cc_946 N_VPWR_c_1462_n N_Q_c_1709_n 0.0151472f $X=11.1 $Y=1.96 $X2=0 $Y2=0
cc_947 N_A_468_47#_c_1643_n N_VGND_c_1790_n 0.00763796f $X=2.315 $Y=0.39 $X2=0
+ $Y2=0
cc_948 N_A_468_47#_c_1632_n N_VGND_c_1790_n 0.0167809f $X=2.525 $Y=0.39 $X2=0
+ $Y2=0
cc_949 N_A_468_47#_M1012_d N_VGND_c_1793_n 0.00387663f $X=2.34 $Y=0.235 $X2=0
+ $Y2=0
cc_950 N_A_468_47#_c_1643_n N_VGND_c_1793_n 0.00579413f $X=2.315 $Y=0.39 $X2=0
+ $Y2=0
cc_951 N_A_468_47#_c_1632_n N_VGND_c_1793_n 0.0133517f $X=2.525 $Y=0.39 $X2=0
+ $Y2=0
cc_952 N_Q_c_1698_n N_VGND_M1023_d 0.00255557f $X=10.415 $Y=0.82 $X2=0 $Y2=0
cc_953 N_Q_c_1703_n N_VGND_M1031_d 0.00384438f $X=11.2 $Y=0.905 $X2=0 $Y2=0
cc_954 N_Q_c_1710_n N_VGND_c_1778_n 0.0357963f $X=9.69 $Y=0.39 $X2=0 $Y2=0
cc_955 N_Q_c_1699_n N_VGND_c_1778_n 0.0125889f $X=9.855 $Y=0.82 $X2=0 $Y2=0
cc_956 N_Q_c_1698_n N_VGND_c_1779_n 0.012101f $X=10.415 $Y=0.82 $X2=0 $Y2=0
cc_957 N_Q_c_1730_n N_VGND_c_1779_n 0.0223967f $X=10.63 $Y=0.39 $X2=0 $Y2=0
cc_958 N_Q_c_1703_n N_VGND_c_1780_n 0.0133599f $X=11.2 $Y=0.905 $X2=0 $Y2=0
cc_959 N_Q_c_1710_n N_VGND_c_1785_n 0.023074f $X=9.69 $Y=0.39 $X2=0 $Y2=0
cc_960 N_Q_c_1698_n N_VGND_c_1785_n 0.00248202f $X=10.415 $Y=0.82 $X2=0 $Y2=0
cc_961 N_Q_c_1698_n N_VGND_c_1787_n 0.00194552f $X=10.415 $Y=0.82 $X2=0 $Y2=0
cc_962 N_Q_c_1730_n N_VGND_c_1787_n 0.023074f $X=10.63 $Y=0.39 $X2=0 $Y2=0
cc_963 N_Q_c_1700_n N_VGND_c_1787_n 0.00233837f $X=10.995 $Y=0.82 $X2=0 $Y2=0
cc_964 N_Q_c_1703_n N_VGND_c_1792_n 0.00361143f $X=11.2 $Y=0.905 $X2=0 $Y2=0
cc_965 N_Q_M1008_s N_VGND_c_1793_n 0.00264276f $X=9.555 $Y=0.235 $X2=0 $Y2=0
cc_966 N_Q_M1030_s N_VGND_c_1793_n 0.00264276f $X=10.495 $Y=0.235 $X2=0 $Y2=0
cc_967 N_Q_c_1710_n N_VGND_c_1793_n 0.0141066f $X=9.69 $Y=0.39 $X2=0 $Y2=0
cc_968 N_Q_c_1698_n N_VGND_c_1793_n 0.0096764f $X=10.415 $Y=0.82 $X2=0 $Y2=0
cc_969 N_Q_c_1730_n N_VGND_c_1793_n 0.0141066f $X=10.63 $Y=0.39 $X2=0 $Y2=0
cc_970 N_Q_c_1700_n N_VGND_c_1793_n 0.00440153f $X=10.995 $Y=0.82 $X2=0 $Y2=0
cc_971 N_Q_c_1703_n N_VGND_c_1793_n 0.00748596f $X=11.2 $Y=0.905 $X2=0 $Y2=0
cc_972 N_VGND_c_1793_n A_689_47# 0.0172576f $X=11.27 $Y=0 $X2=-0.19 $Y2=-0.24
cc_973 N_VGND_c_1793_n A_865_47# 0.00196925f $X=11.27 $Y=0 $X2=-0.19 $Y2=-0.24
cc_974 N_VGND_c_1793_n A_1317_47# 0.00285232f $X=11.27 $Y=0 $X2=-0.19 $Y2=-0.24
cc_975 N_VGND_c_1793_n A_1612_47# 0.0023207f $X=11.27 $Y=0 $X2=-0.19 $Y2=-0.24
