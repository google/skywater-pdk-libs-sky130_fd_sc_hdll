* NGSPICE file created from sky130_fd_sc_hdll__or4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__or4b_1 A B C D_N VGND VNB VPB VPWR X
M1000 a_117_297# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=6.1845e+11p ps=6.42e+06u
M1001 a_225_297# a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=2.961e+11p pd=3.09e+06u as=0p ps=0u
M1002 X a_225_297# VGND VNB nshort w=650000u l=150000u
+  ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u
M1003 VGND A a_225_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_117_297# D_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=4.241e+11p ps=4.1e+06u
M1005 a_504_297# B a_416_297# VPB phighvt w=420000u l=180000u
+  ad=1.344e+11p pd=1.48e+06u as=1.092e+11p ps=1.36e+06u
M1006 a_225_297# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_504_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND C a_225_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_315_297# a_117_297# a_225_297# VPB phighvt w=420000u l=180000u
+  ad=1.365e+11p pd=1.49e+06u as=1.134e+11p ps=1.38e+06u
M1010 a_416_297# C a_315_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_225_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
.ends

