* File: sky130_fd_sc_hdll__dlxtn_4.pex.spice
* Created: Thu Aug 27 19:06:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__DLXTN_4%GATE_N 4 5 7 8 10 13 19 20 24 26
c41 13 0 2.71124e-20 $X=0.52 $Y=0.805
r42 24 27 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r43 24 26 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r44 19 20 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r45 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r46 11 13 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.52 $Y2=0.805
r47 8 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.805
r48 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.445
r49 5 15 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.495 $Y=1.665
+ $X2=0.305 $Y2=1.665
r50 5 7 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.74
+ $X2=0.495 $Y2=2.135
r51 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r52 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r53 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r54 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_4%A_27_47# 1 2 8 9 11 14 18 19 21 24 28 29
+ 30 35 40 42 50 52 53 54 58 61 64 72
c152 54 0 1.08608e-19 $X=3.115 $Y=1.485
c153 53 0 3.37551e-20 $X=3.26 $Y=1.485
r154 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.48
+ $Y=1.74 $X2=3.48 $Y2=1.74
r155 60 61 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.235
+ $X2=0.99 $Y2=1.235
r156 57 60 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=0.805 $Y=1.235
+ $X2=0.965 $Y2=1.235
r157 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.805
+ $Y=1.235 $X2=0.805 $Y2=1.235
r158 53 68 7.5352 $w=3.88e-07 $l=2.55e-07 $layer=LI1_cond $X=3.37 $Y=1.485
+ $X2=3.37 $Y2=1.74
r159 53 72 5.80039 $w=3.88e-07 $l=7e-08 $layer=LI1_cond $X=3.37 $Y=1.485
+ $X2=3.37 $Y2=1.415
r160 52 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.26 $Y=1.485
+ $X2=3.115 $Y2=1.485
r161 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.26 $Y=1.485
+ $X2=3.26 $Y2=1.485
r162 50 54 2.75371 $w=1.4e-07 $l=2.225e-06 $layer=MET1_cond $X=0.89 $Y=1.53
+ $X2=3.115 $Y2=1.53
r163 48 58 12.5266 $w=2.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.775 $Y=1.485
+ $X2=0.775 $Y2=1.235
r164 47 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.745 $Y=1.485
+ $X2=0.89 $Y2=1.485
r165 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.745 $Y=1.485
+ $X2=0.745 $Y2=1.485
r166 40 64 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.025 $Y=0.87
+ $X2=3.025 $Y2=0.705
r167 39 42 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=3 $Y=0.87 $X2=3.26
+ $Y2=0.87
r168 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3 $Y=0.87
+ $X2=3 $Y2=0.87
r169 37 48 15.5329 $w=2.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.775 $Y=1.795
+ $X2=0.775 $Y2=1.485
r170 36 58 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.775 $Y=0.805
+ $X2=0.775 $Y2=1.235
r171 32 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.26 $Y=1.035
+ $X2=3.26 $Y2=0.87
r172 32 72 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.26 $Y=1.035
+ $X2=3.26 $Y2=1.415
r173 31 35 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r174 30 37 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.66 $Y=1.88
+ $X2=0.775 $Y2=1.795
r175 30 31 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.66 $Y=1.88
+ $X2=0.345 $Y2=1.88
r176 28 36 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.66 $Y=0.72
+ $X2=0.775 $Y2=0.805
r177 28 29 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.66 $Y=0.72
+ $X2=0.345 $Y2=0.72
r178 22 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r179 22 24 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r180 19 67 48.3784 $w=2.91e-07 $l=2.76134e-07 $layer=POLY_cond $X=3.425 $Y=1.99
+ $X2=3.48 $Y2=1.74
r181 19 21 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.425 $Y=1.99
+ $X2=3.425 $Y2=2.275
r182 18 64 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.04 $Y=0.415
+ $X2=3.04 $Y2=0.705
r183 12 61 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=1.235
r184 12 14 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=0.445
r185 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.965 $Y=1.74
+ $X2=0.965 $Y2=2.135
r186 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.64 $X2=0.965
+ $Y2=1.74
r187 7 60 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=0.965 $Y=1.37
+ $X2=0.965 $Y2=1.235
r188 7 8 89.5258 $w=2e-07 $l=2.7e-07 $layer=POLY_cond $X=0.965 $Y=1.37 $X2=0.965
+ $Y2=1.64
r189 2 35 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r190 1 24 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_4%D 2 3 5 8 10 14 17
c43 14 0 1.07926e-19 $X=1.725 $Y=1.04
r44 16 17 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.955 $Y=1.04
+ $X2=1.98 $Y2=1.04
r45 13 16 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=1.725 $Y=1.04
+ $X2=1.955 $Y2=1.04
r46 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.725
+ $Y=1.04 $X2=1.725 $Y2=1.04
r47 10 14 4.16546 $w=4.13e-07 $l=1.5e-07 $layer=LI1_cond $X=1.682 $Y=1.19
+ $X2=1.682 $Y2=1.04
r48 6 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.98 $Y=0.875
+ $X2=1.98 $Y2=1.04
r49 6 8 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.98 $Y=0.875 $X2=1.98
+ $Y2=0.445
r50 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.955 $Y=1.77
+ $X2=1.955 $Y2=2.165
r51 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.955 $Y=1.67 $X2=1.955
+ $Y2=1.77
r52 1 16 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.955 $Y=1.205
+ $X2=1.955 $Y2=1.04
r53 1 2 154.183 $w=2e-07 $l=4.65e-07 $layer=POLY_cond $X=1.955 $Y=1.205
+ $X2=1.955 $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_4%A_319_47# 1 2 8 9 11 14 17 19 21 22 23 24
+ 26 33 35
c90 33 0 1.07926e-19 $X=2.405 $Y=0.93
c91 19 0 7.13094e-20 $X=2.12 $Y=0.7
r92 33 36 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.43 $Y=0.93
+ $X2=2.43 $Y2=1.095
r93 33 35 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.43 $Y=0.93
+ $X2=2.43 $Y2=0.765
r94 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.405
+ $Y=0.93 $X2=2.405 $Y2=0.93
r95 26 28 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.72 $Y=0.51
+ $X2=1.72 $Y2=0.7
r96 23 32 8.96999 $w=3.41e-07 $l=2.18746e-07 $layer=LI1_cond $X=2.205 $Y=1.095
+ $X2=2.33 $Y2=0.93
r97 23 24 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.205 $Y=1.095
+ $X2=2.205 $Y2=1.495
r98 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.12 $Y=1.58
+ $X2=2.205 $Y2=1.495
r99 21 22 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.12 $Y=1.58
+ $X2=1.885 $Y2=1.58
r100 20 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.805 $Y=0.7
+ $X2=1.72 $Y2=0.7
r101 19 32 8.22874 $w=3.41e-07 $l=3.18119e-07 $layer=LI1_cond $X=2.12 $Y=0.7
+ $X2=2.33 $Y2=0.93
r102 19 20 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.12 $Y=0.7
+ $X2=1.805 $Y2=0.7
r103 15 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.72 $Y=1.665
+ $X2=1.885 $Y2=1.58
r104 15 17 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.72 $Y=1.665
+ $X2=1.72 $Y2=1.99
r105 14 35 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.45 $Y=0.445
+ $X2=2.45 $Y2=0.765
r106 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.425 $Y=1.77
+ $X2=2.425 $Y2=2.165
r107 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.425 $Y=1.67 $X2=2.425
+ $Y2=1.77
r108 8 36 190.657 $w=2e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=1.67
+ $X2=2.425 $Y2=1.095
r109 2 17 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.595
+ $Y=1.845 $X2=1.72 $Y2=1.99
r110 1 26 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.72 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_4%A_211_363# 1 2 7 8 9 11 12 16 24 26 28 33
+ 35
c102 9 0 3.37551e-20 $X=2.955 $Y=1.99
c103 8 0 1.85442e-19 $X=2.955 $Y=1.89
r104 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.87
+ $Y=1.52 $X2=2.87 $Y2=1.52
r105 30 32 33.2414 $w=2.9e-07 $l=2e-07 $layer=POLY_cond $X=2.895 $Y=1.32
+ $X2=2.895 $Y2=1.52
r106 27 33 13.5463 $w=2.83e-07 $l=3.35e-07 $layer=LI1_cond $X=2.812 $Y=1.855
+ $X2=2.812 $Y2=1.52
r107 26 28 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.755 $Y=1.855
+ $X2=2.61 $Y2=1.855
r108 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.755 $Y=1.855
+ $X2=2.755 $Y2=1.855
r109 24 28 1.56559 $w=1.4e-07 $l=1.265e-06 $layer=MET1_cond $X=1.345 $Y=1.87
+ $X2=2.61 $Y2=1.87
r110 22 35 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=1.2 $Y=1.855
+ $X2=1.2 $Y2=0.51
r111 21 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.2 $Y=1.855
+ $X2=1.345 $Y2=1.855
r112 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=1.855
+ $X2=1.2 $Y2=1.855
r113 14 16 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.47 $Y=1.245
+ $X2=3.47 $Y2=0.415
r114 13 30 18.1727 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=3.055 $Y=1.32
+ $X2=2.895 $Y2=1.32
r115 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.395 $Y=1.32
+ $X2=3.47 $Y2=1.245
r116 12 13 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.395 $Y=1.32
+ $X2=3.055 $Y2=1.32
r117 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.955 $Y=1.99
+ $X2=2.955 $Y2=2.275
r118 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.955 $Y=1.89 $X2=2.955
+ $Y2=1.99
r119 7 32 32.1081 $w=2.9e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.955 $Y=1.685
+ $X2=2.895 $Y2=1.52
r120 7 8 67.9733 $w=2e-07 $l=2.05e-07 $layer=POLY_cond $X=2.955 $Y=1.685
+ $X2=2.955 $Y2=1.89
r121 2 22 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.815 $X2=1.2 $Y2=1.96
r122 1 35 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_4%A_774_21# 1 2 9 11 13 14 16 17 19 20 22 23
+ 25 26 28 29 31 32 34 35 37 38 45 49 52 55 59 60 69
r119 69 70 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=6.855 $Y=1.202
+ $X2=6.88 $Y2=1.202
r120 68 69 57.9703 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=6.41 $Y=1.202
+ $X2=6.855 $Y2=1.202
r121 67 68 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=6.385 $Y=1.202
+ $X2=6.41 $Y2=1.202
r122 66 67 57.9703 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=5.94 $Y=1.202
+ $X2=6.385 $Y2=1.202
r123 65 66 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.915 $Y=1.202
+ $X2=5.94 $Y2=1.202
r124 64 65 57.9703 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=5.47 $Y=1.202
+ $X2=5.915 $Y2=1.202
r125 63 64 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.445 $Y=1.202
+ $X2=5.47 $Y2=1.202
r126 56 63 5.21081 $w=3.7e-07 $l=4e-08 $layer=POLY_cond $X=5.405 $Y=1.202
+ $X2=5.445 $Y2=1.202
r127 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.405
+ $Y=1.16 $X2=5.405 $Y2=1.16
r128 53 60 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=4.86 $Y=1.16
+ $X2=4.765 $Y2=1.16
r129 53 55 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=4.86 $Y=1.16
+ $X2=5.405 $Y2=1.16
r130 52 59 7.52254 $w=2.05e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.765 $Y=1.535
+ $X2=4.75 $Y2=1.7
r131 51 60 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=4.765 $Y=1.325
+ $X2=4.765 $Y2=1.16
r132 51 52 12.2584 $w=1.88e-07 $l=2.1e-07 $layer=LI1_cond $X=4.765 $Y=1.325
+ $X2=4.765 $Y2=1.535
r133 47 60 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=4.765 $Y=0.995
+ $X2=4.765 $Y2=1.16
r134 47 49 24.2249 $w=1.88e-07 $l=4.15e-07 $layer=LI1_cond $X=4.765 $Y=0.995
+ $X2=4.765 $Y2=0.58
r135 43 59 7.52254 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=4.75 $Y=1.865
+ $X2=4.75 $Y2=1.7
r136 43 45 21.2154 $w=2.18e-07 $l=4.05e-07 $layer=LI1_cond $X=4.75 $Y=1.865
+ $X2=4.75 $Y2=2.27
r137 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.225
+ $Y=1.7 $X2=4.225 $Y2=1.7
r138 38 59 0.30096 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.64 $Y=1.7 $X2=4.75
+ $Y2=1.7
r139 38 40 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=4.64 $Y=1.7
+ $X2=4.225 $Y2=1.7
r140 35 70 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.88 $Y=0.995
+ $X2=6.88 $Y2=1.202
r141 35 37 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.88 $Y=0.995
+ $X2=6.88 $Y2=0.56
r142 32 69 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.855 $Y=1.41
+ $X2=6.855 $Y2=1.202
r143 32 34 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.855 $Y=1.41
+ $X2=6.855 $Y2=1.985
r144 29 68 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.41 $Y=0.995
+ $X2=6.41 $Y2=1.202
r145 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.41 $Y=0.995
+ $X2=6.41 $Y2=0.56
r146 26 67 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.385 $Y=1.41
+ $X2=6.385 $Y2=1.202
r147 26 28 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.385 $Y=1.41
+ $X2=6.385 $Y2=1.985
r148 23 66 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.94 $Y=0.995
+ $X2=5.94 $Y2=1.202
r149 23 25 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.94 $Y=0.995
+ $X2=5.94 $Y2=0.56
r150 20 65 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.915 $Y=1.41
+ $X2=5.915 $Y2=1.202
r151 20 22 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.915 $Y=1.41
+ $X2=5.915 $Y2=1.985
r152 17 64 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.47 $Y=0.995
+ $X2=5.47 $Y2=1.202
r153 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.47 $Y=0.995
+ $X2=5.47 $Y2=0.56
r154 14 63 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.445 $Y=1.41
+ $X2=5.445 $Y2=1.202
r155 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.445 $Y=1.41
+ $X2=5.445 $Y2=1.985
r156 11 41 49.5109 $w=4.1e-07 $l=3.55176e-07 $layer=POLY_cond $X=3.97 $Y=1.99
+ $X2=4.115 $Y2=1.7
r157 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.97 $Y=1.99
+ $X2=3.97 $Y2=2.275
r158 7 41 39.7867 $w=4.1e-07 $l=2.38642e-07 $layer=POLY_cond $X=3.945 $Y=1.535
+ $X2=4.115 $Y2=1.7
r159 7 9 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.945 $Y=1.535
+ $X2=3.945 $Y2=0.445
r160 2 59 600 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=1 $X=4.6
+ $Y=1.485 $X2=4.725 $Y2=1.755
r161 2 45 600 $w=1.7e-07 $l=8.45192e-07 $layer=licon1_PDIFF $count=1 $X=4.6
+ $Y=1.485 $X2=4.725 $Y2=2.27
r162 1 49 182 $w=1.7e-07 $l=4.15331e-07 $layer=licon1_NDIFF $count=1 $X=4.6
+ $Y=0.235 $X2=4.755 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_4%A_609_413# 1 2 7 9 10 12 13 14 15 19 24 26
+ 29 32
c78 32 0 1.69345e-19 $X=3.865 $Y=1.16
c79 14 0 1.24894e-19 $X=4.96 $Y=1.202
c80 13 0 1.83267e-19 $X=4.86 $Y=1.16
r81 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.415
+ $Y=1.16 $X2=4.415 $Y2=1.16
r82 27 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.95 $Y=1.16
+ $X2=3.865 $Y2=1.16
r83 27 29 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.95 $Y=1.16
+ $X2=4.415 $Y2=1.16
r84 25 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.865 $Y=1.325
+ $X2=3.865 $Y2=1.16
r85 25 26 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.865 $Y=1.325
+ $X2=3.865 $Y2=2.255
r86 24 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.865 $Y=0.995
+ $X2=3.865 $Y2=1.16
r87 23 24 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.865 $Y=0.535
+ $X2=3.865 $Y2=0.995
r88 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.78 $Y=0.45
+ $X2=3.865 $Y2=0.535
r89 19 21 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.78 $Y=0.45
+ $X2=3.255 $Y2=0.45
r90 15 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.78 $Y=2.34
+ $X2=3.865 $Y2=2.255
r91 15 17 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.78 $Y=2.34 $X2=3.19
+ $Y2=2.34
r92 13 30 77.8133 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=4.86 $Y=1.16
+ $X2=4.415 $Y2=1.16
r93 13 14 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=4.86 $Y=1.16
+ $X2=4.96 $Y2=1.202
r94 10 14 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=4.985 $Y=0.995
+ $X2=4.96 $Y2=1.202
r95 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.985 $Y=0.995
+ $X2=4.985 $Y2=0.56
r96 7 14 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=4.96 $Y=1.41
+ $X2=4.96 $Y2=1.202
r97 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.96 $Y=1.41 $X2=4.96
+ $Y2=1.985
r98 2 17 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=3.045
+ $Y=2.065 $X2=3.19 $Y2=2.34
r99 1 21 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.235 $X2=3.255 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 39 41 44
+ 45 47 48 49 51 69 73 78 84 87 90 94
c113 25 0 1.85442e-19 $X=2.19 $Y=2
c114 21 0 1.08608e-19 $X=0.73 $Y=2.22
r115 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r116 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r117 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r118 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r119 82 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r120 82 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r121 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r122 79 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.315 $Y=2.72
+ $X2=6.19 $Y2=2.72
r123 79 81 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.315 $Y=2.72
+ $X2=6.67 $Y2=2.72
r124 78 93 3.40825 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=7.005 $Y=2.72
+ $X2=7.182 $Y2=2.72
r125 78 81 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.005 $Y=2.72
+ $X2=6.67 $Y2=2.72
r126 77 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r127 77 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r128 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r129 74 87 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.375 $Y=2.72
+ $X2=5.232 $Y2=2.72
r130 74 76 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.375 $Y=2.72
+ $X2=5.75 $Y2=2.72
r131 73 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.065 $Y=2.72
+ $X2=6.19 $Y2=2.72
r132 73 76 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.065 $Y=2.72
+ $X2=5.75 $Y2=2.72
r133 72 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r134 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r135 69 87 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=5.09 $Y=2.72
+ $X2=5.232 $Y2=2.72
r136 69 71 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.09 $Y=2.72
+ $X2=4.83 $Y2=2.72
r137 68 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r138 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r139 65 68 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r140 64 67 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r141 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r142 62 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r143 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r144 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r145 59 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r146 58 61 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r147 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r148 56 84 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r149 56 58 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r150 51 84 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r151 51 53 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r152 49 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r153 49 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r154 47 67 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.12 $Y=2.72
+ $X2=3.91 $Y2=2.72
r155 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.12 $Y=2.72
+ $X2=4.205 $Y2=2.72
r156 46 71 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r157 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.29 $Y=2.72
+ $X2=4.205 $Y2=2.72
r158 44 61 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.07 $Y2=2.72
r159 44 45 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.262 $Y2=2.72
r160 43 64 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.42 $Y=2.72
+ $X2=2.53 $Y2=2.72
r161 43 45 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.42 $Y=2.72
+ $X2=2.262 $Y2=2.72
r162 39 93 3.40825 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=7.09 $Y=2.635
+ $X2=7.182 $Y2=2.72
r163 39 41 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=7.09 $Y=2.635
+ $X2=7.09 $Y2=1.835
r164 35 90 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.19 $Y=2.635
+ $X2=6.19 $Y2=2.72
r165 35 37 36.8782 $w=2.48e-07 $l=8e-07 $layer=LI1_cond $X=6.19 $Y=2.635
+ $X2=6.19 $Y2=1.835
r166 31 87 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=5.232 $Y=2.635
+ $X2=5.232 $Y2=2.72
r167 31 33 36.3929 $w=2.83e-07 $l=9e-07 $layer=LI1_cond $X=5.232 $Y=2.635
+ $X2=5.232 $Y2=1.735
r168 27 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.205 $Y=2.635
+ $X2=4.205 $Y2=2.72
r169 27 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.205 $Y=2.635
+ $X2=4.205 $Y2=2.3
r170 23 45 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.262 $Y=2.635
+ $X2=2.262 $Y2=2.72
r171 23 25 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=2.262 $Y=2.635
+ $X2=2.262 $Y2=2
r172 19 84 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r173 19 21 12.5859 $w=3.78e-07 $l=4.15e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.22
r174 6 41 300 $w=1.7e-07 $l=4.16233e-07 $layer=licon1_PDIFF $count=2 $X=6.945
+ $Y=1.485 $X2=7.09 $Y2=1.835
r175 5 37 300 $w=1.7e-07 $l=4.16233e-07 $layer=licon1_PDIFF $count=2 $X=6.005
+ $Y=1.485 $X2=6.15 $Y2=1.835
r176 4 33 300 $w=1.7e-07 $l=3.20156e-07 $layer=licon1_PDIFF $count=2 $X=5.05
+ $Y=1.485 $X2=5.21 $Y2=1.735
r177 3 29 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=4.06
+ $Y=2.065 $X2=4.205 $Y2=2.3
r178 2 25 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=1.845 $X2=2.19 $Y2=2
r179 1 21 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.815 $X2=0.73 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_4%Q 1 2 3 4 14 17 18 20 21 22 23 24 25 26 27
+ 28 29 30 47 50 68
c50 20 0 1.24894e-19 $X=5.802 $Y=1.16
r51 47 50 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=6.535 $Y=1.16
+ $X2=6.245 $Y2=1.16
r52 30 68 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=7.12 $Y=1.16
+ $X2=7.125 $Y2=1.16
r53 30 65 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=7.12 $Y=1.16
+ $X2=6.805 $Y2=1.16
r54 29 51 7.45556 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.67 $Y=1.16
+ $X2=6.67 $Y2=0.995
r55 29 58 7.45556 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.67 $Y=1.16
+ $X2=6.67 $Y2=1.325
r56 29 47 4.99091 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=6.67 $Y=1.16
+ $X2=6.535 $Y2=1.16
r57 29 65 4.99091 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=6.67 $Y=1.16
+ $X2=6.805 $Y2=1.16
r58 27 28 16.0062 $w=2.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.67 $Y=1.835
+ $X2=6.67 $Y2=2.21
r59 27 58 21.7684 $w=2.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.67 $Y=1.835
+ $X2=6.67 $Y2=1.325
r60 26 51 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.67 $Y=0.85
+ $X2=6.67 $Y2=0.995
r61 25 26 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.67 $Y=0.51
+ $X2=6.67 $Y2=0.85
r62 24 50 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.23 $Y=1.16
+ $X2=6.245 $Y2=1.16
r63 22 23 14.4055 $w=2.98e-07 $l=3.75e-07 $layer=LI1_cond $X=5.745 $Y=1.835
+ $X2=5.745 $Y2=2.21
r64 21 74 10.7101 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=5.745 $Y=0.51
+ $X2=5.745 $Y2=0.745
r65 19 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.895 $Y=1.16
+ $X2=6.23 $Y2=1.16
r66 19 20 0.63164 $w=3.3e-07 $l=9.3e-08 $layer=LI1_cond $X=5.895 $Y=1.16
+ $X2=5.802 $Y2=1.16
r67 17 22 7.29881 $w=2.98e-07 $l=1.9e-07 $layer=LI1_cond $X=5.745 $Y=1.645
+ $X2=5.745 $Y2=1.835
r68 17 18 7.4448 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=5.745 $Y=1.645
+ $X2=5.745 $Y2=1.495
r69 15 20 8.10876 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=5.802 $Y=1.325
+ $X2=5.802 $Y2=1.16
r70 15 18 10.1916 $w=1.83e-07 $l=1.7e-07 $layer=LI1_cond $X=5.802 $Y=1.325
+ $X2=5.802 $Y2=1.495
r71 14 20 8.10876 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=5.802 $Y=0.995
+ $X2=5.802 $Y2=1.16
r72 14 74 14.9877 $w=1.83e-07 $l=2.5e-07 $layer=LI1_cond $X=5.802 $Y=0.995
+ $X2=5.802 $Y2=0.745
r73 4 27 300 $w=1.7e-07 $l=4.16233e-07 $layer=licon1_PDIFF $count=2 $X=6.475
+ $Y=1.485 $X2=6.62 $Y2=1.835
r74 3 22 300 $w=1.7e-07 $l=4.16233e-07 $layer=licon1_PDIFF $count=2 $X=5.535
+ $Y=1.485 $X2=5.68 $Y2=1.835
r75 2 25 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=6.485
+ $Y=0.235 $X2=6.62 $Y2=0.55
r76 1 21 182 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_NDIFF $count=1 $X=5.545
+ $Y=0.235 $X2=5.68 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_4%VGND 1 2 3 4 5 6 21 25 29 31 33 36 37 38
+ 40 45 57 61 66 73 80 86 89 93
c106 93 0 2.71124e-20 $X=7.13 $Y=0
c107 21 0 1.83267e-19 $X=4.205 $Y=0.445
c108 2 0 7.13094e-20 $X=2.055 $Y=0.235
r109 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r110 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r111 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r112 80 83 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=2.165 $Y=0
+ $X2=2.165 $Y2=0.36
r113 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r114 73 76 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.38
r115 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r116 70 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r117 70 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r118 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r119 67 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.315 $Y=0 $X2=6.19
+ $Y2=0
r120 67 69 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.315 $Y=0
+ $X2=6.67 $Y2=0
r121 66 92 3.40825 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=7.005 $Y=0
+ $X2=7.182 $Y2=0
r122 66 69 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.005 $Y=0
+ $X2=6.67 $Y2=0
r123 65 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r124 65 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=5.29
+ $Y2=0
r125 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r126 62 86 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.375 $Y=0
+ $X2=5.232 $Y2=0
r127 62 64 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.375 $Y=0
+ $X2=5.75 $Y2=0
r128 61 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.065 $Y=0 $X2=6.19
+ $Y2=0
r129 61 64 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.065 $Y=0
+ $X2=5.75 $Y2=0
r130 60 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r131 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r132 57 86 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=5.09 $Y=0 $X2=5.232
+ $Y2=0
r133 57 59 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.09 $Y=0 $X2=4.83
+ $Y2=0
r134 56 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r135 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r136 53 56 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.91 $Y2=0
r137 53 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r138 52 55 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r139 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r140 50 80 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.165
+ $Y2=0
r141 50 52 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.355 $Y=0
+ $X2=2.53 $Y2=0
r142 49 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r143 49 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r144 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r145 46 73 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r146 46 48 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.61 $Y2=0
r147 45 80 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=2.165
+ $Y2=0
r148 45 48 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.975 $Y=0
+ $X2=1.61 $Y2=0
r149 40 73 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r150 40 42 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r151 38 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r152 38 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r153 36 55 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.12 $Y=0 $X2=3.91
+ $Y2=0
r154 36 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.12 $Y=0 $X2=4.205
+ $Y2=0
r155 35 59 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.29 $Y=0 $X2=4.83
+ $Y2=0
r156 35 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.29 $Y=0 $X2=4.205
+ $Y2=0
r157 31 92 3.40825 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=7.09 $Y=0.085
+ $X2=7.182 $Y2=0
r158 31 33 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=7.09 $Y=0.085
+ $X2=7.09 $Y2=0.55
r159 27 89 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.19 $Y=0.085
+ $X2=6.19 $Y2=0
r160 27 29 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=6.19 $Y=0.085
+ $X2=6.19 $Y2=0.55
r161 23 86 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=5.232 $Y=0.085
+ $X2=5.232 $Y2=0
r162 23 25 18.803 $w=2.83e-07 $l=4.65e-07 $layer=LI1_cond $X=5.232 $Y=0.085
+ $X2=5.232 $Y2=0.55
r163 19 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.205 $Y=0.085
+ $X2=4.205 $Y2=0
r164 19 21 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.205 $Y=0.085
+ $X2=4.205 $Y2=0.445
r165 6 33 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=6.955
+ $Y=0.235 $X2=7.09 $Y2=0.55
r166 5 29 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=6.015
+ $Y=0.235 $X2=6.15 $Y2=0.55
r167 4 25 182 $w=1.7e-07 $l=3.82721e-07 $layer=licon1_NDIFF $count=1 $X=5.06
+ $Y=0.235 $X2=5.21 $Y2=0.55
r168 3 21 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=4.02
+ $Y=0.235 $X2=4.205 $Y2=0.445
r169 2 83 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.055
+ $Y=0.235 $X2=2.19 $Y2=0.36
r170 1 76 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

