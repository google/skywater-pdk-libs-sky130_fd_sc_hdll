* File: sky130_fd_sc_hdll__dfrtp_1.pex.spice
* Created: Wed Sep  2 08:28:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__DFRTP_1%CLK 1 2 3 5 6 8 13 14
c37 3 0 9.59708e-20 $X=0.495 $Y=1.74
c38 1 0 2.71124e-20 $X=0.305 $Y=1.325
r39 13 14 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.265 $Y=1.16
+ $X2=0.265 $Y2=1.53
r40 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r41 6 18 86.21 $w=2.7e-07 $l=5.0709e-07 $layer=POLY_cond $X=0.52 $Y=0.73
+ $X2=0.352 $Y2=1.16
r42 6 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.445
r43 3 9 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.495 $Y=1.665
+ $X2=0.305 $Y2=1.665
r44 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.74
+ $X2=0.495 $Y2=2.135
r45 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r46 1 18 38.9026 $w=2.7e-07 $l=1.87029e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.352 $Y2=1.16
r47 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.305 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_1%A_27_47# 1 2 8 9 11 14 17 20 22 23 25 26
+ 28 30 31 33 36 40 41 45 49 50 51 54 57 58 59 60 63 69 73 74 80 83 84
c239 84 0 5.71407e-20 $X=2.535 $Y=0.93
c240 74 0 1.3501e-20 $X=6.17 $Y=1.11
c241 60 0 7.20353e-20 $X=2.71 $Y=1.19
c242 59 0 1.58851e-19 $X=5.96 $Y=1.19
c243 40 0 1.21524e-19 $X=6.112 $Y=1.395
c244 30 0 6.96392e-20 $X=6.02 $Y=1.89
c245 26 0 1.56398e-19 $X=3.155 $Y=1.99
c246 23 0 2.20662e-19 $X=2.67 $Y=1.32
r247 83 86 40.2795 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.535 $Y=0.93
+ $X2=2.535 $Y2=1.095
r248 83 85 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.535 $Y=0.93
+ $X2=2.535 $Y2=0.765
r249 83 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.535
+ $Y=0.93 $X2=2.535 $Y2=0.93
r250 79 80 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.235
+ $X2=0.99 $Y2=1.235
r251 76 79 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=0.805 $Y=1.235
+ $X2=0.965 $Y2=1.235
r252 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.17
+ $Y=1.11 $X2=6.17 $Y2=1.11
r253 69 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.105 $Y=1.19
+ $X2=6.105 $Y2=1.19
r254 67 84 11.5244 $w=2.58e-07 $l=2.6e-07 $layer=LI1_cond $X=2.555 $Y=1.19
+ $X2=2.555 $Y2=0.93
r255 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.565 $Y=1.19
+ $X2=2.565 $Y2=1.19
r256 63 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.805
+ $Y=1.235 $X2=0.805 $Y2=1.235
r257 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.745 $Y=1.19
+ $X2=0.745 $Y2=1.19
r258 60 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.71 $Y=1.19
+ $X2=2.565 $Y2=1.19
r259 59 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.96 $Y=1.19
+ $X2=6.105 $Y2=1.19
r260 59 60 4.02227 $w=1.4e-07 $l=3.25e-06 $layer=MET1_cond $X=5.96 $Y=1.19
+ $X2=2.71 $Y2=1.19
r261 58 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.89 $Y=1.19
+ $X2=0.745 $Y2=1.19
r262 57 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.42 $Y=1.19
+ $X2=2.565 $Y2=1.19
r263 57 58 1.89356 $w=1.4e-07 $l=1.53e-06 $layer=MET1_cond $X=2.42 $Y=1.19
+ $X2=0.89 $Y2=1.19
r264 56 63 30.3143 $w=2.28e-07 $l=6.05e-07 $layer=LI1_cond $X=0.775 $Y=1.795
+ $X2=0.775 $Y2=1.19
r265 55 63 19.2909 $w=2.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.775 $Y=0.805
+ $X2=0.775 $Y2=1.19
r266 52 54 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.217 $Y2=1.88
r267 51 56 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.66 $Y=1.88
+ $X2=0.775 $Y2=1.795
r268 51 52 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.66 $Y=1.88
+ $X2=0.345 $Y2=1.88
r269 49 55 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.66 $Y=0.72
+ $X2=0.775 $Y2=0.805
r270 49 50 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.66 $Y=0.72
+ $X2=0.345 $Y2=0.72
r271 43 50 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.217 $Y=0.635
+ $X2=0.345 $Y2=0.72
r272 43 45 5.64923 $w=2.53e-07 $l=1.25e-07 $layer=LI1_cond $X=0.217 $Y=0.635
+ $X2=0.217 $Y2=0.51
r273 41 73 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=6.17 $Y=1.08 $X2=6.17
+ $Y2=1.11
r274 41 42 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=6.17 $Y=1.08
+ $X2=6.17 $Y2=0.945
r275 39 73 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=6.17 $Y=1.245
+ $X2=6.17 $Y2=1.11
r276 39 40 37.4821 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=6.112 $Y=1.245
+ $X2=6.112 $Y2=1.395
r277 36 42 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.11 $Y=0.415
+ $X2=6.11 $Y2=0.945
r278 31 33 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.02 $Y=1.99
+ $X2=6.02 $Y2=2.275
r279 30 31 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=6.02 $Y=1.89 $X2=6.02
+ $Y2=1.99
r280 30 40 164.131 $w=2e-07 $l=4.95e-07 $layer=POLY_cond $X=6.02 $Y=1.89
+ $X2=6.02 $Y2=1.395
r281 26 28 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.155 $Y=1.99
+ $X2=3.155 $Y2=2.275
r282 25 26 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.155 $Y=1.89 $X2=3.155
+ $Y2=1.99
r283 24 25 164.131 $w=2e-07 $l=4.95e-07 $layer=POLY_cond $X=3.155 $Y=1.395
+ $X2=3.155 $Y2=1.89
r284 22 24 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=3.055 $Y=1.32
+ $X2=3.155 $Y2=1.395
r285 22 23 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=3.055 $Y=1.32
+ $X2=2.67 $Y2=1.32
r286 20 85 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.595 $Y=0.415
+ $X2=2.595 $Y2=0.765
r287 17 23 27.7801 $w=1.5e-07 $l=1.35403e-07 $layer=POLY_cond $X=2.567 $Y=1.245
+ $X2=2.67 $Y2=1.32
r288 17 86 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=2.567 $Y=1.245
+ $X2=2.567 $Y2=1.095
r289 12 80 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=1.235
r290 12 14 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=0.445
r291 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.965 $Y=1.74
+ $X2=0.965 $Y2=2.135
r292 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.64 $X2=0.965
+ $Y2=1.74
r293 7 79 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=0.965 $Y=1.37
+ $X2=0.965 $Y2=1.235
r294 7 8 89.5258 $w=2e-07 $l=2.7e-07 $layer=POLY_cond $X=0.965 $Y=1.37 $X2=0.965
+ $Y2=1.64
r295 2 54 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r296 1 45 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_1%D 2 3 5 8 14 18 21
c51 2 0 1.2021e-19 $X=2.09 $Y=1.89
r52 20 21 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.09 $Y=1.465
+ $X2=2.115 $Y2=1.465
r53 17 20 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=1.82 $Y=1.465
+ $X2=2.09 $Y2=1.465
r54 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.82
+ $Y=1.465 $X2=1.82 $Y2=1.465
r55 14 18 1.72767 $w=4.48e-07 $l=6.5e-08 $layer=LI1_cond $X=1.68 $Y=1.53
+ $X2=1.68 $Y2=1.465
r56 6 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.115 $Y=1.3
+ $X2=2.115 $Y2=1.465
r57 6 8 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=2.115 $Y=1.3
+ $X2=2.115 $Y2=0.445
r58 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.09 $Y=1.99 $X2=2.09
+ $Y2=2.275
r59 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.09 $Y=1.89 $X2=2.09
+ $Y2=1.99
r60 1 20 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.09 $Y=1.63 $X2=2.09
+ $Y2=1.465
r61 1 2 86.2101 $w=2e-07 $l=2.6e-07 $layer=POLY_cond $X=2.09 $Y=1.63 $X2=2.09
+ $Y2=1.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_1%A_211_363# 1 2 7 9 12 14 16 17 19 21 24 25
+ 27 28 32 35 36 37 38 47 55 63 65 73
c215 73 0 1.2021e-19 $X=2.94 $Y=1.77
c216 63 0 2.86831e-20 $X=6.495 $Y=1.74
c217 55 0 8.91419e-20 $X=3.135 $Y=0.9
c218 38 0 5.71407e-20 $X=2.955 $Y=1.87
c219 36 0 9.59708e-20 $X=1.345 $Y=1.87
c220 35 0 1.17518e-19 $X=2.665 $Y=1.87
c221 24 0 1.38067e-19 $X=5.69 $Y=0.87
c222 17 0 5.51005e-20 $X=6.56 $Y=1.99
r223 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.495
+ $Y=1.74 $X2=6.495 $Y2=1.74
r224 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.595
+ $Y=1.74 $X2=2.595 $Y2=1.74
r225 47 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.555 $Y=1.87
+ $X2=6.555 $Y2=1.87
r226 45 73 3.84148 $w=3.88e-07 $l=1.3e-07 $layer=LI1_cond $X=2.81 $Y=1.77
+ $X2=2.94 $Y2=1.77
r227 45 52 6.35321 $w=3.88e-07 $l=2.15e-07 $layer=LI1_cond $X=2.81 $Y=1.77
+ $X2=2.595 $Y2=1.77
r228 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.81 $Y=1.87
+ $X2=2.81 $Y2=1.87
r229 41 65 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.2 $Y=1.87
+ $X2=1.2 $Y2=0.51
r230 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=1.87 $X2=1.2
+ $Y2=1.87
r231 38 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.955 $Y=1.87
+ $X2=2.81 $Y2=1.87
r232 37 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.41 $Y=1.87
+ $X2=6.555 $Y2=1.87
r233 37 38 4.27598 $w=1.4e-07 $l=3.455e-06 $layer=MET1_cond $X=6.41 $Y=1.87
+ $X2=2.955 $Y2=1.87
r234 36 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=1.87
+ $X2=1.2 $Y2=1.87
r235 35 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.665 $Y=1.87
+ $X2=2.81 $Y2=1.87
r236 35 36 1.63366 $w=1.4e-07 $l=1.32e-06 $layer=MET1_cond $X=2.665 $Y=1.87
+ $X2=1.345 $Y2=1.87
r237 33 55 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=3.045 $Y=0.9
+ $X2=3.135 $Y2=0.9
r238 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.045
+ $Y=0.9 $X2=3.045 $Y2=0.9
r239 29 32 5.5003 $w=2.18e-07 $l=1.05e-07 $layer=LI1_cond $X=2.94 $Y=0.875
+ $X2=3.045 $Y2=0.875
r240 27 63 15.4023 $w=3.52e-07 $l=4.16233e-07 $layer=LI1_cond $X=6.145 $Y=1.58
+ $X2=6.495 $Y2=1.725
r241 27 28 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.145 $Y=1.58
+ $X2=5.775 $Y2=1.58
r242 25 57 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.69 $Y=0.87
+ $X2=5.565 $Y2=0.87
r243 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.69
+ $Y=0.87 $X2=5.69 $Y2=0.87
r244 22 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.69 $Y=1.495
+ $X2=5.775 $Y2=1.58
r245 22 24 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=5.69 $Y=1.495
+ $X2=5.69 $Y2=0.87
r246 21 73 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.94 $Y=1.575
+ $X2=2.94 $Y2=1.77
r247 20 29 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.94 $Y=0.985
+ $X2=2.94 $Y2=0.875
r248 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.94 $Y=0.985
+ $X2=2.94 $Y2=1.575
r249 17 62 47.761 $w=3.01e-07 $l=2.80624e-07 $layer=POLY_cond $X=6.56 $Y=1.99
+ $X2=6.495 $Y2=1.74
r250 17 19 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.56 $Y=1.99
+ $X2=6.56 $Y2=2.275
r251 14 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.565 $Y=0.705
+ $X2=5.565 $Y2=0.87
r252 14 16 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.565 $Y=0.705
+ $X2=5.565 $Y2=0.415
r253 10 55 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.135 $Y=0.765
+ $X2=3.135 $Y2=0.9
r254 10 12 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.135 $Y=0.765
+ $X2=3.135 $Y2=0.415
r255 7 51 46.5577 $w=3.26e-07 $l=2.54951e-07 $layer=POLY_cond $X=2.61 $Y=1.99
+ $X2=2.62 $Y2=1.74
r256 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.61 $Y=1.99
+ $X2=2.61 $Y2=2.275
r257 2 41 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.815 $X2=1.2 $Y2=1.96
r258 1 65 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_1%A_751_289# 1 2 7 9 12 14 20 22 24 25 26 29
+ 34 36 37
c111 37 0 2.78699e-20 $X=5.24 $Y=1.61
c112 36 0 2.40285e-19 $X=5.195 $Y=0.835
c113 26 0 6.86107e-20 $X=5.325 $Y=1.92
c114 22 0 4.17692e-20 $X=5.24 $Y=1.525
r115 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.73 $Y=2.005
+ $X2=5.73 $Y2=2.3
r116 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.645 $Y=1.92
+ $X2=5.73 $Y2=2.005
r117 25 26 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.645 $Y=1.92
+ $X2=5.325 $Y2=1.92
r118 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.24 $Y=1.835
+ $X2=5.325 $Y2=1.92
r119 23 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.24 $Y=1.695
+ $X2=5.24 $Y2=1.61
r120 23 24 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.24 $Y=1.695
+ $X2=5.24 $Y2=1.835
r121 22 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.24 $Y=1.525
+ $X2=5.24 $Y2=1.61
r122 22 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.24 $Y=1.525
+ $X2=5.24 $Y2=0.835
r123 20 36 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=5.195 $Y=0.705
+ $X2=5.195 $Y2=0.835
r124 19 34 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=5.195 $Y=0.36
+ $X2=5.3 $Y2=0.36
r125 19 20 11.5244 $w=2.58e-07 $l=2.6e-07 $layer=LI1_cond $X=5.195 $Y=0.445
+ $X2=5.195 $Y2=0.705
r126 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.89
+ $Y=1.61 $X2=3.89 $Y2=1.61
r127 14 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=1.61
+ $X2=5.24 $Y2=1.61
r128 14 16 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=5.155 $Y=1.61
+ $X2=3.89 $Y2=1.61
r129 10 17 38.8084 $w=2.75e-07 $l=1.80748e-07 $layer=POLY_cond $X=3.95 $Y=1.445
+ $X2=3.917 $Y2=1.61
r130 10 12 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=3.95 $Y=1.445
+ $X2=3.95 $Y2=0.445
r131 7 17 72.3531 $w=2.75e-07 $l=4.09829e-07 $layer=POLY_cond $X=3.855 $Y=1.99
+ $X2=3.917 $Y2=1.61
r132 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.855 $Y=1.99
+ $X2=3.855 $Y2=2.275
r133 2 29 600 $w=1.7e-07 $l=7.32871e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=1.645 $X2=5.73 $Y2=2.3
r134 1 34 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=5.145
+ $Y=0.235 $X2=5.3 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_1%RESET_B 3 5 6 8 11 14 15 17 18 21 23 24 25
+ 28 30 33 42
c141 28 0 1.04922e-19 $X=4.37 $Y=0.93
c142 23 0 1.21524e-19 $X=7.575 $Y=0.85
c143 21 0 6.89774e-20 $X=4.55 $Y=0.85
c144 15 0 1.5899e-19 $X=7.66 $Y=1.99
c145 6 0 6.86107e-20 $X=4.39 $Y=1.99
r146 34 42 7.77899 $w=3.98e-07 $l=2.7e-07 $layer=LI1_cond $X=7.705 $Y=1.12
+ $X2=7.705 $Y2=0.85
r147 33 36 40.3353 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.7 $Y=1.12
+ $X2=7.7 $Y2=1.285
r148 33 35 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.7 $Y=1.12
+ $X2=7.7 $Y2=0.955
r149 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.695
+ $Y=1.12 $X2=7.695 $Y2=1.12
r150 28 31 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.395 $Y=0.93
+ $X2=4.395 $Y2=1.095
r151 28 30 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.395 $Y=0.93
+ $X2=4.395 $Y2=0.765
r152 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.37
+ $Y=0.93 $X2=4.37 $Y2=0.93
r153 25 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.72 $Y=0.85
+ $X2=7.72 $Y2=0.85
r154 23 25 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.575 $Y=0.85
+ $X2=7.72 $Y2=0.85
r155 23 24 3.50247 $w=1.4e-07 $l=2.83e-06 $layer=MET1_cond $X=7.575 $Y=0.85
+ $X2=4.745 $Y2=0.85
r156 21 29 1.13912 $w=8.38e-07 $l=8e-08 $layer=LI1_cond $X=4.225 $Y=0.85
+ $X2=4.225 $Y2=0.93
r157 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.55 $Y=0.85
+ $X2=4.55 $Y2=0.85
r158 18 24 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=4.63 $Y=0.85
+ $X2=4.745 $Y2=0.85
r159 18 20 0.0513283 $w=2.3e-07 $l=8e-08 $layer=MET1_cond $X=4.63 $Y=0.85
+ $X2=4.55 $Y2=0.85
r160 15 17 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.66 $Y=1.99
+ $X2=7.66 $Y2=2.275
r161 14 15 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.66 $Y=1.89 $X2=7.66
+ $Y2=1.99
r162 14 36 200.604 $w=2e-07 $l=6.05e-07 $layer=POLY_cond $X=7.66 $Y=1.89
+ $X2=7.66 $Y2=1.285
r163 11 35 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=7.635 $Y=0.445
+ $X2=7.635 $Y2=0.955
r164 6 8 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=4.39 $Y=1.99
+ $X2=4.39 $Y2=2.275
r165 5 6 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.39 $Y=1.89 $X2=4.39
+ $Y2=1.99
r166 5 31 263.604 $w=2e-07 $l=7.95e-07 $layer=POLY_cond $X=4.39 $Y=1.89 $X2=4.39
+ $Y2=1.095
r167 3 30 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.31 $Y=0.445
+ $X2=4.31 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_1%A_534_47# 1 2 9 11 13 15 16 20 25 27 28 29
+ 34 35
c128 35 0 6.89774e-20 $X=4.9 $Y=1.17
c129 29 0 8.91419e-20 $X=3.6 $Y=1.27
c130 11 0 1.35364e-19 $X=5.385 $Y=1.495
c131 9 0 1.38067e-19 $X=5.07 $Y=0.555
r132 35 40 51.3607 $w=3.05e-07 $l=3.25e-07 $layer=POLY_cond $X=4.955 $Y=1.17
+ $X2=4.955 $Y2=1.495
r133 34 37 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.9 $Y=1.17 $X2=4.9
+ $Y2=1.27
r134 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.9
+ $Y=1.17 $X2=4.9 $Y2=1.17
r135 30 32 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.28 $Y=1.27
+ $X2=3.515 $Y2=1.27
r136 29 32 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=1.27
+ $X2=3.515 $Y2=1.27
r137 28 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.815 $Y=1.27
+ $X2=4.9 $Y2=1.27
r138 28 29 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=4.815 $Y=1.27
+ $X2=3.6 $Y2=1.27
r139 27 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=1.185
+ $X2=3.515 $Y2=1.27
r140 26 27 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.515 $Y=0.475
+ $X2=3.515 $Y2=1.185
r141 24 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.28 $Y=1.355
+ $X2=3.28 $Y2=1.27
r142 24 25 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.28 $Y=1.355
+ $X2=3.28 $Y2=2.135
r143 20 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.43 $Y=0.39
+ $X2=3.515 $Y2=0.475
r144 20 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.43 $Y=0.39
+ $X2=2.86 $Y2=0.39
r145 16 25 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.195 $Y=2.3
+ $X2=3.28 $Y2=2.135
r146 16 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.195 $Y=2.3
+ $X2=2.85 $Y2=2.3
r147 13 15 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=5.475 $Y=1.57
+ $X2=5.475 $Y2=2.065
r148 12 40 19.3576 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.145 $Y=1.495
+ $X2=4.955 $Y2=1.495
r149 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.385 $Y=1.495
+ $X2=5.475 $Y2=1.57
r150 11 12 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=5.385 $Y=1.495
+ $X2=5.145 $Y2=1.495
r151 7 35 38.5368 $w=3.05e-07 $l=2.14942e-07 $layer=POLY_cond $X=5.07 $Y=1.005
+ $X2=4.955 $Y2=1.17
r152 7 9 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=5.07 $Y=1.005
+ $X2=5.07 $Y2=0.555
r153 2 18 600 $w=1.7e-07 $l=3.31625e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=2.065 $X2=2.85 $Y2=2.33
r154 1 22 182 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_NDIFF $count=1 $X=2.67
+ $Y=0.235 $X2=2.86 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_1%A_1323_21# 1 2 9 12 13 15 16 18 19 21 24
+ 29 30 33 35 36 37 38 40 43 46 47 50 52
c134 52 0 2.86831e-20 $X=6.97 $Y=0.98
c135 12 0 1.3501e-20 $X=6.97 $Y=1.89
r136 46 47 8.82932 $w=2.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.145 $Y=0.695
+ $X2=7.145 $Y2=0.865
r137 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.905
+ $Y=1.16 $X2=8.905 $Y2=1.16
r138 41 50 2.08613 $w=2.1e-07 $l=3.94018e-07 $layer=LI1_cond $X=8.635 $Y=1.18
+ $X2=8.29 $Y2=1.075
r139 41 43 14.2597 $w=2.08e-07 $l=2.7e-07 $layer=LI1_cond $X=8.635 $Y=1.18
+ $X2=8.905 $Y2=1.18
r140 39 50 4.34585 $w=2.57e-07 $l=3.26994e-07 $layer=LI1_cond $X=8.525 $Y=1.295
+ $X2=8.29 $Y2=1.075
r141 39 40 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=8.525 $Y=1.295
+ $X2=8.525 $Y2=1.915
r142 38 50 4.34585 $w=2.57e-07 $l=1.72e-07 $layer=LI1_cond $X=8.462 $Y=1.075
+ $X2=8.29 $Y2=1.075
r143 37 49 2.61083 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=8.462 $Y=0.465
+ $X2=8.462 $Y2=0.38
r144 37 38 20.3765 $w=3.43e-07 $l=6.1e-07 $layer=LI1_cond $X=8.462 $Y=0.465
+ $X2=8.462 $Y2=1.075
r145 35 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.44 $Y=2
+ $X2=8.525 $Y2=1.915
r146 35 36 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=8.44 $Y=2 $X2=7.98
+ $Y2=2
r147 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.895 $Y=2.085
+ $X2=7.98 $Y2=2
r148 31 33 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.895 $Y=2.085
+ $X2=7.895 $Y2=2.21
r149 29 49 5.28309 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=8.29 $Y=0.38
+ $X2=8.462 $Y2=0.38
r150 29 30 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=8.29 $Y=0.38
+ $X2=7.335 $Y2=0.38
r151 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.25 $Y=0.465
+ $X2=7.335 $Y2=0.38
r152 27 46 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.25 $Y=0.465
+ $X2=7.25 $Y2=0.695
r153 25 52 13.2835 $w=2.54e-07 $l=7e-08 $layer=POLY_cond $X=7.04 $Y=0.98
+ $X2=6.97 $Y2=0.98
r154 24 47 4.90855 $w=2.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.09 $Y=0.98
+ $X2=7.09 $Y2=0.865
r155 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.04
+ $Y=0.98 $X2=7.04 $Y2=0.98
r156 19 44 39.7049 $w=4.06e-07 $l=2.29783e-07 $layer=POLY_cond $X=9.155 $Y=0.995
+ $X2=9 $Y2=1.16
r157 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.155 $Y=0.995
+ $X2=9.155 $Y2=0.56
r158 16 44 44.8379 $w=4.06e-07 $l=3.08221e-07 $layer=POLY_cond $X=9.13 $Y=1.41
+ $X2=9 $Y2=1.16
r159 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.13 $Y=1.41
+ $X2=9.13 $Y2=1.985
r160 13 15 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.97 $Y=1.99
+ $X2=6.97 $Y2=2.275
r161 12 13 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=6.97 $Y=1.89 $X2=6.97
+ $Y2=1.99
r162 11 52 8.45288 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=6.97 $Y=1.145
+ $X2=6.97 $Y2=0.98
r163 11 12 247.025 $w=2e-07 $l=7.45e-07 $layer=POLY_cond $X=6.97 $Y=1.145
+ $X2=6.97 $Y2=1.89
r164 7 52 53.1339 $w=2.54e-07 $l=3.52987e-07 $layer=POLY_cond $X=6.69 $Y=0.815
+ $X2=6.97 $Y2=0.98
r165 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.69 $Y=0.815
+ $X2=6.69 $Y2=0.445
r166 2 33 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.75
+ $Y=2.065 $X2=7.895 $Y2=2.21
r167 1 49 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=8.24
+ $Y=0.235 $X2=8.375 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_1%A_1128_47# 1 2 7 9 12 14 18 23 24 25 27 30
+ 33
c105 24 0 5.51005e-20 $X=6.835 $Y=1.4
c106 23 0 1.99514e-19 $X=6.57 $Y=1.315
c107 18 0 1.5899e-19 $X=6.835 $Y=2.295
r108 35 36 5.0779 $w=2.18e-07 $l=8.5e-08 $layer=LI1_cond $X=6.945 $Y=1.66
+ $X2=6.945 $Y2=1.745
r109 33 35 13.6198 $w=2.18e-07 $l=2.6e-07 $layer=LI1_cond $X=6.945 $Y=1.4
+ $X2=6.945 $Y2=1.66
r110 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.105
+ $Y=1.66 $X2=8.105 $Y2=1.66
r111 28 35 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=7.055 $Y=1.66
+ $X2=6.945 $Y2=1.66
r112 28 30 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=7.055 $Y=1.66
+ $X2=8.105 $Y2=1.66
r113 27 36 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.92 $Y=2.125
+ $X2=6.92 $Y2=1.745
r114 24 33 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=6.835 $Y=1.4
+ $X2=6.945 $Y2=1.4
r115 24 25 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.835 $Y=1.4
+ $X2=6.655 $Y2=1.4
r116 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.57 $Y=1.315
+ $X2=6.655 $Y2=1.4
r117 22 23 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=6.57 $Y=0.535
+ $X2=6.57 $Y2=1.315
r118 18 27 7.85115 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=6.835 $Y=2.295
+ $X2=6.92 $Y2=2.125
r119 18 20 19.3204 $w=3.38e-07 $l=5.7e-07 $layer=LI1_cond $X=6.835 $Y=2.295
+ $X2=6.265 $Y2=2.295
r120 14 22 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.485 $Y=0.395
+ $X2=6.57 $Y2=0.535
r121 14 16 24.0778 $w=2.78e-07 $l=5.85e-07 $layer=LI1_cond $X=6.485 $Y=0.395
+ $X2=5.9 $Y2=0.395
r122 10 31 39.6178 $w=2.46e-07 $l=1.92678e-07 $layer=POLY_cond $X=8.165 $Y=1.495
+ $X2=8.105 $Y2=1.66
r123 10 12 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=8.165 $Y=1.495
+ $X2=8.165 $Y2=0.445
r124 7 31 68.2186 $w=2.46e-07 $l=3.47059e-07 $layer=POLY_cond $X=8.14 $Y=1.99
+ $X2=8.105 $Y2=1.66
r125 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=8.14 $Y=1.99
+ $X2=8.14 $Y2=2.275
r126 2 20 600 $w=1.7e-07 $l=3.38748e-07 $layer=licon1_PDIFF $count=1 $X=6.11
+ $Y=2.065 $X2=6.265 $Y2=2.335
r127 1 16 182 $w=1.7e-07 $l=3.245e-07 $layer=licon1_NDIFF $count=1 $X=5.64
+ $Y=0.235 $X2=5.9 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_1%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 42 46 49
+ 50 52 53 55 56 58 59 61 76 87 92 93 96 99 102
r148 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r149 102 105 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=8.35 $Y=2.34
+ $X2=8.35 $Y2=2.72
r150 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r151 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r152 93 106 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=8.51 $Y2=2.72
r153 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r154 90 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.51 $Y2=2.72
r155 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r156 87 105 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.16 $Y=2.72
+ $X2=8.35 $Y2=2.72
r157 87 89 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=8.16 $Y=2.72
+ $X2=8.05 $Y2=2.72
r158 86 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r159 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r160 83 86 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=7.13 $Y2=2.72
r161 83 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r162 82 85 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.75 $Y=2.72
+ $X2=7.13 $Y2=2.72
r163 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r164 80 99 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=5.425 $Y=2.72
+ $X2=5.215 $Y2=2.72
r165 80 82 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.425 $Y=2.72
+ $X2=5.75 $Y2=2.72
r166 79 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r167 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r168 76 99 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=5.005 $Y=2.72
+ $X2=5.215 $Y2=2.72
r169 76 78 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.005 $Y=2.72
+ $X2=4.83 $Y2=2.72
r170 75 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r171 74 75 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r172 72 75 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.91 $Y2=2.72
r173 71 74 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.91 $Y2=2.72
r174 71 72 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r175 69 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r176 69 97 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r177 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r178 66 96 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r179 66 68 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r180 61 96 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r181 61 63 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r182 59 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r183 59 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r184 57 92 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.98 $Y=2.72
+ $X2=9.43 $Y2=2.72
r185 57 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.98 $Y=2.72
+ $X2=8.895 $Y2=2.72
r186 55 85 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.34 $Y=2.72
+ $X2=7.13 $Y2=2.72
r187 55 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.34 $Y=2.72
+ $X2=7.465 $Y2=2.72
r188 54 89 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r189 54 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.59 $Y=2.72
+ $X2=7.465 $Y2=2.72
r190 52 74 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.99 $Y=2.72 $X2=3.91
+ $Y2=2.72
r191 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.99 $Y=2.72
+ $X2=4.155 $Y2=2.72
r192 51 78 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.32 $Y=2.72
+ $X2=4.83 $Y2=2.72
r193 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=2.72
+ $X2=4.155 $Y2=2.72
r194 49 68 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.77 $Y=2.72
+ $X2=1.61 $Y2=2.72
r195 49 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.77 $Y=2.72
+ $X2=1.855 $Y2=2.72
r196 48 71 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.94 $Y=2.72
+ $X2=2.07 $Y2=2.72
r197 48 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.72
+ $X2=1.855 $Y2=2.72
r198 44 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.895 $Y=2.635
+ $X2=8.895 $Y2=2.72
r199 44 46 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.895 $Y=2.635
+ $X2=8.895 $Y2=2
r200 43 105 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.54 $Y=2.72
+ $X2=8.35 $Y2=2.72
r201 42 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.81 $Y=2.72
+ $X2=8.895 $Y2=2.72
r202 42 43 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.81 $Y=2.72
+ $X2=8.54 $Y2=2.72
r203 38 56 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.465 $Y=2.635
+ $X2=7.465 $Y2=2.72
r204 38 40 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=7.465 $Y=2.635
+ $X2=7.465 $Y2=2.34
r205 34 99 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=5.215 $Y=2.635
+ $X2=5.215 $Y2=2.72
r206 34 36 8.09454 $w=4.18e-07 $l=2.95e-07 $layer=LI1_cond $X=5.215 $Y=2.635
+ $X2=5.215 $Y2=2.34
r207 30 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=2.635
+ $X2=4.155 $Y2=2.72
r208 30 32 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.155 $Y=2.635
+ $X2=4.155 $Y2=2.29
r209 26 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=2.635
+ $X2=1.855 $Y2=2.72
r210 26 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.855 $Y=2.635
+ $X2=1.855 $Y2=2.34
r211 22 96 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r212 22 24 12.5859 $w=3.78e-07 $l=4.15e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.22
r213 7 46 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=8.77
+ $Y=1.485 $X2=8.895 $Y2=2
r214 6 102 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=8.23
+ $Y=2.065 $X2=8.375 $Y2=2.34
r215 5 40 600 $w=1.7e-07 $l=4.83322e-07 $layer=licon1_PDIFF $count=1 $X=7.06
+ $Y=2.065 $X2=7.425 $Y2=2.34
r216 4 36 600 $w=1.7e-07 $l=7.77592e-07 $layer=licon1_PDIFF $count=1 $X=5.065
+ $Y=1.645 $X2=5.24 $Y2=2.34
r217 3 32 600 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_PDIFF $count=1 $X=3.945
+ $Y=2.065 $X2=4.155 $Y2=2.29
r218 2 28 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=1.73
+ $Y=2.065 $X2=1.855 $Y2=2.34
r219 1 24 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.815 $X2=0.73 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_1%A_436_413# 1 2 8 12
c32 8 0 1.03144e-19 $X=2.16 $Y=1.835
r33 9 12 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.16 $Y=0.39 $X2=2.33
+ $Y2=0.39
r34 8 15 24.9307 $w=2.37e-07 $l=5.06636e-07 $layer=LI1_cond $X=2.16 $Y=1.835
+ $X2=2.247 $Y2=2.3
r35 7 9 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.475 $X2=2.16
+ $Y2=0.39
r36 7 8 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.16 $Y=0.475
+ $X2=2.16 $Y2=1.835
r37 2 15 600 $w=1.7e-07 $l=3.02738e-07 $layer=licon1_PDIFF $count=1 $X=2.18
+ $Y=2.065 $X2=2.335 $Y2=2.3
r38 1 12 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.19
+ $Y=0.235 $X2=2.33 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_1%A_649_413# 1 2 9 11 12 15
c37 12 0 3.1525e-19 $X=3.705 $Y=1.95
r38 13 15 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.625 $Y=2.035
+ $X2=4.625 $Y2=2.21
r39 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.54 $Y=1.95
+ $X2=4.625 $Y2=2.035
r40 11 12 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=4.54 $Y=1.95
+ $X2=3.705 $Y2=1.95
r41 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.62 $Y=2.035
+ $X2=3.705 $Y2=1.95
r42 7 9 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.62 $Y=2.035
+ $X2=3.62 $Y2=2.21
r43 2 15 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.48
+ $Y=2.065 $X2=4.625 $Y2=2.21
r44 1 9 600 $w=1.7e-07 $l=4.41588e-07 $layer=licon1_PDIFF $count=1 $X=3.245
+ $Y=2.065 $X2=3.62 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_1%Q 1 2 7 8 9 14 18
r15 24 26 23.3929 $w=3.33e-07 $l=6.8e-07 $layer=LI1_cond $X=9.407 $Y=1.62
+ $X2=9.407 $Y2=2.3
r16 9 24 3.09612 $w=3.33e-07 $l=9e-08 $layer=LI1_cond $X=9.407 $Y=1.53 $X2=9.407
+ $Y2=1.62
r17 8 9 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=9.407 $Y=1.19
+ $X2=9.407 $Y2=1.53
r18 8 18 11.1804 $w=3.33e-07 $l=3.25e-07 $layer=LI1_cond $X=9.407 $Y=1.19
+ $X2=9.407 $Y2=0.865
r19 7 18 0.516019 $w=3.33e-07 $l=1.5e-08 $layer=LI1_cond $X=9.407 $Y=0.85
+ $X2=9.407 $Y2=0.865
r20 7 14 14.7926 $w=3.33e-07 $l=4.3e-07 $layer=LI1_cond $X=9.407 $Y=0.85
+ $X2=9.407 $Y2=0.42
r21 2 26 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=9.22
+ $Y=1.485 $X2=9.365 $Y2=2.3
r22 2 24 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.22
+ $Y=1.485 $X2=9.365 $Y2=1.62
r23 1 14 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=9.23
+ $Y=0.235 $X2=9.365 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_1%VGND 1 2 3 4 5 16 20 24 28 32 35 36 38 39
+ 40 42 47 66 67 71 77 80
c138 67 0 2.71124e-20 $X=9.43 $Y=0
r139 80 81 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r140 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r141 72 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r142 71 74 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.38
r143 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r144 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r145 64 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=9.43
+ $Y2=0
r146 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r147 61 64 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.51 $Y2=0
r148 60 63 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=7.13 $Y=0 $X2=8.51
+ $Y2=0
r149 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r150 58 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r151 58 81 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=4.83 $Y2=0
r152 57 58 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r153 55 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.855 $Y=0 $X2=4.69
+ $Y2=0
r154 55 57 118.412 $w=1.68e-07 $l=1.815e-06 $layer=LI1_cond $X=4.855 $Y=0
+ $X2=6.67 $Y2=0
r155 54 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r156 53 54 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r157 51 54 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=4.37
+ $Y2=0
r158 51 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r159 50 53 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=4.37
+ $Y2=0
r160 50 51 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r161 48 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=1.74
+ $Y2=0
r162 48 50 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=0
+ $X2=2.07 $Y2=0
r163 47 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.525 $Y=0 $X2=4.69
+ $Y2=0
r164 47 53 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.525 $Y=0
+ $X2=4.37 $Y2=0
r165 42 71 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r166 42 44 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r167 40 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r168 40 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r169 38 63 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.81 $Y=0 $X2=8.51
+ $Y2=0
r170 38 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.81 $Y=0 $X2=8.895
+ $Y2=0
r171 37 66 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.98 $Y=0 $X2=9.43
+ $Y2=0
r172 37 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.98 $Y=0 $X2=8.895
+ $Y2=0
r173 35 57 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=6.825 $Y=0
+ $X2=6.67 $Y2=0
r174 35 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.825 $Y=0 $X2=6.91
+ $Y2=0
r175 34 60 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.995 $Y=0
+ $X2=7.13 $Y2=0
r176 34 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.995 $Y=0 $X2=6.91
+ $Y2=0
r177 30 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.895 $Y=0.085
+ $X2=8.895 $Y2=0
r178 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.895 $Y=0.085
+ $X2=8.895 $Y2=0.39
r179 26 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.91 $Y=0.085
+ $X2=6.91 $Y2=0
r180 26 28 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.91 $Y=0.085
+ $X2=6.91 $Y2=0.36
r181 22 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.69 $Y=0.085
+ $X2=4.69 $Y2=0
r182 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.69 $Y=0.085
+ $X2=4.69 $Y2=0.38
r183 18 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=0.085
+ $X2=1.74 $Y2=0
r184 18 20 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.74 $Y=0.085
+ $X2=1.74 $Y2=0.36
r185 17 71 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r186 16 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=0 $X2=1.74
+ $Y2=0
r187 16 17 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.575 $Y=0
+ $X2=0.895 $Y2=0
r188 5 32 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=8.77
+ $Y=0.235 $X2=8.895 $Y2=0.39
r189 4 28 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=6.765
+ $Y=0.235 $X2=6.91 $Y2=0.36
r190 3 24 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=4.385
+ $Y=0.235 $X2=4.69 $Y2=0.38
r191 2 20 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.74 $Y2=0.36
r192 1 74 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

