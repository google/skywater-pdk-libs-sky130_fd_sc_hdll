# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__einvp_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__einvp_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.020000 1.020000 9.050000 1.275000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  1.057500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.330000 1.615000 ;
    END
  END TE
  PIN VGND
    ANTENNADIFFAREA  1.014000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VPWR
    ANTENNADIFFAREA  1.360400 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  PIN Z
    ANTENNADIFFAREA  1.992000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.370000 0.635000 9.095000 0.850000 ;
        RECT 5.370000 0.850000 5.800000 1.445000 ;
        RECT 5.370000 1.445000 8.570000 1.615000 ;
        RECT 5.370000 1.615000 5.750000 2.125000 ;
        RECT 6.310000 1.615000 6.690000 2.125000 ;
        RECT 7.250000 1.615000 7.630000 2.125000 ;
        RECT 8.190000 1.615000 8.570000 2.125000 ;
    END
  END Z
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.745000 0.825000 ;
      RECT 0.085000  1.785000 0.925000 1.955000 ;
      RECT 0.085000  1.955000 0.345000 2.465000 ;
      RECT 0.500000  0.825000 0.745000 0.995000 ;
      RECT 0.500000  0.995000 5.200000 1.325000 ;
      RECT 0.500000  1.325000 0.925000 1.785000 ;
      RECT 0.515000  0.085000 0.895000 0.485000 ;
      RECT 0.515000  2.125000 0.925000 2.635000 ;
      RECT 1.135000  0.255000 1.305000 0.655000 ;
      RECT 1.135000  0.655000 5.200000 0.825000 ;
      RECT 1.175000  1.555000 5.200000 1.725000 ;
      RECT 1.175000  1.725000 1.385000 2.465000 ;
      RECT 1.475000  0.085000 1.855000 0.485000 ;
      RECT 1.605000  1.895000 1.935000 2.635000 ;
      RECT 2.075000  0.255000 2.245000 0.655000 ;
      RECT 2.155000  1.725000 2.325000 2.465000 ;
      RECT 2.415000  0.085000 2.795000 0.485000 ;
      RECT 2.545000  1.895000 2.875000 2.635000 ;
      RECT 3.015000  0.255000 3.185000 0.655000 ;
      RECT 3.095000  1.725000 3.265000 2.465000 ;
      RECT 3.355000  0.085000 3.735000 0.485000 ;
      RECT 3.485000  1.895000 3.815000 2.635000 ;
      RECT 3.955000  0.255000 4.125000 0.655000 ;
      RECT 4.035000  1.725000 4.205000 2.465000 ;
      RECT 4.295000  0.085000 4.685000 0.485000 ;
      RECT 4.425000  1.895000 4.755000 2.635000 ;
      RECT 4.855000  0.255000 9.095000 0.465000 ;
      RECT 4.855000  0.465000 5.200000 0.655000 ;
      RECT 4.975000  1.725000 5.200000 2.295000 ;
      RECT 4.975000  2.295000 9.095000 2.465000 ;
      RECT 5.970000  1.785000 6.140000 2.295000 ;
      RECT 6.910000  1.785000 7.080000 2.295000 ;
      RECT 7.850000  1.785000 8.020000 2.295000 ;
      RECT 8.790000  1.445000 9.095000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__einvp_8
END LIBRARY
