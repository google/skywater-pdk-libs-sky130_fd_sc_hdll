* File: sky130_fd_sc_hdll__buf_12.pxi.spice
* Created: Thu Aug 27 18:59:54 2020
* 
x_PM_SKY130_FD_SC_HDLL__BUF_12%A N_A_c_128_n N_A_M1001_g N_A_M1002_g N_A_c_129_n
+ N_A_M1011_g N_A_M1021_g N_A_c_130_n N_A_M1019_g N_A_M1022_g N_A_c_131_n
+ N_A_M1027_g N_A_M1031_g A A A A N_A_c_127_n A A A A
+ PM_SKY130_FD_SC_HDLL__BUF_12%A
x_PM_SKY130_FD_SC_HDLL__BUF_12%A_117_297# N_A_117_297#_M1002_s
+ N_A_117_297#_M1022_s N_A_117_297#_M1001_s N_A_117_297#_M1019_s
+ N_A_117_297#_M1006_g N_A_117_297#_c_227_n N_A_117_297#_M1000_g
+ N_A_117_297#_M1007_g N_A_117_297#_c_228_n N_A_117_297#_M1003_g
+ N_A_117_297#_M1010_g N_A_117_297#_c_229_n N_A_117_297#_M1004_g
+ N_A_117_297#_M1012_g N_A_117_297#_c_230_n N_A_117_297#_M1005_g
+ N_A_117_297#_M1014_g N_A_117_297#_c_231_n N_A_117_297#_M1008_g
+ N_A_117_297#_M1015_g N_A_117_297#_c_232_n N_A_117_297#_M1009_g
+ N_A_117_297#_M1017_g N_A_117_297#_c_233_n N_A_117_297#_M1013_g
+ N_A_117_297#_M1018_g N_A_117_297#_c_234_n N_A_117_297#_M1016_g
+ N_A_117_297#_M1024_g N_A_117_297#_c_235_n N_A_117_297#_M1020_g
+ N_A_117_297#_M1026_g N_A_117_297#_c_236_n N_A_117_297#_M1023_g
+ N_A_117_297#_M1028_g N_A_117_297#_c_237_n N_A_117_297#_M1025_g
+ N_A_117_297#_c_238_n N_A_117_297#_M1030_g N_A_117_297#_M1029_g
+ N_A_117_297#_c_247_n N_A_117_297#_c_250_n N_A_117_297#_c_218_n
+ N_A_117_297#_c_219_n N_A_117_297#_c_239_n N_A_117_297#_c_240_n
+ N_A_117_297#_c_266_n N_A_117_297#_c_269_n N_A_117_297#_c_220_n
+ N_A_117_297#_c_241_n N_A_117_297#_c_221_n N_A_117_297#_c_222_n
+ N_A_117_297#_c_223_n N_A_117_297#_c_243_n N_A_117_297#_c_224_n
+ N_A_117_297#_c_225_n N_A_117_297#_c_226_n
+ PM_SKY130_FD_SC_HDLL__BUF_12%A_117_297#
x_PM_SKY130_FD_SC_HDLL__BUF_12%VPWR N_VPWR_M1001_d N_VPWR_M1011_d N_VPWR_M1027_d
+ N_VPWR_M1003_d N_VPWR_M1005_d N_VPWR_M1009_d N_VPWR_M1016_d N_VPWR_M1023_d
+ N_VPWR_M1030_d N_VPWR_c_501_n N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n
+ N_VPWR_c_505_n N_VPWR_c_506_n N_VPWR_c_507_n N_VPWR_c_508_n N_VPWR_c_509_n
+ N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_512_n N_VPWR_c_513_n N_VPWR_c_514_n
+ VPWR VPWR N_VPWR_c_515_n N_VPWR_c_516_n N_VPWR_c_517_n N_VPWR_c_518_n
+ N_VPWR_c_500_n N_VPWR_c_520_n N_VPWR_c_521_n N_VPWR_c_522_n N_VPWR_c_523_n
+ N_VPWR_c_524_n N_VPWR_c_525_n N_VPWR_c_526_n N_VPWR_c_527_n N_VPWR_c_528_n
+ VPWR VPWR PM_SKY130_FD_SC_HDLL__BUF_12%VPWR
x_PM_SKY130_FD_SC_HDLL__BUF_12%X N_X_M1006_s N_X_M1010_s N_X_M1014_s N_X_M1017_s
+ N_X_M1024_s N_X_M1028_s N_X_M1000_s N_X_M1004_s N_X_M1008_s N_X_M1013_s
+ N_X_M1020_s N_X_M1025_s N_X_c_663_n N_X_c_664_n N_X_c_649_n N_X_c_650_n
+ N_X_c_656_n N_X_c_657_n N_X_c_682_n N_X_c_683_n N_X_c_651_n N_X_c_658_n
+ N_X_c_693_n N_X_c_694_n N_X_c_652_n N_X_c_659_n N_X_c_704_n N_X_c_706_n
+ N_X_c_708_n N_X_c_711_n N_X_c_714_n N_X_c_653_n N_X_c_660_n N_X_c_654_n
+ N_X_c_661_n X N_X_c_725_n X X N_X_c_655_n PM_SKY130_FD_SC_HDLL__BUF_12%X
x_PM_SKY130_FD_SC_HDLL__BUF_12%VGND N_VGND_M1002_d N_VGND_M1021_d N_VGND_M1031_d
+ N_VGND_M1007_d N_VGND_M1012_d N_VGND_M1015_d N_VGND_M1018_d N_VGND_M1026_d
+ N_VGND_M1029_d N_VGND_c_833_n N_VGND_c_834_n N_VGND_c_835_n N_VGND_c_836_n
+ N_VGND_c_837_n N_VGND_c_838_n N_VGND_c_839_n N_VGND_c_840_n N_VGND_c_841_n
+ N_VGND_c_842_n N_VGND_c_843_n N_VGND_c_844_n N_VGND_c_845_n VGND VGND
+ N_VGND_c_846_n N_VGND_c_847_n N_VGND_c_848_n N_VGND_c_849_n N_VGND_c_850_n
+ N_VGND_c_851_n N_VGND_c_852_n N_VGND_c_853_n N_VGND_c_854_n N_VGND_c_855_n
+ N_VGND_c_856_n N_VGND_c_857_n N_VGND_c_858_n N_VGND_c_859_n N_VGND_c_860_n
+ PM_SKY130_FD_SC_HDLL__BUF_12%VGND
cc_1 VNB N_A_M1002_g 0.0240984f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_2 VNB N_A_M1021_g 0.0178804f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_3 VNB N_A_M1022_g 0.0183641f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_4 VNB N_A_M1031_g 0.0175026f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_5 VNB A 0.00806404f $X=-0.19 $Y=-0.24 $X2=1.52 $Y2=1.105
cc_6 VNB N_A_c_127_n 0.111751f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.212
cc_7 VNB N_A_117_297#_M1006_g 0.0180221f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_8 VNB N_A_117_297#_M1007_g 0.0181352f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_9 VNB N_A_117_297#_M1010_g 0.0181597f $X=-0.19 $Y=-0.24 $X2=0.195 $Y2=1.105
cc_10 VNB N_A_117_297#_M1012_g 0.0181597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_117_297#_M1014_g 0.0181597f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.212
cc_12 VNB N_A_117_297#_M1015_g 0.0181537f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.212
cc_13 VNB N_A_117_297#_M1017_g 0.0176554f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=1.175
cc_14 VNB N_A_117_297#_M1018_g 0.017151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_117_297#_M1024_g 0.017151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_117_297#_M1026_g 0.017151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_117_297#_M1028_g 0.0176309f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_117_297#_M1029_g 0.0241263f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_117_297#_c_218_n 0.00380791f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_117_297#_c_219_n 0.00138237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_117_297#_c_220_n 0.00166201f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_117_297#_c_221_n 0.00305801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_117_297#_c_222_n 0.00103736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_117_297#_c_223_n 0.00274061f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_117_297#_c_224_n 0.00114159f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_117_297#_c_225_n 0.00142427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_117_297#_c_226_n 0.301905f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_500_n 0.345644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_X_c_649_n 0.00380791f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.212
cc_30 VNB N_X_c_650_n 0.00129721f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=1.212
cc_31 VNB N_X_c_651_n 0.00380791f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=1.175
cc_32 VNB N_X_c_652_n 0.00337105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_X_c_653_n 0.00114174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_X_c_654_n 0.00114174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_X_c_655_n 0.00163811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_833_n 0.0115514f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_834_n 0.0192014f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.105
cc_38 VNB N_VGND_c_835_n 0.00205913f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_836_n 3.19622e-19 $X=-0.19 $Y=-0.24 $X2=0.385 $Y2=1.16
cc_40 VNB N_VGND_c_837_n 3.19622e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.212
cc_41 VNB N_VGND_c_838_n 3.19622e-19 $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=1.212
cc_42 VNB N_VGND_c_839_n 3.19622e-19 $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.212
cc_43 VNB N_VGND_c_840_n 0.0126624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_841_n 3.19622e-19 $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.19
cc_45 VNB N_VGND_c_842_n 0.0126632f $X=-0.19 $Y=-0.24 $X2=1.115 $Y2=1.175
cc_46 VNB N_VGND_c_843_n 3.19622e-19 $X=-0.19 $Y=-0.24 $X2=1.575 $Y2=1.19
cc_47 VNB N_VGND_c_844_n 0.0132691f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_845_n 0.00669629f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_846_n 0.0145015f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_847_n 0.013707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_848_n 0.0134547f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_849_n 0.0126449f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_850_n 0.0126449f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_851_n 0.0128037f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_852_n 0.399748f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_853_n 0.00574292f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_854_n 0.00503278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_855_n 0.00503278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_856_n 0.00503278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_857_n 0.00503278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_858_n 0.00503278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_859_n 0.00503278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_860_n 0.00577057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VPB N_A_c_128_n 0.0208995f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_65 VPB N_A_c_129_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_66 VPB N_A_c_130_n 0.0158856f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_67 VPB N_A_c_131_n 0.0159691f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_68 VPB N_A_c_127_n 0.0387716f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.212
cc_69 VPB N_A_117_297#_c_227_n 0.0164045f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_70 VPB N_A_117_297#_c_228_n 0.0154215f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_71 VPB N_A_117_297#_c_229_n 0.0157197f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=1.105
cc_72 VPB N_A_117_297#_c_230_n 0.0154404f $X=-0.19 $Y=1.305 $X2=0.385 $Y2=1.16
cc_73 VPB N_A_117_297#_c_231_n 0.0157197f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.212
cc_74 VPB N_A_117_297#_c_232_n 0.0154404f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_117_297#_c_233_n 0.0155735f $X=-0.19 $Y=1.305 $X2=1.115 $Y2=1.19
cc_76 VPB N_A_117_297#_c_234_n 0.015148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_117_297#_c_235_n 0.0154273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_117_297#_c_236_n 0.015148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_117_297#_c_237_n 0.0154273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_117_297#_c_238_n 0.0198847f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_117_297#_c_239_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_117_297#_c_240_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_117_297#_c_241_n 8.69551e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_117_297#_c_222_n 0.00256049f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_117_297#_c_243_n 0.00177041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_117_297#_c_226_n 0.0763953f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_501_n 0.0110239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_502_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.105
cc_89 VPB N_VPWR_c_503_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_504_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_505_n 0.00418552f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.212
cc_92 VPB N_VPWR_c_506_n 3.32195e-19 $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.212
cc_93 VPB N_VPWR_c_507_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=1.505 $Y2=1.16
cc_94 VPB N_VPWR_c_508_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_509_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.19
cc_96 VPB N_VPWR_c_510_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=1.115 $Y2=1.175
cc_97 VPB N_VPWR_c_511_n 0.0140826f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=1.175
cc_98 VPB N_VPWR_c_512_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_513_n 0.0140698f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_514_n 0.00691506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_515_n 0.0176752f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_516_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_517_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_518_n 0.0128037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_500_n 0.0552802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_520_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_521_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_522_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_523_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_524_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_525_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_526_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_527_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_528_n 0.00580385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_X_c_656_n 0.00254663f $X=-0.19 $Y=1.305 $X2=1.505 $Y2=1.16
cc_116 VPB N_X_c_657_n 0.00144538f $X=-0.19 $Y=1.305 $X2=1.505 $Y2=1.16
cc_117 VPB N_X_c_658_n 0.00254663f $X=-0.19 $Y=1.305 $X2=1.115 $Y2=1.19
cc_118 VPB N_X_c_659_n 0.00241328f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_X_c_660_n 0.00108853f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_X_c_661_n 0.00108853f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_X_c_655_n 0.00194871f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 N_A_M1031_g N_A_117_297#_M1006_g 0.0204987f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_123 N_A_c_131_n N_A_117_297#_c_227_n 0.0219169f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A_c_128_n N_A_117_297#_c_247_n 0.0202434f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A_c_129_n N_A_117_297#_c_247_n 0.0115459f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A_c_130_n N_A_117_297#_c_247_n 7.68612e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A_M1021_g N_A_117_297#_c_250_n 0.00442074f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_128 N_A_M1021_g N_A_117_297#_c_218_n 0.0111137f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_129 N_A_M1022_g N_A_117_297#_c_218_n 0.012417f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_130 A N_A_117_297#_c_218_n 0.0545404f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_131 N_A_c_127_n N_A_117_297#_c_218_n 0.00342143f $X=1.905 $Y=1.212 $X2=0
+ $Y2=0
cc_132 N_A_M1002_g N_A_117_297#_c_219_n 0.00124214f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_133 A N_A_117_297#_c_219_n 0.0138098f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_134 N_A_c_127_n N_A_117_297#_c_219_n 0.00308294f $X=1.905 $Y=1.212 $X2=0
+ $Y2=0
cc_135 N_A_c_129_n N_A_117_297#_c_239_n 0.0137916f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A_c_130_n N_A_117_297#_c_239_n 0.0101048f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_137 A N_A_117_297#_c_239_n 0.0394547f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_138 N_A_c_127_n N_A_117_297#_c_239_n 0.00720931f $X=1.905 $Y=1.212 $X2=0
+ $Y2=0
cc_139 N_A_c_128_n N_A_117_297#_c_240_n 0.0101861f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_c_129_n N_A_117_297#_c_240_n 0.00107777f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_141 A N_A_117_297#_c_240_n 0.0305808f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_142 N_A_c_127_n N_A_117_297#_c_240_n 0.0074788f $X=1.905 $Y=1.212 $X2=0 $Y2=0
cc_143 N_A_c_129_n N_A_117_297#_c_266_n 8.07084e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_130_n N_A_117_297#_c_266_n 0.0141618f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_c_131_n N_A_117_297#_c_266_n 0.0116562f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_M1031_g N_A_117_297#_c_269_n 0.00438651f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_147 N_A_M1031_g N_A_117_297#_c_220_n 0.0123787f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_148 A N_A_117_297#_c_220_n 0.00394409f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_149 N_A_c_127_n N_A_117_297#_c_220_n 2.2583e-19 $X=1.905 $Y=1.212 $X2=0 $Y2=0
cc_150 N_A_c_131_n N_A_117_297#_c_241_n 0.0150852f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_c_127_n N_A_117_297#_c_241_n 3.58038e-19 $X=1.905 $Y=1.212 $X2=0
+ $Y2=0
cc_152 N_A_M1031_g N_A_117_297#_c_221_n 0.00420813f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_153 N_A_c_131_n N_A_117_297#_c_222_n 8.37329e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_154 A N_A_117_297#_c_222_n 0.00181689f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_155 N_A_c_127_n N_A_117_297#_c_222_n 0.00368389f $X=1.905 $Y=1.212 $X2=0
+ $Y2=0
cc_156 N_A_c_130_n N_A_117_297#_c_243_n 0.00259297f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_c_131_n N_A_117_297#_c_243_n 0.00128924f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_158 A N_A_117_297#_c_243_n 0.0286323f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_159 N_A_c_127_n N_A_117_297#_c_243_n 0.00751302f $X=1.905 $Y=1.212 $X2=0
+ $Y2=0
cc_160 A N_A_117_297#_c_224_n 0.0138008f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_161 N_A_c_127_n N_A_117_297#_c_224_n 0.00308219f $X=1.905 $Y=1.212 $X2=0
+ $Y2=0
cc_162 A N_A_117_297#_c_225_n 0.01199f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_163 N_A_c_127_n N_A_117_297#_c_225_n 0.00195556f $X=1.905 $Y=1.212 $X2=0
+ $Y2=0
cc_164 N_A_c_127_n N_A_117_297#_c_226_n 0.0204987f $X=1.905 $Y=1.212 $X2=0 $Y2=0
cc_165 N_A_c_128_n N_VPWR_c_502_n 0.00643281f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_166 A N_VPWR_c_502_n 0.00528751f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_167 N_A_c_127_n N_VPWR_c_502_n 0.0030441f $X=1.905 $Y=1.212 $X2=0 $Y2=0
cc_168 N_A_c_129_n N_VPWR_c_503_n 0.0052072f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_c_130_n N_VPWR_c_503_n 0.004751f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_c_130_n N_VPWR_c_504_n 0.00597712f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_c_131_n N_VPWR_c_504_n 0.00673617f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A_c_131_n N_VPWR_c_505_n 0.0052072f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_c_128_n N_VPWR_c_500_n 0.010906f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_c_129_n N_VPWR_c_500_n 0.0118438f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_c_130_n N_VPWR_c_500_n 0.00999457f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A_c_131_n N_VPWR_c_500_n 0.011869f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A_c_128_n N_VPWR_c_520_n 0.00597712f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A_c_129_n N_VPWR_c_520_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_M1002_g N_VGND_c_834_n 0.00330805f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_180 A N_VGND_c_834_n 0.00908165f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_181 N_A_c_127_n N_VGND_c_834_n 0.00551024f $X=1.905 $Y=1.212 $X2=0 $Y2=0
cc_182 N_A_M1002_g N_VGND_c_835_n 6.39981e-19 $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_183 N_A_M1021_g N_VGND_c_835_n 0.0109953f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_184 N_A_M1022_g N_VGND_c_835_n 0.00162962f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_185 N_A_M1022_g N_VGND_c_836_n 6.55283e-19 $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_186 N_A_M1031_g N_VGND_c_836_n 0.011037f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_187 N_A_M1002_g N_VGND_c_846_n 0.00585385f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_188 N_A_M1021_g N_VGND_c_846_n 0.0020416f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_189 N_A_M1022_g N_VGND_c_847_n 0.00439206f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_190 N_A_M1031_g N_VGND_c_847_n 0.0020416f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_191 N_A_M1002_g N_VGND_c_852_n 0.0116684f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_192 N_A_M1021_g N_VGND_c_852_n 0.00288181f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_193 N_A_M1022_g N_VGND_c_852_n 0.00613946f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_194 N_A_M1031_g N_VGND_c_852_n 0.00288181f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_195 N_A_117_297#_c_239_n N_VPWR_M1011_d 0.00199888f $X=1.455 $Y=1.53 $X2=0
+ $Y2=0
cc_196 N_A_117_297#_c_241_n N_VPWR_M1027_d 0.00365803f $X=2.04 $Y=1.53 $X2=0
+ $Y2=0
cc_197 N_A_117_297#_c_247_n N_VPWR_c_502_n 0.0470327f $X=0.73 $Y=1.63 $X2=0
+ $Y2=0
cc_198 N_A_117_297#_c_247_n N_VPWR_c_503_n 0.0385613f $X=0.73 $Y=1.63 $X2=0
+ $Y2=0
cc_199 N_A_117_297#_c_239_n N_VPWR_c_503_n 0.0112848f $X=1.455 $Y=1.53 $X2=0
+ $Y2=0
cc_200 N_A_117_297#_c_266_n N_VPWR_c_503_n 0.0470327f $X=1.67 $Y=1.63 $X2=0
+ $Y2=0
cc_201 N_A_117_297#_c_266_n N_VPWR_c_504_n 0.0223557f $X=1.67 $Y=1.63 $X2=0
+ $Y2=0
cc_202 N_A_117_297#_c_227_n N_VPWR_c_505_n 0.00446011f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_203 N_A_117_297#_c_266_n N_VPWR_c_505_n 0.0385613f $X=1.67 $Y=1.63 $X2=0
+ $Y2=0
cc_204 N_A_117_297#_c_241_n N_VPWR_c_505_n 0.0118234f $X=2.04 $Y=1.53 $X2=0
+ $Y2=0
cc_205 N_A_117_297#_c_223_n N_VPWR_c_505_n 2.86056e-19 $X=4.75 $Y=1.16 $X2=0
+ $Y2=0
cc_206 N_A_117_297#_c_227_n N_VPWR_c_506_n 7.31091e-19 $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_207 N_A_117_297#_c_228_n N_VPWR_c_506_n 0.0156322f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_208 N_A_117_297#_c_229_n N_VPWR_c_506_n 0.0117392f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_209 N_A_117_297#_c_230_n N_VPWR_c_506_n 6.61031e-19 $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_210 N_A_117_297#_c_229_n N_VPWR_c_507_n 6.99539e-19 $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_211 N_A_117_297#_c_230_n N_VPWR_c_507_n 0.0154534f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_212 N_A_117_297#_c_231_n N_VPWR_c_507_n 0.0117392f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_213 N_A_117_297#_c_232_n N_VPWR_c_507_n 6.61031e-19 $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_214 N_A_117_297#_c_231_n N_VPWR_c_508_n 6.99539e-19 $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_215 N_A_117_297#_c_232_n N_VPWR_c_508_n 0.0154534f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_216 N_A_117_297#_c_233_n N_VPWR_c_508_n 0.0117392f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_217 N_A_117_297#_c_234_n N_VPWR_c_508_n 6.61031e-19 $X=5.665 $Y=1.41 $X2=0
+ $Y2=0
cc_218 N_A_117_297#_c_233_n N_VPWR_c_509_n 0.00622633f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_219 N_A_117_297#_c_234_n N_VPWR_c_509_n 0.00427505f $X=5.665 $Y=1.41 $X2=0
+ $Y2=0
cc_220 N_A_117_297#_c_233_n N_VPWR_c_510_n 6.99539e-19 $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_221 N_A_117_297#_c_234_n N_VPWR_c_510_n 0.0154534f $X=5.665 $Y=1.41 $X2=0
+ $Y2=0
cc_222 N_A_117_297#_c_235_n N_VPWR_c_510_n 0.0117392f $X=6.135 $Y=1.41 $X2=0
+ $Y2=0
cc_223 N_A_117_297#_c_236_n N_VPWR_c_510_n 6.61031e-19 $X=6.605 $Y=1.41 $X2=0
+ $Y2=0
cc_224 N_A_117_297#_c_226_n N_VPWR_c_510_n 9.18523e-19 $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_225 N_A_117_297#_c_235_n N_VPWR_c_511_n 0.00622633f $X=6.135 $Y=1.41 $X2=0
+ $Y2=0
cc_226 N_A_117_297#_c_236_n N_VPWR_c_511_n 0.00427505f $X=6.605 $Y=1.41 $X2=0
+ $Y2=0
cc_227 N_A_117_297#_c_235_n N_VPWR_c_512_n 6.99539e-19 $X=6.135 $Y=1.41 $X2=0
+ $Y2=0
cc_228 N_A_117_297#_c_236_n N_VPWR_c_512_n 0.0154534f $X=6.605 $Y=1.41 $X2=0
+ $Y2=0
cc_229 N_A_117_297#_c_237_n N_VPWR_c_512_n 0.0117392f $X=7.075 $Y=1.41 $X2=0
+ $Y2=0
cc_230 N_A_117_297#_c_238_n N_VPWR_c_512_n 6.61031e-19 $X=7.545 $Y=1.41 $X2=0
+ $Y2=0
cc_231 N_A_117_297#_c_226_n N_VPWR_c_512_n 9.18523e-19 $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_232 N_A_117_297#_c_237_n N_VPWR_c_513_n 0.00622633f $X=7.075 $Y=1.41 $X2=0
+ $Y2=0
cc_233 N_A_117_297#_c_238_n N_VPWR_c_513_n 0.00427505f $X=7.545 $Y=1.41 $X2=0
+ $Y2=0
cc_234 N_A_117_297#_c_237_n N_VPWR_c_514_n 8.37274e-19 $X=7.075 $Y=1.41 $X2=0
+ $Y2=0
cc_235 N_A_117_297#_c_238_n N_VPWR_c_514_n 0.022204f $X=7.545 $Y=1.41 $X2=0
+ $Y2=0
cc_236 N_A_117_297#_c_227_n N_VPWR_c_515_n 0.00702461f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_237 N_A_117_297#_c_228_n N_VPWR_c_515_n 0.00427505f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_238 N_A_117_297#_c_229_n N_VPWR_c_516_n 0.00622633f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_239 N_A_117_297#_c_230_n N_VPWR_c_516_n 0.00427505f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_240 N_A_117_297#_c_231_n N_VPWR_c_517_n 0.00622633f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_241 N_A_117_297#_c_232_n N_VPWR_c_517_n 0.00427505f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_242 N_A_117_297#_M1001_s N_VPWR_c_500_n 0.00231261f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_243 N_A_117_297#_M1019_s N_VPWR_c_500_n 0.00231261f $X=1.525 $Y=1.485 $X2=0
+ $Y2=0
cc_244 N_A_117_297#_c_227_n N_VPWR_c_500_n 0.0126126f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_245 N_A_117_297#_c_228_n N_VPWR_c_500_n 0.00740765f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_246 N_A_117_297#_c_229_n N_VPWR_c_500_n 0.010479f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_247 N_A_117_297#_c_230_n N_VPWR_c_500_n 0.00740765f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_248 N_A_117_297#_c_231_n N_VPWR_c_500_n 0.010479f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_249 N_A_117_297#_c_232_n N_VPWR_c_500_n 0.00740765f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_250 N_A_117_297#_c_233_n N_VPWR_c_500_n 0.010479f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_251 N_A_117_297#_c_234_n N_VPWR_c_500_n 0.00740765f $X=5.665 $Y=1.41 $X2=0
+ $Y2=0
cc_252 N_A_117_297#_c_235_n N_VPWR_c_500_n 0.010479f $X=6.135 $Y=1.41 $X2=0
+ $Y2=0
cc_253 N_A_117_297#_c_236_n N_VPWR_c_500_n 0.00740765f $X=6.605 $Y=1.41 $X2=0
+ $Y2=0
cc_254 N_A_117_297#_c_237_n N_VPWR_c_500_n 0.010479f $X=7.075 $Y=1.41 $X2=0
+ $Y2=0
cc_255 N_A_117_297#_c_238_n N_VPWR_c_500_n 0.00740765f $X=7.545 $Y=1.41 $X2=0
+ $Y2=0
cc_256 N_A_117_297#_c_247_n N_VPWR_c_500_n 0.0140101f $X=0.73 $Y=1.63 $X2=0
+ $Y2=0
cc_257 N_A_117_297#_c_266_n N_VPWR_c_500_n 0.0140101f $X=1.67 $Y=1.63 $X2=0
+ $Y2=0
cc_258 N_A_117_297#_c_247_n N_VPWR_c_520_n 0.0223557f $X=0.73 $Y=1.63 $X2=0
+ $Y2=0
cc_259 N_A_117_297#_M1006_g N_X_c_663_n 0.00462807f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_260 N_A_117_297#_c_227_n N_X_c_664_n 0.00771865f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A_117_297#_c_228_n N_X_c_664_n 0.00657309f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A_117_297#_M1007_g N_X_c_649_n 0.0115761f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_263 N_A_117_297#_M1010_g N_X_c_649_n 0.0120362f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_264 N_A_117_297#_c_223_n N_X_c_649_n 0.0538798f $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_265 N_A_117_297#_c_226_n N_X_c_649_n 0.00342143f $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_266 N_A_117_297#_M1006_g N_X_c_650_n 0.00167159f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_267 N_A_117_297#_c_220_n N_X_c_650_n 0.00988205f $X=2.04 $Y=0.82 $X2=0 $Y2=0
cc_268 N_A_117_297#_c_223_n N_X_c_650_n 0.0136633f $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_269 N_A_117_297#_c_226_n N_X_c_650_n 0.00308294f $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_270 N_A_117_297#_c_228_n N_X_c_656_n 0.0146085f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_271 N_A_117_297#_c_229_n N_X_c_656_n 0.0163255f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_272 N_A_117_297#_c_223_n N_X_c_656_n 0.0473195f $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_273 N_A_117_297#_c_226_n N_X_c_656_n 0.0106248f $X=7.545 $Y=1.217 $X2=0 $Y2=0
cc_274 N_A_117_297#_c_227_n N_X_c_657_n 0.00162552f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_275 N_A_117_297#_c_241_n N_X_c_657_n 0.00995523f $X=2.04 $Y=1.53 $X2=0 $Y2=0
cc_276 N_A_117_297#_c_223_n N_X_c_657_n 0.012145f $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_277 N_A_117_297#_c_226_n N_X_c_657_n 0.00418485f $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_278 N_A_117_297#_M1010_g N_X_c_682_n 0.00462807f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_279 N_A_117_297#_c_229_n N_X_c_683_n 0.00702928f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_280 N_A_117_297#_c_230_n N_X_c_683_n 0.00657309f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_281 N_A_117_297#_M1012_g N_X_c_651_n 0.0120914f $X=3.76 $Y=0.56 $X2=0 $Y2=0
cc_282 N_A_117_297#_M1014_g N_X_c_651_n 0.0120914f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_283 N_A_117_297#_c_223_n N_X_c_651_n 0.0538798f $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_284 N_A_117_297#_c_226_n N_X_c_651_n 0.00342143f $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_285 N_A_117_297#_c_230_n N_X_c_658_n 0.0149392f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_286 N_A_117_297#_c_231_n N_X_c_658_n 0.0163685f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_287 N_A_117_297#_c_223_n N_X_c_658_n 0.0473195f $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_288 N_A_117_297#_c_226_n N_X_c_658_n 0.0106248f $X=7.545 $Y=1.217 $X2=0 $Y2=0
cc_289 N_A_117_297#_M1014_g N_X_c_693_n 0.00462807f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_290 N_A_117_297#_c_231_n N_X_c_694_n 0.00702928f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_291 N_A_117_297#_c_232_n N_X_c_694_n 0.00657309f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_292 N_A_117_297#_M1015_g N_X_c_652_n 0.0120914f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_293 N_A_117_297#_M1017_g N_X_c_652_n 0.00943266f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_294 N_A_117_297#_c_223_n N_X_c_652_n 0.027297f $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_295 N_A_117_297#_c_226_n N_X_c_652_n 0.00336301f $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_296 N_A_117_297#_c_232_n N_X_c_659_n 0.0149392f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_297 N_A_117_297#_c_233_n N_X_c_659_n 0.0103795f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_298 N_A_117_297#_c_223_n N_X_c_659_n 0.0239764f $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_299 N_A_117_297#_c_226_n N_X_c_659_n 0.00950791f $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_300 N_A_117_297#_M1017_g N_X_c_704_n 0.00464678f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_301 N_A_117_297#_c_226_n N_X_c_704_n 4.53201e-19 $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_302 N_A_117_297#_M1024_g N_X_c_706_n 0.00464678f $X=6.11 $Y=0.56 $X2=0 $Y2=0
cc_303 N_A_117_297#_c_226_n N_X_c_706_n 4.53201e-19 $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_304 N_A_117_297#_c_235_n N_X_c_708_n 0.00704883f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_305 N_A_117_297#_c_236_n N_X_c_708_n 0.00659264f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_306 N_A_117_297#_c_226_n N_X_c_708_n 5.47843e-19 $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_307 N_A_117_297#_M1028_g N_X_c_711_n 0.00471006f $X=7.05 $Y=0.56 $X2=0 $Y2=0
cc_308 N_A_117_297#_M1029_g N_X_c_711_n 0.0017519f $X=7.57 $Y=0.56 $X2=0 $Y2=0
cc_309 N_A_117_297#_c_226_n N_X_c_711_n 5.90215e-19 $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_310 N_A_117_297#_c_237_n N_X_c_714_n 0.00704883f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_311 N_A_117_297#_c_238_n N_X_c_714_n 0.00289674f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_312 N_A_117_297#_c_226_n N_X_c_714_n 5.50932e-19 $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_313 N_A_117_297#_c_223_n N_X_c_653_n 0.0136633f $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_314 N_A_117_297#_c_226_n N_X_c_653_n 0.00308294f $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_315 N_A_117_297#_c_223_n N_X_c_660_n 0.012145f $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_316 N_A_117_297#_c_226_n N_X_c_660_n 0.00418485f $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_317 N_A_117_297#_c_223_n N_X_c_654_n 0.0136633f $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_318 N_A_117_297#_c_226_n N_X_c_654_n 0.00308294f $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_319 N_A_117_297#_c_223_n N_X_c_661_n 0.012145f $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_320 N_A_117_297#_c_226_n N_X_c_661_n 0.00418485f $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_321 N_A_117_297#_c_233_n N_X_c_725_n 0.00704883f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_322 N_A_117_297#_c_234_n N_X_c_725_n 0.00659264f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_323 N_A_117_297#_c_226_n N_X_c_725_n 5.47843e-19 $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_324 N_A_117_297#_M1015_g N_X_c_655_n 3.38631e-19 $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_325 N_A_117_297#_M1017_g N_X_c_655_n 0.00666252f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_326 N_A_117_297#_c_233_n N_X_c_655_n 0.00711085f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_327 N_A_117_297#_M1018_g N_X_c_655_n 0.0149581f $X=5.64 $Y=0.56 $X2=0 $Y2=0
cc_328 N_A_117_297#_c_234_n N_X_c_655_n 0.0146251f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_329 N_A_117_297#_M1024_g N_X_c_655_n 0.0149581f $X=6.11 $Y=0.56 $X2=0 $Y2=0
cc_330 N_A_117_297#_c_235_n N_X_c_655_n 0.0163897f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_331 N_A_117_297#_M1026_g N_X_c_655_n 0.0149581f $X=6.58 $Y=0.56 $X2=0 $Y2=0
cc_332 N_A_117_297#_c_236_n N_X_c_655_n 0.014573f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_333 N_A_117_297#_M1028_g N_X_c_655_n 0.014543f $X=7.05 $Y=0.56 $X2=0 $Y2=0
cc_334 N_A_117_297#_c_237_n N_X_c_655_n 0.015948f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_335 N_A_117_297#_c_238_n N_X_c_655_n 0.00320702f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_336 N_A_117_297#_M1029_g N_X_c_655_n 0.00549657f $X=7.57 $Y=0.56 $X2=0 $Y2=0
cc_337 N_A_117_297#_c_223_n N_X_c_655_n 0.0105888f $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_338 N_A_117_297#_c_226_n N_X_c_655_n 0.146392f $X=7.545 $Y=1.217 $X2=0 $Y2=0
cc_339 N_A_117_297#_c_218_n N_VGND_M1021_d 0.00213931f $X=1.585 $Y=0.82 $X2=0
+ $Y2=0
cc_340 N_A_117_297#_c_220_n N_VGND_M1031_d 0.00349935f $X=2.04 $Y=0.82 $X2=0
+ $Y2=0
cc_341 N_A_117_297#_c_250_n N_VGND_c_835_n 0.0231432f $X=0.73 $Y=0.56 $X2=0
+ $Y2=0
cc_342 N_A_117_297#_c_218_n N_VGND_c_835_n 0.0219272f $X=1.585 $Y=0.82 $X2=0
+ $Y2=0
cc_343 N_A_117_297#_M1006_g N_VGND_c_836_n 0.00850423f $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_344 N_A_117_297#_M1007_g N_VGND_c_836_n 5.8773e-19 $X=2.82 $Y=0.56 $X2=0
+ $Y2=0
cc_345 N_A_117_297#_c_269_n N_VGND_c_836_n 0.0227699f $X=1.67 $Y=0.56 $X2=0
+ $Y2=0
cc_346 N_A_117_297#_c_220_n N_VGND_c_836_n 0.0190274f $X=2.04 $Y=0.82 $X2=0
+ $Y2=0
cc_347 N_A_117_297#_c_223_n N_VGND_c_836_n 0.00197677f $X=4.75 $Y=1.16 $X2=0
+ $Y2=0
cc_348 N_A_117_297#_M1006_g N_VGND_c_837_n 5.66132e-19 $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_349 N_A_117_297#_M1007_g N_VGND_c_837_n 0.00806522f $X=2.82 $Y=0.56 $X2=0
+ $Y2=0
cc_350 N_A_117_297#_M1010_g N_VGND_c_837_n 0.00842615f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_351 N_A_117_297#_M1012_g N_VGND_c_837_n 5.8773e-19 $X=3.76 $Y=0.56 $X2=0
+ $Y2=0
cc_352 N_A_117_297#_M1010_g N_VGND_c_838_n 5.66132e-19 $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_353 N_A_117_297#_M1012_g N_VGND_c_838_n 0.00806522f $X=3.76 $Y=0.56 $X2=0
+ $Y2=0
cc_354 N_A_117_297#_M1014_g N_VGND_c_838_n 0.00842615f $X=4.23 $Y=0.56 $X2=0
+ $Y2=0
cc_355 N_A_117_297#_M1015_g N_VGND_c_838_n 5.8773e-19 $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_356 N_A_117_297#_M1014_g N_VGND_c_839_n 5.66132e-19 $X=4.23 $Y=0.56 $X2=0
+ $Y2=0
cc_357 N_A_117_297#_M1015_g N_VGND_c_839_n 0.00806522f $X=4.7 $Y=0.56 $X2=0
+ $Y2=0
cc_358 N_A_117_297#_M1017_g N_VGND_c_839_n 0.00842615f $X=5.17 $Y=0.56 $X2=0
+ $Y2=0
cc_359 N_A_117_297#_M1018_g N_VGND_c_839_n 5.8773e-19 $X=5.64 $Y=0.56 $X2=0
+ $Y2=0
cc_360 N_A_117_297#_M1017_g N_VGND_c_840_n 0.0035053f $X=5.17 $Y=0.56 $X2=0
+ $Y2=0
cc_361 N_A_117_297#_M1018_g N_VGND_c_840_n 0.00350562f $X=5.64 $Y=0.56 $X2=0
+ $Y2=0
cc_362 N_A_117_297#_M1017_g N_VGND_c_841_n 5.66132e-19 $X=5.17 $Y=0.56 $X2=0
+ $Y2=0
cc_363 N_A_117_297#_M1018_g N_VGND_c_841_n 0.00806522f $X=5.64 $Y=0.56 $X2=0
+ $Y2=0
cc_364 N_A_117_297#_M1024_g N_VGND_c_841_n 0.00842615f $X=6.11 $Y=0.56 $X2=0
+ $Y2=0
cc_365 N_A_117_297#_M1026_g N_VGND_c_841_n 5.8773e-19 $X=6.58 $Y=0.56 $X2=0
+ $Y2=0
cc_366 N_A_117_297#_c_226_n N_VGND_c_841_n 5.8778e-19 $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_367 N_A_117_297#_M1024_g N_VGND_c_842_n 0.00350562f $X=6.11 $Y=0.56 $X2=0
+ $Y2=0
cc_368 N_A_117_297#_M1026_g N_VGND_c_842_n 0.00350562f $X=6.58 $Y=0.56 $X2=0
+ $Y2=0
cc_369 N_A_117_297#_M1024_g N_VGND_c_843_n 5.66132e-19 $X=6.11 $Y=0.56 $X2=0
+ $Y2=0
cc_370 N_A_117_297#_M1026_g N_VGND_c_843_n 0.00806522f $X=6.58 $Y=0.56 $X2=0
+ $Y2=0
cc_371 N_A_117_297#_M1028_g N_VGND_c_843_n 0.00845883f $X=7.05 $Y=0.56 $X2=0
+ $Y2=0
cc_372 N_A_117_297#_M1029_g N_VGND_c_843_n 5.50819e-19 $X=7.57 $Y=0.56 $X2=0
+ $Y2=0
cc_373 N_A_117_297#_c_226_n N_VGND_c_843_n 5.8778e-19 $X=7.545 $Y=1.217 $X2=0
+ $Y2=0
cc_374 N_A_117_297#_M1028_g N_VGND_c_844_n 0.00350562f $X=7.05 $Y=0.56 $X2=0
+ $Y2=0
cc_375 N_A_117_297#_M1029_g N_VGND_c_844_n 0.00271402f $X=7.57 $Y=0.56 $X2=0
+ $Y2=0
cc_376 N_A_117_297#_M1028_g N_VGND_c_845_n 7.5279e-19 $X=7.05 $Y=0.56 $X2=0
+ $Y2=0
cc_377 N_A_117_297#_M1029_g N_VGND_c_845_n 0.0177043f $X=7.57 $Y=0.56 $X2=0
+ $Y2=0
cc_378 N_A_117_297#_c_250_n N_VGND_c_846_n 0.0115672f $X=0.73 $Y=0.56 $X2=0
+ $Y2=0
cc_379 N_A_117_297#_c_218_n N_VGND_c_846_n 0.00193889f $X=1.585 $Y=0.82 $X2=0
+ $Y2=0
cc_380 N_A_117_297#_c_218_n N_VGND_c_847_n 0.00248202f $X=1.585 $Y=0.82 $X2=0
+ $Y2=0
cc_381 N_A_117_297#_c_269_n N_VGND_c_847_n 0.0112022f $X=1.67 $Y=0.56 $X2=0
+ $Y2=0
cc_382 N_A_117_297#_c_220_n N_VGND_c_847_n 0.00193889f $X=2.04 $Y=0.82 $X2=0
+ $Y2=0
cc_383 N_A_117_297#_M1006_g N_VGND_c_848_n 0.0046653f $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_384 N_A_117_297#_M1007_g N_VGND_c_848_n 0.00350562f $X=2.82 $Y=0.56 $X2=0
+ $Y2=0
cc_385 N_A_117_297#_M1010_g N_VGND_c_849_n 0.00350562f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_386 N_A_117_297#_M1012_g N_VGND_c_849_n 0.00350562f $X=3.76 $Y=0.56 $X2=0
+ $Y2=0
cc_387 N_A_117_297#_M1014_g N_VGND_c_850_n 0.00350562f $X=4.23 $Y=0.56 $X2=0
+ $Y2=0
cc_388 N_A_117_297#_M1015_g N_VGND_c_850_n 0.00350562f $X=4.7 $Y=0.56 $X2=0
+ $Y2=0
cc_389 N_A_117_297#_M1002_s N_VGND_c_852_n 0.00486275f $X=0.595 $Y=0.235 $X2=0
+ $Y2=0
cc_390 N_A_117_297#_M1022_s N_VGND_c_852_n 0.00334116f $X=1.535 $Y=0.235 $X2=0
+ $Y2=0
cc_391 N_A_117_297#_M1006_g N_VGND_c_852_n 0.00809951f $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_392 N_A_117_297#_M1007_g N_VGND_c_852_n 0.00431759f $X=2.82 $Y=0.56 $X2=0
+ $Y2=0
cc_393 N_A_117_297#_M1010_g N_VGND_c_852_n 0.00431759f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_394 N_A_117_297#_M1012_g N_VGND_c_852_n 0.00431759f $X=3.76 $Y=0.56 $X2=0
+ $Y2=0
cc_395 N_A_117_297#_M1014_g N_VGND_c_852_n 0.00431759f $X=4.23 $Y=0.56 $X2=0
+ $Y2=0
cc_396 N_A_117_297#_M1015_g N_VGND_c_852_n 0.00431759f $X=4.7 $Y=0.56 $X2=0
+ $Y2=0
cc_397 N_A_117_297#_M1017_g N_VGND_c_852_n 0.00431701f $X=5.17 $Y=0.56 $X2=0
+ $Y2=0
cc_398 N_A_117_297#_M1018_g N_VGND_c_852_n 0.00431759f $X=5.64 $Y=0.56 $X2=0
+ $Y2=0
cc_399 N_A_117_297#_M1024_g N_VGND_c_852_n 0.00431759f $X=6.11 $Y=0.56 $X2=0
+ $Y2=0
cc_400 N_A_117_297#_M1026_g N_VGND_c_852_n 0.00431759f $X=6.58 $Y=0.56 $X2=0
+ $Y2=0
cc_401 N_A_117_297#_M1028_g N_VGND_c_852_n 0.00443737f $X=7.05 $Y=0.56 $X2=0
+ $Y2=0
cc_402 N_A_117_297#_M1029_g N_VGND_c_852_n 0.00522073f $X=7.57 $Y=0.56 $X2=0
+ $Y2=0
cc_403 N_A_117_297#_c_250_n N_VGND_c_852_n 0.0064623f $X=0.73 $Y=0.56 $X2=0
+ $Y2=0
cc_404 N_A_117_297#_c_218_n N_VGND_c_852_n 0.0104775f $X=1.585 $Y=0.82 $X2=0
+ $Y2=0
cc_405 N_A_117_297#_c_269_n N_VGND_c_852_n 0.00644569f $X=1.67 $Y=0.56 $X2=0
+ $Y2=0
cc_406 N_A_117_297#_c_220_n N_VGND_c_852_n 0.00526647f $X=2.04 $Y=0.82 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_500_n N_X_M1000_s 0.00656398f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_408 N_VPWR_c_500_n N_X_M1004_s 0.00656398f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_409 N_VPWR_c_500_n N_X_M1008_s 0.00656398f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_410 N_VPWR_c_500_n N_X_M1013_s 0.00656398f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_411 N_VPWR_c_500_n N_X_M1020_s 0.00656398f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_412 N_VPWR_c_500_n N_X_M1025_s 0.00656398f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_413 N_VPWR_c_505_n N_X_c_664_n 0.0301172f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_414 N_VPWR_c_506_n N_X_c_664_n 0.0470327f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_415 N_VPWR_c_515_n N_X_c_664_n 0.0118139f $X=2.865 $Y=2.72 $X2=0 $Y2=0
cc_416 N_VPWR_c_500_n N_X_c_664_n 0.00646998f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_417 N_VPWR_M1003_d N_X_c_656_n 0.00209407f $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_418 N_VPWR_c_506_n N_X_c_656_n 0.0172025f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_419 N_VPWR_c_506_n N_X_c_683_n 0.0385613f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_420 N_VPWR_c_507_n N_X_c_683_n 0.0470327f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_421 N_VPWR_c_516_n N_X_c_683_n 0.0118139f $X=3.805 $Y=2.72 $X2=0 $Y2=0
cc_422 N_VPWR_c_500_n N_X_c_683_n 0.00646998f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_423 N_VPWR_M1005_d N_X_c_658_n 0.00209407f $X=3.875 $Y=1.485 $X2=0 $Y2=0
cc_424 N_VPWR_c_507_n N_X_c_658_n 0.0172025f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_425 N_VPWR_c_507_n N_X_c_694_n 0.0385613f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_426 N_VPWR_c_508_n N_X_c_694_n 0.0470327f $X=4.96 $Y=2 $X2=0 $Y2=0
cc_427 N_VPWR_c_517_n N_X_c_694_n 0.0118139f $X=4.745 $Y=2.72 $X2=0 $Y2=0
cc_428 N_VPWR_c_500_n N_X_c_694_n 0.00646998f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_429 N_VPWR_M1009_d N_X_c_659_n 0.00209407f $X=4.815 $Y=1.485 $X2=0 $Y2=0
cc_430 N_VPWR_c_508_n N_X_c_659_n 0.0172025f $X=4.96 $Y=2 $X2=0 $Y2=0
cc_431 N_VPWR_c_510_n N_X_c_708_n 0.0385613f $X=5.9 $Y=2 $X2=0 $Y2=0
cc_432 N_VPWR_c_511_n N_X_c_708_n 0.0118139f $X=6.625 $Y=2.72 $X2=0 $Y2=0
cc_433 N_VPWR_c_512_n N_X_c_708_n 0.0470327f $X=6.84 $Y=2 $X2=0 $Y2=0
cc_434 N_VPWR_c_500_n N_X_c_708_n 0.00646998f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_435 N_VPWR_c_512_n N_X_c_714_n 0.0385613f $X=6.84 $Y=2 $X2=0 $Y2=0
cc_436 N_VPWR_c_513_n N_X_c_714_n 0.0118139f $X=7.565 $Y=2.72 $X2=0 $Y2=0
cc_437 N_VPWR_c_514_n N_X_c_714_n 0.0634568f $X=7.78 $Y=1.66 $X2=0 $Y2=0
cc_438 N_VPWR_c_500_n N_X_c_714_n 0.00646998f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_439 N_VPWR_c_508_n N_X_c_725_n 0.0385613f $X=4.96 $Y=2 $X2=0 $Y2=0
cc_440 N_VPWR_c_509_n N_X_c_725_n 0.0118139f $X=5.685 $Y=2.72 $X2=0 $Y2=0
cc_441 N_VPWR_c_510_n N_X_c_725_n 0.0470327f $X=5.9 $Y=2 $X2=0 $Y2=0
cc_442 N_VPWR_c_500_n N_X_c_725_n 0.00646998f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_443 N_VPWR_M1016_d N_X_c_655_n 0.00218693f $X=5.755 $Y=1.485 $X2=0 $Y2=0
cc_444 N_VPWR_M1023_d N_X_c_655_n 0.00218693f $X=6.695 $Y=1.485 $X2=0 $Y2=0
cc_445 N_VPWR_c_510_n N_X_c_655_n 0.0190013f $X=5.9 $Y=2 $X2=0 $Y2=0
cc_446 N_VPWR_c_512_n N_X_c_655_n 0.0190013f $X=6.84 $Y=2 $X2=0 $Y2=0
cc_447 N_VPWR_c_514_n N_X_c_655_n 0.0107588f $X=7.78 $Y=1.66 $X2=0 $Y2=0
cc_448 N_VPWR_c_514_n N_VGND_c_845_n 0.0107865f $X=7.78 $Y=1.66 $X2=0 $Y2=0
cc_449 N_X_c_649_n N_VGND_M1007_d 0.00213931f $X=3.465 $Y=0.82 $X2=0 $Y2=0
cc_450 N_X_c_651_n N_VGND_M1012_d 0.00213931f $X=4.405 $Y=0.82 $X2=0 $Y2=0
cc_451 N_X_c_652_n N_VGND_M1015_d 0.00213931f $X=5.21 $Y=0.82 $X2=0 $Y2=0
cc_452 N_X_c_655_n N_VGND_M1018_d 0.00223254f $X=7.31 $Y=1.175 $X2=0 $Y2=0
cc_453 N_X_c_655_n N_VGND_M1026_d 0.00223254f $X=7.31 $Y=1.175 $X2=0 $Y2=0
cc_454 N_X_c_663_n N_VGND_c_836_n 0.0189749f $X=2.61 $Y=0.56 $X2=0 $Y2=0
cc_455 N_X_c_649_n N_VGND_c_837_n 0.0203425f $X=3.465 $Y=0.82 $X2=0 $Y2=0
cc_456 N_X_c_682_n N_VGND_c_837_n 0.0189749f $X=3.55 $Y=0.56 $X2=0 $Y2=0
cc_457 N_X_c_651_n N_VGND_c_838_n 0.0203425f $X=4.405 $Y=0.82 $X2=0 $Y2=0
cc_458 N_X_c_693_n N_VGND_c_838_n 0.0189749f $X=4.49 $Y=0.56 $X2=0 $Y2=0
cc_459 N_X_c_652_n N_VGND_c_839_n 0.0203425f $X=5.21 $Y=0.82 $X2=0 $Y2=0
cc_460 N_X_c_704_n N_VGND_c_839_n 0.0189749f $X=5.43 $Y=0.56 $X2=0 $Y2=0
cc_461 N_X_c_652_n N_VGND_c_840_n 0.0011009f $X=5.21 $Y=0.82 $X2=0 $Y2=0
cc_462 N_X_c_704_n N_VGND_c_840_n 0.0113207f $X=5.43 $Y=0.56 $X2=0 $Y2=0
cc_463 N_X_c_655_n N_VGND_c_840_n 0.00372499f $X=7.31 $Y=1.175 $X2=0 $Y2=0
cc_464 N_X_c_706_n N_VGND_c_841_n 0.0189749f $X=6.37 $Y=0.56 $X2=0 $Y2=0
cc_465 N_X_c_655_n N_VGND_c_841_n 0.0223861f $X=7.31 $Y=1.175 $X2=0 $Y2=0
cc_466 N_X_c_706_n N_VGND_c_842_n 0.0113207f $X=6.37 $Y=0.56 $X2=0 $Y2=0
cc_467 N_X_c_655_n N_VGND_c_842_n 0.00494036f $X=7.31 $Y=1.175 $X2=0 $Y2=0
cc_468 N_X_c_711_n N_VGND_c_843_n 0.0189749f $X=7.31 $Y=0.56 $X2=0 $Y2=0
cc_469 N_X_c_655_n N_VGND_c_843_n 0.0223861f $X=7.31 $Y=1.175 $X2=0 $Y2=0
cc_470 N_X_c_711_n N_VGND_c_844_n 0.0115192f $X=7.31 $Y=0.56 $X2=0 $Y2=0
cc_471 N_X_c_655_n N_VGND_c_844_n 0.00285443f $X=7.31 $Y=1.175 $X2=0 $Y2=0
cc_472 N_X_c_711_n N_VGND_c_845_n 0.0358347f $X=7.31 $Y=0.56 $X2=0 $Y2=0
cc_473 N_X_c_655_n N_VGND_c_845_n 0.0124269f $X=7.31 $Y=1.175 $X2=0 $Y2=0
cc_474 N_X_c_663_n N_VGND_c_848_n 0.0115672f $X=2.61 $Y=0.56 $X2=0 $Y2=0
cc_475 N_X_c_649_n N_VGND_c_848_n 0.00193763f $X=3.465 $Y=0.82 $X2=0 $Y2=0
cc_476 N_X_c_649_n N_VGND_c_849_n 0.00259419f $X=3.465 $Y=0.82 $X2=0 $Y2=0
cc_477 N_X_c_682_n N_VGND_c_849_n 0.0115672f $X=3.55 $Y=0.56 $X2=0 $Y2=0
cc_478 N_X_c_651_n N_VGND_c_849_n 0.00193763f $X=4.405 $Y=0.82 $X2=0 $Y2=0
cc_479 N_X_c_651_n N_VGND_c_850_n 0.00259419f $X=4.405 $Y=0.82 $X2=0 $Y2=0
cc_480 N_X_c_693_n N_VGND_c_850_n 0.0115672f $X=4.49 $Y=0.56 $X2=0 $Y2=0
cc_481 N_X_c_652_n N_VGND_c_850_n 0.00193763f $X=5.21 $Y=0.82 $X2=0 $Y2=0
cc_482 N_X_M1006_s N_VGND_c_852_n 0.00632385f $X=2.425 $Y=0.235 $X2=0 $Y2=0
cc_483 N_X_M1010_s N_VGND_c_852_n 0.00332158f $X=3.365 $Y=0.235 $X2=0 $Y2=0
cc_484 N_X_M1014_s N_VGND_c_852_n 0.00332158f $X=4.305 $Y=0.235 $X2=0 $Y2=0
cc_485 N_X_M1017_s N_VGND_c_852_n 0.00334669f $X=5.245 $Y=0.235 $X2=0 $Y2=0
cc_486 N_X_M1024_s N_VGND_c_852_n 0.00334789f $X=6.185 $Y=0.235 $X2=0 $Y2=0
cc_487 N_X_M1028_s N_VGND_c_852_n 0.00697884f $X=7.125 $Y=0.235 $X2=0 $Y2=0
cc_488 N_X_c_663_n N_VGND_c_852_n 0.0064623f $X=2.61 $Y=0.56 $X2=0 $Y2=0
cc_489 N_X_c_649_n N_VGND_c_852_n 0.0104569f $X=3.465 $Y=0.82 $X2=0 $Y2=0
cc_490 N_X_c_682_n N_VGND_c_852_n 0.0064623f $X=3.55 $Y=0.56 $X2=0 $Y2=0
cc_491 N_X_c_651_n N_VGND_c_852_n 0.0104569f $X=4.405 $Y=0.82 $X2=0 $Y2=0
cc_492 N_X_c_693_n N_VGND_c_852_n 0.0064623f $X=4.49 $Y=0.56 $X2=0 $Y2=0
cc_493 N_X_c_652_n N_VGND_c_852_n 0.00710219f $X=5.21 $Y=0.82 $X2=0 $Y2=0
cc_494 N_X_c_704_n N_VGND_c_852_n 0.00641247f $X=5.43 $Y=0.56 $X2=0 $Y2=0
cc_495 N_X_c_706_n N_VGND_c_852_n 0.00641247f $X=6.37 $Y=0.56 $X2=0 $Y2=0
cc_496 N_X_c_711_n N_VGND_c_852_n 0.00641247f $X=7.31 $Y=0.56 $X2=0 $Y2=0
cc_497 N_X_c_655_n N_VGND_c_852_n 0.0263292f $X=7.31 $Y=1.175 $X2=0 $Y2=0
