* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
M1000 a_444_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.7e+11p pd=5.14e+06u as=9.35e+11p ps=7.87e+06u
M1001 VPWR A1 a_444_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 X a_80_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.5e+11p pd=2.7e+06u as=0p ps=0u
M1003 X a_80_21# VGND VNB nshort w=650000u l=150000u
+  ad=2.795e+11p pd=2.16e+06u as=8.5475e+11p ps=6.53e+06u
M1004 a_444_297# B1 a_80_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.25e+11p ps=2.65e+06u
M1005 VPWR a_80_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_80_21# B1 VGND VNB nshort w=650000u l=150000u
+  ad=3.185e+11p pd=2.28e+06u as=0p ps=0u
M1007 VGND a_80_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_532_47# A1 a_80_21# VNB nshort w=650000u l=150000u
+  ad=2.3725e+11p pd=2.03e+06u as=0p ps=0u
M1009 VGND A2 a_532_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
