* File: sky130_fd_sc_hdll__xor2_1.pex.spice
* Created: Wed Sep  2 08:54:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__XOR2_1%B 1 3 4 6 7 9 10 12 14 18 21 22 28
c76 14 0 7.44272e-20 $X=1.805 $Y=1.445
c77 7 0 1.89107e-19 $X=1.965 $Y=1.41
c78 1 0 1.3377e-19 $X=0.535 $Y=1.41
r79 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.57
+ $Y=1.16 $X2=0.57 $Y2=1.16
r80 22 30 5.34211 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.6 $Y=1.53
+ $X2=0.775 $Y2=1.53
r81 22 28 8.05816 $w=4.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.6 $Y=1.445
+ $X2=0.6 $Y2=1.16
r82 22 30 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.8 $Y=1.53
+ $X2=0.775 $Y2=1.53
r83 21 22 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.72 $Y=1.53 $X2=0.8
+ $Y2=1.53
r84 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.93
+ $Y=1.16 $X2=1.93 $Y2=1.16
r85 15 18 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.805 $Y=1.16
+ $X2=1.93 $Y2=1.16
r86 14 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.805 $Y=1.445
+ $X2=1.72 $Y2=1.53
r87 13 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.805 $Y=1.245
+ $X2=1.805 $Y2=1.16
r88 13 14 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.805 $Y=1.245
+ $X2=1.805 $Y2=1.445
r89 10 19 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.99 $Y=0.995
+ $X2=1.93 $Y2=1.16
r90 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.99 $Y=0.995
+ $X2=1.99 $Y2=0.56
r91 7 19 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.965 $Y=1.41
+ $X2=1.93 $Y2=1.16
r92 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.965 $Y=1.41
+ $X2=1.965 $Y2=1.985
r93 4 27 39.2931 $w=2.55e-07 $l=1.69926e-07 $layer=POLY_cond $X=0.56 $Y=0.995
+ $X2=0.57 $Y2=1.16
r94 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.56 $Y=0.995 $X2=0.56
+ $Y2=0.56
r95 1 27 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=0.535 $Y=1.41
+ $X2=0.57 $Y2=1.16
r96 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.535 $Y=1.41
+ $X2=0.535 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_1%A 1 3 4 6 7 9 10 12 13 20
c43 13 0 1.89107e-19 $X=1.16 $Y=1.19
r44 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.485 $Y=1.202
+ $X2=1.51 $Y2=1.202
r45 18 20 35.5158 $w=3.8e-07 $l=2.8e-07 $layer=POLY_cond $X=1.205 $Y=1.202
+ $X2=1.485 $Y2=1.202
r46 16 18 24.1 $w=3.8e-07 $l=1.9e-07 $layer=POLY_cond $X=1.015 $Y=1.202
+ $X2=1.205 $Y2=1.202
r47 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.99 $Y=1.202
+ $X2=1.015 $Y2=1.202
r48 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.205
+ $Y=1.16 $X2=1.205 $Y2=1.16
r49 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=1.202
r50 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=0.56
r51 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.202
r52 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.985
r53 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.015 $Y=1.41
+ $X2=1.015 $Y2=1.202
r54 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.015 $Y=1.41
+ $X2=1.015 $Y2=1.985
r55 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r56 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995 $X2=0.99
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_1%A_35_297# 1 2 7 9 10 12 15 17 19 20 23 25
+ 29 32 33 35
c79 35 0 7.44272e-20 $X=2.955 $Y=1.202
c80 33 0 1.3377e-19 $X=0.77 $Y=0.74
r81 35 36 3.32873 $w=3.62e-07 $l=2.5e-08 $layer=POLY_cond $X=2.955 $Y=1.202
+ $X2=2.98 $Y2=1.202
r82 30 35 39.279 $w=3.62e-07 $l=2.95e-07 $layer=POLY_cond $X=2.66 $Y=1.202
+ $X2=2.955 $Y2=1.202
r83 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.66
+ $Y=1.16 $X2=2.66 $Y2=1.16
r84 27 29 16.7856 $w=2.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.63 $Y=0.825
+ $X2=2.63 $Y2=1.16
r85 26 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.855 $Y=0.74
+ $X2=0.77 $Y2=0.74
r86 25 27 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.515 $Y=0.74
+ $X2=2.63 $Y2=0.825
r87 25 26 108.299 $w=1.68e-07 $l=1.66e-06 $layer=LI1_cond $X=2.515 $Y=0.74
+ $X2=0.855 $Y2=0.74
r88 21 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=0.655
+ $X2=0.77 $Y2=0.74
r89 21 23 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.77 $Y=0.655
+ $X2=0.77 $Y2=0.5
r90 19 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=0.74
+ $X2=0.77 $Y2=0.74
r91 19 20 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=0.685 $Y=0.74
+ $X2=0.255 $Y2=0.74
r92 15 32 9.32938 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=0.275 $Y=1.975
+ $X2=0.275 $Y2=1.785
r93 15 17 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=0.275 $Y=1.975
+ $X2=0.275 $Y2=2
r94 13 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.255 $Y2=0.74
r95 13 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=1.785
r96 10 36 23.4391 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.98 $Y=0.995
+ $X2=2.98 $Y2=1.202
r97 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.98 $Y=0.995
+ $X2=2.98 $Y2=0.56
r98 7 35 19.0988 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.955 $Y=1.41
+ $X2=2.955 $Y2=1.202
r99 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.955 $Y=1.41
+ $X2=2.955 $Y2=1.985
r100 2 17 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.175
+ $Y=1.485 $X2=0.3 $Y2=2
r101 1 23 182 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_NDIFF $count=1 $X=0.635
+ $Y=0.235 $X2=0.77 $Y2=0.5
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_1%VPWR 1 2 9 13 16 17 19 20 21 37 38
r44 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r45 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r46 34 37 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r47 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r48 32 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r49 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r50 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r51 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r52 24 28 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r53 21 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r54 21 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r55 19 31 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.115 $Y=2.72
+ $X2=2.07 $Y2=2.72
r56 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.115 $Y=2.72 $X2=2.2
+ $Y2=2.72
r57 18 34 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.285 $Y=2.72
+ $X2=2.53 $Y2=2.72
r58 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.285 $Y=2.72 $X2=2.2
+ $Y2=2.72
r59 16 28 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.165 $Y=2.72
+ $X2=1.15 $Y2=2.72
r60 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.165 $Y=2.72
+ $X2=1.25 $Y2=2.72
r61 15 31 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=2.07 $Y2=2.72
r62 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.25 $Y2=2.72
r63 11 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=2.635 $X2=2.2
+ $Y2=2.72
r64 11 13 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.2 $Y=2.635 $X2=2.2
+ $Y2=2.29
r65 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=2.635 $X2=1.25
+ $Y2=2.72
r66 7 9 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.25 $Y=2.635
+ $X2=1.25 $Y2=1.95
r67 2 13 600 $w=1.7e-07 $l=8.745e-07 $layer=licon1_PDIFF $count=1 $X=2.055
+ $Y=1.485 $X2=2.2 $Y2=2.29
r68 1 9 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=1.105
+ $Y=1.485 $X2=1.25 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_1%A_315_297# 1 2 9 14 16
r24 10 14 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.885 $Y=1.87
+ $X2=1.695 $Y2=1.87
r25 9 16 5.87433 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.455 $Y=1.87 $X2=2.655
+ $Y2=1.87
r26 9 10 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.455 $Y=1.87
+ $X2=1.885 $Y2=1.87
r27 2 16 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=2.595
+ $Y=1.485 $X2=2.72 $Y2=1.95
r28 1 14 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=1.575
+ $Y=1.485 $X2=1.72 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_1%X 1 2 7 12 13 27
r25 16 22 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.385 $Y=1.45 $X2=3
+ $Y2=1.45
r26 13 27 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.4 $Y=1.45 $X2=3.405
+ $Y2=1.45
r27 13 16 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.4 $Y=1.45
+ $X2=3.385 $Y2=1.45
r28 13 20 26.11 $w=3.18e-07 $l=7.25e-07 $layer=LI1_cond $X=3.385 $Y=1.575
+ $X2=3.385 $Y2=2.3
r29 13 16 1.44055 $w=3.18e-07 $l=4e-08 $layer=LI1_cond $X=3.385 $Y=1.575
+ $X2=3.385 $Y2=1.535
r30 12 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=1.365 $X2=3
+ $Y2=1.45
r31 11 12 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=3 $Y=0.485 $X2=3
+ $Y2=1.365
r32 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.915 $Y=0.4 $X2=3
+ $Y2=0.485
r33 7 9 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.915 $Y=0.4 $X2=2.7
+ $Y2=0.4
r34 2 20 400 $w=1.7e-07 $l=9.46837e-07 $layer=licon1_PDIFF $count=1 $X=3.045
+ $Y=1.485 $X2=3.33 $Y2=2.3
r35 2 13 400 $w=1.7e-07 $l=3.45977e-07 $layer=licon1_PDIFF $count=1 $X=3.045
+ $Y=1.485 $X2=3.33 $Y2=1.62
r36 1 9 91 $w=1.7e-07 $l=7.12741e-07 $layer=licon1_NDIFF $count=2 $X=2.065
+ $Y=0.235 $X2=2.7 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_1%VGND 1 2 3 10 12 16 18 20 22 24 29 41 45
r48 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r49 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r50 36 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r51 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r52 33 36 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.99
+ $Y2=0
r53 33 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r54 32 35 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.99
+ $Y2=0
r55 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r56 30 41 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.415 $Y=0 $X2=1.225
+ $Y2=0
r57 30 32 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.415 $Y=0 $X2=1.61
+ $Y2=0
r58 29 44 4.33193 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.467
+ $Y2=0
r59 29 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=2.99
+ $Y2=0
r60 28 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r61 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r62 25 38 4.68787 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=0 $X2=0.232
+ $Y2=0
r63 25 27 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.465 $Y=0 $X2=0.69
+ $Y2=0
r64 24 41 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.225
+ $Y2=0
r65 24 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r66 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r67 22 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r68 18 44 3.10591 $w=2.9e-07 $l=1.13666e-07 $layer=LI1_cond $X=3.4 $Y=0.085
+ $X2=3.467 $Y2=0
r69 18 20 13.114 $w=2.88e-07 $l=3.3e-07 $layer=LI1_cond $X=3.4 $Y=0.085 $X2=3.4
+ $Y2=0.415
r70 14 41 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=0.085
+ $X2=1.225 $Y2=0
r71 14 16 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=1.225 $Y=0.085
+ $X2=1.225 $Y2=0.39
r72 10 38 3.0783 $w=3.3e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.3 $Y=0.085
+ $X2=0.232 $Y2=0
r73 10 12 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.3 $Y=0.085
+ $X2=0.3 $Y2=0.39
r74 3 20 91 $w=1.7e-07 $l=3.6404e-07 $layer=licon1_NDIFF $count=2 $X=3.055
+ $Y=0.235 $X2=3.34 $Y2=0.415
r75 2 16 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.25 $Y2=0.39
r76 1 12 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.235 $X2=0.3 $Y2=0.39
.ends

