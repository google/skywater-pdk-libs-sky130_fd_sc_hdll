* NGSPICE file created from sky130_fd_sc_hdll__clkbuf_8.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__clkbuf_8 A VGND VNB VPB VPWR X
M1000 VGND a_118_297# X VNB nshort w=420000u l=150000u
+  ad=7.791e+11p pd=8.75e+06u as=5.754e+11p ps=6.1e+06u
M1001 a_118_297# A VGND VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=0p ps=0u
M1002 VGND A a_118_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR a_118_297# X VPB phighvt w=1e+06u l=180000u
+  ad=1.75e+12p pd=1.55e+07u as=1.2e+12p ps=1.04e+07u
M1004 a_118_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1005 X a_118_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_118_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_118_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_118_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_118_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_118_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_118_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_118_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A a_118_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_118_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_118_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_118_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_118_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_118_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_118_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

