* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__inv_16 A VGND VNB VPB VPWR Y
M1000 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=2.57e+12p pd=2.314e+07u as=2.32e+12p ps=2.064e+07u
M1001 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VGND VNB nshort w=650000u l=150000u
+  ad=1.664e+12p pd=1.552e+07u as=1.8265e+12p ps=1.732e+07u
M1005 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
