* NGSPICE file created from sky130_fd_sc_hdll__o21a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
M1000 VPWR a_83_21# X VPB phighvt w=1e+06u l=180000u
+  ad=1.255e+12p pd=6.51e+06u as=2.9e+11p ps=2.58e+06u
M1001 a_394_297# A2 a_83_21# VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=3.6e+11p ps=2.72e+06u
M1002 VGND a_83_21# X VNB nshort w=650000u l=150000u
+  ad=3.835e+11p pd=3.78e+06u as=1.82e+11p ps=1.86e+06u
M1003 a_302_47# B1 a_83_21# VNB nshort w=650000u l=150000u
+  ad=3.445e+11p pd=3.66e+06u as=1.7225e+11p ps=1.83e+06u
M1004 VGND A2 a_302_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_83_21# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_394_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_302_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

