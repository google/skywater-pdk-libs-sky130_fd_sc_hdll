* File: sky130_fd_sc_hdll__inv_16.pex.spice
* Created: Wed Sep  2 08:32:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__INV_16%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 51 52 54 55 57 58 60 61 63
+ 64 66 67 69 70 72 73 75 76 78 79 81 82 84 85 87 88 90 91 93 94 96 97 98 99 100
+ 101 102 138 145 152 155 158 160 164
r289 158 160 48.2585 $w=2.38e-07 $l=1.005e-06 $layer=LI1_cond $X=3.295 $Y=1.195
+ $X2=4.3 $Y2=1.195
r290 145 146 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=7.61 $Y=1.202
+ $X2=7.635 $Y2=1.202
r291 144 145 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=7.165 $Y=1.202
+ $X2=7.61 $Y2=1.202
r292 143 144 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=7.14 $Y=1.202
+ $X2=7.165 $Y2=1.202
r293 142 143 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=6.695 $Y=1.202
+ $X2=7.14 $Y2=1.202
r294 141 142 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=6.67 $Y=1.202
+ $X2=6.695 $Y2=1.202
r295 140 141 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=6.225 $Y=1.202
+ $X2=6.67 $Y2=1.202
r296 139 140 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=6.2 $Y=1.202
+ $X2=6.225 $Y2=1.202
r297 138 164 53.5406 $w=2.38e-07 $l=1.115e-06 $layer=LI1_cond $X=5.96 $Y=1.195
+ $X2=4.845 $Y2=1.195
r298 137 139 31.6932 $w=3.65e-07 $l=2.4e-07 $layer=POLY_cond $X=5.96 $Y=1.202
+ $X2=6.2 $Y2=1.202
r299 137 138 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=5.96
+ $Y=1.16 $X2=5.96 $Y2=1.16
r300 135 137 27.0712 $w=3.65e-07 $l=2.05e-07 $layer=POLY_cond $X=5.755 $Y=1.202
+ $X2=5.96 $Y2=1.202
r301 134 135 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=5.73 $Y=1.202
+ $X2=5.755 $Y2=1.202
r302 133 134 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=5.285 $Y=1.202
+ $X2=5.73 $Y2=1.202
r303 132 133 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=5.26 $Y=1.202
+ $X2=5.285 $Y2=1.202
r304 131 132 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=4.815 $Y=1.202
+ $X2=5.26 $Y2=1.202
r305 130 131 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=4.79 $Y=1.202
+ $X2=4.815 $Y2=1.202
r306 129 130 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=4.345 $Y=1.202
+ $X2=4.79 $Y2=1.202
r307 128 129 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=4.32 $Y=1.202
+ $X2=4.345 $Y2=1.202
r308 127 128 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=3.875 $Y=1.202
+ $X2=4.32 $Y2=1.202
r309 126 127 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=3.85 $Y=1.202
+ $X2=3.875 $Y2=1.202
r310 125 126 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=3.405 $Y=1.202
+ $X2=3.85 $Y2=1.202
r311 124 125 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=3.38 $Y=1.202
+ $X2=3.405 $Y2=1.202
r312 123 124 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=2.935 $Y=1.202
+ $X2=3.38 $Y2=1.202
r313 122 123 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=2.91 $Y=1.202
+ $X2=2.935 $Y2=1.202
r314 121 122 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=2.465 $Y=1.202
+ $X2=2.91 $Y2=1.202
r315 120 121 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=2.44 $Y=1.202
+ $X2=2.465 $Y2=1.202
r316 119 120 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=1.995 $Y=1.202
+ $X2=2.44 $Y2=1.202
r317 118 119 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=1.97 $Y=1.202
+ $X2=1.995 $Y2=1.202
r318 117 118 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=1.525 $Y=1.202
+ $X2=1.97 $Y2=1.202
r319 116 117 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=1.5 $Y=1.202
+ $X2=1.525 $Y2=1.202
r320 115 116 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=1.055 $Y=1.202
+ $X2=1.5 $Y2=1.202
r321 114 115 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=1.03 $Y=1.202
+ $X2=1.055 $Y2=1.202
r322 113 114 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=0.585 $Y=1.202
+ $X2=1.03 $Y2=1.202
r323 112 113 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.56 $Y=1.202
+ $X2=0.585 $Y2=1.202
r324 110 112 34.9945 $w=3.65e-07 $l=2.65e-07 $layer=POLY_cond $X=0.295 $Y=1.202
+ $X2=0.56 $Y2=1.202
r325 102 164 1.20046 $w=2.38e-07 $l=2.5e-08 $layer=LI1_cond $X=4.82 $Y=1.195
+ $X2=4.845 $Y2=1.195
r326 101 102 24.4894 $w=2.38e-07 $l=5.1e-07 $layer=LI1_cond $X=4.31 $Y=1.195
+ $X2=4.82 $Y2=1.195
r327 101 160 0.480185 $w=2.38e-07 $l=1e-08 $layer=LI1_cond $X=4.31 $Y=1.195
+ $X2=4.3 $Y2=1.195
r328 100 158 0.240092 $w=2.38e-07 $l=5e-09 $layer=LI1_cond $X=3.29 $Y=1.195
+ $X2=3.295 $Y2=1.195
r329 100 155 48.0185 $w=2.38e-07 $l=1e-06 $layer=LI1_cond $X=3.29 $Y=1.195
+ $X2=2.29 $Y2=1.195
r330 99 155 0.960369 $w=2.38e-07 $l=2e-08 $layer=LI1_cond $X=2.27 $Y=1.195
+ $X2=2.29 $Y2=1.195
r331 99 152 48.7387 $w=2.38e-07 $l=1.015e-06 $layer=LI1_cond $X=2.27 $Y=1.195
+ $X2=1.255 $Y2=1.195
r332 98 152 0.240092 $w=2.38e-07 $l=5e-09 $layer=LI1_cond $X=1.25 $Y=1.195
+ $X2=1.255 $Y2=1.195
r333 97 98 48.9788 $w=2.38e-07 $l=1.02e-06 $layer=LI1_cond $X=0.23 $Y=1.195
+ $X2=1.25 $Y2=1.195
r334 97 110 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=0.295
+ $Y=1.16 $X2=0.295 $Y2=1.16
r335 94 146 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.635 $Y=0.995
+ $X2=7.635 $Y2=1.202
r336 94 96 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.635 $Y=0.995
+ $X2=7.635 $Y2=0.56
r337 91 145 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.61 $Y=1.41
+ $X2=7.61 $Y2=1.202
r338 91 93 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.61 $Y=1.41
+ $X2=7.61 $Y2=1.985
r339 88 144 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.165 $Y=0.995
+ $X2=7.165 $Y2=1.202
r340 88 90 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.165 $Y=0.995
+ $X2=7.165 $Y2=0.56
r341 85 143 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.14 $Y=1.41
+ $X2=7.14 $Y2=1.202
r342 85 87 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.14 $Y=1.41
+ $X2=7.14 $Y2=1.985
r343 82 142 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.695 $Y=0.995
+ $X2=6.695 $Y2=1.202
r344 82 84 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.695 $Y=0.995
+ $X2=6.695 $Y2=0.56
r345 79 141 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.67 $Y=1.41
+ $X2=6.67 $Y2=1.202
r346 79 81 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.67 $Y=1.41
+ $X2=6.67 $Y2=1.985
r347 76 140 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.225 $Y=0.995
+ $X2=6.225 $Y2=1.202
r348 76 78 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.225 $Y=0.995
+ $X2=6.225 $Y2=0.56
r349 73 139 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.2 $Y=1.41
+ $X2=6.2 $Y2=1.202
r350 73 75 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.2 $Y=1.41
+ $X2=6.2 $Y2=1.985
r351 70 135 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.755 $Y=0.995
+ $X2=5.755 $Y2=1.202
r352 70 72 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.755 $Y=0.995
+ $X2=5.755 $Y2=0.56
r353 67 134 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.73 $Y=1.41
+ $X2=5.73 $Y2=1.202
r354 67 69 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.73 $Y=1.41
+ $X2=5.73 $Y2=1.985
r355 64 133 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.285 $Y=0.995
+ $X2=5.285 $Y2=1.202
r356 64 66 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.285 $Y=0.995
+ $X2=5.285 $Y2=0.56
r357 61 132 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.26 $Y=1.41
+ $X2=5.26 $Y2=1.202
r358 61 63 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.26 $Y=1.41
+ $X2=5.26 $Y2=1.985
r359 58 131 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.815 $Y=0.995
+ $X2=4.815 $Y2=1.202
r360 58 60 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.815 $Y=0.995
+ $X2=4.815 $Y2=0.56
r361 55 130 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.79 $Y=1.41
+ $X2=4.79 $Y2=1.202
r362 55 57 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.79 $Y=1.41
+ $X2=4.79 $Y2=1.985
r363 52 129 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.345 $Y=0.995
+ $X2=4.345 $Y2=1.202
r364 52 54 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.345 $Y=0.995
+ $X2=4.345 $Y2=0.56
r365 49 128 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.32 $Y=1.41
+ $X2=4.32 $Y2=1.202
r366 49 51 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.32 $Y=1.41
+ $X2=4.32 $Y2=1.985
r367 46 127 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.875 $Y=0.995
+ $X2=3.875 $Y2=1.202
r368 46 48 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.875 $Y=0.995
+ $X2=3.875 $Y2=0.56
r369 43 126 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.85 $Y=1.41
+ $X2=3.85 $Y2=1.202
r370 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.85 $Y=1.41
+ $X2=3.85 $Y2=1.985
r371 40 125 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.405 $Y=0.995
+ $X2=3.405 $Y2=1.202
r372 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.405 $Y=0.995
+ $X2=3.405 $Y2=0.56
r373 37 124 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.202
r374 37 39 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.985
r375 34 123 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.935 $Y=0.995
+ $X2=2.935 $Y2=1.202
r376 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.935 $Y=0.995
+ $X2=2.935 $Y2=0.56
r377 31 122 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.91 $Y=1.41
+ $X2=2.91 $Y2=1.202
r378 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.91 $Y=1.41
+ $X2=2.91 $Y2=1.985
r379 28 121 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.465 $Y=0.995
+ $X2=2.465 $Y2=1.202
r380 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.465 $Y=0.995
+ $X2=2.465 $Y2=0.56
r381 25 120 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.44 $Y=1.41
+ $X2=2.44 $Y2=1.202
r382 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.44 $Y=1.41
+ $X2=2.44 $Y2=1.985
r383 22 119 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.995 $Y=0.995
+ $X2=1.995 $Y2=1.202
r384 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.995 $Y=0.995
+ $X2=1.995 $Y2=0.56
r385 19 118 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.97 $Y=1.41
+ $X2=1.97 $Y2=1.202
r386 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.97 $Y=1.41
+ $X2=1.97 $Y2=1.985
r387 16 117 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.525 $Y=0.995
+ $X2=1.525 $Y2=1.202
r388 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.525 $Y=0.995
+ $X2=1.525 $Y2=0.56
r389 13 116 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.5 $Y=1.41
+ $X2=1.5 $Y2=1.202
r390 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.5 $Y=1.41
+ $X2=1.5 $Y2=1.985
r391 10 115 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=1.055 $Y2=1.202
r392 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=1.055 $Y2=0.56
r393 7 114 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.03 $Y2=1.202
r394 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.03 $Y2=1.985
r395 4 113 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.585 $Y=0.995
+ $X2=0.585 $Y2=1.202
r396 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.585 $Y=0.995
+ $X2=0.585 $Y2=0.56
r397 1 112 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.56 $Y=1.41
+ $X2=0.56 $Y2=1.202
r398 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.56 $Y=1.41
+ $X2=0.56 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_16%VPWR 1 2 3 4 5 6 7 8 9 28 30 36 40 44 48 52
+ 56 60 64 67 68 70 71 73 74 76 77 79 80 82 83 85 86 88 89 90 118 119
r134 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r135 116 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r136 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r137 113 116 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r138 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r139 110 113 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r140 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r141 107 110 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r142 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r143 104 107 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r144 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r145 101 104 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r146 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r147 98 101 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r148 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r149 95 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r150 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r151 92 122 3.63491 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.41 $Y=2.72
+ $X2=0.205 $Y2=2.72
r152 92 94 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.41 $Y=2.72
+ $X2=1.15 $Y2=2.72
r153 90 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r154 90 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r155 88 115 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.76 $Y=2.72
+ $X2=7.59 $Y2=2.72
r156 88 89 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.76 $Y=2.72
+ $X2=7.865 $Y2=2.72
r157 87 118 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=7.97 $Y=2.72
+ $X2=8.05 $Y2=2.72
r158 87 89 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.97 $Y=2.72
+ $X2=7.865 $Y2=2.72
r159 85 112 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.82 $Y=2.72
+ $X2=6.67 $Y2=2.72
r160 85 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.82 $Y=2.72
+ $X2=6.905 $Y2=2.72
r161 84 115 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.99 $Y=2.72
+ $X2=7.59 $Y2=2.72
r162 84 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.99 $Y=2.72
+ $X2=6.905 $Y2=2.72
r163 82 109 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=5.88 $Y=2.72
+ $X2=5.75 $Y2=2.72
r164 82 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.88 $Y=2.72
+ $X2=5.965 $Y2=2.72
r165 81 112 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=6.05 $Y=2.72
+ $X2=6.67 $Y2=2.72
r166 81 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.05 $Y=2.72
+ $X2=5.965 $Y2=2.72
r167 79 106 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.94 $Y=2.72
+ $X2=4.83 $Y2=2.72
r168 79 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.94 $Y=2.72
+ $X2=5.025 $Y2=2.72
r169 78 109 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.11 $Y=2.72
+ $X2=5.75 $Y2=2.72
r170 78 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.11 $Y=2.72
+ $X2=5.025 $Y2=2.72
r171 76 103 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4 $Y=2.72 $X2=3.91
+ $Y2=2.72
r172 76 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4 $Y=2.72 $X2=4.085
+ $Y2=2.72
r173 75 106 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.17 $Y=2.72
+ $X2=4.83 $Y2=2.72
r174 75 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.17 $Y=2.72
+ $X2=4.085 $Y2=2.72
r175 73 100 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.06 $Y=2.72
+ $X2=2.99 $Y2=2.72
r176 73 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=2.72
+ $X2=3.145 $Y2=2.72
r177 72 103 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.23 $Y=2.72
+ $X2=3.91 $Y2=2.72
r178 72 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.23 $Y=2.72
+ $X2=3.145 $Y2=2.72
r179 70 97 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.12 $Y=2.72 $X2=2.07
+ $Y2=2.72
r180 70 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=2.72
+ $X2=2.205 $Y2=2.72
r181 69 100 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.29 $Y=2.72
+ $X2=2.99 $Y2=2.72
r182 69 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=2.72
+ $X2=2.205 $Y2=2.72
r183 67 94 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.18 $Y=2.72 $X2=1.15
+ $Y2=2.72
r184 67 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=2.72
+ $X2=1.265 $Y2=2.72
r185 66 97 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.35 $Y=2.72
+ $X2=2.07 $Y2=2.72
r186 66 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=2.72
+ $X2=1.265 $Y2=2.72
r187 62 89 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.865 $Y=2.635
+ $X2=7.865 $Y2=2.72
r188 62 64 33.5368 $w=2.08e-07 $l=6.35e-07 $layer=LI1_cond $X=7.865 $Y=2.635
+ $X2=7.865 $Y2=2
r189 58 86 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.905 $Y=2.635
+ $X2=6.905 $Y2=2.72
r190 58 60 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.905 $Y=2.635
+ $X2=6.905 $Y2=2
r191 54 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.965 $Y=2.635
+ $X2=5.965 $Y2=2.72
r192 54 56 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.965 $Y=2.635
+ $X2=5.965 $Y2=2
r193 50 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.025 $Y=2.635
+ $X2=5.025 $Y2=2.72
r194 50 52 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.025 $Y=2.635
+ $X2=5.025 $Y2=2
r195 46 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.085 $Y=2.635
+ $X2=4.085 $Y2=2.72
r196 46 48 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.085 $Y=2.635
+ $X2=4.085 $Y2=2
r197 42 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.145 $Y=2.635
+ $X2=3.145 $Y2=2.72
r198 42 44 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.145 $Y=2.635
+ $X2=3.145 $Y2=2
r199 38 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.205 $Y=2.635
+ $X2=2.205 $Y2=2.72
r200 38 40 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.205 $Y=2.635
+ $X2=2.205 $Y2=2
r201 34 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=2.635
+ $X2=1.265 $Y2=2.72
r202 34 36 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.265 $Y=2.635
+ $X2=1.265 $Y2=2
r203 30 33 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=0.305 $Y=1.65
+ $X2=0.305 $Y2=2.34
r204 28 122 3.28028 $w=2.1e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.305 $Y=2.635
+ $X2=0.205 $Y2=2.72
r205 28 33 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.305 $Y=2.635
+ $X2=0.305 $Y2=2.34
r206 9 64 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=7.7
+ $Y=1.485 $X2=7.845 $Y2=2
r207 8 60 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.76
+ $Y=1.485 $X2=6.905 $Y2=2
r208 7 56 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.82
+ $Y=1.485 $X2=5.965 $Y2=2
r209 6 52 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.88
+ $Y=1.485 $X2=5.025 $Y2=2
r210 5 48 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.94
+ $Y=1.485 $X2=4.085 $Y2=2
r211 4 44 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3
+ $Y=1.485 $X2=3.145 $Y2=2
r212 3 40 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.06
+ $Y=1.485 $X2=2.205 $Y2=2
r213 2 36 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.12
+ $Y=1.485 $X2=1.265 $Y2=2
r214 1 33 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.2
+ $Y=1.485 $X2=0.325 $Y2=2.34
r215 1 30 400 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=0.2
+ $Y=1.485 $X2=0.325 $Y2=1.65
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 51
+ 53 55 57 58 59 63 67 69 71 75 79 81 83 87 91 93 95 99 103 105 107 111 115 117
+ 119 123 127 129 131 135 139 143 145 146 148 149 151 152 154 155 157 158 160
+ 163 164 165
r295 164 169 2.39139 $w=4.52e-07 $l=9.5e-08 $layer=LI1_cond $X=7.277 $Y=0.81
+ $X2=7.277 $Y2=0.905
r296 164 165 6.15126 $w=5.23e-07 $l=2.7e-07 $layer=LI1_cond $X=7.277 $Y=0.92
+ $X2=7.277 $Y2=1.19
r297 164 169 0.341737 $w=5.23e-07 $l=1.5e-08 $layer=LI1_cond $X=7.277 $Y=0.92
+ $X2=7.277 $Y2=0.905
r298 161 165 6.94865 $w=5.23e-07 $l=3.05e-07 $layer=LI1_cond $X=7.277 $Y=1.495
+ $X2=7.277 $Y2=1.19
r299 161 163 2.15548 $w=4.52e-07 $l=8.5e-08 $layer=LI1_cond $X=7.277 $Y=1.495
+ $X2=7.277 $Y2=1.58
r300 137 163 2.15548 $w=4.52e-07 $l=1.15888e-07 $layer=LI1_cond $X=7.35 $Y=1.665
+ $X2=7.277 $Y2=1.58
r301 137 139 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=7.35 $Y=1.665
+ $X2=7.35 $Y2=2.34
r302 133 164 2.39139 $w=4.52e-07 $l=1.26333e-07 $layer=LI1_cond $X=7.35 $Y=0.715
+ $X2=7.277 $Y2=0.81
r303 133 135 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.35 $Y=0.715
+ $X2=7.35 $Y2=0.38
r304 132 160 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.6 $Y=1.58
+ $X2=6.41 $Y2=1.58
r305 131 163 5.01601 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=7.015 $Y=1.58
+ $X2=7.277 $Y2=1.58
r306 131 132 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=7.015 $Y=1.58
+ $X2=6.6 $Y2=1.58
r307 130 158 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=6.6 $Y=0.81
+ $X2=6.41 $Y2=0.81
r308 129 164 4.58964 $w=1.9e-07 $l=2.62e-07 $layer=LI1_cond $X=7.015 $Y=0.81
+ $X2=7.277 $Y2=0.81
r309 129 130 24.2249 $w=1.88e-07 $l=4.15e-07 $layer=LI1_cond $X=7.015 $Y=0.81
+ $X2=6.6 $Y2=0.81
r310 125 160 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.41 $Y=1.665
+ $X2=6.41 $Y2=1.58
r311 125 127 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=6.41 $Y=1.665
+ $X2=6.41 $Y2=2.34
r312 121 158 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=6.41 $Y=0.715
+ $X2=6.41 $Y2=0.81
r313 121 123 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.41 $Y=0.715
+ $X2=6.41 $Y2=0.38
r314 120 157 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.66 $Y=1.58
+ $X2=5.47 $Y2=1.58
r315 119 160 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.22 $Y=1.58
+ $X2=6.41 $Y2=1.58
r316 119 120 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.22 $Y=1.58
+ $X2=5.66 $Y2=1.58
r317 118 155 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=5.66 $Y=0.81
+ $X2=5.47 $Y2=0.81
r318 117 158 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=6.22 $Y=0.81
+ $X2=6.41 $Y2=0.81
r319 117 118 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=6.22 $Y=0.81
+ $X2=5.66 $Y2=0.81
r320 113 157 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.47 $Y=1.665
+ $X2=5.47 $Y2=1.58
r321 113 115 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=5.47 $Y=1.665
+ $X2=5.47 $Y2=2.34
r322 109 155 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=5.47 $Y=0.715
+ $X2=5.47 $Y2=0.81
r323 109 111 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.47 $Y=0.715
+ $X2=5.47 $Y2=0.38
r324 108 154 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.72 $Y=1.58
+ $X2=4.53 $Y2=1.58
r325 107 157 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.28 $Y=1.58
+ $X2=5.47 $Y2=1.58
r326 107 108 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.28 $Y=1.58
+ $X2=4.72 $Y2=1.58
r327 106 152 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=4.72 $Y=0.81
+ $X2=4.53 $Y2=0.81
r328 105 155 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=5.28 $Y=0.81
+ $X2=5.47 $Y2=0.81
r329 105 106 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=5.28 $Y=0.81
+ $X2=4.72 $Y2=0.81
r330 101 154 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.53 $Y=1.665
+ $X2=4.53 $Y2=1.58
r331 101 103 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=4.53 $Y=1.665
+ $X2=4.53 $Y2=2.34
r332 97 152 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=4.53 $Y=0.715
+ $X2=4.53 $Y2=0.81
r333 97 99 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.53 $Y=0.715
+ $X2=4.53 $Y2=0.38
r334 96 151 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.78 $Y=1.58
+ $X2=3.59 $Y2=1.58
r335 95 154 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.34 $Y=1.58
+ $X2=4.53 $Y2=1.58
r336 95 96 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.34 $Y=1.58
+ $X2=3.78 $Y2=1.58
r337 94 149 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=3.78 $Y=0.81
+ $X2=3.59 $Y2=0.81
r338 93 152 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=4.34 $Y=0.81
+ $X2=4.53 $Y2=0.81
r339 93 94 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=4.34 $Y=0.81
+ $X2=3.78 $Y2=0.81
r340 89 151 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.59 $Y=1.665
+ $X2=3.59 $Y2=1.58
r341 89 91 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=3.59 $Y=1.665
+ $X2=3.59 $Y2=2.34
r342 85 149 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=3.59 $Y=0.715
+ $X2=3.59 $Y2=0.81
r343 85 87 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.59 $Y=0.715
+ $X2=3.59 $Y2=0.38
r344 84 148 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.84 $Y=1.58
+ $X2=2.65 $Y2=1.58
r345 83 151 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.4 $Y=1.58
+ $X2=3.59 $Y2=1.58
r346 83 84 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.4 $Y=1.58
+ $X2=2.84 $Y2=1.58
r347 82 146 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=2.84 $Y=0.81
+ $X2=2.65 $Y2=0.81
r348 81 149 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=3.4 $Y=0.81
+ $X2=3.59 $Y2=0.81
r349 81 82 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=3.4 $Y=0.81 $X2=2.84
+ $Y2=0.81
r350 77 148 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.65 $Y=1.665
+ $X2=2.65 $Y2=1.58
r351 77 79 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=2.65 $Y=1.665
+ $X2=2.65 $Y2=2.34
r352 73 146 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.65 $Y=0.715
+ $X2=2.65 $Y2=0.81
r353 73 75 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.65 $Y=0.715
+ $X2=2.65 $Y2=0.38
r354 72 145 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.9 $Y=1.58
+ $X2=1.71 $Y2=1.58
r355 71 148 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.46 $Y=1.58
+ $X2=2.65 $Y2=1.58
r356 71 72 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.46 $Y=1.58
+ $X2=1.9 $Y2=1.58
r357 70 143 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=1.9 $Y=0.81
+ $X2=1.71 $Y2=0.81
r358 69 146 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=2.46 $Y=0.81
+ $X2=2.65 $Y2=0.81
r359 69 70 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=2.46 $Y=0.81 $X2=1.9
+ $Y2=0.81
r360 65 145 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=1.58
r361 65 67 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=2.34
r362 61 143 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=1.71 $Y=0.715
+ $X2=1.71 $Y2=0.81
r363 61 63 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.71 $Y=0.715
+ $X2=1.71 $Y2=0.38
r364 60 142 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.96 $Y=1.58
+ $X2=0.77 $Y2=1.58
r365 59 145 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.52 $Y=1.58
+ $X2=1.71 $Y2=1.58
r366 59 60 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.52 $Y=1.58
+ $X2=0.96 $Y2=1.58
r367 57 143 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=1.52 $Y=0.81
+ $X2=1.71 $Y2=0.81
r368 57 58 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=1.52 $Y=0.81
+ $X2=0.96 $Y2=0.81
r369 53 142 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=1.665
+ $X2=0.77 $Y2=1.58
r370 53 55 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.77 $Y=1.665
+ $X2=0.77 $Y2=2.34
r371 49 58 7.85115 $w=1.9e-07 $l=2.32702e-07 $layer=LI1_cond $X=0.77 $Y=0.715
+ $X2=0.96 $Y2=0.81
r372 49 51 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.77 $Y=0.715
+ $X2=0.77 $Y2=0.38
r373 16 163 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=7.23
+ $Y=1.485 $X2=7.375 $Y2=1.65
r374 16 139 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.23
+ $Y=1.485 $X2=7.375 $Y2=2.34
r375 15 160 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=6.29
+ $Y=1.485 $X2=6.435 $Y2=1.65
r376 15 127 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.29
+ $Y=1.485 $X2=6.435 $Y2=2.34
r377 14 157 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=5.35
+ $Y=1.485 $X2=5.495 $Y2=1.65
r378 14 115 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.35
+ $Y=1.485 $X2=5.495 $Y2=2.34
r379 13 154 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=4.41
+ $Y=1.485 $X2=4.555 $Y2=1.65
r380 13 103 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.41
+ $Y=1.485 $X2=4.555 $Y2=2.34
r381 12 151 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=3.47
+ $Y=1.485 $X2=3.615 $Y2=1.65
r382 12 91 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.47
+ $Y=1.485 $X2=3.615 $Y2=2.34
r383 11 148 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=2.53
+ $Y=1.485 $X2=2.675 $Y2=1.65
r384 11 79 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.53
+ $Y=1.485 $X2=2.675 $Y2=2.34
r385 10 145 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.485 $X2=1.735 $Y2=1.65
r386 10 67 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.485 $X2=1.735 $Y2=2.34
r387 9 142 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.485 $X2=0.795 $Y2=1.65
r388 9 55 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.485 $X2=0.795 $Y2=2.34
r389 8 135 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=7.24
+ $Y=0.235 $X2=7.375 $Y2=0.38
r390 7 123 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=6.3
+ $Y=0.235 $X2=6.435 $Y2=0.38
r391 6 111 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.36
+ $Y=0.235 $X2=5.495 $Y2=0.38
r392 5 99 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=4.42
+ $Y=0.235 $X2=4.555 $Y2=0.38
r393 4 87 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.48
+ $Y=0.235 $X2=3.615 $Y2=0.38
r394 3 75 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.54
+ $Y=0.235 $X2=2.675 $Y2=0.38
r395 2 63 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.6
+ $Y=0.235 $X2=1.735 $Y2=0.38
r396 1 51 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.66
+ $Y=0.235 $X2=0.795 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_16%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 50
+ 54 58 62 65 66 68 69 71 72 74 75 77 78 80 81 83 84 86 87 88 116 117
r149 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r150 114 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.05 $Y2=0
r151 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r152 111 114 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r153 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r154 108 111 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r155 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r156 105 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r157 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r158 102 105 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.83 $Y2=0
r159 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r160 99 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.91 $Y2=0
r161 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r162 96 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r163 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r164 93 96 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r165 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r166 90 120 3.78596 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.41 $Y=0
+ $X2=0.205 $Y2=0
r167 90 92 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.41 $Y=0 $X2=1.15
+ $Y2=0
r168 88 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r169 88 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r170 86 113 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.76 $Y=0 $X2=7.59
+ $Y2=0
r171 86 87 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.76 $Y=0 $X2=7.865
+ $Y2=0
r172 85 116 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=7.97 $Y=0 $X2=8.05
+ $Y2=0
r173 85 87 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.97 $Y=0 $X2=7.865
+ $Y2=0
r174 83 110 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.82 $Y=0 $X2=6.67
+ $Y2=0
r175 83 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.82 $Y=0 $X2=6.905
+ $Y2=0
r176 82 113 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.99 $Y=0 $X2=7.59
+ $Y2=0
r177 82 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.99 $Y=0 $X2=6.905
+ $Y2=0
r178 80 107 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=5.88 $Y=0 $X2=5.75
+ $Y2=0
r179 80 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.88 $Y=0 $X2=5.965
+ $Y2=0
r180 79 110 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=6.05 $Y=0 $X2=6.67
+ $Y2=0
r181 79 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.05 $Y=0 $X2=5.965
+ $Y2=0
r182 77 104 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.94 $Y=0 $X2=4.83
+ $Y2=0
r183 77 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.94 $Y=0 $X2=5.025
+ $Y2=0
r184 76 107 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.11 $Y=0 $X2=5.75
+ $Y2=0
r185 76 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.11 $Y=0 $X2=5.025
+ $Y2=0
r186 74 101 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4 $Y=0 $X2=3.91
+ $Y2=0
r187 74 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4 $Y=0 $X2=4.085
+ $Y2=0
r188 73 104 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.17 $Y=0 $X2=4.83
+ $Y2=0
r189 73 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.17 $Y=0 $X2=4.085
+ $Y2=0
r190 71 98 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.06 $Y=0 $X2=2.99
+ $Y2=0
r191 71 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=0 $X2=3.145
+ $Y2=0
r192 70 101 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.23 $Y=0 $X2=3.91
+ $Y2=0
r193 70 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.23 $Y=0 $X2=3.145
+ $Y2=0
r194 68 95 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.12 $Y=0 $X2=2.07
+ $Y2=0
r195 68 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=0 $X2=2.205
+ $Y2=0
r196 67 98 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.29 $Y=0 $X2=2.99
+ $Y2=0
r197 67 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=0 $X2=2.205
+ $Y2=0
r198 65 92 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.18 $Y=0 $X2=1.15
+ $Y2=0
r199 65 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=0 $X2=1.265
+ $Y2=0
r200 64 95 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.35 $Y=0 $X2=2.07
+ $Y2=0
r201 64 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.265
+ $Y2=0
r202 60 87 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.865 $Y=0.085
+ $X2=7.865 $Y2=0
r203 60 62 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=7.865 $Y=0.085
+ $X2=7.865 $Y2=0.38
r204 56 84 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.905 $Y=0.085
+ $X2=6.905 $Y2=0
r205 56 58 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.905 $Y=0.085
+ $X2=6.905 $Y2=0.38
r206 52 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.965 $Y=0.085
+ $X2=5.965 $Y2=0
r207 52 54 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.965 $Y=0.085
+ $X2=5.965 $Y2=0.38
r208 48 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.025 $Y=0.085
+ $X2=5.025 $Y2=0
r209 48 50 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.025 $Y=0.085
+ $X2=5.025 $Y2=0.38
r210 44 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.085 $Y=0.085
+ $X2=4.085 $Y2=0
r211 44 46 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.085 $Y=0.085
+ $X2=4.085 $Y2=0.38
r212 40 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.145 $Y=0.085
+ $X2=3.145 $Y2=0
r213 40 42 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.145 $Y=0.085
+ $X2=3.145 $Y2=0.38
r214 36 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.205 $Y=0.085
+ $X2=2.205 $Y2=0
r215 36 38 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.205 $Y=0.085
+ $X2=2.205 $Y2=0.38
r216 32 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=0.085
+ $X2=1.265 $Y2=0
r217 32 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.265 $Y=0.085
+ $X2=1.265 $Y2=0.38
r218 28 120 3.23192 $w=2.3e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.205 $Y2=0
r219 28 30 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.295 $Y2=0.38
r220 9 62 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=7.71
+ $Y=0.235 $X2=7.845 $Y2=0.38
r221 8 58 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.77
+ $Y=0.235 $X2=6.905 $Y2=0.38
r222 7 54 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.83
+ $Y=0.235 $X2=5.965 $Y2=0.38
r223 6 50 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.89
+ $Y=0.235 $X2=5.025 $Y2=0.38
r224 5 46 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.95
+ $Y=0.235 $X2=4.085 $Y2=0.38
r225 4 42 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.01
+ $Y=0.235 $X2=3.145 $Y2=0.38
r226 3 38 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.235 $X2=2.205 $Y2=0.38
r227 2 34 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.13
+ $Y=0.235 $X2=1.265 $Y2=0.38
r228 1 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.2
+ $Y=0.235 $X2=0.325 $Y2=0.38
.ends

