* File: sky130_fd_sc_hdll__o211a_2.pex.spice
* Created: Wed Sep  2 08:42:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O211A_2%C1 1 3 4 6 7 13
c21 4 0 1.69746e-19 $X=0.525 $Y=0.995
r22 7 13 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=1.16 $X2=0.23
+ $Y2=1.16
r23 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r24 4 10 41.0672 $w=4.66e-07 $l=2.41814e-07 $layer=POLY_cond $X=0.525 $Y=0.995
+ $X2=0.352 $Y2=1.16
r25 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.525 $Y=0.995
+ $X2=0.525 $Y2=0.56
r26 1 10 44.7433 $w=4.66e-07 $l=3.15436e-07 $layer=POLY_cond $X=0.5 $Y=1.41
+ $X2=0.352 $Y2=1.16
r27 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_2%B1 1 3 4 6 7 15
r29 7 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.065 $Y=1.16 $X2=1.155
+ $Y2=1.16
r30 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.065
+ $Y=1.16 $X2=1.065 $Y2=1.16
r31 4 10 45.6331 $w=3.55e-07 $l=2.94534e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=1.077 $Y2=1.16
r32 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.98 $Y=1.41 $X2=0.98
+ $Y2=1.985
r33 1 10 38.8445 $w=3.55e-07 $l=2.17612e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=1.077 $Y2=1.16
r34 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_2%A2 1 3 4 6 7 11 15
r27 11 15 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.81 $Y=1.16
+ $X2=1.64 $Y2=1.16
r28 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.81
+ $Y=1.16 $X2=1.81 $Y2=1.16
r29 7 15 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.635 $Y=1.16 $X2=1.64
+ $Y2=1.16
r30 4 10 40.1071 $w=4.25e-07 $l=2.26164e-07 $layer=POLY_cond $X=1.965 $Y=0.995
+ $X2=1.82 $Y2=1.16
r31 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.965 $Y=0.995
+ $X2=1.965 $Y2=0.56
r32 1 10 44.7315 $w=4.25e-07 $l=3.04138e-07 $layer=POLY_cond $X=1.94 $Y=1.41
+ $X2=1.82 $Y2=1.16
r33 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.94 $Y=1.41 $X2=1.94
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_2%A1 1 3 4 6 7 14
r31 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.415
+ $Y=1.16 $X2=2.415 $Y2=1.16
r32 7 14 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=2.525 $Y=1.16
+ $X2=2.415 $Y2=1.16
r33 4 10 38.5818 $w=3.27e-07 $l=1.67481e-07 $layer=POLY_cond $X=2.425 $Y=0.995
+ $X2=2.43 $Y2=1.16
r34 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.425 $Y=0.995
+ $X2=2.425 $Y2=0.56
r35 1 10 46.5183 $w=3.27e-07 $l=2.87228e-07 $layer=POLY_cond $X=2.35 $Y=1.41
+ $X2=2.43 $Y2=1.16
r36 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.35 $Y=1.41 $X2=2.35
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_2%A_27_47# 1 2 3 10 12 13 15 16 18 19 21 24
+ 27 28 29 32 34 37 38 40 47 49 53
r91 53 54 0.646113 $w=3.73e-07 $l=5e-09 $layer=POLY_cond $X=3.42 $Y=1.202
+ $X2=3.425 $Y2=1.202
r92 50 51 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=2.915 $Y=1.202
+ $X2=2.94 $Y2=1.202
r93 47 48 9.55876 $w=4.85e-07 $l=3.8e-07 $layer=LI1_cond $X=0.265 $Y=0.54
+ $X2=0.645 $Y2=0.54
r94 41 53 5.1689 $w=3.73e-07 $l=4e-08 $layer=POLY_cond $X=3.38 $Y=1.202 $X2=3.42
+ $Y2=1.202
r95 41 51 56.8579 $w=3.73e-07 $l=4.4e-07 $layer=POLY_cond $X=3.38 $Y=1.202
+ $X2=2.94 $Y2=1.202
r96 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.38
+ $Y=1.16 $X2=3.38 $Y2=1.16
r97 38 40 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.025 $Y=1.16
+ $X2=3.38 $Y2=1.16
r98 36 38 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.94 $Y=1.325
+ $X2=3.025 $Y2=1.16
r99 36 37 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.94 $Y=1.325
+ $X2=2.94 $Y2=1.51
r100 35 49 11.1863 $w=2.4e-07 $l=3.55421e-07 $layer=LI1_cond $X=1.82 $Y=1.622
+ $X2=1.472 $Y2=1.637
r101 34 37 6.9898 $w=2.25e-07 $l=1.4854e-07 $layer=LI1_cond $X=2.855 $Y=1.622
+ $X2=2.94 $Y2=1.51
r102 34 35 53.0124 $w=2.23e-07 $l=1.035e-06 $layer=LI1_cond $X=2.855 $Y=1.622
+ $X2=1.82 $Y2=1.622
r103 30 49 2.03437 $w=6.95e-07 $l=1.28e-07 $layer=LI1_cond $X=1.472 $Y=1.765
+ $X2=1.472 $Y2=1.637
r104 30 32 2.15122 $w=6.93e-07 $l=1.25e-07 $layer=LI1_cond $X=1.472 $Y=1.765
+ $X2=1.472 $Y2=1.89
r105 28 49 11.1863 $w=2.4e-07 $l=3.47e-07 $layer=LI1_cond $X=1.125 $Y=1.637
+ $X2=1.472 $Y2=1.637
r106 28 29 16.4958 $w=2.53e-07 $l=3.65e-07 $layer=LI1_cond $X=1.125 $Y=1.637
+ $X2=0.76 $Y2=1.637
r107 27 29 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=0.645 $Y=1.637
+ $X2=0.76 $Y2=1.637
r108 27 43 19.117 $w=2.53e-07 $l=4.23e-07 $layer=LI1_cond $X=0.645 $Y=1.637
+ $X2=0.222 $Y2=1.637
r109 26 48 5.11717 $w=2.3e-07 $l=2.85e-07 $layer=LI1_cond $X=0.645 $Y=0.825
+ $X2=0.645 $Y2=0.54
r110 26 27 34.3228 $w=2.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.645 $Y=0.825
+ $X2=0.645 $Y2=1.51
r111 22 43 0.504477 $w=2.65e-07 $l=1.28e-07 $layer=LI1_cond $X=0.222 $Y=1.765
+ $X2=0.222 $Y2=1.637
r112 22 24 2.39186 $w=2.63e-07 $l=5.5e-08 $layer=LI1_cond $X=0.222 $Y=1.765
+ $X2=0.222 $Y2=1.82
r113 19 54 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.425 $Y=0.995
+ $X2=3.425 $Y2=1.202
r114 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.425 $Y=0.995
+ $X2=3.425 $Y2=0.56
r115 16 53 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.42 $Y=1.41
+ $X2=3.42 $Y2=1.202
r116 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.42 $Y=1.41
+ $X2=3.42 $Y2=1.985
r117 13 51 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.94 $Y=1.41
+ $X2=2.94 $Y2=1.202
r118 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.94 $Y=1.41
+ $X2=2.94 $Y2=1.985
r119 10 50 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.915 $Y=0.995
+ $X2=2.915 $Y2=1.202
r120 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.915 $Y=0.995
+ $X2=2.915 $Y2=0.56
r121 3 32 150 $w=1.7e-07 $l=7.61019e-07 $layer=licon1_PDIFF $count=4 $X=1.07
+ $Y=1.485 $X2=1.655 $Y2=1.89
r122 2 24 300 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.82
r123 1 47 91 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.265 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_2%VPWR 1 2 3 12 16 18 20 22 27 37 38 41 44
+ 47
r53 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r54 47 50 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.635 $Y=2.34
+ $X2=3.635 $Y2=2.72
r55 45 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r56 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r57 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r58 38 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r59 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r60 35 50 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.825 $Y=2.72
+ $X2=3.635 $Y2=2.72
r61 35 37 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.825 $Y=2.72
+ $X2=3.91 $Y2=2.72
r62 34 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r63 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r64 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r65 31 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r66 30 33 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r67 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r68 28 41 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.905 $Y=2.72
+ $X2=0.715 $Y2=2.72
r69 28 30 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.905 $Y=2.72
+ $X2=1.15 $Y2=2.72
r70 27 44 11.015 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=2.375 $Y=2.72
+ $X2=2.615 $Y2=2.72
r71 27 33 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.375 $Y=2.72
+ $X2=2.07 $Y2=2.72
r72 22 41 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.715 $Y2=2.72
r73 22 24 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.23 $Y2=2.72
r74 20 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r75 20 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r76 19 44 11.015 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=2.855 $Y=2.72
+ $X2=2.615 $Y2=2.72
r77 18 50 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.445 $Y=2.72
+ $X2=3.635 $Y2=2.72
r78 18 19 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.445 $Y=2.72
+ $X2=2.855 $Y2=2.72
r79 14 44 1.96841 $w=4.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=2.635
+ $X2=2.615 $Y2=2.72
r80 14 16 15.3248 $w=4.78e-07 $l=6.15e-07 $layer=LI1_cond $X=2.615 $Y=2.635
+ $X2=2.615 $Y2=2.02
r81 10 41 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=2.635
+ $X2=0.715 $Y2=2.72
r82 10 12 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=0.715 $Y=2.635
+ $X2=0.715 $Y2=2.02
r83 3 47 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.51
+ $Y=1.485 $X2=3.66 $Y2=2.34
r84 2 16 300 $w=1.7e-07 $l=6.27077e-07 $layer=licon1_PDIFF $count=2 $X=2.44
+ $Y=1.485 $X2=2.64 $Y2=2.02
r85 1 12 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=1.485 $X2=0.74 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_2%X 1 2 9 11 12 13 16 22 25 27
r44 25 27 2.7744 $w=2.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.9 $Y=0.785 $X2=3.9
+ $Y2=0.85
r45 22 25 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.9 $Y=0.7 $X2=3.9
+ $Y2=0.785
r46 22 27 0.426831 $w=2.68e-07 $l=1e-08 $layer=LI1_cond $X=3.9 $Y=0.86 $X2=3.9
+ $Y2=0.85
r47 21 22 44.6038 $w=2.68e-07 $l=1.045e-06 $layer=LI1_cond $X=3.9 $Y=1.905
+ $X2=3.9 $Y2=0.86
r48 16 19 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=3.135 $Y=0.36
+ $X2=3.135 $Y2=0.7
r49 14 19 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.325 $Y=0.7
+ $X2=3.135 $Y2=0.7
r50 13 22 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.765 $Y=0.7 $X2=3.9
+ $Y2=0.7
r51 13 14 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.765 $Y=0.7
+ $X2=3.325 $Y2=0.7
r52 11 21 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.765 $Y=1.99
+ $X2=3.9 $Y2=1.905
r53 11 12 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.765 $Y=1.99
+ $X2=3.275 $Y2=1.99
r54 7 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.18 $Y=2.075
+ $X2=3.275 $Y2=1.99
r55 7 9 13.134 $w=1.88e-07 $l=2.25e-07 $layer=LI1_cond $X=3.18 $Y=2.075 $X2=3.18
+ $Y2=2.3
r56 2 9 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=3.03
+ $Y=1.485 $X2=3.18 $Y2=2.3
r57 1 19 182 $w=1.7e-07 $l=5.43392e-07 $layer=licon1_NDIFF $count=1 $X=2.99
+ $Y=0.235 $X2=3.16 $Y2=0.7
r58 1 16 182 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_NDIFF $count=1 $X=2.99
+ $Y=0.235 $X2=3.16 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_2%A_206_47# 1 2 11
c20 11 0 1.69746e-19 $X=2.21 $Y=0.73
r21 8 11 60.7081 $w=1.88e-07 $l=1.04e-06 $layer=LI1_cond $X=1.17 $Y=0.73
+ $X2=2.21 $Y2=0.73
r22 2 11 182 $w=1.7e-07 $l=5.73738e-07 $layer=licon1_NDIFF $count=1 $X=2.04
+ $Y=0.235 $X2=2.21 $Y2=0.73
r23 1 8 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.235 $X2=1.17 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211A_2%VGND 1 2 3 12 16 18 20 23 24 25 27 36 41
+ 45
r53 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r54 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r55 39 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r56 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r57 36 44 4.48746 $w=1.7e-07 $l=2.97e-07 $layer=LI1_cond $X=3.545 $Y=0 $X2=3.842
+ $Y2=0
r58 36 38 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.545 $Y=0 $X2=3.45
+ $Y2=0
r59 35 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r60 35 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r61 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r62 32 41 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.87 $Y=0 $X2=1.702
+ $Y2=0
r63 32 34 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.87 $Y=0 $X2=2.53
+ $Y2=0
r64 27 41 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.702
+ $Y2=0
r65 27 29 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=1.535 $Y=0 $X2=0.23
+ $Y2=0
r66 25 42 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r67 25 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r68 23 34 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.53
+ $Y2=0
r69 23 24 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.657
+ $Y2=0
r70 22 38 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=3.45
+ $Y2=0
r71 22 24 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.657
+ $Y2=0
r72 18 44 3.27872 $w=3.3e-07 $l=1.69245e-07 $layer=LI1_cond $X=3.71 $Y=0.085
+ $X2=3.842 $Y2=0
r73 18 20 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.71 $Y=0.085
+ $X2=3.71 $Y2=0.36
r74 14 24 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.657 $Y=0.085
+ $X2=2.657 $Y2=0
r75 14 16 13.486 $w=2.33e-07 $l=2.75e-07 $layer=LI1_cond $X=2.657 $Y=0.085
+ $X2=2.657 $Y2=0.36
r76 10 41 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.702 $Y=0.085
+ $X2=1.702 $Y2=0
r77 10 12 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=1.702 $Y=0.085
+ $X2=1.702 $Y2=0.38
r78 3 20 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.5
+ $Y=0.235 $X2=3.71 $Y2=0.36
r79 2 16 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=2.5
+ $Y=0.235 $X2=2.66 $Y2=0.36
r80 1 12 182 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_NDIFF $count=1 $X=1.575
+ $Y=0.235 $X2=1.705 $Y2=0.38
.ends

