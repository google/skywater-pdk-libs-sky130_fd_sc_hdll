* File: sky130_fd_sc_hdll__or3_2.pex.spice
* Created: Thu Aug 27 19:24:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR3_2%C 1 3 6 8 13
c25 13 0 1.66831e-19 $X=0.51 $Y=1.202
c26 8 0 1.91415e-19 $X=0.23 $Y=1.19
r27 13 14 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=0.51 $Y=1.202
+ $X2=0.535 $Y2=1.202
r28 11 13 33.7665 $w=3.64e-07 $l=2.55e-07 $layer=POLY_cond $X=0.255 $Y=1.202
+ $X2=0.51 $Y2=1.202
r29 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.255
+ $Y=1.16 $X2=0.255 $Y2=1.16
r30 4 14 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.535 $Y=0.995
+ $X2=0.535 $Y2=1.202
r31 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.535 $Y=0.995
+ $X2=0.535 $Y2=0.475
r32 1 13 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.41
+ $X2=0.51 $Y2=1.202
r33 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.51 $Y=1.41 $X2=0.51
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_2%B 2 3 4 6 9 10 11 12 13 14 25 29
c44 11 0 6.13246e-20 $X=0.95 $Y=0.91
c45 2 0 2.76319e-19 $X=0.92 $Y=1.31
r46 20 29 5.36482 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=0.985 $Y=2.27
+ $X2=1.12 $Y2=2.27
r47 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.985
+ $Y=2.28 $X2=0.985 $Y2=2.28
r48 14 29 1.98697 $w=2.88e-07 $l=5e-08 $layer=LI1_cond $X=1.17 $Y=2.27 $X2=1.12
+ $Y2=2.27
r49 13 20 10.7296 $w=2.88e-07 $l=2.7e-07 $layer=LI1_cond $X=0.715 $Y=2.27
+ $X2=0.985 $Y2=2.27
r50 13 25 1.98697 $w=2.88e-07 $l=5e-08 $layer=LI1_cond $X=0.715 $Y=2.27
+ $X2=0.665 $Y2=2.27
r51 12 25 17.2866 $w=2.88e-07 $l=4.35e-07 $layer=LI1_cond $X=0.23 $Y=2.27
+ $X2=0.665 $Y2=2.27
r52 10 11 54.0301 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=0.95 $Y=0.76 $X2=0.95
+ $Y2=0.91
r53 9 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.005 $Y=0.475
+ $X2=1.005 $Y2=0.76
r54 4 19 46.6963 $w=3.06e-07 $l=2.8e-07 $layer=POLY_cond $X=0.92 $Y=2.035
+ $X2=0.995 $Y2=2.28
r55 4 6 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=0.92 $Y=2.035 $X2=0.92
+ $Y2=1.695
r56 3 6 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.92 $Y=1.41 $X2=0.92
+ $Y2=1.695
r57 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.92 $Y=1.31 $X2=0.92
+ $Y2=1.41
r58 2 11 132.631 $w=2e-07 $l=4e-07 $layer=POLY_cond $X=0.92 $Y=1.31 $X2=0.92
+ $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_2%A 1 3 6 8 9 10 16 19 23
c51 16 0 1.66831e-19 $X=1.41 $Y=1.16
r52 17 23 0.623162 $w=3.3e-07 $l=1.63e-07 $layer=LI1_cond $X=0.88 $Y=1.16
+ $X2=0.717 $Y2=1.16
r53 17 19 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=0.88 $Y=1.16
+ $X2=1.15 $Y2=1.16
r54 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.41
+ $Y=1.16 $X2=1.41 $Y2=1.16
r55 10 16 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=1.165 $Y=1.16
+ $X2=1.41 $Y2=1.16
r56 10 19 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.165 $Y=1.16
+ $X2=1.15 $Y2=1.16
r57 8 9 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=0.717 $Y=1.19
+ $X2=0.717 $Y2=1.53
r58 8 23 1.06379 $w=3.23e-07 $l=3e-08 $layer=LI1_cond $X=0.717 $Y=1.19 $X2=0.717
+ $Y2=1.16
r59 4 15 38.578 $w=2.95e-07 $l=1.83916e-07 $layer=POLY_cond $X=1.475 $Y=0.995
+ $X2=1.435 $Y2=1.16
r60 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.475 $Y=0.995
+ $X2=1.475 $Y2=0.475
r61 1 15 48.1208 $w=2.95e-07 $l=2.57391e-07 $layer=POLY_cond $X=1.45 $Y=1.41
+ $X2=1.435 $Y2=1.16
r62 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.45 $Y=1.41 $X2=1.45
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_2%A_30_53# 1 2 3 10 12 13 15 16 18 19 21 24 28
+ 30 31 32 33 36 38 40 43 45 46 47 54 60
c112 45 0 1.24896e-19 $X=2 $Y=1.495
r113 60 61 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=2.65 $Y=1.202
+ $X2=2.675 $Y2=1.202
r114 57 58 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=2.155 $Y=1.202
+ $X2=2.18 $Y2=1.202
r115 55 60 55.1763 $w=3.8e-07 $l=4.35e-07 $layer=POLY_cond $X=2.215 $Y=1.202
+ $X2=2.65 $Y2=1.202
r116 55 58 4.43947 $w=3.8e-07 $l=3.5e-08 $layer=POLY_cond $X=2.215 $Y=1.202
+ $X2=2.18 $Y2=1.202
r117 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.215
+ $Y=1.16 $X2=2.215 $Y2=1.16
r118 51 54 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2 $Y=1.16
+ $X2=2.215 $Y2=1.16
r119 47 49 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.285 $Y=1.58
+ $X2=1.285 $Y2=1.87
r120 44 51 3.11056 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2 $Y=1.325 $X2=2
+ $Y2=1.16
r121 44 45 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=2 $Y=1.325 $X2=2
+ $Y2=1.495
r122 43 51 3.11056 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2 $Y=0.995 $X2=2
+ $Y2=1.16
r123 42 43 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=2 $Y=0.825 $X2=2
+ $Y2=0.995
r124 41 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=1.58
+ $X2=1.285 $Y2=1.58
r125 40 45 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.89 $Y=1.58
+ $X2=2 $Y2=1.495
r126 40 41 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.89 $Y=1.58
+ $X2=1.37 $Y2=1.58
r127 39 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=0.74
+ $X2=1.215 $Y2=0.74
r128 38 42 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.89 $Y=0.74
+ $X2=2 $Y2=0.825
r129 38 39 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.89 $Y=0.74 $X2=1.3
+ $Y2=0.74
r130 34 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=0.655
+ $X2=1.215 $Y2=0.74
r131 34 36 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.215 $Y=0.655
+ $X2=1.215 $Y2=0.47
r132 32 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=1.87
+ $X2=1.285 $Y2=1.87
r133 32 33 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=1.2 $Y=1.87
+ $X2=0.385 $Y2=1.87
r134 30 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=0.74
+ $X2=1.215 $Y2=0.74
r135 30 31 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.13 $Y=0.74
+ $X2=0.36 $Y2=0.74
r136 26 33 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=0.245 $Y=1.785
+ $X2=0.385 $Y2=1.87
r137 26 28 4.11587 $w=2.78e-07 $l=1e-07 $layer=LI1_cond $X=0.245 $Y=1.785
+ $X2=0.245 $Y2=1.685
r138 22 31 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.232 $Y=0.655
+ $X2=0.36 $Y2=0.74
r139 22 24 8.36086 $w=2.53e-07 $l=1.85e-07 $layer=LI1_cond $X=0.232 $Y=0.655
+ $X2=0.232 $Y2=0.47
r140 19 61 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.675 $Y=0.995
+ $X2=2.675 $Y2=1.202
r141 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.675 $Y=0.995
+ $X2=2.675 $Y2=0.56
r142 16 60 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.65 $Y=1.41
+ $X2=2.65 $Y2=1.202
r143 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.65 $Y=1.41
+ $X2=2.65 $Y2=1.985
r144 13 58 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.18 $Y=1.41
+ $X2=2.18 $Y2=1.202
r145 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.18 $Y=1.41
+ $X2=2.18 $Y2=1.985
r146 10 57 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.155 $Y=0.995
+ $X2=2.155 $Y2=1.202
r147 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.155 $Y=0.995
+ $X2=2.155 $Y2=0.56
r148 3 28 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.485 $X2=0.275 $Y2=1.685
r149 2 36 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.265 $X2=1.215 $Y2=0.47
r150 1 24 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.265 $X2=0.275 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_2%VPWR 1 2 9 11 13 17 19 24 30 34
c31 1 0 1.24896e-19 $X=1.54 $Y=1.485
r32 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r33 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r34 28 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r35 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r36 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r37 25 30 10.873 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=1.835 $Y2=2.72
r38 25 27 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r39 24 33 4.38699 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=2.825 $Y=2.72
+ $X2=3.022 $Y2=2.72
r40 24 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.825 $Y=2.72
+ $X2=2.53 $Y2=2.72
r41 19 30 10.873 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=1.6 $Y=2.72 $X2=1.835
+ $Y2=2.72
r42 19 21 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=1.6 $Y=2.72
+ $X2=0.23 $Y2=2.72
r43 17 31 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r44 17 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r45 13 16 27.0228 $w=2.88e-07 $l=6.8e-07 $layer=LI1_cond $X=2.97 $Y=1.62
+ $X2=2.97 $Y2=2.3
r46 11 33 3.05085 $w=2.9e-07 $l=1.07912e-07 $layer=LI1_cond $X=2.97 $Y=2.635
+ $X2=3.022 $Y2=2.72
r47 11 16 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=2.97 $Y=2.635
+ $X2=2.97 $Y2=2.3
r48 7 30 1.91284 $w=4.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.835 $Y=2.635
+ $X2=1.835 $Y2=2.72
r49 7 9 16.1598 $w=4.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.835 $Y=2.635
+ $X2=1.835 $Y2=2
r50 2 16 400 $w=1.7e-07 $l=8.95977e-07 $layer=licon1_PDIFF $count=1 $X=2.74
+ $Y=1.485 $X2=2.91 $Y2=2.3
r51 2 13 400 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=2.74
+ $Y=1.485 $X2=2.91 $Y2=1.62
r52 1 9 300 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=2 $X=1.54
+ $Y=1.485 $X2=1.75 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_2%X 1 2 12 14 15 16
r29 14 16 6.66644 $w=3.23e-07 $l=1.88e-07 $layer=LI1_cond $X=2.492 $Y=1.657
+ $X2=2.492 $Y2=1.845
r30 14 15 7.86522 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=2.492 $Y=1.657
+ $X2=2.492 $Y2=1.495
r31 10 12 4.91041 $w=3.43e-07 $l=1.47e-07 $layer=LI1_cond $X=2.415 $Y=0.587
+ $X2=2.562 $Y2=0.587
r32 7 12 4.404 $w=1.85e-07 $l=1.73e-07 $layer=LI1_cond $X=2.562 $Y=0.76
+ $X2=2.562 $Y2=0.587
r33 7 15 44.0639 $w=1.83e-07 $l=7.35e-07 $layer=LI1_cond $X=2.562 $Y=0.76
+ $X2=2.562 $Y2=1.495
r34 2 16 300 $w=1.7e-07 $l=4.2638e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=1.485 $X2=2.415 $Y2=1.845
r35 1 10 182 $w=1.7e-07 $l=4.37836e-07 $layer=licon1_NDIFF $count=1 $X=2.23
+ $Y=0.235 $X2=2.415 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_2%VGND 1 2 3 12 14 16 18 20 30 36 41 44 47
c51 41 0 6.13246e-20 $X=1.47 $Y=0.2
r52 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r53 43 44 13.9479 $w=5.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.735 $Y=0.2
+ $X2=2.09 $Y2=0.2
r54 39 43 2.62298 $w=5.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.61 $Y=0.2
+ $X2=1.735 $Y2=0.2
r55 39 41 9.43642 $w=5.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.61 $Y=0.2 $X2=1.47
+ $Y2=0.2
r56 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r57 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r58 34 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r59 34 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r60 33 44 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=2.09
+ $Y2=0
r61 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r62 30 46 4.38699 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=2.825 $Y=0 $X2=3.022
+ $Y2=0
r63 30 33 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.825 $Y=0 $X2=2.53
+ $Y2=0
r64 29 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r65 29 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r66 28 41 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=1.47
+ $Y2=0
r67 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r68 26 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=0.72
+ $Y2=0
r69 26 28 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=1.15
+ $Y2=0
r70 20 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.72
+ $Y2=0
r71 20 22 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.23
+ $Y2=0
r72 18 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r73 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r74 14 46 3.05085 $w=2.9e-07 $l=1.07912e-07 $layer=LI1_cond $X=2.97 $Y=0.085
+ $X2=3.022 $Y2=0
r75 14 16 12.5179 $w=2.88e-07 $l=3.15e-07 $layer=LI1_cond $X=2.97 $Y=0.085
+ $X2=2.97 $Y2=0.4
r76 10 36 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0
r77 10 12 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0.4
r78 3 16 91 $w=1.7e-07 $l=2.31571e-07 $layer=licon1_NDIFF $count=2 $X=2.75
+ $Y=0.235 $X2=2.91 $Y2=0.4
r79 2 43 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.55
+ $Y=0.265 $X2=1.735 $Y2=0.4
r80 1 12 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=0.61
+ $Y=0.265 $X2=0.745 $Y2=0.4
.ends

