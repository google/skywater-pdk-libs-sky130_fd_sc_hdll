# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__buf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__buf_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.832500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 1.075000 1.340000 1.275000 ;
    END
  END A
  PIN VGND
    ANTENNADIFFAREA  1.176500 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.980000 0.085000 ;
        RECT 0.515000  0.085000 0.895000 0.565000 ;
        RECT 1.455000  0.085000 1.835000 0.565000 ;
        RECT 2.395000  0.085000 2.775000 0.565000 ;
        RECT 3.335000  0.085000 3.715000 0.565000 ;
        RECT 4.275000  0.085000 4.655000 0.565000 ;
        RECT 5.215000  0.085000 5.595000 0.885000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.720000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.980000 2.805000 ;
        RECT 0.645000 1.835000 0.815000 2.635000 ;
        RECT 1.585000 1.835000 1.755000 2.635000 ;
        RECT 2.395000 1.835000 2.775000 2.635000 ;
        RECT 3.335000 1.835000 3.715000 2.635000 ;
        RECT 4.275000 1.835000 4.655000 2.635000 ;
        RECT 5.215000 1.485000 5.595000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  2.024500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.055000 0.255000 2.225000 0.735000 ;
        RECT 2.055000 0.735000 5.045000 0.905000 ;
        RECT 2.055000 1.445000 5.045000 1.615000 ;
        RECT 2.055000 1.615000 2.225000 2.465000 ;
        RECT 2.995000 0.255000 3.165000 0.735000 ;
        RECT 2.995000 1.615000 3.165000 2.465000 ;
        RECT 3.935000 0.255000 4.105000 0.735000 ;
        RECT 3.935000 1.615000 4.105000 2.465000 ;
        RECT 4.690000 0.905000 5.045000 1.445000 ;
        RECT 4.875000 0.255000 5.045000 0.735000 ;
        RECT 4.875000 1.615000 5.045000 2.465000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.095000 1.445000 1.745000 1.615000 ;
      RECT 0.095000 1.615000 0.425000 2.465000 ;
      RECT 0.175000 0.255000 0.345000 0.735000 ;
      RECT 0.175000 0.735000 1.745000 0.905000 ;
      RECT 0.985000 1.615000 1.365000 2.465000 ;
      RECT 1.115000 0.260000 1.285000 0.735000 ;
      RECT 1.570000 0.905000 1.745000 1.075000 ;
      RECT 1.570000 1.075000 4.495000 1.245000 ;
      RECT 1.570000 1.245000 1.745000 1.445000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__buf_8
END LIBRARY
