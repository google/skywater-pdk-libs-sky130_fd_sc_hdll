* File: sky130_fd_sc_hdll__a222oi_1.pxi.spice
* Created: Wed Sep  2 08:18:23 2020
* 
x_PM_SKY130_FD_SC_HDLL__A222OI_1%C1 N_C1_c_51_n N_C1_M1006_g N_C1_c_52_n
+ N_C1_M1011_g C1 N_C1_c_53_n C1 PM_SKY130_FD_SC_HDLL__A222OI_1%C1
x_PM_SKY130_FD_SC_HDLL__A222OI_1%C2 N_C2_c_75_n N_C2_M1002_g N_C2_c_76_n
+ N_C2_M1001_g C2 PM_SKY130_FD_SC_HDLL__A222OI_1%C2
x_PM_SKY130_FD_SC_HDLL__A222OI_1%B2 N_B2_c_100_n N_B2_M1004_g N_B2_c_101_n
+ N_B2_M1010_g B2 B2 PM_SKY130_FD_SC_HDLL__A222OI_1%B2
x_PM_SKY130_FD_SC_HDLL__A222OI_1%B1 N_B1_c_126_n N_B1_M1003_g N_B1_c_127_n
+ N_B1_M1000_g B1 B1 PM_SKY130_FD_SC_HDLL__A222OI_1%B1
x_PM_SKY130_FD_SC_HDLL__A222OI_1%A1 N_A1_c_153_n N_A1_M1005_g N_A1_c_154_n
+ N_A1_M1009_g A1 A1 PM_SKY130_FD_SC_HDLL__A222OI_1%A1
x_PM_SKY130_FD_SC_HDLL__A222OI_1%A2 N_A2_c_179_n N_A2_M1008_g N_A2_c_180_n
+ N_A2_M1007_g A2 A2 PM_SKY130_FD_SC_HDLL__A222OI_1%A2
x_PM_SKY130_FD_SC_HDLL__A222OI_1%Y N_Y_M1011_s N_Y_M1003_d N_Y_M1006_s
+ N_Y_M1001_d N_Y_c_204_n N_Y_c_209_n N_Y_c_201_n N_Y_c_223_n N_Y_c_205_n
+ N_Y_c_246_p Y Y Y N_Y_c_203_n N_Y_c_229_n PM_SKY130_FD_SC_HDLL__A222OI_1%Y
x_PM_SKY130_FD_SC_HDLL__A222OI_1%A_117_297# N_A_117_297#_M1006_d
+ N_A_117_297#_M1004_d N_A_117_297#_c_264_n N_A_117_297#_c_267_n
+ N_A_117_297#_c_263_n PM_SKY130_FD_SC_HDLL__A222OI_1%A_117_297#
x_PM_SKY130_FD_SC_HDLL__A222OI_1%A_357_297# N_A_357_297#_M1004_s
+ N_A_357_297#_M1000_d N_A_357_297#_M1007_d N_A_357_297#_c_286_n
+ N_A_357_297#_c_293_n N_A_357_297#_c_288_n N_A_357_297#_c_285_n
+ PM_SKY130_FD_SC_HDLL__A222OI_1%A_357_297#
x_PM_SKY130_FD_SC_HDLL__A222OI_1%VPWR N_VPWR_M1009_d N_VPWR_c_318_n
+ N_VPWR_c_319_n N_VPWR_c_320_n VPWR N_VPWR_c_321_n N_VPWR_c_317_n
+ PM_SKY130_FD_SC_HDLL__A222OI_1%VPWR
x_PM_SKY130_FD_SC_HDLL__A222OI_1%VGND N_VGND_M1002_d N_VGND_M1008_d
+ N_VGND_c_360_n N_VGND_c_361_n VGND N_VGND_c_362_n N_VGND_c_363_n
+ N_VGND_c_364_n N_VGND_c_365_n VGND PM_SKY130_FD_SC_HDLL__A222OI_1%VGND
cc_1 VNB N_C1_c_51_n 0.0360048f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_C1_c_52_n 0.0228156f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1
cc_3 VNB N_C1_c_53_n 0.0143108f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.165
cc_4 VNB N_C2_c_75_n 0.019489f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_C2_c_76_n 0.0264956f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1
cc_6 VNB C2 0.0056473f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=1.09
cc_7 VNB N_B2_c_100_n 0.0286409f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_8 VNB N_B2_c_101_n 0.02033f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1
cc_9 VNB B2 0.00502952f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.157
cc_10 VNB N_B1_c_126_n 0.0176754f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_11 VNB N_B1_c_127_n 0.0191979f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1
cc_12 VNB B1 0.00413574f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=1.09
cc_13 VNB N_A1_c_153_n 0.0193283f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_14 VNB N_A1_c_154_n 0.0259719f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1
cc_15 VNB A1 0.00479701f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.157
cc_16 VNB N_A2_c_179_n 0.0231274f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_17 VNB N_A2_c_180_n 0.0263717f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1
cc_18 VNB A2 0.0177156f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=1.09
cc_19 VNB N_Y_c_201_n 0.00745159f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB Y 0.0111672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_203_n 0.0153416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_317_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_360_n 0.0139533f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=1.09
cc_24 VNB N_VGND_c_361_n 0.00282211f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.165
cc_25 VNB N_VGND_c_362_n 0.049783f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_363_n 0.0252541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_364_n 0.0190776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_365_n 0.221894f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_C1_c_51_n 0.0384802f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_30 VPB N_C1_c_53_n 8.73116e-19 $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.165
cc_31 VPB N_C2_c_76_n 0.0302038f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1
cc_32 VPB C2 0.00151749f $X=-0.19 $Y=1.305 $X2=0.155 $Y2=1.09
cc_33 VPB N_B2_c_100_n 0.0313001f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_34 VPB B2 3.97067e-19 $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.157
cc_35 VPB N_B1_c_127_n 0.025175f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1
cc_36 VPB B1 6.68054e-19 $X=-0.19 $Y=1.305 $X2=0.155 $Y2=1.09
cc_37 VPB N_A1_c_154_n 0.0265429f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1
cc_38 VPB A1 0.00103719f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.157
cc_39 VPB N_A2_c_180_n 0.0341616f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1
cc_40 VPB A2 0.00294803f $X=-0.19 $Y=1.305 $X2=0.155 $Y2=1.09
cc_41 VPB N_Y_c_204_n 0.012089f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.157
cc_42 VPB N_Y_c_205_n 0.0337035f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB Y 0.00571367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_117_297#_c_263_n 0.0153507f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.157
cc_45 VPB N_A_357_297#_c_285_n 0.0314516f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_318_n 0.00286f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.555
cc_47 VPB N_VPWR_c_319_n 0.0800165f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.165
cc_48 VPB N_VPWR_c_320_n 0.00513801f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.165
cc_49 VPB N_VPWR_c_321_n 0.0213946f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_317_n 0.0494832f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 N_C1_c_52_n N_C2_c_75_n 0.0390402f $X=0.52 $Y=1 $X2=-0.19 $Y2=-0.24
cc_52 N_C1_c_51_n N_C2_c_76_n 0.0810787f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_53 N_C1_c_53_n N_C2_c_76_n 3.59027e-19 $X=0.38 $Y=1.165 $X2=0 $Y2=0
cc_54 N_C1_c_51_n C2 0.00109125f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_55 N_C1_c_53_n C2 0.0265461f $X=0.38 $Y=1.165 $X2=0 $Y2=0
cc_56 N_C1_c_51_n N_Y_c_204_n 0.0210637f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_57 N_C1_c_53_n N_Y_c_204_n 0.0160037f $X=0.38 $Y=1.165 $X2=0 $Y2=0
cc_58 N_C1_c_52_n N_Y_c_209_n 0.00944548f $X=0.52 $Y=1 $X2=0 $Y2=0
cc_59 N_C1_c_53_n N_Y_c_209_n 0.0106373f $X=0.38 $Y=1.165 $X2=0 $Y2=0
cc_60 N_C1_c_51_n N_Y_c_201_n 0.00731804f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_61 N_C1_c_53_n N_Y_c_201_n 0.0236446f $X=0.38 $Y=1.165 $X2=0 $Y2=0
cc_62 N_C1_c_51_n N_Y_c_205_n 0.00569277f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_63 N_C1_c_53_n N_Y_c_205_n 0.0206893f $X=0.38 $Y=1.165 $X2=0 $Y2=0
cc_64 N_C1_c_51_n N_A_117_297#_c_264_n 0.0114255f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_65 N_C1_c_51_n N_VPWR_c_319_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_66 N_C1_c_51_n N_VPWR_c_317_n 0.0129911f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_67 N_C1_c_52_n N_VGND_c_363_n 0.00426565f $X=0.52 $Y=1 $X2=0 $Y2=0
cc_68 N_C1_c_52_n N_VGND_c_364_n 0.00188599f $X=0.52 $Y=1 $X2=0 $Y2=0
cc_69 N_C1_c_52_n N_VGND_c_365_n 0.00672235f $X=0.52 $Y=1 $X2=0 $Y2=0
cc_70 N_C2_c_76_n N_Y_c_204_n 0.0185743f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_71 C2 N_Y_c_204_n 0.0317688f $X=0.87 $Y=1.09 $X2=0 $Y2=0
cc_72 N_C2_c_75_n N_Y_c_209_n 0.0132688f $X=0.88 $Y=1 $X2=0 $Y2=0
cc_73 N_C2_c_76_n N_Y_c_209_n 0.00404123f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_74 C2 N_Y_c_209_n 0.0293396f $X=0.87 $Y=1.09 $X2=0 $Y2=0
cc_75 N_C2_c_75_n Y 0.00491079f $X=0.88 $Y=1 $X2=0 $Y2=0
cc_76 N_C2_c_76_n Y 0.00696213f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_77 C2 Y 0.0263586f $X=0.87 $Y=1.09 $X2=0 $Y2=0
cc_78 N_C2_c_76_n N_A_117_297#_c_264_n 0.012355f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_79 N_C2_c_76_n N_A_117_297#_c_263_n 0.012437f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_80 N_C2_c_76_n N_VPWR_c_319_n 0.00430943f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_81 N_C2_c_76_n N_VPWR_c_317_n 0.00741278f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_82 N_C2_c_75_n N_VGND_c_363_n 0.00340533f $X=0.88 $Y=1 $X2=0 $Y2=0
cc_83 N_C2_c_75_n N_VGND_c_364_n 0.0108923f $X=0.88 $Y=1 $X2=0 $Y2=0
cc_84 N_C2_c_75_n N_VGND_c_365_n 0.00385622f $X=0.88 $Y=1 $X2=0 $Y2=0
cc_85 N_B2_c_101_n N_B1_c_126_n 0.0390286f $X=2.17 $Y=1 $X2=-0.19 $Y2=-0.24
cc_86 N_B2_c_100_n N_B1_c_127_n 0.0810268f $X=2.145 $Y=1.41 $X2=0 $Y2=0
cc_87 B2 N_B1_c_127_n 3.78404e-19 $X=2.075 $Y=1.175 $X2=0 $Y2=0
cc_88 N_B2_c_100_n B1 0.0010697f $X=2.145 $Y=1.41 $X2=0 $Y2=0
cc_89 B2 B1 0.0263163f $X=2.075 $Y=1.175 $X2=0 $Y2=0
cc_90 N_B2_c_100_n N_Y_c_223_n 0.00469679f $X=2.145 $Y=1.41 $X2=0 $Y2=0
cc_91 N_B2_c_101_n N_Y_c_223_n 0.0130513f $X=2.17 $Y=1 $X2=0 $Y2=0
cc_92 B2 N_Y_c_223_n 0.0225913f $X=2.075 $Y=1.175 $X2=0 $Y2=0
cc_93 N_B2_c_100_n Y 0.00670956f $X=2.145 $Y=1.41 $X2=0 $Y2=0
cc_94 N_B2_c_101_n Y 0.00496145f $X=2.17 $Y=1 $X2=0 $Y2=0
cc_95 B2 Y 0.0204653f $X=2.075 $Y=1.175 $X2=0 $Y2=0
cc_96 N_B2_c_100_n N_A_117_297#_c_267_n 0.0102103f $X=2.145 $Y=1.41 $X2=0 $Y2=0
cc_97 N_B2_c_100_n N_A_117_297#_c_263_n 0.00956552f $X=2.145 $Y=1.41 $X2=0 $Y2=0
cc_98 N_B2_c_100_n N_A_357_297#_c_286_n 0.019582f $X=2.145 $Y=1.41 $X2=0 $Y2=0
cc_99 B2 N_A_357_297#_c_286_n 0.0247563f $X=2.075 $Y=1.175 $X2=0 $Y2=0
cc_100 N_B2_c_100_n N_A_357_297#_c_288_n 0.00135714f $X=2.145 $Y=1.41 $X2=0
+ $Y2=0
cc_101 N_B2_c_100_n N_VPWR_c_319_n 0.00429453f $X=2.145 $Y=1.41 $X2=0 $Y2=0
cc_102 N_B2_c_100_n N_VPWR_c_317_n 0.00742188f $X=2.145 $Y=1.41 $X2=0 $Y2=0
cc_103 N_B2_c_101_n N_VGND_c_362_n 0.00426565f $X=2.17 $Y=1 $X2=0 $Y2=0
cc_104 N_B2_c_101_n N_VGND_c_364_n 0.0100257f $X=2.17 $Y=1 $X2=0 $Y2=0
cc_105 N_B2_c_101_n N_VGND_c_365_n 0.00714369f $X=2.17 $Y=1 $X2=0 $Y2=0
cc_106 N_B1_c_126_n N_A1_c_153_n 0.019471f $X=2.53 $Y=1 $X2=-0.19 $Y2=-0.24
cc_107 N_B1_c_127_n N_A1_c_154_n 0.0422953f $X=2.615 $Y=1.41 $X2=0 $Y2=0
cc_108 B1 N_A1_c_154_n 3.58154e-19 $X=2.47 $Y=1.09 $X2=0 $Y2=0
cc_109 N_B1_c_127_n A1 0.00115665f $X=2.615 $Y=1.41 $X2=0 $Y2=0
cc_110 B1 A1 0.0265603f $X=2.47 $Y=1.09 $X2=0 $Y2=0
cc_111 N_B1_c_126_n N_Y_c_229_n 0.0195444f $X=2.53 $Y=1 $X2=0 $Y2=0
cc_112 N_B1_c_127_n N_Y_c_229_n 0.00320504f $X=2.615 $Y=1.41 $X2=0 $Y2=0
cc_113 B1 N_Y_c_229_n 0.0200574f $X=2.47 $Y=1.09 $X2=0 $Y2=0
cc_114 N_B1_c_127_n N_A_357_297#_c_286_n 0.0201794f $X=2.615 $Y=1.41 $X2=0 $Y2=0
cc_115 B1 N_A_357_297#_c_286_n 0.0183872f $X=2.47 $Y=1.09 $X2=0 $Y2=0
cc_116 N_B1_c_127_n N_A_357_297#_c_288_n 0.00823554f $X=2.615 $Y=1.41 $X2=0
+ $Y2=0
cc_117 B1 N_A_357_297#_c_288_n 0.00268539f $X=2.47 $Y=1.09 $X2=0 $Y2=0
cc_118 N_B1_c_127_n N_VPWR_c_318_n 0.00215136f $X=2.615 $Y=1.41 $X2=0 $Y2=0
cc_119 N_B1_c_127_n N_VPWR_c_319_n 0.00678802f $X=2.615 $Y=1.41 $X2=0 $Y2=0
cc_120 N_B1_c_127_n N_VPWR_c_317_n 0.0120649f $X=2.615 $Y=1.41 $X2=0 $Y2=0
cc_121 N_B1_c_126_n N_VGND_c_362_n 0.00365909f $X=2.53 $Y=1 $X2=0 $Y2=0
cc_122 N_B1_c_126_n N_VGND_c_365_n 0.00542828f $X=2.53 $Y=1 $X2=0 $Y2=0
cc_123 N_A1_c_153_n N_A2_c_179_n 0.0281396f $X=3.06 $Y=1 $X2=-0.19 $Y2=-0.24
cc_124 N_A1_c_154_n N_A2_c_180_n 0.0529493f $X=3.085 $Y=1.41 $X2=0 $Y2=0
cc_125 A1 N_A2_c_180_n 3.77261e-19 $X=3.065 $Y=1.175 $X2=0 $Y2=0
cc_126 N_A1_c_154_n A2 0.00116718f $X=3.085 $Y=1.41 $X2=0 $Y2=0
cc_127 A1 A2 0.0275585f $X=3.065 $Y=1.175 $X2=0 $Y2=0
cc_128 A1 N_Y_c_229_n 0.00364837f $X=3.065 $Y=1.175 $X2=0 $Y2=0
cc_129 N_A1_c_154_n N_A_357_297#_c_293_n 0.0198757f $X=3.085 $Y=1.41 $X2=0 $Y2=0
cc_130 A1 N_A_357_297#_c_293_n 0.0232476f $X=3.065 $Y=1.175 $X2=0 $Y2=0
cc_131 N_A1_c_154_n N_A_357_297#_c_288_n 0.00298027f $X=3.085 $Y=1.41 $X2=0
+ $Y2=0
cc_132 A1 N_A_357_297#_c_288_n 0.00260072f $X=3.065 $Y=1.175 $X2=0 $Y2=0
cc_133 N_A1_c_154_n N_VPWR_c_318_n 0.0134039f $X=3.085 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A1_c_154_n N_VPWR_c_319_n 0.00622633f $X=3.085 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A1_c_154_n N_VPWR_c_317_n 0.0105052f $X=3.085 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A1_c_153_n N_VGND_c_361_n 0.00324506f $X=3.06 $Y=1 $X2=0 $Y2=0
cc_137 N_A1_c_153_n N_VGND_c_362_n 0.00585385f $X=3.06 $Y=1 $X2=0 $Y2=0
cc_138 N_A1_c_153_n N_VGND_c_365_n 0.0112939f $X=3.06 $Y=1 $X2=0 $Y2=0
cc_139 N_A2_c_180_n N_A_357_297#_c_293_n 0.0178854f $X=3.615 $Y=1.41 $X2=0 $Y2=0
cc_140 A2 N_A_357_297#_c_293_n 0.0174219f $X=3.795 $Y=1.07 $X2=0 $Y2=0
cc_141 N_A2_c_180_n N_A_357_297#_c_285_n 0.00730782f $X=3.615 $Y=1.41 $X2=0
+ $Y2=0
cc_142 A2 N_A_357_297#_c_285_n 0.0196866f $X=3.795 $Y=1.07 $X2=0 $Y2=0
cc_143 N_A2_c_180_n N_VPWR_c_318_n 0.00624759f $X=3.615 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A2_c_180_n N_VPWR_c_321_n 0.00702461f $X=3.615 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A2_c_180_n N_VPWR_c_317_n 0.0137565f $X=3.615 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A2_c_179_n N_VGND_c_361_n 0.0240859f $X=3.59 $Y=1 $X2=0 $Y2=0
cc_147 N_A2_c_180_n N_VGND_c_361_n 0.00391379f $X=3.615 $Y=1.41 $X2=0 $Y2=0
cc_148 A2 N_VGND_c_361_n 0.0293508f $X=3.795 $Y=1.07 $X2=0 $Y2=0
cc_149 N_A2_c_179_n N_VGND_c_362_n 0.00154325f $X=3.59 $Y=1 $X2=0 $Y2=0
cc_150 N_A2_c_179_n N_VGND_c_365_n 0.00348588f $X=3.59 $Y=1 $X2=0 $Y2=0
cc_151 N_Y_c_204_n N_A_117_297#_M1006_d 0.00531836f $X=1.405 $Y=1.64 $X2=-0.19
+ $Y2=-0.24
cc_152 N_Y_c_204_n N_A_117_297#_c_264_n 0.0125417f $X=1.405 $Y=1.64 $X2=0 $Y2=0
cc_153 N_Y_c_205_n N_A_117_297#_c_264_n 0.0149584f $X=0.26 $Y=1.765 $X2=0 $Y2=0
cc_154 N_Y_M1001_d N_A_117_297#_c_263_n 0.00668468f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_155 N_Y_c_204_n N_A_117_297#_c_263_n 0.0248992f $X=1.405 $Y=1.64 $X2=0 $Y2=0
cc_156 N_Y_c_204_n N_A_357_297#_c_286_n 0.0270266f $X=1.405 $Y=1.64 $X2=0 $Y2=0
cc_157 N_Y_c_205_n N_VPWR_c_319_n 0.00827745f $X=0.26 $Y=1.765 $X2=0 $Y2=0
cc_158 N_Y_M1006_s N_VPWR_c_317_n 0.00450527f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_159 N_Y_M1001_d N_VPWR_c_317_n 0.00218346f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_160 N_Y_c_205_n N_VPWR_c_317_n 0.00865511f $X=0.26 $Y=1.765 $X2=0 $Y2=0
cc_161 N_Y_c_209_n A_119_47# 0.0036173f $X=1.405 $Y=0.73 $X2=-0.19 $Y2=-0.24
cc_162 N_Y_c_209_n N_VGND_M1002_d 0.012203f $X=1.405 $Y=0.73 $X2=-0.19 $Y2=-0.24
cc_163 N_Y_c_223_n N_VGND_M1002_d 0.0188648f $X=2.41 $Y=0.73 $X2=-0.19 $Y2=-0.24
cc_164 N_Y_c_246_p N_VGND_M1002_d 0.00508744f $X=1.53 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_165 Y N_VGND_M1002_d 0.0026233f $X=1.405 $Y=1.09 $X2=-0.19 $Y2=-0.24
cc_166 N_Y_c_223_n N_VGND_c_362_n 0.0109357f $X=2.41 $Y=0.73 $X2=0 $Y2=0
cc_167 N_Y_c_229_n N_VGND_c_362_n 0.0267539f $X=2.81 $Y=0.38 $X2=0 $Y2=0
cc_168 N_Y_c_209_n N_VGND_c_363_n 0.00722221f $X=1.405 $Y=0.73 $X2=0 $Y2=0
cc_169 N_Y_c_203_n N_VGND_c_363_n 0.0215737f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_170 N_Y_c_209_n N_VGND_c_364_n 0.0304018f $X=1.405 $Y=0.73 $X2=0 $Y2=0
cc_171 N_Y_c_223_n N_VGND_c_364_n 0.00358825f $X=2.41 $Y=0.73 $X2=0 $Y2=0
cc_172 N_Y_c_246_p N_VGND_c_364_n 0.0199692f $X=1.53 $Y=0.73 $X2=0 $Y2=0
cc_173 N_Y_M1011_s N_VGND_c_365_n 0.00256712f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_174 N_Y_M1003_d N_VGND_c_365_n 0.00342247f $X=2.605 $Y=0.235 $X2=0 $Y2=0
cc_175 N_Y_c_209_n N_VGND_c_365_n 0.0147863f $X=1.405 $Y=0.73 $X2=0 $Y2=0
cc_176 N_Y_c_223_n N_VGND_c_365_n 0.0192858f $X=2.41 $Y=0.73 $X2=0 $Y2=0
cc_177 N_Y_c_246_p N_VGND_c_365_n 0.00127592f $X=1.53 $Y=0.73 $X2=0 $Y2=0
cc_178 N_Y_c_203_n N_VGND_c_365_n 0.0125683f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_179 N_Y_c_229_n N_VGND_c_365_n 0.0203845f $X=2.81 $Y=0.38 $X2=0 $Y2=0
cc_180 N_Y_c_223_n A_449_47# 0.00535658f $X=2.41 $Y=0.73 $X2=-0.19 $Y2=-0.24
cc_181 N_A_117_297#_c_263_n N_A_357_297#_M1004_s 0.00736972f $X=2.17 $Y=2.3
+ $X2=-0.19 $Y2=1.305
cc_182 N_A_117_297#_M1004_d N_A_357_297#_c_286_n 0.00809642f $X=2.235 $Y=1.485
+ $X2=0 $Y2=0
cc_183 N_A_117_297#_c_267_n N_A_357_297#_c_286_n 0.0120622f $X=2.38 $Y=2.3 $X2=0
+ $Y2=0
cc_184 N_A_117_297#_c_263_n N_A_357_297#_c_286_n 0.00988445f $X=2.17 $Y=2.3
+ $X2=0 $Y2=0
cc_185 N_A_117_297#_c_267_n N_A_357_297#_c_288_n 0.00707935f $X=2.38 $Y=2.3
+ $X2=0 $Y2=0
cc_186 N_A_117_297#_c_264_n N_VPWR_c_319_n 0.0184162f $X=0.73 $Y=2.3 $X2=0 $Y2=0
cc_187 N_A_117_297#_c_263_n N_VPWR_c_319_n 0.0951894f $X=2.17 $Y=2.3 $X2=0 $Y2=0
cc_188 N_A_117_297#_M1006_d N_VPWR_c_317_n 0.00231261f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_189 N_A_117_297#_M1004_d N_VPWR_c_317_n 0.00436106f $X=2.235 $Y=1.485 $X2=0
+ $Y2=0
cc_190 N_A_117_297#_c_264_n N_VPWR_c_317_n 0.0121547f $X=0.73 $Y=2.3 $X2=0 $Y2=0
cc_191 N_A_117_297#_c_263_n N_VPWR_c_317_n 0.0570174f $X=2.17 $Y=2.3 $X2=0 $Y2=0
cc_192 N_A_357_297#_c_293_n N_VPWR_M1009_d 0.00961877f $X=3.765 $Y=1.617
+ $X2=-0.19 $Y2=1.305
cc_193 N_A_357_297#_c_293_n N_VPWR_c_318_n 0.0210667f $X=3.765 $Y=1.617 $X2=0
+ $Y2=0
cc_194 N_A_357_297#_c_288_n N_VPWR_c_318_n 0.0215026f $X=2.85 $Y=1.665 $X2=0
+ $Y2=0
cc_195 N_A_357_297#_c_288_n N_VPWR_c_319_n 0.0063902f $X=2.85 $Y=1.665 $X2=0
+ $Y2=0
cc_196 N_A_357_297#_c_285_n N_VPWR_c_321_n 0.00753114f $X=3.85 $Y=1.665 $X2=0
+ $Y2=0
cc_197 N_A_357_297#_M1004_s N_VPWR_c_317_n 0.00218346f $X=1.785 $Y=1.485 $X2=0
+ $Y2=0
cc_198 N_A_357_297#_M1000_d N_VPWR_c_317_n 0.00478011f $X=2.705 $Y=1.485 $X2=0
+ $Y2=0
cc_199 N_A_357_297#_M1007_d N_VPWR_c_317_n 0.00460549f $X=3.705 $Y=1.485 $X2=0
+ $Y2=0
cc_200 N_A_357_297#_c_288_n N_VPWR_c_317_n 0.00830125f $X=2.85 $Y=1.665 $X2=0
+ $Y2=0
cc_201 N_A_357_297#_c_285_n N_VPWR_c_317_n 0.00873505f $X=3.85 $Y=1.665 $X2=0
+ $Y2=0
cc_202 A_119_47# N_VGND_c_365_n 0.00248276f $X=0.595 $Y=0.235 $X2=0.26 $Y2=0.51
cc_203 N_VGND_c_365_n A_449_47# 0.00230787f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_204 N_VGND_c_365_n A_627_47# 0.016267f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
