* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nor4bb_1 A B C_N D_N VGND VNB VPB VPWR Y
X0 Y a_216_93# a_422_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 Y a_27_410# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_422_297# a_27_410# a_518_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 VGND a_216_93# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND D_N a_216_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_622_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_518_297# B a_622_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_27_410# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X10 VPWR D_N a_216_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X11 a_27_410# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
