* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nor4bb_1 A B C_N D_N VGND VNB VPB VPWR Y
M1000 VGND C_N a_27_410# VNB nshort w=420000u l=150000u
+  ad=7.674e+11p pd=7.31e+06u as=1.302e+11p ps=1.46e+06u
M1001 Y B VGND VNB nshort w=650000u l=150000u
+  ad=3.9e+11p pd=3.8e+06u as=0p ps=0u
M1002 a_216_93# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.281e+11p pd=1.45e+06u as=0p ps=0u
M1003 Y a_216_93# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_422_297# a_216_93# Y VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=2.7e+11p ps=2.54e+06u
M1006 VGND a_27_410# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_622_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.23625e+11p pd=5.22e+06u as=2.9e+11p ps=2.58e+06u
M1008 VPWR C_N a_27_410# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1009 a_216_93# D_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1010 a_622_297# B a_518_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.4e+11p ps=2.68e+06u
M1011 a_518_297# a_27_410# a_422_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
