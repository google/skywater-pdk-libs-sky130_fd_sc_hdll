* File: sky130_fd_sc_hdll__a211oi_4.spice
* Created: Thu Aug 27 18:51:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a211oi_4.pex.spice"
.subckt sky130_fd_sc_hdll__a211oi_4  VNB VPB A2 A1 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A2_M1003_g N_A_119_47#_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75007.4 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A2_M1011_g N_A_119_47#_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75006.9 A=0.0975 P=1.6 MULT=1
MM1020 N_VGND_M1011_d N_A2_M1020_g N_A_119_47#_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75006.4 A=0.0975 P=1.6 MULT=1
MM1012 N_A_119_47#_M1020_s N_A1_M1012_g N_Y_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.6
+ SB=75006 A=0.0975 P=1.6 MULT=1
MM1025 N_A_119_47#_M1025_d N_A1_M1025_g N_Y_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75005.5 A=0.0975 P=1.6 MULT=1
MM1028 N_A_119_47#_M1025_d N_A1_M1028_g N_Y_M1028_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.5
+ SB=75005.1 A=0.0975 P=1.6 MULT=1
MM1030 N_A_119_47#_M1030_d N_A1_M1030_g N_Y_M1028_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.1
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1031 N_VGND_M1031_d N_A2_M1031_g N_A_119_47#_M1030_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.5
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1031_d N_B1_M1005_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.141375 PD=0.92 PS=1.085 NRD=0 NRS=11.988 M=1 R=4.33333
+ SA=75003.9 SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_B1_M1008_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.141375 PD=0.98 PS=1.085 NRD=0 NRS=16.608 M=1 R=4.33333
+ SA=75004.5 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1008_d N_B1_M1021_g N_Y_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.105625 PD=0.98 PS=0.975 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75005
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_C1_M1001_g N_Y_M1021_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.105625 PD=0.97 PS=0.975 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75005.5
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1001_d N_C1_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75006 SB=75001.6
+ A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_C1_M1013_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75006.4 SB=75001.2
+ A=0.0975 P=1.6 MULT=1
MM1022 N_VGND_M1013_d N_C1_M1022_g N_Y_M1022_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.10725 PD=0.97 PS=0.98 NRD=8.304 NRS=0.912 M=1 R=4.33333 SA=75006.9
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1024 N_VGND_M1024_d N_B1_M1024_g N_Y_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1885 AS=0.10725 PD=1.88 PS=0.98 NRD=0.912 NRS=8.304 M=1 R=4.33333
+ SA=75007.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM16_noxref N_VPWR_M16_noxref_d N_A2_M16_noxref_g N_noxref_7_M16_noxref_s VPB
+ PHIGHVT L=0.18 W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.2 SB=90007.3 A=0.18 P=2.36 MULT=1
MM17_noxref N_noxref_7_M17_noxref_d N_A2_M17_noxref_g N_VPWR_M16_noxref_d VPB
+ PHIGHVT L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.6 SB=90006.9 A=0.18 P=2.36 MULT=1
MM18_noxref N_VPWR_M18_noxref_d N_A2_M18_noxref_g N_noxref_7_M17_noxref_d VPB
+ PHIGHVT L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001.1 SB=90006.4 A=0.18 P=2.36 MULT=1
MM19_noxref N_noxref_7_M19_noxref_d N_A1_M19_noxref_g N_VPWR_M18_noxref_d VPB
+ PHIGHVT L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001.6 SB=90005.9 A=0.18 P=2.36 MULT=1
MM20_noxref N_VPWR_M20_noxref_d N_A1_M20_noxref_g N_noxref_7_M19_noxref_d VPB
+ PHIGHVT L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90002.1 SB=90005.5 A=0.18 P=2.36 MULT=1
MM21_noxref N_noxref_7_M21_noxref_d N_A1_M21_noxref_g N_VPWR_M20_noxref_d VPB
+ PHIGHVT L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90002.5 SB=90005 A=0.18 P=2.36 MULT=1
MM22_noxref N_VPWR_M22_noxref_d N_A1_M22_noxref_g N_noxref_7_M21_noxref_d VPB
+ PHIGHVT L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90003 SB=90004.5 A=0.18 P=2.36 MULT=1
MM23_noxref N_noxref_7_M23_noxref_d N_A2_M23_noxref_g N_VPWR_M22_noxref_d VPB
+ PHIGHVT L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90003.5 SB=90004.1 A=0.18 P=2.36 MULT=1
MM24_noxref N_noxref_9_M24_noxref_d N_B1_M24_noxref_g N_noxref_7_M23_noxref_d
+ VPB PHIGHVT L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653
+ M=1 R=5.55556 SA=90003.9 SB=90003.6 A=0.18 P=2.36 MULT=1
MM25_noxref N_noxref_7_M25_noxref_d N_B1_M25_noxref_g N_noxref_9_M24_noxref_d
+ VPB PHIGHVT L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653
+ M=1 R=5.55556 SA=90004.4 SB=90003.1 A=0.18 P=2.36 MULT=1
MM26_noxref noxref_10 N_B1_M26_noxref_g N_noxref_7_M25_noxref_d VPB PHIGHVT
+ L=0.18 W=1 AD=0.16 AS=0.145 PD=1.32 PS=1.29 NRD=20.6653 NRS=0.9653 M=1
+ R=5.55556 SA=90004.9 SB=90002.6 A=0.18 P=2.36 MULT=1
MM27_noxref N_Y_M27_noxref_d N_C1_M27_noxref_g noxref_10 VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.16 PD=1.3 PS=1.32 NRD=1.9503 NRS=20.6653 M=1 R=5.55556 SA=90005.4
+ SB=90002.1 A=0.18 P=2.36 MULT=1
MM28_noxref N_noxref_9_M28_noxref_d N_C1_M28_noxref_g N_Y_M27_noxref_d VPB
+ PHIGHVT L=0.18 W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1
+ R=5.55556 SA=90005.9 SB=90001.7 A=0.18 P=2.36 MULT=1
MM29_noxref N_Y_M29_noxref_d N_C1_M29_noxref_g N_noxref_9_M28_noxref_d VPB
+ PHIGHVT L=0.18 W=1 AD=0.16 AS=0.15 PD=1.32 PS=1.3 NRD=5.8903 NRS=1.9503 M=1
+ R=5.55556 SA=90006.3 SB=90001.2 A=0.18 P=2.36 MULT=1
MM30_noxref noxref_12 N_C1_M30_noxref_g N_Y_M29_noxref_d VPB PHIGHVT L=0.18 W=1
+ AD=0.165 AS=0.16 PD=1.33 PS=1.32 NRD=21.6503 NRS=1.9503 M=1 R=5.55556
+ SA=90006.8 SB=90000.7 A=0.18 P=2.36 MULT=1
MM31_noxref N_noxref_7_M31_noxref_d N_B1_M31_noxref_g noxref_12 VPB PHIGHVT
+ L=0.18 W=1 AD=0.27 AS=0.165 PD=2.54 PS=1.33 NRD=0.9653 NRS=21.6503 M=1
+ R=5.55556 SA=90007.3 SB=90000.2 A=0.18 P=2.36 MULT=1
DX32_noxref VNB VPB NWDIODE A=13.8993 P=20.53
pX33_noxref noxref_15 Y Y PROBETYPE=1
*
.include "sky130_fd_sc_hdll__a211oi_4.pxi.spice"
*
.ends
*
*
