* File: sky130_fd_sc_hdll__a211oi_4.spice
* Created: Wed Sep  2 08:16:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a211oi_4.pex.spice"
.subckt sky130_fd_sc_hdll__a211oi_4  VNB VPB A2 A1 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A2_M1003_g N_A_119_47#_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75007.4 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A2_M1011_g N_A_119_47#_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75006.9 A=0.0975 P=1.6 MULT=1
MM1020 N_VGND_M1011_d N_A2_M1020_g N_A_119_47#_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75006.4 A=0.0975 P=1.6 MULT=1
MM1012 N_A_119_47#_M1020_s N_A1_M1012_g N_Y_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.6
+ SB=75006 A=0.0975 P=1.6 MULT=1
MM1025 N_A_119_47#_M1025_d N_A1_M1025_g N_Y_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75005.5 A=0.0975 P=1.6 MULT=1
MM1028 N_A_119_47#_M1025_d N_A1_M1028_g N_Y_M1028_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.5
+ SB=75005.1 A=0.0975 P=1.6 MULT=1
MM1030 N_A_119_47#_M1030_d N_A1_M1030_g N_Y_M1028_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.1
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1031 N_VGND_M1031_d N_A2_M1031_g N_A_119_47#_M1030_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.5
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1031_d N_B1_M1005_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.141375 PD=0.92 PS=1.085 NRD=0 NRS=11.988 M=1 R=4.33333
+ SA=75003.9 SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_B1_M1008_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.141375 PD=0.98 PS=1.085 NRD=0 NRS=16.608 M=1 R=4.33333
+ SA=75004.5 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1008_d N_B1_M1021_g N_Y_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.105625 PD=0.98 PS=0.975 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75005
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_C1_M1001_g N_Y_M1021_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.105625 PD=0.97 PS=0.975 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75005.5
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1001_d N_C1_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75006 SB=75001.6
+ A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_C1_M1013_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75006.4 SB=75001.2
+ A=0.0975 P=1.6 MULT=1
MM1022 N_VGND_M1013_d N_C1_M1022_g N_Y_M1022_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.10725 PD=0.97 PS=0.98 NRD=8.304 NRS=0.912 M=1 R=4.33333 SA=75006.9
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1024 N_VGND_M1024_d N_B1_M1024_g N_Y_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1885 AS=0.10725 PD=1.88 PS=0.98 NRD=0.912 NRS=8.304 M=1 R=4.33333
+ SA=75007.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_A_27_297#_M1000_d N_A2_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90007.3 A=0.18 P=2.36 MULT=1
MM1002 N_A_27_297#_M1002_d N_A2_M1002_g N_VPWR_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90006.9 A=0.18 P=2.36 MULT=1
MM1014 N_A_27_297#_M1002_d N_A2_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90006.4 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1014_s N_A1_M1007_g N_A_27_297#_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90005.9 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1010_d N_A1_M1010_g N_A_27_297#_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90005.5 A=0.18 P=2.36 MULT=1
MM1016 N_VPWR_M1010_d N_A1_M1016_g N_A_27_297#_M1016_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90005 A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1018_d N_A1_M1018_g N_A_27_297#_M1016_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90004.5 A=0.18 P=2.36 MULT=1
MM1029 N_A_27_297#_M1029_d N_A2_M1029_g N_VPWR_M1018_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90004.1 A=0.18 P=2.36 MULT=1
MM1017 N_A_27_297#_M1029_d N_B1_M1017_g N_A_869_297#_M1017_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.9 SB=90003.6 A=0.18 P=2.36 MULT=1
MM1023 N_A_27_297#_M1023_d N_B1_M1023_g N_A_869_297#_M1017_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.4 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1009 N_A_27_297#_M1023_d N_B1_M1009_g A_1057_297# VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.16 PD=1.29 PS=1.32 NRD=0.9653 NRS=20.6653 M=1 R=5.55556
+ SA=90004.9 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1015 A_1057_297# N_C1_M1015_g N_Y_M1015_s VPB PHIGHVT L=0.18 W=1 AD=0.16
+ AS=0.15 PD=1.32 PS=1.3 NRD=20.6653 NRS=1.9503 M=1 R=5.55556 SA=90005.4
+ SB=90002.1 A=0.18 P=2.36 MULT=1
MM1006 N_A_869_297#_M1006_d N_C1_M1006_g N_Y_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90005.9
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1019 N_A_869_297#_M1006_d N_C1_M1019_g N_Y_M1019_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.16 PD=1.3 PS=1.32 NRD=1.9503 NRS=5.8903 M=1 R=5.55556 SA=90006.3
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1026 A_1449_297# N_C1_M1026_g N_Y_M1019_s VPB PHIGHVT L=0.18 W=1 AD=0.165
+ AS=0.16 PD=1.33 PS=1.32 NRD=21.6503 NRS=1.9503 M=1 R=5.55556 SA=90006.8
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1027 N_A_27_297#_M1027_d N_B1_M1027_g A_1449_297# VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.165 PD=2.54 PS=1.33 NRD=0.9653 NRS=21.6503 M=1 R=5.55556
+ SA=90007.3 SB=90000.2 A=0.18 P=2.36 MULT=1
DX32_noxref VNB VPB NWDIODE A=13.8993 P=20.53
pX33_noxref noxref_15 Y Y PROBETYPE=1
*
.include "sky130_fd_sc_hdll__a211oi_4.pxi.spice"
*
.ends
*
*
