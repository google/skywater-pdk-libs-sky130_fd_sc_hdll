* File: sky130_fd_sc_hdll__and2_6.spice
* Created: Wed Sep  2 08:21:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and2_6.pex.spice"
.subckt sky130_fd_sc_hdll__and2_6  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1001 A_293_47# N_B_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65 AD=0.078
+ AS=0.2405 PD=0.89 PS=2.04 NRD=11.988 NRS=19.38 M=1 R=4.33333 SA=75000.3
+ SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1008 N_A_117_297#_M1008_d N_A_M1008_g A_293_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.078 PD=0.92 PS=0.89 NRD=0 NRS=11.988 M=1 R=4.33333 SA=75000.7
+ SB=75004 A=0.0975 P=1.6 MULT=1
MM1009 N_A_117_297#_M1008_d N_A_M1009_g A_131_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.091 PD=0.92 PS=0.93 NRD=0 NRS=15.684 M=1 R=4.33333 SA=75001.1
+ SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1012 A_131_47# N_B_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.13975 PD=0.93 PS=1.08 NRD=15.684 NRS=12.912 M=1 R=4.33333 SA=75001.5
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1012_s N_A_117_297#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.13975 AS=0.08775 PD=1.08 PS=0.92 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A_117_297#_M1006_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.5
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1006_d N_A_117_297#_M1010_g N_X_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1014_d N_A_117_297#_M1014_g N_X_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.5
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1014_d N_A_117_297#_M1017_g N_X_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75004
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1019_d N_A_117_297#_M1019_g N_X_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2145 AS=0.08775 PD=1.96 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75004.4
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1007 N_A_117_297#_M1007_d N_B_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90004.4 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_A_117_297#_M1007_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90004 A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1002_d N_A_M1018_g N_A_117_297#_M1018_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1015 N_A_117_297#_M1018_s N_B_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90003 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1015_s N_A_117_297#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_A_117_297#_M1003_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1003_d N_A_117_297#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_A_117_297#_M1011_g N_X_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1011_d N_A_117_297#_M1013_g N_X_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.9 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1016 N_VPWR_M1016_d N_A_117_297#_M1016_g N_X_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.29 AS=0.145 PD=2.58 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.4 SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=9.4695 P=15.01
*
.include "sky130_fd_sc_hdll__and2_6.pxi.spice"
*
.ends
*
*
