* File: sky130_fd_sc_hdll__a21o_8.pex.spice
* Created: Thu Aug 27 18:53:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A21O_8%A2 1 3 4 6 7 9 10 12 14 15 16 18 19 23 26
c88 18 0 1.53044e-19 $X=1.79 $Y=1.46
c89 14 0 1.34369e-19 $X=0.61 $Y=1.46
c90 10 0 1.86168e-19 $X=1.905 $Y=1.41
r91 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.49
+ $Y=1.16 $X2=0.49 $Y2=1.16
r92 26 30 12.7504 $w=2.33e-07 $l=2.6e-07 $layer=LI1_cond $X=0.23 $Y=1.172
+ $X2=0.49 $Y2=1.172
r93 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.16 $X2=1.88 $Y2=1.16
r94 20 23 4.41361 $w=2.33e-07 $l=9e-08 $layer=LI1_cond $X=1.79 $Y=1.172 $X2=1.88
+ $Y2=1.172
r95 19 30 1.7164 $w=2.33e-07 $l=3.5e-08 $layer=LI1_cond $X=0.525 $Y=1.172
+ $X2=0.49 $Y2=1.172
r96 17 20 2.6346 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=1.79 $Y=1.29 $X2=1.79
+ $Y2=1.172
r97 17 18 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.79 $Y=1.29
+ $X2=1.79 $Y2=1.46
r98 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.705 $Y=1.545
+ $X2=1.79 $Y2=1.46
r99 15 16 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=1.705 $Y=1.545
+ $X2=0.695 $Y2=1.545
r100 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.46
+ $X2=0.695 $Y2=1.545
r101 13 19 7.04737 $w=2.35e-07 $l=1.54771e-07 $layer=LI1_cond $X=0.61 $Y=1.29
+ $X2=0.525 $Y2=1.172
r102 13 14 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.61 $Y=1.29
+ $X2=0.61 $Y2=1.46
r103 10 24 51.486 $w=2.55e-07 $l=2.62202e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.88 $Y2=1.16
r104 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r105 7 24 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.82 $Y=0.995
+ $X2=1.88 $Y2=1.16
r106 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.82 $Y=0.995
+ $X2=1.82 $Y2=0.56
r107 4 29 38.5416 $w=3.03e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.58 $Y=0.995
+ $X2=0.49 $Y2=1.16
r108 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.58 $Y=0.995
+ $X2=0.58 $Y2=0.56
r109 1 29 47.6478 $w=3.03e-07 $l=2.52488e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.49 $Y2=1.16
r110 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_8%A1 1 3 4 6 7 9 10 12 13 19 20
r52 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.202
+ $X2=1.435 $Y2=1.202
r53 18 20 5.07368 $w=3.8e-07 $l=4e-08 $layer=POLY_cond $X=1.37 $Y=1.202 $X2=1.41
+ $Y2=1.202
r54 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.37
+ $Y=1.16 $X2=1.37 $Y2=1.16
r55 16 18 48.2 $w=3.8e-07 $l=3.8e-07 $layer=POLY_cond $X=0.99 $Y=1.202 $X2=1.37
+ $Y2=1.202
r56 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r57 13 19 10.7888 $w=2.33e-07 $l=2.2e-07 $layer=LI1_cond $X=1.15 $Y=1.172
+ $X2=1.37 $Y2=1.172
r58 10 21 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r59 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r60 7 20 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.202
r61 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995 $X2=1.41
+ $Y2=0.56
r62 4 16 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r63 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995 $X2=0.99
+ $Y2=0.56
r64 1 15 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r65 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_8%B1 1 3 4 6 7 9 10 12 13 18
c54 1 0 1.53044e-19 $X=2.375 $Y=1.41
r55 18 20 24.3634 $w=3.66e-07 $l=1.85e-07 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=3.03 $Y2=1.202
r56 17 18 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.845 $Y2=1.202
r57 16 17 55.3115 $w=3.66e-07 $l=4.2e-07 $layer=POLY_cond $X=2.4 $Y=1.202
+ $X2=2.82 $Y2=1.202
r58 15 16 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.4 $Y2=1.202
r59 13 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.03
+ $Y=1.16 $X2=3.03 $Y2=1.16
r60 10 18 19.3576 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r61 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r62 7 17 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=1.202
r63 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.82 $Y=0.995 $X2=2.82
+ $Y2=0.56
r64 4 16 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.4 $Y=0.995 $X2=2.4
+ $Y2=1.202
r65 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.4 $Y=0.995 $X2=2.4
+ $Y2=0.56
r66 1 15 19.3576 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r67 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_8%A_213_47# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 51 52 54 55 57 60 62 63
+ 66 71 72 75 76 81 84 86 105
r215 105 106 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=7.1 $Y=1.202
+ $X2=7.125 $Y2=1.202
r216 104 105 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=6.68 $Y=1.202
+ $X2=7.1 $Y2=1.202
r217 103 104 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=6.655 $Y=1.202
+ $X2=6.68 $Y2=1.202
r218 102 103 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=6.185 $Y=1.202
+ $X2=6.655 $Y2=1.202
r219 101 102 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=6.16 $Y=1.202
+ $X2=6.185 $Y2=1.202
r220 98 99 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=5.715 $Y=1.202
+ $X2=5.74 $Y2=1.202
r221 97 98 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=5.245 $Y=1.202
+ $X2=5.715 $Y2=1.202
r222 96 97 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=5.22 $Y=1.202
+ $X2=5.245 $Y2=1.202
r223 95 96 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=4.8 $Y=1.202
+ $X2=5.22 $Y2=1.202
r224 94 95 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=4.775 $Y=1.202
+ $X2=4.8 $Y2=1.202
r225 93 94 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=4.305 $Y=1.202
+ $X2=4.775 $Y2=1.202
r226 92 93 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=4.28 $Y=1.202
+ $X2=4.305 $Y2=1.202
r227 89 90 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=3.835 $Y=1.202
+ $X2=3.86 $Y2=1.202
r228 86 87 6.88461 $w=2.98e-07 $l=1.7e-07 $layer=LI1_cond $X=2.595 $Y=1.96
+ $X2=2.595 $Y2=1.79
r229 82 101 24.8859 $w=3.68e-07 $l=1.9e-07 $layer=POLY_cond $X=5.97 $Y=1.202
+ $X2=6.16 $Y2=1.202
r230 82 99 30.125 $w=3.68e-07 $l=2.3e-07 $layer=POLY_cond $X=5.97 $Y=1.202
+ $X2=5.74 $Y2=1.202
r231 81 82 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=5.97
+ $Y=1.16 $X2=5.97 $Y2=1.16
r232 79 92 45.8424 $w=3.68e-07 $l=3.5e-07 $layer=POLY_cond $X=3.93 $Y=1.202
+ $X2=4.28 $Y2=1.202
r233 79 90 9.16848 $w=3.68e-07 $l=7e-08 $layer=POLY_cond $X=3.93 $Y=1.202
+ $X2=3.86 $Y2=1.202
r234 78 81 97.9577 $w=2.38e-07 $l=2.04e-06 $layer=LI1_cond $X=3.93 $Y=1.155
+ $X2=5.97 $Y2=1.155
r235 78 79 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=3.93
+ $Y=1.16 $X2=3.93 $Y2=1.16
r236 76 78 9.3636 $w=2.38e-07 $l=1.95e-07 $layer=LI1_cond $X=3.735 $Y=1.155
+ $X2=3.93 $Y2=1.155
r237 75 76 7.07814 $w=2.4e-07 $l=1.56844e-07 $layer=LI1_cond $X=3.65 $Y=1.035
+ $X2=3.735 $Y2=1.155
r238 74 75 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.65 $Y=0.885
+ $X2=3.65 $Y2=1.035
r239 73 84 3.9099 $w=2.1e-07 $l=1.5e-07 $layer=LI1_cond $X=2.745 $Y=0.78
+ $X2=2.595 $Y2=0.78
r240 72 74 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.565 $Y=0.78
+ $X2=3.65 $Y2=0.885
r241 72 73 43.3074 $w=2.08e-07 $l=8.2e-07 $layer=LI1_cond $X=3.565 $Y=0.78
+ $X2=2.745 $Y2=0.78
r242 71 87 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=2.57 $Y=1.62
+ $X2=2.57 $Y2=1.79
r243 68 84 2.27033 $w=2.5e-07 $l=1.16833e-07 $layer=LI1_cond $X=2.57 $Y=0.885
+ $X2=2.595 $Y2=0.78
r244 68 71 33.8818 $w=2.48e-07 $l=7.35e-07 $layer=LI1_cond $X=2.57 $Y=0.885
+ $X2=2.57 $Y2=1.62
r245 64 84 2.27033 $w=3e-07 $l=1.05e-07 $layer=LI1_cond $X=2.595 $Y=0.675
+ $X2=2.595 $Y2=0.78
r246 64 66 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=2.595 $Y=0.675
+ $X2=2.595 $Y2=0.42
r247 62 84 3.9099 $w=2.1e-07 $l=1.5e-07 $layer=LI1_cond $X=2.445 $Y=0.78
+ $X2=2.595 $Y2=0.78
r248 62 63 57.039 $w=2.08e-07 $l=1.08e-06 $layer=LI1_cond $X=2.445 $Y=0.78
+ $X2=1.365 $Y2=0.78
r249 58 63 7.26367 $w=2.1e-07 $l=2.11069e-07 $layer=LI1_cond $X=1.2 $Y=0.675
+ $X2=1.365 $Y2=0.78
r250 58 60 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=0.675
+ $X2=1.2 $Y2=0.38
r251 55 106 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.202
r252 55 57 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.985
r253 52 105 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.1 $Y=0.995
+ $X2=7.1 $Y2=1.202
r254 52 54 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.1 $Y=0.995
+ $X2=7.1 $Y2=0.56
r255 49 104 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.68 $Y=0.995
+ $X2=6.68 $Y2=1.202
r256 49 51 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.68 $Y=0.995
+ $X2=6.68 $Y2=0.56
r257 46 103 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.202
r258 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.985
r259 43 102 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.202
r260 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.985
r261 40 101 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=1.202
r262 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=0.56
r263 37 99 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.74 $Y=0.995
+ $X2=5.74 $Y2=1.202
r264 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.74 $Y=0.995
+ $X2=5.74 $Y2=0.56
r265 34 98 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.202
r266 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.985
r267 31 97 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.202
r268 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.985
r269 28 96 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.22 $Y=0.995
+ $X2=5.22 $Y2=1.202
r270 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.22 $Y=0.995
+ $X2=5.22 $Y2=0.56
r271 25 95 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.8 $Y=0.995
+ $X2=4.8 $Y2=1.202
r272 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.8 $Y=0.995
+ $X2=4.8 $Y2=0.56
r273 22 94 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.202
r274 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
r275 19 93 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.202
r276 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.985
r277 16 92 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.28 $Y=0.995
+ $X2=4.28 $Y2=1.202
r278 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.28 $Y=0.995
+ $X2=4.28 $Y2=0.56
r279 13 90 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.86 $Y=0.995
+ $X2=3.86 $Y2=1.202
r280 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.86 $Y=0.995
+ $X2=3.86 $Y2=0.56
r281 10 89 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.202
r282 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.985
r283 3 86 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.96
r284 3 71 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.62
r285 2 66 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=2.475
+ $Y=0.235 $X2=2.61 $Y2=0.42
r286 1 60 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_8%A_27_297# 1 2 3 4 15 19 21 25 28 33 35 36
+ 39 41 43 44
c71 33 0 1.86168e-19 $X=2.14 $Y=1.63
r72 37 39 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=3.08 $Y=2.295
+ $X2=3.08 $Y2=1.87
r73 35 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.915 $Y=2.38
+ $X2=3.08 $Y2=2.295
r74 35 36 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.915 $Y=2.38
+ $X2=2.275 $Y2=2.38
r75 31 44 3.52026 $w=2.65e-07 $l=1.00995e-07 $layer=LI1_cond $X=2.16 $Y=1.8
+ $X2=2.125 $Y2=1.885
r76 31 33 8.51806 $w=2.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.16 $Y=1.8 $X2=2.16
+ $Y2=1.63
r77 30 44 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=1.97
+ $X2=2.125 $Y2=1.885
r78 28 36 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.125 $Y=2.295
+ $X2=2.275 $Y2=2.38
r79 28 30 12.4848 $w=2.98e-07 $l=3.25e-07 $layer=LI1_cond $X=2.125 $Y=2.295
+ $X2=2.125 $Y2=1.97
r80 26 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=1.885
+ $X2=1.2 $Y2=1.885
r81 25 44 2.98021 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.975 $Y=1.885
+ $X2=2.125 $Y2=1.885
r82 25 26 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.975 $Y=1.885
+ $X2=1.365 $Y2=1.885
r83 22 41 3.3845 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=1.885
+ $X2=0.26 $Y2=1.885
r84 21 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=1.885
+ $X2=1.2 $Y2=1.885
r85 21 22 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.035 $Y=1.885
+ $X2=0.425 $Y2=1.885
r86 17 41 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.97
+ $X2=0.26 $Y2=1.885
r87 17 19 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=0.26 $Y=1.97 $X2=0.26
+ $Y2=2
r88 13 41 3.19717 $w=2.95e-07 $l=1.00995e-07 $layer=LI1_cond $X=0.225 $Y=1.8
+ $X2=0.26 $Y2=1.885
r89 13 15 6.20546 $w=2.58e-07 $l=1.4e-07 $layer=LI1_cond $X=0.225 $Y=1.8
+ $X2=0.225 $Y2=1.66
r90 4 39 300 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=1.87
r91 3 33 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.63
r92 3 30 300 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.97
r93 2 43 300 $w=1.7e-07 $l=4.66905e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.885
r94 1 19 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
r95 1 15 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_8%VPWR 1 2 3 4 5 6 7 24 26 30 34 40 44 48 52
+ 57 58 60 61 63 64 66 67 69 70 71 73 98 99 102 105
r123 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r124 103 106 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r125 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r126 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r127 96 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r128 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r129 93 96 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r130 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r131 90 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r132 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r133 87 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r134 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r135 84 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r136 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r137 81 84 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r138 81 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r139 80 83 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r140 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r141 78 105 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=1.67 $Y2=2.72
r142 78 80 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=2.07 $Y2=2.72
r143 73 102 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.73 $Y2=2.72
r144 73 75 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r145 71 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r146 71 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r147 69 95 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=7.215 $Y=2.72
+ $X2=7.13 $Y2=2.72
r148 69 70 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=7.215 $Y=2.72
+ $X2=7.37 $Y2=2.72
r149 68 98 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=7.525 $Y=2.72
+ $X2=7.59 $Y2=2.72
r150 68 70 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=7.525 $Y=2.72
+ $X2=7.37 $Y2=2.72
r151 66 92 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=6.255 $Y=2.72
+ $X2=6.21 $Y2=2.72
r152 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.255 $Y=2.72
+ $X2=6.42 $Y2=2.72
r153 65 95 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=6.585 $Y=2.72
+ $X2=7.13 $Y2=2.72
r154 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.585 $Y=2.72
+ $X2=6.42 $Y2=2.72
r155 63 89 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.315 $Y=2.72
+ $X2=5.29 $Y2=2.72
r156 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.315 $Y=2.72
+ $X2=5.48 $Y2=2.72
r157 62 92 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.645 $Y=2.72
+ $X2=6.21 $Y2=2.72
r158 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.645 $Y=2.72
+ $X2=5.48 $Y2=2.72
r159 60 86 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.375 $Y=2.72
+ $X2=4.37 $Y2=2.72
r160 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.375 $Y=2.72
+ $X2=4.54 $Y2=2.72
r161 59 89 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.705 $Y=2.72
+ $X2=5.29 $Y2=2.72
r162 59 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=2.72
+ $X2=4.54 $Y2=2.72
r163 57 83 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.485 $Y=2.72
+ $X2=3.45 $Y2=2.72
r164 57 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.485 $Y=2.72
+ $X2=3.61 $Y2=2.72
r165 56 86 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.735 $Y=2.72
+ $X2=4.37 $Y2=2.72
r166 56 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.735 $Y=2.72
+ $X2=3.61 $Y2=2.72
r167 52 55 25.2794 $w=3.08e-07 $l=6.8e-07 $layer=LI1_cond $X=7.37 $Y=1.63
+ $X2=7.37 $Y2=2.31
r168 50 70 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.37 $Y=2.635
+ $X2=7.37 $Y2=2.72
r169 50 55 12.0821 $w=3.08e-07 $l=3.25e-07 $layer=LI1_cond $X=7.37 $Y=2.635
+ $X2=7.37 $Y2=2.31
r170 46 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=2.72
r171 46 48 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=1.87
r172 42 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2.72
r173 42 44 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=1.87
r174 38 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=2.635
+ $X2=4.54 $Y2=2.72
r175 38 40 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=4.54 $Y=2.635
+ $X2=4.54 $Y2=1.87
r176 34 37 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=3.61 $Y=1.66
+ $X2=3.61 $Y2=2.34
r177 32 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.61 $Y=2.635
+ $X2=3.61 $Y2=2.72
r178 32 37 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.61 $Y=2.635
+ $X2=3.61 $Y2=2.34
r179 28 105 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.72
r180 28 30 14.0854 $w=2.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.305
r181 27 102 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.865 $Y=2.72
+ $X2=0.73 $Y2=2.72
r182 26 105 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.535 $Y=2.72
+ $X2=1.67 $Y2=2.72
r183 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.535 $Y=2.72
+ $X2=0.865 $Y2=2.72
r184 22 102 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.72
r185 22 24 14.0854 $w=2.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.305
r186 7 55 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=7.215
+ $Y=1.485 $X2=7.36 $Y2=2.31
r187 7 52 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.215
+ $Y=1.485 $X2=7.36 $Y2=1.63
r188 6 48 300 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_PDIFF $count=2 $X=6.275
+ $Y=1.485 $X2=6.42 $Y2=1.87
r189 5 44 300 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_PDIFF $count=2 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=1.87
r190 4 40 300 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_PDIFF $count=2 $X=4.395
+ $Y=1.485 $X2=4.54 $Y2=1.87
r191 3 37 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=3.475
+ $Y=1.485 $X2=3.6 $Y2=2.34
r192 3 34 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=3.475
+ $Y=1.485 $X2=3.6 $Y2=1.66
r193 2 30 600 $w=1.7e-07 $l=8.8955e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.305
r194 1 24 600 $w=1.7e-07 $l=8.8955e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.305
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_8%X 1 2 3 4 5 6 7 8 27 31 35 36 37 38 41 45
+ 49 51 55 59 63 65 69 71 73 77 78 79 80 82 87
r128 84 87 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=6.67 $Y=1.445
+ $X2=6.67 $Y2=1.19
r129 81 87 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=6.67 $Y=0.865
+ $X2=6.67 $Y2=1.19
r130 81 82 3.24686 $w=2.9e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.67 $Y=0.865
+ $X2=6.8 $Y2=0.78
r131 73 75 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.89 $Y=1.62
+ $X2=6.89 $Y2=2.3
r132 71 84 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=6.89 $Y=1.53
+ $X2=6.67 $Y2=1.53
r133 71 73 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=6.89 $Y=1.615
+ $X2=6.89 $Y2=1.62
r134 67 82 3.24686 $w=2.9e-07 $l=1.25499e-07 $layer=LI1_cond $X=6.89 $Y=0.695
+ $X2=6.8 $Y2=0.78
r135 67 69 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.89 $Y=0.695
+ $X2=6.89 $Y2=0.36
r136 66 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.115 $Y=0.78
+ $X2=5.95 $Y2=0.78
r137 65 82 3.3199 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=6.545 $Y=0.78
+ $X2=6.8 $Y2=0.78
r138 65 66 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=6.545 $Y=0.78
+ $X2=6.115 $Y2=0.78
r139 64 80 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.085 $Y=1.53
+ $X2=5.95 $Y2=1.53
r140 63 84 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.545 $Y=1.53
+ $X2=6.67 $Y2=1.53
r141 63 64 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.545 $Y=1.53
+ $X2=6.085 $Y2=1.53
r142 59 61 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.95 $Y=1.62
+ $X2=5.95 $Y2=2.3
r143 57 80 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=1.615
+ $X2=5.95 $Y2=1.53
r144 57 59 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=5.95 $Y=1.615
+ $X2=5.95 $Y2=1.62
r145 53 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=0.695
+ $X2=5.95 $Y2=0.78
r146 53 55 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.95 $Y=0.695
+ $X2=5.95 $Y2=0.36
r147 52 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.175 $Y=0.78
+ $X2=5.01 $Y2=0.78
r148 51 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.785 $Y=0.78
+ $X2=5.95 $Y2=0.78
r149 51 52 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.785 $Y=0.78
+ $X2=5.175 $Y2=0.78
r150 50 78 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.145 $Y=1.53
+ $X2=5.01 $Y2=1.53
r151 49 80 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.815 $Y=1.53
+ $X2=5.95 $Y2=1.53
r152 49 50 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.815 $Y=1.53
+ $X2=5.145 $Y2=1.53
r153 45 47 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.01 $Y=1.62
+ $X2=5.01 $Y2=2.3
r154 43 78 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.01 $Y=1.615
+ $X2=5.01 $Y2=1.53
r155 43 45 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=5.01 $Y=1.615
+ $X2=5.01 $Y2=1.62
r156 39 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.01 $Y=0.695
+ $X2=5.01 $Y2=0.78
r157 39 41 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.01 $Y=0.695
+ $X2=5.01 $Y2=0.36
r158 37 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.845 $Y=0.78
+ $X2=5.01 $Y2=0.78
r159 37 38 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.845 $Y=0.78
+ $X2=4.235 $Y2=0.78
r160 35 78 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.875 $Y=1.53
+ $X2=5.01 $Y2=1.53
r161 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.875 $Y=1.53
+ $X2=4.205 $Y2=1.53
r162 31 33 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.07 $Y=1.62
+ $X2=4.07 $Y2=2.3
r163 29 36 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.07 $Y=1.615
+ $X2=4.205 $Y2=1.53
r164 29 31 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=4.07 $Y=1.615
+ $X2=4.07 $Y2=1.62
r165 25 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.07 $Y=0.695
+ $X2=4.235 $Y2=0.78
r166 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.07 $Y=0.695
+ $X2=4.07 $Y2=0.36
r167 8 75 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=2.3
r168 8 73 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=1.62
r169 7 61 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=2.3
r170 7 59 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=1.62
r171 6 47 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=2.3
r172 6 45 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=1.62
r173 5 33 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=2.3
r174 5 31 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=1.62
r175 4 69 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=6.755
+ $Y=0.235 $X2=6.89 $Y2=0.36
r176 3 55 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=5.815
+ $Y=0.235 $X2=5.95 $Y2=0.36
r177 2 41 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=4.875
+ $Y=0.235 $X2=5.01 $Y2=0.36
r178 1 27 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=3.935
+ $Y=0.235 $X2=4.07 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_8%VGND 1 2 3 4 5 6 7 22 24 28 34 38 42 46 49
+ 50 52 53 55 56 58 59 60 62 84 85 91 96 102
r116 101 102 10.0909 $w=5.88e-07 $l=1.65e-07 $layer=LI1_cond $X=3.57 $Y=0.21
+ $X2=3.735 $Y2=0.21
r117 98 101 2.4327 $w=5.88e-07 $l=1.2e-07 $layer=LI1_cond $X=3.45 $Y=0.21
+ $X2=3.57 $Y2=0.21
r118 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r119 95 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r120 94 98 9.32536 $w=5.88e-07 $l=4.6e-07 $layer=LI1_cond $X=2.99 $Y=0.21
+ $X2=3.45 $Y2=0.21
r121 94 96 8.2664 $w=5.88e-07 $l=7.5e-08 $layer=LI1_cond $X=2.99 $Y=0.21
+ $X2=2.915 $Y2=0.21
r122 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r123 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r124 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r125 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r126 82 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=7.59
+ $Y2=0
r127 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r128 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r129 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r130 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r131 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r132 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r133 73 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.45
+ $Y2=0
r134 72 102 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.37 $Y=0
+ $X2=3.735 $Y2=0
r135 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r136 69 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r137 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r138 66 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r139 65 68 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r140 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r141 63 88 4.56433 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=0.535 $Y=0
+ $X2=0.267 $Y2=0
r142 63 65 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.535 $Y=0
+ $X2=0.69 $Y2=0
r143 62 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=2.11
+ $Y2=0
r144 62 68 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.945 $Y=0
+ $X2=1.61 $Y2=0
r145 60 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r146 60 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r147 58 81 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.225 $Y=0 $X2=7.13
+ $Y2=0
r148 58 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.225 $Y=0 $X2=7.35
+ $Y2=0
r149 57 84 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.475 $Y=0
+ $X2=7.59 $Y2=0
r150 57 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.475 $Y=0 $X2=7.35
+ $Y2=0
r151 55 78 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.285 $Y=0 $X2=6.21
+ $Y2=0
r152 55 56 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.285 $Y=0 $X2=6.42
+ $Y2=0
r153 54 81 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.555 $Y=0
+ $X2=7.13 $Y2=0
r154 54 56 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.555 $Y=0 $X2=6.42
+ $Y2=0
r155 52 75 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=5.345 $Y=0 $X2=5.29
+ $Y2=0
r156 52 53 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.345 $Y=0 $X2=5.48
+ $Y2=0
r157 51 78 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.615 $Y=0
+ $X2=6.21 $Y2=0
r158 51 53 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.615 $Y=0 $X2=5.48
+ $Y2=0
r159 49 72 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.405 $Y=0 $X2=4.37
+ $Y2=0
r160 49 50 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.405 $Y=0 $X2=4.54
+ $Y2=0
r161 48 75 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.675 $Y=0 $X2=5.29
+ $Y2=0
r162 48 50 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.675 $Y=0 $X2=4.54
+ $Y2=0
r163 44 59 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.35 $Y=0.085
+ $X2=7.35 $Y2=0
r164 44 46 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=7.35 $Y=0.085
+ $X2=7.35 $Y2=0.36
r165 40 56 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0
r166 40 42 11.7378 $w=2.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0.36
r167 36 53 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0
r168 36 38 11.7378 $w=2.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.36
r169 32 50 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0
r170 32 34 11.7378 $w=2.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0.36
r171 31 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.11
+ $Y2=0
r172 31 96 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.915
+ $Y2=0
r173 26 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.11 $Y2=0
r174 26 28 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.11 $Y2=0.38
r175 22 88 3.20184 $w=3.3e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.37 $Y=0.085
+ $X2=0.267 $Y2=0
r176 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.37 $Y=0.085
+ $X2=0.37 $Y2=0.38
r177 7 46 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=7.175
+ $Y=0.235 $X2=7.31 $Y2=0.36
r178 6 42 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=6.235
+ $Y=0.235 $X2=6.42 $Y2=0.36
r179 5 38 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=5.295
+ $Y=0.235 $X2=5.48 $Y2=0.36
r180 4 34 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=4.355
+ $Y=0.235 $X2=4.54 $Y2=0.36
r181 3 101 91 $w=1.7e-07 $l=7.43976e-07 $layer=licon1_NDIFF $count=2 $X=2.895
+ $Y=0.235 $X2=3.57 $Y2=0.38
r182 2 28 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.235 $X2=2.11 $Y2=0.38
r183 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.245
+ $Y=0.235 $X2=0.37 $Y2=0.38
.ends

