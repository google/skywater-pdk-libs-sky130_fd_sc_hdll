* File: sky130_fd_sc_hdll__o2bb2a_4.pxi.spice
* Created: Thu Aug 27 19:21:56 2020
* 
x_PM_SKY130_FD_SC_HDLL__O2BB2A_4%B1 N_B1_c_123_n N_B1_M1009_g N_B1_c_124_n
+ N_B1_M1017_g N_B1_c_125_n N_B1_M1014_g N_B1_c_126_n N_B1_M1018_g N_B1_c_131_n
+ N_B1_c_127_n B1 N_B1_c_128_n PM_SKY130_FD_SC_HDLL__O2BB2A_4%B1
x_PM_SKY130_FD_SC_HDLL__O2BB2A_4%B2 N_B2_c_199_n N_B2_M1006_g N_B2_c_203_n
+ N_B2_M1001_g N_B2_c_204_n N_B2_M1023_g N_B2_c_200_n N_B2_M1027_g B2
+ N_B2_c_202_n PM_SKY130_FD_SC_HDLL__O2BB2A_4%B2
x_PM_SKY130_FD_SC_HDLL__O2BB2A_4%A_455_21# N_A_455_21#_M1016_s
+ N_A_455_21#_M1004_s N_A_455_21#_M1019_d N_A_455_21#_c_246_n
+ N_A_455_21#_M1021_g N_A_455_21#_c_256_n N_A_455_21#_M1005_g
+ N_A_455_21#_c_247_n N_A_455_21#_M1022_g N_A_455_21#_c_257_n
+ N_A_455_21#_M1011_g N_A_455_21#_c_248_n N_A_455_21#_c_249_n
+ N_A_455_21#_c_250_n N_A_455_21#_c_251_n N_A_455_21#_c_267_p
+ N_A_455_21#_c_318_p N_A_455_21#_c_276_p N_A_455_21#_c_252_n
+ N_A_455_21#_c_277_p N_A_455_21#_c_253_n N_A_455_21#_c_254_n
+ N_A_455_21#_c_279_p N_A_455_21#_c_255_n
+ PM_SKY130_FD_SC_HDLL__O2BB2A_4%A_455_21#
x_PM_SKY130_FD_SC_HDLL__O2BB2A_4%A1_N N_A1_N_c_367_n N_A1_N_M1004_g
+ N_A1_N_c_368_n N_A1_N_M1000_g N_A1_N_c_369_n N_A1_N_M1026_g N_A1_N_c_370_n
+ N_A1_N_M1010_g N_A1_N_c_374_n N_A1_N_c_375_n A1_N
+ PM_SKY130_FD_SC_HDLL__O2BB2A_4%A1_N
x_PM_SKY130_FD_SC_HDLL__O2BB2A_4%A2_N N_A2_N_c_451_n N_A2_N_M1016_g
+ N_A2_N_c_455_n N_A2_N_M1013_g N_A2_N_c_456_n N_A2_N_M1019_g N_A2_N_c_452_n
+ N_A2_N_M1025_g A2_N N_A2_N_c_453_n N_A2_N_c_454_n A2_N
+ PM_SKY130_FD_SC_HDLL__O2BB2A_4%A2_N
x_PM_SKY130_FD_SC_HDLL__O2BB2A_4%A_211_297# N_A_211_297#_M1021_s
+ N_A_211_297#_M1001_d N_A_211_297#_M1005_s N_A_211_297#_c_497_n
+ N_A_211_297#_M1002_g N_A_211_297#_c_504_n N_A_211_297#_M1003_g
+ N_A_211_297#_c_498_n N_A_211_297#_M1007_g N_A_211_297#_c_505_n
+ N_A_211_297#_M1012_g N_A_211_297#_c_499_n N_A_211_297#_M1008_g
+ N_A_211_297#_c_506_n N_A_211_297#_M1015_g N_A_211_297#_c_507_n
+ N_A_211_297#_M1024_g N_A_211_297#_c_500_n N_A_211_297#_M1020_g
+ N_A_211_297#_c_514_n N_A_211_297#_c_501_n N_A_211_297#_c_553_n
+ N_A_211_297#_c_600_p N_A_211_297#_c_519_n N_A_211_297#_c_529_n
+ N_A_211_297#_c_508_n N_A_211_297#_c_554_n N_A_211_297#_c_509_n
+ N_A_211_297#_c_510_n N_A_211_297#_c_502_n N_A_211_297#_c_503_n
+ PM_SKY130_FD_SC_HDLL__O2BB2A_4%A_211_297#
x_PM_SKY130_FD_SC_HDLL__O2BB2A_4%VPWR N_VPWR_M1009_s N_VPWR_M1014_s
+ N_VPWR_M1011_d N_VPWR_M1013_s N_VPWR_M1026_d N_VPWR_M1012_s N_VPWR_M1024_s
+ N_VPWR_c_652_n N_VPWR_c_653_n N_VPWR_c_654_n N_VPWR_c_655_n N_VPWR_c_656_n
+ N_VPWR_c_657_n N_VPWR_c_658_n N_VPWR_c_659_n N_VPWR_c_660_n N_VPWR_c_661_n
+ N_VPWR_c_662_n N_VPWR_c_663_n N_VPWR_c_664_n N_VPWR_c_665_n N_VPWR_c_666_n
+ VPWR N_VPWR_c_667_n N_VPWR_c_668_n N_VPWR_c_651_n N_VPWR_c_670_n
+ N_VPWR_c_671_n N_VPWR_c_672_n PM_SKY130_FD_SC_HDLL__O2BB2A_4%VPWR
x_PM_SKY130_FD_SC_HDLL__O2BB2A_4%A_117_297# N_A_117_297#_M1009_d
+ N_A_117_297#_M1023_s N_A_117_297#_c_776_n N_A_117_297#_c_777_n
+ N_A_117_297#_c_788_n N_A_117_297#_c_783_n
+ PM_SKY130_FD_SC_HDLL__O2BB2A_4%A_117_297#
x_PM_SKY130_FD_SC_HDLL__O2BB2A_4%X N_X_M1002_d N_X_M1008_d N_X_M1003_d
+ N_X_M1015_d N_X_c_803_n N_X_c_842_n N_X_c_806_n N_X_c_810_n N_X_c_792_n
+ N_X_c_793_n N_X_c_824_n N_X_c_847_n N_X_c_794_n N_X_c_795_n N_X_c_797_n X X
+ N_X_c_800_n PM_SKY130_FD_SC_HDLL__O2BB2A_4%X
x_PM_SKY130_FD_SC_HDLL__O2BB2A_4%A_27_47# N_A_27_47#_M1017_s N_A_27_47#_M1006_d
+ N_A_27_47#_M1018_s N_A_27_47#_M1022_d N_A_27_47#_c_871_n N_A_27_47#_c_872_n
+ N_A_27_47#_c_873_n N_A_27_47#_c_883_n N_A_27_47#_c_874_n N_A_27_47#_c_888_n
+ N_A_27_47#_c_889_n N_A_27_47#_c_875_n N_A_27_47#_c_876_n
+ PM_SKY130_FD_SC_HDLL__O2BB2A_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__O2BB2A_4%VGND N_VGND_M1017_d N_VGND_M1027_s
+ N_VGND_M1000_s N_VGND_M1010_s N_VGND_M1007_s N_VGND_M1020_s N_VGND_c_932_n
+ N_VGND_c_933_n N_VGND_c_934_n N_VGND_c_935_n N_VGND_c_936_n N_VGND_c_937_n
+ N_VGND_c_938_n N_VGND_c_939_n N_VGND_c_940_n N_VGND_c_941_n N_VGND_c_942_n
+ N_VGND_c_943_n N_VGND_c_944_n N_VGND_c_945_n N_VGND_c_946_n VGND
+ N_VGND_c_947_n N_VGND_c_948_n N_VGND_c_949_n N_VGND_c_950_n
+ PM_SKY130_FD_SC_HDLL__O2BB2A_4%VGND
x_PM_SKY130_FD_SC_HDLL__O2BB2A_4%A_787_47# N_A_787_47#_M1000_d
+ N_A_787_47#_M1025_d N_A_787_47#_c_1055_n N_A_787_47#_c_1072_n
+ N_A_787_47#_c_1053_n PM_SKY130_FD_SC_HDLL__O2BB2A_4%A_787_47#
cc_1 VNB N_B1_c_123_n 0.0297078f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_B1_c_124_n 0.0217065f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_3 VNB N_B1_c_125_n 0.0219092f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_4 VNB N_B1_c_126_n 0.0166732f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_5 VNB N_B1_c_127_n 0.00368755f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_6 VNB N_B1_c_128_n 0.0132328f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_7 VNB N_B2_c_199_n 0.0169338f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_8 VNB N_B2_c_200_n 0.0173947f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_9 VNB B2 0.00158382f $X=-0.19 $Y=-0.24 $X2=1.715 $Y2=1.53
cc_10 VNB N_B2_c_202_n 0.0364643f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_455_21#_c_246_n 0.0162503f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_12 VNB N_A_455_21#_c_247_n 0.0200627f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_13 VNB N_A_455_21#_c_248_n 6.87055e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_455_21#_c_249_n 0.00351905f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_455_21#_c_250_n 9.23368e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_455_21#_c_251_n 0.00586918f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_455_21#_c_252_n 0.00116072f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_455_21#_c_253_n 0.00266991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_455_21#_c_254_n 0.00739552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_455_21#_c_255_n 0.056033f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A1_N_c_367_n 0.0302091f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_22 VNB N_A1_N_c_368_n 0.0197012f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_23 VNB N_A1_N_c_369_n 0.023969f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_24 VNB N_A1_N_c_370_n 0.0169407f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_25 VNB A1_N 0.00384344f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_26 VNB N_A2_N_c_451_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_27 VNB N_A2_N_c_452_n 0.0176182f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_28 VNB N_A2_N_c_453_n 0.00334784f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.53
cc_29 VNB N_A2_N_c_454_n 0.034303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_211_297#_c_497_n 0.0166276f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_31 VNB N_A_211_297#_c_498_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_32 VNB N_A_211_297#_c_499_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_211_297#_c_500_n 0.0201731f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.53
cc_34 VNB N_A_211_297#_c_501_n 9.79172e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_211_297#_c_502_n 0.0773349f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_211_297#_c_503_n 0.00158483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_651_n 0.326667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_X_c_792_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0.435 $Y2=1.16
cc_39 VNB N_X_c_793_n 0.00241158f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_40 VNB N_X_c_794_n 0.0146676f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_X_c_795_n 0.00261326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB X 0.0228661f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_27_47#_c_871_n 0.0184392f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.16
cc_44 VNB N_A_27_47#_c_872_n 0.00393701f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_45 VNB N_A_27_47#_c_873_n 0.0101931f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_27_47#_c_874_n 0.00985012f $X=-0.19 $Y=-0.24 $X2=0.435 $Y2=1.16
cc_47 VNB N_A_27_47#_c_875_n 0.0030295f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.53
cc_48 VNB N_A_27_47#_c_876_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_932_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0.435 $Y2=1.16
cc_50 VNB N_VGND_c_933_n 0.0193072f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_51 VNB N_VGND_c_934_n 0.00467885f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.19
cc_52 VNB N_VGND_c_935_n 0.0047052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_936_n 0.0074124f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_937_n 0.00468725f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_938_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_939_n 0.0415597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_940_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_941_n 0.0424806f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_942_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_943_n 0.0201935f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_944_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_945_n 0.0195532f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_946_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_947_n 0.0130943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_948_n 0.378227f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_949_n 0.0219964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_950_n 0.00323927f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_787_47#_c_1053_n 0.00280072f $X=-0.19 $Y=-0.24 $X2=1.715 $Y2=1.53
cc_69 VPB N_B1_c_123_n 0.0301878f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_70 VPB N_B1_c_125_n 0.0247986f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_71 VPB N_B1_c_131_n 0.00826127f $X=-0.19 $Y=1.305 $X2=1.715 $Y2=1.53
cc_72 VPB N_B1_c_127_n 0.00264769f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_73 VPB N_B1_c_128_n 0.0162013f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_74 VPB N_B2_c_203_n 0.015998f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_75 VPB N_B2_c_204_n 0.0159964f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_76 VPB N_B2_c_202_n 0.0193263f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_455_21#_c_256_n 0.0155984f $X=-0.19 $Y=1.305 $X2=1.715 $Y2=1.53
cc_78 VPB N_A_455_21#_c_257_n 0.0196508f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.53
cc_79 VPB N_A_455_21#_c_250_n 0.00307961f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_455_21#_c_255_n 0.0314214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A1_N_c_367_n 0.0319081f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_82 VPB N_A1_N_c_369_n 0.0247986f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_83 VPB N_A1_N_c_374_n 0.00825943f $X=-0.19 $Y=1.305 $X2=1.715 $Y2=1.53
cc_84 VPB N_A1_N_c_375_n 0.00249295f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_85 VPB A1_N 0.00255881f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_86 VPB N_A2_N_c_455_n 0.015997f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_87 VPB N_A2_N_c_456_n 0.015996f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_88 VPB N_A2_N_c_454_n 0.0192992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_211_297#_c_504_n 0.015957f $X=-0.19 $Y=1.305 $X2=1.715 $Y2=1.53
cc_90 VPB N_A_211_297#_c_505_n 0.016165f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.53
cc_91 VPB N_A_211_297#_c_506_n 0.016148f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_92 VPB N_A_211_297#_c_507_n 0.0191635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_211_297#_c_508_n 0.00146248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_211_297#_c_509_n 0.00159726f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_211_297#_c_510_n 0.00703511f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_211_297#_c_502_n 0.0485604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_211_297#_c_503_n 0.00246423f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_652_n 0.010584f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_653_n 0.0049401f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_100 VPB N_VPWR_c_654_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_655_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_656_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_657_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_658_n 0.00518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_659_n 0.0191411f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_660_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_661_n 0.0187819f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_662_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_663_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_664_n 0.00478125f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_665_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_666_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_667_n 0.0416044f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_668_n 0.0128037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_651_n 0.0552102f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_670_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_671_n 0.0200031f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_672_n 0.0219329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_X_c_797_n 0.00245799f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB X 0.00633508f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB X 0.00263649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_X_c_800_n 0.0210463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 N_B1_c_124_n N_B2_c_199_n 0.0233179f $X=0.52 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_124 N_B1_c_123_n N_B2_c_203_n 0.0226077f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_125 N_B1_c_131_n N_B2_c_203_n 0.0169405f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_126 N_B1_c_128_n N_B2_c_203_n 9.80334e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_127 N_B1_c_125_n N_B2_c_204_n 0.0378352f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_128 N_B1_c_131_n N_B2_c_204_n 0.0122542f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_129 N_B1_c_127_n N_B2_c_204_n 0.00101445f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_130 N_B1_c_126_n N_B2_c_200_n 0.0212656f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_131 N_B1_c_123_n B2 7.71575e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_132 N_B1_c_125_n B2 2.06373e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_133 N_B1_c_131_n B2 0.0416942f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_134 N_B1_c_127_n B2 0.0117433f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_135 N_B1_c_128_n B2 0.0145168f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_136 N_B1_c_123_n N_B2_c_202_n 0.0233179f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_137 N_B1_c_125_n N_B2_c_202_n 0.0264727f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_138 N_B1_c_131_n N_B2_c_202_n 0.00803891f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_139 N_B1_c_127_n N_B2_c_202_n 0.00478003f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_140 N_B1_c_128_n N_B2_c_202_n 0.00409926f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_141 N_B1_c_126_n N_A_455_21#_c_246_n 0.0118576f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_142 N_B1_c_125_n N_A_455_21#_c_256_n 0.0361729f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_143 N_B1_c_127_n N_A_455_21#_c_256_n 7.06474e-19 $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_144 N_B1_c_125_n N_A_455_21#_c_255_n 0.0261814f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_145 N_B1_c_127_n N_A_455_21#_c_255_n 0.00111312f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_146 N_B1_c_131_n N_A_211_297#_M1001_d 0.00187091f $X=1.715 $Y=1.53 $X2=0
+ $Y2=0
cc_147 N_B1_c_125_n N_A_211_297#_c_514_n 0.0136241f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_148 N_B1_c_131_n N_A_211_297#_c_514_n 0.0218268f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_149 N_B1_c_127_n N_A_211_297#_c_514_n 0.0201576f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_150 N_B1_c_125_n N_A_211_297#_c_501_n 4.31451e-19 $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_151 N_B1_c_126_n N_A_211_297#_c_501_n 4.40557e-19 $X=1.93 $Y=0.995 $X2=0
+ $Y2=0
cc_152 N_B1_c_131_n N_A_211_297#_c_519_n 0.0135474f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_153 N_B1_c_127_n N_A_211_297#_c_508_n 8.59464e-19 $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_154 N_B1_c_125_n N_A_211_297#_c_503_n 0.00137254f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_155 N_B1_c_127_n N_A_211_297#_c_503_n 0.0402332f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_156 N_B1_c_128_n N_VPWR_M1009_s 0.00304954f $X=0.41 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_157 N_B1_c_127_n N_VPWR_M1014_s 0.00156278f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_158 N_B1_c_123_n N_VPWR_c_653_n 0.00787572f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_159 N_B1_c_128_n N_VPWR_c_653_n 0.0172375f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_160 N_B1_c_125_n N_VPWR_c_654_n 0.00300743f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_161 N_B1_c_123_n N_VPWR_c_667_n 0.00702461f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_162 N_B1_c_125_n N_VPWR_c_667_n 0.00702461f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_163 N_B1_c_123_n N_VPWR_c_651_n 0.0134462f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_164 N_B1_c_125_n N_VPWR_c_651_n 0.006985f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_165 N_B1_c_131_n N_A_117_297#_M1009_d 0.00187091f $X=1.715 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_166 N_B1_c_131_n N_A_117_297#_M1023_s 0.00172342f $X=1.715 $Y=1.53 $X2=0
+ $Y2=0
cc_167 N_B1_c_127_n N_A_117_297#_M1023_s 7.76441e-19 $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_168 N_B1_c_131_n N_A_117_297#_c_776_n 0.0143191f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_169 N_B1_c_123_n N_A_27_47#_c_872_n 5.76707e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_170 N_B1_c_124_n N_A_27_47#_c_872_n 0.0107165f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_171 N_B1_c_131_n N_A_27_47#_c_872_n 0.00780885f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_172 N_B1_c_128_n N_A_27_47#_c_872_n 0.0152041f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_173 N_B1_c_123_n N_A_27_47#_c_873_n 0.00393412f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_174 N_B1_c_128_n N_A_27_47#_c_873_n 0.0296273f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_175 N_B1_c_124_n N_A_27_47#_c_883_n 5.32212e-19 $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_176 N_B1_c_125_n N_A_27_47#_c_874_n 0.00442788f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_177 N_B1_c_126_n N_A_27_47#_c_874_n 0.0085711f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_178 N_B1_c_131_n N_A_27_47#_c_874_n 0.00848512f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_179 N_B1_c_127_n N_A_27_47#_c_874_n 0.0307661f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_180 N_B1_c_126_n N_A_27_47#_c_888_n 0.00373464f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_181 N_B1_c_126_n N_A_27_47#_c_889_n 0.00499625f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_182 N_B1_c_124_n N_VGND_c_932_n 0.00268723f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_183 N_B1_c_126_n N_VGND_c_934_n 0.00358858f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_184 N_B1_c_126_n N_VGND_c_939_n 0.00395719f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_185 N_B1_c_124_n N_VGND_c_948_n 0.00691278f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_186 N_B1_c_126_n N_VGND_c_948_n 0.00575407f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_187 N_B1_c_124_n N_VGND_c_949_n 0.00437852f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_188 N_B2_c_204_n N_A_211_297#_c_514_n 0.0108425f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_189 N_B2_c_203_n N_VPWR_c_667_n 0.00429453f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_190 N_B2_c_204_n N_VPWR_c_667_n 0.00429453f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_191 N_B2_c_203_n N_VPWR_c_651_n 0.00609021f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_192 N_B2_c_204_n N_VPWR_c_651_n 0.00609021f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_193 N_B2_c_203_n N_A_117_297#_c_777_n 0.0143148f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_194 N_B2_c_204_n N_A_117_297#_c_777_n 0.0100164f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_195 N_B2_c_199_n N_A_27_47#_c_872_n 0.00865686f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_196 B2 N_A_27_47#_c_872_n 0.00900407f $X=1.165 $Y=1.105 $X2=0 $Y2=0
cc_197 N_B2_c_199_n N_A_27_47#_c_883_n 0.00644736f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_198 N_B2_c_200_n N_A_27_47#_c_874_n 0.0117475f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_199 B2 N_A_27_47#_c_874_n 0.00552863f $X=1.165 $Y=1.105 $X2=0 $Y2=0
cc_200 N_B2_c_200_n N_A_27_47#_c_889_n 5.51986e-19 $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_201 N_B2_c_199_n N_A_27_47#_c_876_n 0.00119564f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_202 B2 N_A_27_47#_c_876_n 0.0307352f $X=1.165 $Y=1.105 $X2=0 $Y2=0
cc_203 N_B2_c_202_n N_A_27_47#_c_876_n 0.00486271f $X=1.435 $Y=1.202 $X2=0 $Y2=0
cc_204 N_B2_c_199_n N_VGND_c_932_n 0.00268723f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_205 N_B2_c_199_n N_VGND_c_933_n 0.00423334f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_206 N_B2_c_200_n N_VGND_c_933_n 0.00439206f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_207 N_B2_c_200_n N_VGND_c_934_n 0.00276126f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_208 N_B2_c_199_n N_VGND_c_948_n 0.00598581f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_209 N_B2_c_200_n N_VGND_c_948_n 0.00629903f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A_455_21#_c_249_n N_A1_N_c_367_n 0.00183713f $X=3.35 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_211 N_A_455_21#_c_250_n N_A1_N_c_367_n 0.00727379f $X=3.35 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_212 N_A_455_21#_c_267_p N_A1_N_c_367_n 0.0144083f $X=3.945 $Y=1.875 $X2=-0.19
+ $Y2=-0.24
cc_213 N_A_455_21#_c_252_n N_A1_N_c_367_n 0.00141249f $X=3.35 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_214 N_A_455_21#_c_254_n N_A1_N_c_367_n 0.00589039f $X=4.325 $Y=0.775
+ $X2=-0.19 $Y2=-0.24
cc_215 N_A_455_21#_c_255_n N_A1_N_c_367_n 0.00921846f $X=2.845 $Y=1.202
+ $X2=-0.19 $Y2=-0.24
cc_216 N_A_455_21#_c_249_n N_A1_N_c_368_n 0.00257611f $X=3.35 $Y=1.075 $X2=0
+ $Y2=0
cc_217 N_A_455_21#_c_253_n N_A1_N_c_368_n 3.90453e-19 $X=4.54 $Y=0.73 $X2=0
+ $Y2=0
cc_218 N_A_455_21#_c_254_n N_A1_N_c_368_n 0.0137356f $X=4.325 $Y=0.775 $X2=0
+ $Y2=0
cc_219 N_A_455_21#_M1004_s N_A1_N_c_374_n 0.00176577f $X=3.925 $Y=1.485 $X2=0
+ $Y2=0
cc_220 N_A_455_21#_M1019_d N_A1_N_c_374_n 0.00144684f $X=4.865 $Y=1.485 $X2=0
+ $Y2=0
cc_221 N_A_455_21#_c_276_p N_A1_N_c_374_n 0.0338481f $X=4.885 $Y=1.875 $X2=0
+ $Y2=0
cc_222 N_A_455_21#_c_277_p N_A1_N_c_374_n 0.0113442f $X=4.07 $Y=1.875 $X2=0
+ $Y2=0
cc_223 N_A_455_21#_c_254_n N_A1_N_c_374_n 0.00459871f $X=4.325 $Y=0.775 $X2=0
+ $Y2=0
cc_224 N_A_455_21#_c_279_p N_A1_N_c_374_n 0.00973329f $X=5.01 $Y=1.96 $X2=0
+ $Y2=0
cc_225 N_A_455_21#_c_250_n N_A1_N_c_375_n 0.0279483f $X=3.35 $Y=1.785 $X2=0
+ $Y2=0
cc_226 N_A_455_21#_c_267_p N_A1_N_c_375_n 0.0176425f $X=3.945 $Y=1.875 $X2=0
+ $Y2=0
cc_227 N_A_455_21#_c_252_n N_A1_N_c_375_n 0.0142914f $X=3.35 $Y=1.16 $X2=0 $Y2=0
cc_228 N_A_455_21#_c_277_p N_A1_N_c_375_n 9.22875e-19 $X=4.07 $Y=1.875 $X2=0
+ $Y2=0
cc_229 N_A_455_21#_c_254_n N_A1_N_c_375_n 0.0284297f $X=4.325 $Y=0.775 $X2=0
+ $Y2=0
cc_230 N_A_455_21#_M1019_d A1_N 4.95579e-19 $X=4.865 $Y=1.485 $X2=0 $Y2=0
cc_231 N_A_455_21#_c_279_p A1_N 0.00338168f $X=5.01 $Y=1.96 $X2=0 $Y2=0
cc_232 N_A_455_21#_c_253_n N_A2_N_c_451_n 0.00303187f $X=4.54 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_233 N_A_455_21#_c_254_n N_A2_N_c_451_n 0.00762189f $X=4.325 $Y=0.775
+ $X2=-0.19 $Y2=-0.24
cc_234 N_A_455_21#_c_276_p N_A2_N_c_455_n 0.0122287f $X=4.885 $Y=1.875 $X2=0
+ $Y2=0
cc_235 N_A_455_21#_c_276_p N_A2_N_c_456_n 0.012183f $X=4.885 $Y=1.875 $X2=0
+ $Y2=0
cc_236 N_A_455_21#_c_253_n N_A2_N_c_452_n 4.134e-19 $X=4.54 $Y=0.73 $X2=0 $Y2=0
cc_237 N_A_455_21#_c_254_n N_A2_N_c_453_n 0.0384434f $X=4.325 $Y=0.775 $X2=0
+ $Y2=0
cc_238 N_A_455_21#_c_253_n N_A2_N_c_454_n 0.0047334f $X=4.54 $Y=0.73 $X2=0 $Y2=0
cc_239 N_A_455_21#_c_246_n N_A_211_297#_c_501_n 0.00373294f $X=2.35 $Y=0.995
+ $X2=0 $Y2=0
cc_240 N_A_455_21#_c_247_n N_A_211_297#_c_501_n 0.00148773f $X=2.82 $Y=0.995
+ $X2=0 $Y2=0
cc_241 N_A_455_21#_c_249_n N_A_211_297#_c_501_n 0.00547843f $X=3.35 $Y=1.075
+ $X2=0 $Y2=0
cc_242 N_A_455_21#_c_251_n N_A_211_297#_c_501_n 0.00216081f $X=3.445 $Y=0.815
+ $X2=0 $Y2=0
cc_243 N_A_455_21#_c_255_n N_A_211_297#_c_501_n 0.00822246f $X=2.845 $Y=1.202
+ $X2=0 $Y2=0
cc_244 N_A_455_21#_c_246_n N_A_211_297#_c_529_n 0.00217268f $X=2.35 $Y=0.995
+ $X2=0 $Y2=0
cc_245 N_A_455_21#_c_247_n N_A_211_297#_c_529_n 0.0063344f $X=2.82 $Y=0.995
+ $X2=0 $Y2=0
cc_246 N_A_455_21#_c_251_n N_A_211_297#_c_529_n 0.00352442f $X=3.445 $Y=0.815
+ $X2=0 $Y2=0
cc_247 N_A_455_21#_c_257_n N_A_211_297#_c_508_n 0.00602115f $X=2.845 $Y=1.41
+ $X2=0 $Y2=0
cc_248 N_A_455_21#_c_248_n N_A_211_297#_c_508_n 0.00472924f $X=3.255 $Y=1.16
+ $X2=0 $Y2=0
cc_249 N_A_455_21#_c_250_n N_A_211_297#_c_508_n 0.00323411f $X=3.35 $Y=1.785
+ $X2=0 $Y2=0
cc_250 N_A_455_21#_c_255_n N_A_211_297#_c_508_n 0.00797233f $X=2.845 $Y=1.202
+ $X2=0 $Y2=0
cc_251 N_A_455_21#_c_248_n N_A_211_297#_c_510_n 0.0111482f $X=3.255 $Y=1.16
+ $X2=0 $Y2=0
cc_252 N_A_455_21#_c_250_n N_A_211_297#_c_510_n 0.0203587f $X=3.35 $Y=1.785
+ $X2=0 $Y2=0
cc_253 N_A_455_21#_c_267_p N_A_211_297#_c_510_n 0.0100528f $X=3.945 $Y=1.875
+ $X2=0 $Y2=0
cc_254 N_A_455_21#_c_276_p N_A_211_297#_c_510_n 0.00501218f $X=4.885 $Y=1.875
+ $X2=0 $Y2=0
cc_255 N_A_455_21#_c_277_p N_A_211_297#_c_510_n 0.00195488f $X=4.07 $Y=1.875
+ $X2=0 $Y2=0
cc_256 N_A_455_21#_c_254_n N_A_211_297#_c_510_n 0.00861998f $X=4.325 $Y=0.775
+ $X2=0 $Y2=0
cc_257 N_A_455_21#_c_279_p N_A_211_297#_c_510_n 0.00208665f $X=5.01 $Y=1.96
+ $X2=0 $Y2=0
cc_258 N_A_455_21#_c_255_n N_A_211_297#_c_510_n 0.00639596f $X=2.845 $Y=1.202
+ $X2=0 $Y2=0
cc_259 N_A_455_21#_c_256_n N_A_211_297#_c_503_n 0.0180491f $X=2.375 $Y=1.41
+ $X2=0 $Y2=0
cc_260 N_A_455_21#_c_257_n N_A_211_297#_c_503_n 0.0285171f $X=2.845 $Y=1.41
+ $X2=0 $Y2=0
cc_261 N_A_455_21#_c_248_n N_A_211_297#_c_503_n 0.0135723f $X=3.255 $Y=1.16
+ $X2=0 $Y2=0
cc_262 N_A_455_21#_c_250_n N_A_211_297#_c_503_n 0.016852f $X=3.35 $Y=1.785 $X2=0
+ $Y2=0
cc_263 N_A_455_21#_c_318_p N_A_211_297#_c_503_n 0.00825683f $X=3.445 $Y=1.875
+ $X2=0 $Y2=0
cc_264 N_A_455_21#_c_255_n N_A_211_297#_c_503_n 0.0296718f $X=2.845 $Y=1.202
+ $X2=0 $Y2=0
cc_265 N_A_455_21#_c_250_n N_VPWR_M1011_d 0.00936213f $X=3.35 $Y=1.785 $X2=0
+ $Y2=0
cc_266 N_A_455_21#_c_267_p N_VPWR_M1011_d 0.00656708f $X=3.945 $Y=1.875 $X2=0
+ $Y2=0
cc_267 N_A_455_21#_c_318_p N_VPWR_M1011_d 0.00627812f $X=3.445 $Y=1.875 $X2=0
+ $Y2=0
cc_268 N_A_455_21#_c_276_p N_VPWR_M1013_s 0.00333773f $X=4.885 $Y=1.875 $X2=0
+ $Y2=0
cc_269 N_A_455_21#_c_256_n N_VPWR_c_654_n 0.00300743f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_270 N_A_455_21#_c_276_p N_VPWR_c_655_n 0.0134451f $X=4.885 $Y=1.875 $X2=0
+ $Y2=0
cc_271 N_A_455_21#_c_267_p N_VPWR_c_659_n 0.00254499f $X=3.945 $Y=1.875 $X2=0
+ $Y2=0
cc_272 N_A_455_21#_c_276_p N_VPWR_c_659_n 0.00254499f $X=4.885 $Y=1.875 $X2=0
+ $Y2=0
cc_273 N_A_455_21#_c_277_p N_VPWR_c_659_n 0.00431749f $X=4.07 $Y=1.875 $X2=0
+ $Y2=0
cc_274 N_A_455_21#_c_276_p N_VPWR_c_661_n 0.00254499f $X=4.885 $Y=1.875 $X2=0
+ $Y2=0
cc_275 N_A_455_21#_c_279_p N_VPWR_c_661_n 0.0148962f $X=5.01 $Y=1.96 $X2=0 $Y2=0
cc_276 N_A_455_21#_M1004_s N_VPWR_c_651_n 0.00328969f $X=3.925 $Y=1.485 $X2=0
+ $Y2=0
cc_277 N_A_455_21#_M1019_d N_VPWR_c_651_n 0.00310186f $X=4.865 $Y=1.485 $X2=0
+ $Y2=0
cc_278 N_A_455_21#_c_256_n N_VPWR_c_651_n 0.00695682f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_279 N_A_455_21#_c_257_n N_VPWR_c_651_n 0.0102931f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_280 N_A_455_21#_c_267_p N_VPWR_c_651_n 0.00575145f $X=3.945 $Y=1.875 $X2=0
+ $Y2=0
cc_281 N_A_455_21#_c_318_p N_VPWR_c_651_n 7.8019e-19 $X=3.445 $Y=1.875 $X2=0
+ $Y2=0
cc_282 N_A_455_21#_c_276_p N_VPWR_c_651_n 0.0103558f $X=4.885 $Y=1.875 $X2=0
+ $Y2=0
cc_283 N_A_455_21#_c_277_p N_VPWR_c_651_n 0.0074482f $X=4.07 $Y=1.875 $X2=0
+ $Y2=0
cc_284 N_A_455_21#_c_279_p N_VPWR_c_651_n 0.00954569f $X=5.01 $Y=1.96 $X2=0
+ $Y2=0
cc_285 N_A_455_21#_c_256_n N_VPWR_c_671_n 0.00702461f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_286 N_A_455_21#_c_257_n N_VPWR_c_671_n 0.00587432f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_287 N_A_455_21#_c_257_n N_VPWR_c_672_n 0.00685266f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_288 N_A_455_21#_c_267_p N_VPWR_c_672_n 0.0184256f $X=3.945 $Y=1.875 $X2=0
+ $Y2=0
cc_289 N_A_455_21#_c_318_p N_VPWR_c_672_n 0.015863f $X=3.445 $Y=1.875 $X2=0
+ $Y2=0
cc_290 N_A_455_21#_c_246_n N_A_27_47#_c_875_n 0.0109334f $X=2.35 $Y=0.995 $X2=0
+ $Y2=0
cc_291 N_A_455_21#_c_247_n N_A_27_47#_c_875_n 0.0125971f $X=2.82 $Y=0.995 $X2=0
+ $Y2=0
cc_292 N_A_455_21#_c_248_n N_A_27_47#_c_875_n 0.0093048f $X=3.255 $Y=1.16 $X2=0
+ $Y2=0
cc_293 N_A_455_21#_c_255_n N_A_27_47#_c_875_n 0.00643661f $X=2.845 $Y=1.202
+ $X2=0 $Y2=0
cc_294 N_A_455_21#_c_254_n N_VGND_M1000_s 0.00448642f $X=4.325 $Y=0.775 $X2=0
+ $Y2=0
cc_295 N_A_455_21#_c_247_n N_VGND_c_935_n 0.00179926f $X=2.82 $Y=0.995 $X2=0
+ $Y2=0
cc_296 N_A_455_21#_c_254_n N_VGND_c_935_n 0.0131987f $X=4.325 $Y=0.775 $X2=0
+ $Y2=0
cc_297 N_A_455_21#_c_246_n N_VGND_c_939_n 0.00357877f $X=2.35 $Y=0.995 $X2=0
+ $Y2=0
cc_298 N_A_455_21#_c_247_n N_VGND_c_939_n 0.00357877f $X=2.82 $Y=0.995 $X2=0
+ $Y2=0
cc_299 N_A_455_21#_c_251_n N_VGND_c_939_n 0.00323451f $X=3.445 $Y=0.815 $X2=0
+ $Y2=0
cc_300 N_A_455_21#_c_254_n N_VGND_c_939_n 0.00102539f $X=4.325 $Y=0.775 $X2=0
+ $Y2=0
cc_301 N_A_455_21#_c_254_n N_VGND_c_941_n 0.00200011f $X=4.325 $Y=0.775 $X2=0
+ $Y2=0
cc_302 N_A_455_21#_M1016_s N_VGND_c_948_n 0.00301822f $X=4.355 $Y=0.235 $X2=0
+ $Y2=0
cc_303 N_A_455_21#_c_246_n N_VGND_c_948_n 0.00538422f $X=2.35 $Y=0.995 $X2=0
+ $Y2=0
cc_304 N_A_455_21#_c_247_n N_VGND_c_948_n 0.00668309f $X=2.82 $Y=0.995 $X2=0
+ $Y2=0
cc_305 N_A_455_21#_c_251_n N_VGND_c_948_n 0.00534938f $X=3.445 $Y=0.815 $X2=0
+ $Y2=0
cc_306 N_A_455_21#_c_254_n N_VGND_c_948_n 0.00772395f $X=4.325 $Y=0.775 $X2=0
+ $Y2=0
cc_307 N_A_455_21#_c_254_n N_A_787_47#_M1000_d 0.00191752f $X=4.325 $Y=0.775
+ $X2=-0.19 $Y2=-0.24
cc_308 N_A_455_21#_M1016_s N_A_787_47#_c_1055_n 0.00527949f $X=4.355 $Y=0.235
+ $X2=0 $Y2=0
cc_309 N_A_455_21#_c_253_n N_A_787_47#_c_1055_n 0.0201898f $X=4.54 $Y=0.73 $X2=0
+ $Y2=0
cc_310 N_A_455_21#_c_254_n N_A_787_47#_c_1055_n 0.0169115f $X=4.325 $Y=0.775
+ $X2=0 $Y2=0
cc_311 N_A_455_21#_c_253_n N_A_787_47#_c_1053_n 6.50328e-19 $X=4.54 $Y=0.73
+ $X2=0 $Y2=0
cc_312 N_A1_N_c_368_n N_A2_N_c_451_n 0.0269138f $X=3.86 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_313 N_A1_N_c_367_n N_A2_N_c_455_n 0.0362562f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_314 N_A1_N_c_374_n N_A2_N_c_455_n 0.0113465f $X=5.055 $Y=1.53 $X2=0 $Y2=0
cc_315 N_A1_N_c_375_n N_A2_N_c_455_n 9.66622e-19 $X=3.78 $Y=1.16 $X2=0 $Y2=0
cc_316 N_A1_N_c_369_n N_A2_N_c_456_n 0.0225897f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_317 N_A1_N_c_374_n N_A2_N_c_456_n 0.011241f $X=5.055 $Y=1.53 $X2=0 $Y2=0
cc_318 A1_N N_A2_N_c_456_n 0.00102676f $X=5.215 $Y=1.105 $X2=0 $Y2=0
cc_319 N_A1_N_c_370_n N_A2_N_c_452_n 0.0103419f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_320 N_A1_N_c_367_n N_A2_N_c_453_n 0.00123423f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_321 N_A1_N_c_369_n N_A2_N_c_453_n 6.98835e-19 $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_322 N_A1_N_c_374_n N_A2_N_c_453_n 0.0463302f $X=5.055 $Y=1.53 $X2=0 $Y2=0
cc_323 N_A1_N_c_375_n N_A2_N_c_453_n 0.0169406f $X=3.78 $Y=1.16 $X2=0 $Y2=0
cc_324 A1_N N_A2_N_c_453_n 0.0178646f $X=5.215 $Y=1.105 $X2=0 $Y2=0
cc_325 N_A1_N_c_367_n N_A2_N_c_454_n 0.0263659f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_326 N_A1_N_c_369_n N_A2_N_c_454_n 0.0263033f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_327 N_A1_N_c_374_n N_A2_N_c_454_n 0.00798993f $X=5.055 $Y=1.53 $X2=0 $Y2=0
cc_328 N_A1_N_c_375_n N_A2_N_c_454_n 0.002584f $X=3.78 $Y=1.16 $X2=0 $Y2=0
cc_329 A1_N N_A2_N_c_454_n 0.00398164f $X=5.215 $Y=1.105 $X2=0 $Y2=0
cc_330 N_A1_N_c_370_n N_A_211_297#_c_497_n 0.0123221f $X=5.27 $Y=0.995 $X2=0
+ $Y2=0
cc_331 N_A1_N_c_369_n N_A_211_297#_c_504_n 0.022784f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_332 A1_N N_A_211_297#_c_504_n 0.00116599f $X=5.215 $Y=1.105 $X2=0 $Y2=0
cc_333 A1_N N_A_211_297#_c_553_n 0.0128267f $X=5.215 $Y=1.105 $X2=0 $Y2=0
cc_334 A1_N N_A_211_297#_c_554_n 0.00197511f $X=5.215 $Y=1.105 $X2=0 $Y2=0
cc_335 N_A1_N_c_369_n N_A_211_297#_c_509_n 4.80357e-19 $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_336 A1_N N_A_211_297#_c_509_n 0.0232018f $X=5.215 $Y=1.105 $X2=0 $Y2=0
cc_337 N_A1_N_c_374_n N_A_211_297#_c_510_n 0.0425816f $X=5.055 $Y=1.53 $X2=0
+ $Y2=0
cc_338 N_A1_N_c_375_n N_A_211_297#_c_510_n 0.0184566f $X=3.78 $Y=1.16 $X2=0
+ $Y2=0
cc_339 A1_N N_A_211_297#_c_510_n 0.0319874f $X=5.215 $Y=1.105 $X2=0 $Y2=0
cc_340 N_A1_N_c_369_n N_A_211_297#_c_502_n 0.0265038f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_341 A1_N N_A_211_297#_c_502_n 0.00234695f $X=5.215 $Y=1.105 $X2=0 $Y2=0
cc_342 N_A1_N_c_375_n N_VPWR_M1011_d 0.00149204f $X=3.78 $Y=1.16 $X2=0 $Y2=0
cc_343 N_A1_N_c_374_n N_VPWR_M1013_s 0.00187547f $X=5.055 $Y=1.53 $X2=0 $Y2=0
cc_344 A1_N N_VPWR_M1026_d 0.00157591f $X=5.215 $Y=1.105 $X2=0 $Y2=0
cc_345 N_A1_N_c_369_n N_VPWR_c_656_n 0.00314922f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_346 A1_N N_VPWR_c_656_n 0.00550954f $X=5.215 $Y=1.105 $X2=0 $Y2=0
cc_347 N_A1_N_c_367_n N_VPWR_c_659_n 0.0053025f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_348 N_A1_N_c_369_n N_VPWR_c_661_n 0.00702461f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_349 N_A1_N_c_367_n N_VPWR_c_651_n 0.00825795f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_350 N_A1_N_c_369_n N_VPWR_c_651_n 0.0124596f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_351 N_A1_N_c_367_n N_VPWR_c_672_n 0.00514457f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_352 N_A1_N_c_368_n N_VGND_c_935_n 0.00723564f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_353 N_A1_N_c_369_n N_VGND_c_936_n 2.29798e-19 $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_354 N_A1_N_c_370_n N_VGND_c_936_n 0.00276034f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_355 A1_N N_VGND_c_936_n 0.0057781f $X=5.215 $Y=1.105 $X2=0 $Y2=0
cc_356 N_A1_N_c_368_n N_VGND_c_941_n 0.00400663f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_357 N_A1_N_c_370_n N_VGND_c_941_n 0.00585385f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_358 N_A1_N_c_368_n N_VGND_c_948_n 0.00693457f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_359 N_A1_N_c_370_n N_VGND_c_948_n 0.0107097f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_360 N_A1_N_c_368_n N_A_787_47#_c_1055_n 0.00459931f $X=3.86 $Y=0.995 $X2=0
+ $Y2=0
cc_361 N_A1_N_c_369_n N_A_787_47#_c_1053_n 0.00235048f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_362 N_A1_N_c_374_n N_A_787_47#_c_1053_n 0.00369961f $X=5.055 $Y=1.53 $X2=0
+ $Y2=0
cc_363 A1_N N_A_787_47#_c_1053_n 0.00959459f $X=5.215 $Y=1.105 $X2=0 $Y2=0
cc_364 N_A2_N_c_453_n N_A_211_297#_c_510_n 0.0051473f $X=4.545 $Y=1.16 $X2=0
+ $Y2=0
cc_365 N_A2_N_c_455_n N_VPWR_c_655_n 0.00300743f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_366 N_A2_N_c_456_n N_VPWR_c_655_n 0.00300743f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_367 N_A2_N_c_455_n N_VPWR_c_659_n 0.0053025f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_368 N_A2_N_c_456_n N_VPWR_c_661_n 0.0053025f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_369 N_A2_N_c_455_n N_VPWR_c_651_n 0.00697807f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_370 N_A2_N_c_456_n N_VPWR_c_651_n 0.00693014f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_371 N_A2_N_c_451_n N_VGND_c_941_n 0.00368123f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_372 N_A2_N_c_452_n N_VGND_c_941_n 0.00368123f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_373 N_A2_N_c_451_n N_VGND_c_948_n 0.00552518f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_374 N_A2_N_c_452_n N_VGND_c_948_n 0.00564339f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_375 N_A2_N_c_451_n N_A_787_47#_c_1055_n 0.00888424f $X=4.28 $Y=0.995 $X2=0
+ $Y2=0
cc_376 N_A2_N_c_452_n N_A_787_47#_c_1055_n 0.0105389f $X=4.8 $Y=0.995 $X2=0
+ $Y2=0
cc_377 N_A2_N_c_453_n N_A_787_47#_c_1055_n 0.00402166f $X=4.545 $Y=1.16 $X2=0
+ $Y2=0
cc_378 N_A_211_297#_c_514_n N_VPWR_M1014_s 0.00737637f $X=2.265 $Y=1.87 $X2=0
+ $Y2=0
cc_379 N_A_211_297#_c_508_n N_VPWR_M1011_d 0.00200003f $X=2.975 $Y=1.51 $X2=0
+ $Y2=0
cc_380 N_A_211_297#_c_510_n N_VPWR_M1011_d 0.00598364f $X=5.665 $Y=1.52 $X2=0
+ $Y2=0
cc_381 N_A_211_297#_c_510_n N_VPWR_M1026_d 0.00193338f $X=5.665 $Y=1.52 $X2=0
+ $Y2=0
cc_382 N_A_211_297#_c_514_n N_VPWR_c_654_n 0.0139109f $X=2.265 $Y=1.87 $X2=0
+ $Y2=0
cc_383 N_A_211_297#_c_504_n N_VPWR_c_656_n 0.00300743f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_384 N_A_211_297#_c_510_n N_VPWR_c_656_n 0.0080935f $X=5.665 $Y=1.52 $X2=0
+ $Y2=0
cc_385 N_A_211_297#_c_505_n N_VPWR_c_657_n 0.00300743f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_386 N_A_211_297#_c_506_n N_VPWR_c_657_n 0.00300743f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_387 N_A_211_297#_c_507_n N_VPWR_c_658_n 0.00479105f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_388 N_A_211_297#_c_504_n N_VPWR_c_663_n 0.00702461f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_389 N_A_211_297#_c_505_n N_VPWR_c_663_n 0.00702461f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_390 N_A_211_297#_c_506_n N_VPWR_c_665_n 0.00702461f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_391 N_A_211_297#_c_507_n N_VPWR_c_665_n 0.00702461f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_392 N_A_211_297#_M1001_d N_VPWR_c_651_n 0.00232092f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_393 N_A_211_297#_M1005_s N_VPWR_c_651_n 0.0024101f $X=2.465 $Y=1.485 $X2=0
+ $Y2=0
cc_394 N_A_211_297#_c_504_n N_VPWR_c_651_n 0.0124344f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_395 N_A_211_297#_c_505_n N_VPWR_c_651_n 0.00693457f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_396 N_A_211_297#_c_506_n N_VPWR_c_651_n 0.00693457f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_397 N_A_211_297#_c_507_n N_VPWR_c_651_n 0.0134606f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_398 N_A_211_297#_c_514_n N_VPWR_c_651_n 0.00856702f $X=2.265 $Y=1.87 $X2=0
+ $Y2=0
cc_399 N_A_211_297#_c_503_n N_VPWR_c_651_n 0.0205991f $X=2.61 $Y=1.96 $X2=0
+ $Y2=0
cc_400 N_A_211_297#_c_503_n N_VPWR_c_671_n 0.0181679f $X=2.61 $Y=1.96 $X2=0
+ $Y2=0
cc_401 N_A_211_297#_c_510_n N_VPWR_c_672_n 0.0108166f $X=5.665 $Y=1.52 $X2=0
+ $Y2=0
cc_402 N_A_211_297#_c_503_n N_VPWR_c_672_n 0.0220731f $X=2.61 $Y=1.96 $X2=0
+ $Y2=0
cc_403 N_A_211_297#_c_514_n N_A_117_297#_M1023_s 0.00367036f $X=2.265 $Y=1.87
+ $X2=0 $Y2=0
cc_404 N_A_211_297#_M1001_d N_A_117_297#_c_777_n 0.00352392f $X=1.055 $Y=1.485
+ $X2=0 $Y2=0
cc_405 N_A_211_297#_c_514_n N_A_117_297#_c_777_n 0.00608347f $X=2.265 $Y=1.87
+ $X2=0 $Y2=0
cc_406 N_A_211_297#_c_519_n N_A_117_297#_c_777_n 0.0127274f $X=1.2 $Y=1.87 $X2=0
+ $Y2=0
cc_407 N_A_211_297#_c_514_n N_A_117_297#_c_783_n 0.0130645f $X=2.265 $Y=1.87
+ $X2=0 $Y2=0
cc_408 N_A_211_297#_c_554_n N_X_M1003_d 0.00240549f $X=5.81 $Y=1.53 $X2=0 $Y2=0
cc_409 N_A_211_297#_c_509_n N_X_M1003_d 0.0025736f $X=5.81 $Y=1.53 $X2=0 $Y2=0
cc_410 N_A_211_297#_c_497_n N_X_c_803_n 0.00494802f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_411 N_A_211_297#_c_498_n N_X_c_803_n 0.0066581f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_412 N_A_211_297#_c_499_n N_X_c_803_n 5.38967e-19 $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_413 N_A_211_297#_c_505_n N_X_c_806_n 0.0133996f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_414 N_A_211_297#_c_506_n N_X_c_806_n 0.0134427f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_415 N_A_211_297#_c_600_p N_X_c_806_n 0.0164753f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_416 N_A_211_297#_c_502_n N_X_c_806_n 0.00503753f $X=7.125 $Y=1.202 $X2=0
+ $Y2=0
cc_417 N_A_211_297#_c_600_p N_X_c_810_n 0.00153327f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_418 N_A_211_297#_c_554_n N_X_c_810_n 0.00402205f $X=5.81 $Y=1.53 $X2=0 $Y2=0
cc_419 N_A_211_297#_c_509_n N_X_c_810_n 0.0116255f $X=5.81 $Y=1.53 $X2=0 $Y2=0
cc_420 N_A_211_297#_c_502_n N_X_c_810_n 0.00213176f $X=7.125 $Y=1.202 $X2=0
+ $Y2=0
cc_421 N_A_211_297#_c_498_n N_X_c_792_n 0.00901745f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_422 N_A_211_297#_c_499_n N_X_c_792_n 0.00901745f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_423 N_A_211_297#_c_600_p N_X_c_792_n 0.0392656f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_424 N_A_211_297#_c_502_n N_X_c_792_n 0.00345541f $X=7.125 $Y=1.202 $X2=0
+ $Y2=0
cc_425 N_A_211_297#_c_497_n N_X_c_793_n 0.002651f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_426 N_A_211_297#_c_498_n N_X_c_793_n 0.00116579f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_427 N_A_211_297#_c_553_n N_X_c_793_n 0.0226678f $X=6.005 $Y=1.16 $X2=0 $Y2=0
cc_428 N_A_211_297#_c_600_p N_X_c_793_n 0.00865078f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_429 N_A_211_297#_c_554_n N_X_c_793_n 9.68005e-19 $X=5.81 $Y=1.53 $X2=0 $Y2=0
cc_430 N_A_211_297#_c_502_n N_X_c_793_n 0.00357692f $X=7.125 $Y=1.202 $X2=0
+ $Y2=0
cc_431 N_A_211_297#_c_498_n N_X_c_824_n 5.19459e-19 $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_432 N_A_211_297#_c_499_n N_X_c_824_n 0.00633209f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_433 N_A_211_297#_c_500_n N_X_c_794_n 0.0140462f $X=7.15 $Y=0.995 $X2=0 $Y2=0
cc_434 N_A_211_297#_c_600_p N_X_c_794_n 0.00208021f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_435 N_A_211_297#_c_499_n N_X_c_795_n 0.00119508f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_436 N_A_211_297#_c_600_p N_X_c_795_n 0.0303261f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_437 N_A_211_297#_c_502_n N_X_c_795_n 0.00485798f $X=7.125 $Y=1.202 $X2=0
+ $Y2=0
cc_438 N_A_211_297#_c_506_n N_X_c_797_n 0.00188142f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_439 N_A_211_297#_c_507_n N_X_c_797_n 2.29143e-19 $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_440 N_A_211_297#_c_600_p N_X_c_797_n 0.0200073f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_441 N_A_211_297#_c_502_n N_X_c_797_n 0.00661719f $X=7.125 $Y=1.202 $X2=0
+ $Y2=0
cc_442 N_A_211_297#_c_500_n X 0.0182171f $X=7.15 $Y=0.995 $X2=0 $Y2=0
cc_443 N_A_211_297#_c_600_p X 0.00871662f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_444 N_A_211_297#_c_507_n X 0.0217101f $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_445 N_A_211_297#_c_600_p X 0.00495201f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_446 N_A_211_297#_c_502_n X 9.89874e-19 $X=7.125 $Y=1.202 $X2=0 $Y2=0
cc_447 N_A_211_297#_c_529_n N_A_27_47#_c_874_n 0.00727438f $X=2.61 $Y=0.73 $X2=0
+ $Y2=0
cc_448 N_A_211_297#_M1021_s N_A_27_47#_c_875_n 0.00399909f $X=2.425 $Y=0.235
+ $X2=0 $Y2=0
cc_449 N_A_211_297#_c_529_n N_A_27_47#_c_875_n 0.020134f $X=2.61 $Y=0.73 $X2=0
+ $Y2=0
cc_450 N_A_211_297#_c_503_n N_A_27_47#_c_875_n 0.00345006f $X=2.61 $Y=1.96 $X2=0
+ $Y2=0
cc_451 N_A_211_297#_c_497_n N_VGND_c_936_n 0.00275355f $X=5.69 $Y=0.995 $X2=0
+ $Y2=0
cc_452 N_A_211_297#_c_510_n N_VGND_c_936_n 0.00390271f $X=5.665 $Y=1.52 $X2=0
+ $Y2=0
cc_453 N_A_211_297#_c_498_n N_VGND_c_937_n 0.00410249f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_454 N_A_211_297#_c_499_n N_VGND_c_937_n 0.00276126f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_455 N_A_211_297#_c_500_n N_VGND_c_938_n 0.00438629f $X=7.15 $Y=0.995 $X2=0
+ $Y2=0
cc_456 N_A_211_297#_c_497_n N_VGND_c_943_n 0.00542163f $X=5.69 $Y=0.995 $X2=0
+ $Y2=0
cc_457 N_A_211_297#_c_498_n N_VGND_c_943_n 0.00424138f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_458 N_A_211_297#_c_499_n N_VGND_c_945_n 0.00424138f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_459 N_A_211_297#_c_500_n N_VGND_c_945_n 0.00437852f $X=7.15 $Y=0.995 $X2=0
+ $Y2=0
cc_460 N_A_211_297#_M1021_s N_VGND_c_948_n 0.00256987f $X=2.425 $Y=0.235 $X2=0
+ $Y2=0
cc_461 N_A_211_297#_c_497_n N_VGND_c_948_n 0.00965669f $X=5.69 $Y=0.995 $X2=0
+ $Y2=0
cc_462 N_A_211_297#_c_498_n N_VGND_c_948_n 0.00609398f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_463 N_A_211_297#_c_499_n N_VGND_c_948_n 0.00608656f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_464 N_A_211_297#_c_500_n N_VGND_c_948_n 0.00722755f $X=7.15 $Y=0.995 $X2=0
+ $Y2=0
cc_465 N_A_211_297#_c_510_n N_A_787_47#_c_1053_n 0.00144574f $X=5.665 $Y=1.52
+ $X2=0 $Y2=0
cc_466 N_VPWR_c_651_n N_A_117_297#_M1009_d 0.00297222f $X=7.59 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_467 N_VPWR_c_651_n N_A_117_297#_M1023_s 0.00241598f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_468 N_VPWR_c_667_n N_A_117_297#_c_777_n 0.0386815f $X=2.015 $Y=2.72 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_651_n N_A_117_297#_c_777_n 0.0239184f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_667_n N_A_117_297#_c_788_n 0.015002f $X=2.015 $Y=2.72 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_651_n N_A_117_297#_c_788_n 0.00962794f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_472 N_VPWR_c_667_n N_A_117_297#_c_783_n 0.0143006f $X=2.015 $Y=2.72 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_651_n N_A_117_297#_c_783_n 0.00938288f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_474 N_VPWR_c_651_n N_X_M1003_d 0.0031047f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_475 N_VPWR_c_651_n N_X_M1015_d 0.0031047f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_476 N_VPWR_c_663_n N_X_c_842_n 0.0149311f $X=6.295 $Y=2.72 $X2=0 $Y2=0
cc_477 N_VPWR_c_651_n N_X_c_842_n 0.00955092f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_478 N_VPWR_M1012_s N_X_c_806_n 0.0047345f $X=6.275 $Y=1.485 $X2=0 $Y2=0
cc_479 N_VPWR_c_657_n N_X_c_806_n 0.011587f $X=6.42 $Y=2.33 $X2=0 $Y2=0
cc_480 N_VPWR_c_651_n N_X_c_806_n 0.0142452f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_481 N_VPWR_c_665_n N_X_c_847_n 0.0149311f $X=7.235 $Y=2.72 $X2=0 $Y2=0
cc_482 N_VPWR_c_651_n N_X_c_847_n 0.00955092f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_483 N_VPWR_M1024_s X 0.00150236f $X=7.215 $Y=1.485 $X2=0 $Y2=0
cc_484 N_VPWR_c_658_n X 0.0110395f $X=7.36 $Y=1.99 $X2=0 $Y2=0
cc_485 N_VPWR_M1024_s N_X_c_800_n 0.001627f $X=7.215 $Y=1.485 $X2=0 $Y2=0
cc_486 N_VPWR_c_658_n N_X_c_800_n 0.00712278f $X=7.36 $Y=1.99 $X2=0 $Y2=0
cc_487 N_X_c_792_n N_VGND_M1007_s 0.00251047f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_488 N_X_c_794_n N_VGND_M1020_s 0.00320332f $X=7.405 $Y=0.815 $X2=0 $Y2=0
cc_489 N_X_c_793_n N_VGND_c_936_n 0.00750114f $X=6.115 $Y=0.815 $X2=0 $Y2=0
cc_490 N_X_c_803_n N_VGND_c_937_n 0.0171386f $X=5.95 $Y=0.39 $X2=0 $Y2=0
cc_491 N_X_c_792_n N_VGND_c_937_n 0.0127273f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_492 N_X_c_794_n N_VGND_c_938_n 0.013002f $X=7.405 $Y=0.815 $X2=0 $Y2=0
cc_493 N_X_c_803_n N_VGND_c_943_n 0.0198028f $X=5.95 $Y=0.39 $X2=0 $Y2=0
cc_494 N_X_c_792_n N_VGND_c_943_n 0.00266636f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_495 N_X_c_792_n N_VGND_c_945_n 0.00198695f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_496 N_X_c_824_n N_VGND_c_945_n 0.0205249f $X=6.89 $Y=0.39 $X2=0 $Y2=0
cc_497 N_X_c_794_n N_VGND_c_945_n 0.00254521f $X=7.405 $Y=0.815 $X2=0 $Y2=0
cc_498 N_X_c_794_n N_VGND_c_947_n 0.004465f $X=7.405 $Y=0.815 $X2=0 $Y2=0
cc_499 N_X_M1002_d N_VGND_c_948_n 0.00256339f $X=5.765 $Y=0.235 $X2=0 $Y2=0
cc_500 N_X_M1008_d N_VGND_c_948_n 0.00305225f $X=6.705 $Y=0.235 $X2=0 $Y2=0
cc_501 N_X_c_803_n N_VGND_c_948_n 0.0139751f $X=5.95 $Y=0.39 $X2=0 $Y2=0
cc_502 N_X_c_792_n N_VGND_c_948_n 0.00972452f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_503 N_X_c_824_n N_VGND_c_948_n 0.0141809f $X=6.89 $Y=0.39 $X2=0 $Y2=0
cc_504 N_X_c_794_n N_VGND_c_948_n 0.013148f $X=7.405 $Y=0.815 $X2=0 $Y2=0
cc_505 N_A_27_47#_c_872_n N_VGND_M1017_d 0.00162089f $X=0.985 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_506 N_A_27_47#_c_874_n N_VGND_M1027_s 0.00255557f $X=1.925 $Y=0.82 $X2=0
+ $Y2=0
cc_507 N_A_27_47#_c_872_n N_VGND_c_932_n 0.0122559f $X=0.985 $Y=0.815 $X2=0
+ $Y2=0
cc_508 N_A_27_47#_c_872_n N_VGND_c_933_n 0.00198695f $X=0.985 $Y=0.815 $X2=0
+ $Y2=0
cc_509 N_A_27_47#_c_883_n N_VGND_c_933_n 0.0231806f $X=1.2 $Y=0.39 $X2=0 $Y2=0
cc_510 N_A_27_47#_c_874_n N_VGND_c_933_n 0.00248202f $X=1.925 $Y=0.82 $X2=0
+ $Y2=0
cc_511 N_A_27_47#_c_874_n N_VGND_c_934_n 0.012101f $X=1.925 $Y=0.82 $X2=0 $Y2=0
cc_512 N_A_27_47#_c_888_n N_VGND_c_934_n 0.0172916f $X=2.075 $Y=0.475 $X2=0
+ $Y2=0
cc_513 N_A_27_47#_c_889_n N_VGND_c_934_n 0.00582645f $X=2.14 $Y=0.73 $X2=0 $Y2=0
cc_514 N_A_27_47#_c_875_n N_VGND_c_935_n 0.0130087f $X=3.08 $Y=0.39 $X2=0 $Y2=0
cc_515 N_A_27_47#_c_874_n N_VGND_c_939_n 0.00194552f $X=1.925 $Y=0.82 $X2=0
+ $Y2=0
cc_516 N_A_27_47#_c_888_n N_VGND_c_939_n 0.0186086f $X=2.075 $Y=0.475 $X2=0
+ $Y2=0
cc_517 N_A_27_47#_c_875_n N_VGND_c_939_n 0.0587424f $X=3.08 $Y=0.39 $X2=0 $Y2=0
cc_518 N_A_27_47#_M1017_s N_VGND_c_948_n 0.00258952f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_519 N_A_27_47#_M1006_d N_VGND_c_948_n 0.00304426f $X=1.015 $Y=0.235 $X2=0
+ $Y2=0
cc_520 N_A_27_47#_M1018_s N_VGND_c_948_n 0.00215206f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_521 N_A_27_47#_M1022_d N_VGND_c_948_n 0.00250339f $X=2.895 $Y=0.235 $X2=0
+ $Y2=0
cc_522 N_A_27_47#_c_871_n N_VGND_c_948_n 0.0126169f $X=0.26 $Y=0.39 $X2=0 $Y2=0
cc_523 N_A_27_47#_c_872_n N_VGND_c_948_n 0.0094839f $X=0.985 $Y=0.815 $X2=0
+ $Y2=0
cc_524 N_A_27_47#_c_883_n N_VGND_c_948_n 0.0143352f $X=1.2 $Y=0.39 $X2=0 $Y2=0
cc_525 N_A_27_47#_c_874_n N_VGND_c_948_n 0.0096764f $X=1.925 $Y=0.82 $X2=0 $Y2=0
cc_526 N_A_27_47#_c_888_n N_VGND_c_948_n 0.0111017f $X=2.075 $Y=0.475 $X2=0
+ $Y2=0
cc_527 N_A_27_47#_c_875_n N_VGND_c_948_n 0.0366908f $X=3.08 $Y=0.39 $X2=0 $Y2=0
cc_528 N_A_27_47#_c_871_n N_VGND_c_949_n 0.0217962f $X=0.26 $Y=0.39 $X2=0 $Y2=0
cc_529 N_A_27_47#_c_872_n N_VGND_c_949_n 0.00254521f $X=0.985 $Y=0.815 $X2=0
+ $Y2=0
cc_530 N_VGND_c_948_n N_A_787_47#_M1000_d 0.00218617f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_531 N_VGND_c_948_n N_A_787_47#_M1025_d 0.00325021f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_532 N_VGND_c_935_n N_A_787_47#_c_1055_n 0.0132045f $X=3.6 $Y=0.39 $X2=0 $Y2=0
cc_533 N_VGND_c_941_n N_A_787_47#_c_1055_n 0.0450213f $X=5.395 $Y=0 $X2=0 $Y2=0
cc_534 N_VGND_c_948_n N_A_787_47#_c_1055_n 0.0366514f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_535 N_VGND_c_941_n N_A_787_47#_c_1072_n 0.0120493f $X=5.395 $Y=0 $X2=0 $Y2=0
cc_536 N_VGND_c_948_n N_A_787_47#_c_1072_n 0.00934683f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_537 N_VGND_c_936_n N_A_787_47#_c_1053_n 5.82165e-19 $X=5.48 $Y=0.39 $X2=0
+ $Y2=0
