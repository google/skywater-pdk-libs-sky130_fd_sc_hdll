* File: sky130_fd_sc_hdll__o2bb2ai_1.spice
* Created: Wed Sep  2 08:46:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o2bb2ai_1.pex.spice"
.subckt sky130_fd_sc_hdll__o2bb2ai_1  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1006 A_122_47# N_A1_N_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.21125 PD=0.92 PS=1.95 NRD=14.76 NRS=11.076 M=1 R=4.33333
+ SA=75000.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1004 N_A_120_297#_M1004_d N_A2_N_M1004_g A_122_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=14.76 M=1 R=4.33333 SA=75000.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_A_396_47#_M1005_d N_A_120_297#_M1005_g N_Y_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.1105 AS=0.1755 PD=0.99 PS=1.84 NRD=11.988 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_B2_M1009_g N_A_396_47#_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.1105 PD=0.92 PS=0.99 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1001 N_A_396_47#_M1001_d N_B1_M1001_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_A_120_297#_M1000_d N_A1_N_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.285 PD=1.29 PS=2.57 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A2_N_M1008_g N_A_120_297#_M1000_d VPB PHIGHVT L=0.18 W=1
+ AD=0.36 AS=0.145 PD=1.72 PS=1.29 NRD=8.8453 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90002 A=0.18 P=2.36 MULT=1
MM1002 N_Y_M1002_d N_A_120_297#_M1002_g N_VPWR_M1008_d VPB PHIGHVT L=0.18 W=1
+ AD=0.155 AS=0.36 PD=1.31 PS=1.72 NRD=0.9653 NRS=8.8453 M=1 R=5.55556
+ SA=90001.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1007 A_492_297# N_B2_M1007_g N_Y_M1002_d VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.155 PD=1.29 PS=1.31 NRD=17.7103 NRS=4.9053 M=1 R=5.55556 SA=90002.1
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_B1_M1003_g A_492_297# VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=17.7103 M=1 R=5.55556 SA=90002.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hdll__o2bb2ai_1.pxi.spice"
*
.ends
*
*
