* File: sky130_fd_sc_hdll__nor4_6.pxi.spice
* Created: Wed Sep  2 08:41:19 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR4_6%A N_A_c_166_n N_A_M1000_g N_A_c_159_n N_A_M1006_g
+ N_A_c_160_n N_A_M1011_g N_A_c_167_n N_A_M1005_g N_A_c_168_n N_A_M1014_g
+ N_A_c_161_n N_A_M1019_g N_A_c_162_n N_A_M1021_g N_A_c_169_n N_A_M1020_g
+ N_A_c_170_n N_A_M1030_g N_A_c_163_n N_A_M1026_g N_A_c_164_n N_A_M1034_g
+ N_A_c_171_n N_A_M1042_g A N_A_c_175_p N_A_c_165_n
+ PM_SKY130_FD_SC_HDLL__NOR4_6%A
x_PM_SKY130_FD_SC_HDLL__NOR4_6%B N_B_c_272_n N_B_M1009_g N_B_c_265_n N_B_M1003_g
+ N_B_c_266_n N_B_M1008_g N_B_c_273_n N_B_M1017_g N_B_c_274_n N_B_M1024_g
+ N_B_c_267_n N_B_M1012_g N_B_c_268_n N_B_M1022_g N_B_c_275_n N_B_M1033_g
+ N_B_c_276_n N_B_M1035_g N_B_c_269_n N_B_M1036_g N_B_c_270_n N_B_M1046_g
+ N_B_c_277_n N_B_M1040_g B N_B_c_281_n N_B_c_271_n
+ PM_SKY130_FD_SC_HDLL__NOR4_6%B
x_PM_SKY130_FD_SC_HDLL__NOR4_6%C N_C_c_384_n N_C_M1001_g N_C_c_377_n N_C_M1010_g
+ N_C_c_378_n N_C_M1013_g N_C_c_385_n N_C_M1007_g N_C_c_386_n N_C_M1015_g
+ N_C_c_379_n N_C_M1028_g N_C_c_380_n N_C_M1038_g N_C_c_387_n N_C_M1016_g
+ N_C_c_388_n N_C_M1043_g N_C_c_381_n N_C_M1039_g N_C_c_382_n N_C_M1044_g
+ N_C_c_389_n N_C_M1045_g C N_C_c_393_p N_C_c_383_n C
+ PM_SKY130_FD_SC_HDLL__NOR4_6%C
x_PM_SKY130_FD_SC_HDLL__NOR4_6%D N_D_c_497_n N_D_M1002_g N_D_c_489_n N_D_M1004_g
+ N_D_c_490_n N_D_M1023_g N_D_c_498_n N_D_M1018_g N_D_c_499_n N_D_M1027_g
+ N_D_c_491_n N_D_M1025_g N_D_c_492_n N_D_M1032_g N_D_c_500_n N_D_M1029_g
+ N_D_c_501_n N_D_M1031_g N_D_c_493_n N_D_M1041_g N_D_c_494_n N_D_M1047_g
+ N_D_c_502_n N_D_M1037_g D N_D_c_495_n N_D_c_496_n
+ PM_SKY130_FD_SC_HDLL__NOR4_6%D
x_PM_SKY130_FD_SC_HDLL__NOR4_6%A_27_297# N_A_27_297#_M1000_s N_A_27_297#_M1005_s
+ N_A_27_297#_M1020_s N_A_27_297#_M1042_s N_A_27_297#_M1017_d
+ N_A_27_297#_M1033_d N_A_27_297#_M1040_d N_A_27_297#_c_604_n
+ N_A_27_297#_c_605_n N_A_27_297#_c_606_n N_A_27_297#_c_641_p
+ N_A_27_297#_c_607_n N_A_27_297#_c_643_p N_A_27_297#_c_608_n
+ N_A_27_297#_c_609_n N_A_27_297#_c_645_p N_A_27_297#_c_631_n
+ N_A_27_297#_c_673_p N_A_27_297#_c_633_n N_A_27_297#_c_677_p
+ N_A_27_297#_c_610_n N_A_27_297#_c_611_n N_A_27_297#_c_612_n
+ N_A_27_297#_c_613_n N_A_27_297#_c_649_p N_A_27_297#_c_650_p
+ PM_SKY130_FD_SC_HDLL__NOR4_6%A_27_297#
x_PM_SKY130_FD_SC_HDLL__NOR4_6%VPWR N_VPWR_M1000_d N_VPWR_M1014_d N_VPWR_M1030_d
+ N_VPWR_c_693_n N_VPWR_c_694_n N_VPWR_c_695_n N_VPWR_c_696_n N_VPWR_c_697_n
+ VPWR N_VPWR_c_698_n N_VPWR_c_692_n N_VPWR_c_700_n N_VPWR_c_701_n
+ N_VPWR_c_702_n VPWR PM_SKY130_FD_SC_HDLL__NOR4_6%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR4_6%A_685_297# N_A_685_297#_M1009_s
+ N_A_685_297#_M1024_s N_A_685_297#_M1035_s N_A_685_297#_M1001_s
+ N_A_685_297#_M1015_s N_A_685_297#_M1043_s N_A_685_297#_c_830_n
+ N_A_685_297#_c_831_n N_A_685_297#_c_832_n N_A_685_297#_c_833_n
+ N_A_685_297#_c_834_n N_A_685_297#_c_835_n N_A_685_297#_c_836_n
+ N_A_685_297#_c_837_n N_A_685_297#_c_838_n N_A_685_297#_c_839_n
+ N_A_685_297#_c_840_n PM_SKY130_FD_SC_HDLL__NOR4_6%A_685_297#
x_PM_SKY130_FD_SC_HDLL__NOR4_6%A_1263_297# N_A_1263_297#_M1001_d
+ N_A_1263_297#_M1007_d N_A_1263_297#_M1016_d N_A_1263_297#_M1045_d
+ N_A_1263_297#_M1018_s N_A_1263_297#_M1029_s N_A_1263_297#_M1037_s
+ N_A_1263_297#_c_920_n N_A_1263_297#_c_925_n N_A_1263_297#_c_921_n
+ N_A_1263_297#_c_983_n N_A_1263_297#_c_927_n N_A_1263_297#_c_988_n
+ N_A_1263_297#_c_929_n N_A_1263_297#_c_922_n N_A_1263_297#_c_933_n
+ N_A_1263_297#_c_999_p N_A_1263_297#_c_935_n N_A_1263_297#_c_1003_p
+ N_A_1263_297#_c_937_n N_A_1263_297#_c_923_n N_A_1263_297#_c_924_n
+ N_A_1263_297#_c_965_n N_A_1263_297#_c_967_n N_A_1263_297#_c_969_n
+ N_A_1263_297#_c_971_n N_A_1263_297#_c_973_n
+ PM_SKY130_FD_SC_HDLL__NOR4_6%A_1263_297#
x_PM_SKY130_FD_SC_HDLL__NOR4_6%Y N_Y_M1006_s N_Y_M1019_s N_Y_M1026_s N_Y_M1003_s
+ N_Y_M1012_s N_Y_M1036_s N_Y_M1010_s N_Y_M1028_s N_Y_M1039_s N_Y_M1004_d
+ N_Y_M1025_d N_Y_M1041_d N_Y_M1002_d N_Y_M1027_d N_Y_M1031_d N_Y_c_1037_n
+ N_Y_c_1011_n N_Y_c_1012_n N_Y_c_1048_n N_Y_c_1013_n N_Y_c_1056_n N_Y_c_1014_n
+ N_Y_c_1062_n N_Y_c_1015_n N_Y_c_1082_n N_Y_c_1016_n N_Y_c_1090_n N_Y_c_1017_n
+ N_Y_c_1111_n N_Y_c_1018_n N_Y_c_1118_n N_Y_c_1019_n N_Y_c_1126_n N_Y_c_1020_n
+ N_Y_c_1132_n N_Y_c_1033_n N_Y_c_1021_n N_Y_c_1160_n N_Y_c_1034_n N_Y_c_1022_n
+ N_Y_c_1172_n N_Y_c_1023_n N_Y_c_1024_n N_Y_c_1025_n N_Y_c_1026_n N_Y_c_1027_n
+ N_Y_c_1028_n N_Y_c_1029_n N_Y_c_1030_n N_Y_c_1031_n N_Y_c_1035_n N_Y_c_1032_n
+ N_Y_c_1036_n N_Y_c_1188_n N_Y_c_1190_n Y PM_SKY130_FD_SC_HDLL__NOR4_6%Y
x_PM_SKY130_FD_SC_HDLL__NOR4_6%VGND N_VGND_M1006_d N_VGND_M1011_d N_VGND_M1021_d
+ N_VGND_M1034_d N_VGND_M1008_d N_VGND_M1022_d N_VGND_M1046_d N_VGND_M1013_d
+ N_VGND_M1038_d N_VGND_M1044_d N_VGND_M1023_s N_VGND_M1032_s N_VGND_M1047_s
+ N_VGND_c_1318_n N_VGND_c_1319_n N_VGND_c_1320_n N_VGND_c_1321_n
+ N_VGND_c_1322_n N_VGND_c_1323_n N_VGND_c_1324_n N_VGND_c_1325_n
+ N_VGND_c_1326_n N_VGND_c_1327_n N_VGND_c_1328_n N_VGND_c_1329_n
+ N_VGND_c_1330_n N_VGND_c_1331_n N_VGND_c_1332_n N_VGND_c_1333_n
+ N_VGND_c_1334_n N_VGND_c_1335_n N_VGND_c_1336_n N_VGND_c_1337_n
+ N_VGND_c_1338_n N_VGND_c_1339_n N_VGND_c_1340_n N_VGND_c_1341_n
+ N_VGND_c_1342_n N_VGND_c_1343_n N_VGND_c_1344_n N_VGND_c_1345_n
+ N_VGND_c_1346_n N_VGND_c_1347_n VGND N_VGND_c_1348_n N_VGND_c_1349_n
+ N_VGND_c_1350_n N_VGND_c_1351_n N_VGND_c_1352_n N_VGND_c_1353_n
+ N_VGND_c_1354_n N_VGND_c_1355_n PM_SKY130_FD_SC_HDLL__NOR4_6%VGND
cc_1 VNB N_A_c_159_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_2 VNB N_A_c_160_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_3 VNB N_A_c_161_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=0.995
cc_4 VNB N_A_c_162_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=0.995
cc_5 VNB N_A_c_163_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=2.42 $Y2=0.995
cc_6 VNB N_A_c_164_n 0.0168874f $X=-0.19 $Y=-0.24 $X2=2.84 $Y2=0.995
cc_7 VNB N_A_c_165_n 0.126213f $X=-0.19 $Y=-0.24 $X2=2.84 $Y2=1.202
cc_8 VNB N_B_c_265_n 0.0168874f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_9 VNB N_B_c_266_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_10 VNB N_B_c_267_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=0.995
cc_11 VNB N_B_c_268_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=0.995
cc_12 VNB N_B_c_269_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=2.42 $Y2=0.995
cc_13 VNB N_B_c_270_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=2.84 $Y2=0.995
cc_14 VNB N_B_c_271_n 0.124727f $X=-0.19 $Y=-0.24 $X2=2.84 $Y2=1.202
cc_15 VNB N_C_c_377_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_16 VNB N_C_c_378_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_17 VNB N_C_c_379_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=0.995
cc_18 VNB N_C_c_380_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=0.995
cc_19 VNB N_C_c_381_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=2.42 $Y2=0.995
cc_20 VNB N_C_c_382_n 0.0168874f $X=-0.19 $Y=-0.24 $X2=2.84 $Y2=0.995
cc_21 VNB N_C_c_383_n 0.124713f $X=-0.19 $Y=-0.24 $X2=2.84 $Y2=1.202
cc_22 VNB N_D_c_489_n 0.0168874f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_23 VNB N_D_c_490_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_24 VNB N_D_c_491_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=0.995
cc_25 VNB N_D_c_492_n 0.0166924f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=0.995
cc_26 VNB N_D_c_493_n 0.0163356f $X=-0.19 $Y=-0.24 $X2=2.42 $Y2=0.995
cc_27 VNB N_D_c_494_n 0.0209805f $X=-0.19 $Y=-0.24 $X2=2.84 $Y2=0.995
cc_28 VNB N_D_c_495_n 0.00174962f $X=-0.19 $Y=-0.24 $X2=2.71 $Y2=1.202
cc_29 VNB N_D_c_496_n 0.125306f $X=-0.19 $Y=-0.24 $X2=2.84 $Y2=1.202
cc_30 VNB N_VPWR_c_692_n 0.516438f $X=-0.19 $Y=-0.24 $X2=2.865 $Y2=1.985
cc_31 VNB N_Y_c_1011_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=2.395 $Y2=1.202
cc_32 VNB N_Y_c_1012_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=2.42 $Y2=1.202
cc_33 VNB N_Y_c_1013_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=2.865 $Y2=1.202
cc_34 VNB N_Y_c_1014_n 0.005207f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_Y_c_1015_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_Y_c_1016_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_Y_c_1017_n 0.0132852f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_Y_c_1018_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_Y_c_1019_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_Y_c_1020_n 0.00528638f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_Y_c_1021_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_Y_c_1022_n 0.00344273f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_Y_c_1023_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_Y_c_1024_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_Y_c_1025_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_Y_c_1026_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_Y_c_1027_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_Y_c_1028_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_Y_c_1029_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_Y_c_1030_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_Y_c_1031_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_Y_c_1032_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_1318_n 0.0116364f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.202
cc_54 VNB N_VGND_c_1319_n 0.0348682f $X=-0.19 $Y=-0.24 $X2=0.67 $Y2=1.16
cc_55 VNB N_VGND_c_1320_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=1.202
cc_56 VNB N_VGND_c_1321_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=1.202
cc_57 VNB N_VGND_c_1322_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=2.395 $Y2=1.202
cc_58 VNB N_VGND_c_1323_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=2.71 $Y2=1.16
cc_59 VNB N_VGND_c_1324_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=2.865 $Y2=1.202
cc_60 VNB N_VGND_c_1325_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1326_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1327_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1328_n 0.00413904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1329_n 0.00413904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1330_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1331_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1332_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1333_n 0.00466649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1334_n 0.0122696f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1335_n 0.0338006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1336_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1337_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1338_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1339_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1340_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1341_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1342_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1343_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1344_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1345_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1346_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1347_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1348_n 0.0186336f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1349_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1350_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1351_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1352_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1353_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1354_n 0.0222052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1355_n 0.564485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VPB N_A_c_166_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_92 VPB N_A_c_167_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_93 VPB N_A_c_168_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_94 VPB N_A_c_169_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_95 VPB N_A_c_170_n 0.0159747f $X=-0.19 $Y=1.305 $X2=2.395 $Y2=1.41
cc_96 VPB N_A_c_171_n 0.0161064f $X=-0.19 $Y=1.305 $X2=2.865 $Y2=1.41
cc_97 VPB N_A_c_165_n 0.0742474f $X=-0.19 $Y=1.305 $X2=2.84 $Y2=1.202
cc_98 VPB N_B_c_272_n 0.0164231f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_99 VPB N_B_c_273_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_100 VPB N_B_c_274_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_101 VPB N_B_c_275_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_102 VPB N_B_c_276_n 0.0159747f $X=-0.19 $Y=1.305 $X2=2.395 $Y2=1.41
cc_103 VPB N_B_c_277_n 0.0203443f $X=-0.19 $Y=1.305 $X2=2.865 $Y2=1.41
cc_104 VPB N_B_c_271_n 0.0751311f $X=-0.19 $Y=1.305 $X2=2.84 $Y2=1.202
cc_105 VPB N_C_c_384_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_106 VPB N_C_c_385_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_107 VPB N_C_c_386_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_108 VPB N_C_c_387_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_109 VPB N_C_c_388_n 0.0159747f $X=-0.19 $Y=1.305 $X2=2.395 $Y2=1.41
cc_110 VPB N_C_c_389_n 0.0164231f $X=-0.19 $Y=1.305 $X2=2.865 $Y2=1.41
cc_111 VPB N_C_c_383_n 0.0751311f $X=-0.19 $Y=1.305 $X2=2.84 $Y2=1.202
cc_112 VPB N_D_c_497_n 0.0164231f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_113 VPB N_D_c_498_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_114 VPB N_D_c_499_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_115 VPB N_D_c_500_n 0.0159542f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_116 VPB N_D_c_501_n 0.015773f $X=-0.19 $Y=1.305 $X2=2.395 $Y2=1.41
cc_117 VPB N_D_c_502_n 0.0199561f $X=-0.19 $Y=1.305 $X2=2.865 $Y2=1.41
cc_118 VPB N_D_c_496_n 0.0757423f $X=-0.19 $Y=1.305 $X2=2.84 $Y2=1.202
cc_119 VPB N_A_27_297#_c_604_n 0.0116935f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_120 VPB N_A_27_297#_c_605_n 0.0315052f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.985
cc_121 VPB N_A_27_297#_c_606_n 0.00203429f $X=-0.19 $Y=1.305 $X2=2.395 $Y2=1.985
cc_122 VPB N_A_27_297#_c_607_n 0.00193318f $X=-0.19 $Y=1.305 $X2=2.84 $Y2=0.56
cc_123 VPB N_A_27_297#_c_608_n 0.00204701f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_27_297#_c_609_n 0.00416602f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.202
cc_125 VPB N_A_27_297#_c_610_n 0.00180756f $X=-0.19 $Y=1.305 $X2=2.71 $Y2=1.16
cc_126 VPB N_A_27_297#_c_611_n 0.00482315f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_27_297#_c_612_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_27_297#_c_613_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_693_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.985
cc_130 VPB N_VPWR_c_694_n 0.0195604f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=0.995
cc_131 VPB N_VPWR_c_695_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=0.56
cc_132 VPB N_VPWR_c_696_n 0.0195604f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_133 VPB N_VPWR_c_697_n 0.00516582f $X=-0.19 $Y=1.305 $X2=2.395 $Y2=1.985
cc_134 VPB N_VPWR_c_698_n 0.221759f $X=-0.19 $Y=1.305 $X2=2.865 $Y2=1.985
cc_135 VPB N_VPWR_c_692_n 0.0578198f $X=-0.19 $Y=1.305 $X2=2.865 $Y2=1.985
cc_136 VPB N_VPWR_c_700_n 0.0241054f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_137 VPB N_VPWR_c_701_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.67 $Y2=1.16
cc_138 VPB N_VPWR_c_702_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_139 VPB N_A_685_297#_c_830_n 0.00193318f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=0.56
cc_140 VPB N_A_685_297#_c_831_n 0.00193318f $X=-0.19 $Y=1.305 $X2=2.395 $Y2=1.41
cc_141 VPB N_A_685_297#_c_832_n 0.0215869f $X=-0.19 $Y=1.305 $X2=2.42 $Y2=0.56
cc_142 VPB N_A_685_297#_c_833_n 0.00193318f $X=-0.19 $Y=1.305 $X2=2.84 $Y2=0.56
cc_143 VPB N_A_685_297#_c_834_n 0.00193318f $X=-0.19 $Y=1.305 $X2=1.525
+ $Y2=1.105
cc_144 VPB N_A_685_297#_c_835_n 0.00174485f $X=-0.19 $Y=1.305 $X2=0.67 $Y2=1.16
cc_145 VPB N_A_685_297#_c_836_n 0.00149756f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.202
cc_146 VPB N_A_685_297#_c_837_n 0.00149756f $X=-0.19 $Y=1.305 $X2=1.455
+ $Y2=1.202
cc_147 VPB N_A_685_297#_c_838_n 0.00149756f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=1.202
cc_148 VPB N_A_685_297#_c_839_n 0.00149756f $X=-0.19 $Y=1.305 $X2=2.395
+ $Y2=1.202
cc_149 VPB N_A_685_297#_c_840_n 0.00175152f $X=-0.19 $Y=1.305 $X2=2.71 $Y2=1.202
cc_150 VPB N_A_1263_297#_c_920_n 0.00482315f $X=-0.19 $Y=1.305 $X2=1.925
+ $Y2=1.985
cc_151 VPB N_A_1263_297#_c_921_n 0.00180756f $X=-0.19 $Y=1.305 $X2=2.395
+ $Y2=1.985
cc_152 VPB N_A_1263_297#_c_922_n 0.00442576f $X=-0.19 $Y=1.305 $X2=0.67 $Y2=1.16
cc_153 VPB N_A_1263_297#_c_923_n 0.00719505f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_1263_297#_c_924_n 0.0351112f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_Y_c_1033_n 0.00193318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_Y_c_1034_n 0.00222931f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_Y_c_1035_n 0.00175152f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_Y_c_1036_n 0.00149756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 N_A_c_171_n N_B_c_272_n 0.00971598f $X=2.865 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_160 N_A_c_164_n N_B_c_265_n 0.0179509f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_c_175_p N_B_c_281_n 0.00795414f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A_c_165_n N_B_c_281_n 8.31714e-19 $X=2.84 $Y=1.202 $X2=0 $Y2=0
cc_163 N_A_c_175_p N_B_c_271_n 8.31714e-19 $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A_c_165_n N_B_c_271_n 0.0237215f $X=2.84 $Y=1.202 $X2=0 $Y2=0
cc_165 N_A_c_166_n N_A_27_297#_c_606_n 0.0181833f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_c_167_n N_A_27_297#_c_606_n 0.0156273f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_c_175_p N_A_27_297#_c_606_n 0.0417725f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A_c_165_n N_A_27_297#_c_606_n 0.00871881f $X=2.84 $Y=1.202 $X2=0 $Y2=0
cc_169 N_A_c_168_n N_A_27_297#_c_607_n 0.0156273f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_c_169_n N_A_27_297#_c_607_n 0.0156273f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_c_175_p N_A_27_297#_c_607_n 0.0486996f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A_c_165_n N_A_27_297#_c_607_n 0.00885494f $X=2.84 $Y=1.202 $X2=0 $Y2=0
cc_173 N_A_c_170_n N_A_27_297#_c_608_n 0.0156273f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_c_171_n N_A_27_297#_c_608_n 0.0164448f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_c_175_p N_A_27_297#_c_608_n 0.0417725f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A_c_165_n N_A_27_297#_c_608_n 0.00859761f $X=2.84 $Y=1.202 $X2=0 $Y2=0
cc_177 N_A_c_175_p N_A_27_297#_c_612_n 0.0204509f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_c_165_n N_A_27_297#_c_612_n 0.00635938f $X=2.84 $Y=1.202 $X2=0 $Y2=0
cc_179 N_A_c_175_p N_A_27_297#_c_613_n 0.0204509f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_c_165_n N_A_27_297#_c_613_n 0.00635938f $X=2.84 $Y=1.202 $X2=0 $Y2=0
cc_181 N_A_c_166_n N_VPWR_c_693_n 0.00300743f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A_c_167_n N_VPWR_c_693_n 0.00300743f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A_c_167_n N_VPWR_c_694_n 0.00702461f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A_c_168_n N_VPWR_c_694_n 0.00702461f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A_c_168_n N_VPWR_c_695_n 0.00300743f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_186 N_A_c_169_n N_VPWR_c_695_n 0.00300743f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_187 N_A_c_169_n N_VPWR_c_696_n 0.00702461f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A_c_170_n N_VPWR_c_696_n 0.00702461f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A_c_170_n N_VPWR_c_697_n 0.00300743f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_190 N_A_c_171_n N_VPWR_c_697_n 0.00300743f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_191 N_A_c_171_n N_VPWR_c_698_n 0.00702461f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_192 N_A_c_166_n N_VPWR_c_692_n 0.0133387f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A_c_167_n N_VPWR_c_692_n 0.0124092f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A_c_168_n N_VPWR_c_692_n 0.0124092f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A_c_169_n N_VPWR_c_692_n 0.0124092f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A_c_170_n N_VPWR_c_692_n 0.0124092f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A_c_171_n N_VPWR_c_692_n 0.0124344f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_c_166_n N_VPWR_c_700_n 0.00702461f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A_c_159_n N_Y_c_1037_n 0.00539651f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_c_160_n N_Y_c_1037_n 0.00671723f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_c_161_n N_Y_c_1037_n 5.24636e-19 $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_c_160_n N_Y_c_1011_n 0.00929182f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A_c_161_n N_Y_c_1011_n 0.00929182f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A_c_175_p N_Y_c_1011_n 0.0435408f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A_c_165_n N_Y_c_1011_n 0.00468948f $X=2.84 $Y=1.202 $X2=0 $Y2=0
cc_206 N_A_c_159_n N_Y_c_1012_n 0.00262807f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A_c_160_n N_Y_c_1012_n 0.00113286f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A_c_175_p N_Y_c_1012_n 0.0266272f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A_c_165_n N_Y_c_1012_n 0.00230339f $X=2.84 $Y=1.202 $X2=0 $Y2=0
cc_210 N_A_c_160_n N_Y_c_1048_n 5.24636e-19 $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A_c_161_n N_Y_c_1048_n 0.00671723f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A_c_162_n N_Y_c_1048_n 0.00671723f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A_c_163_n N_Y_c_1048_n 5.24636e-19 $X=2.42 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A_c_162_n N_Y_c_1013_n 0.00929182f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A_c_163_n N_Y_c_1013_n 0.00929182f $X=2.42 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A_c_175_p N_Y_c_1013_n 0.0435408f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A_c_165_n N_Y_c_1013_n 0.00468948f $X=2.84 $Y=1.202 $X2=0 $Y2=0
cc_218 N_A_c_162_n N_Y_c_1056_n 5.24636e-19 $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A_c_163_n N_Y_c_1056_n 0.00671723f $X=2.42 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_c_164_n N_Y_c_1056_n 0.00671723f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A_c_164_n N_Y_c_1014_n 0.00972073f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A_c_175_p N_Y_c_1014_n 0.00550176f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A_c_165_n N_Y_c_1014_n 0.00164699f $X=2.84 $Y=1.202 $X2=0 $Y2=0
cc_224 N_A_c_164_n N_Y_c_1062_n 5.24636e-19 $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A_c_161_n N_Y_c_1023_n 0.00113286f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A_c_162_n N_Y_c_1023_n 0.00113286f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A_c_175_p N_Y_c_1023_n 0.0266272f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_228 N_A_c_165_n N_Y_c_1023_n 0.00230339f $X=2.84 $Y=1.202 $X2=0 $Y2=0
cc_229 N_A_c_163_n N_Y_c_1024_n 0.00113286f $X=2.42 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A_c_164_n N_Y_c_1024_n 0.00113286f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A_c_175_p N_Y_c_1024_n 0.0266272f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_232 N_A_c_165_n N_Y_c_1024_n 0.00230339f $X=2.84 $Y=1.202 $X2=0 $Y2=0
cc_233 N_A_c_159_n N_VGND_c_1319_n 0.0036824f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A_c_159_n N_VGND_c_1320_n 0.00541359f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A_c_160_n N_VGND_c_1320_n 0.00423334f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A_c_160_n N_VGND_c_1321_n 0.00166854f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A_c_161_n N_VGND_c_1321_n 0.00166854f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_238 N_A_c_161_n N_VGND_c_1322_n 0.00423334f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A_c_162_n N_VGND_c_1322_n 0.00423334f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A_c_162_n N_VGND_c_1323_n 0.00166854f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A_c_163_n N_VGND_c_1323_n 0.00166854f $X=2.42 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_c_163_n N_VGND_c_1324_n 0.00423334f $X=2.42 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A_c_164_n N_VGND_c_1324_n 0.00423334f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_c_164_n N_VGND_c_1325_n 0.00166854f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A_c_159_n N_VGND_c_1355_n 0.0105165f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_c_160_n N_VGND_c_1355_n 0.00595861f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A_c_161_n N_VGND_c_1355_n 0.00595861f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A_c_162_n N_VGND_c_1355_n 0.00595861f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A_c_163_n N_VGND_c_1355_n 0.00595861f $X=2.42 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A_c_164_n N_VGND_c_1355_n 0.00596967f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_251 N_B_c_272_n N_A_27_297#_c_609_n 2.98195e-19 $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_252 N_B_c_272_n N_A_27_297#_c_631_n 0.0143578f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_253 N_B_c_273_n N_A_27_297#_c_631_n 0.01161f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_254 N_B_c_274_n N_A_27_297#_c_633_n 0.01161f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_255 N_B_c_275_n N_A_27_297#_c_633_n 0.01161f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_256 N_B_c_276_n N_A_27_297#_c_610_n 0.01161f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_257 N_B_c_277_n N_A_27_297#_c_610_n 0.01161f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_258 N_B_c_272_n N_VPWR_c_698_n 0.00429453f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_259 N_B_c_273_n N_VPWR_c_698_n 0.00429453f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_260 N_B_c_274_n N_VPWR_c_698_n 0.00429453f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_261 N_B_c_275_n N_VPWR_c_698_n 0.00429453f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_262 N_B_c_276_n N_VPWR_c_698_n 0.00429453f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_263 N_B_c_277_n N_VPWR_c_698_n 0.00429453f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_264 N_B_c_272_n N_VPWR_c_692_n 0.00609021f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_265 N_B_c_273_n N_VPWR_c_692_n 0.00606499f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_266 N_B_c_274_n N_VPWR_c_692_n 0.00606499f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_267 N_B_c_275_n N_VPWR_c_692_n 0.00606499f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_268 N_B_c_276_n N_VPWR_c_692_n 0.00606499f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_269 N_B_c_277_n N_VPWR_c_692_n 0.00734734f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_270 N_B_c_273_n N_A_685_297#_c_830_n 0.0128188f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_271 N_B_c_274_n N_A_685_297#_c_830_n 0.0128795f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_272 N_B_c_281_n N_A_685_297#_c_830_n 0.0486996f $X=5.53 $Y=1.16 $X2=0 $Y2=0
cc_273 N_B_c_271_n N_A_685_297#_c_830_n 0.00844349f $X=5.66 $Y=1.202 $X2=0 $Y2=0
cc_274 N_B_c_275_n N_A_685_297#_c_831_n 0.0128795f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_275 N_B_c_276_n N_A_685_297#_c_831_n 0.0128795f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_276 N_B_c_281_n N_A_685_297#_c_831_n 0.0486996f $X=5.53 $Y=1.16 $X2=0 $Y2=0
cc_277 N_B_c_271_n N_A_685_297#_c_831_n 0.00844349f $X=5.66 $Y=1.202 $X2=0 $Y2=0
cc_278 N_B_c_277_n N_A_685_297#_c_832_n 0.0157575f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_279 N_B_c_281_n N_A_685_297#_c_832_n 0.00830509f $X=5.53 $Y=1.16 $X2=0 $Y2=0
cc_280 N_B_c_271_n N_A_685_297#_c_832_n 9.00973e-19 $X=5.66 $Y=1.202 $X2=0 $Y2=0
cc_281 N_B_c_272_n N_A_685_297#_c_835_n 2.98195e-19 $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_282 N_B_c_281_n N_A_685_297#_c_835_n 0.0204252f $X=5.53 $Y=1.16 $X2=0 $Y2=0
cc_283 N_B_c_271_n N_A_685_297#_c_835_n 0.00675794f $X=5.66 $Y=1.202 $X2=0 $Y2=0
cc_284 N_B_c_281_n N_A_685_297#_c_836_n 0.0204252f $X=5.53 $Y=1.16 $X2=0 $Y2=0
cc_285 N_B_c_271_n N_A_685_297#_c_836_n 0.00675794f $X=5.66 $Y=1.202 $X2=0 $Y2=0
cc_286 N_B_c_281_n N_A_685_297#_c_837_n 0.0204252f $X=5.53 $Y=1.16 $X2=0 $Y2=0
cc_287 N_B_c_271_n N_A_685_297#_c_837_n 0.00675794f $X=5.66 $Y=1.202 $X2=0 $Y2=0
cc_288 N_B_c_265_n N_Y_c_1056_n 5.24636e-19 $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_289 N_B_c_265_n N_Y_c_1014_n 0.0104562f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_290 N_B_c_281_n N_Y_c_1014_n 0.00550176f $X=5.53 $Y=1.16 $X2=0 $Y2=0
cc_291 N_B_c_271_n N_Y_c_1014_n 0.00224539f $X=5.66 $Y=1.202 $X2=0 $Y2=0
cc_292 N_B_c_265_n N_Y_c_1062_n 0.00671723f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_293 N_B_c_266_n N_Y_c_1062_n 0.00671723f $X=3.78 $Y=0.995 $X2=0 $Y2=0
cc_294 N_B_c_267_n N_Y_c_1062_n 5.24636e-19 $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_295 N_B_c_266_n N_Y_c_1015_n 0.00929182f $X=3.78 $Y=0.995 $X2=0 $Y2=0
cc_296 N_B_c_267_n N_Y_c_1015_n 0.00929182f $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_297 N_B_c_281_n N_Y_c_1015_n 0.0435408f $X=5.53 $Y=1.16 $X2=0 $Y2=0
cc_298 N_B_c_271_n N_Y_c_1015_n 0.00468948f $X=5.66 $Y=1.202 $X2=0 $Y2=0
cc_299 N_B_c_266_n N_Y_c_1082_n 5.24636e-19 $X=3.78 $Y=0.995 $X2=0 $Y2=0
cc_300 N_B_c_267_n N_Y_c_1082_n 0.00671723f $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_301 N_B_c_268_n N_Y_c_1082_n 0.00671723f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_302 N_B_c_269_n N_Y_c_1082_n 5.24636e-19 $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_303 N_B_c_268_n N_Y_c_1016_n 0.00929182f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_304 N_B_c_269_n N_Y_c_1016_n 0.00929182f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_305 N_B_c_281_n N_Y_c_1016_n 0.0435408f $X=5.53 $Y=1.16 $X2=0 $Y2=0
cc_306 N_B_c_271_n N_Y_c_1016_n 0.00468948f $X=5.66 $Y=1.202 $X2=0 $Y2=0
cc_307 N_B_c_268_n N_Y_c_1090_n 5.24636e-19 $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_308 N_B_c_269_n N_Y_c_1090_n 0.00671723f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_309 N_B_c_270_n N_Y_c_1090_n 0.0109565f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_310 N_B_c_270_n N_Y_c_1017_n 0.0114284f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_311 N_B_c_281_n N_Y_c_1017_n 0.00550176f $X=5.53 $Y=1.16 $X2=0 $Y2=0
cc_312 N_B_c_271_n N_Y_c_1017_n 0.00164699f $X=5.66 $Y=1.202 $X2=0 $Y2=0
cc_313 N_B_c_265_n N_Y_c_1025_n 0.00113286f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_314 N_B_c_266_n N_Y_c_1025_n 0.00113286f $X=3.78 $Y=0.995 $X2=0 $Y2=0
cc_315 N_B_c_281_n N_Y_c_1025_n 0.0266272f $X=5.53 $Y=1.16 $X2=0 $Y2=0
cc_316 N_B_c_271_n N_Y_c_1025_n 0.00230339f $X=5.66 $Y=1.202 $X2=0 $Y2=0
cc_317 N_B_c_267_n N_Y_c_1026_n 0.00113286f $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_318 N_B_c_268_n N_Y_c_1026_n 0.00113286f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_319 N_B_c_281_n N_Y_c_1026_n 0.0266272f $X=5.53 $Y=1.16 $X2=0 $Y2=0
cc_320 N_B_c_271_n N_Y_c_1026_n 0.00230339f $X=5.66 $Y=1.202 $X2=0 $Y2=0
cc_321 N_B_c_269_n N_Y_c_1027_n 0.00113286f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_322 N_B_c_270_n N_Y_c_1027_n 0.00113286f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_323 N_B_c_281_n N_Y_c_1027_n 0.0266272f $X=5.53 $Y=1.16 $X2=0 $Y2=0
cc_324 N_B_c_271_n N_Y_c_1027_n 0.00230339f $X=5.66 $Y=1.202 $X2=0 $Y2=0
cc_325 N_B_c_265_n N_VGND_c_1325_n 0.00166854f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_326 N_B_c_265_n N_VGND_c_1326_n 0.00423334f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_327 N_B_c_266_n N_VGND_c_1326_n 0.00423334f $X=3.78 $Y=0.995 $X2=0 $Y2=0
cc_328 N_B_c_266_n N_VGND_c_1327_n 0.00166854f $X=3.78 $Y=0.995 $X2=0 $Y2=0
cc_329 N_B_c_267_n N_VGND_c_1327_n 0.00166854f $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_330 N_B_c_268_n N_VGND_c_1328_n 0.00166854f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_331 N_B_c_269_n N_VGND_c_1328_n 0.00166738f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_332 N_B_c_267_n N_VGND_c_1336_n 0.00423334f $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_333 N_B_c_268_n N_VGND_c_1336_n 0.00423334f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_334 N_B_c_269_n N_VGND_c_1353_n 0.00423334f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_335 N_B_c_270_n N_VGND_c_1353_n 0.00423334f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_336 N_B_c_270_n N_VGND_c_1354_n 0.00336547f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_337 N_B_c_265_n N_VGND_c_1355_n 0.00596967f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_338 N_B_c_266_n N_VGND_c_1355_n 0.00595861f $X=3.78 $Y=0.995 $X2=0 $Y2=0
cc_339 N_B_c_267_n N_VGND_c_1355_n 0.00595861f $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_340 N_B_c_268_n N_VGND_c_1355_n 0.00595861f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_341 N_B_c_269_n N_VGND_c_1355_n 0.00595861f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_342 N_B_c_270_n N_VGND_c_1355_n 0.0070399f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_343 N_C_c_389_n N_D_c_497_n 0.0095757f $X=9.025 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_344 N_C_c_382_n N_D_c_489_n 0.0179509f $X=9 $Y=0.995 $X2=0 $Y2=0
cc_345 N_C_c_393_p N_D_c_495_n 0.00959259f $X=8.87 $Y=1.16 $X2=0 $Y2=0
cc_346 N_C_c_383_n N_D_c_495_n 9.65453e-19 $X=9 $Y=1.202 $X2=0 $Y2=0
cc_347 N_C_c_393_p N_D_c_496_n 2.28928e-19 $X=8.87 $Y=1.16 $X2=0 $Y2=0
cc_348 N_C_c_383_n N_D_c_496_n 0.0230009f $X=9 $Y=1.202 $X2=0 $Y2=0
cc_349 N_C_c_384_n N_VPWR_c_698_n 0.00429453f $X=6.675 $Y=1.41 $X2=0 $Y2=0
cc_350 N_C_c_385_n N_VPWR_c_698_n 0.00429453f $X=7.145 $Y=1.41 $X2=0 $Y2=0
cc_351 N_C_c_386_n N_VPWR_c_698_n 0.00429453f $X=7.615 $Y=1.41 $X2=0 $Y2=0
cc_352 N_C_c_387_n N_VPWR_c_698_n 0.00429453f $X=8.085 $Y=1.41 $X2=0 $Y2=0
cc_353 N_C_c_388_n N_VPWR_c_698_n 0.00429453f $X=8.555 $Y=1.41 $X2=0 $Y2=0
cc_354 N_C_c_389_n N_VPWR_c_698_n 0.00429453f $X=9.025 $Y=1.41 $X2=0 $Y2=0
cc_355 N_C_c_384_n N_VPWR_c_692_n 0.00734734f $X=6.675 $Y=1.41 $X2=0 $Y2=0
cc_356 N_C_c_385_n N_VPWR_c_692_n 0.00606499f $X=7.145 $Y=1.41 $X2=0 $Y2=0
cc_357 N_C_c_386_n N_VPWR_c_692_n 0.00606499f $X=7.615 $Y=1.41 $X2=0 $Y2=0
cc_358 N_C_c_387_n N_VPWR_c_692_n 0.00606499f $X=8.085 $Y=1.41 $X2=0 $Y2=0
cc_359 N_C_c_388_n N_VPWR_c_692_n 0.00606499f $X=8.555 $Y=1.41 $X2=0 $Y2=0
cc_360 N_C_c_389_n N_VPWR_c_692_n 0.00609021f $X=9.025 $Y=1.41 $X2=0 $Y2=0
cc_361 N_C_c_384_n N_A_685_297#_c_832_n 0.0157575f $X=6.675 $Y=1.41 $X2=0 $Y2=0
cc_362 N_C_c_393_p N_A_685_297#_c_832_n 0.00830509f $X=8.87 $Y=1.16 $X2=0 $Y2=0
cc_363 N_C_c_383_n N_A_685_297#_c_832_n 9.00973e-19 $X=9 $Y=1.202 $X2=0 $Y2=0
cc_364 N_C_c_385_n N_A_685_297#_c_833_n 0.0128795f $X=7.145 $Y=1.41 $X2=0 $Y2=0
cc_365 N_C_c_386_n N_A_685_297#_c_833_n 0.0128795f $X=7.615 $Y=1.41 $X2=0 $Y2=0
cc_366 N_C_c_393_p N_A_685_297#_c_833_n 0.0486996f $X=8.87 $Y=1.16 $X2=0 $Y2=0
cc_367 N_C_c_383_n N_A_685_297#_c_833_n 0.00844349f $X=9 $Y=1.202 $X2=0 $Y2=0
cc_368 N_C_c_387_n N_A_685_297#_c_834_n 0.0128795f $X=8.085 $Y=1.41 $X2=0 $Y2=0
cc_369 N_C_c_388_n N_A_685_297#_c_834_n 0.0128188f $X=8.555 $Y=1.41 $X2=0 $Y2=0
cc_370 N_C_c_393_p N_A_685_297#_c_834_n 0.0486996f $X=8.87 $Y=1.16 $X2=0 $Y2=0
cc_371 N_C_c_383_n N_A_685_297#_c_834_n 0.00844349f $X=9 $Y=1.202 $X2=0 $Y2=0
cc_372 N_C_c_393_p N_A_685_297#_c_838_n 0.0204252f $X=8.87 $Y=1.16 $X2=0 $Y2=0
cc_373 N_C_c_383_n N_A_685_297#_c_838_n 0.00675794f $X=9 $Y=1.202 $X2=0 $Y2=0
cc_374 N_C_c_393_p N_A_685_297#_c_839_n 0.0204252f $X=8.87 $Y=1.16 $X2=0 $Y2=0
cc_375 N_C_c_383_n N_A_685_297#_c_839_n 0.00675794f $X=9 $Y=1.202 $X2=0 $Y2=0
cc_376 N_C_c_389_n N_A_685_297#_c_840_n 2.98817e-19 $X=9.025 $Y=1.41 $X2=0 $Y2=0
cc_377 N_C_c_393_p N_A_685_297#_c_840_n 0.0204252f $X=8.87 $Y=1.16 $X2=0 $Y2=0
cc_378 N_C_c_383_n N_A_685_297#_c_840_n 0.00675794f $X=9 $Y=1.202 $X2=0 $Y2=0
cc_379 N_C_c_384_n N_A_1263_297#_c_925_n 0.01161f $X=6.675 $Y=1.41 $X2=0 $Y2=0
cc_380 N_C_c_385_n N_A_1263_297#_c_925_n 0.01161f $X=7.145 $Y=1.41 $X2=0 $Y2=0
cc_381 N_C_c_386_n N_A_1263_297#_c_927_n 0.01161f $X=7.615 $Y=1.41 $X2=0 $Y2=0
cc_382 N_C_c_387_n N_A_1263_297#_c_927_n 0.01161f $X=8.085 $Y=1.41 $X2=0 $Y2=0
cc_383 N_C_c_388_n N_A_1263_297#_c_929_n 0.01161f $X=8.555 $Y=1.41 $X2=0 $Y2=0
cc_384 N_C_c_389_n N_A_1263_297#_c_929_n 0.0143578f $X=9.025 $Y=1.41 $X2=0 $Y2=0
cc_385 N_C_c_389_n N_A_1263_297#_c_922_n 2.65342e-19 $X=9.025 $Y=1.41 $X2=0
+ $Y2=0
cc_386 N_C_c_377_n N_Y_c_1017_n 0.0114284f $X=6.7 $Y=0.995 $X2=0 $Y2=0
cc_387 N_C_c_393_p N_Y_c_1017_n 0.00550176f $X=8.87 $Y=1.16 $X2=0 $Y2=0
cc_388 N_C_c_383_n N_Y_c_1017_n 0.00164699f $X=9 $Y=1.202 $X2=0 $Y2=0
cc_389 N_C_c_377_n N_Y_c_1111_n 0.0109565f $X=6.7 $Y=0.995 $X2=0 $Y2=0
cc_390 N_C_c_378_n N_Y_c_1111_n 0.00671723f $X=7.12 $Y=0.995 $X2=0 $Y2=0
cc_391 N_C_c_379_n N_Y_c_1111_n 5.24636e-19 $X=7.64 $Y=0.995 $X2=0 $Y2=0
cc_392 N_C_c_378_n N_Y_c_1018_n 0.00929182f $X=7.12 $Y=0.995 $X2=0 $Y2=0
cc_393 N_C_c_379_n N_Y_c_1018_n 0.00929182f $X=7.64 $Y=0.995 $X2=0 $Y2=0
cc_394 N_C_c_393_p N_Y_c_1018_n 0.0435408f $X=8.87 $Y=1.16 $X2=0 $Y2=0
cc_395 N_C_c_383_n N_Y_c_1018_n 0.00468948f $X=9 $Y=1.202 $X2=0 $Y2=0
cc_396 N_C_c_378_n N_Y_c_1118_n 5.24636e-19 $X=7.12 $Y=0.995 $X2=0 $Y2=0
cc_397 N_C_c_379_n N_Y_c_1118_n 0.00671723f $X=7.64 $Y=0.995 $X2=0 $Y2=0
cc_398 N_C_c_380_n N_Y_c_1118_n 0.00671723f $X=8.06 $Y=0.995 $X2=0 $Y2=0
cc_399 N_C_c_381_n N_Y_c_1118_n 5.24636e-19 $X=8.58 $Y=0.995 $X2=0 $Y2=0
cc_400 N_C_c_380_n N_Y_c_1019_n 0.00929182f $X=8.06 $Y=0.995 $X2=0 $Y2=0
cc_401 N_C_c_381_n N_Y_c_1019_n 0.00929182f $X=8.58 $Y=0.995 $X2=0 $Y2=0
cc_402 N_C_c_393_p N_Y_c_1019_n 0.0435408f $X=8.87 $Y=1.16 $X2=0 $Y2=0
cc_403 N_C_c_383_n N_Y_c_1019_n 0.00468948f $X=9 $Y=1.202 $X2=0 $Y2=0
cc_404 N_C_c_380_n N_Y_c_1126_n 5.24636e-19 $X=8.06 $Y=0.995 $X2=0 $Y2=0
cc_405 N_C_c_381_n N_Y_c_1126_n 0.00671723f $X=8.58 $Y=0.995 $X2=0 $Y2=0
cc_406 N_C_c_382_n N_Y_c_1126_n 0.00671723f $X=9 $Y=0.995 $X2=0 $Y2=0
cc_407 N_C_c_382_n N_Y_c_1020_n 0.0104562f $X=9 $Y=0.995 $X2=0 $Y2=0
cc_408 N_C_c_393_p N_Y_c_1020_n 0.00550176f $X=8.87 $Y=1.16 $X2=0 $Y2=0
cc_409 N_C_c_383_n N_Y_c_1020_n 0.00224539f $X=9 $Y=1.202 $X2=0 $Y2=0
cc_410 N_C_c_382_n N_Y_c_1132_n 5.24636e-19 $X=9 $Y=0.995 $X2=0 $Y2=0
cc_411 N_C_c_377_n N_Y_c_1028_n 0.00113286f $X=6.7 $Y=0.995 $X2=0 $Y2=0
cc_412 N_C_c_378_n N_Y_c_1028_n 0.00113286f $X=7.12 $Y=0.995 $X2=0 $Y2=0
cc_413 N_C_c_393_p N_Y_c_1028_n 0.0266272f $X=8.87 $Y=1.16 $X2=0 $Y2=0
cc_414 N_C_c_383_n N_Y_c_1028_n 0.00230339f $X=9 $Y=1.202 $X2=0 $Y2=0
cc_415 N_C_c_379_n N_Y_c_1029_n 0.00113286f $X=7.64 $Y=0.995 $X2=0 $Y2=0
cc_416 N_C_c_380_n N_Y_c_1029_n 0.00113286f $X=8.06 $Y=0.995 $X2=0 $Y2=0
cc_417 N_C_c_393_p N_Y_c_1029_n 0.0266272f $X=8.87 $Y=1.16 $X2=0 $Y2=0
cc_418 N_C_c_383_n N_Y_c_1029_n 0.00230339f $X=9 $Y=1.202 $X2=0 $Y2=0
cc_419 N_C_c_381_n N_Y_c_1030_n 0.00113286f $X=8.58 $Y=0.995 $X2=0 $Y2=0
cc_420 N_C_c_382_n N_Y_c_1030_n 0.00113286f $X=9 $Y=0.995 $X2=0 $Y2=0
cc_421 N_C_c_393_p N_Y_c_1030_n 0.0266272f $X=8.87 $Y=1.16 $X2=0 $Y2=0
cc_422 N_C_c_383_n N_Y_c_1030_n 0.00230339f $X=9 $Y=1.202 $X2=0 $Y2=0
cc_423 N_C_c_378_n N_VGND_c_1329_n 0.00166738f $X=7.12 $Y=0.995 $X2=0 $Y2=0
cc_424 N_C_c_379_n N_VGND_c_1329_n 0.00166854f $X=7.64 $Y=0.995 $X2=0 $Y2=0
cc_425 N_C_c_380_n N_VGND_c_1330_n 0.00166854f $X=8.06 $Y=0.995 $X2=0 $Y2=0
cc_426 N_C_c_381_n N_VGND_c_1330_n 0.00166854f $X=8.58 $Y=0.995 $X2=0 $Y2=0
cc_427 N_C_c_382_n N_VGND_c_1331_n 0.00166854f $X=9 $Y=0.995 $X2=0 $Y2=0
cc_428 N_C_c_377_n N_VGND_c_1338_n 0.00423334f $X=6.7 $Y=0.995 $X2=0 $Y2=0
cc_429 N_C_c_378_n N_VGND_c_1338_n 0.00423334f $X=7.12 $Y=0.995 $X2=0 $Y2=0
cc_430 N_C_c_379_n N_VGND_c_1340_n 0.00423334f $X=7.64 $Y=0.995 $X2=0 $Y2=0
cc_431 N_C_c_380_n N_VGND_c_1340_n 0.00423334f $X=8.06 $Y=0.995 $X2=0 $Y2=0
cc_432 N_C_c_381_n N_VGND_c_1342_n 0.00423334f $X=8.58 $Y=0.995 $X2=0 $Y2=0
cc_433 N_C_c_382_n N_VGND_c_1342_n 0.00423334f $X=9 $Y=0.995 $X2=0 $Y2=0
cc_434 N_C_c_377_n N_VGND_c_1354_n 0.00336547f $X=6.7 $Y=0.995 $X2=0 $Y2=0
cc_435 N_C_c_377_n N_VGND_c_1355_n 0.0070399f $X=6.7 $Y=0.995 $X2=0 $Y2=0
cc_436 N_C_c_378_n N_VGND_c_1355_n 0.00595861f $X=7.12 $Y=0.995 $X2=0 $Y2=0
cc_437 N_C_c_379_n N_VGND_c_1355_n 0.00595861f $X=7.64 $Y=0.995 $X2=0 $Y2=0
cc_438 N_C_c_380_n N_VGND_c_1355_n 0.00595861f $X=8.06 $Y=0.995 $X2=0 $Y2=0
cc_439 N_C_c_381_n N_VGND_c_1355_n 0.00595861f $X=8.58 $Y=0.995 $X2=0 $Y2=0
cc_440 N_C_c_382_n N_VGND_c_1355_n 0.00596967f $X=9 $Y=0.995 $X2=0 $Y2=0
cc_441 N_D_c_497_n N_VPWR_c_698_n 0.00429453f $X=9.495 $Y=1.41 $X2=0 $Y2=0
cc_442 N_D_c_498_n N_VPWR_c_698_n 0.00429453f $X=9.965 $Y=1.41 $X2=0 $Y2=0
cc_443 N_D_c_499_n N_VPWR_c_698_n 0.00429453f $X=10.435 $Y=1.41 $X2=0 $Y2=0
cc_444 N_D_c_500_n N_VPWR_c_698_n 0.00429453f $X=10.905 $Y=1.41 $X2=0 $Y2=0
cc_445 N_D_c_501_n N_VPWR_c_698_n 0.00429453f $X=11.375 $Y=1.41 $X2=0 $Y2=0
cc_446 N_D_c_502_n N_VPWR_c_698_n 0.00429453f $X=11.845 $Y=1.41 $X2=0 $Y2=0
cc_447 N_D_c_497_n N_VPWR_c_692_n 0.00609021f $X=9.495 $Y=1.41 $X2=0 $Y2=0
cc_448 N_D_c_498_n N_VPWR_c_692_n 0.00606499f $X=9.965 $Y=1.41 $X2=0 $Y2=0
cc_449 N_D_c_499_n N_VPWR_c_692_n 0.00606499f $X=10.435 $Y=1.41 $X2=0 $Y2=0
cc_450 N_D_c_500_n N_VPWR_c_692_n 0.00606499f $X=10.905 $Y=1.41 $X2=0 $Y2=0
cc_451 N_D_c_501_n N_VPWR_c_692_n 0.00606499f $X=11.375 $Y=1.41 $X2=0 $Y2=0
cc_452 N_D_c_502_n N_VPWR_c_692_n 0.00704277f $X=11.845 $Y=1.41 $X2=0 $Y2=0
cc_453 N_D_c_497_n N_A_1263_297#_c_922_n 2.65342e-19 $X=9.495 $Y=1.41 $X2=0
+ $Y2=0
cc_454 N_D_c_497_n N_A_1263_297#_c_933_n 0.0143578f $X=9.495 $Y=1.41 $X2=0 $Y2=0
cc_455 N_D_c_498_n N_A_1263_297#_c_933_n 0.01161f $X=9.965 $Y=1.41 $X2=0 $Y2=0
cc_456 N_D_c_499_n N_A_1263_297#_c_935_n 0.01161f $X=10.435 $Y=1.41 $X2=0 $Y2=0
cc_457 N_D_c_500_n N_A_1263_297#_c_935_n 0.01161f $X=10.905 $Y=1.41 $X2=0 $Y2=0
cc_458 N_D_c_501_n N_A_1263_297#_c_937_n 0.0112917f $X=11.375 $Y=1.41 $X2=0
+ $Y2=0
cc_459 N_D_c_502_n N_A_1263_297#_c_937_n 0.0119418f $X=11.845 $Y=1.41 $X2=0
+ $Y2=0
cc_460 N_D_c_502_n N_A_1263_297#_c_924_n 0.00612903f $X=11.845 $Y=1.41 $X2=0
+ $Y2=0
cc_461 N_D_c_489_n N_Y_c_1126_n 5.24636e-19 $X=9.52 $Y=0.995 $X2=0 $Y2=0
cc_462 N_D_c_489_n N_Y_c_1020_n 0.00922411f $X=9.52 $Y=0.995 $X2=0 $Y2=0
cc_463 N_D_c_495_n N_Y_c_1020_n 0.011918f $X=10.92 $Y=1.16 $X2=0 $Y2=0
cc_464 N_D_c_496_n N_Y_c_1020_n 0.00141784f $X=11.82 $Y=1.202 $X2=0 $Y2=0
cc_465 N_D_c_489_n N_Y_c_1132_n 0.00671723f $X=9.52 $Y=0.995 $X2=0 $Y2=0
cc_466 N_D_c_490_n N_Y_c_1132_n 0.00671723f $X=9.94 $Y=0.995 $X2=0 $Y2=0
cc_467 N_D_c_491_n N_Y_c_1132_n 5.24636e-19 $X=10.46 $Y=0.995 $X2=0 $Y2=0
cc_468 N_D_c_498_n N_Y_c_1033_n 0.0128188f $X=9.965 $Y=1.41 $X2=0 $Y2=0
cc_469 N_D_c_499_n N_Y_c_1033_n 0.0128795f $X=10.435 $Y=1.41 $X2=0 $Y2=0
cc_470 N_D_c_495_n N_Y_c_1033_n 0.0486996f $X=10.92 $Y=1.16 $X2=0 $Y2=0
cc_471 N_D_c_496_n N_Y_c_1033_n 0.00844349f $X=11.82 $Y=1.202 $X2=0 $Y2=0
cc_472 N_D_c_490_n N_Y_c_1021_n 0.00929182f $X=9.94 $Y=0.995 $X2=0 $Y2=0
cc_473 N_D_c_491_n N_Y_c_1021_n 0.00929182f $X=10.46 $Y=0.995 $X2=0 $Y2=0
cc_474 N_D_c_495_n N_Y_c_1021_n 0.0435408f $X=10.92 $Y=1.16 $X2=0 $Y2=0
cc_475 N_D_c_496_n N_Y_c_1021_n 0.00468948f $X=11.82 $Y=1.202 $X2=0 $Y2=0
cc_476 N_D_c_490_n N_Y_c_1160_n 5.24636e-19 $X=9.94 $Y=0.995 $X2=0 $Y2=0
cc_477 N_D_c_491_n N_Y_c_1160_n 0.00671723f $X=10.46 $Y=0.995 $X2=0 $Y2=0
cc_478 N_D_c_492_n N_Y_c_1160_n 0.00671723f $X=10.88 $Y=0.995 $X2=0 $Y2=0
cc_479 N_D_c_493_n N_Y_c_1160_n 5.24636e-19 $X=11.4 $Y=0.995 $X2=0 $Y2=0
cc_480 N_D_c_500_n N_Y_c_1034_n 0.0128795f $X=10.905 $Y=1.41 $X2=0 $Y2=0
cc_481 N_D_c_501_n N_Y_c_1034_n 0.0132089f $X=11.375 $Y=1.41 $X2=0 $Y2=0
cc_482 N_D_c_495_n N_Y_c_1034_n 0.0203546f $X=10.92 $Y=1.16 $X2=0 $Y2=0
cc_483 N_D_c_496_n N_Y_c_1034_n 0.00871238f $X=11.82 $Y=1.202 $X2=0 $Y2=0
cc_484 N_D_c_492_n N_Y_c_1022_n 0.00929182f $X=10.88 $Y=0.995 $X2=0 $Y2=0
cc_485 N_D_c_493_n N_Y_c_1022_n 0.0106784f $X=11.4 $Y=0.995 $X2=0 $Y2=0
cc_486 N_D_c_495_n N_Y_c_1022_n 0.0177573f $X=10.92 $Y=1.16 $X2=0 $Y2=0
cc_487 N_D_c_496_n N_Y_c_1022_n 0.00537693f $X=11.82 $Y=1.202 $X2=0 $Y2=0
cc_488 N_D_c_492_n N_Y_c_1172_n 5.23845e-19 $X=10.88 $Y=0.995 $X2=0 $Y2=0
cc_489 N_D_c_493_n N_Y_c_1172_n 0.00671723f $X=11.4 $Y=0.995 $X2=0 $Y2=0
cc_490 N_D_c_494_n N_Y_c_1172_n 0.00777777f $X=11.82 $Y=0.995 $X2=0 $Y2=0
cc_491 N_D_c_489_n N_Y_c_1031_n 0.00113286f $X=9.52 $Y=0.995 $X2=0 $Y2=0
cc_492 N_D_c_490_n N_Y_c_1031_n 0.00113286f $X=9.94 $Y=0.995 $X2=0 $Y2=0
cc_493 N_D_c_495_n N_Y_c_1031_n 0.0266272f $X=10.92 $Y=1.16 $X2=0 $Y2=0
cc_494 N_D_c_496_n N_Y_c_1031_n 0.00230339f $X=11.82 $Y=1.202 $X2=0 $Y2=0
cc_495 N_D_c_497_n N_Y_c_1035_n 2.98817e-19 $X=9.495 $Y=1.41 $X2=0 $Y2=0
cc_496 N_D_c_495_n N_Y_c_1035_n 0.0204252f $X=10.92 $Y=1.16 $X2=0 $Y2=0
cc_497 N_D_c_496_n N_Y_c_1035_n 0.00675794f $X=11.82 $Y=1.202 $X2=0 $Y2=0
cc_498 N_D_c_491_n N_Y_c_1032_n 0.00113286f $X=10.46 $Y=0.995 $X2=0 $Y2=0
cc_499 N_D_c_492_n N_Y_c_1032_n 0.00113286f $X=10.88 $Y=0.995 $X2=0 $Y2=0
cc_500 N_D_c_495_n N_Y_c_1032_n 0.0266272f $X=10.92 $Y=1.16 $X2=0 $Y2=0
cc_501 N_D_c_496_n N_Y_c_1032_n 0.00230339f $X=11.82 $Y=1.202 $X2=0 $Y2=0
cc_502 N_D_c_495_n N_Y_c_1036_n 0.0204252f $X=10.92 $Y=1.16 $X2=0 $Y2=0
cc_503 N_D_c_496_n N_Y_c_1036_n 0.00675794f $X=11.82 $Y=1.202 $X2=0 $Y2=0
cc_504 N_D_c_493_n N_Y_c_1188_n 7.13294e-19 $X=11.4 $Y=0.995 $X2=0 $Y2=0
cc_505 N_D_c_494_n N_Y_c_1188_n 0.00292444f $X=11.82 $Y=0.995 $X2=0 $Y2=0
cc_506 N_D_c_500_n N_Y_c_1190_n 5.27206e-19 $X=10.905 $Y=1.41 $X2=0 $Y2=0
cc_507 N_D_c_501_n N_Y_c_1190_n 0.00780896f $X=11.375 $Y=1.41 $X2=0 $Y2=0
cc_508 N_D_c_502_n N_Y_c_1190_n 0.0116317f $X=11.845 $Y=1.41 $X2=0 $Y2=0
cc_509 N_D_c_492_n Y 4.16977e-19 $X=10.88 $Y=0.995 $X2=0 $Y2=0
cc_510 N_D_c_500_n Y 2.01376e-19 $X=10.905 $Y=1.41 $X2=0 $Y2=0
cc_511 N_D_c_501_n Y 0.00134899f $X=11.375 $Y=1.41 $X2=0 $Y2=0
cc_512 N_D_c_493_n Y 0.00281406f $X=11.4 $Y=0.995 $X2=0 $Y2=0
cc_513 N_D_c_494_n Y 0.0053721f $X=11.82 $Y=0.995 $X2=0 $Y2=0
cc_514 N_D_c_502_n Y 0.00264009f $X=11.845 $Y=1.41 $X2=0 $Y2=0
cc_515 N_D_c_495_n Y 0.00917996f $X=10.92 $Y=1.16 $X2=0 $Y2=0
cc_516 N_D_c_496_n Y 0.0539813f $X=11.82 $Y=1.202 $X2=0 $Y2=0
cc_517 N_D_c_489_n N_VGND_c_1331_n 0.00166854f $X=9.52 $Y=0.995 $X2=0 $Y2=0
cc_518 N_D_c_490_n N_VGND_c_1332_n 0.00166854f $X=9.94 $Y=0.995 $X2=0 $Y2=0
cc_519 N_D_c_491_n N_VGND_c_1332_n 0.00166854f $X=10.46 $Y=0.995 $X2=0 $Y2=0
cc_520 N_D_c_492_n N_VGND_c_1333_n 0.00166854f $X=10.88 $Y=0.995 $X2=0 $Y2=0
cc_521 N_D_c_493_n N_VGND_c_1333_n 0.00296353f $X=11.4 $Y=0.995 $X2=0 $Y2=0
cc_522 N_D_c_494_n N_VGND_c_1335_n 0.00651338f $X=11.82 $Y=0.995 $X2=0 $Y2=0
cc_523 N_D_c_489_n N_VGND_c_1344_n 0.00423334f $X=9.52 $Y=0.995 $X2=0 $Y2=0
cc_524 N_D_c_490_n N_VGND_c_1344_n 0.00423334f $X=9.94 $Y=0.995 $X2=0 $Y2=0
cc_525 N_D_c_491_n N_VGND_c_1346_n 0.00423334f $X=10.46 $Y=0.995 $X2=0 $Y2=0
cc_526 N_D_c_492_n N_VGND_c_1346_n 0.00423334f $X=10.88 $Y=0.995 $X2=0 $Y2=0
cc_527 N_D_c_493_n N_VGND_c_1348_n 0.00423334f $X=11.4 $Y=0.995 $X2=0 $Y2=0
cc_528 N_D_c_494_n N_VGND_c_1348_n 0.00450273f $X=11.82 $Y=0.995 $X2=0 $Y2=0
cc_529 N_D_c_489_n N_VGND_c_1355_n 0.00596967f $X=9.52 $Y=0.995 $X2=0 $Y2=0
cc_530 N_D_c_490_n N_VGND_c_1355_n 0.00595861f $X=9.94 $Y=0.995 $X2=0 $Y2=0
cc_531 N_D_c_491_n N_VGND_c_1355_n 0.00595861f $X=10.46 $Y=0.995 $X2=0 $Y2=0
cc_532 N_D_c_492_n N_VGND_c_1355_n 0.00595861f $X=10.88 $Y=0.995 $X2=0 $Y2=0
cc_533 N_D_c_493_n N_VGND_c_1355_n 0.00595861f $X=11.4 $Y=0.995 $X2=0 $Y2=0
cc_534 N_D_c_494_n N_VGND_c_1355_n 0.00846284f $X=11.82 $Y=0.995 $X2=0 $Y2=0
cc_535 N_A_27_297#_c_606_n N_VPWR_M1000_d 0.00187091f $X=1.095 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_536 N_A_27_297#_c_607_n N_VPWR_M1014_d 0.00187091f $X=2.035 $Y=1.54 $X2=0
+ $Y2=0
cc_537 N_A_27_297#_c_608_n N_VPWR_M1030_d 0.00187091f $X=2.975 $Y=1.54 $X2=0
+ $Y2=0
cc_538 N_A_27_297#_c_606_n N_VPWR_c_693_n 0.0143191f $X=1.095 $Y=1.54 $X2=0
+ $Y2=0
cc_539 N_A_27_297#_c_641_p N_VPWR_c_694_n 0.0149311f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_540 N_A_27_297#_c_607_n N_VPWR_c_695_n 0.0143191f $X=2.035 $Y=1.54 $X2=0
+ $Y2=0
cc_541 N_A_27_297#_c_643_p N_VPWR_c_696_n 0.0149311f $X=2.16 $Y=2.3 $X2=0 $Y2=0
cc_542 N_A_27_297#_c_608_n N_VPWR_c_697_n 0.0143191f $X=2.975 $Y=1.54 $X2=0
+ $Y2=0
cc_543 N_A_27_297#_c_645_p N_VPWR_c_698_n 0.015002f $X=3.1 $Y=2.295 $X2=0 $Y2=0
cc_544 N_A_27_297#_c_631_n N_VPWR_c_698_n 0.0386815f $X=3.915 $Y=2.38 $X2=0
+ $Y2=0
cc_545 N_A_27_297#_c_633_n N_VPWR_c_698_n 0.0386815f $X=4.855 $Y=2.38 $X2=0
+ $Y2=0
cc_546 N_A_27_297#_c_610_n N_VPWR_c_698_n 0.057821f $X=5.795 $Y=2.38 $X2=0 $Y2=0
cc_547 N_A_27_297#_c_649_p N_VPWR_c_698_n 0.0149886f $X=4.04 $Y=2.38 $X2=0 $Y2=0
cc_548 N_A_27_297#_c_650_p N_VPWR_c_698_n 0.0149886f $X=4.98 $Y=2.38 $X2=0 $Y2=0
cc_549 N_A_27_297#_M1000_s N_VPWR_c_692_n 0.00303344f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_550 N_A_27_297#_M1005_s N_VPWR_c_692_n 0.00370124f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_551 N_A_27_297#_M1020_s N_VPWR_c_692_n 0.00370124f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_552 N_A_27_297#_M1042_s N_VPWR_c_692_n 0.00297222f $X=2.955 $Y=1.485 $X2=0
+ $Y2=0
cc_553 N_A_27_297#_M1017_d N_VPWR_c_692_n 0.00231264f $X=3.895 $Y=1.485 $X2=0
+ $Y2=0
cc_554 N_A_27_297#_M1033_d N_VPWR_c_692_n 0.00231264f $X=4.835 $Y=1.485 $X2=0
+ $Y2=0
cc_555 N_A_27_297#_M1040_d N_VPWR_c_692_n 0.00217519f $X=5.775 $Y=1.485 $X2=0
+ $Y2=0
cc_556 N_A_27_297#_c_605_n N_VPWR_c_692_n 0.0110914f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_557 N_A_27_297#_c_641_p N_VPWR_c_692_n 0.00955092f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_558 N_A_27_297#_c_643_p N_VPWR_c_692_n 0.00955092f $X=2.16 $Y=2.3 $X2=0 $Y2=0
cc_559 N_A_27_297#_c_645_p N_VPWR_c_692_n 0.00962794f $X=3.1 $Y=2.295 $X2=0
+ $Y2=0
cc_560 N_A_27_297#_c_631_n N_VPWR_c_692_n 0.0239144f $X=3.915 $Y=2.38 $X2=0
+ $Y2=0
cc_561 N_A_27_297#_c_633_n N_VPWR_c_692_n 0.0239144f $X=4.855 $Y=2.38 $X2=0
+ $Y2=0
cc_562 N_A_27_297#_c_610_n N_VPWR_c_692_n 0.0350785f $X=5.795 $Y=2.38 $X2=0
+ $Y2=0
cc_563 N_A_27_297#_c_649_p N_VPWR_c_692_n 0.00962421f $X=4.04 $Y=2.38 $X2=0
+ $Y2=0
cc_564 N_A_27_297#_c_650_p N_VPWR_c_692_n 0.00962421f $X=4.98 $Y=2.38 $X2=0
+ $Y2=0
cc_565 N_A_27_297#_c_605_n N_VPWR_c_700_n 0.0190242f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_566 N_A_27_297#_c_631_n N_A_685_297#_M1009_s 0.00352392f $X=3.915 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_567 N_A_27_297#_c_633_n N_A_685_297#_M1024_s 0.00352392f $X=4.855 $Y=2.38
+ $X2=0 $Y2=0
cc_568 N_A_27_297#_c_610_n N_A_685_297#_M1035_s 0.00352392f $X=5.795 $Y=2.38
+ $X2=0 $Y2=0
cc_569 N_A_27_297#_M1017_d N_A_685_297#_c_830_n 0.00187091f $X=3.895 $Y=1.485
+ $X2=0 $Y2=0
cc_570 N_A_27_297#_c_631_n N_A_685_297#_c_830_n 0.00385532f $X=3.915 $Y=2.38
+ $X2=0 $Y2=0
cc_571 N_A_27_297#_c_673_p N_A_685_297#_c_830_n 0.0143018f $X=4.04 $Y=1.96 $X2=0
+ $Y2=0
cc_572 N_A_27_297#_c_633_n N_A_685_297#_c_830_n 0.00385532f $X=4.855 $Y=2.38
+ $X2=0 $Y2=0
cc_573 N_A_27_297#_M1033_d N_A_685_297#_c_831_n 0.00187091f $X=4.835 $Y=1.485
+ $X2=0 $Y2=0
cc_574 N_A_27_297#_c_633_n N_A_685_297#_c_831_n 0.00385532f $X=4.855 $Y=2.38
+ $X2=0 $Y2=0
cc_575 N_A_27_297#_c_677_p N_A_685_297#_c_831_n 0.0143018f $X=4.98 $Y=1.96 $X2=0
+ $Y2=0
cc_576 N_A_27_297#_c_610_n N_A_685_297#_c_831_n 0.00385532f $X=5.795 $Y=2.38
+ $X2=0 $Y2=0
cc_577 N_A_27_297#_M1040_d N_A_685_297#_c_832_n 0.00295666f $X=5.775 $Y=1.485
+ $X2=0 $Y2=0
cc_578 N_A_27_297#_c_610_n N_A_685_297#_c_832_n 0.00385532f $X=5.795 $Y=2.38
+ $X2=0 $Y2=0
cc_579 N_A_27_297#_c_611_n N_A_685_297#_c_832_n 0.0205983f $X=5.92 $Y=1.96 $X2=0
+ $Y2=0
cc_580 N_A_27_297#_c_609_n N_A_685_297#_c_835_n 0.00226124f $X=3.1 $Y=1.625
+ $X2=0 $Y2=0
cc_581 N_A_27_297#_c_631_n N_A_685_297#_c_835_n 0.013395f $X=3.915 $Y=2.38 $X2=0
+ $Y2=0
cc_582 N_A_27_297#_c_633_n N_A_685_297#_c_836_n 0.013395f $X=4.855 $Y=2.38 $X2=0
+ $Y2=0
cc_583 N_A_27_297#_c_610_n N_A_685_297#_c_837_n 0.013395f $X=5.795 $Y=2.38 $X2=0
+ $Y2=0
cc_584 N_A_27_297#_c_611_n N_A_1263_297#_c_920_n 0.0376802f $X=5.92 $Y=1.96
+ $X2=0 $Y2=0
cc_585 N_A_27_297#_c_610_n N_A_1263_297#_c_921_n 0.0147157f $X=5.795 $Y=2.38
+ $X2=0 $Y2=0
cc_586 N_A_27_297#_c_608_n N_Y_c_1014_n 0.00286947f $X=2.975 $Y=1.54 $X2=0 $Y2=0
cc_587 N_A_27_297#_c_609_n N_Y_c_1014_n 0.00936521f $X=3.1 $Y=1.625 $X2=0 $Y2=0
cc_588 N_A_27_297#_c_604_n N_VGND_c_1319_n 0.0119289f $X=0.26 $Y=1.625 $X2=0
+ $Y2=0
cc_589 N_A_27_297#_c_606_n N_VGND_c_1319_n 3.19131e-19 $X=1.095 $Y=1.54 $X2=0
+ $Y2=0
cc_590 N_VPWR_c_692_n N_A_685_297#_M1009_s 0.00232895f $X=12.19 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_591 N_VPWR_c_692_n N_A_685_297#_M1024_s 0.00232895f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_592 N_VPWR_c_692_n N_A_685_297#_M1035_s 0.00232895f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_593 N_VPWR_c_692_n N_A_685_297#_M1001_s 0.00232895f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_594 N_VPWR_c_692_n N_A_685_297#_M1015_s 0.00232895f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_595 N_VPWR_c_692_n N_A_685_297#_M1043_s 0.00232895f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_596 N_VPWR_c_692_n N_A_1263_297#_M1001_d 0.00217519f $X=12.19 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_597 N_VPWR_c_692_n N_A_1263_297#_M1007_d 0.00231264f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_598 N_VPWR_c_692_n N_A_1263_297#_M1016_d 0.00231264f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_599 N_VPWR_c_692_n N_A_1263_297#_M1045_d 0.00231264f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_600 N_VPWR_c_692_n N_A_1263_297#_M1018_s 0.00231264f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_601 N_VPWR_c_692_n N_A_1263_297#_M1029_s 0.00231264f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_602 N_VPWR_c_692_n N_A_1263_297#_M1037_s 0.00242118f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_603 N_VPWR_c_698_n N_A_1263_297#_c_925_n 0.0386815f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_604 N_VPWR_c_692_n N_A_1263_297#_c_925_n 0.0239144f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_605 N_VPWR_c_698_n N_A_1263_297#_c_921_n 0.0191395f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_606 N_VPWR_c_692_n N_A_1263_297#_c_921_n 0.0111641f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_607 N_VPWR_c_698_n N_A_1263_297#_c_927_n 0.0386815f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_608 N_VPWR_c_692_n N_A_1263_297#_c_927_n 0.0239144f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_609 N_VPWR_c_698_n N_A_1263_297#_c_929_n 0.0386815f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_610 N_VPWR_c_692_n N_A_1263_297#_c_929_n 0.0239144f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_611 N_VPWR_c_698_n N_A_1263_297#_c_933_n 0.0386815f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_612 N_VPWR_c_692_n N_A_1263_297#_c_933_n 0.0239144f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_613 N_VPWR_c_698_n N_A_1263_297#_c_935_n 0.0386815f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_614 N_VPWR_c_692_n N_A_1263_297#_c_935_n 0.0239144f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_615 N_VPWR_c_698_n N_A_1263_297#_c_937_n 0.0407825f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_616 N_VPWR_c_692_n N_A_1263_297#_c_937_n 0.0257767f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_617 N_VPWR_c_698_n N_A_1263_297#_c_923_n 0.0175728f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_618 N_VPWR_c_692_n N_A_1263_297#_c_923_n 0.00962271f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_619 N_VPWR_c_698_n N_A_1263_297#_c_965_n 0.0149886f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_620 N_VPWR_c_692_n N_A_1263_297#_c_965_n 0.00962421f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_621 N_VPWR_c_698_n N_A_1263_297#_c_967_n 0.0149886f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_622 N_VPWR_c_692_n N_A_1263_297#_c_967_n 0.00962421f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_623 N_VPWR_c_698_n N_A_1263_297#_c_969_n 0.015002f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_624 N_VPWR_c_692_n N_A_1263_297#_c_969_n 0.00961749f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_625 N_VPWR_c_698_n N_A_1263_297#_c_971_n 0.0149886f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_626 N_VPWR_c_692_n N_A_1263_297#_c_971_n 0.00962421f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_627 N_VPWR_c_698_n N_A_1263_297#_c_973_n 0.0149886f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_628 N_VPWR_c_692_n N_A_1263_297#_c_973_n 0.00962421f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_629 N_VPWR_c_692_n N_Y_M1002_d 0.00232895f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_630 N_VPWR_c_692_n N_Y_M1027_d 0.00232895f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_631 N_VPWR_c_692_n N_Y_M1031_d 0.00232895f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_632 N_A_685_297#_c_832_n N_A_1263_297#_M1001_d 0.00295666f $X=6.785 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_633 N_A_685_297#_c_833_n N_A_1263_297#_M1007_d 0.00187091f $X=7.725 $Y=1.54
+ $X2=0 $Y2=0
cc_634 N_A_685_297#_c_834_n N_A_1263_297#_M1016_d 0.00187091f $X=8.665 $Y=1.54
+ $X2=0 $Y2=0
cc_635 N_A_685_297#_c_832_n N_A_1263_297#_c_920_n 0.0205983f $X=6.785 $Y=1.54
+ $X2=0 $Y2=0
cc_636 N_A_685_297#_M1001_s N_A_1263_297#_c_925_n 0.00352392f $X=6.765 $Y=1.485
+ $X2=0 $Y2=0
cc_637 N_A_685_297#_c_832_n N_A_1263_297#_c_925_n 0.00385532f $X=6.785 $Y=1.54
+ $X2=0 $Y2=0
cc_638 N_A_685_297#_c_833_n N_A_1263_297#_c_925_n 0.00385532f $X=7.725 $Y=1.54
+ $X2=0 $Y2=0
cc_639 N_A_685_297#_c_838_n N_A_1263_297#_c_925_n 0.013395f $X=6.91 $Y=1.62
+ $X2=0 $Y2=0
cc_640 N_A_685_297#_c_833_n N_A_1263_297#_c_983_n 0.0143018f $X=7.725 $Y=1.54
+ $X2=0 $Y2=0
cc_641 N_A_685_297#_M1015_s N_A_1263_297#_c_927_n 0.00352392f $X=7.705 $Y=1.485
+ $X2=0 $Y2=0
cc_642 N_A_685_297#_c_833_n N_A_1263_297#_c_927_n 0.00385532f $X=7.725 $Y=1.54
+ $X2=0 $Y2=0
cc_643 N_A_685_297#_c_834_n N_A_1263_297#_c_927_n 0.00385532f $X=8.665 $Y=1.54
+ $X2=0 $Y2=0
cc_644 N_A_685_297#_c_839_n N_A_1263_297#_c_927_n 0.013395f $X=7.85 $Y=1.62
+ $X2=0 $Y2=0
cc_645 N_A_685_297#_c_834_n N_A_1263_297#_c_988_n 0.0143018f $X=8.665 $Y=1.54
+ $X2=0 $Y2=0
cc_646 N_A_685_297#_M1043_s N_A_1263_297#_c_929_n 0.00352392f $X=8.645 $Y=1.485
+ $X2=0 $Y2=0
cc_647 N_A_685_297#_c_834_n N_A_1263_297#_c_929_n 0.00385532f $X=8.665 $Y=1.54
+ $X2=0 $Y2=0
cc_648 N_A_685_297#_c_840_n N_A_1263_297#_c_929_n 0.013395f $X=8.79 $Y=1.62
+ $X2=0 $Y2=0
cc_649 N_A_685_297#_c_840_n N_A_1263_297#_c_922_n 0.00209545f $X=8.79 $Y=1.62
+ $X2=0 $Y2=0
cc_650 N_A_685_297#_c_832_n N_Y_c_1017_n 0.0315746f $X=6.785 $Y=1.54 $X2=0 $Y2=0
cc_651 N_A_1263_297#_c_933_n N_Y_M1002_d 0.00352392f $X=10.075 $Y=2.38 $X2=0
+ $Y2=0
cc_652 N_A_1263_297#_c_935_n N_Y_M1027_d 0.00352392f $X=11.015 $Y=2.38 $X2=0
+ $Y2=0
cc_653 N_A_1263_297#_c_937_n N_Y_M1031_d 0.00352392f $X=12.005 $Y=2.38 $X2=0
+ $Y2=0
cc_654 N_A_1263_297#_c_922_n N_Y_c_1020_n 0.00929029f $X=9.26 $Y=1.62 $X2=0
+ $Y2=0
cc_655 N_A_1263_297#_M1018_s N_Y_c_1033_n 0.00187091f $X=10.055 $Y=1.485 $X2=0
+ $Y2=0
cc_656 N_A_1263_297#_c_933_n N_Y_c_1033_n 0.00385532f $X=10.075 $Y=2.38 $X2=0
+ $Y2=0
cc_657 N_A_1263_297#_c_999_p N_Y_c_1033_n 0.0143018f $X=10.2 $Y=1.96 $X2=0 $Y2=0
cc_658 N_A_1263_297#_c_935_n N_Y_c_1033_n 0.00385532f $X=11.015 $Y=2.38 $X2=0
+ $Y2=0
cc_659 N_A_1263_297#_M1029_s N_Y_c_1034_n 0.00187091f $X=10.995 $Y=1.485 $X2=0
+ $Y2=0
cc_660 N_A_1263_297#_c_935_n N_Y_c_1034_n 0.00385532f $X=11.015 $Y=2.38 $X2=0
+ $Y2=0
cc_661 N_A_1263_297#_c_1003_p N_Y_c_1034_n 0.0143018f $X=11.14 $Y=1.96 $X2=0
+ $Y2=0
cc_662 N_A_1263_297#_c_937_n N_Y_c_1034_n 0.00342456f $X=12.005 $Y=2.38 $X2=0
+ $Y2=0
cc_663 N_A_1263_297#_c_922_n N_Y_c_1035_n 0.00209545f $X=9.26 $Y=1.62 $X2=0
+ $Y2=0
cc_664 N_A_1263_297#_c_933_n N_Y_c_1035_n 0.013395f $X=10.075 $Y=2.38 $X2=0
+ $Y2=0
cc_665 N_A_1263_297#_c_935_n N_Y_c_1036_n 0.013395f $X=11.015 $Y=2.38 $X2=0
+ $Y2=0
cc_666 N_A_1263_297#_c_937_n N_Y_c_1190_n 0.0203261f $X=12.005 $Y=2.38 $X2=0
+ $Y2=0
cc_667 N_A_1263_297#_c_924_n N_Y_c_1190_n 0.0522181f $X=12.09 $Y=1.62 $X2=0
+ $Y2=0
cc_668 N_A_1263_297#_c_924_n N_VGND_c_1335_n 0.0102366f $X=12.09 $Y=1.62 $X2=0
+ $Y2=0
cc_669 N_Y_c_1011_n N_VGND_M1011_d 0.00274794f $X=1.525 $Y=0.815 $X2=0 $Y2=0
cc_670 N_Y_c_1013_n N_VGND_M1021_d 0.00274794f $X=2.465 $Y=0.815 $X2=0 $Y2=0
cc_671 N_Y_c_1014_n N_VGND_M1034_d 0.00274794f $X=3.405 $Y=0.815 $X2=0 $Y2=0
cc_672 N_Y_c_1015_n N_VGND_M1008_d 0.00274794f $X=4.345 $Y=0.815 $X2=0 $Y2=0
cc_673 N_Y_c_1016_n N_VGND_M1022_d 0.00274794f $X=5.285 $Y=0.815 $X2=0 $Y2=0
cc_674 N_Y_c_1017_n N_VGND_M1046_d 0.0127463f $X=6.745 $Y=0.815 $X2=0 $Y2=0
cc_675 N_Y_c_1018_n N_VGND_M1013_d 0.00274794f $X=7.685 $Y=0.815 $X2=0 $Y2=0
cc_676 N_Y_c_1019_n N_VGND_M1038_d 0.00274794f $X=8.625 $Y=0.815 $X2=0 $Y2=0
cc_677 N_Y_c_1020_n N_VGND_M1044_d 0.00274794f $X=9.565 $Y=0.815 $X2=0 $Y2=0
cc_678 N_Y_c_1021_n N_VGND_M1023_s 0.00274794f $X=10.505 $Y=0.815 $X2=0 $Y2=0
cc_679 N_Y_c_1022_n N_VGND_M1032_s 0.00274794f $X=11.445 $Y=0.815 $X2=0 $Y2=0
cc_680 N_Y_c_1012_n N_VGND_c_1319_n 0.0083648f $X=0.915 $Y=0.815 $X2=0 $Y2=0
cc_681 N_Y_c_1037_n N_VGND_c_1320_n 0.0188551f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_682 N_Y_c_1011_n N_VGND_c_1320_n 0.00198695f $X=1.525 $Y=0.815 $X2=0 $Y2=0
cc_683 N_Y_c_1011_n N_VGND_c_1321_n 0.0201123f $X=1.525 $Y=0.815 $X2=0 $Y2=0
cc_684 N_Y_c_1011_n N_VGND_c_1322_n 0.00198695f $X=1.525 $Y=0.815 $X2=0 $Y2=0
cc_685 N_Y_c_1048_n N_VGND_c_1322_n 0.0188551f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_686 N_Y_c_1013_n N_VGND_c_1322_n 0.00198695f $X=2.465 $Y=0.815 $X2=0 $Y2=0
cc_687 N_Y_c_1013_n N_VGND_c_1323_n 0.0201123f $X=2.465 $Y=0.815 $X2=0 $Y2=0
cc_688 N_Y_c_1013_n N_VGND_c_1324_n 0.00198695f $X=2.465 $Y=0.815 $X2=0 $Y2=0
cc_689 N_Y_c_1056_n N_VGND_c_1324_n 0.0188551f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_690 N_Y_c_1014_n N_VGND_c_1324_n 0.00198695f $X=3.405 $Y=0.815 $X2=0 $Y2=0
cc_691 N_Y_c_1014_n N_VGND_c_1325_n 0.0201123f $X=3.405 $Y=0.815 $X2=0 $Y2=0
cc_692 N_Y_c_1014_n N_VGND_c_1326_n 0.00198695f $X=3.405 $Y=0.815 $X2=0 $Y2=0
cc_693 N_Y_c_1062_n N_VGND_c_1326_n 0.0188551f $X=3.57 $Y=0.39 $X2=0 $Y2=0
cc_694 N_Y_c_1015_n N_VGND_c_1326_n 0.00198695f $X=4.345 $Y=0.815 $X2=0 $Y2=0
cc_695 N_Y_c_1015_n N_VGND_c_1327_n 0.0201123f $X=4.345 $Y=0.815 $X2=0 $Y2=0
cc_696 N_Y_c_1016_n N_VGND_c_1328_n 0.0201123f $X=5.285 $Y=0.815 $X2=0 $Y2=0
cc_697 N_Y_c_1018_n N_VGND_c_1329_n 0.0201123f $X=7.685 $Y=0.815 $X2=0 $Y2=0
cc_698 N_Y_c_1019_n N_VGND_c_1330_n 0.0201123f $X=8.625 $Y=0.815 $X2=0 $Y2=0
cc_699 N_Y_c_1020_n N_VGND_c_1331_n 0.0201123f $X=9.565 $Y=0.815 $X2=0 $Y2=0
cc_700 N_Y_c_1021_n N_VGND_c_1332_n 0.0201123f $X=10.505 $Y=0.815 $X2=0 $Y2=0
cc_701 N_Y_c_1022_n N_VGND_c_1333_n 0.0201123f $X=11.445 $Y=0.815 $X2=0 $Y2=0
cc_702 N_Y_c_1172_n N_VGND_c_1335_n 0.0361363f $X=11.61 $Y=0.39 $X2=0 $Y2=0
cc_703 N_Y_c_1188_n N_VGND_c_1335_n 0.0145666f $X=11.64 $Y=0.815 $X2=0 $Y2=0
cc_704 N_Y_c_1015_n N_VGND_c_1336_n 0.00198695f $X=4.345 $Y=0.815 $X2=0 $Y2=0
cc_705 N_Y_c_1082_n N_VGND_c_1336_n 0.0188551f $X=4.51 $Y=0.39 $X2=0 $Y2=0
cc_706 N_Y_c_1016_n N_VGND_c_1336_n 0.00198695f $X=5.285 $Y=0.815 $X2=0 $Y2=0
cc_707 N_Y_c_1017_n N_VGND_c_1338_n 0.00198695f $X=6.745 $Y=0.815 $X2=0 $Y2=0
cc_708 N_Y_c_1111_n N_VGND_c_1338_n 0.0188551f $X=6.91 $Y=0.39 $X2=0 $Y2=0
cc_709 N_Y_c_1018_n N_VGND_c_1338_n 0.00198695f $X=7.685 $Y=0.815 $X2=0 $Y2=0
cc_710 N_Y_c_1018_n N_VGND_c_1340_n 0.00198695f $X=7.685 $Y=0.815 $X2=0 $Y2=0
cc_711 N_Y_c_1118_n N_VGND_c_1340_n 0.0188551f $X=7.85 $Y=0.39 $X2=0 $Y2=0
cc_712 N_Y_c_1019_n N_VGND_c_1340_n 0.00198695f $X=8.625 $Y=0.815 $X2=0 $Y2=0
cc_713 N_Y_c_1019_n N_VGND_c_1342_n 0.00198695f $X=8.625 $Y=0.815 $X2=0 $Y2=0
cc_714 N_Y_c_1126_n N_VGND_c_1342_n 0.0188551f $X=8.79 $Y=0.39 $X2=0 $Y2=0
cc_715 N_Y_c_1020_n N_VGND_c_1342_n 0.00198695f $X=9.565 $Y=0.815 $X2=0 $Y2=0
cc_716 N_Y_c_1020_n N_VGND_c_1344_n 0.00198695f $X=9.565 $Y=0.815 $X2=0 $Y2=0
cc_717 N_Y_c_1132_n N_VGND_c_1344_n 0.0188551f $X=9.73 $Y=0.39 $X2=0 $Y2=0
cc_718 N_Y_c_1021_n N_VGND_c_1344_n 0.00198695f $X=10.505 $Y=0.815 $X2=0 $Y2=0
cc_719 N_Y_c_1021_n N_VGND_c_1346_n 0.00198695f $X=10.505 $Y=0.815 $X2=0 $Y2=0
cc_720 N_Y_c_1160_n N_VGND_c_1346_n 0.0188551f $X=10.67 $Y=0.39 $X2=0 $Y2=0
cc_721 N_Y_c_1022_n N_VGND_c_1346_n 0.00198695f $X=11.445 $Y=0.815 $X2=0 $Y2=0
cc_722 N_Y_c_1022_n N_VGND_c_1348_n 0.00198695f $X=11.445 $Y=0.815 $X2=0 $Y2=0
cc_723 N_Y_c_1172_n N_VGND_c_1348_n 0.0229947f $X=11.61 $Y=0.39 $X2=0 $Y2=0
cc_724 N_Y_c_1016_n N_VGND_c_1353_n 0.00198695f $X=5.285 $Y=0.815 $X2=0 $Y2=0
cc_725 N_Y_c_1090_n N_VGND_c_1353_n 0.0188551f $X=5.45 $Y=0.39 $X2=0 $Y2=0
cc_726 N_Y_c_1017_n N_VGND_c_1353_n 0.00198695f $X=6.745 $Y=0.815 $X2=0 $Y2=0
cc_727 N_Y_c_1017_n N_VGND_c_1354_n 0.0606502f $X=6.745 $Y=0.815 $X2=0 $Y2=0
cc_728 N_Y_M1006_s N_VGND_c_1355_n 0.00215201f $X=0.615 $Y=0.235 $X2=0 $Y2=0
cc_729 N_Y_M1019_s N_VGND_c_1355_n 0.00215201f $X=1.555 $Y=0.235 $X2=0 $Y2=0
cc_730 N_Y_M1026_s N_VGND_c_1355_n 0.00215201f $X=2.495 $Y=0.235 $X2=0 $Y2=0
cc_731 N_Y_M1003_s N_VGND_c_1355_n 0.00215201f $X=3.435 $Y=0.235 $X2=0 $Y2=0
cc_732 N_Y_M1012_s N_VGND_c_1355_n 0.00215201f $X=4.375 $Y=0.235 $X2=0 $Y2=0
cc_733 N_Y_M1036_s N_VGND_c_1355_n 0.00215201f $X=5.315 $Y=0.235 $X2=0 $Y2=0
cc_734 N_Y_M1010_s N_VGND_c_1355_n 0.00215201f $X=6.775 $Y=0.235 $X2=0 $Y2=0
cc_735 N_Y_M1028_s N_VGND_c_1355_n 0.00215201f $X=7.715 $Y=0.235 $X2=0 $Y2=0
cc_736 N_Y_M1039_s N_VGND_c_1355_n 0.00215201f $X=8.655 $Y=0.235 $X2=0 $Y2=0
cc_737 N_Y_M1004_d N_VGND_c_1355_n 0.00215201f $X=9.595 $Y=0.235 $X2=0 $Y2=0
cc_738 N_Y_M1025_d N_VGND_c_1355_n 0.00215201f $X=10.535 $Y=0.235 $X2=0 $Y2=0
cc_739 N_Y_M1041_d N_VGND_c_1355_n 0.00215201f $X=11.475 $Y=0.235 $X2=0 $Y2=0
cc_740 N_Y_c_1037_n N_VGND_c_1355_n 0.0122069f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_741 N_Y_c_1011_n N_VGND_c_1355_n 0.00874058f $X=1.525 $Y=0.815 $X2=0 $Y2=0
cc_742 N_Y_c_1048_n N_VGND_c_1355_n 0.0122069f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_743 N_Y_c_1013_n N_VGND_c_1355_n 0.00874058f $X=2.465 $Y=0.815 $X2=0 $Y2=0
cc_744 N_Y_c_1056_n N_VGND_c_1355_n 0.0122069f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_745 N_Y_c_1014_n N_VGND_c_1355_n 0.00874058f $X=3.405 $Y=0.815 $X2=0 $Y2=0
cc_746 N_Y_c_1062_n N_VGND_c_1355_n 0.0122069f $X=3.57 $Y=0.39 $X2=0 $Y2=0
cc_747 N_Y_c_1015_n N_VGND_c_1355_n 0.00874058f $X=4.345 $Y=0.815 $X2=0 $Y2=0
cc_748 N_Y_c_1082_n N_VGND_c_1355_n 0.0122069f $X=4.51 $Y=0.39 $X2=0 $Y2=0
cc_749 N_Y_c_1016_n N_VGND_c_1355_n 0.00874058f $X=5.285 $Y=0.815 $X2=0 $Y2=0
cc_750 N_Y_c_1090_n N_VGND_c_1355_n 0.0122069f $X=5.45 $Y=0.39 $X2=0 $Y2=0
cc_751 N_Y_c_1017_n N_VGND_c_1355_n 0.0107088f $X=6.745 $Y=0.815 $X2=0 $Y2=0
cc_752 N_Y_c_1111_n N_VGND_c_1355_n 0.0122069f $X=6.91 $Y=0.39 $X2=0 $Y2=0
cc_753 N_Y_c_1018_n N_VGND_c_1355_n 0.00874058f $X=7.685 $Y=0.815 $X2=0 $Y2=0
cc_754 N_Y_c_1118_n N_VGND_c_1355_n 0.0122069f $X=7.85 $Y=0.39 $X2=0 $Y2=0
cc_755 N_Y_c_1019_n N_VGND_c_1355_n 0.00874058f $X=8.625 $Y=0.815 $X2=0 $Y2=0
cc_756 N_Y_c_1126_n N_VGND_c_1355_n 0.0122069f $X=8.79 $Y=0.39 $X2=0 $Y2=0
cc_757 N_Y_c_1020_n N_VGND_c_1355_n 0.00874058f $X=9.565 $Y=0.815 $X2=0 $Y2=0
cc_758 N_Y_c_1132_n N_VGND_c_1355_n 0.0122069f $X=9.73 $Y=0.39 $X2=0 $Y2=0
cc_759 N_Y_c_1021_n N_VGND_c_1355_n 0.00874058f $X=10.505 $Y=0.815 $X2=0 $Y2=0
cc_760 N_Y_c_1160_n N_VGND_c_1355_n 0.0122069f $X=10.67 $Y=0.39 $X2=0 $Y2=0
cc_761 N_Y_c_1022_n N_VGND_c_1355_n 0.00874058f $X=11.445 $Y=0.815 $X2=0 $Y2=0
cc_762 N_Y_c_1172_n N_VGND_c_1355_n 0.014258f $X=11.61 $Y=0.39 $X2=0 $Y2=0
