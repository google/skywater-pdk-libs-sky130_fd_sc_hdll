# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a21bo_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21bo_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.885000 0.995000 3.085000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.375000 0.995000 3.665000 1.615000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225000 0.995000 1.695000 1.325000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.547000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 0.715000 0.900000 0.885000 ;
        RECT 0.110000 0.885000 0.380000 1.835000 ;
        RECT 0.110000 1.835000 0.900000 2.005000 ;
        RECT 0.520000 0.315000 0.900000 0.715000 ;
        RECT 0.645000 2.005000 0.900000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.085000 0.345000 0.545000 ;
      RECT 0.090000  2.255000 0.425000 2.635000 ;
      RECT 0.620000  1.075000 0.950000 1.495000 ;
      RECT 0.620000  1.495000 1.385000 1.665000 ;
      RECT 1.070000  0.085000 1.400000 0.785000 ;
      RECT 1.140000  2.275000 1.470000 2.635000 ;
      RECT 1.215000  1.665000 1.385000 1.895000 ;
      RECT 1.215000  1.895000 2.375000 2.105000 ;
      RECT 1.555000  1.555000 2.035000 1.725000 ;
      RECT 1.605000  0.655000 2.035000 0.825000 ;
      RECT 1.865000  0.825000 2.035000 0.995000 ;
      RECT 1.865000  0.995000 2.325000 1.325000 ;
      RECT 1.865000  1.325000 2.035000 1.555000 ;
      RECT 2.125000  0.085000 2.455000 0.465000 ;
      RECT 2.125000  2.105000 2.375000 2.465000 ;
      RECT 2.205000  1.505000 2.715000 1.675000 ;
      RECT 2.205000  1.675000 2.375000 1.895000 ;
      RECT 2.495000  0.635000 2.940000 0.825000 ;
      RECT 2.495000  0.825000 2.715000 1.505000 ;
      RECT 2.545000  1.845000 3.875000 2.015000 ;
      RECT 2.545000  2.015000 2.925000 2.465000 ;
      RECT 3.155000  2.185000 3.325000 2.635000 ;
      RECT 3.495000  0.085000 3.875000 0.825000 ;
      RECT 3.495000  2.015000 3.875000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21bo_2
