* File: sky130_fd_sc_hdll__decap_8.pxi.spice
* Created: Wed Sep  2 08:27:53 2020
* 
x_PM_SKY130_FD_SC_HDLL__DECAP_8%VGND N_VGND_M1001_s N_VGND_M1000_g N_VGND_c_16_n
+ N_VGND_c_17_n VGND N_VGND_c_18_n N_VGND_c_19_n N_VGND_c_20_n
+ PM_SKY130_FD_SC_HDLL__DECAP_8%VGND
x_PM_SKY130_FD_SC_HDLL__DECAP_8%VPWR N_VPWR_M1000_s N_VPWR_M1001_g N_VPWR_c_42_n
+ N_VPWR_c_43_n VPWR N_VPWR_c_38_n N_VPWR_c_39_n N_VPWR_c_40_n N_VPWR_c_41_n
+ PM_SKY130_FD_SC_HDLL__DECAP_8%VPWR
cc_1 VNB N_VGND_c_16_n 0.0184325f $X=-0.19 $Y=-0.24 $X2=3.125 $Y2=0.385
cc_2 VNB N_VGND_c_17_n 0.0803708f $X=-0.19 $Y=-0.24 $X2=1.735 $Y2=0.385
cc_3 VNB N_VGND_c_18_n 0.0461317f $X=-0.19 $Y=-0.24 $X2=1.715 $Y2=1.87
cc_4 VNB N_VGND_c_19_n 0.0439751f $X=-0.19 $Y=-0.24 $X2=3.42 $Y2=0.475
cc_5 VNB N_VGND_c_20_n 0.19806f $X=-0.19 $Y=-0.24 $X2=3.45 $Y2=0
cc_6 VNB N_VPWR_c_38_n 0.112251f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_VPWR_c_39_n 0.171259f $X=-0.19 $Y=-0.24 $X2=1.55 $Y2=1.29
cc_8 VNB N_VPWR_c_40_n 0.0178259f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=0
cc_9 VNB N_VPWR_c_41_n 0.155873f $X=-0.19 $Y=-0.24 $X2=3.42 $Y2=0.475
cc_10 VPB N_VGND_c_17_n 0.0068688f $X=-0.19 $Y=1.305 $X2=1.735 $Y2=0.385
cc_11 VPB N_VGND_c_18_n 0.23585f $X=-0.19 $Y=1.305 $X2=1.715 $Y2=1.87
cc_12 VPB N_VPWR_c_42_n 0.0157765f $X=-0.19 $Y=1.305 $X2=3.125 $Y2=0.385
cc_13 VPB N_VPWR_c_43_n 0.0597303f $X=-0.19 $Y=1.305 $X2=1.735 $Y2=0.385
cc_14 VPB N_VPWR_c_40_n 0.083571f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=0
cc_15 VPB N_VPWR_c_41_n 0.0421815f $X=-0.19 $Y=1.305 $X2=3.42 $Y2=0.475
cc_16 N_VGND_c_17_n N_VPWR_c_42_n 0.0859391f $X=1.735 $Y=0.385 $X2=0 $Y2=0
cc_17 N_VGND_c_18_n N_VPWR_c_42_n 0.158744f $X=1.715 $Y=1.87 $X2=0 $Y2=0
cc_18 N_VGND_c_17_n N_VPWR_c_43_n 0.0561345f $X=1.735 $Y=0.385 $X2=0 $Y2=0
cc_19 N_VGND_c_18_n N_VPWR_c_43_n 0.0493583f $X=1.715 $Y=1.87 $X2=0 $Y2=0
cc_20 N_VGND_c_16_n N_VPWR_c_38_n 0.0203068f $X=3.125 $Y=0.385 $X2=0 $Y2=0
cc_21 N_VGND_c_17_n N_VPWR_c_38_n 0.150639f $X=1.735 $Y=0.385 $X2=0 $Y2=0
cc_22 N_VGND_c_18_n N_VPWR_c_38_n 0.0905513f $X=1.715 $Y=1.87 $X2=0 $Y2=0
cc_23 N_VGND_c_16_n N_VPWR_c_39_n 0.123224f $X=3.125 $Y=0.385 $X2=0 $Y2=0
cc_24 N_VGND_c_17_n N_VPWR_c_39_n 0.00648593f $X=1.735 $Y=0.385 $X2=0 $Y2=0
cc_25 N_VGND_c_18_n N_VPWR_c_39_n 0.0987678f $X=1.715 $Y=1.87 $X2=0 $Y2=0
cc_26 N_VGND_c_19_n N_VPWR_c_39_n 0.0237188f $X=3.42 $Y=0.475 $X2=0 $Y2=0
cc_27 N_VGND_c_16_n N_VPWR_c_40_n 0.102789f $X=3.125 $Y=0.385 $X2=0 $Y2=0
cc_28 N_VGND_c_17_n N_VPWR_c_40_n 0.0327855f $X=1.735 $Y=0.385 $X2=0 $Y2=0
cc_29 N_VGND_c_18_n N_VPWR_c_40_n 0.202395f $X=1.715 $Y=1.87 $X2=0 $Y2=0
cc_30 N_VGND_c_19_n N_VPWR_c_40_n 0.0425904f $X=3.42 $Y=0.475 $X2=0 $Y2=0
