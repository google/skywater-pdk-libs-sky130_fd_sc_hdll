* NGSPICE file created from sky130_fd_sc_hdll__and4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
M1000 a_503_47# a_27_47# a_184_21# VNB nshort w=420000u l=150000u
+  ad=1.449e+11p pd=1.53e+06u as=1.092e+11p ps=1.36e+06u
M1001 VPWR D a_184_21# VPB phighvt w=420000u l=180000u
+  ad=1.299e+12p pd=9.38e+06u as=2.562e+11p ps=2.9e+06u
M1002 VPWR A_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1003 a_184_21# C VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_602_47# a_545_280# a_503_47# VNB nshort w=420000u l=150000u
+  ad=1.407e+11p pd=1.51e+06u as=0p ps=0u
M1005 VGND D a_699_47# VNB nshort w=420000u l=150000u
+  ad=6.1255e+11p pd=5.76e+06u as=1.134e+11p ps=1.38e+06u
M1006 a_699_47# C a_602_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_545_280# B_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1008 a_184_21# a_27_47# VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_545_280# a_184_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_184_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1011 VGND A_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1012 VGND a_184_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1013 X a_184_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_545_280# B_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1015 X a_184_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

