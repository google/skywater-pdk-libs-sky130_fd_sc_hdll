# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__or4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.840000 0.995000 3.595000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.705000 2.125000 3.395000 2.455000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.995000 0.830000 1.695000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 0.995000 1.340000 1.325000 ;
    END
  END D_N
  PIN VGND
    ANTENNADIFFAREA  0.812100 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  0.859325 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.155000 0.415000 4.455000 0.760000 ;
        RECT 4.155000 1.495000 4.455000 2.465000 ;
        RECT 4.260000 0.760000 4.455000 1.495000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.450000 0.405000 0.825000 ;
      RECT 0.085000  0.825000 0.260000 1.865000 ;
      RECT 0.085000  1.865000 2.040000 2.035000 ;
      RECT 0.085000  2.035000 0.345000 2.455000 ;
      RECT 0.515000  2.205000 0.895000 2.635000 ;
      RECT 0.710000  0.085000 0.880000 0.825000 ;
      RECT 1.045000  1.525000 1.700000 1.695000 ;
      RECT 1.180000  0.450000 1.350000 0.655000 ;
      RECT 1.180000  0.655000 1.700000 0.825000 ;
      RECT 1.510000  0.825000 1.700000 1.075000 ;
      RECT 1.510000  1.075000 1.955000 1.245000 ;
      RECT 1.510000  1.245000 1.700000 1.525000 ;
      RECT 1.595000  0.085000 1.970000 0.485000 ;
      RECT 1.635000  2.205000 2.430000 2.375000 ;
      RECT 1.870000  1.415000 2.570000 1.585000 ;
      RECT 1.870000  1.585000 2.040000 1.865000 ;
      RECT 2.190000  0.305000 2.360000 0.655000 ;
      RECT 2.190000  0.655000 3.935000 0.825000 ;
      RECT 2.260000  1.785000 3.395000 1.955000 ;
      RECT 2.260000  1.955000 2.430000 2.205000 ;
      RECT 2.400000  0.995000 2.570000 1.415000 ;
      RECT 2.545000  0.085000 2.925000 0.485000 ;
      RECT 3.145000  0.305000 3.315000 0.655000 ;
      RECT 3.225000  1.495000 3.935000 1.665000 ;
      RECT 3.225000  1.665000 3.395000 1.785000 ;
      RECT 3.485000  0.085000 3.915000 0.485000 ;
      RECT 3.615000  1.835000 3.895000 2.635000 ;
      RECT 3.765000  0.825000 3.935000 0.995000 ;
      RECT 3.765000  0.995000 4.040000 1.325000 ;
      RECT 3.765000  1.325000 3.935000 1.495000 ;
      RECT 4.650000  0.085000 4.820000 0.915000 ;
      RECT 4.650000  1.440000 4.820000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4bb_2
