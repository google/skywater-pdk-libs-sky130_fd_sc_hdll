* File: sky130_fd_sc_hdll__a31o_1.spice
* Created: Wed Sep  2 08:19:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a31o_1.pex.spice"
.subckt sky130_fd_sc_hdll__a31o_1  VNB VPB A3 A2 A1 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_80_21#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.125125 AS=0.17225 PD=1.035 PS=1.83 NRD=14.76 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1008 A_217_47# N_A3_M1008_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65 AD=0.1235
+ AS=0.125125 PD=1.03 PS=1.035 NRD=24.912 NRS=4.608 M=1 R=4.33333 SA=75000.7
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1006 A_323_47# N_A2_M1006_g A_217_47# VNB NSHORT L=0.15 W=0.65 AD=0.1235
+ AS=0.1235 PD=1.03 PS=1.03 NRD=24.912 NRS=24.912 M=1 R=4.33333 SA=75001.3
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1007 N_A_80_21#_M1007_d N_A1_M1007_g A_323_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.1235 PD=1.03 PS=1.03 NRD=10.152 NRS=24.912 M=1 R=4.33333
+ SA=75001.8 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_B1_M1000_g N_A_80_21#_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2405 AS=0.1235 PD=2.04 PS=1.03 NRD=13.836 NRS=8.304 M=1 R=4.33333
+ SA=75002.3 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_80_21#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1775 AS=0.275 PD=1.355 PS=2.55 NRD=7.8603 NRS=1.9503 M=1 R=5.55556
+ SA=90000.2 SB=90002.4 A=0.18 P=2.36 MULT=1
MM1005 N_A_225_297#_M1005_d N_A3_M1005_g N_VPWR_M1003_d VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.1775 PD=1.35 PS=1.355 NRD=6.8753 NRS=6.8753 M=1 R=5.55556
+ SA=90000.7 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A2_M1001_g N_A_225_297#_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=6.8753 NRS=6.8753 M=1 R=5.55556
+ SA=90001.2 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1002 N_A_225_297#_M1002_d N_A1_M1002_g N_VPWR_M1001_d VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=6.8753 NRS=6.8753 M=1 R=5.55556
+ SA=90001.8 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1009 N_A_80_21#_M1009_d N_B1_M1009_g N_A_225_297#_M1002_d VPB PHIGHVT L=0.18
+ W=1 AD=0.33 AS=0.175 PD=2.66 PS=1.35 NRD=12.7853 NRS=6.8753 M=1 R=5.55556
+ SA=90002.3 SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
c_52 VPB 0 1.20528e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__a31o_1.pxi.spice"
*
.ends
*
*
