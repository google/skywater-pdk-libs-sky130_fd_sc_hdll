* File: sky130_fd_sc_hdll__nor4_6.pex.spice
* Created: Thu Aug 27 19:17:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR4_6%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 37 54 55
r106 55 56 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=2.84 $Y=1.202
+ $X2=2.865 $Y2=1.202
r107 53 55 16.9351 $w=3.7e-07 $l=1.3e-07 $layer=POLY_cond $X=2.71 $Y=1.202
+ $X2=2.84 $Y2=1.202
r108 53 54 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=2.71
+ $Y=1.16 $X2=2.71 $Y2=1.16
r109 51 53 37.7784 $w=3.7e-07 $l=2.9e-07 $layer=POLY_cond $X=2.42 $Y=1.202
+ $X2=2.71 $Y2=1.202
r110 50 51 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=2.395 $Y=1.202
+ $X2=2.42 $Y2=1.202
r111 49 50 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=1.925 $Y=1.202
+ $X2=2.395 $Y2=1.202
r112 48 49 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.9 $Y=1.202
+ $X2=1.925 $Y2=1.202
r113 47 48 54.7135 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=1.48 $Y=1.202
+ $X2=1.9 $Y2=1.202
r114 46 47 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.48 $Y2=1.202
r115 45 46 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.455 $Y2=1.202
r116 44 45 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.96 $Y=1.202
+ $X2=0.985 $Y2=1.202
r117 42 44 37.7784 $w=3.7e-07 $l=2.9e-07 $layer=POLY_cond $X=0.67 $Y=1.202
+ $X2=0.96 $Y2=1.202
r118 42 43 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=0.67
+ $Y=1.16 $X2=0.67 $Y2=1.16
r119 40 42 16.9351 $w=3.7e-07 $l=1.3e-07 $layer=POLY_cond $X=0.54 $Y=1.202
+ $X2=0.67 $Y2=1.202
r120 39 40 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.54 $Y2=1.202
r121 37 54 58.0952 $w=2.08e-07 $l=1.1e-06 $layer=LI1_cond $X=1.61 $Y=1.18
+ $X2=2.71 $Y2=1.18
r122 37 43 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=1.61 $Y=1.18
+ $X2=0.67 $Y2=1.18
r123 34 56 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.865 $Y=1.41
+ $X2=2.865 $Y2=1.202
r124 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.865 $Y=1.41
+ $X2=2.865 $Y2=1.985
r125 31 55 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.84 $Y=0.995
+ $X2=2.84 $Y2=1.202
r126 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.84 $Y=0.995
+ $X2=2.84 $Y2=0.56
r127 28 51 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.42 $Y=0.995
+ $X2=2.42 $Y2=1.202
r128 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.42 $Y=0.995
+ $X2=2.42 $Y2=0.56
r129 25 50 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.202
r130 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.985
r131 22 49 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r132 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r133 19 48 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.9 $Y=0.995
+ $X2=1.9 $Y2=1.202
r134 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.9 $Y=0.995
+ $X2=1.9 $Y2=0.56
r135 16 47 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.48 $Y=0.995
+ $X2=1.48 $Y2=1.202
r136 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.48 $Y=0.995
+ $X2=1.48 $Y2=0.56
r137 13 46 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r138 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r139 10 45 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r140 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r141 7 44 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=0.96 $Y2=1.202
r142 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=0.96 $Y2=0.56
r143 4 40 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.54 $Y2=1.202
r144 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.54 $Y2=0.56
r145 1 39 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r146 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_6%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 37 54 55
r112 55 56 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.66 $Y=1.202
+ $X2=5.685 $Y2=1.202
r113 53 55 16.9351 $w=3.7e-07 $l=1.3e-07 $layer=POLY_cond $X=5.53 $Y=1.202
+ $X2=5.66 $Y2=1.202
r114 53 54 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=5.53
+ $Y=1.16 $X2=5.53 $Y2=1.16
r115 51 53 37.7784 $w=3.7e-07 $l=2.9e-07 $layer=POLY_cond $X=5.24 $Y=1.202
+ $X2=5.53 $Y2=1.202
r116 50 51 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.215 $Y=1.202
+ $X2=5.24 $Y2=1.202
r117 49 50 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=4.745 $Y=1.202
+ $X2=5.215 $Y2=1.202
r118 48 49 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=4.72 $Y=1.202
+ $X2=4.745 $Y2=1.202
r119 47 48 54.7135 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.3 $Y=1.202
+ $X2=4.72 $Y2=1.202
r120 46 47 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=4.275 $Y=1.202
+ $X2=4.3 $Y2=1.202
r121 45 46 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=3.805 $Y=1.202
+ $X2=4.275 $Y2=1.202
r122 44 45 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=3.78 $Y=1.202
+ $X2=3.805 $Y2=1.202
r123 42 44 37.7784 $w=3.7e-07 $l=2.9e-07 $layer=POLY_cond $X=3.49 $Y=1.202
+ $X2=3.78 $Y2=1.202
r124 42 43 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=3.49
+ $Y=1.16 $X2=3.49 $Y2=1.16
r125 40 42 16.9351 $w=3.7e-07 $l=1.3e-07 $layer=POLY_cond $X=3.36 $Y=1.202
+ $X2=3.49 $Y2=1.202
r126 39 40 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=3.335 $Y=1.202
+ $X2=3.36 $Y2=1.202
r127 37 54 61.2641 $w=2.08e-07 $l=1.16e-06 $layer=LI1_cond $X=4.37 $Y=1.18
+ $X2=5.53 $Y2=1.18
r128 37 43 46.4762 $w=2.08e-07 $l=8.8e-07 $layer=LI1_cond $X=4.37 $Y=1.18
+ $X2=3.49 $Y2=1.18
r129 34 56 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.685 $Y=1.41
+ $X2=5.685 $Y2=1.202
r130 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.685 $Y=1.41
+ $X2=5.685 $Y2=1.985
r131 31 55 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.66 $Y=0.995
+ $X2=5.66 $Y2=1.202
r132 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.66 $Y=0.995
+ $X2=5.66 $Y2=0.56
r133 28 51 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=1.202
r134 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=0.56
r135 25 50 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.215 $Y=1.41
+ $X2=5.215 $Y2=1.202
r136 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.215 $Y=1.41
+ $X2=5.215 $Y2=1.985
r137 22 49 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.745 $Y=1.41
+ $X2=4.745 $Y2=1.202
r138 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.745 $Y=1.41
+ $X2=4.745 $Y2=1.985
r139 19 48 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.72 $Y=0.995
+ $X2=4.72 $Y2=1.202
r140 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.72 $Y=0.995
+ $X2=4.72 $Y2=0.56
r141 16 47 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.3 $Y=0.995
+ $X2=4.3 $Y2=1.202
r142 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.3 $Y=0.995
+ $X2=4.3 $Y2=0.56
r143 13 46 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.275 $Y=1.41
+ $X2=4.275 $Y2=1.202
r144 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.275 $Y=1.41
+ $X2=4.275 $Y2=1.985
r145 10 45 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.805 $Y=1.41
+ $X2=3.805 $Y2=1.202
r146 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.805 $Y=1.41
+ $X2=3.805 $Y2=1.985
r147 7 44 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.78 $Y=0.995
+ $X2=3.78 $Y2=1.202
r148 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.78 $Y=0.995
+ $X2=3.78 $Y2=0.56
r149 4 40 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.36 $Y=0.995
+ $X2=3.36 $Y2=1.202
r150 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.36 $Y=0.995
+ $X2=3.36 $Y2=0.56
r151 1 39 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.335 $Y=1.41
+ $X2=3.335 $Y2=1.202
r152 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.335 $Y=1.41
+ $X2=3.335 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_6%C 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 37 54 55 60
r112 55 56 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=9 $Y=1.202
+ $X2=9.025 $Y2=1.202
r113 53 55 16.9351 $w=3.7e-07 $l=1.3e-07 $layer=POLY_cond $X=8.87 $Y=1.202 $X2=9
+ $Y2=1.202
r114 53 54 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=8.87
+ $Y=1.16 $X2=8.87 $Y2=1.16
r115 51 53 37.7784 $w=3.7e-07 $l=2.9e-07 $layer=POLY_cond $X=8.58 $Y=1.202
+ $X2=8.87 $Y2=1.202
r116 50 51 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=8.555 $Y=1.202
+ $X2=8.58 $Y2=1.202
r117 49 50 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=8.085 $Y=1.202
+ $X2=8.555 $Y2=1.202
r118 48 49 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=8.06 $Y=1.202
+ $X2=8.085 $Y2=1.202
r119 47 48 54.7135 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=7.64 $Y=1.202
+ $X2=8.06 $Y2=1.202
r120 46 47 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=7.615 $Y=1.202
+ $X2=7.64 $Y2=1.202
r121 45 46 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=7.145 $Y=1.202
+ $X2=7.615 $Y2=1.202
r122 44 45 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=7.12 $Y=1.202
+ $X2=7.145 $Y2=1.202
r123 43 60 64.1688 $w=2.08e-07 $l=1.215e-06 $layer=LI1_cond $X=6.83 $Y=1.18
+ $X2=8.045 $Y2=1.18
r124 42 44 37.7784 $w=3.7e-07 $l=2.9e-07 $layer=POLY_cond $X=6.83 $Y=1.202
+ $X2=7.12 $Y2=1.202
r125 42 43 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=6.83
+ $Y=1.16 $X2=6.83 $Y2=1.16
r126 40 42 16.9351 $w=3.7e-07 $l=1.3e-07 $layer=POLY_cond $X=6.7 $Y=1.202
+ $X2=6.83 $Y2=1.202
r127 39 40 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=6.675 $Y=1.202
+ $X2=6.7 $Y2=1.202
r128 37 54 43.3074 $w=2.08e-07 $l=8.2e-07 $layer=LI1_cond $X=8.05 $Y=1.18
+ $X2=8.87 $Y2=1.18
r129 37 60 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=8.05 $Y=1.18
+ $X2=8.045 $Y2=1.18
r130 34 56 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.025 $Y=1.41
+ $X2=9.025 $Y2=1.202
r131 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.025 $Y=1.41
+ $X2=9.025 $Y2=1.985
r132 31 55 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9 $Y=0.995 $X2=9
+ $Y2=1.202
r133 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9 $Y=0.995 $X2=9
+ $Y2=0.56
r134 28 51 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.58 $Y=0.995
+ $X2=8.58 $Y2=1.202
r135 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.58 $Y=0.995
+ $X2=8.58 $Y2=0.56
r136 25 50 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.555 $Y=1.41
+ $X2=8.555 $Y2=1.202
r137 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.555 $Y=1.41
+ $X2=8.555 $Y2=1.985
r138 22 49 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.085 $Y=1.41
+ $X2=8.085 $Y2=1.202
r139 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.085 $Y=1.41
+ $X2=8.085 $Y2=1.985
r140 19 48 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.06 $Y=0.995
+ $X2=8.06 $Y2=1.202
r141 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.06 $Y=0.995
+ $X2=8.06 $Y2=0.56
r142 16 47 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.64 $Y=0.995
+ $X2=7.64 $Y2=1.202
r143 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.64 $Y=0.995
+ $X2=7.64 $Y2=0.56
r144 13 46 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.615 $Y=1.41
+ $X2=7.615 $Y2=1.202
r145 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.615 $Y=1.41
+ $X2=7.615 $Y2=1.985
r146 10 45 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.145 $Y=1.41
+ $X2=7.145 $Y2=1.202
r147 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.145 $Y=1.41
+ $X2=7.145 $Y2=1.985
r148 7 44 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.12 $Y=0.995
+ $X2=7.12 $Y2=1.202
r149 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.12 $Y=0.995
+ $X2=7.12 $Y2=0.56
r150 4 40 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.7 $Y=0.995
+ $X2=6.7 $Y2=1.202
r151 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.7 $Y=0.995 $X2=6.7
+ $Y2=0.56
r152 1 39 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.675 $Y=1.41
+ $X2=6.675 $Y2=1.202
r153 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.675 $Y=1.41
+ $X2=6.675 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_6%D 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 37 52 55
r115 55 56 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=11.82 $Y=1.202
+ $X2=11.845 $Y2=1.202
r116 54 55 54.7135 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=11.4 $Y=1.202
+ $X2=11.82 $Y2=1.202
r117 53 54 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=11.375 $Y=1.202
+ $X2=11.4 $Y2=1.202
r118 51 53 59.273 $w=3.7e-07 $l=4.55e-07 $layer=POLY_cond $X=10.92 $Y=1.202
+ $X2=11.375 $Y2=1.202
r119 51 52 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=10.92
+ $Y=1.16 $X2=10.92 $Y2=1.16
r120 49 51 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=10.905 $Y=1.202
+ $X2=10.92 $Y2=1.202
r121 48 49 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=10.88 $Y=1.202
+ $X2=10.905 $Y2=1.202
r122 47 48 54.7135 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=10.46 $Y=1.202
+ $X2=10.88 $Y2=1.202
r123 46 47 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=10.435 $Y=1.202
+ $X2=10.46 $Y2=1.202
r124 45 46 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=9.965 $Y=1.202
+ $X2=10.435 $Y2=1.202
r125 44 45 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=9.94 $Y=1.202
+ $X2=9.965 $Y2=1.202
r126 42 44 49.5027 $w=3.7e-07 $l=3.8e-07 $layer=POLY_cond $X=9.56 $Y=1.202
+ $X2=9.94 $Y2=1.202
r127 42 43 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=9.56
+ $Y=1.16 $X2=9.56 $Y2=1.16
r128 40 42 5.21081 $w=3.7e-07 $l=4e-08 $layer=POLY_cond $X=9.52 $Y=1.202
+ $X2=9.56 $Y2=1.202
r129 39 40 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=9.495 $Y=1.202
+ $X2=9.52 $Y2=1.202
r130 37 52 30.1039 $w=2.08e-07 $l=5.7e-07 $layer=LI1_cond $X=10.35 $Y=1.18
+ $X2=10.92 $Y2=1.18
r131 37 43 41.7229 $w=2.08e-07 $l=7.9e-07 $layer=LI1_cond $X=10.35 $Y=1.18
+ $X2=9.56 $Y2=1.18
r132 34 56 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=11.845 $Y=1.41
+ $X2=11.845 $Y2=1.202
r133 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.845 $Y=1.41
+ $X2=11.845 $Y2=1.985
r134 31 55 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.82 $Y=0.995
+ $X2=11.82 $Y2=1.202
r135 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.82 $Y=0.995
+ $X2=11.82 $Y2=0.56
r136 28 54 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.4 $Y=0.995
+ $X2=11.4 $Y2=1.202
r137 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.4 $Y=0.995
+ $X2=11.4 $Y2=0.56
r138 25 53 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=11.375 $Y=1.41
+ $X2=11.375 $Y2=1.202
r139 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.375 $Y=1.41
+ $X2=11.375 $Y2=1.985
r140 22 49 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.905 $Y=1.41
+ $X2=10.905 $Y2=1.202
r141 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.905 $Y=1.41
+ $X2=10.905 $Y2=1.985
r142 19 48 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.88 $Y=0.995
+ $X2=10.88 $Y2=1.202
r143 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.88 $Y=0.995
+ $X2=10.88 $Y2=0.56
r144 16 47 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.46 $Y=0.995
+ $X2=10.46 $Y2=1.202
r145 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.46 $Y=0.995
+ $X2=10.46 $Y2=0.56
r146 13 46 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.435 $Y=1.41
+ $X2=10.435 $Y2=1.202
r147 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.435 $Y=1.41
+ $X2=10.435 $Y2=1.985
r148 10 45 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.965 $Y=1.41
+ $X2=9.965 $Y2=1.202
r149 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.965 $Y=1.41
+ $X2=9.965 $Y2=1.985
r150 7 44 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.94 $Y=0.995
+ $X2=9.94 $Y2=1.202
r151 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.94 $Y=0.995
+ $X2=9.94 $Y2=0.56
r152 4 40 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.52 $Y=0.995
+ $X2=9.52 $Y2=1.202
r153 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.52 $Y=0.995
+ $X2=9.52 $Y2=0.56
r154 1 39 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.495 $Y=1.41
+ $X2=9.495 $Y2=1.202
r155 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.495 $Y=1.41
+ $X2=9.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_6%A_27_297# 1 2 3 4 5 6 7 22 24 26 30 32 36
+ 38 40 41 42 46 48 52 54 58 63 65 70 71
r88 56 58 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=5.94 $Y=2.295
+ $X2=5.94 $Y2=1.96
r89 55 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.105 $Y=2.38
+ $X2=4.98 $Y2=2.38
r90 54 56 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=5.795 $Y=2.38
+ $X2=5.94 $Y2=2.295
r91 54 55 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.795 $Y=2.38
+ $X2=5.105 $Y2=2.38
r92 50 71 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.295
+ $X2=4.98 $Y2=2.38
r93 50 52 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.98 $Y=2.295
+ $X2=4.98 $Y2=1.96
r94 49 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.165 $Y=2.38
+ $X2=4.04 $Y2=2.38
r95 48 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.855 $Y=2.38
+ $X2=4.98 $Y2=2.38
r96 48 49 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.855 $Y=2.38
+ $X2=4.165 $Y2=2.38
r97 44 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=2.295
+ $X2=4.04 $Y2=2.38
r98 44 46 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.04 $Y=2.295
+ $X2=4.04 $Y2=1.96
r99 43 69 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.225 $Y=2.38
+ $X2=3.1 $Y2=2.38
r100 42 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.915 $Y=2.38
+ $X2=4.04 $Y2=2.38
r101 42 43 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.915 $Y=2.38
+ $X2=3.225 $Y2=2.38
r102 41 69 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=2.295 $X2=3.1
+ $Y2=2.38
r103 40 67 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=1.625 $X2=3.1
+ $Y2=1.54
r104 40 41 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=3.1 $Y=1.625
+ $X2=3.1 $Y2=2.295
r105 39 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=1.54
+ $X2=2.16 $Y2=1.54
r106 38 67 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.975 $Y=1.54
+ $X2=3.1 $Y2=1.54
r107 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.975 $Y=1.54
+ $X2=2.285 $Y2=1.54
r108 34 65 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=1.625
+ $X2=2.16 $Y2=1.54
r109 34 36 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.16 $Y=1.625
+ $X2=2.16 $Y2=2.3
r110 33 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=1.54
+ $X2=1.22 $Y2=1.54
r111 32 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=1.54
+ $X2=2.16 $Y2=1.54
r112 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.035 $Y=1.54
+ $X2=1.345 $Y2=1.54
r113 28 63 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=1.625
+ $X2=1.22 $Y2=1.54
r114 28 30 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.22 $Y=1.625
+ $X2=1.22 $Y2=2.3
r115 27 61 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.405 $Y=1.54
+ $X2=0.26 $Y2=1.54
r116 26 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=1.54
+ $X2=1.22 $Y2=1.54
r117 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=1.54
+ $X2=0.405 $Y2=1.54
r118 22 61 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.26 $Y2=1.54
r119 22 24 26.8241 $w=2.88e-07 $l=6.75e-07 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.26 $Y2=2.3
r120 7 58 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.775
+ $Y=1.485 $X2=5.92 $Y2=1.96
r121 6 52 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.835
+ $Y=1.485 $X2=4.98 $Y2=1.96
r122 5 46 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.895
+ $Y=1.485 $X2=4.04 $Y2=1.96
r123 4 69 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.485 $X2=3.1 $Y2=2.3
r124 4 67 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.485 $X2=3.1 $Y2=1.62
r125 3 65 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=1.62
r126 3 36 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=2.3
r127 2 63 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.62
r128 2 30 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.3
r129 1 61 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r130 1 24 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_6%VPWR 1 2 3 14 16 20 22 26 28 35 36 39 42 45
+ 50
r138 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r139 43 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r140 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r141 40 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r142 40 50 0.125198 $w=4.8e-07 $l=4.4e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.25 $Y2=2.72
r143 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r144 35 36 0.885714 $w=1.7e-07 $l=1.785e-06 $layer=mcon $count=10 $X=12.19
+ $Y=2.72 $X2=12.19 $Y2=2.72
r145 33 36 2.61778 $w=4.8e-07 $l=9.2e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=12.19 $Y2=2.72
r146 33 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r147 32 35 600.214 $w=1.68e-07 $l=9.2e-06 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=12.19 $Y2=2.72
r148 32 33 0.885714 $w=1.7e-07 $l=1.785e-06 $layer=mcon $count=10 $X=2.99
+ $Y=2.72 $X2=2.99 $Y2=2.72
r149 30 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.755 $Y=2.72
+ $X2=2.63 $Y2=2.72
r150 30 32 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.755 $Y=2.72
+ $X2=2.99 $Y2=2.72
r151 28 50 0.00426813 $w=4.8e-07 $l=1.5e-08 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.25 $Y2=2.72
r152 24 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=2.635
+ $X2=2.63 $Y2=2.72
r153 24 26 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.63 $Y=2.635
+ $X2=2.63 $Y2=1.96
r154 23 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=1.69 $Y2=2.72
r155 22 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.505 $Y=2.72
+ $X2=2.63 $Y2=2.72
r156 22 23 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.505 $Y=2.72
+ $X2=1.815 $Y2=2.72
r157 18 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=2.635
+ $X2=1.69 $Y2=2.72
r158 18 20 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.69 $Y=2.635
+ $X2=1.69 $Y2=1.96
r159 17 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=0.75 $Y2=2.72
r160 16 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.565 $Y=2.72
+ $X2=1.69 $Y2=2.72
r161 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.565 $Y=2.72
+ $X2=0.875 $Y2=2.72
r162 12 39 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r163 12 14 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=1.96
r164 3 26 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.485
+ $Y=1.485 $X2=2.63 $Y2=1.96
r165 2 20 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=1.96
r166 1 14 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_6%A_685_297# 1 2 3 4 5 6 21 25 29 33 37 42 44
+ 46 48 50 52
r90 38 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.975 $Y=1.54
+ $X2=7.85 $Y2=1.54
r91 37 52 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.665 $Y=1.54
+ $X2=8.79 $Y2=1.54
r92 37 38 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.665 $Y=1.54
+ $X2=7.975 $Y2=1.54
r93 34 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.035 $Y=1.54
+ $X2=6.91 $Y2=1.54
r94 33 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.725 $Y=1.54
+ $X2=7.85 $Y2=1.54
r95 33 34 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.725 $Y=1.54
+ $X2=7.035 $Y2=1.54
r96 30 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.575 $Y=1.54
+ $X2=5.45 $Y2=1.54
r97 29 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.785 $Y=1.54
+ $X2=6.91 $Y2=1.54
r98 29 30 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=6.785 $Y=1.54
+ $X2=5.575 $Y2=1.54
r99 26 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.635 $Y=1.54
+ $X2=4.51 $Y2=1.54
r100 25 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.325 $Y=1.54
+ $X2=5.45 $Y2=1.54
r101 25 26 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.325 $Y=1.54
+ $X2=4.635 $Y2=1.54
r102 22 42 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.695 $Y=1.54
+ $X2=3.57 $Y2=1.54
r103 21 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.385 $Y=1.54
+ $X2=4.51 $Y2=1.54
r104 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.385 $Y=1.54
+ $X2=3.695 $Y2=1.54
r105 6 52 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=8.645
+ $Y=1.485 $X2=8.79 $Y2=1.62
r106 5 50 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=7.705
+ $Y=1.485 $X2=7.85 $Y2=1.62
r107 4 48 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.765
+ $Y=1.485 $X2=6.91 $Y2=1.62
r108 3 46 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=5.305
+ $Y=1.485 $X2=5.45 $Y2=1.62
r109 2 44 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=4.365
+ $Y=1.485 $X2=4.51 $Y2=1.62
r110 1 42 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.425
+ $Y=1.485 $X2=3.57 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_6%A_1263_297# 1 2 3 4 5 6 7 24 26 27 30 32 36
+ 38 42 44 48 50 54 56 58 60 62 63 65 66 67
r91 58 69 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.13 $Y=2.295
+ $X2=12.13 $Y2=2.38
r92 58 60 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=12.13 $Y=2.295
+ $X2=12.13 $Y2=1.62
r93 57 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.265 $Y=2.38
+ $X2=11.14 $Y2=2.38
r94 56 69 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.005 $Y=2.38
+ $X2=12.13 $Y2=2.38
r95 56 57 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=12.005 $Y=2.38
+ $X2=11.265 $Y2=2.38
r96 52 67 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.14 $Y=2.295
+ $X2=11.14 $Y2=2.38
r97 52 54 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=11.14 $Y=2.295
+ $X2=11.14 $Y2=1.96
r98 51 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.325 $Y=2.38
+ $X2=10.2 $Y2=2.38
r99 50 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.015 $Y=2.38
+ $X2=11.14 $Y2=2.38
r100 50 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.015 $Y=2.38
+ $X2=10.325 $Y2=2.38
r101 46 66 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.2 $Y=2.295
+ $X2=10.2 $Y2=2.38
r102 46 48 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=10.2 $Y=2.295
+ $X2=10.2 $Y2=1.96
r103 45 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.385 $Y=2.38
+ $X2=9.26 $Y2=2.38
r104 44 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.075 $Y=2.38
+ $X2=10.2 $Y2=2.38
r105 44 45 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.075 $Y=2.38
+ $X2=9.385 $Y2=2.38
r106 40 65 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.26 $Y=2.295
+ $X2=9.26 $Y2=2.38
r107 40 42 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=9.26 $Y=2.295
+ $X2=9.26 $Y2=1.62
r108 39 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.445 $Y=2.38
+ $X2=8.32 $Y2=2.38
r109 38 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.135 $Y=2.38
+ $X2=9.26 $Y2=2.38
r110 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.135 $Y=2.38
+ $X2=8.445 $Y2=2.38
r111 34 63 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.32 $Y=2.295
+ $X2=8.32 $Y2=2.38
r112 34 36 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=8.32 $Y=2.295
+ $X2=8.32 $Y2=1.96
r113 33 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.505 $Y=2.38
+ $X2=7.38 $Y2=2.38
r114 32 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.195 $Y=2.38
+ $X2=8.32 $Y2=2.38
r115 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.195 $Y=2.38
+ $X2=7.505 $Y2=2.38
r116 28 62 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.38 $Y=2.295
+ $X2=7.38 $Y2=2.38
r117 28 30 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=7.38 $Y=2.295
+ $X2=7.38 $Y2=1.96
r118 26 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.255 $Y=2.38
+ $X2=7.38 $Y2=2.38
r119 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.255 $Y=2.38
+ $X2=6.565 $Y2=2.38
r120 22 27 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=6.42 $Y=2.295
+ $X2=6.565 $Y2=2.38
r121 22 24 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=6.42 $Y=2.295
+ $X2=6.42 $Y2=1.96
r122 7 69 400 $w=1.7e-07 $l=8.89129e-07 $layer=licon1_PDIFF $count=1 $X=11.935
+ $Y=1.485 $X2=12.09 $Y2=2.3
r123 7 60 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=11.935
+ $Y=1.485 $X2=12.09 $Y2=1.62
r124 6 54 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=10.995
+ $Y=1.485 $X2=11.14 $Y2=1.96
r125 5 48 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=10.055
+ $Y=1.485 $X2=10.2 $Y2=1.96
r126 4 65 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=9.115
+ $Y=1.485 $X2=9.26 $Y2=2.3
r127 4 42 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.115
+ $Y=1.485 $X2=9.26 $Y2=1.62
r128 3 36 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=8.175
+ $Y=1.485 $X2=8.32 $Y2=1.96
r129 2 30 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=7.235
+ $Y=1.485 $X2=7.38 $Y2=1.96
r130 1 24 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=6.315
+ $Y=1.485 $X2=6.44 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_6%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 48 50
+ 51 54 56 60 62 66 68 72 74 78 80 84 86 90 92 96 98 102 106 108 112 116 118 122
+ 126 127 128 129 130 131 132 133 134 136 137 139 141 144 145
r307 142 145 7.8307 $w=3.88e-07 $l=2.65e-07 $layer=LI1_cond $X=11.64 $Y=1.455
+ $X2=11.64 $Y2=1.19
r308 142 144 2.47594 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=11.64 $Y=1.455
+ $X2=11.64 $Y2=1.54
r309 140 145 8.4217 $w=3.88e-07 $l=2.85e-07 $layer=LI1_cond $X=11.64 $Y=0.905
+ $X2=11.64 $Y2=1.19
r310 140 141 2.61037 $w=3.9e-07 $l=9e-08 $layer=LI1_cond $X=11.64 $Y=0.905
+ $X2=11.64 $Y2=0.815
r311 120 141 2.61037 $w=3.9e-07 $l=9e-08 $layer=LI1_cond $X=11.64 $Y=0.725
+ $X2=11.64 $Y2=0.815
r312 120 122 9.89919 $w=3.88e-07 $l=3.35e-07 $layer=LI1_cond $X=11.64 $Y=0.725
+ $X2=11.64 $Y2=0.39
r313 119 137 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=10.835 $Y=0.815
+ $X2=10.67 $Y2=0.815
r314 118 141 4.22815 $w=1.8e-07 $l=1.95e-07 $layer=LI1_cond $X=11.445 $Y=0.815
+ $X2=11.64 $Y2=0.815
r315 118 119 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=11.445 $Y=0.815
+ $X2=10.835 $Y2=0.815
r316 117 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.795 $Y=1.54
+ $X2=10.67 $Y2=1.54
r317 116 144 4.4465 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=11.445 $Y=1.54
+ $X2=11.64 $Y2=1.54
r318 116 117 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=11.445 $Y=1.54
+ $X2=10.795 $Y2=1.54
r319 110 137 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=10.67 $Y=0.725
+ $X2=10.67 $Y2=0.815
r320 110 112 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=10.67 $Y=0.725
+ $X2=10.67 $Y2=0.39
r321 109 134 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=9.895 $Y=0.815
+ $X2=9.73 $Y2=0.815
r322 108 137 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=10.505 $Y=0.815
+ $X2=10.67 $Y2=0.815
r323 108 109 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=10.505 $Y=0.815
+ $X2=9.895 $Y2=0.815
r324 107 136 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.855 $Y=1.54
+ $X2=9.73 $Y2=1.54
r325 106 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.545 $Y=1.54
+ $X2=10.67 $Y2=1.54
r326 106 107 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.545 $Y=1.54
+ $X2=9.855 $Y2=1.54
r327 100 134 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=9.73 $Y=0.725
+ $X2=9.73 $Y2=0.815
r328 100 102 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.73 $Y=0.725
+ $X2=9.73 $Y2=0.39
r329 99 133 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=8.955 $Y=0.815
+ $X2=8.79 $Y2=0.815
r330 98 134 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=9.565 $Y=0.815
+ $X2=9.73 $Y2=0.815
r331 98 99 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=9.565 $Y=0.815
+ $X2=8.955 $Y2=0.815
r332 94 133 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=8.79 $Y=0.725
+ $X2=8.79 $Y2=0.815
r333 94 96 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.79 $Y=0.725
+ $X2=8.79 $Y2=0.39
r334 93 132 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=8.015 $Y=0.815
+ $X2=7.85 $Y2=0.815
r335 92 133 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=8.625 $Y=0.815
+ $X2=8.79 $Y2=0.815
r336 92 93 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=8.625 $Y=0.815
+ $X2=8.015 $Y2=0.815
r337 88 132 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=7.85 $Y=0.725
+ $X2=7.85 $Y2=0.815
r338 88 90 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.85 $Y=0.725
+ $X2=7.85 $Y2=0.39
r339 87 131 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.075 $Y=0.815
+ $X2=6.91 $Y2=0.815
r340 86 132 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.685 $Y=0.815
+ $X2=7.85 $Y2=0.815
r341 86 87 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=7.685 $Y=0.815
+ $X2=7.075 $Y2=0.815
r342 82 131 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=6.91 $Y=0.725
+ $X2=6.91 $Y2=0.815
r343 82 84 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.91 $Y=0.725
+ $X2=6.91 $Y2=0.39
r344 81 130 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.615 $Y=0.815
+ $X2=5.45 $Y2=0.815
r345 80 131 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.745 $Y=0.815
+ $X2=6.91 $Y2=0.815
r346 80 81 69.6263 $w=1.78e-07 $l=1.13e-06 $layer=LI1_cond $X=6.745 $Y=0.815
+ $X2=5.615 $Y2=0.815
r347 76 130 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.45 $Y=0.725
+ $X2=5.45 $Y2=0.815
r348 76 78 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.45 $Y=0.725
+ $X2=5.45 $Y2=0.39
r349 75 129 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.675 $Y=0.815
+ $X2=4.51 $Y2=0.815
r350 74 130 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.285 $Y=0.815
+ $X2=5.45 $Y2=0.815
r351 74 75 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=5.285 $Y=0.815
+ $X2=4.675 $Y2=0.815
r352 70 129 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.51 $Y=0.725
+ $X2=4.51 $Y2=0.815
r353 70 72 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.51 $Y=0.725
+ $X2=4.51 $Y2=0.39
r354 69 128 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.735 $Y=0.815
+ $X2=3.57 $Y2=0.815
r355 68 129 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.345 $Y=0.815
+ $X2=4.51 $Y2=0.815
r356 68 69 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=4.345 $Y=0.815
+ $X2=3.735 $Y2=0.815
r357 64 128 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.57 $Y=0.725
+ $X2=3.57 $Y2=0.815
r358 64 66 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.57 $Y=0.725
+ $X2=3.57 $Y2=0.39
r359 63 127 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=0.815
+ $X2=2.63 $Y2=0.815
r360 62 128 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=0.815
+ $X2=3.57 $Y2=0.815
r361 62 63 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=3.405 $Y=0.815
+ $X2=2.795 $Y2=0.815
r362 58 127 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.63 $Y=0.725
+ $X2=2.63 $Y2=0.815
r363 58 60 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.63 $Y=0.725
+ $X2=2.63 $Y2=0.39
r364 57 126 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=0.815
+ $X2=1.69 $Y2=0.815
r365 56 127 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=0.815
+ $X2=2.63 $Y2=0.815
r366 56 57 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=2.465 $Y=0.815
+ $X2=1.855 $Y2=0.815
r367 52 126 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.69 $Y=0.725
+ $X2=1.69 $Y2=0.815
r368 52 54 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.69 $Y=0.725
+ $X2=1.69 $Y2=0.39
r369 50 126 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.525 $Y=0.815
+ $X2=1.69 $Y2=0.815
r370 50 51 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=1.525 $Y=0.815
+ $X2=0.915 $Y2=0.815
r371 46 51 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.75 $Y=0.725
+ $X2=0.915 $Y2=0.815
r372 46 48 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.75 $Y=0.725
+ $X2=0.75 $Y2=0.39
r373 15 144 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=11.465
+ $Y=1.485 $X2=11.61 $Y2=1.62
r374 14 139 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=10.525
+ $Y=1.485 $X2=10.67 $Y2=1.62
r375 13 136 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=9.585
+ $Y=1.485 $X2=9.73 $Y2=1.62
r376 12 122 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=11.475
+ $Y=0.235 $X2=11.61 $Y2=0.39
r377 11 112 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=10.535
+ $Y=0.235 $X2=10.67 $Y2=0.39
r378 10 102 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=9.595
+ $Y=0.235 $X2=9.73 $Y2=0.39
r379 9 96 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=8.655
+ $Y=0.235 $X2=8.79 $Y2=0.39
r380 8 90 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=7.715
+ $Y=0.235 $X2=7.85 $Y2=0.39
r381 7 84 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.775
+ $Y=0.235 $X2=6.91 $Y2=0.39
r382 6 78 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.315
+ $Y=0.235 $X2=5.45 $Y2=0.39
r383 5 72 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.375
+ $Y=0.235 $X2=4.51 $Y2=0.39
r384 4 66 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.435
+ $Y=0.235 $X2=3.57 $Y2=0.39
r385 3 60 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.495
+ $Y=0.235 $X2=2.63 $Y2=0.39
r386 2 54 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.555
+ $Y=0.235 $X2=1.69 $Y2=0.39
r387 1 48 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.615
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_6%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 40 42 44
+ 48 50 54 56 60 62 66 70 74 78 82 86 90 92 94 97 98 100 101 103 104 106 107 109
+ 110 112 113 114 140 148 151 154 157 162 165 168
r207 167 168 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r208 164 165 9.8562 $w=6.38e-07 $l=1.35e-07 $layer=LI1_cond $X=6.44 $Y=0.235
+ $X2=6.575 $Y2=0.235
r209 160 164 4.29841 $w=6.38e-07 $l=2.3e-07 $layer=LI1_cond $X=6.21 $Y=0.235
+ $X2=6.44 $Y2=0.235
r210 160 162 15.2759 $w=6.38e-07 $l=4.25e-07 $layer=LI1_cond $X=6.21 $Y=0.235
+ $X2=5.785 $Y2=0.235
r211 160 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r212 157 158 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r213 155 158 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.91 $Y2=0
r214 154 155 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r215 152 155 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=2.99 $Y2=0
r216 151 152 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r217 149 152 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.07 $Y2=0
r218 148 149 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r219 143 168 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.19 $Y2=0
r220 142 143 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r221 140 167 3.95357 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=12.005 $Y=0
+ $X2=12.212 $Y2=0
r222 140 142 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=12.005 $Y=0
+ $X2=11.73 $Y2=0
r223 139 143 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.73 $Y2=0
r224 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r225 136 139 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.81 $Y2=0
r226 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r227 133 136 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.89 $Y2=0
r228 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r229 130 133 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.97 $Y2=0
r230 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r231 127 130 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r232 127 161 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=6.21 $Y2=0
r233 126 165 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=7.13 $Y=0
+ $X2=6.575 $Y2=0
r234 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r235 123 161 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.21 $Y2=0
r236 122 162 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=5.75 $Y=0
+ $X2=5.785 $Y2=0
r237 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r238 119 123 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r239 119 158 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=3.91 $Y2=0
r240 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r241 116 157 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.175 $Y=0
+ $X2=4.04 $Y2=0
r242 116 118 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.175 $Y=0
+ $X2=4.83 $Y2=0
r243 114 149 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=1.15 $Y2=0
r244 114 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r245 112 138 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=11.005 $Y=0
+ $X2=10.81 $Y2=0
r246 112 113 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.005 $Y=0
+ $X2=11.14 $Y2=0
r247 111 142 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=11.275 $Y=0
+ $X2=11.73 $Y2=0
r248 111 113 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.275 $Y=0
+ $X2=11.14 $Y2=0
r249 109 135 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=10.065 $Y=0
+ $X2=9.89 $Y2=0
r250 109 110 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.065 $Y=0
+ $X2=10.2 $Y2=0
r251 108 138 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=10.335 $Y=0
+ $X2=10.81 $Y2=0
r252 108 110 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.335 $Y=0
+ $X2=10.2 $Y2=0
r253 106 132 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=9.125 $Y=0
+ $X2=8.97 $Y2=0
r254 106 107 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=9.125 $Y=0
+ $X2=9.26 $Y2=0
r255 105 135 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=9.395 $Y=0
+ $X2=9.89 $Y2=0
r256 105 107 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=9.395 $Y=0
+ $X2=9.26 $Y2=0
r257 103 129 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=8.185 $Y=0
+ $X2=8.05 $Y2=0
r258 103 104 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.185 $Y=0
+ $X2=8.32 $Y2=0
r259 102 132 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=8.455 $Y=0
+ $X2=8.97 $Y2=0
r260 102 104 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.455 $Y=0
+ $X2=8.32 $Y2=0
r261 100 126 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.245 $Y=0
+ $X2=7.13 $Y2=0
r262 100 101 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.245 $Y=0
+ $X2=7.38 $Y2=0
r263 99 129 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=7.515 $Y=0
+ $X2=8.05 $Y2=0
r264 99 101 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.515 $Y=0
+ $X2=7.38 $Y2=0
r265 97 118 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.845 $Y=0
+ $X2=4.83 $Y2=0
r266 97 98 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.845 $Y=0 $X2=4.98
+ $Y2=0
r267 96 122 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.115 $Y=0
+ $X2=5.75 $Y2=0
r268 96 98 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.115 $Y=0 $X2=4.98
+ $Y2=0
r269 92 167 3.18959 $w=2.5e-07 $l=1.19143e-07 $layer=LI1_cond $X=12.13 $Y=0.085
+ $X2=12.212 $Y2=0
r270 92 94 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=12.13 $Y=0.085
+ $X2=12.13 $Y2=0.39
r271 88 113 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.14 $Y=0.085
+ $X2=11.14 $Y2=0
r272 88 90 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=11.14 $Y=0.085
+ $X2=11.14 $Y2=0.39
r273 84 110 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.2 $Y=0.085
+ $X2=10.2 $Y2=0
r274 84 86 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.2 $Y=0.085
+ $X2=10.2 $Y2=0.39
r275 80 107 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.26 $Y=0.085
+ $X2=9.26 $Y2=0
r276 80 82 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.26 $Y=0.085
+ $X2=9.26 $Y2=0.39
r277 76 104 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.32 $Y=0.085
+ $X2=8.32 $Y2=0
r278 76 78 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.32 $Y=0.085
+ $X2=8.32 $Y2=0.39
r279 72 101 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.38 $Y=0.085
+ $X2=7.38 $Y2=0
r280 72 74 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.38 $Y=0.085
+ $X2=7.38 $Y2=0.39
r281 68 98 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0
r282 68 70 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0.39
r283 64 157 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0
r284 64 66 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0.39
r285 63 154 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.235 $Y=0 $X2=3.1
+ $Y2=0
r286 62 157 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.905 $Y=0
+ $X2=4.04 $Y2=0
r287 62 63 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.905 $Y=0
+ $X2=3.235 $Y2=0
r288 58 154 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=0.085
+ $X2=3.1 $Y2=0
r289 58 60 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.1 $Y=0.085
+ $X2=3.1 $Y2=0.39
r290 57 151 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.295 $Y=0
+ $X2=2.16 $Y2=0
r291 56 154 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.965 $Y=0 $X2=3.1
+ $Y2=0
r292 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.965 $Y=0
+ $X2=2.295 $Y2=0
r293 52 151 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0
r294 52 54 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0.39
r295 51 148 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.355 $Y=0
+ $X2=1.22 $Y2=0
r296 50 151 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=2.16 $Y2=0
r297 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=1.355 $Y2=0
r298 46 148 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r299 46 48 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.39
r300 45 145 4.45492 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.415 $Y=0
+ $X2=0.207 $Y2=0
r301 44 148 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.085 $Y=0
+ $X2=1.22 $Y2=0
r302 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.085 $Y=0
+ $X2=0.415 $Y2=0
r303 40 145 3.06275 $w=3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.207 $Y2=0
r304 40 42 11.7165 $w=2.98e-07 $l=3.05e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.265 $Y2=0.39
r305 13 94 91 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_NDIFF $count=2 $X=11.895
+ $Y=0.235 $X2=12.09 $Y2=0.39
r306 12 90 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=10.955
+ $Y=0.235 $X2=11.14 $Y2=0.39
r307 11 86 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=10.015
+ $Y=0.235 $X2=10.2 $Y2=0.39
r308 10 82 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=9.075
+ $Y=0.235 $X2=9.26 $Y2=0.39
r309 9 78 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=8.135
+ $Y=0.235 $X2=8.32 $Y2=0.39
r310 8 74 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=7.195
+ $Y=0.235 $X2=7.38 $Y2=0.39
r311 7 164 91 $w=1.7e-07 $l=7.78653e-07 $layer=licon1_NDIFF $count=2 $X=5.735
+ $Y=0.235 $X2=6.44 $Y2=0.39
r312 6 70 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.795
+ $Y=0.235 $X2=4.98 $Y2=0.39
r313 5 66 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=3.855
+ $Y=0.235 $X2=4.04 $Y2=0.39
r314 4 60 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.235 $X2=3.1 $Y2=0.39
r315 3 54 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.16 $Y2=0.39
r316 2 48 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.235 $X2=1.22 $Y2=0.39
r317 1 42 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

