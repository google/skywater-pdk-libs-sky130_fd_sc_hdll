* NGSPICE file created from sky130_fd_sc_hdll__xor3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__xor3_1 A B C VGND VNB VPB VPWR X
M1000 VGND A a_991_365# VNB nshort w=640000u l=150000u
+  ad=9.7095e+11p pd=6.94e+06u as=4.498e+11p ps=3.99e+06u
M1001 a_276_93# C VPWR VPB phighvt w=640000u l=180000u
+  ad=1.856e+11p pd=1.86e+06u as=1.3094e+12p ps=8.68e+06u
M1002 a_276_93# C VGND VNB nshort w=420000u l=150000u
+  ad=1.974e+11p pd=1.78e+06u as=0p ps=0u
M1003 a_875_297# B VGND VNB nshort w=650000u l=150000u
+  ad=1.653e+11p pd=1.82e+06u as=0p ps=0u
M1004 a_424_49# B a_991_365# VNB nshort w=640000u l=150000u
+  ad=5.931e+11p pd=4.52e+06u as=0p ps=0u
M1005 a_116_21# C a_406_325# VPB phighvt w=840000u l=180000u
+  ad=3.36e+11p pd=2.48e+06u as=7.824e+11p ps=5.28e+06u
M1006 a_875_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.126e+11p pd=2.64e+06u as=0p ps=0u
M1007 a_116_21# C a_424_49# VNB nshort w=640000u l=150000u
+  ad=2.88e+11p pd=2.18e+06u as=0p ps=0u
M1008 a_1276_297# a_875_297# a_424_49# VNB nshort w=420000u l=150000u
+  ad=5.677e+11p pd=4.42e+06u as=0p ps=0u
M1009 a_406_325# B a_1276_297# VNB nshort w=640000u l=150000u
+  ad=6.5745e+11p pd=4.66e+06u as=0p ps=0u
M1010 a_991_365# a_875_297# a_424_49# VPB phighvt w=840000u l=180000u
+  ad=7.234e+11p pd=5.3e+06u as=7.558e+11p ps=5.2e+06u
M1011 a_406_325# B a_991_365# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_424_49# B a_1276_297# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=7.998e+11p ps=5.68e+06u
M1013 a_1276_297# a_991_365# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_991_365# a_875_297# a_406_325# VNB nshort w=600000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1276_297# a_875_297# a_406_325# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A a_991_365# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_424_49# a_276_93# a_116_21# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_116_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.82e+11p ps=1.86e+06u
M1019 VPWR a_116_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1020 a_406_325# a_276_93# a_116_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1276_297# a_991_365# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

