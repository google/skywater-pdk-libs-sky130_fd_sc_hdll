* File: sky130_fd_sc_hdll__a22oi_2.pxi.spice
* Created: Thu Aug 27 18:54:29 2020
* 
x_PM_SKY130_FD_SC_HDLL__A22OI_2%B2 N_B2_c_70_n N_B2_M1000_g N_B2_c_66_n
+ N_B2_M1001_g N_B2_c_71_n N_B2_M1008_g N_B2_c_67_n N_B2_M1011_g B2 B2
+ N_B2_c_68_n B2 PM_SKY130_FD_SC_HDLL__A22OI_2%B2
x_PM_SKY130_FD_SC_HDLL__A22OI_2%B1 N_B1_c_108_n N_B1_M1004_g N_B1_c_112_n
+ N_B1_M1009_g N_B1_c_113_n N_B1_M1014_g N_B1_c_109_n N_B1_M1012_g B1 B1
+ N_B1_c_110_n B1 B1 PM_SKY130_FD_SC_HDLL__A22OI_2%B1
x_PM_SKY130_FD_SC_HDLL__A22OI_2%A1 N_A1_c_163_n N_A1_M1003_g N_A1_c_159_n
+ N_A1_M1002_g N_A1_c_164_n N_A1_M1006_g N_A1_c_160_n N_A1_M1007_g A1 A1
+ N_A1_c_161_n A1 A1 PM_SKY130_FD_SC_HDLL__A22OI_2%A1
x_PM_SKY130_FD_SC_HDLL__A22OI_2%A2 N_A2_c_211_n N_A2_M1005_g N_A2_c_215_n
+ N_A2_M1010_g N_A2_c_216_n N_A2_M1015_g N_A2_c_212_n N_A2_M1013_g A2 A2
+ N_A2_c_214_n A2 PM_SKY130_FD_SC_HDLL__A22OI_2%A2
x_PM_SKY130_FD_SC_HDLL__A22OI_2%Y N_Y_M1004_d N_Y_M1002_s N_Y_M1000_d
+ N_Y_M1008_d N_Y_M1014_d N_Y_c_254_n N_Y_c_261_n N_Y_c_255_n N_Y_c_267_n
+ N_Y_c_272_n N_Y_c_276_n N_Y_c_251_n N_Y_c_256_n Y Y Y Y Y N_Y_c_259_n
+ PM_SKY130_FD_SC_HDLL__A22OI_2%Y
x_PM_SKY130_FD_SC_HDLL__A22OI_2%A_117_297# N_A_117_297#_M1000_s
+ N_A_117_297#_M1009_s N_A_117_297#_M1003_d N_A_117_297#_M1006_d
+ N_A_117_297#_M1015_d N_A_117_297#_c_344_n N_A_117_297#_c_345_n
+ N_A_117_297#_c_346_n N_A_117_297#_c_384_n N_A_117_297#_c_339_n
+ N_A_117_297#_c_350_n N_A_117_297#_c_349_n N_A_117_297#_c_353_n
+ N_A_117_297#_c_340_n N_A_117_297#_c_360_n N_A_117_297#_c_341_n
+ N_A_117_297#_c_342_n N_A_117_297#_c_406_p N_A_117_297#_c_343_n
+ PM_SKY130_FD_SC_HDLL__A22OI_2%A_117_297#
x_PM_SKY130_FD_SC_HDLL__A22OI_2%VPWR N_VPWR_M1003_s N_VPWR_M1010_s
+ N_VPWR_c_424_n N_VPWR_c_425_n N_VPWR_c_426_n N_VPWR_c_427_n N_VPWR_c_428_n
+ N_VPWR_c_429_n VPWR VPWR VPWR N_VPWR_c_430_n N_VPWR_c_423_n
+ PM_SKY130_FD_SC_HDLL__A22OI_2%VPWR
x_PM_SKY130_FD_SC_HDLL__A22OI_2%A_27_47# N_A_27_47#_M1001_d N_A_27_47#_M1011_d
+ N_A_27_47#_M1012_s N_A_27_47#_c_485_n N_A_27_47#_c_489_n N_A_27_47#_c_486_n
+ N_A_27_47#_c_508_p N_A_27_47#_c_487_n PM_SKY130_FD_SC_HDLL__A22OI_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__A22OI_2%VGND N_VGND_M1001_s N_VGND_M1005_s
+ N_VGND_c_522_n N_VGND_c_523_n N_VGND_c_524_n VGND VGND N_VGND_c_526_n
+ N_VGND_c_527_n N_VGND_c_528_n N_VGND_c_529_n
+ PM_SKY130_FD_SC_HDLL__A22OI_2%VGND
x_PM_SKY130_FD_SC_HDLL__A22OI_2%A_507_47# N_A_507_47#_M1002_d
+ N_A_507_47#_M1007_d N_A_507_47#_M1013_d N_A_507_47#_c_584_n
+ N_A_507_47#_c_590_n N_A_507_47#_c_585_n N_A_507_47#_c_591_n
+ N_A_507_47#_c_586_n PM_SKY130_FD_SC_HDLL__A22OI_2%A_507_47#
cc_1 VNB N_B2_c_66_n 0.0219558f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB N_B2_c_67_n 0.0167331f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB N_B2_c_68_n 0.0500592f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_4 VNB B2 0.0105733f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_5 VNB N_B1_c_108_n 0.0171642f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_6 VNB N_B1_c_109_n 0.0208617f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_7 VNB N_B1_c_110_n 0.0385596f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_8 VNB B1 0.00568899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A1_c_159_n 0.0203777f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_10 VNB N_A1_c_160_n 0.0176098f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_11 VNB N_A1_c_161_n 0.0475229f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_12 VNB A1 0.00568036f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A2_c_211_n 0.017839f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_14 VNB N_A2_c_212_n 0.0226943f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_15 VNB A2 0.0131271f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_16 VNB N_A2_c_214_n 0.0442787f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_17 VNB N_Y_c_251_n 0.0092054f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB Y 0.00170628f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB Y 0.00786012f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_423_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_485_n 0.0161681f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_22 VNB N_A_27_47#_c_486_n 0.00783052f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_23 VNB N_A_27_47#_c_487_n 0.00293729f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_24 VNB N_VGND_c_522_n 5.44809e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_25 VNB N_VGND_c_523_n 0.0707198f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_26 VNB N_VGND_c_524_n 0.00508852f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_27 VNB VGND 0.00573949f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_28 VNB N_VGND_c_526_n 0.0144524f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_29 VNB N_VGND_c_527_n 0.0195794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_528_n 0.265131f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_529_n 0.00280658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_507_47#_c_584_n 0.00289221f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_33 VNB N_A_507_47#_c_585_n 0.0110523f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_34 VNB N_A_507_47#_c_586_n 0.0182437f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_35 VPB N_B2_c_70_n 0.0210029f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_36 VPB N_B2_c_71_n 0.0163884f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_37 VPB N_B2_c_68_n 0.0260351f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_38 VPB N_B1_c_112_n 0.0163826f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_39 VPB N_B1_c_113_n 0.0195908f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_40 VPB N_B1_c_110_n 0.0205108f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_41 VPB N_A1_c_163_n 0.0195195f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_42 VPB N_A1_c_164_n 0.0171107f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_43 VPB N_A1_c_161_n 0.0241803f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_44 VPB N_A2_c_215_n 0.0171107f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_45 VPB N_A2_c_216_n 0.0210029f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_46 VPB N_A2_c_214_n 0.0231908f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_47 VPB N_Y_c_254_n 0.0305923f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_48 VPB N_Y_c_255_n 0.00982506f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_49 VPB N_Y_c_256_n 0.00171921f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB Y 0.00190162f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB Y 0.00355713f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_Y_c_259_n 0.00599414f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_117_297#_c_339_n 0.0105087f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_117_297#_c_340_n 0.00196636f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_117_297#_c_341_n 0.0109515f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_117_297#_c_342_n 0.0321265f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_117_297#_c_343_n 0.00625553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_424_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_59 VPB N_VPWR_c_425_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_60 VPB N_VPWR_c_426_n 0.0743192f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_427_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.202
cc_62 VPB N_VPWR_c_428_n 0.0228593f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_63 VPB N_VPWR_c_429_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_64 VPB N_VPWR_c_430_n 0.0240648f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_423_n 0.0536741f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 N_B2_c_67_n N_B1_c_108_n 0.0234135f $X=0.99 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_67 N_B2_c_71_n N_B1_c_112_n 0.0225713f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_68 N_B2_c_68_n N_B1_c_110_n 0.0234135f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_69 N_B2_c_68_n B1 0.00711339f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_70 B2 B1 0.014751f $X=0.695 $Y=1.19 $X2=0 $Y2=0
cc_71 N_B2_c_70_n N_Y_c_254_n 0.00606201f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_72 N_B2_c_70_n N_Y_c_261_n 0.0158832f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_73 N_B2_c_71_n N_Y_c_261_n 0.00993063f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_74 N_B2_c_68_n N_Y_c_261_n 0.0065164f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_75 B2 N_Y_c_261_n 0.0248494f $X=0.695 $Y=1.19 $X2=0 $Y2=0
cc_76 N_B2_c_68_n N_Y_c_255_n 0.00169719f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_77 B2 N_Y_c_255_n 0.0137141f $X=0.695 $Y=1.19 $X2=0 $Y2=0
cc_78 N_B2_c_70_n N_Y_c_267_n 5.07942e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_79 N_B2_c_71_n N_Y_c_267_n 0.00905045f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_80 N_B2_c_71_n N_Y_c_256_n 0.00280691f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_81 N_B2_c_70_n N_A_117_297#_c_344_n 0.00778357f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_82 N_B2_c_71_n N_A_117_297#_c_345_n 0.0104149f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_83 N_B2_c_70_n N_A_117_297#_c_346_n 0.00305463f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_84 N_B2_c_70_n N_VPWR_c_426_n 0.00596194f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_85 N_B2_c_71_n N_VPWR_c_426_n 0.00429453f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_86 N_B2_c_70_n N_VPWR_c_423_n 0.0110796f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_87 N_B2_c_71_n N_VPWR_c_423_n 0.00609118f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_88 N_B2_c_66_n N_A_27_47#_c_485_n 0.00634847f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_89 N_B2_c_66_n N_A_27_47#_c_489_n 0.0114189f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_90 N_B2_c_67_n N_A_27_47#_c_489_n 0.0127252f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_91 N_B2_c_68_n N_A_27_47#_c_489_n 0.00570291f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_92 B2 N_A_27_47#_c_489_n 0.0240276f $X=0.695 $Y=1.19 $X2=0 $Y2=0
cc_93 N_B2_c_68_n N_A_27_47#_c_486_n 0.0017342f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_94 B2 N_A_27_47#_c_486_n 0.012897f $X=0.695 $Y=1.19 $X2=0 $Y2=0
cc_95 N_B2_c_67_n N_VGND_c_523_n 0.00431606f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_96 N_B2_c_66_n N_VGND_c_526_n 0.00200664f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_97 N_B2_c_66_n N_VGND_c_528_n 0.00372264f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_98 N_B2_c_67_n N_VGND_c_528_n 0.0059003f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_99 N_B2_c_66_n N_VGND_c_529_n 0.011864f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_100 N_B2_c_67_n N_VGND_c_529_n 0.00317372f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_101 N_B1_c_110_n N_A1_c_161_n 0.00371462f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_102 N_B1_c_110_n A1 5.28075e-19 $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_103 N_B1_c_112_n N_Y_c_267_n 0.0068728f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_104 N_B1_c_113_n N_Y_c_267_n 5.41141e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_105 N_B1_c_112_n N_Y_c_272_n 0.0115007f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_106 N_B1_c_113_n N_Y_c_272_n 0.00988775f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_107 N_B1_c_110_n N_Y_c_272_n 0.00637297f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_108 B1 N_Y_c_272_n 0.0207635f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_109 N_B1_c_108_n N_Y_c_276_n 0.00257667f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_110 N_B1_c_109_n N_Y_c_276_n 0.00405728f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_111 N_B1_c_110_n N_Y_c_276_n 0.0045813f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_112 B1 N_Y_c_276_n 0.014583f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_113 N_B1_c_112_n N_Y_c_256_n 5.95141e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_114 B1 N_Y_c_256_n 0.0191343f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_115 N_B1_c_109_n Y 0.00637354f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_116 N_B1_c_113_n Y 0.00124298f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_117 N_B1_c_108_n Y 6.45771e-19 $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_118 N_B1_c_112_n Y 3.6902e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_119 N_B1_c_113_n Y 0.00318468f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_120 N_B1_c_109_n Y 0.00656444f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B1_c_110_n Y 0.0216169f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_122 B1 Y 0.0151116f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_123 N_B1_c_112_n N_Y_c_259_n 5.76782e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_124 N_B1_c_113_n N_Y_c_259_n 0.00884964f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_125 N_B1_c_112_n N_A_117_297#_c_345_n 0.0111434f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_126 N_B1_c_113_n N_A_117_297#_c_339_n 0.0124578f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_127 N_B1_c_113_n N_A_117_297#_c_349_n 0.00324063f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_128 N_B1_c_112_n N_VPWR_c_426_n 0.00429453f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_129 N_B1_c_113_n N_VPWR_c_426_n 0.00429453f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_130 N_B1_c_112_n N_VPWR_c_423_n 0.00609118f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_131 N_B1_c_113_n N_VPWR_c_423_n 0.00739666f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_132 B1 N_A_27_47#_c_489_n 0.0144906f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_133 N_B1_c_108_n N_A_27_47#_c_487_n 0.0131478f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_134 N_B1_c_109_n N_A_27_47#_c_487_n 0.0105232f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_135 B1 N_A_27_47#_c_487_n 0.00395343f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_136 N_B1_c_108_n N_VGND_c_523_n 0.00357877f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_137 N_B1_c_109_n N_VGND_c_523_n 0.00357877f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_138 N_B1_c_108_n N_VGND_c_528_n 0.00554393f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_139 N_B1_c_109_n N_VGND_c_528_n 0.00680287f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A1_c_160_n N_A2_c_211_n 0.0190866f $X=3.39 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_141 N_A1_c_164_n N_A2_c_215_n 0.0217731f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A1_c_161_n A2 7.73302e-19 $X=3.365 $Y=1.202 $X2=0 $Y2=0
cc_143 A1 A2 0.0147576f $X=3.415 $Y=1.19 $X2=0 $Y2=0
cc_144 N_A1_c_161_n N_A2_c_214_n 0.0190866f $X=3.365 $Y=1.202 $X2=0 $Y2=0
cc_145 A1 N_A2_c_214_n 7.8169e-19 $X=3.415 $Y=1.19 $X2=0 $Y2=0
cc_146 N_A1_c_159_n N_Y_c_251_n 0.0108195f $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A1_c_161_n N_Y_c_251_n 0.00734086f $X=3.365 $Y=1.202 $X2=0 $Y2=0
cc_148 A1 N_Y_c_251_n 0.0319615f $X=3.415 $Y=1.19 $X2=0 $Y2=0
cc_149 N_A1_c_163_n Y 0.00215082f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A1_c_159_n Y 0.0041059f $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A1_c_161_n Y 0.00686246f $X=3.365 $Y=1.202 $X2=0 $Y2=0
cc_152 A1 Y 0.012447f $X=3.415 $Y=1.19 $X2=0 $Y2=0
cc_153 N_A1_c_163_n N_A_117_297#_c_350_n 0.00215639f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_154 N_A1_c_163_n N_A_117_297#_c_349_n 0.00859039f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_155 N_A1_c_164_n N_A_117_297#_c_349_n 5.97821e-19 $X=3.365 $Y=1.41 $X2=0
+ $Y2=0
cc_156 N_A1_c_163_n N_A_117_297#_c_353_n 0.0140468f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A1_c_164_n N_A_117_297#_c_353_n 0.0102366f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A1_c_161_n N_A_117_297#_c_353_n 0.0065164f $X=3.365 $Y=1.202 $X2=0
+ $Y2=0
cc_159 A1 N_A_117_297#_c_353_n 0.0295688f $X=3.415 $Y=1.19 $X2=0 $Y2=0
cc_160 N_A1_c_163_n N_A_117_297#_c_340_n 6.12117e-19 $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_161 N_A1_c_161_n N_A_117_297#_c_340_n 0.00273196f $X=3.365 $Y=1.202 $X2=0
+ $Y2=0
cc_162 A1 N_A_117_297#_c_340_n 0.0100453f $X=3.415 $Y=1.19 $X2=0 $Y2=0
cc_163 N_A1_c_163_n N_A_117_297#_c_360_n 6.72814e-19 $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_164 N_A1_c_164_n N_A_117_297#_c_360_n 0.0254977f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A1_c_164_n N_A_117_297#_c_343_n 0.00481936f $X=3.365 $Y=1.41 $X2=0
+ $Y2=0
cc_166 A1 N_A_117_297#_c_343_n 0.0080638f $X=3.415 $Y=1.19 $X2=0 $Y2=0
cc_167 N_A1_c_163_n N_VPWR_c_424_n 0.00523952f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A1_c_164_n N_VPWR_c_424_n 0.00477849f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A1_c_163_n N_VPWR_c_426_n 0.00672099f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A1_c_164_n N_VPWR_c_428_n 0.00597712f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A1_c_163_n N_VPWR_c_423_n 0.0130892f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A1_c_164_n N_VPWR_c_423_n 0.0102887f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A1_c_160_n N_VGND_c_522_n 0.00114049f $X=3.39 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A1_c_159_n N_VGND_c_523_n 0.00357877f $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A1_c_160_n N_VGND_c_523_n 0.00357877f $X=3.39 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A1_c_159_n N_VGND_c_528_n 0.00668309f $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A1_c_160_n N_VGND_c_528_n 0.00565902f $X=3.39 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A1_c_159_n N_A_507_47#_c_584_n 0.0101441f $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A1_c_160_n N_A_507_47#_c_584_n 0.0152957f $X=3.39 $Y=0.995 $X2=0 $Y2=0
cc_180 A1 N_A_507_47#_c_584_n 0.00554306f $X=3.415 $Y=1.19 $X2=0 $Y2=0
cc_181 N_A1_c_160_n N_A_507_47#_c_590_n 0.00384138f $X=3.39 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A1_c_160_n N_A_507_47#_c_591_n 0.00182231f $X=3.39 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A2_c_215_n N_A_117_297#_c_360_n 0.0107419f $X=3.935 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A2_c_216_n N_A_117_297#_c_360_n 6.47444e-19 $X=4.405 $Y=1.41 $X2=0
+ $Y2=0
cc_185 N_A2_c_215_n N_A_117_297#_c_341_n 0.0140468f $X=3.935 $Y=1.41 $X2=0 $Y2=0
cc_186 N_A2_c_216_n N_A_117_297#_c_341_n 0.0125026f $X=4.405 $Y=1.41 $X2=0 $Y2=0
cc_187 A2 N_A_117_297#_c_341_n 0.0408255f $X=4.3 $Y=1.105 $X2=0 $Y2=0
cc_188 N_A2_c_214_n N_A_117_297#_c_341_n 0.00631727f $X=4.405 $Y=1.202 $X2=0
+ $Y2=0
cc_189 N_A2_c_215_n N_A_117_297#_c_342_n 6.74705e-19 $X=3.935 $Y=1.41 $X2=0
+ $Y2=0
cc_190 N_A2_c_216_n N_A_117_297#_c_342_n 0.0132104f $X=4.405 $Y=1.41 $X2=0 $Y2=0
cc_191 N_A2_c_215_n N_A_117_297#_c_343_n 6.12117e-19 $X=3.935 $Y=1.41 $X2=0
+ $Y2=0
cc_192 A2 N_A_117_297#_c_343_n 0.00441973f $X=4.3 $Y=1.105 $X2=0 $Y2=0
cc_193 N_A2_c_215_n N_VPWR_c_425_n 0.00524193f $X=3.935 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A2_c_216_n N_VPWR_c_425_n 0.00477849f $X=4.405 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A2_c_215_n N_VPWR_c_428_n 0.00673617f $X=3.935 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A2_c_216_n N_VPWR_c_430_n 0.00597712f $X=4.405 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A2_c_215_n N_VPWR_c_423_n 0.0120877f $X=3.935 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A2_c_216_n N_VPWR_c_423_n 0.0110244f $X=4.405 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A2_c_211_n N_VGND_c_522_n 0.00728397f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A2_c_212_n N_VGND_c_522_n 0.00778384f $X=4.43 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A2_c_211_n N_VGND_c_523_n 0.00416467f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A2_c_212_n N_VGND_c_527_n 0.00416467f $X=4.43 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A2_c_211_n N_VGND_c_528_n 0.00507032f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A2_c_212_n N_VGND_c_528_n 0.00592483f $X=4.43 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A2_c_211_n N_A_507_47#_c_585_n 0.0115761f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A2_c_212_n N_A_507_47#_c_585_n 0.0124346f $X=4.43 $Y=0.995 $X2=0 $Y2=0
cc_207 A2 N_A_507_47#_c_585_n 0.0416051f $X=4.3 $Y=1.105 $X2=0 $Y2=0
cc_208 N_A2_c_214_n N_A_507_47#_c_585_n 0.00451459f $X=4.405 $Y=1.202 $X2=0
+ $Y2=0
cc_209 A2 N_A_507_47#_c_591_n 7.63207e-19 $X=4.3 $Y=1.105 $X2=0 $Y2=0
cc_210 N_Y_c_261_n N_A_117_297#_M1000_s 0.00342165f $X=0.985 $Y=1.57 $X2=-0.19
+ $Y2=-0.24
cc_211 N_Y_c_272_n N_A_117_297#_M1009_s 0.00343916f $X=1.925 $Y=1.57 $X2=0 $Y2=0
cc_212 N_Y_c_254_n N_A_117_297#_c_344_n 0.0354254f $X=0.26 $Y=1.8 $X2=0 $Y2=0
cc_213 N_Y_c_261_n N_A_117_297#_c_344_n 0.0191122f $X=0.985 $Y=1.57 $X2=0 $Y2=0
cc_214 N_Y_c_267_n N_A_117_297#_c_344_n 0.0233631f $X=1.2 $Y=1.66 $X2=0 $Y2=0
cc_215 N_Y_M1008_d N_A_117_297#_c_345_n 0.00352392f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_216 N_Y_c_261_n N_A_117_297#_c_345_n 0.00249206f $X=0.985 $Y=1.57 $X2=0 $Y2=0
cc_217 N_Y_c_267_n N_A_117_297#_c_345_n 0.0195208f $X=1.2 $Y=1.66 $X2=0 $Y2=0
cc_218 N_Y_c_272_n N_A_117_297#_c_345_n 0.00361673f $X=1.925 $Y=1.57 $X2=0 $Y2=0
cc_219 N_Y_c_254_n N_A_117_297#_c_346_n 0.0137304f $X=0.26 $Y=1.8 $X2=0 $Y2=0
cc_220 N_Y_c_267_n N_A_117_297#_c_384_n 0.0183625f $X=1.2 $Y=1.66 $X2=0 $Y2=0
cc_221 N_Y_c_272_n N_A_117_297#_c_384_n 0.0136007f $X=1.925 $Y=1.57 $X2=0 $Y2=0
cc_222 N_Y_c_259_n N_A_117_297#_c_384_n 0.0226368f $X=2.14 $Y=1.66 $X2=0 $Y2=0
cc_223 N_Y_M1014_d N_A_117_297#_c_339_n 0.00510164f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_224 N_Y_c_272_n N_A_117_297#_c_339_n 0.00249206f $X=1.925 $Y=1.57 $X2=0 $Y2=0
cc_225 N_Y_c_259_n N_A_117_297#_c_339_n 0.0285489f $X=2.14 $Y=1.66 $X2=0 $Y2=0
cc_226 N_Y_c_259_n N_A_117_297#_c_349_n 0.03244f $X=2.14 $Y=1.66 $X2=0 $Y2=0
cc_227 N_Y_c_251_n N_A_117_297#_c_340_n 0.00209868f $X=3.13 $Y=0.76 $X2=0 $Y2=0
cc_228 Y N_A_117_297#_c_340_n 0.0131731f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_229 N_Y_c_254_n N_VPWR_c_426_n 0.0174931f $X=0.26 $Y=1.8 $X2=0 $Y2=0
cc_230 N_Y_M1000_d N_VPWR_c_423_n 0.00430086f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_231 N_Y_M1008_d N_VPWR_c_423_n 0.00232895f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_232 N_Y_M1014_d N_VPWR_c_423_n 0.00218346f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_233 N_Y_c_254_n N_VPWR_c_423_n 0.00955092f $X=0.26 $Y=1.8 $X2=0 $Y2=0
cc_234 Y N_A_27_47#_M1012_s 0.00293402f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_235 N_Y_c_261_n N_A_27_47#_c_489_n 0.00240635f $X=0.985 $Y=1.57 $X2=0 $Y2=0
cc_236 N_Y_c_256_n N_A_27_47#_c_489_n 0.00113658f $X=1.175 $Y=1.57 $X2=0 $Y2=0
cc_237 N_Y_c_255_n N_A_27_47#_c_486_n 0.00196792f $X=0.345 $Y=1.57 $X2=0 $Y2=0
cc_238 N_Y_M1004_d N_A_27_47#_c_487_n 0.00509721f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_239 N_Y_c_276_n N_A_27_47#_c_487_n 0.0252434f $X=1.93 $Y=0.76 $X2=0 $Y2=0
cc_240 Y N_A_27_47#_c_487_n 0.0250128f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_241 N_Y_c_251_n N_VGND_c_523_n 0.00226279f $X=3.13 $Y=0.76 $X2=0 $Y2=0
cc_242 Y N_VGND_c_523_n 0.00103015f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_243 N_Y_M1004_d N_VGND_c_528_n 0.00297142f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_244 N_Y_M1002_s N_VGND_c_528_n 0.00256987f $X=2.995 $Y=0.235 $X2=0 $Y2=0
cc_245 N_Y_c_251_n N_VGND_c_528_n 0.00510281f $X=3.13 $Y=0.76 $X2=0 $Y2=0
cc_246 Y N_VGND_c_528_n 0.00246963f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_247 N_Y_c_251_n N_A_507_47#_M1002_d 0.00821042f $X=3.13 $Y=0.76 $X2=-0.19
+ $Y2=-0.24
cc_248 N_Y_M1002_s N_A_507_47#_c_584_n 0.00400706f $X=2.995 $Y=0.235 $X2=0 $Y2=0
cc_249 N_Y_c_251_n N_A_507_47#_c_584_n 0.0457715f $X=3.13 $Y=0.76 $X2=0 $Y2=0
cc_250 N_A_117_297#_c_353_n N_VPWR_M1003_s 0.00337913f $X=3.385 $Y=1.57
+ $X2=-0.19 $Y2=1.305
cc_251 N_A_117_297#_c_341_n N_VPWR_M1010_s 0.00337913f $X=4.425 $Y=1.57 $X2=0
+ $Y2=0
cc_252 N_A_117_297#_c_350_n N_VPWR_c_424_n 0.0109394f $X=2.7 $Y=2.295 $X2=0
+ $Y2=0
cc_253 N_A_117_297#_c_349_n N_VPWR_c_424_n 0.0278277f $X=2.66 $Y=1.66 $X2=0
+ $Y2=0
cc_254 N_A_117_297#_c_353_n N_VPWR_c_424_n 0.0136682f $X=3.385 $Y=1.57 $X2=0
+ $Y2=0
cc_255 N_A_117_297#_c_360_n N_VPWR_c_424_n 0.0486716f $X=3.7 $Y=1.66 $X2=0 $Y2=0
cc_256 N_A_117_297#_c_360_n N_VPWR_c_425_n 0.0398994f $X=3.7 $Y=1.66 $X2=0 $Y2=0
cc_257 N_A_117_297#_c_341_n N_VPWR_c_425_n 0.0136682f $X=4.425 $Y=1.57 $X2=0
+ $Y2=0
cc_258 N_A_117_297#_c_342_n N_VPWR_c_425_n 0.0477793f $X=4.64 $Y=1.66 $X2=0
+ $Y2=0
cc_259 N_A_117_297#_c_345_n N_VPWR_c_426_n 0.0415032f $X=1.585 $Y=2.38 $X2=0
+ $Y2=0
cc_260 N_A_117_297#_c_346_n N_VPWR_c_426_n 0.018821f $X=0.815 $Y=2.38 $X2=0
+ $Y2=0
cc_261 N_A_117_297#_c_339_n N_VPWR_c_426_n 0.0485782f $X=2.575 $Y=2.38 $X2=0
+ $Y2=0
cc_262 N_A_117_297#_c_350_n N_VPWR_c_426_n 0.0155188f $X=2.7 $Y=2.295 $X2=0
+ $Y2=0
cc_263 N_A_117_297#_c_406_p N_VPWR_c_426_n 0.0119021f $X=1.67 $Y=2.38 $X2=0
+ $Y2=0
cc_264 N_A_117_297#_c_360_n N_VPWR_c_428_n 0.0294205f $X=3.7 $Y=1.66 $X2=0 $Y2=0
cc_265 N_A_117_297#_c_342_n N_VPWR_c_430_n 0.0244686f $X=4.64 $Y=1.66 $X2=0
+ $Y2=0
cc_266 N_A_117_297#_M1000_s N_VPWR_c_423_n 0.00231266f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_267 N_A_117_297#_M1009_s N_VPWR_c_423_n 0.00231272f $X=1.525 $Y=1.485 $X2=0
+ $Y2=0
cc_268 N_A_117_297#_M1003_d N_VPWR_c_423_n 0.00217521f $X=2.535 $Y=1.485 $X2=0
+ $Y2=0
cc_269 N_A_117_297#_M1006_d N_VPWR_c_423_n 0.00312363f $X=3.455 $Y=1.485 $X2=0
+ $Y2=0
cc_270 N_A_117_297#_M1015_d N_VPWR_c_423_n 0.00217517f $X=4.495 $Y=1.485 $X2=0
+ $Y2=0
cc_271 N_A_117_297#_c_345_n N_VPWR_c_423_n 0.0268781f $X=1.585 $Y=2.38 $X2=0
+ $Y2=0
cc_272 N_A_117_297#_c_346_n N_VPWR_c_423_n 0.0111382f $X=0.815 $Y=2.38 $X2=0
+ $Y2=0
cc_273 N_A_117_297#_c_339_n N_VPWR_c_423_n 0.0296368f $X=2.575 $Y=2.38 $X2=0
+ $Y2=0
cc_274 N_A_117_297#_c_350_n N_VPWR_c_423_n 0.00946403f $X=2.7 $Y=2.295 $X2=0
+ $Y2=0
cc_275 N_A_117_297#_c_360_n N_VPWR_c_423_n 0.0179337f $X=3.7 $Y=1.66 $X2=0 $Y2=0
cc_276 N_A_117_297#_c_342_n N_VPWR_c_423_n 0.0141694f $X=4.64 $Y=1.66 $X2=0
+ $Y2=0
cc_277 N_A_117_297#_c_406_p N_VPWR_c_423_n 0.00653671f $X=1.67 $Y=2.38 $X2=0
+ $Y2=0
cc_278 N_A_117_297#_c_341_n N_A_507_47#_c_585_n 0.00625864f $X=4.425 $Y=1.57
+ $X2=0 $Y2=0
cc_279 N_A_117_297#_c_343_n N_A_507_47#_c_591_n 0.0051163f $X=3.625 $Y=1.57
+ $X2=0 $Y2=0
cc_280 N_A_27_47#_c_489_n N_VGND_M1001_s 0.00445216f $X=1.115 $Y=0.765 $X2=-0.19
+ $Y2=-0.24
cc_281 N_A_27_47#_c_489_n N_VGND_c_523_n 0.00281019f $X=1.115 $Y=0.765 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_508_p N_VGND_c_523_n 0.0113602f $X=1.285 $Y=0.38 $X2=0 $Y2=0
cc_283 N_A_27_47#_c_487_n N_VGND_c_523_n 0.0592143f $X=2.14 $Y=0.42 $X2=0 $Y2=0
cc_284 N_A_27_47#_c_485_n N_VGND_c_526_n 0.0173223f $X=0.22 $Y=0.68 $X2=0 $Y2=0
cc_285 N_A_27_47#_c_489_n N_VGND_c_526_n 0.00219121f $X=1.115 $Y=0.765 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_M1001_d N_VGND_c_528_n 0.00295891f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_M1011_d N_VGND_c_528_n 0.00238334f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_M1012_s N_VGND_c_528_n 0.00209344f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_485_n N_VGND_c_528_n 0.00951769f $X=0.22 $Y=0.68 $X2=0 $Y2=0
cc_290 N_A_27_47#_c_489_n N_VGND_c_528_n 0.0110524f $X=1.115 $Y=0.765 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_508_p N_VGND_c_528_n 0.00652422f $X=1.285 $Y=0.38 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_487_n N_VGND_c_528_n 0.0368686f $X=2.14 $Y=0.42 $X2=0 $Y2=0
cc_293 N_A_27_47#_c_485_n N_VGND_c_529_n 0.0195878f $X=0.22 $Y=0.68 $X2=0 $Y2=0
cc_294 N_A_27_47#_c_489_n N_VGND_c_529_n 0.0216074f $X=1.115 $Y=0.765 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_487_n N_A_507_47#_c_584_n 0.0214677f $X=2.14 $Y=0.42 $X2=0
+ $Y2=0
cc_296 N_VGND_c_528_n N_A_507_47#_M1002_d 0.00250339f $X=4.83 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_297 N_VGND_c_528_n N_A_507_47#_M1007_d 0.00318642f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_298 N_VGND_c_528_n N_A_507_47#_M1013_d 0.00230841f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_299 N_VGND_c_523_n N_A_507_47#_c_584_n 0.0770817f $X=3.98 $Y=0 $X2=0 $Y2=0
cc_300 N_VGND_c_528_n N_A_507_47#_c_584_n 0.0471488f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_301 N_VGND_M1005_s N_A_507_47#_c_585_n 0.0052865f $X=3.985 $Y=0.235 $X2=0
+ $Y2=0
cc_302 N_VGND_c_522_n N_A_507_47#_c_585_n 0.020293f $X=4.17 $Y=0.4 $X2=0 $Y2=0
cc_303 N_VGND_c_523_n N_A_507_47#_c_585_n 0.00256227f $X=3.98 $Y=0 $X2=0 $Y2=0
cc_304 N_VGND_c_527_n N_A_507_47#_c_585_n 0.00256227f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_305 N_VGND_c_528_n N_A_507_47#_c_585_n 0.0108045f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_306 N_VGND_c_527_n N_A_507_47#_c_586_n 0.0220856f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_307 N_VGND_c_528_n N_A_507_47#_c_586_n 0.0122041f $X=4.83 $Y=0 $X2=0 $Y2=0
