* File: sky130_fd_sc_hdll__mux2_8.pxi.spice
* Created: Wed Sep  2 08:34:44 2020
* 
x_PM_SKY130_FD_SC_HDLL__MUX2_8%A_79_21# N_A_79_21#_M1003_d N_A_79_21#_M1017_d
+ N_A_79_21#_M1002_s N_A_79_21#_M1016_s N_A_79_21#_c_122_n N_A_79_21#_M1006_g
+ N_A_79_21#_c_139_n N_A_79_21#_M1000_g N_A_79_21#_c_123_n N_A_79_21#_M1009_g
+ N_A_79_21#_c_140_n N_A_79_21#_M1001_g N_A_79_21#_c_124_n N_A_79_21#_M1010_g
+ N_A_79_21#_c_141_n N_A_79_21#_M1004_g N_A_79_21#_c_125_n N_A_79_21#_M1020_g
+ N_A_79_21#_c_142_n N_A_79_21#_M1008_g N_A_79_21#_c_126_n N_A_79_21#_M1026_g
+ N_A_79_21#_c_143_n N_A_79_21#_M1014_g N_A_79_21#_c_127_n N_A_79_21#_M1027_g
+ N_A_79_21#_c_144_n N_A_79_21#_M1018_g N_A_79_21#_c_128_n N_A_79_21#_M1029_g
+ N_A_79_21#_c_145_n N_A_79_21#_M1021_g N_A_79_21#_c_146_n N_A_79_21#_M1028_g
+ N_A_79_21#_c_129_n N_A_79_21#_M1030_g N_A_79_21#_c_279_p N_A_79_21#_c_130_n
+ N_A_79_21#_c_131_n N_A_79_21#_c_152_p N_A_79_21#_c_302_p N_A_79_21#_c_231_p
+ N_A_79_21#_c_153_p N_A_79_21#_c_186_p N_A_79_21#_c_132_n N_A_79_21#_c_133_n
+ N_A_79_21#_c_134_n N_A_79_21#_c_135_n N_A_79_21#_c_136_n N_A_79_21#_c_137_n
+ N_A_79_21#_c_138_n PM_SKY130_FD_SC_HDLL__MUX2_8%A_79_21#
x_PM_SKY130_FD_SC_HDLL__MUX2_8%S N_S_c_400_n N_S_M1022_g N_S_c_401_n N_S_M1007_g
+ N_S_c_402_n N_S_M1033_g N_S_c_403_n N_S_M1023_g N_S_c_404_n N_S_M1032_g
+ N_S_c_405_n N_S_M1019_g N_S_c_406_n N_S_c_437_n N_S_c_440_n N_S_c_441_n
+ N_S_c_407_n N_S_c_414_n N_S_c_415_n S N_S_c_408_n
+ PM_SKY130_FD_SC_HDLL__MUX2_8%S
x_PM_SKY130_FD_SC_HDLL__MUX2_8%A1 N_A1_c_548_n N_A1_M1003_g N_A1_c_549_n
+ N_A1_M1005_g N_A1_c_555_n N_A1_M1016_g N_A1_c_556_n N_A1_M1024_g N_A1_c_550_n
+ N_A1_c_551_n A1 N_A1_c_558_n N_A1_c_552_n N_A1_c_553_n
+ PM_SKY130_FD_SC_HDLL__MUX2_8%A1
x_PM_SKY130_FD_SC_HDLL__MUX2_8%A0 N_A0_c_651_n N_A0_M1002_g N_A0_c_652_n
+ N_A0_M1012_g N_A0_c_644_n N_A0_M1017_g N_A0_c_645_n N_A0_c_646_n N_A0_M1031_g
+ N_A0_c_647_n N_A0_c_672_n N_A0_c_648_n N_A0_c_677_n N_A0_c_649_n A0
+ N_A0_c_650_n N_A0_c_683_n A0 N_A0_c_684_n PM_SKY130_FD_SC_HDLL__MUX2_8%A0
x_PM_SKY130_FD_SC_HDLL__MUX2_8%A_1369_199# N_A_1369_199#_M1032_d
+ N_A_1369_199#_M1019_d N_A_1369_199#_c_764_n N_A_1369_199#_M1013_g
+ N_A_1369_199#_c_765_n N_A_1369_199#_M1011_g N_A_1369_199#_c_766_n
+ N_A_1369_199#_M1025_g N_A_1369_199#_c_767_n N_A_1369_199#_M1015_g
+ N_A_1369_199#_c_768_n N_A_1369_199#_c_778_n N_A_1369_199#_c_781_n
+ N_A_1369_199#_c_769_n N_A_1369_199#_c_806_n N_A_1369_199#_c_871_p
+ N_A_1369_199#_c_810_n N_A_1369_199#_c_851_p N_A_1369_199#_c_878_p
+ N_A_1369_199#_c_814_n N_A_1369_199#_c_853_p N_A_1369_199#_c_816_n
+ PM_SKY130_FD_SC_HDLL__MUX2_8%A_1369_199#
x_PM_SKY130_FD_SC_HDLL__MUX2_8%VPWR N_VPWR_M1000_d N_VPWR_M1001_d N_VPWR_M1008_d
+ N_VPWR_M1018_d N_VPWR_M1028_d N_VPWR_M1033_s N_VPWR_M1015_d N_VPWR_c_890_n
+ N_VPWR_c_891_n N_VPWR_c_892_n N_VPWR_c_893_n N_VPWR_c_894_n N_VPWR_c_895_n
+ N_VPWR_c_896_n N_VPWR_c_897_n VPWR N_VPWR_c_898_n N_VPWR_c_899_n
+ N_VPWR_c_900_n N_VPWR_c_901_n N_VPWR_c_902_n N_VPWR_c_903_n N_VPWR_c_889_n
+ N_VPWR_c_905_n N_VPWR_c_906_n N_VPWR_c_907_n N_VPWR_c_908_n N_VPWR_c_909_n
+ PM_SKY130_FD_SC_HDLL__MUX2_8%VPWR
x_PM_SKY130_FD_SC_HDLL__MUX2_8%X N_X_M1006_d N_X_M1010_d N_X_M1026_d N_X_M1029_d
+ N_X_M1000_s N_X_M1004_s N_X_M1014_s N_X_M1021_s N_X_c_1032_n N_X_c_1033_n
+ N_X_c_1034_n N_X_c_1038_n N_X_c_1119_p N_X_c_1042_n N_X_c_1044_n N_X_c_1048_n
+ N_X_c_1052_n N_X_c_1053_n N_X_c_1055_n N_X_c_1061_n N_X_c_1125_p N_X_c_1067_n
+ N_X_c_1071_n N_X_c_1073_n N_X_c_1075_n N_X_c_1077_n N_X_c_1079_n X
+ PM_SKY130_FD_SC_HDLL__MUX2_8%X
x_PM_SKY130_FD_SC_HDLL__MUX2_8%A_870_297# N_A_870_297#_M1022_d
+ N_A_870_297#_M1012_d N_A_870_297#_c_1147_n
+ PM_SKY130_FD_SC_HDLL__MUX2_8%A_870_297#
x_PM_SKY130_FD_SC_HDLL__MUX2_8%A_1420_297# N_A_1420_297#_M1013_s
+ N_A_1420_297#_M1024_d N_A_1420_297#_c_1163_n
+ PM_SKY130_FD_SC_HDLL__MUX2_8%A_1420_297#
x_PM_SKY130_FD_SC_HDLL__MUX2_8%VGND N_VGND_M1006_s N_VGND_M1009_s N_VGND_M1020_s
+ N_VGND_M1027_s N_VGND_M1030_s N_VGND_M1023_d N_VGND_M1025_d N_VGND_c_1179_n
+ N_VGND_c_1180_n N_VGND_c_1181_n VGND N_VGND_c_1182_n N_VGND_c_1183_n
+ N_VGND_c_1184_n N_VGND_c_1185_n N_VGND_c_1186_n N_VGND_c_1187_n
+ N_VGND_c_1188_n N_VGND_c_1189_n N_VGND_c_1190_n N_VGND_c_1191_n
+ N_VGND_c_1192_n N_VGND_c_1193_n N_VGND_c_1194_n N_VGND_c_1195_n
+ PM_SKY130_FD_SC_HDLL__MUX2_8%VGND
x_PM_SKY130_FD_SC_HDLL__MUX2_8%A_872_47# N_A_872_47#_M1007_s N_A_872_47#_M1005_s
+ N_A_872_47#_c_1334_n PM_SKY130_FD_SC_HDLL__MUX2_8%A_872_47#
x_PM_SKY130_FD_SC_HDLL__MUX2_8%A_1422_47# N_A_1422_47#_M1011_s
+ N_A_1422_47#_M1031_s N_A_1422_47#_c_1355_n
+ PM_SKY130_FD_SC_HDLL__MUX2_8%A_1422_47#
cc_1 VNB N_A_79_21#_c_122_n 0.0215258f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_123_n 0.0166773f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_3 VNB N_A_79_21#_c_124_n 0.0167353f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_4 VNB N_A_79_21#_c_125_n 0.0167427f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.995
cc_5 VNB N_A_79_21#_c_126_n 0.0167427f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=0.995
cc_6 VNB N_A_79_21#_c_127_n 0.0167427f $X=-0.19 $Y=-0.24 $X2=2.82 $Y2=0.995
cc_7 VNB N_A_79_21#_c_128_n 0.0171735f $X=-0.19 $Y=-0.24 $X2=3.29 $Y2=0.995
cc_8 VNB N_A_79_21#_c_129_n 0.01648f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.995
cc_9 VNB N_A_79_21#_c_130_n 0.00157396f $X=-0.19 $Y=-0.24 $X2=3.89 $Y2=1.075
cc_10 VNB N_A_79_21#_c_131_n 3.47426e-19 $X=-0.19 $Y=-0.24 $X2=3.89 $Y2=1.835
cc_11 VNB N_A_79_21#_c_132_n 0.00102315f $X=-0.19 $Y=-0.24 $X2=3.89 $Y2=1.16
cc_12 VNB N_A_79_21#_c_133_n 0.00991546f $X=-0.19 $Y=-0.24 $X2=8.09 $Y2=0.85
cc_13 VNB N_A_79_21#_c_134_n 0.00119944f $X=-0.19 $Y=-0.24 $X2=5.4 $Y2=0.85
cc_14 VNB N_A_79_21#_c_135_n 0.00487674f $X=-0.19 $Y=-0.24 $X2=8.235 $Y2=0.85
cc_15 VNB N_A_79_21#_c_136_n 0.16124f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.202
cc_16 VNB N_A_79_21#_c_137_n 0.0012422f $X=-0.19 $Y=-0.24 $X2=5.255 $Y2=0.72
cc_17 VNB N_A_79_21#_c_138_n 0.0016504f $X=-0.19 $Y=-0.24 $X2=8.26 $Y2=0.72
cc_18 VNB N_S_c_400_n 0.02574f $X=-0.19 $Y=-0.24 $X2=4.805 $Y2=0.235
cc_19 VNB N_S_c_401_n 0.0177581f $X=-0.19 $Y=-0.24 $X2=8.665 $Y2=1.485
cc_20 VNB N_S_c_402_n 0.0226618f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_S_c_403_n 0.0220282f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_S_c_404_n 0.022747f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_23 VNB N_S_c_405_n 0.0381652f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_24 VNB N_S_c_406_n 6.24445e-19 $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_25 VNB N_S_c_407_n 0.00418629f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_26 VNB N_S_c_408_n 0.00450635f $X=-0.19 $Y=-0.24 $X2=2.82 $Y2=0.995
cc_27 VNB N_A1_c_548_n 0.0151583f $X=-0.19 $Y=-0.24 $X2=4.805 $Y2=0.235
cc_28 VNB N_A1_c_549_n 0.0519005f $X=-0.19 $Y=-0.24 $X2=8.665 $Y2=1.485
cc_29 VNB N_A1_c_550_n 0.0108181f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_30 VNB N_A1_c_551_n 0.00223999f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_31 VNB N_A1_c_552_n 0.064466f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_32 VNB N_A1_c_553_n 0.00306074f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_33 VNB N_A0_c_644_n 0.0297217f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A0_c_645_n 0.0297823f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A0_c_646_n 0.0189956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A0_c_647_n 0.00244117f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_37 VNB N_A0_c_648_n 0.00256383f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_38 VNB N_A0_c_649_n 0.00397827f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_39 VNB N_A0_c_650_n 0.0502369f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_40 VNB N_A_1369_199#_c_764_n 0.0288786f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_1369_199#_c_765_n 0.0190435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_1369_199#_c_766_n 0.0234282f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_43 VNB N_A_1369_199#_c_767_n 0.0274913f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_44 VNB N_A_1369_199#_c_768_n 4.7857e-19 $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_45 VNB N_A_1369_199#_c_769_n 0.00135754f $X=-0.19 $Y=-0.24 $X2=1.435
+ $Y2=1.985
cc_46 VNB N_VPWR_c_889_n 0.440529f $X=-0.19 $Y=-0.24 $X2=7.93 $Y2=0.72
cc_47 VNB X 0.00208947f $X=-0.19 $Y=-0.24 $X2=3.975 $Y2=1.92
cc_48 VNB N_VGND_c_1179_n 0.0102396f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_49 VNB N_VGND_c_1180_n 0.0133473f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_50 VNB N_VGND_c_1181_n 0.00281836f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_51 VNB N_VGND_c_1182_n 0.0129637f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_52 VNB N_VGND_c_1183_n 0.012495f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=0.995
cc_53 VNB N_VGND_c_1184_n 0.0123761f $X=-0.19 $Y=-0.24 $X2=2.375 $Y2=1.985
cc_54 VNB N_VGND_c_1185_n 0.0132631f $X=-0.19 $Y=-0.24 $X2=2.845 $Y2=1.985
cc_55 VNB N_VGND_c_1186_n 0.0616f $X=-0.19 $Y=-0.24 $X2=3.315 $Y2=1.41
cc_56 VNB N_VGND_c_1187_n 0.0700793f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.985
cc_57 VNB N_VGND_c_1188_n 0.0159282f $X=-0.19 $Y=-0.24 $X2=3.54 $Y2=1.16
cc_58 VNB N_VGND_c_1189_n 0.489909f $X=-0.19 $Y=-0.24 $X2=3.54 $Y2=1.16
cc_59 VNB N_VGND_c_1190_n 0.00537041f $X=-0.19 $Y=-0.24 $X2=4.94 $Y2=0.72
cc_60 VNB N_VGND_c_1191_n 0.00537882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1192_n 0.00537882f $X=-0.19 $Y=-0.24 $X2=5.4 $Y2=0.85
cc_62 VNB N_VGND_c_1193_n 0.00845922f $X=-0.19 $Y=-0.24 $X2=8.235 $Y2=0.85
cc_63 VNB N_VGND_c_1194_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=1.25 $Y2=1.202
cc_64 VNB N_VGND_c_1195_n 0.00860652f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_65 VPB N_A_79_21#_c_139_n 0.0202186f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_66 VPB N_A_79_21#_c_140_n 0.0157869f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_67 VPB N_A_79_21#_c_141_n 0.0160885f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_68 VPB N_A_79_21#_c_142_n 0.0158129f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_69 VPB N_A_79_21#_c_143_n 0.0160921f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_70 VPB N_A_79_21#_c_144_n 0.0158129f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_71 VPB N_A_79_21#_c_145_n 0.016086f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.41
cc_72 VPB N_A_79_21#_c_146_n 0.0155343f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_73 VPB N_A_79_21#_c_131_n 0.00108787f $X=-0.19 $Y=1.305 $X2=3.89 $Y2=1.835
cc_74 VPB N_A_79_21#_c_136_n 0.104523f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.202
cc_75 VPB N_S_c_400_n 0.0297946f $X=-0.19 $Y=1.305 $X2=4.805 $Y2=0.235
cc_76 VPB N_S_c_402_n 0.0257407f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_S_c_405_n 0.032677f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_78 VPB N_S_c_406_n 0.00664512f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_79 VPB N_S_c_407_n 0.00320975f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_80 VPB N_S_c_414_n 0.0225454f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=0.995
cc_81 VPB N_S_c_415_n 0.00137569f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=0.56
cc_82 VPB S 0.00104623f $X=-0.19 $Y=1.305 $X2=2.35 $Y2=0.995
cc_83 VPB N_S_c_408_n 0.00706769f $X=-0.19 $Y=1.305 $X2=2.82 $Y2=0.995
cc_84 VPB N_A1_c_549_n 0.0172424f $X=-0.19 $Y=1.305 $X2=8.665 $Y2=1.485
cc_85 VPB N_A1_c_555_n 0.0206328f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A1_c_556_n 0.0161215f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A1_c_551_n 2.57451e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_88 VPB N_A1_c_558_n 0.00204052f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=0.995
cc_89 VPB N_A1_c_552_n 0.0174194f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=0.56
cc_90 VPB N_A1_c_553_n 3.16598e-19 $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_91 VPB N_A0_c_651_n 0.0210142f $X=-0.19 $Y=1.305 $X2=4.805 $Y2=0.235
cc_92 VPB N_A0_c_652_n 0.0163411f $X=-0.19 $Y=1.305 $X2=8.665 $Y2=1.485
cc_93 VPB N_A0_c_644_n 0.00550272f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A0_c_645_n 0.0148999f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A0_c_649_n 0.0016233f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=0.995
cc_96 VPB N_A0_c_650_n 0.0175401f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_97 VPB N_A_1369_199#_c_764_n 0.0322252f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_1369_199#_c_767_n 0.0263082f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_99 VPB N_A_1369_199#_c_768_n 0.00628483f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_100 VPB N_A_1369_199#_c_769_n 0.00175739f $X=-0.19 $Y=1.305 $X2=1.435
+ $Y2=1.985
cc_101 VPB N_VPWR_c_890_n 0.010306f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_102 VPB N_VPWR_c_891_n 0.0266961f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_103 VPB N_VPWR_c_892_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_104 VPB N_VPWR_c_893_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=1.88 $Y2=0.56
cc_105 VPB N_VPWR_c_894_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_106 VPB N_VPWR_c_895_n 0.00474148f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_107 VPB N_VPWR_c_896_n 0.060035f $X=-0.19 $Y=1.305 $X2=2.82 $Y2=0.995
cc_108 VPB N_VPWR_c_897_n 0.0032427f $X=-0.19 $Y=1.305 $X2=2.82 $Y2=0.56
cc_109 VPB N_VPWR_c_898_n 0.0137063f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.985
cc_110 VPB N_VPWR_c_899_n 0.0140826f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.41
cc_111 VPB N_VPWR_c_900_n 0.0140826f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.985
cc_112 VPB N_VPWR_c_901_n 0.0141085f $X=-0.19 $Y=1.305 $X2=1.25 $Y2=1.16
cc_113 VPB N_VPWR_c_902_n 0.0670602f $X=-0.19 $Y=1.305 $X2=3.975 $Y2=0.72
cc_114 VPB N_VPWR_c_903_n 0.0157945f $X=-0.19 $Y=1.305 $X2=8.15 $Y2=0.72
cc_115 VPB N_VPWR_c_889_n 0.0489137f $X=-0.19 $Y=1.305 $X2=7.93 $Y2=0.72
cc_116 VPB N_VPWR_c_905_n 0.00503453f $X=-0.19 $Y=1.305 $X2=5.255 $Y2=0.85
cc_117 VPB N_VPWR_c_906_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_907_n 0.00503453f $X=-0.19 $Y=1.305 $X2=8.235 $Y2=0.85
cc_119 VPB N_VPWR_c_908_n 0.0054644f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_120 VPB N_VPWR_c_909_n 0.00872118f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_121 VPB X 0.00264212f $X=-0.19 $Y=1.305 $X2=3.975 $Y2=1.92
cc_122 N_A_79_21#_c_146_n N_S_c_400_n 0.0362983f $X=3.785 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_123 N_A_79_21#_c_130_n N_S_c_400_n 4.63096e-19 $X=3.89 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_124 N_A_79_21#_c_131_n N_S_c_400_n 0.00493132f $X=3.89 $Y=1.835 $X2=-0.19
+ $Y2=-0.24
cc_125 N_A_79_21#_c_152_p N_S_c_400_n 0.00333858f $X=5.17 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_126 N_A_79_21#_c_153_p N_S_c_400_n 0.0167671f $X=8.81 $Y=1.92 $X2=-0.19
+ $Y2=-0.24
cc_127 N_A_79_21#_c_132_n N_S_c_400_n 0.00115091f $X=3.89 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_128 N_A_79_21#_c_136_n N_S_c_400_n 0.0244902f $X=3.785 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_129 N_A_79_21#_c_129_n N_S_c_401_n 0.020266f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_79_21#_c_130_n N_S_c_401_n 0.00369234f $X=3.89 $Y=1.075 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_152_p N_S_c_401_n 0.0121866f $X=5.17 $Y=0.72 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_153_p N_S_c_402_n 0.015004f $X=8.81 $Y=1.92 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_133_n N_S_c_402_n 8.26873e-19 $X=8.09 $Y=0.85 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_133_n N_S_c_403_n 0.00341729f $X=8.09 $Y=0.85 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_146_n N_S_c_406_n 2.01092e-19 $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_130_n N_S_c_406_n 0.00579357f $X=3.89 $Y=1.075 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_131_n N_S_c_406_n 0.0184028f $X=3.89 $Y=1.835 $X2=0 $Y2=0
cc_138 N_A_79_21#_c_152_p N_S_c_406_n 0.0132818f $X=5.17 $Y=0.72 $X2=0 $Y2=0
cc_139 N_A_79_21#_c_132_n N_S_c_406_n 0.0139493f $X=3.89 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A_79_21#_c_136_n N_S_c_406_n 5.44659e-19 $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_141 N_A_79_21#_M1002_s N_S_c_437_n 0.00339645f $X=5.625 $Y=1.485 $X2=0 $Y2=0
cc_142 N_A_79_21#_c_153_p N_S_c_437_n 0.106911f $X=8.81 $Y=1.92 $X2=0 $Y2=0
cc_143 N_A_79_21#_c_137_n N_S_c_437_n 0.0025162f $X=5.255 $Y=0.72 $X2=0 $Y2=0
cc_144 N_A_79_21#_c_153_p N_S_c_440_n 0.0136945f $X=8.81 $Y=1.92 $X2=0 $Y2=0
cc_145 N_A_79_21#_c_153_p N_S_c_441_n 0.0244507f $X=8.81 $Y=1.92 $X2=0 $Y2=0
cc_146 N_A_79_21#_c_133_n N_S_c_407_n 0.00337413f $X=8.09 $Y=0.85 $X2=0 $Y2=0
cc_147 N_A_79_21#_c_153_p N_S_c_414_n 0.0277242f $X=8.81 $Y=1.92 $X2=0 $Y2=0
cc_148 N_A_79_21#_c_153_p N_S_c_415_n 0.00208167f $X=8.81 $Y=1.92 $X2=0 $Y2=0
cc_149 N_A_79_21#_c_152_p N_A1_c_548_n 0.00865779f $X=5.17 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_150 N_A_79_21#_c_134_n N_A1_c_548_n 6.81815e-19 $X=5.4 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_151 N_A_79_21#_c_137_n N_A1_c_548_n 9.64511e-19 $X=5.255 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_152 N_A_79_21#_c_152_p N_A1_c_549_n 0.00806459f $X=5.17 $Y=0.72 $X2=0 $Y2=0
cc_153 N_A_79_21#_c_134_n N_A1_c_549_n 0.00405063f $X=5.4 $Y=0.85 $X2=0 $Y2=0
cc_154 N_A_79_21#_c_137_n N_A1_c_549_n 0.0108837f $X=5.255 $Y=0.72 $X2=0 $Y2=0
cc_155 N_A_79_21#_c_153_p N_A1_c_555_n 0.0122583f $X=8.81 $Y=1.92 $X2=0 $Y2=0
cc_156 N_A_79_21#_c_153_p N_A1_c_556_n 0.00331994f $X=8.81 $Y=1.92 $X2=0 $Y2=0
cc_157 N_A_79_21#_c_152_p N_A1_c_550_n 0.00587314f $X=5.17 $Y=0.72 $X2=0 $Y2=0
cc_158 N_A_79_21#_c_153_p N_A1_c_550_n 3.94934e-19 $X=8.81 $Y=1.92 $X2=0 $Y2=0
cc_159 N_A_79_21#_c_186_p N_A1_c_550_n 0.00193289f $X=8.15 $Y=0.72 $X2=0 $Y2=0
cc_160 N_A_79_21#_c_133_n N_A1_c_550_n 0.214283f $X=8.09 $Y=0.85 $X2=0 $Y2=0
cc_161 N_A_79_21#_c_134_n N_A1_c_550_n 0.0276841f $X=5.4 $Y=0.85 $X2=0 $Y2=0
cc_162 N_A_79_21#_c_135_n N_A1_c_550_n 0.0322629f $X=8.235 $Y=0.85 $X2=0 $Y2=0
cc_163 N_A_79_21#_c_137_n N_A1_c_550_n 8.22363e-19 $X=5.255 $Y=0.72 $X2=0 $Y2=0
cc_164 N_A_79_21#_c_138_n N_A1_c_550_n 0.00118207f $X=8.26 $Y=0.72 $X2=0 $Y2=0
cc_165 N_A_79_21#_c_152_p N_A1_c_551_n 0.00576993f $X=5.17 $Y=0.72 $X2=0 $Y2=0
cc_166 N_A_79_21#_c_152_p N_A1_c_558_n 0.012318f $X=5.17 $Y=0.72 $X2=0 $Y2=0
cc_167 N_A_79_21#_c_153_p N_A0_c_651_n 0.0123212f $X=8.81 $Y=1.92 $X2=-0.19
+ $Y2=-0.24
cc_168 N_A_79_21#_c_153_p N_A0_c_652_n 0.0102783f $X=8.81 $Y=1.92 $X2=0 $Y2=0
cc_169 N_A_79_21#_c_186_p N_A0_c_644_n 0.00263741f $X=8.15 $Y=0.72 $X2=0 $Y2=0
cc_170 N_A_79_21#_c_133_n N_A0_c_644_n 0.00400797f $X=8.09 $Y=0.85 $X2=0 $Y2=0
cc_171 N_A_79_21#_c_135_n N_A0_c_644_n 5.80314e-19 $X=8.235 $Y=0.85 $X2=0 $Y2=0
cc_172 N_A_79_21#_c_138_n N_A0_c_644_n 3.96886e-19 $X=8.26 $Y=0.72 $X2=0 $Y2=0
cc_173 N_A_79_21#_c_186_p N_A0_c_645_n 0.00653842f $X=8.15 $Y=0.72 $X2=0 $Y2=0
cc_174 N_A_79_21#_c_133_n N_A0_c_645_n 0.00324605f $X=8.09 $Y=0.85 $X2=0 $Y2=0
cc_175 N_A_79_21#_c_135_n N_A0_c_645_n 0.00137995f $X=8.235 $Y=0.85 $X2=0 $Y2=0
cc_176 N_A_79_21#_c_186_p N_A0_c_646_n 0.00209249f $X=8.15 $Y=0.72 $X2=0 $Y2=0
cc_177 N_A_79_21#_c_135_n N_A0_c_646_n 6.63251e-19 $X=8.235 $Y=0.85 $X2=0 $Y2=0
cc_178 N_A_79_21#_c_138_n N_A0_c_646_n 0.0135454f $X=8.26 $Y=0.72 $X2=0 $Y2=0
cc_179 N_A_79_21#_c_133_n N_A0_c_647_n 0.0106236f $X=8.09 $Y=0.85 $X2=0 $Y2=0
cc_180 N_A_79_21#_c_134_n N_A0_c_647_n 0.00192884f $X=5.4 $Y=0.85 $X2=0 $Y2=0
cc_181 N_A_79_21#_c_137_n N_A0_c_647_n 0.00585177f $X=5.255 $Y=0.72 $X2=0 $Y2=0
cc_182 N_A_79_21#_c_186_p N_A0_c_672_n 0.0104433f $X=8.15 $Y=0.72 $X2=0 $Y2=0
cc_183 N_A_79_21#_c_133_n N_A0_c_672_n 0.0390798f $X=8.09 $Y=0.85 $X2=0 $Y2=0
cc_184 N_A_79_21#_c_133_n N_A0_c_648_n 0.0104819f $X=8.09 $Y=0.85 $X2=0 $Y2=0
cc_185 N_A_79_21#_c_135_n N_A0_c_648_n 0.00131668f $X=8.235 $Y=0.85 $X2=0 $Y2=0
cc_186 N_A_79_21#_c_138_n N_A0_c_648_n 0.00134402f $X=8.26 $Y=0.72 $X2=0 $Y2=0
cc_187 N_A_79_21#_c_133_n N_A0_c_677_n 0.00590559f $X=8.09 $Y=0.85 $X2=0 $Y2=0
cc_188 N_A_79_21#_c_134_n N_A0_c_677_n 0.00137765f $X=5.4 $Y=0.85 $X2=0 $Y2=0
cc_189 N_A_79_21#_c_137_n N_A0_c_677_n 0.00999032f $X=5.255 $Y=0.72 $X2=0 $Y2=0
cc_190 N_A_79_21#_c_186_p N_A0_c_649_n 0.006437f $X=8.15 $Y=0.72 $X2=0 $Y2=0
cc_191 N_A_79_21#_c_133_n N_A0_c_649_n 0.00376919f $X=8.09 $Y=0.85 $X2=0 $Y2=0
cc_192 N_A_79_21#_c_133_n N_A0_c_650_n 0.00897501f $X=8.09 $Y=0.85 $X2=0 $Y2=0
cc_193 N_A_79_21#_c_133_n N_A0_c_683_n 0.0199367f $X=8.09 $Y=0.85 $X2=0 $Y2=0
cc_194 N_A_79_21#_c_133_n N_A0_c_684_n 0.00670453f $X=8.09 $Y=0.85 $X2=0 $Y2=0
cc_195 N_A_79_21#_c_153_p N_A_1369_199#_c_764_n 0.0166371f $X=8.81 $Y=1.92 $X2=0
+ $Y2=0
cc_196 N_A_79_21#_c_133_n N_A_1369_199#_c_764_n 0.0027076f $X=8.09 $Y=0.85 $X2=0
+ $Y2=0
cc_197 N_A_79_21#_c_133_n N_A_1369_199#_c_765_n 0.00273034f $X=8.09 $Y=0.85
+ $X2=0 $Y2=0
cc_198 N_A_79_21#_c_133_n N_A_1369_199#_c_768_n 0.00169401f $X=8.09 $Y=0.85
+ $X2=0 $Y2=0
cc_199 N_A_79_21#_M1016_s N_A_1369_199#_c_778_n 0.00471432f $X=8.665 $Y=1.485
+ $X2=0 $Y2=0
cc_200 N_A_79_21#_c_153_p N_A_1369_199#_c_778_n 0.108892f $X=8.81 $Y=1.92 $X2=0
+ $Y2=0
cc_201 N_A_79_21#_c_138_n N_A_1369_199#_c_778_n 0.00351082f $X=8.26 $Y=0.72
+ $X2=0 $Y2=0
cc_202 N_A_79_21#_c_153_p N_A_1369_199#_c_781_n 0.0127022f $X=8.81 $Y=1.92 $X2=0
+ $Y2=0
cc_203 N_A_79_21#_c_131_n N_VPWR_M1028_d 0.00351098f $X=3.89 $Y=1.835 $X2=0
+ $Y2=0
cc_204 N_A_79_21#_c_231_p N_VPWR_M1028_d 5.35521e-19 $X=3.975 $Y=1.92 $X2=0
+ $Y2=0
cc_205 N_A_79_21#_c_153_p N_VPWR_M1028_d 0.00649549f $X=8.81 $Y=1.92 $X2=0 $Y2=0
cc_206 N_A_79_21#_c_153_p N_VPWR_M1033_s 0.00617601f $X=8.81 $Y=1.92 $X2=0 $Y2=0
cc_207 N_A_79_21#_c_139_n N_VPWR_c_891_n 0.011965f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A_79_21#_c_140_n N_VPWR_c_891_n 5.64468e-19 $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_209 N_A_79_21#_c_139_n N_VPWR_c_892_n 6.33692e-19 $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_210 N_A_79_21#_c_140_n N_VPWR_c_892_n 0.0141913f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A_79_21#_c_141_n N_VPWR_c_892_n 0.0107665f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A_79_21#_c_142_n N_VPWR_c_892_n 5.96427e-19 $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_213 N_A_79_21#_c_141_n N_VPWR_c_893_n 6.33692e-19 $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_214 N_A_79_21#_c_142_n N_VPWR_c_893_n 0.0141913f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A_79_21#_c_143_n N_VPWR_c_893_n 0.0107665f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A_79_21#_c_144_n N_VPWR_c_893_n 5.96427e-19 $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_217 N_A_79_21#_c_143_n N_VPWR_c_894_n 6.33692e-19 $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_218 N_A_79_21#_c_144_n N_VPWR_c_894_n 0.0141913f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_219 N_A_79_21#_c_145_n N_VPWR_c_894_n 0.0107665f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_220 N_A_79_21#_c_146_n N_VPWR_c_894_n 5.96427e-19 $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_221 N_A_79_21#_c_153_p N_VPWR_c_895_n 0.0127213f $X=8.81 $Y=1.92 $X2=0 $Y2=0
cc_222 N_A_79_21#_c_153_p N_VPWR_c_896_n 0.00942317f $X=8.81 $Y=1.92 $X2=0 $Y2=0
cc_223 N_A_79_21#_c_139_n N_VPWR_c_898_n 0.00622633f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_224 N_A_79_21#_c_140_n N_VPWR_c_898_n 0.00427505f $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_225 N_A_79_21#_c_141_n N_VPWR_c_899_n 0.00622633f $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_226 N_A_79_21#_c_142_n N_VPWR_c_899_n 0.00427505f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_227 N_A_79_21#_c_143_n N_VPWR_c_900_n 0.00622633f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_228 N_A_79_21#_c_144_n N_VPWR_c_900_n 0.00427505f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_229 N_A_79_21#_c_145_n N_VPWR_c_901_n 0.00622633f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_230 N_A_79_21#_c_146_n N_VPWR_c_901_n 0.00429282f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_231 N_A_79_21#_c_153_p N_VPWR_c_902_n 0.00221628f $X=8.81 $Y=1.92 $X2=0 $Y2=0
cc_232 N_A_79_21#_M1002_s N_VPWR_c_889_n 0.00235479f $X=5.625 $Y=1.485 $X2=0
+ $Y2=0
cc_233 N_A_79_21#_M1016_s N_VPWR_c_889_n 0.00235479f $X=8.665 $Y=1.485 $X2=0
+ $Y2=0
cc_234 N_A_79_21#_c_139_n N_VPWR_c_889_n 0.0104011f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A_79_21#_c_140_n N_VPWR_c_889_n 0.00732977f $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_236 N_A_79_21#_c_141_n N_VPWR_c_889_n 0.0104011f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_237 N_A_79_21#_c_142_n N_VPWR_c_889_n 0.00732977f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_238 N_A_79_21#_c_143_n N_VPWR_c_889_n 0.0104011f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_239 N_A_79_21#_c_144_n N_VPWR_c_889_n 0.00732977f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_240 N_A_79_21#_c_145_n N_VPWR_c_889_n 0.0104011f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_241 N_A_79_21#_c_146_n N_VPWR_c_889_n 0.00732982f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_242 N_A_79_21#_c_231_p N_VPWR_c_889_n 8.63719e-19 $X=3.975 $Y=1.92 $X2=0
+ $Y2=0
cc_243 N_A_79_21#_c_153_p N_VPWR_c_889_n 0.0321736f $X=8.81 $Y=1.92 $X2=0 $Y2=0
cc_244 N_A_79_21#_c_145_n N_VPWR_c_908_n 5.36535e-19 $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_245 N_A_79_21#_c_146_n N_VPWR_c_908_n 0.00964424f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_246 N_A_79_21#_c_231_p N_VPWR_c_908_n 0.00639725f $X=3.975 $Y=1.92 $X2=0
+ $Y2=0
cc_247 N_A_79_21#_c_153_p N_VPWR_c_908_n 0.00829338f $X=8.81 $Y=1.92 $X2=0 $Y2=0
cc_248 N_A_79_21#_c_122_n N_X_c_1032_n 0.00420101f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A_79_21#_c_140_n N_X_c_1033_n 0.00514591f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_250 N_A_79_21#_c_123_n N_X_c_1034_n 0.0142863f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A_79_21#_c_124_n N_X_c_1034_n 0.0123454f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A_79_21#_c_279_p N_X_c_1034_n 0.0212919f $X=3.805 $Y=1.16 $X2=0 $Y2=0
cc_253 N_A_79_21#_c_136_n N_X_c_1034_n 0.00348793f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_254 N_A_79_21#_c_140_n N_X_c_1038_n 0.0204305f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_255 N_A_79_21#_c_141_n N_X_c_1038_n 0.0178982f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_256 N_A_79_21#_c_279_p N_X_c_1038_n 0.0174713f $X=3.805 $Y=1.16 $X2=0 $Y2=0
cc_257 N_A_79_21#_c_136_n N_X_c_1038_n 0.00626154f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_258 N_A_79_21#_c_141_n N_X_c_1042_n 0.00530373f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A_79_21#_c_142_n N_X_c_1042_n 0.00490547f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A_79_21#_c_125_n N_X_c_1044_n 0.0123454f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A_79_21#_c_126_n N_X_c_1044_n 0.0126234f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_262 N_A_79_21#_c_279_p N_X_c_1044_n 0.0314632f $X=3.805 $Y=1.16 $X2=0 $Y2=0
cc_263 N_A_79_21#_c_136_n N_X_c_1044_n 0.00348793f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_264 N_A_79_21#_c_142_n N_X_c_1048_n 0.0163691f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A_79_21#_c_143_n N_X_c_1048_n 0.0178982f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A_79_21#_c_279_p N_X_c_1048_n 0.0264364f $X=3.805 $Y=1.16 $X2=0 $Y2=0
cc_267 N_A_79_21#_c_136_n N_X_c_1048_n 0.00626154f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_268 N_A_79_21#_c_126_n N_X_c_1052_n 0.00391984f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_269 N_A_79_21#_c_143_n N_X_c_1053_n 0.00530373f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_270 N_A_79_21#_c_144_n N_X_c_1053_n 0.00490547f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_271 N_A_79_21#_c_127_n N_X_c_1055_n 0.0126234f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A_79_21#_c_128_n N_X_c_1055_n 0.012122f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A_79_21#_c_129_n N_X_c_1055_n 0.0013291f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A_79_21#_c_279_p N_X_c_1055_n 0.0406499f $X=3.805 $Y=1.16 $X2=0 $Y2=0
cc_275 N_A_79_21#_c_302_p N_X_c_1055_n 0.0148586f $X=3.975 $Y=0.72 $X2=0 $Y2=0
cc_276 N_A_79_21#_c_136_n N_X_c_1055_n 0.00760536f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_277 N_A_79_21#_c_144_n N_X_c_1061_n 0.016326f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_278 N_A_79_21#_c_145_n N_X_c_1061_n 0.0174108f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_279 N_A_79_21#_c_146_n N_X_c_1061_n 0.00141217f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_280 N_A_79_21#_c_279_p N_X_c_1061_n 0.0345056f $X=3.805 $Y=1.16 $X2=0 $Y2=0
cc_281 N_A_79_21#_c_131_n N_X_c_1061_n 0.013418f $X=3.89 $Y=1.835 $X2=0 $Y2=0
cc_282 N_A_79_21#_c_136_n N_X_c_1061_n 0.0103736f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_283 N_A_79_21#_c_145_n N_X_c_1067_n 0.00530373f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_284 N_A_79_21#_c_146_n N_X_c_1067_n 0.00626371f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_285 N_A_79_21#_c_131_n N_X_c_1067_n 0.00624815f $X=3.89 $Y=1.835 $X2=0 $Y2=0
cc_286 N_A_79_21#_c_231_p N_X_c_1067_n 0.0133617f $X=3.975 $Y=1.92 $X2=0 $Y2=0
cc_287 N_A_79_21#_c_122_n N_X_c_1071_n 0.00543425f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_288 N_A_79_21#_c_123_n N_X_c_1071_n 0.00178664f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_289 N_A_79_21#_c_279_p N_X_c_1073_n 0.00897186f $X=3.805 $Y=1.16 $X2=0 $Y2=0
cc_290 N_A_79_21#_c_136_n N_X_c_1073_n 0.00314844f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_291 N_A_79_21#_c_279_p N_X_c_1075_n 0.00806916f $X=3.805 $Y=1.16 $X2=0 $Y2=0
cc_292 N_A_79_21#_c_136_n N_X_c_1075_n 0.00424973f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_293 N_A_79_21#_c_279_p N_X_c_1077_n 0.00902757f $X=3.805 $Y=1.16 $X2=0 $Y2=0
cc_294 N_A_79_21#_c_136_n N_X_c_1077_n 0.0031577f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_295 N_A_79_21#_c_279_p N_X_c_1079_n 0.00806916f $X=3.805 $Y=1.16 $X2=0 $Y2=0
cc_296 N_A_79_21#_c_136_n N_X_c_1079_n 0.00424973f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_297 N_A_79_21#_c_122_n X 0.00495928f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_298 N_A_79_21#_c_139_n X 0.00246557f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_299 N_A_79_21#_c_123_n X 0.00351321f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_300 N_A_79_21#_c_140_n X 0.00250116f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_301 N_A_79_21#_c_279_p X 0.0107158f $X=3.805 $Y=1.16 $X2=0 $Y2=0
cc_302 N_A_79_21#_c_136_n X 0.0473071f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_303 N_A_79_21#_c_153_p N_A_870_297#_M1022_d 0.0300118f $X=8.81 $Y=1.92
+ $X2=-0.19 $Y2=-0.24
cc_304 N_A_79_21#_c_153_p N_A_870_297#_M1012_d 0.00384167f $X=8.81 $Y=1.92 $X2=0
+ $Y2=0
cc_305 N_A_79_21#_M1002_s N_A_870_297#_c_1147_n 0.00402806f $X=5.625 $Y=1.485
+ $X2=0 $Y2=0
cc_306 N_A_79_21#_c_153_p N_A_870_297#_c_1147_n 0.0719292f $X=8.81 $Y=1.92 $X2=0
+ $Y2=0
cc_307 N_A_79_21#_c_153_p N_A_1420_297#_M1013_s 0.0368158f $X=8.81 $Y=1.92
+ $X2=-0.19 $Y2=-0.24
cc_308 N_A_79_21#_M1016_s N_A_1420_297#_c_1163_n 0.00402806f $X=8.665 $Y=1.485
+ $X2=0 $Y2=0
cc_309 N_A_79_21#_c_153_p N_A_1420_297#_c_1163_n 0.0844077f $X=8.81 $Y=1.92
+ $X2=0 $Y2=0
cc_310 N_A_79_21#_c_130_n N_VGND_M1030_s 9.61388e-19 $X=3.89 $Y=1.075 $X2=0
+ $Y2=0
cc_311 N_A_79_21#_c_152_p N_VGND_M1030_s 0.00701181f $X=5.17 $Y=0.72 $X2=0 $Y2=0
cc_312 N_A_79_21#_c_302_p N_VGND_M1030_s 3.513e-19 $X=3.975 $Y=0.72 $X2=0 $Y2=0
cc_313 N_A_79_21#_c_122_n N_VGND_c_1180_n 0.00896034f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_314 N_A_79_21#_c_123_n N_VGND_c_1180_n 4.98922e-19 $X=0.94 $Y=0.995 $X2=0
+ $Y2=0
cc_315 N_A_79_21#_c_133_n N_VGND_c_1181_n 0.00128242f $X=8.09 $Y=0.85 $X2=0
+ $Y2=0
cc_316 N_A_79_21#_c_122_n N_VGND_c_1182_n 0.0046653f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_317 N_A_79_21#_c_123_n N_VGND_c_1182_n 0.00340075f $X=0.94 $Y=0.995 $X2=0
+ $Y2=0
cc_318 N_A_79_21#_c_124_n N_VGND_c_1183_n 0.00340075f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_319 N_A_79_21#_c_125_n N_VGND_c_1183_n 0.00340075f $X=1.88 $Y=0.995 $X2=0
+ $Y2=0
cc_320 N_A_79_21#_c_126_n N_VGND_c_1184_n 0.00340075f $X=2.35 $Y=0.995 $X2=0
+ $Y2=0
cc_321 N_A_79_21#_c_127_n N_VGND_c_1184_n 0.00340075f $X=2.82 $Y=0.995 $X2=0
+ $Y2=0
cc_322 N_A_79_21#_c_128_n N_VGND_c_1185_n 0.00340075f $X=3.29 $Y=0.995 $X2=0
+ $Y2=0
cc_323 N_A_79_21#_c_129_n N_VGND_c_1185_n 0.00273179f $X=3.81 $Y=0.995 $X2=0
+ $Y2=0
cc_324 N_A_79_21#_c_152_p N_VGND_c_1186_n 0.00261734f $X=5.17 $Y=0.72 $X2=0
+ $Y2=0
cc_325 N_A_79_21#_M1003_d N_VGND_c_1189_n 0.00219239f $X=4.805 $Y=0.235 $X2=0
+ $Y2=0
cc_326 N_A_79_21#_M1017_d N_VGND_c_1189_n 0.00246014f $X=7.745 $Y=0.235 $X2=0
+ $Y2=0
cc_327 N_A_79_21#_c_122_n N_VGND_c_1189_n 0.00801876f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_328 N_A_79_21#_c_123_n N_VGND_c_1189_n 0.00407108f $X=0.94 $Y=0.995 $X2=0
+ $Y2=0
cc_329 N_A_79_21#_c_124_n N_VGND_c_1189_n 0.00411893f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_330 N_A_79_21#_c_125_n N_VGND_c_1189_n 0.00411893f $X=1.88 $Y=0.995 $X2=0
+ $Y2=0
cc_331 N_A_79_21#_c_126_n N_VGND_c_1189_n 0.00407108f $X=2.35 $Y=0.995 $X2=0
+ $Y2=0
cc_332 N_A_79_21#_c_127_n N_VGND_c_1189_n 0.00407108f $X=2.82 $Y=0.995 $X2=0
+ $Y2=0
cc_333 N_A_79_21#_c_128_n N_VGND_c_1189_n 0.00423871f $X=3.29 $Y=0.995 $X2=0
+ $Y2=0
cc_334 N_A_79_21#_c_129_n N_VGND_c_1189_n 0.00522073f $X=3.81 $Y=0.995 $X2=0
+ $Y2=0
cc_335 N_A_79_21#_c_152_p N_VGND_c_1189_n 0.00646026f $X=5.17 $Y=0.72 $X2=0
+ $Y2=0
cc_336 N_A_79_21#_c_302_p N_VGND_c_1189_n 8.18865e-19 $X=3.975 $Y=0.72 $X2=0
+ $Y2=0
cc_337 N_A_79_21#_c_133_n N_VGND_c_1189_n 0.123536f $X=8.09 $Y=0.85 $X2=0 $Y2=0
cc_338 N_A_79_21#_c_134_n N_VGND_c_1189_n 0.0146876f $X=5.4 $Y=0.85 $X2=0 $Y2=0
cc_339 N_A_79_21#_c_135_n N_VGND_c_1189_n 0.017167f $X=8.235 $Y=0.85 $X2=0 $Y2=0
cc_340 N_A_79_21#_c_122_n N_VGND_c_1190_n 4.98468e-19 $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_341 N_A_79_21#_c_123_n N_VGND_c_1190_n 0.00701096f $X=0.94 $Y=0.995 $X2=0
+ $Y2=0
cc_342 N_A_79_21#_c_124_n N_VGND_c_1190_n 0.00752754f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_343 N_A_79_21#_c_125_n N_VGND_c_1190_n 5.94835e-19 $X=1.88 $Y=0.995 $X2=0
+ $Y2=0
cc_344 N_A_79_21#_c_124_n N_VGND_c_1191_n 5.82991e-19 $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_345 N_A_79_21#_c_125_n N_VGND_c_1191_n 0.00732961f $X=1.88 $Y=0.995 $X2=0
+ $Y2=0
cc_346 N_A_79_21#_c_126_n N_VGND_c_1191_n 0.00725547f $X=2.35 $Y=0.995 $X2=0
+ $Y2=0
cc_347 N_A_79_21#_c_127_n N_VGND_c_1191_n 5.13099e-19 $X=2.82 $Y=0.995 $X2=0
+ $Y2=0
cc_348 N_A_79_21#_c_126_n N_VGND_c_1192_n 4.98468e-19 $X=2.35 $Y=0.995 $X2=0
+ $Y2=0
cc_349 N_A_79_21#_c_127_n N_VGND_c_1192_n 0.00701096f $X=2.82 $Y=0.995 $X2=0
+ $Y2=0
cc_350 N_A_79_21#_c_128_n N_VGND_c_1192_n 0.00755689f $X=3.29 $Y=0.995 $X2=0
+ $Y2=0
cc_351 N_A_79_21#_c_129_n N_VGND_c_1192_n 5.60961e-19 $X=3.81 $Y=0.995 $X2=0
+ $Y2=0
cc_352 N_A_79_21#_c_128_n N_VGND_c_1193_n 6.19306e-19 $X=3.29 $Y=0.995 $X2=0
+ $Y2=0
cc_353 N_A_79_21#_c_129_n N_VGND_c_1193_n 0.00995499f $X=3.81 $Y=0.995 $X2=0
+ $Y2=0
cc_354 N_A_79_21#_c_152_p N_VGND_c_1193_n 0.013548f $X=5.17 $Y=0.72 $X2=0 $Y2=0
cc_355 N_A_79_21#_c_302_p N_VGND_c_1193_n 0.00898811f $X=3.975 $Y=0.72 $X2=0
+ $Y2=0
cc_356 N_A_79_21#_c_152_p N_A_872_47#_M1007_s 0.00864706f $X=5.17 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_357 N_A_79_21#_c_133_n N_A_872_47#_M1005_s 0.00191061f $X=8.09 $Y=0.85 $X2=0
+ $Y2=0
cc_358 N_A_79_21#_c_134_n N_A_872_47#_M1005_s 8.4102e-19 $X=5.4 $Y=0.85 $X2=0
+ $Y2=0
cc_359 N_A_79_21#_c_137_n N_A_872_47#_M1005_s 0.00278902f $X=5.255 $Y=0.72 $X2=0
+ $Y2=0
cc_360 N_A_79_21#_M1003_d N_A_872_47#_c_1334_n 0.00313811f $X=4.805 $Y=0.235
+ $X2=0 $Y2=0
cc_361 N_A_79_21#_c_152_p N_A_872_47#_c_1334_n 0.0384733f $X=5.17 $Y=0.72 $X2=0
+ $Y2=0
cc_362 N_A_79_21#_c_133_n N_A_872_47#_c_1334_n 0.00324871f $X=8.09 $Y=0.85 $X2=0
+ $Y2=0
cc_363 N_A_79_21#_c_134_n N_A_872_47#_c_1334_n 0.00241642f $X=5.4 $Y=0.85 $X2=0
+ $Y2=0
cc_364 N_A_79_21#_c_137_n N_A_872_47#_c_1334_n 0.00715296f $X=5.255 $Y=0.72
+ $X2=0 $Y2=0
cc_365 N_A_79_21#_c_133_n N_A_1422_47#_M1011_s 8.05638e-19 $X=8.09 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_366 N_A_79_21#_c_135_n N_A_1422_47#_M1031_s 0.00643896f $X=8.235 $Y=0.85
+ $X2=0 $Y2=0
cc_367 N_A_79_21#_c_138_n N_A_1422_47#_M1031_s 0.00681307f $X=8.26 $Y=0.72 $X2=0
+ $Y2=0
cc_368 N_A_79_21#_M1017_d N_A_1422_47#_c_1355_n 0.00507522f $X=7.745 $Y=0.235
+ $X2=0 $Y2=0
cc_369 N_A_79_21#_c_186_p N_A_1422_47#_c_1355_n 0.0202345f $X=8.15 $Y=0.72 $X2=0
+ $Y2=0
cc_370 N_A_79_21#_c_133_n N_A_1422_47#_c_1355_n 0.00467975f $X=8.09 $Y=0.85
+ $X2=0 $Y2=0
cc_371 N_A_79_21#_c_135_n N_A_1422_47#_c_1355_n 0.00257421f $X=8.235 $Y=0.85
+ $X2=0 $Y2=0
cc_372 N_A_79_21#_c_138_n N_A_1422_47#_c_1355_n 0.0102322f $X=8.26 $Y=0.72 $X2=0
+ $Y2=0
cc_373 N_S_c_401_n N_A1_c_548_n 0.0249936f $X=4.285 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_374 N_S_c_400_n N_A1_c_549_n 0.019159f $X=4.26 $Y=1.41 $X2=0 $Y2=0
cc_375 N_S_c_406_n N_A1_c_549_n 9.99501e-19 $X=4.23 $Y=1.16 $X2=0 $Y2=0
cc_376 N_S_c_437_n N_A1_c_549_n 0.0150307f $X=6.17 $Y=1.58 $X2=0 $Y2=0
cc_377 N_S_c_414_n N_A1_c_555_n 0.00257014f $X=9.745 $Y=1.53 $X2=0 $Y2=0
cc_378 N_S_c_414_n N_A1_c_556_n 0.0014559f $X=9.745 $Y=1.53 $X2=0 $Y2=0
cc_379 N_S_c_402_n N_A1_c_550_n 0.00108992f $X=6.475 $Y=1.41 $X2=0 $Y2=0
cc_380 N_S_c_437_n N_A1_c_550_n 0.0352437f $X=6.17 $Y=1.58 $X2=0 $Y2=0
cc_381 N_S_c_407_n N_A1_c_550_n 0.0210814f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_382 N_S_c_414_n N_A1_c_550_n 0.190979f $X=9.745 $Y=1.53 $X2=0 $Y2=0
cc_383 N_S_c_415_n N_A1_c_550_n 0.0255809f $X=6.4 $Y=1.53 $X2=0 $Y2=0
cc_384 N_S_c_400_n N_A1_c_551_n 0.00411408f $X=4.26 $Y=1.41 $X2=0 $Y2=0
cc_385 N_S_c_406_n N_A1_c_551_n 0.0070044f $X=4.23 $Y=1.16 $X2=0 $Y2=0
cc_386 N_S_c_437_n N_A1_c_551_n 0.00658346f $X=6.17 $Y=1.58 $X2=0 $Y2=0
cc_387 N_S_c_414_n A1 0.032133f $X=9.745 $Y=1.53 $X2=0 $Y2=0
cc_388 N_S_c_400_n N_A1_c_558_n 0.00136567f $X=4.26 $Y=1.41 $X2=0 $Y2=0
cc_389 N_S_c_406_n N_A1_c_558_n 0.0105012f $X=4.23 $Y=1.16 $X2=0 $Y2=0
cc_390 N_S_c_437_n N_A1_c_558_n 0.0155823f $X=6.17 $Y=1.58 $X2=0 $Y2=0
cc_391 N_S_c_414_n N_A1_c_552_n 0.00234049f $X=9.745 $Y=1.53 $X2=0 $Y2=0
cc_392 N_S_c_414_n N_A1_c_553_n 0.00263898f $X=9.745 $Y=1.53 $X2=0 $Y2=0
cc_393 N_S_c_437_n N_A0_c_651_n 0.0141724f $X=6.17 $Y=1.58 $X2=-0.19 $Y2=-0.24
cc_394 N_S_c_402_n N_A0_c_652_n 0.0399529f $X=6.475 $Y=1.41 $X2=0 $Y2=0
cc_395 N_S_c_437_n N_A0_c_652_n 0.0122397f $X=6.17 $Y=1.58 $X2=0 $Y2=0
cc_396 N_S_c_407_n N_A0_c_652_n 0.00190613f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_397 N_S_c_415_n N_A0_c_652_n 0.00153225f $X=6.4 $Y=1.53 $X2=0 $Y2=0
cc_398 N_S_c_414_n N_A0_c_644_n 0.00839646f $X=9.745 $Y=1.53 $X2=0 $Y2=0
cc_399 N_S_c_402_n N_A0_c_647_n 3.0536e-19 $X=6.475 $Y=1.41 $X2=0 $Y2=0
cc_400 N_S_c_403_n N_A0_c_647_n 0.0029333f $X=6.5 $Y=0.995 $X2=0 $Y2=0
cc_401 N_S_c_437_n N_A0_c_647_n 0.0140154f $X=6.17 $Y=1.58 $X2=0 $Y2=0
cc_402 N_S_c_407_n N_A0_c_647_n 0.0124522f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_403 N_S_c_402_n N_A0_c_672_n 0.00143275f $X=6.475 $Y=1.41 $X2=0 $Y2=0
cc_404 N_S_c_403_n N_A0_c_672_n 0.0135968f $X=6.5 $Y=0.995 $X2=0 $Y2=0
cc_405 N_S_c_414_n N_A0_c_649_n 0.00247602f $X=9.745 $Y=1.53 $X2=0 $Y2=0
cc_406 N_S_c_402_n N_A0_c_650_n 0.0259529f $X=6.475 $Y=1.41 $X2=0 $Y2=0
cc_407 N_S_c_437_n N_A0_c_650_n 0.00328398f $X=6.17 $Y=1.58 $X2=0 $Y2=0
cc_408 N_S_c_407_n N_A0_c_650_n 0.00579164f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_409 N_S_c_407_n N_A0_c_683_n 0.0253672f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_410 N_S_c_402_n N_A0_c_684_n 6.68847e-19 $X=6.475 $Y=1.41 $X2=0 $Y2=0
cc_411 N_S_c_408_n N_A_1369_199#_M1019_d 0.00576286f $X=10.15 $Y=1.16 $X2=0
+ $Y2=0
cc_412 N_S_c_402_n N_A_1369_199#_c_764_n 0.0569691f $X=6.475 $Y=1.41 $X2=0 $Y2=0
cc_413 N_S_c_441_n N_A_1369_199#_c_764_n 2.37626e-19 $X=6.377 $Y=1.495 $X2=0
+ $Y2=0
cc_414 N_S_c_407_n N_A_1369_199#_c_764_n 0.00178586f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_415 N_S_c_414_n N_A_1369_199#_c_764_n 0.00259714f $X=9.745 $Y=1.53 $X2=0
+ $Y2=0
cc_416 N_S_c_403_n N_A_1369_199#_c_765_n 0.0226554f $X=6.5 $Y=0.995 $X2=0 $Y2=0
cc_417 N_S_c_404_n N_A_1369_199#_c_766_n 0.0195231f $X=10.04 $Y=0.995 $X2=0
+ $Y2=0
cc_418 N_S_c_405_n N_A_1369_199#_c_767_n 0.0485577f $X=10.065 $Y=1.41 $X2=0
+ $Y2=0
cc_419 N_S_c_414_n N_A_1369_199#_c_767_n 0.00251865f $X=9.745 $Y=1.53 $X2=0
+ $Y2=0
cc_420 N_S_c_408_n N_A_1369_199#_c_767_n 0.00334991f $X=10.15 $Y=1.16 $X2=0
+ $Y2=0
cc_421 N_S_c_402_n N_A_1369_199#_c_768_n 0.00168674f $X=6.475 $Y=1.41 $X2=0
+ $Y2=0
cc_422 N_S_c_407_n N_A_1369_199#_c_768_n 0.0214562f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_423 N_S_c_414_n N_A_1369_199#_c_768_n 0.00590283f $X=9.745 $Y=1.53 $X2=0
+ $Y2=0
cc_424 N_S_c_415_n N_A_1369_199#_c_768_n 2.34085e-19 $X=6.4 $Y=1.53 $X2=0 $Y2=0
cc_425 N_S_c_414_n N_A_1369_199#_c_778_n 0.09431f $X=9.745 $Y=1.53 $X2=0 $Y2=0
cc_426 N_S_c_402_n N_A_1369_199#_c_781_n 2.40885e-19 $X=6.475 $Y=1.41 $X2=0
+ $Y2=0
cc_427 N_S_c_441_n N_A_1369_199#_c_781_n 0.00215289f $X=6.377 $Y=1.495 $X2=0
+ $Y2=0
cc_428 N_S_c_414_n N_A_1369_199#_c_781_n 0.00687607f $X=9.745 $Y=1.53 $X2=0
+ $Y2=0
cc_429 N_S_c_415_n N_A_1369_199#_c_781_n 2.67241e-19 $X=6.4 $Y=1.53 $X2=0 $Y2=0
cc_430 N_S_c_404_n N_A_1369_199#_c_769_n 0.00338504f $X=10.04 $Y=0.995 $X2=0
+ $Y2=0
cc_431 N_S_c_405_n N_A_1369_199#_c_769_n 6.76724e-19 $X=10.065 $Y=1.41 $X2=0
+ $Y2=0
cc_432 N_S_c_414_n N_A_1369_199#_c_769_n 0.0129437f $X=9.745 $Y=1.53 $X2=0 $Y2=0
cc_433 S N_A_1369_199#_c_769_n 0.00138473f $X=9.805 $Y=1.445 $X2=0 $Y2=0
cc_434 N_S_c_408_n N_A_1369_199#_c_769_n 0.0386674f $X=10.15 $Y=1.16 $X2=0 $Y2=0
cc_435 N_S_c_404_n N_A_1369_199#_c_806_n 0.0128687f $X=10.04 $Y=0.995 $X2=0
+ $Y2=0
cc_436 N_S_c_405_n N_A_1369_199#_c_806_n 0.00497414f $X=10.065 $Y=1.41 $X2=0
+ $Y2=0
cc_437 S N_A_1369_199#_c_806_n 0.00268678f $X=9.805 $Y=1.445 $X2=0 $Y2=0
cc_438 N_S_c_408_n N_A_1369_199#_c_806_n 0.0280671f $X=10.15 $Y=1.16 $X2=0 $Y2=0
cc_439 N_S_c_405_n N_A_1369_199#_c_810_n 0.0119825f $X=10.065 $Y=1.41 $X2=0
+ $Y2=0
cc_440 N_S_c_414_n N_A_1369_199#_c_810_n 0.00427154f $X=9.745 $Y=1.53 $X2=0
+ $Y2=0
cc_441 S N_A_1369_199#_c_810_n 0.00838822f $X=9.805 $Y=1.445 $X2=0 $Y2=0
cc_442 N_S_c_408_n N_A_1369_199#_c_810_n 0.0122662f $X=10.15 $Y=1.16 $X2=0 $Y2=0
cc_443 N_S_c_405_n N_A_1369_199#_c_814_n 0.0033249f $X=10.065 $Y=1.41 $X2=0
+ $Y2=0
cc_444 N_S_c_408_n N_A_1369_199#_c_814_n 0.00162807f $X=10.15 $Y=1.16 $X2=0
+ $Y2=0
cc_445 N_S_c_414_n N_A_1369_199#_c_816_n 0.014464f $X=9.745 $Y=1.53 $X2=0 $Y2=0
cc_446 S N_A_1369_199#_c_816_n 0.00226297f $X=9.805 $Y=1.445 $X2=0 $Y2=0
cc_447 N_S_c_408_n N_A_1369_199#_c_816_n 0.00617552f $X=10.15 $Y=1.16 $X2=0
+ $Y2=0
cc_448 N_S_c_414_n N_VPWR_M1033_s 0.00304429f $X=9.745 $Y=1.53 $X2=0 $Y2=0
cc_449 N_S_c_414_n N_VPWR_M1015_d 0.00101493f $X=9.745 $Y=1.53 $X2=0 $Y2=0
cc_450 S N_VPWR_M1015_d 0.00250029f $X=9.805 $Y=1.445 $X2=0 $Y2=0
cc_451 N_S_c_408_n N_VPWR_M1015_d 0.00149719f $X=10.15 $Y=1.16 $X2=0 $Y2=0
cc_452 N_S_c_402_n N_VPWR_c_895_n 0.00572314f $X=6.475 $Y=1.41 $X2=0 $Y2=0
cc_453 N_S_c_400_n N_VPWR_c_896_n 0.00480135f $X=4.26 $Y=1.41 $X2=0 $Y2=0
cc_454 N_S_c_402_n N_VPWR_c_896_n 0.00514401f $X=6.475 $Y=1.41 $X2=0 $Y2=0
cc_455 N_S_c_405_n N_VPWR_c_903_n 0.00311736f $X=10.065 $Y=1.41 $X2=0 $Y2=0
cc_456 N_S_c_400_n N_VPWR_c_889_n 0.00687434f $X=4.26 $Y=1.41 $X2=0 $Y2=0
cc_457 N_S_c_402_n N_VPWR_c_889_n 0.00708101f $X=6.475 $Y=1.41 $X2=0 $Y2=0
cc_458 N_S_c_405_n N_VPWR_c_889_n 0.00464062f $X=10.065 $Y=1.41 $X2=0 $Y2=0
cc_459 N_S_c_400_n N_VPWR_c_908_n 0.0103214f $X=4.26 $Y=1.41 $X2=0 $Y2=0
cc_460 N_S_c_405_n N_VPWR_c_909_n 0.0110499f $X=10.065 $Y=1.41 $X2=0 $Y2=0
cc_461 N_S_c_437_n N_A_870_297#_M1022_d 0.0313719f $X=6.17 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_462 N_S_c_437_n N_A_870_297#_M1012_d 4.70802e-19 $X=6.17 $Y=1.58 $X2=0 $Y2=0
cc_463 N_S_c_441_n N_A_870_297#_M1012_d 0.00174089f $X=6.377 $Y=1.495 $X2=0
+ $Y2=0
cc_464 N_S_c_400_n N_A_870_297#_c_1147_n 0.00361488f $X=4.26 $Y=1.41 $X2=0 $Y2=0
cc_465 N_S_c_402_n N_A_870_297#_c_1147_n 0.00270409f $X=6.475 $Y=1.41 $X2=0
+ $Y2=0
cc_466 N_S_c_403_n N_VGND_c_1181_n 0.00838946f $X=6.5 $Y=0.995 $X2=0 $Y2=0
cc_467 N_S_c_401_n N_VGND_c_1186_n 0.00423128f $X=4.285 $Y=0.995 $X2=0 $Y2=0
cc_468 N_S_c_403_n N_VGND_c_1186_n 0.00426565f $X=6.5 $Y=0.995 $X2=0 $Y2=0
cc_469 N_S_c_404_n N_VGND_c_1188_n 0.00199063f $X=10.04 $Y=0.995 $X2=0 $Y2=0
cc_470 N_S_c_401_n N_VGND_c_1189_n 0.00579723f $X=4.285 $Y=0.995 $X2=0 $Y2=0
cc_471 N_S_c_403_n N_VGND_c_1189_n 0.00725515f $X=6.5 $Y=0.995 $X2=0 $Y2=0
cc_472 N_S_c_404_n N_VGND_c_1189_n 0.00369877f $X=10.04 $Y=0.995 $X2=0 $Y2=0
cc_473 N_S_c_401_n N_VGND_c_1193_n 0.00315076f $X=4.285 $Y=0.995 $X2=0 $Y2=0
cc_474 N_S_c_404_n N_VGND_c_1195_n 0.0128194f $X=10.04 $Y=0.995 $X2=0 $Y2=0
cc_475 N_S_c_401_n N_A_872_47#_c_1334_n 0.00148617f $X=4.285 $Y=0.995 $X2=0
+ $Y2=0
cc_476 N_A1_c_550_n N_A0_c_644_n 8.79477e-19 $X=8.765 $Y=1.19 $X2=0 $Y2=0
cc_477 N_A1_c_550_n N_A0_c_645_n 0.00619051f $X=8.765 $Y=1.19 $X2=0 $Y2=0
cc_478 A1 N_A0_c_645_n 3.99038e-19 $X=8.885 $Y=1.105 $X2=0 $Y2=0
cc_479 N_A1_c_552_n N_A0_c_645_n 0.0248654f $X=9.045 $Y=1.202 $X2=0 $Y2=0
cc_480 N_A1_c_553_n N_A0_c_645_n 0.00157713f $X=8.97 $Y=1.19 $X2=0 $Y2=0
cc_481 N_A1_c_549_n N_A0_c_647_n 0.00352824f $X=5.15 $Y=0.96 $X2=0 $Y2=0
cc_482 N_A1_c_550_n N_A0_c_647_n 0.0150163f $X=8.765 $Y=1.19 $X2=0 $Y2=0
cc_483 N_A1_c_558_n N_A0_c_647_n 0.00495414f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_484 N_A1_c_550_n N_A0_c_672_n 0.00322056f $X=8.765 $Y=1.19 $X2=0 $Y2=0
cc_485 N_A1_c_549_n N_A0_c_677_n 0.0044939f $X=5.15 $Y=0.96 $X2=0 $Y2=0
cc_486 N_A1_c_550_n N_A0_c_649_n 0.0217372f $X=8.765 $Y=1.19 $X2=0 $Y2=0
cc_487 N_A1_c_552_n N_A0_c_649_n 0.00134463f $X=9.045 $Y=1.202 $X2=0 $Y2=0
cc_488 N_A1_c_549_n N_A0_c_650_n 0.0238871f $X=5.15 $Y=0.96 $X2=0 $Y2=0
cc_489 N_A1_c_550_n N_A0_c_650_n 0.0090165f $X=8.765 $Y=1.19 $X2=0 $Y2=0
cc_490 N_A1_c_551_n N_A0_c_650_n 4.08231e-19 $X=4.96 $Y=1.19 $X2=0 $Y2=0
cc_491 N_A1_c_558_n N_A0_c_650_n 9.59785e-19 $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_492 N_A1_c_550_n N_A0_c_683_n 0.00238349f $X=8.765 $Y=1.19 $X2=0 $Y2=0
cc_493 N_A1_c_550_n N_A_1369_199#_c_764_n 0.00301433f $X=8.765 $Y=1.19 $X2=0
+ $Y2=0
cc_494 N_A1_c_556_n N_A_1369_199#_c_767_n 0.0371628f $X=9.045 $Y=1.41 $X2=0
+ $Y2=0
cc_495 N_A1_c_552_n N_A_1369_199#_c_767_n 0.0240223f $X=9.045 $Y=1.202 $X2=0
+ $Y2=0
cc_496 N_A1_c_553_n N_A_1369_199#_c_767_n 0.00207545f $X=8.97 $Y=1.19 $X2=0
+ $Y2=0
cc_497 N_A1_c_550_n N_A_1369_199#_c_768_n 0.013453f $X=8.765 $Y=1.19 $X2=0 $Y2=0
cc_498 N_A1_c_555_n N_A_1369_199#_c_778_n 0.015572f $X=8.575 $Y=1.41 $X2=0 $Y2=0
cc_499 N_A1_c_556_n N_A_1369_199#_c_778_n 0.0129019f $X=9.045 $Y=1.41 $X2=0
+ $Y2=0
cc_500 N_A1_c_550_n N_A_1369_199#_c_778_n 0.00926239f $X=8.765 $Y=1.19 $X2=0
+ $Y2=0
cc_501 A1 N_A_1369_199#_c_778_n 0.00120239f $X=8.885 $Y=1.105 $X2=0 $Y2=0
cc_502 N_A1_c_552_n N_A_1369_199#_c_778_n 0.00487258f $X=9.045 $Y=1.202 $X2=0
+ $Y2=0
cc_503 N_A1_c_553_n N_A_1369_199#_c_778_n 0.0165311f $X=8.97 $Y=1.19 $X2=0 $Y2=0
cc_504 N_A1_c_556_n N_A_1369_199#_c_769_n 0.00137111f $X=9.045 $Y=1.41 $X2=0
+ $Y2=0
cc_505 A1 N_A_1369_199#_c_769_n 0.00134071f $X=8.885 $Y=1.105 $X2=0 $Y2=0
cc_506 N_A1_c_552_n N_A_1369_199#_c_769_n 0.00100599f $X=9.045 $Y=1.202 $X2=0
+ $Y2=0
cc_507 N_A1_c_553_n N_A_1369_199#_c_769_n 0.017533f $X=8.97 $Y=1.19 $X2=0 $Y2=0
cc_508 N_A1_c_555_n N_VPWR_c_902_n 0.00439333f $X=8.575 $Y=1.41 $X2=0 $Y2=0
cc_509 N_A1_c_556_n N_VPWR_c_902_n 0.00439333f $X=9.045 $Y=1.41 $X2=0 $Y2=0
cc_510 N_A1_c_555_n N_VPWR_c_889_n 0.00745558f $X=8.575 $Y=1.41 $X2=0 $Y2=0
cc_511 N_A1_c_556_n N_VPWR_c_889_n 0.00610813f $X=9.045 $Y=1.41 $X2=0 $Y2=0
cc_512 N_A1_c_555_n N_A_1420_297#_c_1163_n 0.0138826f $X=8.575 $Y=1.41 $X2=0
+ $Y2=0
cc_513 N_A1_c_556_n N_A_1420_297#_c_1163_n 0.0114f $X=9.045 $Y=1.41 $X2=0 $Y2=0
cc_514 N_A1_c_548_n N_VGND_c_1186_n 0.00366111f $X=4.73 $Y=0.96 $X2=0 $Y2=0
cc_515 N_A1_c_549_n N_VGND_c_1186_n 0.00366111f $X=5.15 $Y=0.96 $X2=0 $Y2=0
cc_516 N_A1_c_548_n N_VGND_c_1189_n 0.00532774f $X=4.73 $Y=0.96 $X2=0 $Y2=0
cc_517 N_A1_c_549_n N_VGND_c_1189_n 0.00647726f $X=5.15 $Y=0.96 $X2=0 $Y2=0
cc_518 N_A1_c_548_n N_A_872_47#_c_1334_n 0.00788636f $X=4.73 $Y=0.96 $X2=0 $Y2=0
cc_519 N_A1_c_549_n N_A_872_47#_c_1334_n 0.00783835f $X=5.15 $Y=0.96 $X2=0 $Y2=0
cc_520 N_A1_c_552_n N_A_1422_47#_c_1355_n 0.00254434f $X=9.045 $Y=1.202 $X2=0
+ $Y2=0
cc_521 N_A0_c_644_n N_A_1369_199#_c_764_n 0.0121015f $X=7.67 $Y=0.96 $X2=0 $Y2=0
cc_522 N_A0_c_672_n N_A_1369_199#_c_764_n 0.00558508f $X=7.325 $Y=0.73 $X2=0
+ $Y2=0
cc_523 N_A0_c_649_n N_A_1369_199#_c_764_n 0.0021752f $X=7.41 $Y=1.16 $X2=0 $Y2=0
cc_524 N_A0_c_644_n N_A_1369_199#_c_765_n 0.0206937f $X=7.67 $Y=0.96 $X2=0 $Y2=0
cc_525 N_A0_c_672_n N_A_1369_199#_c_765_n 0.0118644f $X=7.325 $Y=0.73 $X2=0
+ $Y2=0
cc_526 N_A0_c_648_n N_A_1369_199#_c_765_n 0.0032974f $X=7.41 $Y=0.995 $X2=0
+ $Y2=0
cc_527 N_A0_c_644_n N_A_1369_199#_c_768_n 7.22657e-19 $X=7.67 $Y=0.96 $X2=0
+ $Y2=0
cc_528 N_A0_c_672_n N_A_1369_199#_c_768_n 0.0125369f $X=7.325 $Y=0.73 $X2=0
+ $Y2=0
cc_529 N_A0_c_649_n N_A_1369_199#_c_768_n 0.0143594f $X=7.41 $Y=1.16 $X2=0 $Y2=0
cc_530 N_A0_c_644_n N_A_1369_199#_c_778_n 0.00270982f $X=7.67 $Y=0.96 $X2=0
+ $Y2=0
cc_531 N_A0_c_645_n N_A_1369_199#_c_778_n 0.0142315f $X=8.115 $Y=1.142 $X2=0
+ $Y2=0
cc_532 N_A0_c_649_n N_A_1369_199#_c_778_n 0.0248142f $X=7.41 $Y=1.16 $X2=0 $Y2=0
cc_533 N_A0_c_651_n N_VPWR_c_896_n 0.00439333f $X=5.535 $Y=1.41 $X2=0 $Y2=0
cc_534 N_A0_c_652_n N_VPWR_c_896_n 0.00439333f $X=6.005 $Y=1.41 $X2=0 $Y2=0
cc_535 N_A0_c_651_n N_VPWR_c_889_n 0.00745558f $X=5.535 $Y=1.41 $X2=0 $Y2=0
cc_536 N_A0_c_652_n N_VPWR_c_889_n 0.00610813f $X=6.005 $Y=1.41 $X2=0 $Y2=0
cc_537 N_A0_c_651_n N_A_870_297#_c_1147_n 0.0138826f $X=5.535 $Y=1.41 $X2=0
+ $Y2=0
cc_538 N_A0_c_652_n N_A_870_297#_c_1147_n 0.00977237f $X=6.005 $Y=1.41 $X2=0
+ $Y2=0
cc_539 N_A0_c_672_n N_VGND_M1023_d 0.00774541f $X=7.325 $Y=0.73 $X2=0 $Y2=0
cc_540 N_A0_c_644_n N_VGND_c_1181_n 0.00114889f $X=7.67 $Y=0.96 $X2=0 $Y2=0
cc_541 N_A0_c_672_n N_VGND_c_1181_n 0.0179073f $X=7.325 $Y=0.73 $X2=0 $Y2=0
cc_542 N_A0_c_672_n N_VGND_c_1186_n 0.00374524f $X=7.325 $Y=0.73 $X2=0 $Y2=0
cc_543 N_A0_c_677_n N_VGND_c_1186_n 0.00480391f $X=5.8 $Y=0.62 $X2=0 $Y2=0
cc_544 N_A0_c_683_n N_VGND_c_1186_n 0.0184623f $X=6.195 $Y=0.62 $X2=0 $Y2=0
cc_545 N_A0_c_644_n N_VGND_c_1187_n 0.00366111f $X=7.67 $Y=0.96 $X2=0 $Y2=0
cc_546 N_A0_c_646_n N_VGND_c_1187_n 0.00366111f $X=8.19 $Y=0.96 $X2=0 $Y2=0
cc_547 N_A0_c_672_n N_VGND_c_1187_n 0.00258949f $X=7.325 $Y=0.73 $X2=0 $Y2=0
cc_548 N_A0_c_644_n N_VGND_c_1189_n 0.00595908f $X=7.67 $Y=0.96 $X2=0 $Y2=0
cc_549 N_A0_c_646_n N_VGND_c_1189_n 0.0067042f $X=8.19 $Y=0.96 $X2=0 $Y2=0
cc_550 N_A0_c_672_n N_VGND_c_1189_n 0.00614972f $X=7.325 $Y=0.73 $X2=0 $Y2=0
cc_551 N_A0_c_677_n N_VGND_c_1189_n 0.00317366f $X=5.8 $Y=0.62 $X2=0 $Y2=0
cc_552 N_A0_c_683_n N_VGND_c_1189_n 0.00930158f $X=6.195 $Y=0.62 $X2=0 $Y2=0
cc_553 N_A0_c_647_n N_A_872_47#_M1005_s 0.00139381f $X=5.665 $Y=1.16 $X2=0 $Y2=0
cc_554 N_A0_c_677_n N_A_872_47#_M1005_s 0.011809f $X=5.8 $Y=0.62 $X2=0 $Y2=0
cc_555 N_A0_c_683_n N_A_872_47#_M1005_s 0.020124f $X=6.195 $Y=0.62 $X2=0 $Y2=0
cc_556 N_A0_c_684_n N_A_872_47#_M1005_s 0.00452131f $X=6.39 $Y=0.62 $X2=0 $Y2=0
cc_557 N_A0_c_677_n N_A_872_47#_c_1334_n 0.00279235f $X=5.8 $Y=0.62 $X2=0 $Y2=0
cc_558 N_A0_c_650_n N_A_872_47#_c_1334_n 0.00254434f $X=6.005 $Y=1.202 $X2=0
+ $Y2=0
cc_559 N_A0_c_672_n N_A_1422_47#_M1011_s 0.0096978f $X=7.325 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_560 N_A0_c_648_n N_A_1422_47#_M1011_s 0.00200006f $X=7.41 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_561 N_A0_c_644_n N_A_1422_47#_c_1355_n 0.0123986f $X=7.67 $Y=0.96 $X2=0 $Y2=0
cc_562 N_A0_c_646_n N_A_1422_47#_c_1355_n 0.00837958f $X=8.19 $Y=0.96 $X2=0
+ $Y2=0
cc_563 N_A0_c_672_n N_A_1422_47#_c_1355_n 0.0203831f $X=7.325 $Y=0.73 $X2=0
+ $Y2=0
cc_564 N_A0_c_649_n N_A_1422_47#_c_1355_n 0.00241368f $X=7.41 $Y=1.16 $X2=0
+ $Y2=0
cc_565 N_A_1369_199#_c_810_n N_VPWR_M1015_d 0.00602617f $X=10.215 $Y=2 $X2=0
+ $Y2=0
cc_566 N_A_1369_199#_c_764_n N_VPWR_c_895_n 0.00585347f $X=7.01 $Y=1.41 $X2=0
+ $Y2=0
cc_567 N_A_1369_199#_c_764_n N_VPWR_c_902_n 0.00490942f $X=7.01 $Y=1.41 $X2=0
+ $Y2=0
cc_568 N_A_1369_199#_c_767_n N_VPWR_c_902_n 0.00502091f $X=9.515 $Y=1.41 $X2=0
+ $Y2=0
cc_569 N_A_1369_199#_c_810_n N_VPWR_c_902_n 3.16703e-19 $X=10.215 $Y=2 $X2=0
+ $Y2=0
cc_570 N_A_1369_199#_c_851_p N_VPWR_c_902_n 0.00316861f $X=9.635 $Y=2 $X2=0
+ $Y2=0
cc_571 N_A_1369_199#_c_810_n N_VPWR_c_903_n 0.00238051f $X=10.215 $Y=2 $X2=0
+ $Y2=0
cc_572 N_A_1369_199#_c_853_p N_VPWR_c_903_n 0.011801f $X=10.3 $Y=2.3 $X2=0 $Y2=0
cc_573 N_A_1369_199#_M1019_d N_VPWR_c_889_n 0.00380573f $X=10.155 $Y=1.485 $X2=0
+ $Y2=0
cc_574 N_A_1369_199#_c_764_n N_VPWR_c_889_n 0.0080133f $X=7.01 $Y=1.41 $X2=0
+ $Y2=0
cc_575 N_A_1369_199#_c_767_n N_VPWR_c_889_n 0.0068565f $X=9.515 $Y=1.41 $X2=0
+ $Y2=0
cc_576 N_A_1369_199#_c_810_n N_VPWR_c_889_n 0.0067711f $X=10.215 $Y=2 $X2=0
+ $Y2=0
cc_577 N_A_1369_199#_c_851_p N_VPWR_c_889_n 0.00495396f $X=9.635 $Y=2 $X2=0
+ $Y2=0
cc_578 N_A_1369_199#_c_853_p N_VPWR_c_889_n 0.00646745f $X=10.3 $Y=2.3 $X2=0
+ $Y2=0
cc_579 N_A_1369_199#_c_767_n N_VPWR_c_909_n 0.00638092f $X=9.515 $Y=1.41 $X2=0
+ $Y2=0
cc_580 N_A_1369_199#_c_810_n N_VPWR_c_909_n 0.0236534f $X=10.215 $Y=2 $X2=0
+ $Y2=0
cc_581 N_A_1369_199#_c_853_p N_VPWR_c_909_n 0.0156776f $X=10.3 $Y=2.3 $X2=0
+ $Y2=0
cc_582 N_A_1369_199#_c_778_n N_A_1420_297#_M1013_s 0.0380172f $X=9.415 $Y=1.58
+ $X2=-0.19 $Y2=-0.24
cc_583 N_A_1369_199#_c_778_n N_A_1420_297#_M1024_d 0.00642019f $X=9.415 $Y=1.58
+ $X2=0 $Y2=0
cc_584 N_A_1369_199#_c_764_n N_A_1420_297#_c_1163_n 0.00430899f $X=7.01 $Y=1.41
+ $X2=0 $Y2=0
cc_585 N_A_1369_199#_c_767_n N_A_1420_297#_c_1163_n 0.00245323f $X=9.515 $Y=1.41
+ $X2=0 $Y2=0
cc_586 N_A_1369_199#_c_778_n N_A_1420_297#_c_1163_n 0.00891681f $X=9.415 $Y=1.58
+ $X2=0 $Y2=0
cc_587 N_A_1369_199#_c_851_p N_A_1420_297#_c_1163_n 0.00140438f $X=9.635 $Y=2
+ $X2=0 $Y2=0
cc_588 N_A_1369_199#_c_769_n N_VGND_M1025_d 8.04056e-19 $X=9.5 $Y=1.16 $X2=0
+ $Y2=0
cc_589 N_A_1369_199#_c_806_n N_VGND_M1025_d 0.00860919f $X=10.215 $Y=0.73 $X2=0
+ $Y2=0
cc_590 N_A_1369_199#_c_871_p N_VGND_M1025_d 2.40435e-19 $X=9.635 $Y=0.73 $X2=0
+ $Y2=0
cc_591 N_A_1369_199#_c_765_n N_VGND_c_1181_n 0.00859749f $X=7.035 $Y=0.995 $X2=0
+ $Y2=0
cc_592 N_A_1369_199#_c_765_n N_VGND_c_1187_n 0.00340533f $X=7.035 $Y=0.995 $X2=0
+ $Y2=0
cc_593 N_A_1369_199#_c_766_n N_VGND_c_1187_n 0.00426418f $X=9.49 $Y=0.995 $X2=0
+ $Y2=0
cc_594 N_A_1369_199#_c_806_n N_VGND_c_1187_n 5.06102e-19 $X=10.215 $Y=0.73 $X2=0
+ $Y2=0
cc_595 N_A_1369_199#_c_871_p N_VGND_c_1187_n 0.00342461f $X=9.635 $Y=0.73 $X2=0
+ $Y2=0
cc_596 N_A_1369_199#_c_806_n N_VGND_c_1188_n 0.00238481f $X=10.215 $Y=0.73 $X2=0
+ $Y2=0
cc_597 N_A_1369_199#_c_878_p N_VGND_c_1188_n 0.00921316f $X=10.3 $Y=0.46 $X2=0
+ $Y2=0
cc_598 N_A_1369_199#_M1032_d N_VGND_c_1189_n 0.00434565f $X=10.115 $Y=0.235
+ $X2=0 $Y2=0
cc_599 N_A_1369_199#_c_765_n N_VGND_c_1189_n 0.00426385f $X=7.035 $Y=0.995 $X2=0
+ $Y2=0
cc_600 N_A_1369_199#_c_766_n N_VGND_c_1189_n 0.00760146f $X=9.49 $Y=0.995 $X2=0
+ $Y2=0
cc_601 N_A_1369_199#_c_806_n N_VGND_c_1189_n 0.00698367f $X=10.215 $Y=0.73 $X2=0
+ $Y2=0
cc_602 N_A_1369_199#_c_871_p N_VGND_c_1189_n 0.00580088f $X=9.635 $Y=0.73 $X2=0
+ $Y2=0
cc_603 N_A_1369_199#_c_878_p N_VGND_c_1189_n 0.00629232f $X=10.3 $Y=0.46 $X2=0
+ $Y2=0
cc_604 N_A_1369_199#_c_766_n N_VGND_c_1195_n 0.00913205f $X=9.49 $Y=0.995 $X2=0
+ $Y2=0
cc_605 N_A_1369_199#_c_806_n N_VGND_c_1195_n 0.0229285f $X=10.215 $Y=0.73 $X2=0
+ $Y2=0
cc_606 N_A_1369_199#_c_878_p N_VGND_c_1195_n 0.0126914f $X=10.3 $Y=0.46 $X2=0
+ $Y2=0
cc_607 N_A_1369_199#_c_765_n N_A_1422_47#_c_1355_n 0.00179047f $X=7.035 $Y=0.995
+ $X2=0 $Y2=0
cc_608 N_VPWR_c_889_n N_X_M1000_s 0.00508986f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_609 N_VPWR_c_889_n N_X_M1004_s 0.00647849f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_610 N_VPWR_c_889_n N_X_M1014_s 0.00647849f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_611 N_VPWR_c_889_n N_X_M1021_s 0.00647849f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_612 N_VPWR_c_892_n N_X_c_1033_n 0.0417031f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_613 N_VPWR_c_898_n N_X_c_1033_n 0.0133725f $X=0.985 $Y=2.72 $X2=0 $Y2=0
cc_614 N_VPWR_c_889_n N_X_c_1033_n 0.00801045f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_615 N_VPWR_M1001_d N_X_c_1038_n 0.00385063f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_616 N_VPWR_c_892_n N_X_c_1038_n 0.0209383f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_617 N_VPWR_c_892_n N_X_c_1042_n 0.0336646f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_618 N_VPWR_c_893_n N_X_c_1042_n 0.0410603f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_619 N_VPWR_c_899_n N_X_c_1042_n 0.0118139f $X=1.925 $Y=2.72 $X2=0 $Y2=0
cc_620 N_VPWR_c_889_n N_X_c_1042_n 0.00646998f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_621 N_VPWR_M1008_d N_X_c_1048_n 0.00385063f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_622 N_VPWR_c_893_n N_X_c_1048_n 0.0209383f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_623 N_VPWR_c_893_n N_X_c_1053_n 0.0336646f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_624 N_VPWR_c_894_n N_X_c_1053_n 0.0410603f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_625 N_VPWR_c_900_n N_X_c_1053_n 0.0118139f $X=2.865 $Y=2.72 $X2=0 $Y2=0
cc_626 N_VPWR_c_889_n N_X_c_1053_n 0.00646998f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_627 N_VPWR_M1018_d N_X_c_1061_n 0.00385063f $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_628 N_VPWR_c_894_n N_X_c_1061_n 0.0209383f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_629 N_VPWR_c_894_n N_X_c_1067_n 0.0336646f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_630 N_VPWR_c_901_n N_X_c_1067_n 0.0118139f $X=3.805 $Y=2.72 $X2=0 $Y2=0
cc_631 N_VPWR_c_889_n N_X_c_1067_n 0.00646998f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_632 N_VPWR_c_908_n N_X_c_1067_n 0.0156776f $X=4.02 $Y=2.34 $X2=0 $Y2=0
cc_633 N_VPWR_c_889_n N_A_870_297#_M1022_d 0.01034f $X=10.35 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_634 N_VPWR_c_889_n N_A_870_297#_M1012_d 0.00233855f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_635 N_VPWR_c_895_n N_A_870_297#_c_1147_n 0.00923188f $X=6.76 $Y=2.34 $X2=0
+ $Y2=0
cc_636 N_VPWR_c_896_n N_A_870_297#_c_1147_n 0.0828059f $X=6.675 $Y=2.72 $X2=0
+ $Y2=0
cc_637 N_VPWR_c_889_n N_A_870_297#_c_1147_n 0.0625997f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_638 N_VPWR_c_908_n N_A_870_297#_c_1147_n 0.00665437f $X=4.02 $Y=2.34 $X2=0
+ $Y2=0
cc_639 N_VPWR_c_889_n N_A_1420_297#_M1013_s 0.0114104f $X=10.35 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_640 N_VPWR_c_889_n N_A_1420_297#_M1024_d 0.00233855f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_641 N_VPWR_c_895_n N_A_1420_297#_c_1163_n 0.0123628f $X=6.76 $Y=2.34 $X2=0
+ $Y2=0
cc_642 N_VPWR_c_902_n N_A_1420_297#_c_1163_n 0.113775f $X=9.665 $Y=2.72 $X2=0
+ $Y2=0
cc_643 N_VPWR_c_889_n N_A_1420_297#_c_1163_n 0.0854635f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_644 N_VPWR_c_909_n N_A_1420_297#_c_1163_n 0.0114572f $X=9.83 $Y=2.34 $X2=0
+ $Y2=0
cc_645 N_X_c_1034_n N_VGND_M1009_s 0.00472004f $X=1.585 $Y=0.72 $X2=0 $Y2=0
cc_646 N_X_c_1044_n N_VGND_M1020_s 0.00439476f $X=2.525 $Y=0.72 $X2=0 $Y2=0
cc_647 N_X_c_1055_n N_VGND_M1027_s 0.00439476f $X=3.465 $Y=0.72 $X2=0 $Y2=0
cc_648 N_X_c_1032_n N_VGND_c_1180_n 0.0150877f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_649 N_X_c_1032_n N_VGND_c_1182_n 0.0144177f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_650 N_X_c_1034_n N_VGND_c_1182_n 0.00195705f $X=1.585 $Y=0.72 $X2=0 $Y2=0
cc_651 N_X_c_1034_n N_VGND_c_1183_n 0.00325972f $X=1.585 $Y=0.72 $X2=0 $Y2=0
cc_652 N_X_c_1119_p N_VGND_c_1183_n 0.00904465f $X=1.67 $Y=0.46 $X2=0 $Y2=0
cc_653 N_X_c_1044_n N_VGND_c_1183_n 0.00244629f $X=2.525 $Y=0.72 $X2=0 $Y2=0
cc_654 N_X_c_1044_n N_VGND_c_1184_n 0.0032663f $X=2.525 $Y=0.72 $X2=0 $Y2=0
cc_655 N_X_c_1052_n N_VGND_c_1184_n 0.01143f $X=2.61 $Y=0.42 $X2=0 $Y2=0
cc_656 N_X_c_1055_n N_VGND_c_1184_n 0.00245287f $X=3.465 $Y=0.72 $X2=0 $Y2=0
cc_657 N_X_c_1055_n N_VGND_c_1185_n 0.00325972f $X=3.465 $Y=0.72 $X2=0 $Y2=0
cc_658 N_X_c_1125_p N_VGND_c_1185_n 0.00920056f $X=3.55 $Y=0.46 $X2=0 $Y2=0
cc_659 N_X_M1006_d N_VGND_c_1189_n 0.00480647f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_660 N_X_M1010_d N_VGND_c_1189_n 0.0031153f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_661 N_X_M1026_d N_VGND_c_1189_n 0.00307738f $X=2.425 $Y=0.235 $X2=0 $Y2=0
cc_662 N_X_M1029_d N_VGND_c_1189_n 0.00687576f $X=3.365 $Y=0.235 $X2=0 $Y2=0
cc_663 N_X_c_1032_n N_VGND_c_1189_n 0.00801045f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_664 N_X_c_1034_n N_VGND_c_1189_n 0.01012f $X=1.585 $Y=0.72 $X2=0 $Y2=0
cc_665 N_X_c_1119_p N_VGND_c_1189_n 0.00628881f $X=1.67 $Y=0.46 $X2=0 $Y2=0
cc_666 N_X_c_1044_n N_VGND_c_1189_n 0.0115126f $X=2.525 $Y=0.72 $X2=0 $Y2=0
cc_667 N_X_c_1052_n N_VGND_c_1189_n 0.00643448f $X=2.61 $Y=0.42 $X2=0 $Y2=0
cc_668 N_X_c_1055_n N_VGND_c_1189_n 0.0115126f $X=3.465 $Y=0.72 $X2=0 $Y2=0
cc_669 N_X_c_1125_p N_VGND_c_1189_n 0.00628881f $X=3.55 $Y=0.46 $X2=0 $Y2=0
cc_670 N_X_c_1071_n N_VGND_c_1189_n 0.00148162f $X=0.735 $Y=0.72 $X2=0 $Y2=0
cc_671 N_X_c_1034_n N_VGND_c_1190_n 0.0197774f $X=1.585 $Y=0.72 $X2=0 $Y2=0
cc_672 N_X_c_1119_p N_VGND_c_1190_n 0.0104056f $X=1.67 $Y=0.46 $X2=0 $Y2=0
cc_673 N_X_c_1044_n N_VGND_c_1191_n 0.0197774f $X=2.525 $Y=0.72 $X2=0 $Y2=0
cc_674 N_X_c_1052_n N_VGND_c_1191_n 0.0128539f $X=2.61 $Y=0.42 $X2=0 $Y2=0
cc_675 N_X_c_1055_n N_VGND_c_1192_n 0.0197774f $X=3.465 $Y=0.72 $X2=0 $Y2=0
cc_676 N_X_c_1125_p N_VGND_c_1192_n 0.0104056f $X=3.55 $Y=0.46 $X2=0 $Y2=0
cc_677 N_X_c_1125_p N_VGND_c_1193_n 0.0126914f $X=3.55 $Y=0.46 $X2=0 $Y2=0
cc_678 N_VGND_c_1189_n N_A_872_47#_M1007_s 0.00237915f $X=10.35 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_679 N_VGND_c_1189_n N_A_872_47#_M1005_s 0.00934106f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_680 N_VGND_c_1186_n N_A_872_47#_c_1334_n 0.0523253f $X=6.66 $Y=0 $X2=0 $Y2=0
cc_681 N_VGND_c_1189_n N_A_872_47#_c_1334_n 0.032796f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_682 N_VGND_c_1189_n N_A_1422_47#_M1011_s 0.00339599f $X=10.35 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_683 N_VGND_c_1189_n N_A_1422_47#_M1031_s 0.0386173f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_684 N_VGND_c_1181_n N_A_1422_47#_c_1355_n 0.012994f $X=6.825 $Y=0.38 $X2=0
+ $Y2=0
cc_685 N_VGND_c_1187_n N_A_1422_47#_c_1355_n 0.0647469f $X=9.665 $Y=0 $X2=0
+ $Y2=0
cc_686 N_VGND_c_1189_n N_A_1422_47#_c_1355_n 0.0247721f $X=10.35 $Y=0 $X2=0
+ $Y2=0
