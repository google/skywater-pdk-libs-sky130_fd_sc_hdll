* File: sky130_fd_sc_hdll__and2_6.pex.spice
* Created: Thu Aug 27 18:57:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND2_6%B 1 3 4 6 7 9 10 12 13 14 15 16 18 19 24 28
c81 18 0 1.22108e-19 $X=1.795 $Y=1.465
c82 15 0 1.48863e-19 $X=1.705 $Y=1.55
c83 10 0 1.60887e-19 $X=1.905 $Y=1.41
c84 7 0 7.31881e-20 $X=1.82 $Y=0.995
r85 24 27 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=1.16
+ $X2=1.835 $Y2=1.325
r86 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.16 $X2=1.88 $Y2=1.16
r87 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.49
+ $Y=1.16 $X2=0.49 $Y2=1.16
r88 19 28 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.435 $Y=1.16
+ $X2=0.23 $Y2=1.16
r89 19 21 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=0.435 $Y=1.16 $X2=0.525
+ $Y2=1.16
r90 18 27 8.62626 $w=1.78e-07 $l=1.4e-07 $layer=LI1_cond $X=1.795 $Y=1.465
+ $X2=1.795 $Y2=1.325
r91 15 18 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.705 $Y=1.55
+ $X2=1.795 $Y2=1.465
r92 15 16 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=1.705 $Y=1.55
+ $X2=0.615 $Y2=1.55
r93 14 16 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.525 $Y=1.465
+ $X2=0.615 $Y2=1.55
r94 13 21 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=1.325
+ $X2=0.525 $Y2=1.16
r95 13 14 8.62626 $w=1.78e-07 $l=1.4e-07 $layer=LI1_cond $X=0.525 $Y=1.325
+ $X2=0.525 $Y2=1.465
r96 10 25 49.2447 $w=2.79e-07 $l=2.54951e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.895 $Y2=1.16
r97 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r98 7 25 38.7444 $w=2.79e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.82 $Y=0.995
+ $X2=1.895 $Y2=1.16
r99 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.82 $Y=0.995 $X2=1.82
+ $Y2=0.56
r100 4 22 38.5416 $w=3.03e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.58 $Y=0.995
+ $X2=0.49 $Y2=1.16
r101 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.58 $Y=0.995
+ $X2=0.58 $Y2=0.56
r102 1 22 47.6478 $w=3.03e-07 $l=2.52488e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.49 $Y2=1.16
r103 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_6%A 1 3 4 6 7 9 10 12 13 19 20
r48 20 21 5.70789 $w=3.8e-07 $l=4.5e-08 $layer=POLY_cond $X=1.39 $Y=1.202
+ $X2=1.435 $Y2=1.202
r49 18 20 2.53684 $w=3.8e-07 $l=2e-08 $layer=POLY_cond $X=1.37 $Y=1.202 $X2=1.39
+ $Y2=1.202
r50 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.37
+ $Y=1.16 $X2=1.37 $Y2=1.16
r51 16 18 50.7368 $w=3.8e-07 $l=4e-07 $layer=POLY_cond $X=0.97 $Y=1.202 $X2=1.37
+ $Y2=1.202
r52 15 16 0.634211 $w=3.8e-07 $l=5e-09 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.97 $Y2=1.202
r53 13 19 8.45125 $w=2.98e-07 $l=2.2e-07 $layer=LI1_cond $X=1.15 $Y=1.145
+ $X2=1.37 $Y2=1.145
r54 10 21 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r55 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r56 7 20 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.39 $Y=0.995
+ $X2=1.39 $Y2=1.202
r57 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.39 $Y=0.995 $X2=1.39
+ $Y2=0.56
r58 4 16 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.97 $Y=0.995
+ $X2=0.97 $Y2=1.202
r59 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.97 $Y=0.995 $X2=0.97
+ $Y2=0.56
r60 1 15 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r61 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_6%A_117_297# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 39 40 42 43 45 48 52 54 55 58 61 63 69 73 75 76
+ 89
c165 89 0 7.45138e-20 $X=4.7 $Y=1.202
c166 75 0 1.60887e-19 $X=1.67 $Y=1.96
c167 10 0 1.96457e-19 $X=2.375 $Y=1.41
r168 89 90 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=4.7 $Y=1.202
+ $X2=4.725 $Y2=1.202
r169 88 89 54.7135 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.28 $Y=1.202
+ $X2=4.7 $Y2=1.202
r170 87 88 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=4.255 $Y=1.202
+ $X2=4.28 $Y2=1.202
r171 84 85 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=3.76 $Y=1.202
+ $X2=3.785 $Y2=1.202
r172 83 84 54.7135 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.34 $Y=1.202
+ $X2=3.76 $Y2=1.202
r173 82 83 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=3.315 $Y=1.202
+ $X2=3.34 $Y2=1.202
r174 81 82 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=3.315 $Y2=1.202
r175 80 81 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.845 $Y2=1.202
r176 77 78 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.4 $Y2=1.202
r177 70 87 14.9811 $w=3.7e-07 $l=1.15e-07 $layer=POLY_cond $X=4.14 $Y=1.202
+ $X2=4.255 $Y2=1.202
r178 70 85 46.2459 $w=3.7e-07 $l=3.55e-07 $layer=POLY_cond $X=4.14 $Y=1.202
+ $X2=3.785 $Y2=1.202
r179 69 70 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=4.14
+ $Y=1.16 $X2=4.14 $Y2=1.16
r180 67 80 49.5027 $w=3.7e-07 $l=3.8e-07 $layer=POLY_cond $X=2.44 $Y=1.202
+ $X2=2.82 $Y2=1.202
r181 67 78 5.21081 $w=3.7e-07 $l=4e-08 $layer=POLY_cond $X=2.44 $Y=1.202 $X2=2.4
+ $Y2=1.202
r182 66 69 89.7835 $w=2.08e-07 $l=1.7e-06 $layer=LI1_cond $X=2.44 $Y=1.16
+ $X2=4.14 $Y2=1.16
r183 66 67 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=2.44
+ $Y=1.16 $X2=2.44 $Y2=1.16
r184 64 76 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=1.16
+ $X2=2.22 $Y2=1.16
r185 64 66 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=2.305 $Y=1.16
+ $X2=2.44 $Y2=1.16
r186 62 76 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.22 $Y=1.265
+ $X2=2.22 $Y2=1.16
r187 62 63 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.22 $Y=1.265
+ $X2=2.22 $Y2=1.805
r188 61 76 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.22 $Y=1.055
+ $X2=2.22 $Y2=1.16
r189 60 61 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.22 $Y=0.825
+ $X2=2.22 $Y2=1.055
r190 59 75 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.805 $Y=1.89
+ $X2=1.67 $Y2=1.89
r191 58 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.135 $Y=1.89
+ $X2=2.22 $Y2=1.805
r192 58 59 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.135 $Y=1.89
+ $X2=1.805 $Y2=1.89
r193 54 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.135 $Y=0.74
+ $X2=2.22 $Y2=0.825
r194 54 55 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=2.135 $Y=0.74
+ $X2=1.345 $Y2=0.74
r195 50 55 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.18 $Y=0.655
+ $X2=1.345 $Y2=0.74
r196 50 52 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.18 $Y=0.655
+ $X2=1.18 $Y2=0.38
r197 49 73 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.865 $Y=1.89
+ $X2=0.715 $Y2=1.89
r198 48 75 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.535 $Y=1.89
+ $X2=1.67 $Y2=1.89
r199 48 49 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.535 $Y=1.89
+ $X2=0.865 $Y2=1.89
r200 43 90 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.202
r201 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.985
r202 40 89 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.7 $Y=0.995
+ $X2=4.7 $Y2=1.202
r203 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.7 $Y=0.995
+ $X2=4.7 $Y2=0.56
r204 37 88 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.28 $Y=0.995
+ $X2=4.28 $Y2=1.202
r205 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.28 $Y=0.995
+ $X2=4.28 $Y2=0.56
r206 34 87 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.202
r207 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.985
r208 31 85 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.202
r209 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r210 28 84 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.76 $Y=0.995
+ $X2=3.76 $Y2=1.202
r211 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.76 $Y=0.995
+ $X2=3.76 $Y2=0.56
r212 25 83 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.34 $Y=0.995
+ $X2=3.34 $Y2=1.202
r213 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.34 $Y=0.995
+ $X2=3.34 $Y2=0.56
r214 22 82 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.202
r215 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r216 19 81 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r217 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r218 16 80 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=1.202
r219 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=0.56
r220 13 78 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.4 $Y=0.995
+ $X2=2.4 $Y2=1.202
r221 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.4 $Y=0.995
+ $X2=2.4 $Y2=0.56
r222 10 77 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r223 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r224 3 75 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.96
r225 2 73 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.96
r226 1 52 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.045
+ $Y=0.235 $X2=1.18 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_6%VPWR 1 2 3 4 5 6 19 21 25 29 31 35 37 41 43
+ 47 49 51 56 63 64 70 73 76 79 82
r92 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r93 80 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r94 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r95 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r96 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r97 74 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r98 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r99 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r100 64 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r101 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r102 61 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=2.72
+ $X2=4.96 $Y2=2.72
r103 61 63 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=2.72
+ $X2=5.29 $Y2=2.72
r104 60 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r105 60 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r106 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r107 57 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.2 $Y2=2.72
r108 57 59 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.61 $Y2=2.72
r109 56 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=2.72
+ $X2=2.14 $Y2=2.72
r110 56 59 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.975 $Y=2.72
+ $X2=1.61 $Y2=2.72
r111 55 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r112 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r113 52 67 4.49698 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r114 52 54 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.69 $Y2=2.72
r115 51 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=1.2 $Y2=2.72
r116 51 54 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=0.69 $Y2=2.72
r117 49 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r118 49 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r119 45 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=2.72
r120 45 47 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=1.89
r121 44 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=2.72
+ $X2=4.02 $Y2=2.72
r122 43 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=2.72
+ $X2=4.96 $Y2=2.72
r123 43 44 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.795 $Y=2.72
+ $X2=4.185 $Y2=2.72
r124 39 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=2.72
r125 39 41 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=1.89
r126 38 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=2.72
+ $X2=3.08 $Y2=2.72
r127 37 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=2.72
+ $X2=4.02 $Y2=2.72
r128 37 38 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.855 $Y=2.72
+ $X2=3.245 $Y2=2.72
r129 33 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2.72
r130 33 35 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=1.89
r131 32 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=2.72
+ $X2=2.14 $Y2=2.72
r132 31 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=3.08 $Y2=2.72
r133 31 32 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=2.305 $Y2=2.72
r134 27 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.72
r135 27 29 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.245
r136 23 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.72
r137 23 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.34
r138 19 67 3.0207 $w=3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.197 $Y2=2.72
r139 19 21 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.245 $Y2=2
r140 6 47 300 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=1.89
r141 5 41 300 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=1.89
r142 4 35 300 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=1.89
r143 3 29 600 $w=1.7e-07 $l=8.29337e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2.245
r144 2 25 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.34
r145 1 21 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_6%X 1 2 3 4 5 6 21 25 29 30 31 32 35 39 43 45
+ 49 53 57 58 60 62 63
c85 30 0 7.31881e-20 $X=2.745 $Y=0.8
r86 61 63 6.1 $w=4.98e-07 $l=2.55e-07 $layer=LI1_cond $X=4.725 $Y=1.445
+ $X2=4.725 $Y2=1.19
r87 61 62 2.50573 $w=3.85e-07 $l=1.11018e-07 $layer=LI1_cond $X=4.725 $Y=1.445
+ $X2=4.665 $Y2=1.53
r88 59 63 7.29608 $w=4.98e-07 $l=3.05e-07 $layer=LI1_cond $X=4.725 $Y=0.885
+ $X2=4.725 $Y2=1.19
r89 59 60 2.50573 $w=3.85e-07 $l=1.11018e-07 $layer=LI1_cond $X=4.725 $Y=0.885
+ $X2=4.665 $Y2=0.8
r90 53 55 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.49 $Y=1.62
+ $X2=4.49 $Y2=2.3
r91 51 62 2.50573 $w=3.85e-07 $l=2.13307e-07 $layer=LI1_cond $X=4.49 $Y=1.615
+ $X2=4.665 $Y2=1.53
r92 51 53 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=4.49 $Y=1.615
+ $X2=4.49 $Y2=1.62
r93 47 60 2.50573 $w=3.85e-07 $l=2.13307e-07 $layer=LI1_cond $X=4.49 $Y=0.715
+ $X2=4.665 $Y2=0.8
r94 47 49 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.49 $Y=0.715
+ $X2=4.49 $Y2=0.42
r95 46 58 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.685 $Y=1.53
+ $X2=3.55 $Y2=1.53
r96 45 62 4.39717 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=4.355 $Y=1.53
+ $X2=4.665 $Y2=1.53
r97 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.355 $Y=1.53
+ $X2=3.685 $Y2=1.53
r98 44 57 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.685 $Y=0.8
+ $X2=3.55 $Y2=0.8
r99 43 60 4.39717 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=4.355 $Y=0.8
+ $X2=4.665 $Y2=0.8
r100 43 44 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.355 $Y=0.8
+ $X2=3.685 $Y2=0.8
r101 39 41 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.55 $Y=1.62
+ $X2=3.55 $Y2=2.3
r102 37 58 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=1.615
+ $X2=3.55 $Y2=1.53
r103 37 39 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=3.55 $Y=1.615
+ $X2=3.55 $Y2=1.62
r104 33 57 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=0.715
+ $X2=3.55 $Y2=0.8
r105 33 35 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.55 $Y=0.715
+ $X2=3.55 $Y2=0.42
r106 31 58 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.415 $Y=1.53
+ $X2=3.55 $Y2=1.53
r107 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.415 $Y=1.53
+ $X2=2.745 $Y2=1.53
r108 29 57 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.415 $Y=0.8
+ $X2=3.55 $Y2=0.8
r109 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.415 $Y=0.8
+ $X2=2.745 $Y2=0.8
r110 25 27 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.61 $Y=1.62
+ $X2=2.61 $Y2=2.3
r111 23 32 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.61 $Y=1.615
+ $X2=2.745 $Y2=1.53
r112 23 25 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=2.61 $Y=1.615
+ $X2=2.61 $Y2=1.62
r113 19 30 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.61 $Y=0.715
+ $X2=2.745 $Y2=0.8
r114 19 21 6.61588 $w=2.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.61 $Y=0.715
+ $X2=2.61 $Y2=0.56
r115 6 55 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=2.3
r116 6 53 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=1.62
r117 5 41 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2.3
r118 5 39 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.62
r119 4 27 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.3
r120 4 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.62
r121 3 49 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=4.355
+ $Y=0.235 $X2=4.49 $Y2=0.42
r122 2 35 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=3.415
+ $Y=0.235 $X2=3.55 $Y2=0.42
r123 1 21 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=2.61 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_6%VGND 1 2 3 4 5 16 18 22 24 28 30 34 36 40
+ 42 44 54 55 61 64 67 70
r81 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r82 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r83 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r84 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r85 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r86 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r87 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r88 55 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r89 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r90 52 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=0 $X2=4.96
+ $Y2=0
r91 52 54 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=0 $X2=5.29
+ $Y2=0
r92 51 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r93 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r94 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r95 47 50 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r96 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r97 45 58 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r98 45 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r99 44 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=2.105
+ $Y2=0
r100 44 50 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=1.61
+ $Y2=0
r101 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r102 42 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r103 38 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0
r104 38 40 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0.44
r105 37 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=0 $X2=4.02
+ $Y2=0
r106 36 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=4.96
+ $Y2=0
r107 36 37 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.795 $Y=0
+ $X2=4.185 $Y2=0
r108 32 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0
r109 32 34 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0.44
r110 31 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=0 $X2=3.08
+ $Y2=0
r111 30 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=0 $X2=4.02
+ $Y2=0
r112 30 31 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.855 $Y=0
+ $X2=3.245 $Y2=0
r113 26 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0
r114 26 28 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.44
r115 25 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.105
+ $Y2=0
r116 24 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=3.08
+ $Y2=0
r117 24 25 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=2.915 $Y=0
+ $X2=2.27 $Y2=0
r118 20 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0
r119 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0.36
r120 16 58 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r121 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r122 5 40 182 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.235 $X2=4.96 $Y2=0.44
r123 4 34 182 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_NDIFF $count=1 $X=3.835
+ $Y=0.235 $X2=4.02 $Y2=0.44
r124 3 28 182 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.44
r125 2 22 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.235 $X2=2.105 $Y2=0.36
r126 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

