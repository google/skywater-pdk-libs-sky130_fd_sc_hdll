* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__inputiso1p_1 A SLEEP VGND VNB VPB VPWR X
M1000 a_44_297# A VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=3.517e+11p ps=3.53e+06u
M1001 VPWR SLEEP a_134_297# VPB phighvt w=420000u l=180000u
+  ad=3.057e+11p pd=2.71e+06u as=1.218e+11p ps=1.42e+06u
M1002 X a_44_297# VGND VNB nshort w=650000u l=150000u
+  ad=2.405e+11p pd=2.04e+06u as=0p ps=0u
M1003 VGND SLEEP a_44_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_134_297# A a_44_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1005 X a_44_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=4.1e+11p pd=2.82e+06u as=0p ps=0u
.ends
