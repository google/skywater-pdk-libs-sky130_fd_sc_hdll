* File: sky130_fd_sc_hdll__a22oi_4.pex.spice
* Created: Wed Sep  2 08:19:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A22OI_4%B2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39 44
c83 19 0 1.70485e-19 $X=1.905 $Y=1.41
r84 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=1.93 $Y2=1.202
r85 37 39 14.9005 $w=3.72e-07 $l=1.15e-07 $layer=POLY_cond $X=1.79 $Y=1.202
+ $X2=1.905 $Y2=1.202
r86 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.79
+ $Y=1.16 $X2=1.79 $Y2=1.16
r87 35 37 45.9973 $w=3.72e-07 $l=3.55e-07 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.79 $Y2=1.202
r88 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.202
+ $X2=1.435 $Y2=1.202
r89 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=1.41 $Y2=1.202
r90 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.202
+ $X2=0.965 $Y2=1.202
r91 31 44 29.6682 $w=1.98e-07 $l=5.35e-07 $layer=LI1_cond $X=0.62 $Y=1.175
+ $X2=1.155 $Y2=1.175
r92 30 32 41.4624 $w=3.72e-07 $l=3.2e-07 $layer=POLY_cond $X=0.62 $Y=1.202
+ $X2=0.94 $Y2=1.202
r93 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.62
+ $Y=1.16 $X2=0.62 $Y2=1.16
r94 28 30 16.1962 $w=3.72e-07 $l=1.25e-07 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.62 $Y2=1.202
r95 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r96 25 38 34.3818 $w=1.98e-07 $l=6.2e-07 $layer=LI1_cond $X=1.17 $Y=1.175
+ $X2=1.79 $Y2=1.175
r97 25 44 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=1.17 $Y=1.175
+ $X2=1.155 $Y2=1.175
r98 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r99 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r100 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r101 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r102 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r103 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r104 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.202
r105 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=0.56
r106 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r107 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r108 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=1.202
r109 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=0.56
r110 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r111 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r112 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.202
r113 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_4%B1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 37 40 42
c70 1 0 1.56657e-19 $X=2.35 $Y=0.995
r71 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.845
+ $Y=1.16 $X2=3.845 $Y2=1.16
r72 37 39 7.8587 $w=3.68e-07 $l=6e-08 $layer=POLY_cond $X=3.785 $Y=1.202
+ $X2=3.845 $Y2=1.202
r73 36 37 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=3.76 $Y=1.202
+ $X2=3.785 $Y2=1.202
r74 35 36 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=3.315 $Y=1.202
+ $X2=3.76 $Y2=1.202
r75 34 35 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.202
+ $X2=3.315 $Y2=1.202
r76 33 42 6.65455 $w=1.98e-07 $l=1.2e-07 $layer=LI1_cond $X=3.115 $Y=1.175
+ $X2=2.995 $Y2=1.175
r77 32 34 22.9212 $w=3.68e-07 $l=1.75e-07 $layer=POLY_cond $X=3.115 $Y=1.202
+ $X2=3.29 $Y2=1.202
r78 32 33 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.115
+ $Y=1.16 $X2=3.115 $Y2=1.16
r79 30 32 35.3641 $w=3.68e-07 $l=2.7e-07 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=3.115 $Y2=1.202
r80 29 30 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.845 $Y2=1.202
r81 28 29 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.82 $Y2=1.202
r82 27 28 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.202
+ $X2=2.375 $Y2=1.202
r83 25 40 21.9045 $w=1.98e-07 $l=3.95e-07 $layer=LI1_cond $X=3.45 $Y=1.175
+ $X2=3.845 $Y2=1.175
r84 25 33 18.5773 $w=1.98e-07 $l=3.35e-07 $layer=LI1_cond $X=3.45 $Y=1.175
+ $X2=3.115 $Y2=1.175
r85 22 37 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.202
r86 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r87 19 36 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.76 $Y=0.995
+ $X2=3.76 $Y2=1.202
r88 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.76 $Y=0.995
+ $X2=3.76 $Y2=0.56
r89 16 35 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.202
r90 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r91 13 34 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=1.202
r92 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=0.56
r93 10 30 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r94 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r95 7 29 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=1.202
r96 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.82 $Y=0.995 $X2=2.82
+ $Y2=0.56
r97 4 28 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r98 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r99 1 27 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.202
r100 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_4%A1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39 43
r62 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.185 $Y=1.202
+ $X2=6.21 $Y2=1.202
r63 37 39 22.6747 $w=3.72e-07 $l=1.75e-07 $layer=POLY_cond $X=6.01 $Y=1.202
+ $X2=6.185 $Y2=1.202
r64 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.01
+ $Y=1.16 $X2=6.01 $Y2=1.16
r65 35 37 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=5.715 $Y=1.202
+ $X2=6.01 $Y2=1.202
r66 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.69 $Y=1.202
+ $X2=5.715 $Y2=1.202
r67 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=5.245 $Y=1.202
+ $X2=5.69 $Y2=1.202
r68 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.22 $Y=1.202
+ $X2=5.245 $Y2=1.202
r69 30 32 49.2366 $w=3.72e-07 $l=3.8e-07 $layer=POLY_cond $X=4.84 $Y=1.202
+ $X2=5.22 $Y2=1.202
r70 30 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.84
+ $Y=1.16 $X2=4.84 $Y2=1.16
r71 28 30 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=4.775 $Y=1.202
+ $X2=4.84 $Y2=1.202
r72 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.75 $Y=1.202
+ $X2=4.775 $Y2=1.202
r73 25 38 37.2338 $w=2.08e-07 $l=7.05e-07 $layer=LI1_cond $X=5.305 $Y=1.18
+ $X2=6.01 $Y2=1.18
r74 25 43 24.5584 $w=2.08e-07 $l=4.65e-07 $layer=LI1_cond $X=5.305 $Y=1.18
+ $X2=4.84 $Y2=1.18
r75 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.21 $Y=0.995
+ $X2=6.21 $Y2=1.202
r76 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.21 $Y=0.995
+ $X2=6.21 $Y2=0.56
r77 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.202
r78 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.985
r79 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.202
r80 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.985
r81 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=1.202
r82 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=0.56
r83 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.202
r84 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.985
r85 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.22 $Y=0.995
+ $X2=5.22 $Y2=1.202
r86 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.22 $Y=0.995 $X2=5.22
+ $Y2=0.56
r87 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.202
r88 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
r89 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.75 $Y=0.995
+ $X2=4.75 $Y2=1.202
r90 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.75 $Y=0.995 $X2=4.75
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_4%A2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39 42
r75 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.065 $Y=1.202
+ $X2=8.09 $Y2=1.202
r76 37 39 22.6747 $w=3.72e-07 $l=1.75e-07 $layer=POLY_cond $X=7.89 $Y=1.202
+ $X2=8.065 $Y2=1.202
r77 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.89
+ $Y=1.16 $X2=7.89 $Y2=1.16
r78 35 37 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=7.595 $Y=1.202
+ $X2=7.89 $Y2=1.202
r79 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.57 $Y=1.202
+ $X2=7.595 $Y2=1.202
r80 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=7.125 $Y=1.202
+ $X2=7.57 $Y2=1.202
r81 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.1 $Y=1.202
+ $X2=7.125 $Y2=1.202
r82 30 32 49.2366 $w=3.72e-07 $l=3.8e-07 $layer=POLY_cond $X=6.72 $Y=1.202
+ $X2=7.1 $Y2=1.202
r83 30 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.72
+ $Y=1.16 $X2=6.72 $Y2=1.16
r84 28 30 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=6.655 $Y=1.202
+ $X2=6.72 $Y2=1.202
r85 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.63 $Y=1.202
+ $X2=6.655 $Y2=1.202
r86 25 38 15.8442 $w=2.08e-07 $l=3e-07 $layer=LI1_cond $X=7.59 $Y=1.18 $X2=7.89
+ $Y2=1.18
r87 25 42 47.2684 $w=2.08e-07 $l=8.95e-07 $layer=LI1_cond $X=7.59 $Y=1.18
+ $X2=6.695 $Y2=1.18
r88 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.09 $Y=0.995
+ $X2=8.09 $Y2=1.202
r89 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.09 $Y=0.995
+ $X2=8.09 $Y2=0.56
r90 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.065 $Y=1.41
+ $X2=8.065 $Y2=1.202
r91 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.065 $Y=1.41
+ $X2=8.065 $Y2=1.985
r92 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.595 $Y=1.41
+ $X2=7.595 $Y2=1.202
r93 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.595 $Y=1.41
+ $X2=7.595 $Y2=1.985
r94 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.57 $Y=0.995
+ $X2=7.57 $Y2=1.202
r95 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.57 $Y=0.995
+ $X2=7.57 $Y2=0.56
r96 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.202
r97 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.985
r98 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.1 $Y=0.995 $X2=7.1
+ $Y2=1.202
r99 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.1 $Y=0.995 $X2=7.1
+ $Y2=0.56
r100 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.202
r101 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.985
r102 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=1.202
r103 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_4%A_27_297# 1 2 3 4 5 6 7 8 9 28 30 32 36 38
+ 42 44 48 50 52 53 54 58 60 64 66 70 72 74 76 80 81 82 88 90 92
r116 74 94 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.3 $Y=1.625 $X2=8.3
+ $Y2=1.54
r117 74 76 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=8.3 $Y=1.625
+ $X2=8.3 $Y2=2.3
r118 73 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.485 $Y=1.54
+ $X2=7.36 $Y2=1.54
r119 72 94 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.175 $Y=1.54
+ $X2=8.3 $Y2=1.54
r120 72 73 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.175 $Y=1.54
+ $X2=7.485 $Y2=1.54
r121 68 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=1.625
+ $X2=7.36 $Y2=1.54
r122 68 70 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=7.36 $Y=1.625
+ $X2=7.36 $Y2=2.3
r123 67 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.545 $Y=1.54
+ $X2=6.42 $Y2=1.54
r124 66 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.235 $Y=1.54
+ $X2=7.36 $Y2=1.54
r125 66 67 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.235 $Y=1.54
+ $X2=6.545 $Y2=1.54
r126 62 90 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=1.625
+ $X2=6.42 $Y2=1.54
r127 62 64 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=6.42 $Y=1.625
+ $X2=6.42 $Y2=2.3
r128 61 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.605 $Y=1.54
+ $X2=5.48 $Y2=1.54
r129 60 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.295 $Y=1.54
+ $X2=6.42 $Y2=1.54
r130 60 61 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.295 $Y=1.54
+ $X2=5.605 $Y2=1.54
r131 56 88 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=1.625
+ $X2=5.48 $Y2=1.54
r132 56 58 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.48 $Y=1.625
+ $X2=5.48 $Y2=2.3
r133 55 84 9.25644 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=4.665 $Y=1.54
+ $X2=4.28 $Y2=1.54
r134 54 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.355 $Y=1.54
+ $X2=5.48 $Y2=1.54
r135 54 55 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.355 $Y=1.54
+ $X2=4.665 $Y2=1.54
r136 53 86 2.04363 $w=7.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.28 $Y=2.295
+ $X2=4.28 $Y2=2.38
r137 52 84 2.04363 $w=7.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.28 $Y=1.625
+ $X2=4.28 $Y2=1.54
r138 52 53 10.4074 $w=7.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.28 $Y=1.625
+ $X2=4.28 $Y2=2.295
r139 51 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.205 $Y=2.38
+ $X2=3.08 $Y2=2.38
r140 50 86 9.25644 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=3.895 $Y=2.38
+ $X2=4.28 $Y2=2.38
r141 50 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.895 $Y=2.38
+ $X2=3.205 $Y2=2.38
r142 46 82 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.295
+ $X2=3.08 $Y2=2.38
r143 46 48 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.08 $Y=2.295
+ $X2=3.08 $Y2=1.96
r144 45 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.265 $Y=2.38
+ $X2=2.14 $Y2=2.38
r145 44 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.955 $Y=2.38
+ $X2=3.08 $Y2=2.38
r146 44 45 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.955 $Y=2.38
+ $X2=2.265 $Y2=2.38
r147 40 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.295
+ $X2=2.14 $Y2=2.38
r148 40 42 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.14 $Y=2.295
+ $X2=2.14 $Y2=1.96
r149 39 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.325 $Y=2.38
+ $X2=1.2 $Y2=2.38
r150 38 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.015 $Y=2.38
+ $X2=2.14 $Y2=2.38
r151 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.015 $Y=2.38
+ $X2=1.325 $Y2=2.38
r152 34 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.295
+ $X2=1.2 $Y2=2.38
r153 34 36 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.2 $Y=2.295
+ $X2=1.2 $Y2=1.96
r154 33 79 5.18513 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.425 $Y=2.38
+ $X2=0.257 $Y2=2.38
r155 32 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.075 $Y=2.38
+ $X2=1.2 $Y2=2.38
r156 32 33 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.075 $Y=2.38
+ $X2=0.425 $Y2=2.38
r157 28 79 2.62343 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.257 $Y=2.295
+ $X2=0.257 $Y2=2.38
r158 28 30 22.5328 $w=3.33e-07 $l=6.55e-07 $layer=LI1_cond $X=0.257 $Y=2.295
+ $X2=0.257 $Y2=1.64
r159 9 94 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.155
+ $Y=1.485 $X2=8.3 $Y2=1.62
r160 9 76 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=8.155
+ $Y=1.485 $X2=8.3 $Y2=2.3
r161 8 92 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.215
+ $Y=1.485 $X2=7.36 $Y2=1.62
r162 8 70 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=7.215
+ $Y=1.485 $X2=7.36 $Y2=2.3
r163 7 90 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.275
+ $Y=1.485 $X2=6.42 $Y2=1.62
r164 7 64 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=6.275
+ $Y=1.485 $X2=6.42 $Y2=2.3
r165 6 88 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=1.62
r166 6 58 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=2.3
r167 5 86 200 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=3 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=2.3
r168 5 84 200 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=3 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=1.62
r169 4 48 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=1.96
r170 3 42 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.96
r171 2 36 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.96
r172 1 79 400 $w=1.7e-07 $l=8.95321e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.32
r173 1 30 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.64
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_4%Y 1 2 3 4 5 6 7 8 29 31 32 41 43 47 49 53
+ 55 56 57
c99 32 0 1.70485e-19 $X=2.545 $Y=1.445
r100 57 60 18.7929 $w=1.78e-07 $l=3.05e-07 $layer=LI1_cond $X=1.16 $Y=1.535
+ $X2=0.855 $Y2=1.535
r101 56 60 3.69874 $w=1.8e-07 $l=1.05e-07 $layer=LI1_cond $X=0.75 $Y=1.535
+ $X2=0.855 $Y2=1.535
r102 47 57 23.7222 $w=1.78e-07 $l=3.85e-07 $layer=LI1_cond $X=1.545 $Y=1.535
+ $X2=1.16 $Y2=1.535
r103 47 49 6.72674 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=1.545 $Y=1.535
+ $X2=1.67 $Y2=1.535
r104 44 53 4.43084 $w=1.8e-07 $l=1.7e-07 $layer=LI1_cond $X=2.735 $Y=1.535
+ $X2=2.565 $Y2=1.535
r105 43 55 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.425 $Y=1.535
+ $X2=3.55 $Y2=1.535
r106 43 44 42.5152 $w=1.78e-07 $l=6.9e-07 $layer=LI1_cond $X=3.425 $Y=1.535
+ $X2=2.735 $Y2=1.535
r107 39 41 45.1374 $w=2.38e-07 $l=9.4e-07 $layer=LI1_cond $X=5.01 $Y=0.765
+ $X2=5.95 $Y2=0.765
r108 37 39 70.1069 $w=2.38e-07 $l=1.46e-06 $layer=LI1_cond $X=3.55 $Y=0.765
+ $X2=5.01 $Y2=0.765
r109 35 51 3.84807 $w=2.4e-07 $l=1.5e-07 $layer=LI1_cond $X=2.695 $Y=0.765
+ $X2=2.545 $Y2=0.765
r110 35 37 41.0558 $w=2.38e-07 $l=8.55e-07 $layer=LI1_cond $X=2.695 $Y=0.765
+ $X2=3.55 $Y2=0.765
r111 32 53 1.86605 $w=3e-07 $l=9.94987e-08 $layer=LI1_cond $X=2.545 $Y=1.445
+ $X2=2.565 $Y2=1.535
r112 31 51 3.07845 $w=3e-07 $l=1.2e-07 $layer=LI1_cond $X=2.545 $Y=0.885
+ $X2=2.545 $Y2=0.765
r113 31 32 21.5123 $w=2.98e-07 $l=5.6e-07 $layer=LI1_cond $X=2.545 $Y=0.885
+ $X2=2.545 $Y2=1.445
r114 30 49 6.72674 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=1.795 $Y=1.535
+ $X2=1.67 $Y2=1.535
r115 29 53 4.43084 $w=1.8e-07 $l=1.7e-07 $layer=LI1_cond $X=2.395 $Y=1.535
+ $X2=2.565 $Y2=1.535
r116 29 30 36.9697 $w=1.78e-07 $l=6e-07 $layer=LI1_cond $X=2.395 $Y=1.535
+ $X2=1.795 $Y2=1.535
r117 8 55 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.62
r118 7 53 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.62
r119 6 49 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.62
r120 5 56 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.62
r121 4 41 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=5.765
+ $Y=0.235 $X2=5.95 $Y2=0.73
r122 3 39 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=4.825
+ $Y=0.235 $X2=5.01 $Y2=0.73
r123 2 37 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.73
r124 1 51 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_4%VPWR 1 2 3 4 15 19 23 27 30 31 33 34 36 37
+ 39 40 41 60 61
r102 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r103 58 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r104 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r105 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r106 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r107 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r108 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r109 49 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r110 48 49 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r111 44 48 300.107 $w=1.68e-07 $l=4.6e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=4.83 $Y2=2.72
r112 41 49 1.30889 $w=4.8e-07 $l=4.6e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=4.83 $Y2=2.72
r113 41 44 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r114 39 57 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.705 $Y=2.72
+ $X2=7.59 $Y2=2.72
r115 39 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.705 $Y=2.72
+ $X2=7.83 $Y2=2.72
r116 38 60 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=7.955 $Y=2.72
+ $X2=8.51 $Y2=2.72
r117 38 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.955 $Y=2.72
+ $X2=7.83 $Y2=2.72
r118 36 54 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=6.765 $Y=2.72
+ $X2=6.67 $Y2=2.72
r119 36 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.765 $Y=2.72
+ $X2=6.89 $Y2=2.72
r120 35 57 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=7.015 $Y=2.72
+ $X2=7.59 $Y2=2.72
r121 35 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.015 $Y=2.72
+ $X2=6.89 $Y2=2.72
r122 33 51 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.825 $Y=2.72
+ $X2=5.75 $Y2=2.72
r123 33 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.825 $Y=2.72
+ $X2=5.95 $Y2=2.72
r124 32 54 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=6.075 $Y=2.72
+ $X2=6.67 $Y2=2.72
r125 32 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.075 $Y=2.72
+ $X2=5.95 $Y2=2.72
r126 30 48 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.885 $Y=2.72
+ $X2=4.83 $Y2=2.72
r127 30 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.885 $Y=2.72
+ $X2=5.01 $Y2=2.72
r128 29 51 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.135 $Y=2.72
+ $X2=5.75 $Y2=2.72
r129 29 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.135 $Y=2.72
+ $X2=5.01 $Y2=2.72
r130 25 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.83 $Y=2.635
+ $X2=7.83 $Y2=2.72
r131 25 27 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=7.83 $Y=2.635
+ $X2=7.83 $Y2=1.96
r132 21 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=2.635
+ $X2=6.89 $Y2=2.72
r133 21 23 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=6.89 $Y=2.635
+ $X2=6.89 $Y2=1.96
r134 17 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=2.635
+ $X2=5.95 $Y2=2.72
r135 17 19 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.95 $Y=2.635
+ $X2=5.95 $Y2=1.96
r136 13 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.01 $Y=2.635
+ $X2=5.01 $Y2=2.72
r137 13 15 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.01 $Y=2.635
+ $X2=5.01 $Y2=1.96
r138 4 27 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=7.685
+ $Y=1.485 $X2=7.83 $Y2=1.96
r139 3 23 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=1.96
r140 2 19 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=1.96
r141 1 15 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_4%A_27_47# 1 2 3 4 5 18 20 21 24 26 28 29 34
+ 36
c72 29 0 1.56657e-19 $X=2.075 $Y=0.725
r73 32 34 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=3.08 $Y=0.365
+ $X2=4.02 $Y2=0.365
r74 30 38 4.05488 $w=2.2e-07 $l=1.5e-07 $layer=LI1_cond $X=2.225 $Y=0.365
+ $X2=2.075 $Y2=0.365
r75 30 32 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=2.225 $Y=0.365
+ $X2=3.08 $Y2=0.365
r76 29 40 2.76965 $w=3e-07 $l=9e-08 $layer=LI1_cond $X=2.075 $Y=0.725 $X2=2.075
+ $Y2=0.815
r77 28 38 2.97358 $w=3e-07 $l=1.1e-07 $layer=LI1_cond $X=2.075 $Y=0.475
+ $X2=2.075 $Y2=0.365
r78 28 29 9.60369 $w=2.98e-07 $l=2.5e-07 $layer=LI1_cond $X=2.075 $Y=0.475
+ $X2=2.075 $Y2=0.725
r79 27 36 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.365 $Y=0.815
+ $X2=1.175 $Y2=0.815
r80 26 40 4.61608 $w=1.8e-07 $l=1.5e-07 $layer=LI1_cond $X=1.925 $Y=0.815
+ $X2=2.075 $Y2=0.815
r81 26 27 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.925 $Y=0.815
+ $X2=1.365 $Y2=0.815
r82 22 36 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=1.175 $Y=0.725
+ $X2=1.175 $Y2=0.815
r83 22 24 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.175 $Y=0.725
+ $X2=1.175 $Y2=0.39
r84 20 36 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=0.985 $Y=0.815
+ $X2=1.175 $Y2=0.815
r85 20 21 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=0.985 $Y=0.815
+ $X2=0.425 $Y2=0.815
r86 16 21 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.26 $Y=0.725
+ $X2=0.425 $Y2=0.815
r87 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.26 $Y=0.725
+ $X2=0.26 $Y2=0.39
r88 5 34 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=3.835
+ $Y=0.235 $X2=4.02 $Y2=0.39
r89 4 32 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.39
r90 3 40 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.73
r91 3 38 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.39
r92 2 24 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.39
r93 1 18 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_4%VGND 1 2 3 4 17 19 23 27 31 34 35 37 38 39
+ 52 53 56 59 62
r113 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r114 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r115 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r116 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r117 50 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.51
+ $Y2=0
r118 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r119 47 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.59
+ $Y2=0
r120 46 47 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r121 44 47 1.30889 $w=4.8e-07 $l=4.6e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=6.67
+ $Y2=0
r122 44 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r123 43 46 300.107 $w=1.68e-07 $l=4.6e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=6.67
+ $Y2=0
r124 43 44 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r125 41 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=0 $X2=1.67
+ $Y2=0
r126 41 43 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.755 $Y=0
+ $X2=2.07 $Y2=0
r127 39 57 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r128 39 62 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r129 37 49 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.59 $Y2=0
r130 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.745 $Y=0 $X2=7.83
+ $Y2=0
r131 36 52 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=7.915 $Y=0
+ $X2=8.51 $Y2=0
r132 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.915 $Y=0 $X2=7.83
+ $Y2=0
r133 34 46 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.805 $Y=0
+ $X2=6.67 $Y2=0
r134 34 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.805 $Y=0 $X2=6.89
+ $Y2=0
r135 33 49 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=6.975 $Y=0 $X2=7.59
+ $Y2=0
r136 33 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.975 $Y=0 $X2=6.89
+ $Y2=0
r137 29 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.83 $Y=0.085
+ $X2=7.83 $Y2=0
r138 29 31 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.83 $Y=0.085
+ $X2=7.83 $Y2=0.39
r139 25 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=0.085
+ $X2=6.89 $Y2=0
r140 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.89 $Y=0.085
+ $X2=6.89 $Y2=0.39
r141 21 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0
r142 21 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0.39
r143 20 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.73
+ $Y2=0
r144 19 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=0 $X2=1.67
+ $Y2=0
r145 19 20 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.585 $Y=0
+ $X2=0.815 $Y2=0
r146 15 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r147 15 17 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.39
r148 4 31 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=7.645
+ $Y=0.235 $X2=7.83 $Y2=0.39
r149 3 27 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=6.705
+ $Y=0.235 $X2=6.89 $Y2=0.39
r150 2 23 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.39
r151 1 17 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_4%A_883_47# 1 2 3 4 5 16 22 23 24 28 30 34
+ 40
r68 32 34 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=8.275 $Y=0.725
+ $X2=8.275 $Y2=0.39
r69 31 40 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=7.525 $Y=0.815
+ $X2=7.335 $Y2=0.815
r70 30 32 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=8.085 $Y=0.815
+ $X2=8.275 $Y2=0.725
r71 30 31 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=8.085 $Y=0.815
+ $X2=7.525 $Y2=0.815
r72 26 40 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=7.335 $Y=0.725
+ $X2=7.335 $Y2=0.815
r73 26 28 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.335 $Y=0.725
+ $X2=7.335 $Y2=0.39
r74 25 39 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=6.585 $Y=0.815
+ $X2=6.46 $Y2=0.815
r75 24 40 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=7.145 $Y=0.815
+ $X2=7.335 $Y2=0.815
r76 24 25 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=7.145 $Y=0.815
+ $X2=6.585 $Y2=0.815
r77 23 39 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=6.46 $Y=0.725 $X2=6.46
+ $Y2=0.815
r78 22 37 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=6.46 $Y=0.475
+ $X2=6.46 $Y2=0.365
r79 22 23 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=6.46 $Y=0.475
+ $X2=6.46 $Y2=0.725
r80 18 21 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=4.54 $Y=0.365
+ $X2=5.48 $Y2=0.365
r81 16 37 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=6.335 $Y=0.365
+ $X2=6.46 $Y2=0.365
r82 16 21 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=6.335 $Y=0.365
+ $X2=5.48 $Y2=0.365
r83 5 34 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=8.165
+ $Y=0.235 $X2=8.3 $Y2=0.39
r84 4 28 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=7.175
+ $Y=0.235 $X2=7.36 $Y2=0.39
r85 3 39 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=6.285
+ $Y=0.235 $X2=6.42 $Y2=0.73
r86 3 37 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.285
+ $Y=0.235 $X2=6.42 $Y2=0.39
r87 2 21 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=5.295
+ $Y=0.235 $X2=5.48 $Y2=0.39
r88 1 18 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=4.415
+ $Y=0.235 $X2=4.54 $Y2=0.39
.ends

