* File: sky130_fd_sc_hdll__and3_2.pex.spice
* Created: Wed Sep  2 08:22:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND3_2%A 1 3 6 8
r26 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r27 8 12 9.27941 $w=3.83e-07 $l=3.1e-07 $layer=LI1_cond $X=0.277 $Y=0.85
+ $X2=0.277 $Y2=1.16
r28 4 11 39.2698 $w=3.83e-07 $l=2.31571e-07 $layer=POLY_cond $X=0.535 $Y=0.995
+ $X2=0.375 $Y2=1.16
r29 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.535 $Y=0.995
+ $X2=0.535 $Y2=0.475
r30 1 11 53.9003 $w=3.83e-07 $l=3.79473e-07 $layer=POLY_cond $X=0.505 $Y=1.48
+ $X2=0.375 $Y2=1.16
r31 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.505 $Y=1.48
+ $X2=0.505 $Y2=1.765
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_2%B 1 3 6 8 9 17
r44 13 17 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=1.03 $Y=2.295
+ $X2=1.15 $Y2=2.295
r45 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.03
+ $Y=2.3 $X2=1.03 $Y2=2.3
r46 9 17 3.38954 $w=3.38e-07 $l=1e-07 $layer=LI1_cond $X=1.25 $Y=2.295 $X2=1.15
+ $Y2=2.295
r47 6 12 38.3834 $w=3.29e-07 $l=2.27321e-07 $layer=POLY_cond $X=0.975 $Y=2.105
+ $X2=1.045 $Y2=2.3
r48 6 8 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=0.975 $Y=2.105
+ $X2=0.975 $Y2=1.765
r49 5 8 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.975 $Y=1.48
+ $X2=0.975 $Y2=1.765
r50 1 5 44 $w=2.41e-07 $l=2.56905e-07 $layer=POLY_cond $X=0.895 $Y=1.26
+ $X2=0.975 $Y2=1.48
r51 1 3 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=0.895 $Y=1.26
+ $X2=0.895 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_2%C 3 5 7 8 9
c45 5 0 9.98623e-20 $X=1.5 $Y=1.41
r46 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.41
+ $Y=1.16 $X2=1.41 $Y2=1.16
r47 9 20 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=1.19 $Y=0.51 $X2=1.19
+ $Y2=0.75
r48 8 14 6.62115 $w=5.58e-07 $l=3.1e-07 $layer=LI1_cond $X=1.345 $Y=0.85
+ $X2=1.345 $Y2=1.16
r49 8 20 5.85187 $w=5.58e-07 $l=1e-07 $layer=LI1_cond $X=1.345 $Y=0.85 $X2=1.345
+ $Y2=0.75
r50 5 13 47.4309 $w=3.07e-07 $l=2.77489e-07 $layer=POLY_cond $X=1.5 $Y=1.41
+ $X2=1.442 $Y2=1.16
r51 5 7 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.5 $Y=1.41 $X2=1.5
+ $Y2=1.695
r52 1 13 38.5336 $w=3.07e-07 $l=2.05925e-07 $layer=POLY_cond $X=1.35 $Y=0.995
+ $X2=1.442 $Y2=1.16
r53 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.35 $Y=0.995 $X2=1.35
+ $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_2%A_29_311# 1 2 3 10 12 13 15 16 18 19 21 24
+ 26 30 31 33 34 36 40 43 44 52
c105 34 0 9.98623e-20 $X=1.18 $Y=1.51
r106 52 53 3.8871 $w=3.72e-07 $l=3e-08 $layer=POLY_cond $X=2.515 $Y=1.202
+ $X2=2.545 $Y2=1.202
r107 51 52 59.6021 $w=3.72e-07 $l=4.6e-07 $layer=POLY_cond $X=2.055 $Y=1.202
+ $X2=2.515 $Y2=1.202
r108 50 51 1.2957 $w=3.72e-07 $l=1e-08 $layer=POLY_cond $X=2.045 $Y=1.202
+ $X2=2.055 $Y2=1.202
r109 44 47 8.25918 $w=2.98e-07 $l=2.15e-07 $layer=LI1_cond $X=1.33 $Y=1.51
+ $X2=1.33 $Y2=1.725
r110 41 50 11.6613 $w=3.72e-07 $l=9e-08 $layer=POLY_cond $X=1.955 $Y=1.202
+ $X2=2.045 $Y2=1.202
r111 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.955
+ $Y=1.16 $X2=1.955 $Y2=1.16
r112 38 40 13.2781 $w=2.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.925 $Y=1.425
+ $X2=1.925 $Y2=1.16
r113 37 44 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.48 $Y=1.51 $X2=1.33
+ $Y2=1.51
r114 36 38 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.81 $Y=1.51
+ $X2=1.925 $Y2=1.425
r115 36 37 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.81 $Y=1.51
+ $X2=1.48 $Y2=1.51
r116 35 43 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=0.895 $Y=1.51
+ $X2=0.792 $Y2=1.51
r117 34 44 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.18 $Y=1.51 $X2=1.33
+ $Y2=1.51
r118 34 35 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.18 $Y=1.51
+ $X2=0.895 $Y2=1.51
r119 33 43 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.792 $Y=1.425
+ $X2=0.792 $Y2=1.51
r120 32 33 46.2572 $w=2.03e-07 $l=8.55e-07 $layer=LI1_cond $X=0.792 $Y=0.57
+ $X2=0.792 $Y2=1.425
r121 30 43 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=0.69 $Y=1.51
+ $X2=0.792 $Y2=1.51
r122 30 31 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.69 $Y=1.51
+ $X2=0.355 $Y2=1.51
r123 26 32 6.96198 $w=2.65e-07 $l=1.76791e-07 $layer=LI1_cond $X=0.69 $Y=0.437
+ $X2=0.792 $Y2=0.57
r124 26 28 18.0477 $w=2.63e-07 $l=4.15e-07 $layer=LI1_cond $X=0.69 $Y=0.437
+ $X2=0.275 $Y2=0.437
r125 22 31 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.227 $Y=1.595
+ $X2=0.355 $Y2=1.51
r126 22 24 7.45698 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.227 $Y=1.595
+ $X2=0.227 $Y2=1.76
r127 19 53 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.545 $Y=0.995
+ $X2=2.545 $Y2=1.202
r128 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.545 $Y=0.995
+ $X2=2.545 $Y2=0.56
r129 16 52 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.515 $Y=1.41
+ $X2=2.515 $Y2=1.202
r130 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.515 $Y=1.41
+ $X2=2.515 $Y2=1.985
r131 13 51 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.055 $Y=0.995
+ $X2=2.055 $Y2=1.202
r132 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.055 $Y=0.995
+ $X2=2.055 $Y2=0.56
r133 10 50 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.045 $Y=1.41
+ $X2=2.045 $Y2=1.202
r134 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.045 $Y=1.41
+ $X2=2.045 $Y2=1.985
r135 3 47 600 $w=1.7e-07 $l=2.72029e-07 $layer=licon1_PDIFF $count=1 $X=1.065
+ $Y=1.555 $X2=1.265 $Y2=1.725
r136 2 24 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.555 $X2=0.27 $Y2=1.76
r137 1 28 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.265 $X2=0.275 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_2%VPWR 1 2 3 11 14 16 18 23 26 27 28 34 39 45
r55 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r56 39 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r57 37 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r58 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r59 34 44 4.0276 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.79 $Y=2.72
+ $X2=3.005 $Y2=2.72
r60 34 36 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.79 $Y=2.72
+ $X2=2.53 $Y2=2.72
r61 33 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r62 33 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r63 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r64 30 39 9.33093 $w=1.7e-07 $l=3.83e-07 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=0.382 $Y2=2.72
r65 30 32 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=1.61 $Y2=2.72
r66 28 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r67 28 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r68 26 32 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.705 $Y=2.72
+ $X2=1.61 $Y2=2.72
r69 26 27 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=1.705 $Y=2.72
+ $X2=1.812 $Y2=2.72
r70 25 36 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.92 $Y=2.72
+ $X2=2.53 $Y2=2.72
r71 25 27 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=1.92 $Y=2.72
+ $X2=1.812 $Y2=2.72
r72 16 44 3.18462 $w=2.6e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.92 $Y=2.635
+ $X2=3.005 $Y2=2.72
r73 16 18 29.9192 $w=2.58e-07 $l=6.75e-07 $layer=LI1_cond $X=2.92 $Y=2.635
+ $X2=2.92 $Y2=1.96
r74 12 27 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.812 $Y=2.635
+ $X2=1.812 $Y2=2.72
r75 12 14 36.4494 $w=2.13e-07 $l=6.8e-07 $layer=LI1_cond $X=1.812 $Y=2.635
+ $X2=1.812 $Y2=1.955
r76 11 39 15.9 $w=7.01e-07 $l=7.09415e-07 $layer=LI1_cond $X=0.645 $Y=2.13
+ $X2=0.382 $Y2=2.72
r77 10 23 5.54545 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=0.645 $Y=1.86
+ $X2=0.74 $Y2=1.86
r78 10 11 8.40323 $w=2.38e-07 $l=1.75e-07 $layer=LI1_cond $X=0.645 $Y=1.955
+ $X2=0.645 $Y2=2.13
r79 3 18 300 $w=1.7e-07 $l=5.94874e-07 $layer=licon1_PDIFF $count=2 $X=2.605
+ $Y=1.485 $X2=2.875 $Y2=1.96
r80 2 14 300 $w=1.7e-07 $l=5.69473e-07 $layer=licon1_PDIFF $count=2 $X=1.59
+ $Y=1.485 $X2=1.81 $Y2=1.955
r81 1 23 600 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.555 $X2=0.74 $Y2=1.85
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_2%X 1 2 11 12 13 24 25 31
r30 25 32 11.2043 $w=3.58e-07 $l=3.5e-07 $layer=LI1_cond $X=2.44 $Y=1.795
+ $X2=2.44 $Y2=1.445
r31 24 25 4.89848 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=1.96
+ $X2=2.395 $Y2=1.795
r32 22 31 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.345 $Y=0.715
+ $X2=2.345 $Y2=0.925
r33 21 22 9.3792 $w=4.43e-07 $l=1.85e-07 $layer=LI1_cond $X=2.207 $Y=0.53
+ $X2=2.207 $Y2=0.715
r34 13 32 7.08564 $w=6.63e-07 $l=2.55e-07 $layer=LI1_cond $X=2.592 $Y=1.19
+ $X2=2.592 $Y2=1.445
r35 13 31 12.3779 $w=6.63e-07 $l=2.65e-07 $layer=LI1_cond $X=2.592 $Y=1.19
+ $X2=2.592 $Y2=0.925
r36 12 24 6.64488 $w=4.48e-07 $l=2.5e-07 $layer=LI1_cond $X=2.395 $Y=2.21
+ $X2=2.395 $Y2=1.96
r37 11 21 0.517952 $w=4.43e-07 $l=2e-08 $layer=LI1_cond $X=2.207 $Y=0.51
+ $X2=2.207 $Y2=0.53
r38 2 24 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.135
+ $Y=1.485 $X2=2.28 $Y2=1.96
r39 1 21 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=2.13
+ $Y=0.235 $X2=2.265 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_2%VGND 1 2 9 11 13 15 17 25 31 35
r35 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r36 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r37 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r38 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r39 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r40 26 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.65
+ $Y2=0
r41 26 28 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=2.53
+ $Y2=0
r42 25 34 4.06435 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.957
+ $Y2=0
r43 25 28 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.53
+ $Y2=0
r44 24 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r45 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r46 19 23 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r47 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=0 $X2=1.65
+ $Y2=0
r48 17 23 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.485 $Y=0 $X2=1.15
+ $Y2=0
r49 15 24 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r50 15 19 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r51 11 34 3.25769 $w=2.75e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.832 $Y=0.085
+ $X2=2.957 $Y2=0
r52 11 13 18.02 $w=2.73e-07 $l=4.3e-07 $layer=LI1_cond $X=2.832 $Y=0.085
+ $X2=2.832 $Y2=0.515
r53 7 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=0.085 $X2=1.65
+ $Y2=0
r54 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.65 $Y=0.085 $X2=1.65
+ $Y2=0.495
r55 2 13 182 $w=1.7e-07 $l=3.50999e-07 $layer=licon1_NDIFF $count=1 $X=2.62
+ $Y=0.235 $X2=2.78 $Y2=0.515
r56 1 9 182 $w=1.7e-07 $l=3.23497e-07 $layer=licon1_NDIFF $count=1 $X=1.425
+ $Y=0.265 $X2=1.65 $Y2=0.495
.ends

