* File: sky130_fd_sc_hdll__a21oi_2.pxi.spice
* Created: Wed Sep  2 08:17:48 2020
* 
x_PM_SKY130_FD_SC_HDLL__A21OI_2%A2 N_A2_c_50_n N_A2_M1000_g N_A2_M1003_g
+ N_A2_c_52_n N_A2_M1007_g N_A2_c_53_n N_A2_M1011_g N_A2_c_62_p N_A2_c_54_n A2
+ N_A2_c_55_n PM_SKY130_FD_SC_HDLL__A21OI_2%A2
x_PM_SKY130_FD_SC_HDLL__A21OI_2%A1 N_A1_c_126_n N_A1_M1008_g N_A1_c_130_n
+ N_A1_M1001_g N_A1_c_131_n N_A1_M1006_g N_A1_c_127_n N_A1_M1005_g A1
+ N_A1_c_128_n N_A1_c_129_n A1 PM_SKY130_FD_SC_HDLL__A21OI_2%A1
x_PM_SKY130_FD_SC_HDLL__A21OI_2%B1 N_B1_M1002_g N_B1_c_178_n N_B1_M1009_g
+ N_B1_M1004_g N_B1_c_179_n N_B1_M1010_g N_B1_c_175_n B1 B1 N_B1_c_177_n
+ PM_SKY130_FD_SC_HDLL__A21OI_2%B1
x_PM_SKY130_FD_SC_HDLL__A21OI_2%A_27_297# N_A_27_297#_M1000_s
+ N_A_27_297#_M1001_s N_A_27_297#_M1011_s N_A_27_297#_M1010_d
+ N_A_27_297#_c_225_n N_A_27_297#_c_226_n N_A_27_297#_c_234_n
+ N_A_27_297#_c_260_p N_A_27_297#_c_237_n N_A_27_297#_c_239_n
+ N_A_27_297#_c_241_n N_A_27_297#_c_227_n N_A_27_297#_c_242_n
+ N_A_27_297#_c_228_n N_A_27_297#_c_243_n
+ PM_SKY130_FD_SC_HDLL__A21OI_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A21OI_2%VPWR N_VPWR_M1000_d N_VPWR_M1006_d
+ N_VPWR_c_288_n N_VPWR_c_289_n N_VPWR_c_290_n VPWR N_VPWR_c_291_n
+ N_VPWR_c_292_n N_VPWR_c_287_n N_VPWR_c_294_n
+ PM_SKY130_FD_SC_HDLL__A21OI_2%VPWR
x_PM_SKY130_FD_SC_HDLL__A21OI_2%Y N_Y_M1008_s N_Y_M1002_s N_Y_M1009_s
+ N_Y_c_343_n N_Y_c_346_n N_Y_c_342_n N_Y_c_350_n N_Y_c_364_n N_Y_c_366_n Y
+ N_Y_c_367_n PM_SKY130_FD_SC_HDLL__A21OI_2%Y
x_PM_SKY130_FD_SC_HDLL__A21OI_2%VGND N_VGND_M1003_d N_VGND_M1007_d
+ N_VGND_M1004_d N_VGND_c_390_n N_VGND_c_391_n N_VGND_c_392_n N_VGND_c_393_n
+ VGND N_VGND_c_394_n N_VGND_c_395_n N_VGND_c_396_n N_VGND_c_397_n
+ PM_SKY130_FD_SC_HDLL__A21OI_2%VGND
cc_1 VNB N_A2_c_50_n 0.0319731f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_2 VNB N_A2_M1003_g 0.0239603f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.56
cc_3 VNB N_A2_c_52_n 0.0165896f $X=-0.19 $Y=-0.24 $X2=1.86 $Y2=0.995
cc_4 VNB N_A2_c_53_n 0.0222715f $X=-0.19 $Y=-0.24 $X2=1.945 $Y2=1.41
cc_5 VNB N_A2_c_54_n 0.00370446f $X=-0.19 $Y=-0.24 $X2=1.92 $Y2=1.16
cc_6 VNB N_A2_c_55_n 0.0165013f $X=-0.19 $Y=-0.24 $X2=0.4 $Y2=1.16
cc_7 VNB N_A1_c_126_n 0.0173559f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_8 VNB N_A1_c_127_n 0.0166612f $X=-0.19 $Y=-0.24 $X2=1.86 $Y2=0.56
cc_9 VNB N_A1_c_128_n 0.00471933f $X=-0.19 $Y=-0.24 $X2=1.92 $Y2=1.16
cc_10 VNB N_A1_c_129_n 0.0345699f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B1_M1002_g 0.0181604f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.985
cc_12 VNB N_B1_M1004_g 0.0230561f $X=-0.19 $Y=-0.24 $X2=1.86 $Y2=0.56
cc_13 VNB N_B1_c_175_n 0.0322809f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.585
cc_14 VNB B1 0.0229957f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B1_c_177_n 0.0271178f $X=-0.19 $Y=-0.24 $X2=0.4 $Y2=1.16
cc_16 VNB N_VPWR_c_287_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_390_n 0.0110651f $X=-0.19 $Y=-0.24 $X2=1.86 $Y2=0.56
cc_18 VNB N_VGND_c_391_n 0.030651f $X=-0.19 $Y=-0.24 $X2=1.945 $Y2=1.985
cc_19 VNB N_VGND_c_392_n 0.0166826f $X=-0.19 $Y=-0.24 $X2=1.755 $Y2=1.585
cc_20 VNB N_VGND_c_393_n 0.0287266f $X=-0.19 $Y=-0.24 $X2=1.942 $Y2=1.495
cc_21 VNB N_VGND_c_394_n 0.0409256f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_395_n 0.0212545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_396_n 0.00922167f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_397_n 0.2058f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VPB N_A2_c_50_n 0.0313087f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_26 VPB N_A2_c_53_n 0.0247855f $X=-0.19 $Y=1.305 $X2=1.945 $Y2=1.41
cc_27 VPB N_A2_c_54_n 0.00327823f $X=-0.19 $Y=1.305 $X2=1.92 $Y2=1.16
cc_28 VPB N_A2_c_55_n 0.00908318f $X=-0.19 $Y=1.305 $X2=0.4 $Y2=1.16
cc_29 VPB N_A1_c_130_n 0.0163995f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.015
cc_30 VPB N_A1_c_131_n 0.016507f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_A1_c_128_n 2.50904e-19 $X=-0.19 $Y=1.305 $X2=1.92 $Y2=1.16
cc_32 VPB N_A1_c_129_n 0.0196114f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_B1_c_178_n 0.0163998f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.56
cc_34 VPB N_B1_c_179_n 0.0188133f $X=-0.19 $Y=1.305 $X2=1.945 $Y2=1.985
cc_35 VPB N_B1_c_175_n 0.0210614f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.585
cc_36 VPB B1 0.0213099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_B1_c_177_n 0.00963904f $X=-0.19 $Y=1.305 $X2=0.4 $Y2=1.16
cc_38 VPB N_A_27_297#_c_225_n 0.0113777f $X=-0.19 $Y=1.305 $X2=1.945 $Y2=1.985
cc_39 VPB N_A_27_297#_c_226_n 0.0134872f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.585
cc_40 VPB N_A_27_297#_c_227_n 0.00795084f $X=-0.19 $Y=1.305 $X2=0.42 $Y2=1.16
cc_41 VPB N_A_27_297#_c_228_n 0.0192574f $X=-0.19 $Y=1.305 $X2=0.42 $Y2=1.585
cc_42 VPB N_VPWR_c_288_n 0.00474148f $X=-0.19 $Y=1.305 $X2=1.86 $Y2=0.56
cc_43 VPB N_VPWR_c_289_n 0.0174821f $X=-0.19 $Y=1.305 $X2=1.945 $Y2=1.985
cc_44 VPB N_VPWR_c_290_n 0.00324214f $X=-0.19 $Y=1.305 $X2=1.945 $Y2=1.985
cc_45 VPB N_VPWR_c_291_n 0.0150764f $X=-0.19 $Y=1.305 $X2=1.942 $Y2=1.495
cc_46 VPB N_VPWR_c_292_n 0.0479263f $X=-0.19 $Y=1.305 $X2=0.42 $Y2=1.53
cc_47 VPB N_VPWR_c_287_n 0.0530135f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_294_n 0.00556536f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_Y_c_342_n 0.00118595f $X=-0.19 $Y=1.305 $X2=1.942 $Y2=1.495
cc_50 N_A2_M1003_g N_A1_c_126_n 0.0290468f $X=0.54 $Y=0.56 $X2=-0.19 $Y2=-0.24
cc_51 N_A2_c_50_n N_A1_c_130_n 0.0375701f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_52 N_A2_c_62_p N_A1_c_130_n 0.0119274f $X=1.755 $Y=1.585 $X2=0 $Y2=0
cc_53 N_A2_c_55_n N_A1_c_130_n 0.00232217f $X=0.4 $Y=1.16 $X2=0 $Y2=0
cc_54 N_A2_c_53_n N_A1_c_131_n 0.0396504f $X=1.945 $Y=1.41 $X2=0 $Y2=0
cc_55 N_A2_c_62_p N_A1_c_131_n 0.0123811f $X=1.755 $Y=1.585 $X2=0 $Y2=0
cc_56 N_A2_c_54_n N_A1_c_131_n 0.00200016f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_57 N_A2_c_52_n N_A1_c_127_n 0.0388415f $X=1.86 $Y=0.995 $X2=0 $Y2=0
cc_58 N_A2_c_50_n N_A1_c_128_n 3.2034e-19 $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_59 N_A2_M1003_g N_A1_c_128_n 2.52545e-19 $X=0.54 $Y=0.56 $X2=0 $Y2=0
cc_60 N_A2_c_53_n N_A1_c_128_n 8.49791e-19 $X=1.945 $Y=1.41 $X2=0 $Y2=0
cc_61 N_A2_c_62_p N_A1_c_128_n 0.0446363f $X=1.755 $Y=1.585 $X2=0 $Y2=0
cc_62 N_A2_c_54_n N_A1_c_128_n 0.0202035f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A2_c_55_n N_A1_c_128_n 0.0223121f $X=0.4 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A2_c_50_n N_A1_c_129_n 0.0290468f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_65 N_A2_c_53_n N_A1_c_129_n 0.0425455f $X=1.945 $Y=1.41 $X2=0 $Y2=0
cc_66 N_A2_c_62_p N_A1_c_129_n 0.00639214f $X=1.755 $Y=1.585 $X2=0 $Y2=0
cc_67 N_A2_c_54_n N_A1_c_129_n 0.00290823f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A2_c_55_n N_A1_c_129_n 0.00332724f $X=0.4 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A2_c_52_n N_B1_M1002_g 0.0183355f $X=1.86 $Y=0.995 $X2=0 $Y2=0
cc_70 N_A2_c_53_n N_B1_M1002_g 0.0221345f $X=1.945 $Y=1.41 $X2=0 $Y2=0
cc_71 N_A2_c_53_n N_B1_c_178_n 0.0236146f $X=1.945 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A2_c_62_p N_B1_c_178_n 0.00170522f $X=1.755 $Y=1.585 $X2=0 $Y2=0
cc_73 N_A2_c_54_n N_B1_c_178_n 7.24621e-19 $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A2_c_53_n N_B1_c_175_n 0.00370749f $X=1.945 $Y=1.41 $X2=0 $Y2=0
cc_75 N_A2_c_54_n N_B1_c_175_n 0.00260883f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A2_c_55_n N_A_27_297#_M1000_s 0.0118476f $X=0.4 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_77 N_A2_c_62_p N_A_27_297#_M1001_s 0.00358863f $X=1.755 $Y=1.585 $X2=0 $Y2=0
cc_78 N_A2_c_62_p N_A_27_297#_M1011_s 0.00264939f $X=1.755 $Y=1.585 $X2=0 $Y2=0
cc_79 N_A2_c_50_n N_A_27_297#_c_225_n 4.88387e-19 $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A2_c_55_n N_A_27_297#_c_225_n 0.0189341f $X=0.4 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A2_c_50_n N_A_27_297#_c_234_n 0.0132291f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A2_c_62_p N_A_27_297#_c_234_n 0.0235789f $X=1.755 $Y=1.585 $X2=0 $Y2=0
cc_83 N_A2_c_55_n N_A_27_297#_c_234_n 0.0158987f $X=0.4 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A2_c_53_n N_A_27_297#_c_237_n 0.010823f $X=1.945 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A2_c_62_p N_A_27_297#_c_237_n 0.0362212f $X=1.755 $Y=1.585 $X2=0 $Y2=0
cc_86 N_A2_c_53_n N_A_27_297#_c_239_n 7.36455e-19 $X=1.945 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A2_c_62_p N_A_27_297#_c_239_n 0.00473113f $X=1.755 $Y=1.585 $X2=0 $Y2=0
cc_88 N_A2_c_53_n N_A_27_297#_c_241_n 0.00418949f $X=1.945 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A2_c_53_n N_A_27_297#_c_242_n 0.00227366f $X=1.945 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A2_c_62_p N_A_27_297#_c_243_n 0.0131878f $X=1.755 $Y=1.585 $X2=0 $Y2=0
cc_91 N_A2_c_62_p N_VPWR_M1000_d 0.00797279f $X=1.755 $Y=1.585 $X2=-0.19
+ $Y2=-0.24
cc_92 N_A2_c_55_n N_VPWR_M1000_d 9.5006e-19 $X=0.4 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_93 N_A2_c_62_p N_VPWR_M1006_d 0.0069012f $X=1.755 $Y=1.585 $X2=0 $Y2=0
cc_94 N_A2_c_53_n N_VPWR_c_288_n 0.0039542f $X=1.945 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A2_c_50_n N_VPWR_c_291_n 0.0032362f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A2_c_53_n N_VPWR_c_292_n 0.0051032f $X=1.945 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A2_c_50_n N_VPWR_c_287_n 0.00474648f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A2_c_53_n N_VPWR_c_287_n 0.00678224f $X=1.945 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A2_c_50_n N_VPWR_c_294_n 0.0104644f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A2_c_52_n N_Y_c_343_n 0.0122033f $X=1.86 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A2_c_53_n N_Y_c_343_n 0.00405236f $X=1.945 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A2_c_54_n N_Y_c_343_n 0.0169781f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A2_c_52_n N_Y_c_346_n 0.001021f $X=1.86 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A2_c_53_n N_Y_c_346_n 7.1307e-19 $X=1.945 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A2_c_54_n N_Y_c_346_n 0.0143619f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A2_c_54_n N_Y_c_342_n 0.00756296f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A2_M1003_g N_Y_c_350_n 0.0016586f $X=0.54 $Y=0.56 $X2=0 $Y2=0
cc_108 N_A2_c_50_n N_VGND_c_391_n 0.00369598f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A2_M1003_g N_VGND_c_391_n 0.0113338f $X=0.54 $Y=0.56 $X2=0 $Y2=0
cc_110 N_A2_c_55_n N_VGND_c_391_n 0.0219794f $X=0.4 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A2_M1003_g N_VGND_c_394_n 0.00585385f $X=0.54 $Y=0.56 $X2=0 $Y2=0
cc_112 N_A2_c_52_n N_VGND_c_394_n 0.0035176f $X=1.86 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A2_c_52_n N_VGND_c_396_n 0.0088425f $X=1.86 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A2_M1003_g N_VGND_c_397_n 0.0117318f $X=0.54 $Y=0.56 $X2=0 $Y2=0
cc_115 N_A2_c_52_n N_VGND_c_397_n 0.00395487f $X=1.86 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A1_c_130_n N_A_27_297#_c_234_n 0.013666f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A1_c_131_n N_A_27_297#_c_237_n 0.0117763f $X=1.475 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A1_c_131_n N_A_27_297#_c_241_n 7.50844e-19 $X=1.475 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A1_c_131_n N_VPWR_c_288_n 0.00426997f $X=1.475 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A1_c_130_n N_VPWR_c_289_n 0.00464324f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A1_c_131_n N_VPWR_c_289_n 0.0052046f $X=1.475 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A1_c_130_n N_VPWR_c_287_n 0.00525281f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A1_c_131_n N_VPWR_c_287_n 0.00687867f $X=1.475 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A1_c_130_n N_VPWR_c_294_n 0.00738999f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A1_c_131_n N_VPWR_c_294_n 0.00104319f $X=1.475 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A1_c_127_n N_Y_c_343_n 0.00946148f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A1_c_128_n N_Y_c_343_n 0.00980958f $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A1_c_126_n N_Y_c_350_n 0.0113796f $X=0.97 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A1_c_128_n N_Y_c_350_n 0.0236315f $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A1_c_129_n N_Y_c_350_n 0.0045174f $X=1.475 $Y=1.202 $X2=0 $Y2=0
cc_131 N_A1_c_126_n N_VGND_c_394_n 0.00526178f $X=0.97 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A1_c_127_n N_VGND_c_394_n 0.00422112f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A1_c_127_n N_VGND_c_396_n 0.00175799f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A1_c_126_n N_VGND_c_397_n 0.00964811f $X=0.97 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A1_c_127_n N_VGND_c_397_n 0.00591585f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_136 B1 N_A_27_297#_M1010_d 0.00744486f $X=3.08 $Y=1.105 $X2=0 $Y2=0
cc_137 N_B1_c_178_n N_A_27_297#_c_239_n 0.00277027f $X=2.415 $Y=1.41 $X2=0 $Y2=0
cc_138 N_B1_c_178_n N_A_27_297#_c_241_n 0.00408605f $X=2.415 $Y=1.41 $X2=0 $Y2=0
cc_139 N_B1_c_179_n N_A_27_297#_c_241_n 7.22416e-19 $X=2.885 $Y=1.41 $X2=0 $Y2=0
cc_140 N_B1_c_178_n N_A_27_297#_c_227_n 0.0133041f $X=2.415 $Y=1.41 $X2=0 $Y2=0
cc_141 N_B1_c_179_n N_A_27_297#_c_227_n 0.0165004f $X=2.885 $Y=1.41 $X2=0 $Y2=0
cc_142 B1 N_A_27_297#_c_227_n 0.00141565f $X=3.08 $Y=1.105 $X2=0 $Y2=0
cc_143 N_B1_c_178_n N_A_27_297#_c_242_n 4.8481e-19 $X=2.415 $Y=1.41 $X2=0 $Y2=0
cc_144 N_B1_c_179_n N_A_27_297#_c_228_n 0.0139373f $X=2.885 $Y=1.41 $X2=0 $Y2=0
cc_145 B1 N_A_27_297#_c_228_n 0.0272893f $X=3.08 $Y=1.105 $X2=0 $Y2=0
cc_146 N_B1_c_177_n N_A_27_297#_c_228_n 7.9185e-19 $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_147 N_B1_c_178_n N_VPWR_c_292_n 0.00429425f $X=2.415 $Y=1.41 $X2=0 $Y2=0
cc_148 N_B1_c_179_n N_VPWR_c_292_n 0.00429453f $X=2.885 $Y=1.41 $X2=0 $Y2=0
cc_149 N_B1_c_178_n N_VPWR_c_287_n 0.00609019f $X=2.415 $Y=1.41 $X2=0 $Y2=0
cc_150 N_B1_c_179_n N_VPWR_c_287_n 0.0072432f $X=2.885 $Y=1.41 $X2=0 $Y2=0
cc_151 N_B1_M1002_g N_Y_c_343_n 0.0102052f $X=2.39 $Y=0.56 $X2=0 $Y2=0
cc_152 N_B1_M1002_g N_Y_c_346_n 0.00682767f $X=2.39 $Y=0.56 $X2=0 $Y2=0
cc_153 N_B1_M1004_g N_Y_c_346_n 0.0109984f $X=2.86 $Y=0.56 $X2=0 $Y2=0
cc_154 N_B1_c_175_n N_Y_c_346_n 0.00955154f $X=2.985 $Y=1.16 $X2=0 $Y2=0
cc_155 B1 N_Y_c_346_n 0.0506466f $X=3.08 $Y=1.105 $X2=0 $Y2=0
cc_156 N_B1_c_178_n N_Y_c_342_n 9.14539e-19 $X=2.415 $Y=1.41 $X2=0 $Y2=0
cc_157 N_B1_c_179_n N_Y_c_342_n 0.0179927f $X=2.885 $Y=1.41 $X2=0 $Y2=0
cc_158 N_B1_c_175_n N_Y_c_342_n 0.00323496f $X=2.985 $Y=1.16 $X2=0 $Y2=0
cc_159 N_B1_M1002_g N_Y_c_364_n 0.00204408f $X=2.39 $Y=0.56 $X2=0 $Y2=0
cc_160 N_B1_M1004_g N_Y_c_364_n 0.00270876f $X=2.86 $Y=0.56 $X2=0 $Y2=0
cc_161 N_B1_c_175_n N_Y_c_366_n 0.0269209f $X=2.985 $Y=1.16 $X2=0 $Y2=0
cc_162 N_B1_M1004_g N_Y_c_367_n 0.00637454f $X=2.86 $Y=0.56 $X2=0 $Y2=0
cc_163 N_B1_M1004_g N_VGND_c_393_n 0.0161391f $X=2.86 $Y=0.56 $X2=0 $Y2=0
cc_164 B1 N_VGND_c_393_n 0.0300461f $X=3.08 $Y=1.105 $X2=0 $Y2=0
cc_165 N_B1_c_177_n N_VGND_c_393_n 0.00141736f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_166 N_B1_M1002_g N_VGND_c_395_n 0.00422057f $X=2.39 $Y=0.56 $X2=0 $Y2=0
cc_167 N_B1_M1004_g N_VGND_c_395_n 0.00465454f $X=2.86 $Y=0.56 $X2=0 $Y2=0
cc_168 N_B1_M1002_g N_VGND_c_396_n 0.00323317f $X=2.39 $Y=0.56 $X2=0 $Y2=0
cc_169 N_B1_M1002_g N_VGND_c_397_n 0.00595814f $X=2.39 $Y=0.56 $X2=0 $Y2=0
cc_170 N_B1_M1004_g N_VGND_c_397_n 0.00935497f $X=2.86 $Y=0.56 $X2=0 $Y2=0
cc_171 N_A_27_297#_c_234_n N_VPWR_M1000_d 0.00395992f $X=1.15 $Y=1.98 $X2=-0.19
+ $Y2=1.305
cc_172 N_A_27_297#_c_237_n N_VPWR_M1006_d 0.00362947f $X=2.015 $Y=1.94 $X2=0
+ $Y2=0
cc_173 N_A_27_297#_c_260_p N_VPWR_c_288_n 0.0127516f $X=1.235 $Y=2.3 $X2=0 $Y2=0
cc_174 N_A_27_297#_c_237_n N_VPWR_c_288_n 0.0130459f $X=2.015 $Y=1.94 $X2=0
+ $Y2=0
cc_175 N_A_27_297#_c_241_n N_VPWR_c_288_n 0.00541825f $X=2.18 $Y=2.285 $X2=0
+ $Y2=0
cc_176 N_A_27_297#_c_242_n N_VPWR_c_288_n 0.0115829f $X=2.345 $Y=2.375 $X2=0
+ $Y2=0
cc_177 N_A_27_297#_c_234_n N_VPWR_c_289_n 0.00362125f $X=1.15 $Y=1.98 $X2=0
+ $Y2=0
cc_178 N_A_27_297#_c_260_p N_VPWR_c_289_n 0.0117203f $X=1.235 $Y=2.3 $X2=0 $Y2=0
cc_179 N_A_27_297#_c_237_n N_VPWR_c_289_n 0.00367471f $X=2.015 $Y=1.94 $X2=0
+ $Y2=0
cc_180 N_A_27_297#_c_226_n N_VPWR_c_291_n 0.0179971f $X=0.275 $Y=2.3 $X2=0 $Y2=0
cc_181 N_A_27_297#_c_234_n N_VPWR_c_291_n 0.00258044f $X=1.15 $Y=1.98 $X2=0
+ $Y2=0
cc_182 N_A_27_297#_c_237_n N_VPWR_c_292_n 0.0027955f $X=2.015 $Y=1.94 $X2=0
+ $Y2=0
cc_183 N_A_27_297#_c_227_n N_VPWR_c_292_n 0.0630289f $X=3.085 $Y=2.375 $X2=0
+ $Y2=0
cc_184 N_A_27_297#_c_242_n N_VPWR_c_292_n 0.0189647f $X=2.345 $Y=2.375 $X2=0
+ $Y2=0
cc_185 N_A_27_297#_M1000_s N_VPWR_c_287_n 0.00251264f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_186 N_A_27_297#_M1001_s N_VPWR_c_287_n 0.00288166f $X=1.085 $Y=1.485 $X2=0
+ $Y2=0
cc_187 N_A_27_297#_M1011_s N_VPWR_c_287_n 0.00231261f $X=2.035 $Y=1.485 $X2=0
+ $Y2=0
cc_188 N_A_27_297#_M1010_d N_VPWR_c_287_n 0.0030031f $X=2.975 $Y=1.485 $X2=0
+ $Y2=0
cc_189 N_A_27_297#_c_226_n N_VPWR_c_287_n 0.00990273f $X=0.275 $Y=2.3 $X2=0
+ $Y2=0
cc_190 N_A_27_297#_c_234_n N_VPWR_c_287_n 0.0119994f $X=1.15 $Y=1.98 $X2=0 $Y2=0
cc_191 N_A_27_297#_c_260_p N_VPWR_c_287_n 0.00645162f $X=1.235 $Y=2.3 $X2=0
+ $Y2=0
cc_192 N_A_27_297#_c_237_n N_VPWR_c_287_n 0.0131151f $X=2.015 $Y=1.94 $X2=0
+ $Y2=0
cc_193 N_A_27_297#_c_227_n N_VPWR_c_287_n 0.0377824f $X=3.085 $Y=2.375 $X2=0
+ $Y2=0
cc_194 N_A_27_297#_c_242_n N_VPWR_c_287_n 0.0123455f $X=2.345 $Y=2.375 $X2=0
+ $Y2=0
cc_195 N_A_27_297#_c_234_n N_VPWR_c_294_n 0.0200578f $X=1.15 $Y=1.98 $X2=0 $Y2=0
cc_196 N_A_27_297#_c_260_p N_VPWR_c_294_n 0.01124f $X=1.235 $Y=2.3 $X2=0 $Y2=0
cc_197 N_A_27_297#_c_227_n N_Y_M1009_s 0.00353015f $X=3.085 $Y=2.375 $X2=0 $Y2=0
cc_198 N_A_27_297#_c_227_n N_Y_c_342_n 0.0184099f $X=3.085 $Y=2.375 $X2=0 $Y2=0
cc_199 N_A_27_297#_c_228_n N_Y_c_342_n 0.02034f $X=3.22 $Y=1.96 $X2=0 $Y2=0
cc_200 N_VPWR_c_287_n N_Y_M1009_s 0.00232895f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_201 N_Y_c_343_n N_VGND_M1007_d 0.00933387f $X=2.41 $Y=0.7 $X2=0 $Y2=0
cc_202 N_Y_c_350_n N_VGND_c_391_n 0.0150491f $X=1.235 $Y=0.36 $X2=0 $Y2=0
cc_203 N_Y_c_346_n N_VGND_c_393_n 0.00249031f $X=2.637 $Y=1.103 $X2=0 $Y2=0
cc_204 N_Y_c_364_n N_VGND_c_393_n 0.0110879f $X=2.65 $Y=0.76 $X2=0 $Y2=0
cc_205 N_Y_c_367_n N_VGND_c_393_n 0.0220779f $X=2.65 $Y=0.42 $X2=0 $Y2=0
cc_206 N_Y_c_343_n N_VGND_c_394_n 0.00790063f $X=2.41 $Y=0.7 $X2=0 $Y2=0
cc_207 N_Y_c_350_n N_VGND_c_394_n 0.0240714f $X=1.235 $Y=0.36 $X2=0 $Y2=0
cc_208 N_Y_c_343_n N_VGND_c_395_n 0.00188038f $X=2.41 $Y=0.7 $X2=0 $Y2=0
cc_209 N_Y_c_364_n N_VGND_c_395_n 0.0020837f $X=2.65 $Y=0.76 $X2=0 $Y2=0
cc_210 N_Y_c_367_n N_VGND_c_395_n 0.0201743f $X=2.65 $Y=0.42 $X2=0 $Y2=0
cc_211 N_Y_c_343_n N_VGND_c_396_n 0.0218271f $X=2.41 $Y=0.7 $X2=0 $Y2=0
cc_212 N_Y_M1008_s N_VGND_c_397_n 0.00310795f $X=1.045 $Y=0.235 $X2=0 $Y2=0
cc_213 N_Y_M1002_s N_VGND_c_397_n 0.00280994f $X=2.465 $Y=0.235 $X2=0 $Y2=0
cc_214 N_Y_c_343_n N_VGND_c_397_n 0.017943f $X=2.41 $Y=0.7 $X2=0 $Y2=0
cc_215 N_Y_c_350_n N_VGND_c_397_n 0.0147877f $X=1.235 $Y=0.36 $X2=0 $Y2=0
cc_216 N_Y_c_364_n N_VGND_c_397_n 0.00379118f $X=2.65 $Y=0.76 $X2=0 $Y2=0
cc_217 N_Y_c_367_n N_VGND_c_397_n 0.011813f $X=2.65 $Y=0.42 $X2=0 $Y2=0
cc_218 N_Y_c_343_n A_315_47# 0.00529826f $X=2.41 $Y=0.7 $X2=-0.19 $Y2=1.305
cc_219 N_VGND_c_397_n A_123_47# 0.0119688f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
cc_220 N_VGND_c_397_n A_315_47# 0.00239227f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
