* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nand2_2 A B VGND VNB VPB VPWR Y
M1000 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=8.3e+11p pd=7.66e+06u as=5.8e+11p ps=5.16e+06u
M1001 a_27_47# B VGND VNB nshort w=650000u l=150000u
+  ad=5.135e+11p pd=5.48e+06u as=2.405e+11p ps=2.04e+06u
M1002 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=2.405e+11p pd=2.04e+06u as=0p ps=0u
M1003 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
