* File: sky130_fd_sc_hdll__buf_1.pxi.spice
* Created: Wed Sep  2 08:24:09 2020
* 
x_PM_SKY130_FD_SC_HDLL__BUF_1%A N_A_c_39_n N_A_c_40_n N_A_M1000_g N_A_M1002_g A
+ N_A_c_38_n PM_SKY130_FD_SC_HDLL__BUF_1%A
x_PM_SKY130_FD_SC_HDLL__BUF_1%A_27_47# N_A_27_47#_M1002_s N_A_27_47#_M1000_s
+ N_A_27_47#_c_69_n N_A_27_47#_M1001_g N_A_27_47#_M1003_g N_A_27_47#_c_85_n
+ N_A_27_47#_c_120_p N_A_27_47#_c_71_n N_A_27_47#_c_72_n N_A_27_47#_c_76_n
+ N_A_27_47#_c_77_n N_A_27_47#_c_78_n N_A_27_47#_c_73_n N_A_27_47#_c_74_n
+ PM_SKY130_FD_SC_HDLL__BUF_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__BUF_1%VPWR N_VPWR_M1000_d N_VPWR_c_130_n VPWR VPWR
+ N_VPWR_c_131_n N_VPWR_c_132_n N_VPWR_c_129_n N_VPWR_c_134_n
+ PM_SKY130_FD_SC_HDLL__BUF_1%VPWR
x_PM_SKY130_FD_SC_HDLL__BUF_1%X N_X_M1003_d N_X_M1001_d N_X_c_154_n N_X_c_151_n
+ X X X N_X_c_153_n PM_SKY130_FD_SC_HDLL__BUF_1%X
x_PM_SKY130_FD_SC_HDLL__BUF_1%VGND N_VGND_M1002_d N_VGND_c_176_n VGND VGND
+ N_VGND_c_177_n VGND N_VGND_c_178_n N_VGND_c_179_n N_VGND_c_180_n
+ PM_SKY130_FD_SC_HDLL__BUF_1%VGND
cc_1 VNB N_A_M1002_g 0.0317693f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.495
cc_2 VNB A 0.0179991f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.105
cc_3 VNB N_A_c_38_n 0.0266942f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=1.16
cc_4 VNB N_A_27_47#_c_69_n 0.0184581f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.495
cc_5 VNB N_A_27_47#_M1003_g 0.0326284f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=1.16
cc_6 VNB N_A_27_47#_c_71_n 0.00556178f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_72_n 0.00375621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_73_n 0.00314921f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_74_n 0.00420848f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_VPWR_c_129_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_X_c_151_n 0.0256935f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.105
cc_12 VNB X 0.0136052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_X_c_153_n 0.0115694f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_VGND_c_176_n 0.00276307f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_15 VNB N_VGND_c_177_n 0.0154145f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=1.16
cc_16 VNB N_VGND_c_178_n 0.0290065f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_179_n 0.140082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_180_n 0.00560016f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VPB N_A_c_39_n 0.0164699f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.52
cc_20 VPB N_A_c_40_n 0.0263798f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.62
cc_21 VPB A 0.0064129f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.105
cc_22 VPB N_A_c_38_n 0.00348369f $X=-0.19 $Y=1.305 $X2=0.46 $Y2=1.16
cc_23 VPB N_A_27_47#_c_69_n 0.0427866f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.495
cc_24 VPB N_A_27_47#_c_76_n 0.00500472f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_25 VPB N_A_27_47#_c_77_n 0.00847174f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_26 VPB N_A_27_47#_c_78_n 0.0013355f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_A_27_47#_c_73_n 6.56842e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB N_VPWR_c_130_n 0.0028167f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_29 VPB N_VPWR_c_131_n 0.0161285f $X=-0.19 $Y=1.305 $X2=0.46 $Y2=1.16
cc_30 VPB N_VPWR_c_132_n 0.0290102f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_129_n 0.059866f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_134_n 0.00566735f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_X_c_154_n 0.0121424f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_X_c_151_n 0.011831f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.105
cc_35 VPB X 0.0292376f $X=-0.19 $Y=1.305 $X2=0.46 $Y2=1.16
cc_36 N_A_c_39_n N_A_27_47#_c_69_n 0.00935647f $X=0.495 $Y=1.52 $X2=0 $Y2=0
cc_37 N_A_c_40_n N_A_27_47#_c_69_n 0.0107646f $X=0.495 $Y=1.62 $X2=0 $Y2=0
cc_38 A N_A_27_47#_c_69_n 2.83759e-19 $X=0.305 $Y=1.105 $X2=0 $Y2=0
cc_39 N_A_c_38_n N_A_27_47#_c_69_n 0.0189172f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_40 N_A_M1002_g N_A_27_47#_M1003_g 0.023845f $X=0.52 $Y=0.495 $X2=0 $Y2=0
cc_41 N_A_c_40_n N_A_27_47#_c_85_n 0.00627093f $X=0.495 $Y=1.62 $X2=0 $Y2=0
cc_42 N_A_M1002_g N_A_27_47#_c_71_n 0.0138654f $X=0.52 $Y=0.495 $X2=0 $Y2=0
cc_43 A N_A_27_47#_c_71_n 0.0145322f $X=0.305 $Y=1.105 $X2=0 $Y2=0
cc_44 N_A_c_38_n N_A_27_47#_c_71_n 6.71548e-19 $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_45 A N_A_27_47#_c_72_n 0.0143235f $X=0.305 $Y=1.105 $X2=0 $Y2=0
cc_46 N_A_c_40_n N_A_27_47#_c_76_n 0.018909f $X=0.495 $Y=1.62 $X2=0 $Y2=0
cc_47 A N_A_27_47#_c_76_n 0.0141328f $X=0.305 $Y=1.105 $X2=0 $Y2=0
cc_48 N_A_c_38_n N_A_27_47#_c_76_n 3.19113e-19 $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_49 A N_A_27_47#_c_77_n 0.0154163f $X=0.305 $Y=1.105 $X2=0 $Y2=0
cc_50 N_A_c_39_n N_A_27_47#_c_78_n 0.00348557f $X=0.495 $Y=1.52 $X2=0 $Y2=0
cc_51 N_A_c_38_n N_A_27_47#_c_73_n 0.00348557f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_52 N_A_M1002_g N_A_27_47#_c_74_n 0.00348557f $X=0.52 $Y=0.495 $X2=0 $Y2=0
cc_53 A N_A_27_47#_c_74_n 0.0287477f $X=0.305 $Y=1.105 $X2=0 $Y2=0
cc_54 N_A_c_40_n N_VPWR_c_130_n 0.0157173f $X=0.495 $Y=1.62 $X2=0 $Y2=0
cc_55 N_A_c_40_n N_VPWR_c_131_n 0.0046653f $X=0.495 $Y=1.62 $X2=0 $Y2=0
cc_56 N_A_c_40_n N_VPWR_c_129_n 0.00885548f $X=0.495 $Y=1.62 $X2=0 $Y2=0
cc_57 N_A_c_40_n N_X_c_154_n 6.23649e-19 $X=0.495 $Y=1.62 $X2=0 $Y2=0
cc_58 N_A_M1002_g X 5.4697e-19 $X=0.52 $Y=0.495 $X2=0 $Y2=0
cc_59 N_A_M1002_g N_VGND_c_176_n 0.0107485f $X=0.52 $Y=0.495 $X2=0 $Y2=0
cc_60 N_A_M1002_g N_VGND_c_177_n 0.00226008f $X=0.52 $Y=0.495 $X2=0 $Y2=0
cc_61 N_A_M1002_g N_VGND_c_179_n 0.00393085f $X=0.52 $Y=0.495 $X2=0 $Y2=0
cc_62 N_A_27_47#_c_76_n N_VPWR_M1000_d 0.00212434f $X=0.72 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_63 N_A_27_47#_c_69_n N_VPWR_c_130_n 0.00345026f $X=0.985 $Y=1.62 $X2=0 $Y2=0
cc_64 N_A_27_47#_c_85_n N_VPWR_c_130_n 0.0422302f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_65 N_A_27_47#_c_76_n N_VPWR_c_130_n 0.0214008f $X=0.72 $Y=1.62 $X2=0 $Y2=0
cc_66 N_A_27_47#_c_85_n N_VPWR_c_131_n 0.0125171f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_67 N_A_27_47#_c_69_n N_VPWR_c_132_n 0.00687021f $X=0.985 $Y=1.62 $X2=0 $Y2=0
cc_68 N_A_27_47#_M1000_s N_VPWR_c_129_n 0.0053343f $X=0.135 $Y=1.695 $X2=0 $Y2=0
cc_69 N_A_27_47#_c_69_n N_VPWR_c_129_n 0.0134108f $X=0.985 $Y=1.62 $X2=0 $Y2=0
cc_70 N_A_27_47#_c_85_n N_VPWR_c_129_n 0.00685509f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_71 N_A_27_47#_c_69_n N_X_c_154_n 0.00618152f $X=0.985 $Y=1.62 $X2=0 $Y2=0
cc_72 N_A_27_47#_c_76_n N_X_c_154_n 0.0111516f $X=0.72 $Y=1.62 $X2=0 $Y2=0
cc_73 N_A_27_47#_M1003_g N_X_c_151_n 0.0157458f $X=1.01 $Y=0.495 $X2=0 $Y2=0
cc_74 N_A_27_47#_c_78_n N_X_c_151_n 0.00530245f $X=0.805 $Y=1.535 $X2=0 $Y2=0
cc_75 N_A_27_47#_c_73_n N_X_c_151_n 0.0237746f $X=0.95 $Y=1.225 $X2=0 $Y2=0
cc_76 N_A_27_47#_c_74_n N_X_c_151_n 0.0120117f $X=0.877 $Y=1.06 $X2=0 $Y2=0
cc_77 N_A_27_47#_M1003_g X 0.006285f $X=1.01 $Y=0.495 $X2=0 $Y2=0
cc_78 N_A_27_47#_c_69_n X 0.0088978f $X=0.985 $Y=1.62 $X2=0 $Y2=0
cc_79 N_A_27_47#_M1003_g N_X_c_153_n 0.00357209f $X=1.01 $Y=0.495 $X2=0 $Y2=0
cc_80 N_A_27_47#_c_71_n N_X_c_153_n 0.00478763f $X=0.72 $Y=0.72 $X2=0 $Y2=0
cc_81 N_A_27_47#_c_71_n N_VGND_M1002_d 0.00305131f $X=0.72 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_82 N_A_27_47#_c_69_n N_VGND_c_176_n 2.27088e-19 $X=0.985 $Y=1.62 $X2=0 $Y2=0
cc_83 N_A_27_47#_M1003_g N_VGND_c_176_n 0.00425261f $X=1.01 $Y=0.495 $X2=0 $Y2=0
cc_84 N_A_27_47#_c_120_p N_VGND_c_176_n 0.0149682f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_85 N_A_27_47#_c_71_n N_VGND_c_176_n 0.0233571f $X=0.72 $Y=0.72 $X2=0 $Y2=0
cc_86 N_A_27_47#_c_120_p N_VGND_c_177_n 0.0116326f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_87 N_A_27_47#_c_71_n N_VGND_c_177_n 0.00259539f $X=0.72 $Y=0.72 $X2=0 $Y2=0
cc_88 N_A_27_47#_M1003_g N_VGND_c_178_n 0.0055654f $X=1.01 $Y=0.495 $X2=0 $Y2=0
cc_89 N_A_27_47#_M1002_s N_VGND_c_179_n 0.00431832f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_90 N_A_27_47#_M1003_g N_VGND_c_179_n 0.011535f $X=1.01 $Y=0.495 $X2=0 $Y2=0
cc_91 N_A_27_47#_c_120_p N_VGND_c_179_n 0.00643448f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_71_n N_VGND_c_179_n 0.00640917f $X=0.72 $Y=0.72 $X2=0 $Y2=0
cc_93 N_VPWR_c_129_n N_X_M1001_d 0.00217517f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_94 N_VPWR_c_130_n X 0.0471129f $X=0.73 $Y=1.96 $X2=0 $Y2=0
cc_95 N_VPWR_c_132_n X 0.0210947f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_96 N_VPWR_c_129_n X 0.0125182f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_97 X N_VGND_c_178_n 0.0209687f $X=1.155 $Y=0.425 $X2=0 $Y2=0
cc_98 N_X_M1003_d N_VGND_c_179_n 0.00210122f $X=1.085 $Y=0.235 $X2=0 $Y2=0
cc_99 X N_VGND_c_179_n 0.0125012f $X=1.155 $Y=0.425 $X2=0 $Y2=0
