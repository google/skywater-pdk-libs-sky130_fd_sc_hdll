* File: sky130_fd_sc_hdll__mux2i_1.spice
* Created: Thu Aug 27 19:11:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__mux2i_1.pex.spice"
.subckt sky130_fd_sc_hdll__mux2i_1  VNB VPB A0 A1 S Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* S	S
* A1	A1
* A0	A0
* VPB	VPB
* VNB	VNB
MM1005 N_Y_M1005_d N_A0_M1005_g N_A_27_47#_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.2145 PD=0.92 PS=1.96 NRD=0 NRS=11.988 M=1 R=4.33333 SA=75000.3
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1002 N_A_207_47#_M1002_d N_A1_M1002_g N_Y_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A_303_205#_M1008_g N_A_27_47#_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1009 N_A_207_47#_M1009_d N_S_M1009_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1885 AS=0.08775 PD=1.88 PS=0.92 NRD=4.608 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_S_M1003_g N_A_303_205#_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.2275 PD=1.82 PS=2 NRD=0 NRS=11.988 M=1 R=4.33333 SA=75000.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_Y_M1000_d N_A0_M1000_g N_A_27_297#_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002 A=0.18 P=2.36 MULT=1
MM1007 A_215_297# N_A1_M1007_g N_Y_M1000_d VPB PHIGHVT L=0.18 W=1 AD=0.225
+ AS=0.145 PD=1.45 PS=1.29 NRD=33.4703 NRS=0.9653 M=1 R=5.55556 SA=90000.7
+ SB=90001.5 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A_303_205#_M1006_g A_215_297# VPB PHIGHVT L=0.18 W=1
+ AD=0.275 AS=0.225 PD=1.55 PS=1.45 NRD=26.5753 NRS=33.4703 M=1 R=5.55556
+ SA=90001.3 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1001 N_A_27_297#_M1001_d N_S_M1001_g N_VPWR_M1006_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.275 PD=2.54 PS=1.55 NRD=0.9653 NRS=26.5753 M=1 R=5.55556 SA=90002
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_S_M1004_g N_A_303_205#_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.3 PD=2.54 PS=2.6 NRD=0.9653 NRS=4.9053 M=1 R=5.55556 SA=90000.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.2546 P=12.25
c_63 VPB 0 1.72057e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__mux2i_1.pxi.spice"
*
.ends
*
*
