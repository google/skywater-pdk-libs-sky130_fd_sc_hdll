# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__or4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.815000 0.995000 3.570000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.680000 2.125000 3.370000 2.455000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.810000 1.695000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.980000 0.995000 1.335000 1.325000 ;
    END
  END D_N
  PIN VGND
    ANTENNADIFFAREA  0.620550 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  0.564325 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  0.463750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.130000 0.415000 4.455000 0.760000 ;
        RECT 4.130000 1.495000 4.455000 2.465000 ;
        RECT 4.235000 0.760000 4.455000 1.495000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.450000 0.400000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.865000 ;
      RECT 0.085000  1.865000 2.015000 2.035000 ;
      RECT 0.085000  2.035000 0.345000 2.455000 ;
      RECT 0.515000  2.205000 0.895000 2.635000 ;
      RECT 0.705000  0.085000 0.875000 0.825000 ;
      RECT 1.040000  1.525000 1.675000 1.695000 ;
      RECT 1.175000  0.450000 1.345000 0.655000 ;
      RECT 1.175000  0.655000 1.675000 0.825000 ;
      RECT 1.505000  0.825000 1.675000 1.075000 ;
      RECT 1.505000  1.075000 2.155000 1.245000 ;
      RECT 1.505000  1.245000 1.675000 1.525000 ;
      RECT 1.570000  0.085000 1.945000 0.485000 ;
      RECT 1.610000  2.205000 2.405000 2.375000 ;
      RECT 1.845000  1.415000 2.545000 1.585000 ;
      RECT 1.845000  1.585000 2.015000 1.865000 ;
      RECT 2.165000  0.305000 2.335000 0.655000 ;
      RECT 2.165000  0.655000 3.910000 0.825000 ;
      RECT 2.235000  1.785000 3.370000 1.955000 ;
      RECT 2.235000  1.955000 2.405000 2.205000 ;
      RECT 2.375000  0.995000 2.545000 1.415000 ;
      RECT 2.520000  0.085000 2.900000 0.485000 ;
      RECT 3.120000  0.305000 3.290000 0.655000 ;
      RECT 3.200000  1.495000 3.910000 1.665000 ;
      RECT 3.200000  1.665000 3.370000 1.785000 ;
      RECT 3.460000  0.085000 3.890000 0.485000 ;
      RECT 3.590000  1.835000 3.870000 2.635000 ;
      RECT 3.740000  0.825000 3.910000 0.995000 ;
      RECT 3.740000  0.995000 4.030000 1.325000 ;
      RECT 3.740000  1.325000 3.910000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4bb_1
END LIBRARY
