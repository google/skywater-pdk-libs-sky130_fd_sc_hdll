* File: sky130_fd_sc_hdll__nand3_1.spice
* Created: Wed Sep  2 08:37:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nand3_1.pex.spice"
.subckt sky130_fd_sc_hdll__nand3_1  VNB VPB C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1005 A_119_47# N_C_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.2015 PD=0.92 PS=1.92 NRD=14.76 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1001 A_203_47# N_B_M1001_g A_119_47# VNB NSHORT L=0.15 W=0.65 AD=0.1235
+ AS=0.08775 PD=1.03 PS=0.92 NRD=24.912 NRS=14.76 M=1 R=4.33333 SA=75000.7
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g A_203_47# VNB NSHORT L=0.15 W=0.65 AD=0.2015
+ AS=0.1235 PD=1.92 PS=1.03 NRD=8.304 NRS=24.912 M=1 R=4.33333 SA=75001.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_Y_M1003_d N_C_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_B_M1000_g N_Y_M1003_d VPB PHIGHVT L=0.18 W=1 AD=0.175
+ AS=0.145 PD=1.35 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.6
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g N_VPWR_M1000_d VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.175 PD=2.54 PS=1.35 NRD=0.9653 NRS=12.7853 M=1 R=5.55556 SA=90001.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
*
.include "sky130_fd_sc_hdll__nand3_1.pxi.spice"
*
.ends
*
*
