* File: sky130_fd_sc_hdll__nor3b_1.spice
* Created: Wed Sep  2 08:40:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nor3b_1.pex.spice"
.subckt sky130_fd_sc_hdll__nor3b_1  VNB VPB B A C_N Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* C_N	C_N
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_91_199#_M1005_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.2535 PD=0.97 PS=2.08 NRD=0 NRS=23.076 M=1 R=4.33333 SA=75000.3
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_B_M1004_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.8
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A_M1006_g N_Y_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.154299 AS=0.08775 PD=1.31822 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1000 N_A_91_199#_M1000_d N_C_N_M1000_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0997009 PD=1.36 PS=0.851776 NRD=0 NRS=32.136 M=1 R=2.8
+ SA=75001.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_169_297# N_A_91_199#_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.33 PD=1.29 PS=2.66 NRD=17.7103 NRS=12.7853 M=1 R=5.55556
+ SA=90000.2 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1001 A_263_297# N_B_M1001_g A_169_297# VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=17.7103 NRS=17.7103 M=1 R=5.55556 SA=90000.7
+ SB=90000.9 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g A_263_297# VPB PHIGHVT L=0.18 W=1 AD=0.215282
+ AS=0.145 PD=1.90845 PS=1.29 NRD=0.9653 NRS=17.7103 M=1 R=5.55556 SA=90001.2
+ SB=90000.4 A=0.18 P=2.36 MULT=1
MM1003 N_A_91_199#_M1003_d N_C_N_M1003_g N_VPWR_M1007_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.0904183 PD=1.38 PS=0.801549 NRD=2.3443 NRS=75.1752 M=1
+ R=2.33333 SA=90001.7 SB=90000.2 A=0.0756 P=1.2 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
pX9_noxref noxref_12 A A PROBETYPE=1
*
.include "sky130_fd_sc_hdll__nor3b_1.pxi.spice"
*
.ends
*
*
