* File: sky130_fd_sc_hdll__a21bo_1.pxi.spice
* Created: Thu Aug 27 18:52:03 2020
* 
x_PM_SKY130_FD_SC_HDLL__A21BO_1%B1_N N_B1_N_c_62_n N_B1_N_c_63_n N_B1_N_c_67_n
+ N_B1_N_M1002_g N_B1_N_c_64_n N_B1_N_M1004_g N_B1_N_c_68_n B1_N B1_N B1_N B1_N
+ N_B1_N_c_66_n PM_SKY130_FD_SC_HDLL__A21BO_1%B1_N
x_PM_SKY130_FD_SC_HDLL__A21BO_1%A_27_413# N_A_27_413#_M1004_s
+ N_A_27_413#_M1002_s N_A_27_413#_c_99_n N_A_27_413#_c_106_n N_A_27_413#_M1008_g
+ N_A_27_413#_M1003_g N_A_27_413#_c_101_n N_A_27_413#_c_108_n
+ N_A_27_413#_c_102_n N_A_27_413#_c_109_n N_A_27_413#_c_103_n
+ N_A_27_413#_c_104_n PM_SKY130_FD_SC_HDLL__A21BO_1%A_27_413#
x_PM_SKY130_FD_SC_HDLL__A21BO_1%A1 N_A1_c_166_n N_A1_M1001_g N_A1_c_167_n
+ N_A1_M1007_g A1 A1 PM_SKY130_FD_SC_HDLL__A21BO_1%A1
x_PM_SKY130_FD_SC_HDLL__A21BO_1%A2 N_A2_c_201_n N_A2_M1006_g N_A2_c_202_n
+ N_A2_M1000_g A2 A2 PM_SKY130_FD_SC_HDLL__A21BO_1%A2
x_PM_SKY130_FD_SC_HDLL__A21BO_1%A_235_297# N_A_235_297#_M1003_d
+ N_A_235_297#_M1008_s N_A_235_297#_c_231_n N_A_235_297#_M1009_g
+ N_A_235_297#_c_232_n N_A_235_297#_M1005_g N_A_235_297#_c_237_n
+ N_A_235_297#_c_233_n N_A_235_297#_c_261_n N_A_235_297#_c_234_n
+ N_A_235_297#_c_235_n N_A_235_297#_c_256_n
+ PM_SKY130_FD_SC_HDLL__A21BO_1%A_235_297#
x_PM_SKY130_FD_SC_HDLL__A21BO_1%VPWR N_VPWR_M1002_d N_VPWR_M1007_d
+ N_VPWR_M1009_s N_VPWR_c_304_n N_VPWR_c_305_n N_VPWR_c_306_n N_VPWR_c_307_n
+ N_VPWR_c_308_n VPWR N_VPWR_c_309_n N_VPWR_c_310_n N_VPWR_c_311_n
+ N_VPWR_c_303_n N_VPWR_c_313_n N_VPWR_c_314_n
+ PM_SKY130_FD_SC_HDLL__A21BO_1%VPWR
x_PM_SKY130_FD_SC_HDLL__A21BO_1%A_326_297# N_A_326_297#_M1008_d
+ N_A_326_297#_M1000_d N_A_326_297#_c_364_n N_A_326_297#_c_370_n
+ N_A_326_297#_c_369_n PM_SKY130_FD_SC_HDLL__A21BO_1%A_326_297#
x_PM_SKY130_FD_SC_HDLL__A21BO_1%X N_X_M1005_d N_X_M1009_d X X X X X X
+ PM_SKY130_FD_SC_HDLL__A21BO_1%X
x_PM_SKY130_FD_SC_HDLL__A21BO_1%VGND N_VGND_M1004_d N_VGND_M1006_d
+ N_VGND_c_397_n VGND N_VGND_c_398_n N_VGND_c_399_n N_VGND_c_400_n
+ N_VGND_c_401_n N_VGND_c_402_n N_VGND_c_403_n
+ PM_SKY130_FD_SC_HDLL__A21BO_1%VGND
cc_1 VNB N_B1_N_c_62_n 0.0415819f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=0.83
cc_2 VNB N_B1_N_c_63_n 0.0206114f $X=-0.19 $Y=-0.24 $X2=0.375 $Y2=0.83
cc_3 VNB N_B1_N_c_64_n 0.021468f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=0.755
cc_4 VNB B1_N 0.0223982f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.425
cc_5 VNB N_B1_N_c_66_n 0.0388369f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_6 VNB N_A_27_413#_c_99_n 0.0196424f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=0.445
cc_7 VNB N_A_27_413#_M1003_g 0.028759f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_8 VNB N_A_27_413#_c_101_n 0.00552114f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_9 VNB N_A_27_413#_c_102_n 0.00594942f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_10 VNB N_A_27_413#_c_103_n 0.00385036f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_413#_c_104_n 0.0100652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A1_c_166_n 0.0170109f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=0.83
cc_13 VNB N_A1_c_167_n 0.0194605f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_14 VNB A1 0.00594606f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=0.445
cc_15 VNB N_A2_c_201_n 0.0227665f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=0.83
cc_16 VNB N_A2_c_202_n 0.0248506f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_17 VNB A2 0.00534236f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=0.445
cc_18 VNB N_A_235_297#_c_231_n 0.0266449f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=0.445
cc_19 VNB N_A_235_297#_c_232_n 0.023154f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.902
cc_20 VNB N_A_235_297#_c_233_n 0.00434152f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_235_297#_c_234_n 0.00777387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_235_297#_c_235_n 0.0113775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_303_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB X 0.0457123f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=0.445
cc_25 VNB N_VGND_c_397_n 0.00726972f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=0.905
cc_26 VNB N_VGND_c_398_n 0.0309477f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_27 VNB N_VGND_c_399_n 0.0238369f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_400_n 0.226103f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.53
cc_29 VNB N_VGND_c_401_n 0.00471252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_402_n 0.0347596f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_403_n 0.021931f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_B1_N_c_67_n 0.0217834f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_33 VPB N_B1_N_c_68_n 0.0376976f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.815
cc_34 VPB N_B1_N_c_66_n 0.0498728f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_35 VPB N_A_27_413#_c_99_n 0.0197919f $X=-0.19 $Y=1.305 $X2=0.865 $Y2=0.445
cc_36 VPB N_A_27_413#_c_106_n 0.0191189f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=0.905
cc_37 VPB N_A_27_413#_c_101_n 0.00531579f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_38 VPB N_A_27_413#_c_108_n 0.0151468f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_413#_c_109_n 0.0271708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_413#_c_103_n 5.81433e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_413#_c_104_n 0.0205145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A1_c_167_n 0.0229547f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_43 VPB A1 0.00256806f $X=-0.19 $Y=1.305 $X2=0.865 $Y2=0.445
cc_44 VPB N_A2_c_202_n 0.0296209f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_45 VPB A2 0.00276991f $X=-0.19 $Y=1.305 $X2=0.865 $Y2=0.445
cc_46 VPB N_A_235_297#_c_231_n 0.0339304f $X=-0.19 $Y=1.305 $X2=0.865 $Y2=0.445
cc_47 VPB N_A_235_297#_c_237_n 0.0112798f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_48 VPB N_A_235_297#_c_234_n 0.00199182f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_235_297#_c_235_n 0.00251691f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_304_n 0.00640047f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.902
cc_51 VPB N_VPWR_c_305_n 4.20076e-19 $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_52 VPB N_VPWR_c_306_n 0.0179977f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_307_n 0.0175141f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_308_n 0.00545601f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_309_n 0.014663f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.16
cc_56 VPB N_VPWR_c_310_n 0.0290331f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_311_n 0.0243997f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_303_n 0.0639438f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_313_n 0.00618204f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_314_n 0.00503278f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB X 0.0469905f $X=-0.19 $Y=1.305 $X2=0.865 $Y2=0.445
cc_62 N_B1_N_c_64_n N_A_27_413#_M1003_g 0.0127677f $X=0.865 $Y=0.755 $X2=0 $Y2=0
cc_63 N_B1_N_c_67_n N_A_27_413#_c_108_n 0.00503067f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_64 N_B1_N_c_68_n N_A_27_413#_c_108_n 0.00171886f $X=0.24 $Y=1.815 $X2=0 $Y2=0
cc_65 N_B1_N_c_62_n N_A_27_413#_c_102_n 0.0198067f $X=0.79 $Y=0.83 $X2=0 $Y2=0
cc_66 N_B1_N_c_64_n N_A_27_413#_c_102_n 0.00755763f $X=0.865 $Y=0.755 $X2=0
+ $Y2=0
cc_67 B1_N N_A_27_413#_c_102_n 0.099627f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_68 N_B1_N_c_66_n N_A_27_413#_c_102_n 0.0129125f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_69 N_B1_N_c_67_n N_A_27_413#_c_109_n 0.00670118f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_70 N_B1_N_c_68_n N_A_27_413#_c_109_n 0.0311722f $X=0.24 $Y=1.815 $X2=0 $Y2=0
cc_71 B1_N N_A_27_413#_c_109_n 0.016773f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_72 N_B1_N_c_62_n N_A_27_413#_c_103_n 0.00372807f $X=0.79 $Y=0.83 $X2=0 $Y2=0
cc_73 N_B1_N_c_62_n N_A_27_413#_c_104_n 0.0103536f $X=0.79 $Y=0.83 $X2=0 $Y2=0
cc_74 B1_N N_A_27_413#_c_104_n 2.94496e-19 $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_75 N_B1_N_c_66_n N_A_27_413#_c_104_n 0.010691f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_76 N_B1_N_c_67_n N_A_235_297#_c_237_n 0.00383723f $X=0.495 $Y=1.99 $X2=0
+ $Y2=0
cc_77 N_B1_N_c_68_n N_A_235_297#_c_237_n 5.92587e-19 $X=0.24 $Y=1.815 $X2=0
+ $Y2=0
cc_78 N_B1_N_c_62_n N_A_235_297#_c_233_n 2.66874e-19 $X=0.79 $Y=0.83 $X2=0 $Y2=0
cc_79 N_B1_N_c_67_n N_VPWR_c_304_n 0.0135794f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_80 N_B1_N_c_67_n N_VPWR_c_309_n 0.00315243f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_81 N_B1_N_c_68_n N_VPWR_c_309_n 3.38344e-19 $X=0.24 $Y=1.815 $X2=0 $Y2=0
cc_82 N_B1_N_c_67_n N_VPWR_c_303_n 0.00477468f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_83 N_B1_N_c_64_n N_VGND_c_397_n 0.0102408f $X=0.865 $Y=0.755 $X2=0 $Y2=0
cc_84 N_B1_N_c_62_n N_VGND_c_398_n 6.22378e-19 $X=0.79 $Y=0.83 $X2=0 $Y2=0
cc_85 N_B1_N_c_63_n N_VGND_c_398_n 0.00357448f $X=0.375 $Y=0.83 $X2=0 $Y2=0
cc_86 N_B1_N_c_64_n N_VGND_c_398_n 0.00579368f $X=0.865 $Y=0.755 $X2=0 $Y2=0
cc_87 B1_N N_VGND_c_398_n 0.0113151f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_88 N_B1_N_c_63_n N_VGND_c_400_n 0.00411268f $X=0.375 $Y=0.83 $X2=0 $Y2=0
cc_89 N_B1_N_c_64_n N_VGND_c_400_n 0.0125963f $X=0.865 $Y=0.755 $X2=0 $Y2=0
cc_90 B1_N N_VGND_c_400_n 0.00846606f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_91 N_A_27_413#_M1003_g N_A1_c_166_n 0.0155617f $X=1.565 $Y=0.56 $X2=-0.19
+ $Y2=-0.24
cc_92 N_A_27_413#_c_106_n N_A1_c_167_n 0.0208939f $X=1.54 $Y=1.41 $X2=0 $Y2=0
cc_93 N_A_27_413#_c_101_n N_A1_c_167_n 0.0155617f $X=1.54 $Y=1.297 $X2=0 $Y2=0
cc_94 N_A_27_413#_c_106_n A1 9.77397e-19 $X=1.54 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A_27_413#_M1003_g A1 9.95408e-19 $X=1.565 $Y=0.56 $X2=0 $Y2=0
cc_96 N_A_27_413#_c_101_n A1 5.83568e-19 $X=1.54 $Y=1.297 $X2=0 $Y2=0
cc_97 N_A_27_413#_c_99_n N_A_235_297#_c_237_n 0.0100166f $X=1.44 $Y=1.285 $X2=0
+ $Y2=0
cc_98 N_A_27_413#_c_106_n N_A_235_297#_c_237_n 0.0150761f $X=1.54 $Y=1.41 $X2=0
+ $Y2=0
cc_99 N_A_27_413#_c_101_n N_A_235_297#_c_237_n 0.00177768f $X=1.54 $Y=1.297
+ $X2=0 $Y2=0
cc_100 N_A_27_413#_c_109_n N_A_235_297#_c_237_n 0.0175151f $X=0.74 $Y=1.845
+ $X2=0 $Y2=0
cc_101 N_A_27_413#_c_103_n N_A_235_297#_c_237_n 0.0416984f $X=0.85 $Y=1.35 $X2=0
+ $Y2=0
cc_102 N_A_27_413#_c_104_n N_A_235_297#_c_237_n 0.0011422f $X=0.85 $Y=1.285
+ $X2=0 $Y2=0
cc_103 N_A_27_413#_M1003_g N_A_235_297#_c_233_n 0.00742211f $X=1.565 $Y=0.56
+ $X2=0 $Y2=0
cc_104 N_A_27_413#_c_102_n N_A_235_297#_c_233_n 0.00513721f $X=0.6 $Y=0.45 $X2=0
+ $Y2=0
cc_105 N_A_27_413#_c_99_n N_A_235_297#_c_235_n 0.0130044f $X=1.44 $Y=1.285 $X2=0
+ $Y2=0
cc_106 N_A_27_413#_M1003_g N_A_235_297#_c_235_n 0.00607897f $X=1.565 $Y=0.56
+ $X2=0 $Y2=0
cc_107 N_A_27_413#_c_101_n N_A_235_297#_c_235_n 0.0130528f $X=1.54 $Y=1.297
+ $X2=0 $Y2=0
cc_108 N_A_27_413#_c_102_n N_A_235_297#_c_235_n 0.00633431f $X=0.6 $Y=0.45 $X2=0
+ $Y2=0
cc_109 N_A_27_413#_c_103_n N_A_235_297#_c_235_n 0.0146395f $X=0.85 $Y=1.35 $X2=0
+ $Y2=0
cc_110 N_A_27_413#_M1003_g N_A_235_297#_c_256_n 0.0138831f $X=1.565 $Y=0.56
+ $X2=0 $Y2=0
cc_111 N_A_27_413#_c_106_n N_VPWR_c_304_n 0.0023773f $X=1.54 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A_27_413#_c_108_n N_VPWR_c_304_n 0.0161453f $X=0.26 $Y=2.27 $X2=0 $Y2=0
cc_113 N_A_27_413#_c_109_n N_VPWR_c_304_n 0.0272795f $X=0.74 $Y=1.845 $X2=0
+ $Y2=0
cc_114 N_A_27_413#_c_106_n N_VPWR_c_305_n 0.00120762f $X=1.54 $Y=1.41 $X2=0
+ $Y2=0
cc_115 N_A_27_413#_c_108_n N_VPWR_c_309_n 0.0135192f $X=0.26 $Y=2.27 $X2=0 $Y2=0
cc_116 N_A_27_413#_c_109_n N_VPWR_c_309_n 0.00270664f $X=0.74 $Y=1.845 $X2=0
+ $Y2=0
cc_117 N_A_27_413#_c_106_n N_VPWR_c_310_n 0.00681403f $X=1.54 $Y=1.41 $X2=0
+ $Y2=0
cc_118 N_A_27_413#_c_109_n N_VPWR_c_310_n 8.42227e-19 $X=0.74 $Y=1.845 $X2=0
+ $Y2=0
cc_119 N_A_27_413#_M1002_s N_VPWR_c_303_n 0.00245295f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_120 N_A_27_413#_c_106_n N_VPWR_c_303_n 0.0134342f $X=1.54 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_27_413#_c_108_n N_VPWR_c_303_n 0.0088929f $X=0.26 $Y=2.27 $X2=0 $Y2=0
cc_122 N_A_27_413#_c_109_n N_VPWR_c_303_n 0.00734704f $X=0.74 $Y=1.845 $X2=0
+ $Y2=0
cc_123 N_A_27_413#_c_99_n N_VGND_c_397_n 0.00408228f $X=1.44 $Y=1.285 $X2=0
+ $Y2=0
cc_124 N_A_27_413#_M1003_g N_VGND_c_397_n 0.00529755f $X=1.565 $Y=0.56 $X2=0
+ $Y2=0
cc_125 N_A_27_413#_c_102_n N_VGND_c_397_n 0.0337402f $X=0.6 $Y=0.45 $X2=0 $Y2=0
cc_126 N_A_27_413#_c_102_n N_VGND_c_398_n 0.0164742f $X=0.6 $Y=0.45 $X2=0 $Y2=0
cc_127 N_A_27_413#_M1004_s N_VGND_c_400_n 0.00303425f $X=0.475 $Y=0.235 $X2=0
+ $Y2=0
cc_128 N_A_27_413#_M1003_g N_VGND_c_400_n 0.00584613f $X=1.565 $Y=0.56 $X2=0
+ $Y2=0
cc_129 N_A_27_413#_c_102_n N_VGND_c_400_n 0.0106271f $X=0.6 $Y=0.45 $X2=0 $Y2=0
cc_130 N_A_27_413#_M1003_g N_VGND_c_402_n 0.00359757f $X=1.565 $Y=0.56 $X2=0
+ $Y2=0
cc_131 N_A1_c_166_n N_A2_c_201_n 0.0337816f $X=1.985 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_132 N_A1_c_167_n N_A2_c_202_n 0.0577418f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_133 A1 N_A2_c_202_n 0.00406308f $X=1.96 $Y=1.105 $X2=0 $Y2=0
cc_134 N_A1_c_167_n A2 5.75391e-19 $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_135 A1 A2 0.0484944f $X=1.96 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A1_c_167_n N_A_235_297#_c_237_n 9.85492e-19 $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_137 A1 N_A_235_297#_c_237_n 0.00779391f $X=1.96 $Y=1.105 $X2=0 $Y2=0
cc_138 N_A1_c_166_n N_A_235_297#_c_233_n 0.00376119f $X=1.985 $Y=0.995 $X2=0
+ $Y2=0
cc_139 A1 N_A_235_297#_c_233_n 0.00414057f $X=1.96 $Y=1.105 $X2=0 $Y2=0
cc_140 N_A1_c_166_n N_A_235_297#_c_261_n 0.00959075f $X=1.985 $Y=0.995 $X2=0
+ $Y2=0
cc_141 N_A1_c_167_n N_A_235_297#_c_261_n 7.06693e-19 $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_142 A1 N_A_235_297#_c_261_n 0.0232212f $X=1.96 $Y=1.105 $X2=0 $Y2=0
cc_143 N_A1_c_167_n N_A_235_297#_c_235_n 0.00112086f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_144 A1 N_A_235_297#_c_235_n 0.0263202f $X=1.96 $Y=1.105 $X2=0 $Y2=0
cc_145 N_A1_c_166_n N_A_235_297#_c_256_n 0.00900002f $X=1.985 $Y=0.995 $X2=0
+ $Y2=0
cc_146 A1 N_A_235_297#_c_256_n 0.00265009f $X=1.96 $Y=1.105 $X2=0 $Y2=0
cc_147 A1 N_VPWR_M1007_d 0.00239384f $X=1.96 $Y=1.105 $X2=0 $Y2=0
cc_148 N_A1_c_167_n N_VPWR_c_305_n 0.0123487f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A1_c_167_n N_VPWR_c_310_n 0.00335922f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A1_c_167_n N_VPWR_c_303_n 0.00406774f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A1_c_167_n N_A_326_297#_c_364_n 0.0122453f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_152 A1 N_A_326_297#_c_364_n 0.0232788f $X=1.96 $Y=1.105 $X2=0 $Y2=0
cc_153 N_A1_c_166_n N_VGND_c_400_n 0.00588898f $X=1.985 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A1_c_166_n N_VGND_c_402_n 0.00412344f $X=1.985 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A2_c_202_n N_A_235_297#_c_231_n 0.00379134f $X=2.49 $Y=1.41 $X2=0 $Y2=0
cc_156 A2 N_A_235_297#_c_231_n 0.00510617f $X=2.51 $Y=1.105 $X2=0 $Y2=0
cc_157 N_A2_c_201_n N_A_235_297#_c_261_n 0.016895f $X=2.465 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A2_c_202_n N_A_235_297#_c_261_n 7.41797e-19 $X=2.49 $Y=1.41 $X2=0 $Y2=0
cc_159 A2 N_A_235_297#_c_261_n 0.0173214f $X=2.51 $Y=1.105 $X2=0 $Y2=0
cc_160 N_A2_c_202_n N_A_235_297#_c_234_n 0.00126328f $X=2.49 $Y=1.41 $X2=0 $Y2=0
cc_161 A2 N_A_235_297#_c_234_n 0.0112959f $X=2.51 $Y=1.105 $X2=0 $Y2=0
cc_162 N_A2_c_201_n N_A_235_297#_c_256_n 0.00181733f $X=2.465 $Y=0.995 $X2=0
+ $Y2=0
cc_163 N_A2_c_202_n N_VPWR_c_305_n 0.00886786f $X=2.49 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A2_c_202_n N_VPWR_c_306_n 0.00717608f $X=2.49 $Y=1.41 $X2=0 $Y2=0
cc_165 A2 N_VPWR_c_306_n 0.00547566f $X=2.51 $Y=1.105 $X2=0 $Y2=0
cc_166 N_A2_c_202_n N_VPWR_c_307_n 0.00482324f $X=2.49 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A2_c_202_n N_VPWR_c_303_n 0.00683347f $X=2.49 $Y=1.41 $X2=0 $Y2=0
cc_168 A2 N_A_326_297#_M1000_d 0.00260575f $X=2.51 $Y=1.105 $X2=0 $Y2=0
cc_169 N_A2_c_202_n N_A_326_297#_c_364_n 0.0140813f $X=2.49 $Y=1.41 $X2=0 $Y2=0
cc_170 A2 N_A_326_297#_c_364_n 0.0103421f $X=2.51 $Y=1.105 $X2=0 $Y2=0
cc_171 A2 N_A_326_297#_c_369_n 0.00572486f $X=2.51 $Y=1.105 $X2=0 $Y2=0
cc_172 N_A2_c_201_n N_VGND_c_400_n 0.00735404f $X=2.465 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A2_c_201_n N_VGND_c_402_n 0.0042361f $X=2.465 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A2_c_201_n N_VGND_c_403_n 0.0144211f $X=2.465 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A_235_297#_c_237_n N_VPWR_c_304_n 0.016227f $X=1.3 $Y=1.63 $X2=0 $Y2=0
cc_176 N_A_235_297#_c_231_n N_VPWR_c_306_n 0.0049899f $X=3.485 $Y=1.41 $X2=0
+ $Y2=0
cc_177 N_A_235_297#_c_234_n N_VPWR_c_306_n 0.00557927f $X=3.45 $Y=1.16 $X2=0
+ $Y2=0
cc_178 N_A_235_297#_c_237_n N_VPWR_c_310_n 0.0198101f $X=1.3 $Y=1.63 $X2=0 $Y2=0
cc_179 N_A_235_297#_c_231_n N_VPWR_c_311_n 0.00702461f $X=3.485 $Y=1.41 $X2=0
+ $Y2=0
cc_180 N_A_235_297#_M1008_s N_VPWR_c_303_n 0.00221957f $X=1.175 $Y=1.485 $X2=0
+ $Y2=0
cc_181 N_A_235_297#_c_231_n N_VPWR_c_303_n 0.0148765f $X=3.485 $Y=1.41 $X2=0
+ $Y2=0
cc_182 N_A_235_297#_c_237_n N_VPWR_c_303_n 0.0124356f $X=1.3 $Y=1.63 $X2=0 $Y2=0
cc_183 N_A_235_297#_c_235_n N_A_326_297#_c_370_n 0.00191131f $X=1.595 $Y=1.195
+ $X2=0 $Y2=0
cc_184 N_A_235_297#_c_231_n X 0.0255501f $X=3.485 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A_235_297#_c_232_n X 0.0291825f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_235_297#_c_261_n X 0.0154713f $X=3.285 $Y=0.72 $X2=0 $Y2=0
cc_187 N_A_235_297#_c_234_n X 0.0389767f $X=3.45 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A_235_297#_c_261_n N_VGND_M1006_d 0.0374112f $X=3.285 $Y=0.72 $X2=0
+ $Y2=0
cc_189 N_A_235_297#_c_234_n N_VGND_M1006_d 0.00277153f $X=3.45 $Y=1.16 $X2=0
+ $Y2=0
cc_190 N_A_235_297#_c_235_n N_VGND_c_397_n 0.0127167f $X=1.595 $Y=1.195 $X2=0
+ $Y2=0
cc_191 N_A_235_297#_c_232_n N_VGND_c_399_n 0.00466641f $X=3.51 $Y=0.995 $X2=0
+ $Y2=0
cc_192 N_A_235_297#_c_261_n N_VGND_c_399_n 0.00314428f $X=3.285 $Y=0.72 $X2=0
+ $Y2=0
cc_193 N_A_235_297#_M1003_d N_VGND_c_400_n 0.00215535f $X=1.64 $Y=0.235 $X2=0
+ $Y2=0
cc_194 N_A_235_297#_c_232_n N_VGND_c_400_n 0.00963052f $X=3.51 $Y=0.995 $X2=0
+ $Y2=0
cc_195 N_A_235_297#_c_261_n N_VGND_c_400_n 0.0268783f $X=3.285 $Y=0.72 $X2=0
+ $Y2=0
cc_196 N_A_235_297#_c_256_n N_VGND_c_400_n 0.0173085f $X=1.775 $Y=0.38 $X2=0
+ $Y2=0
cc_197 N_A_235_297#_c_261_n N_VGND_c_402_n 0.0105706f $X=3.285 $Y=0.72 $X2=0
+ $Y2=0
cc_198 N_A_235_297#_c_256_n N_VGND_c_402_n 0.0263384f $X=1.775 $Y=0.38 $X2=0
+ $Y2=0
cc_199 N_A_235_297#_c_232_n N_VGND_c_403_n 0.0106637f $X=3.51 $Y=0.995 $X2=0
+ $Y2=0
cc_200 N_A_235_297#_c_261_n N_VGND_c_403_n 0.0560776f $X=3.285 $Y=0.72 $X2=0
+ $Y2=0
cc_201 N_A_235_297#_c_261_n A_412_47# 0.00758801f $X=3.285 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_202 N_VPWR_c_303_n N_A_326_297#_M1008_d 0.00449267f $X=3.91 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_203 N_VPWR_c_303_n N_A_326_297#_M1000_d 0.00410926f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_204 N_VPWR_M1007_d N_A_326_297#_c_364_n 0.0058462f $X=2.1 $Y=1.485 $X2=0
+ $Y2=0
cc_205 N_VPWR_c_305_n N_A_326_297#_c_364_n 0.0204605f $X=2.25 $Y=2.24 $X2=0
+ $Y2=0
cc_206 N_VPWR_c_307_n N_A_326_297#_c_364_n 0.00262603f $X=3.075 $Y=2.72 $X2=0
+ $Y2=0
cc_207 N_VPWR_c_310_n N_A_326_297#_c_364_n 0.00192591f $X=2.035 $Y=2.72 $X2=0
+ $Y2=0
cc_208 N_VPWR_c_303_n N_A_326_297#_c_364_n 0.0103798f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_209 N_VPWR_c_310_n N_A_326_297#_c_370_n 0.0116843f $X=2.035 $Y=2.72 $X2=0
+ $Y2=0
cc_210 N_VPWR_c_303_n N_A_326_297#_c_370_n 0.00680917f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_211 N_VPWR_c_305_n N_A_326_297#_c_369_n 0.0180488f $X=2.25 $Y=2.24 $X2=0
+ $Y2=0
cc_212 N_VPWR_c_306_n N_A_326_297#_c_369_n 0.0387968f $X=3.25 $Y=1.66 $X2=0
+ $Y2=0
cc_213 N_VPWR_c_307_n N_A_326_297#_c_369_n 0.0110892f $X=3.075 $Y=2.72 $X2=0
+ $Y2=0
cc_214 N_VPWR_c_303_n N_A_326_297#_c_369_n 0.00643678f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_215 N_VPWR_c_303_n N_X_M1009_d 0.00802392f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_216 N_VPWR_c_311_n X 0.0184162f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_217 N_VPWR_c_303_n X 0.0106557f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_218 X N_VGND_c_399_n 0.0184162f $X=3.78 $Y=0.425 $X2=0 $Y2=0
cc_219 N_X_M1005_d N_VGND_c_400_n 0.00759479f $X=3.585 $Y=0.235 $X2=0 $Y2=0
cc_220 X N_VGND_c_400_n 0.0106557f $X=3.78 $Y=0.425 $X2=0 $Y2=0
cc_221 X N_VGND_c_403_n 0.00903964f $X=3.78 $Y=0.425 $X2=0 $Y2=0
cc_222 N_VGND_c_400_n A_412_47# 0.00380637f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
