* File: sky130_fd_sc_hdll__nand4b_1.pxi.spice
* Created: Thu Aug 27 19:14:40 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND4B_1%A_N N_A_N_c_51_n N_A_N_M1001_g N_A_N_c_52_n
+ N_A_N_M1002_g A_N A_N PM_SKY130_FD_SC_HDLL__NAND4B_1%A_N
x_PM_SKY130_FD_SC_HDLL__NAND4B_1%D N_D_c_78_n N_D_M1008_g N_D_c_79_n N_D_M1009_g
+ D D PM_SKY130_FD_SC_HDLL__NAND4B_1%D
x_PM_SKY130_FD_SC_HDLL__NAND4B_1%C N_C_c_109_n N_C_M1007_g N_C_c_110_n
+ N_C_M1006_g C C PM_SKY130_FD_SC_HDLL__NAND4B_1%C
x_PM_SKY130_FD_SC_HDLL__NAND4B_1%B N_B_c_144_n N_B_M1004_g N_B_c_145_n
+ N_B_M1000_g B B PM_SKY130_FD_SC_HDLL__NAND4B_1%B
x_PM_SKY130_FD_SC_HDLL__NAND4B_1%A_40_93# N_A_40_93#_M1001_s N_A_40_93#_M1002_s
+ N_A_40_93#_c_180_n N_A_40_93#_M1005_g N_A_40_93#_c_181_n N_A_40_93#_M1003_g
+ N_A_40_93#_c_182_n N_A_40_93#_c_193_n N_A_40_93#_c_203_n N_A_40_93#_c_183_n
+ N_A_40_93#_c_184_n N_A_40_93#_c_188_n N_A_40_93#_c_199_n N_A_40_93#_c_185_n
+ PM_SKY130_FD_SC_HDLL__NAND4B_1%A_40_93#
x_PM_SKY130_FD_SC_HDLL__NAND4B_1%VPWR N_VPWR_M1002_d N_VPWR_M1006_d
+ N_VPWR_M1003_d N_VPWR_c_262_n N_VPWR_c_263_n N_VPWR_c_264_n N_VPWR_c_265_n
+ N_VPWR_c_266_n N_VPWR_c_267_n N_VPWR_c_268_n N_VPWR_c_269_n VPWR
+ N_VPWR_c_270_n N_VPWR_c_261_n PM_SKY130_FD_SC_HDLL__NAND4B_1%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND4B_1%Y N_Y_M1005_d N_Y_M1008_d N_Y_M1000_d
+ N_Y_c_310_n N_Y_c_312_n N_Y_c_316_n N_Y_c_318_n N_Y_c_308_n N_Y_c_305_n
+ N_Y_c_323_n N_Y_c_306_n Y N_Y_c_307_n PM_SKY130_FD_SC_HDLL__NAND4B_1%Y
x_PM_SKY130_FD_SC_HDLL__NAND4B_1%VGND N_VGND_M1001_d N_VGND_c_355_n VGND
+ N_VGND_c_356_n N_VGND_c_357_n N_VGND_c_358_n
+ PM_SKY130_FD_SC_HDLL__NAND4B_1%VGND
cc_1 VNB N_A_N_c_51_n 0.0219089f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=0.995
cc_2 VNB N_A_N_c_52_n 0.0285844f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.41
cc_3 VNB A_N 0.00282596f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_4 VNB N_D_c_78_n 0.0264207f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=0.995
cc_5 VNB N_D_c_79_n 0.0197201f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.41
cc_6 VNB D 0.00207248f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_7 VNB N_C_c_109_n 0.0161784f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=0.995
cc_8 VNB N_C_c_110_n 0.0206045f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.41
cc_9 VNB C 0.00319507f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_10 VNB N_B_c_144_n 0.0163265f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=0.995
cc_11 VNB N_B_c_145_n 0.0206111f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.41
cc_12 VNB B 0.00323605f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_13 VNB N_A_40_93#_c_180_n 0.0195248f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_14 VNB N_A_40_93#_c_181_n 0.0254907f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_15 VNB N_A_40_93#_c_182_n 0.0224554f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=1.16
cc_16 VNB N_A_40_93#_c_183_n 9.39379e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_40_93#_c_184_n 0.0208983f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_40_93#_c_185_n 0.00208581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_261_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_305_n 0.0235709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_306_n 0.00710642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_Y_c_307_n 0.0161093f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_355_n 0.0113245f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_356_n 0.0583061f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_357_n 0.185936f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_358_n 0.0269741f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VPB N_A_N_c_52_n 0.035521f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.41
cc_28 VPB A_N 0.00205184f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_29 VPB N_D_c_78_n 0.0323882f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=0.995
cc_30 VPB D 3.01511e-19 $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_31 VPB N_C_c_110_n 0.0251745f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.41
cc_32 VPB C 6.65656e-19 $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_33 VPB N_B_c_145_n 0.0251353f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.41
cc_34 VPB B 8.1666e-19 $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_35 VPB N_A_40_93#_c_181_n 0.0283409f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_36 VPB N_A_40_93#_c_182_n 0.0149907f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=1.16
cc_37 VPB N_A_40_93#_c_188_n 0.0232716f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_40_93#_c_185_n 9.473e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_262_n 0.0232531f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_40 VPB N_VPWR_c_263_n 0.00524573f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_264_n 0.0104574f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_265_n 0.0279645f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_266_n 0.0261689f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_267_n 0.00477947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_268_n 0.0190531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_269_n 0.00525886f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_270_n 0.0244675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_261_n 0.05603f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_Y_c_308_n 0.00907079f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_Y_c_305_n 0.010274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 N_A_N_c_52_n N_D_c_78_n 0.034704f $X=0.62 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_52 A_N N_D_c_78_n 0.00226422f $X=0.605 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_53 N_A_N_c_51_n N_D_c_79_n 0.0164844f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_54 N_A_N_c_52_n D 2.99721e-19 $X=0.62 $Y=1.41 $X2=0 $Y2=0
cc_55 A_N D 0.0243847f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_56 N_A_N_c_51_n N_A_40_93#_c_182_n 0.00526949f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_57 N_A_N_c_52_n N_A_40_93#_c_182_n 0.0153742f $X=0.62 $Y=1.41 $X2=0 $Y2=0
cc_58 A_N N_A_40_93#_c_182_n 0.0251136f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_59 N_A_N_c_51_n N_A_40_93#_c_193_n 0.0106906f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_60 N_A_N_c_51_n N_A_40_93#_c_184_n 4.38141e-19 $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_61 N_A_N_c_52_n N_A_40_93#_c_184_n 0.00540014f $X=0.62 $Y=1.41 $X2=0 $Y2=0
cc_62 A_N N_A_40_93#_c_184_n 0.0252267f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_63 N_A_N_c_52_n N_A_40_93#_c_188_n 0.00518047f $X=0.62 $Y=1.41 $X2=0 $Y2=0
cc_64 A_N N_A_40_93#_c_188_n 0.00344351f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_65 N_A_N_c_51_n N_A_40_93#_c_199_n 9.1283e-19 $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_66 N_A_N_c_52_n N_VPWR_c_262_n 0.00545995f $X=0.62 $Y=1.41 $X2=0 $Y2=0
cc_67 A_N N_VPWR_c_262_n 0.00505451f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_68 N_A_N_c_52_n N_VPWR_c_266_n 0.00393512f $X=0.62 $Y=1.41 $X2=0 $Y2=0
cc_69 N_A_N_c_52_n N_VPWR_c_261_n 0.00500987f $X=0.62 $Y=1.41 $X2=0 $Y2=0
cc_70 N_A_N_c_51_n N_VGND_c_355_n 0.00387685f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_71 N_A_N_c_51_n N_VGND_c_357_n 0.00512902f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_72 N_A_N_c_51_n N_VGND_c_358_n 0.00392914f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_73 N_D_c_79_n N_C_c_109_n 0.0424006f $X=1.18 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_74 N_D_c_78_n N_C_c_110_n 0.0361505f $X=1.155 $Y=1.41 $X2=0 $Y2=0
cc_75 D N_C_c_110_n 0.00101956f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_76 N_D_c_78_n C 9.80911e-19 $X=1.155 $Y=1.41 $X2=0 $Y2=0
cc_77 N_D_c_79_n C 0.00160005f $X=1.18 $Y=0.995 $X2=0 $Y2=0
cc_78 D C 0.0270082f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_79 N_D_c_78_n N_A_40_93#_c_193_n 0.00442168f $X=1.155 $Y=1.41 $X2=0 $Y2=0
cc_80 N_D_c_79_n N_A_40_93#_c_193_n 0.00826642f $X=1.18 $Y=0.995 $X2=0 $Y2=0
cc_81 D N_A_40_93#_c_193_n 0.0117288f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_82 N_D_c_79_n N_A_40_93#_c_203_n 2.09696e-19 $X=1.18 $Y=0.995 $X2=0 $Y2=0
cc_83 N_D_c_79_n N_A_40_93#_c_199_n 0.00987447f $X=1.18 $Y=0.995 $X2=0 $Y2=0
cc_84 D N_A_40_93#_c_199_n 0.00779052f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_85 N_D_c_78_n N_VPWR_c_262_n 0.00998255f $X=1.155 $Y=1.41 $X2=0 $Y2=0
cc_86 N_D_c_78_n N_VPWR_c_268_n 0.00597712f $X=1.155 $Y=1.41 $X2=0 $Y2=0
cc_87 N_D_c_78_n N_VPWR_c_261_n 0.0113021f $X=1.155 $Y=1.41 $X2=0 $Y2=0
cc_88 N_D_c_78_n N_Y_c_310_n 0.00452336f $X=1.155 $Y=1.41 $X2=0 $Y2=0
cc_89 D N_Y_c_310_n 0.010089f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_90 N_D_c_78_n N_Y_c_312_n 0.0120097f $X=1.155 $Y=1.41 $X2=0 $Y2=0
cc_91 N_D_c_79_n N_VGND_c_355_n 0.0116446f $X=1.18 $Y=0.995 $X2=0 $Y2=0
cc_92 N_D_c_79_n N_VGND_c_356_n 0.00415631f $X=1.18 $Y=0.995 $X2=0 $Y2=0
cc_93 N_D_c_79_n N_VGND_c_357_n 0.00706529f $X=1.18 $Y=0.995 $X2=0 $Y2=0
cc_94 N_C_c_109_n N_B_c_144_n 0.034466f $X=1.595 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_95 C N_B_c_144_n 6.57426e-19 $X=1.525 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_96 N_C_c_110_n N_B_c_145_n 0.0468539f $X=1.625 $Y=1.41 $X2=0 $Y2=0
cc_97 C N_B_c_145_n 3.39346e-19 $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_98 N_C_c_109_n B 6.62669e-19 $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_99 N_C_c_110_n B 0.00191591f $X=1.625 $Y=1.41 $X2=0 $Y2=0
cc_100 C B 0.0438224f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_101 N_C_c_109_n N_A_40_93#_c_203_n 0.0103767f $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_102 N_C_c_110_n N_A_40_93#_c_203_n 0.00117431f $X=1.625 $Y=1.41 $X2=0 $Y2=0
cc_103 C N_A_40_93#_c_203_n 0.0132366f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_104 N_C_c_109_n N_A_40_93#_c_199_n 0.00410404f $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_105 C N_A_40_93#_c_199_n 0.00431714f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_106 N_C_c_110_n N_VPWR_c_263_n 0.00311303f $X=1.625 $Y=1.41 $X2=0 $Y2=0
cc_107 N_C_c_110_n N_VPWR_c_268_n 0.00673617f $X=1.625 $Y=1.41 $X2=0 $Y2=0
cc_108 N_C_c_110_n N_VPWR_c_261_n 0.0117925f $X=1.625 $Y=1.41 $X2=0 $Y2=0
cc_109 N_C_c_110_n N_Y_c_310_n 5.7874e-19 $X=1.625 $Y=1.41 $X2=0 $Y2=0
cc_110 C N_Y_c_310_n 0.00304392f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_111 N_C_c_110_n N_Y_c_312_n 0.0100689f $X=1.625 $Y=1.41 $X2=0 $Y2=0
cc_112 N_C_c_110_n N_Y_c_316_n 0.0147181f $X=1.625 $Y=1.41 $X2=0 $Y2=0
cc_113 C N_Y_c_316_n 0.0137982f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_114 N_C_c_110_n N_Y_c_318_n 5.94842e-19 $X=1.625 $Y=1.41 $X2=0 $Y2=0
cc_115 N_C_c_109_n N_VGND_c_356_n 0.00390868f $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_116 N_C_c_109_n N_VGND_c_357_n 0.00563134f $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_117 C A_334_47# 0.00138412f $X=1.525 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_118 N_B_c_144_n N_A_40_93#_c_180_n 0.0331984f $X=2.08 $Y=0.995 $X2=0 $Y2=0
cc_119 B N_A_40_93#_c_180_n 6.62814e-19 $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_120 N_B_c_145_n N_A_40_93#_c_181_n 0.0339219f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_121 B N_A_40_93#_c_181_n 3.16969e-19 $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_122 N_B_c_144_n N_A_40_93#_c_203_n 0.0112915f $X=2.08 $Y=0.995 $X2=0 $Y2=0
cc_123 N_B_c_145_n N_A_40_93#_c_203_n 0.00168052f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_124 B N_A_40_93#_c_203_n 0.0131757f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_125 N_B_c_144_n N_A_40_93#_c_183_n 0.00407484f $X=2.08 $Y=0.995 $X2=0 $Y2=0
cc_126 B N_A_40_93#_c_183_n 0.0179859f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_127 N_B_c_145_n N_A_40_93#_c_185_n 0.00197607f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_128 B N_A_40_93#_c_185_n 0.0258731f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_129 N_B_c_145_n N_VPWR_c_263_n 0.00308286f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_130 N_B_c_145_n N_VPWR_c_270_n 0.00673617f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_131 N_B_c_145_n N_VPWR_c_261_n 0.0118287f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_132 N_B_c_145_n N_Y_c_312_n 5.89583e-19 $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_133 N_B_c_145_n N_Y_c_316_n 0.0138057f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_134 B N_Y_c_316_n 0.0167037f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_135 N_B_c_145_n N_Y_c_318_n 0.0101423f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_136 N_B_c_145_n N_Y_c_323_n 0.00255341f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_137 B N_Y_c_323_n 0.00284414f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_138 N_B_c_144_n N_VGND_c_356_n 0.00390868f $X=2.08 $Y=0.995 $X2=0 $Y2=0
cc_139 N_B_c_144_n N_VGND_c_357_n 0.00579024f $X=2.08 $Y=0.995 $X2=0 $Y2=0
cc_140 B A_334_47# 0.00123785f $X=1.985 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_141 B A_431_47# 0.001186f $X=1.985 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_142 N_A_40_93#_c_193_n N_VPWR_c_262_n 0.00529132f $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A_40_93#_c_188_n N_VPWR_c_262_n 0.00114497f $X=0.385 $Y=1.76 $X2=0
+ $Y2=0
cc_144 N_A_40_93#_c_181_n N_VPWR_c_265_n 0.0175891f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_40_93#_c_181_n N_VPWR_c_270_n 0.00688798f $X=2.585 $Y=1.41 $X2=0
+ $Y2=0
cc_146 N_A_40_93#_c_181_n N_VPWR_c_261_n 0.0134952f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_40_93#_c_188_n N_VPWR_c_261_n 0.0159191f $X=0.385 $Y=1.76 $X2=0 $Y2=0
cc_148 N_A_40_93#_c_199_n N_Y_c_310_n 0.00119657f $X=1.285 $Y=0.51 $X2=0 $Y2=0
cc_149 N_A_40_93#_c_181_n N_Y_c_318_n 0.0169775f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_40_93#_c_181_n N_Y_c_308_n 0.0179968f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_40_93#_c_185_n N_Y_c_308_n 0.0132319f $X=2.62 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_40_93#_c_180_n N_Y_c_305_n 0.00301227f $X=2.56 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_40_93#_c_181_n N_Y_c_305_n 0.0137127f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_40_93#_c_183_n N_Y_c_305_n 0.00826683f $X=2.497 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_40_93#_c_185_n N_Y_c_305_n 0.0254799f $X=2.62 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_40_93#_c_181_n N_Y_c_323_n 2.74535e-19 $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_40_93#_c_185_n N_Y_c_323_n 0.00682585f $X=2.62 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A_40_93#_c_180_n N_Y_c_307_n 0.0149034f $X=2.56 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A_40_93#_c_203_n N_Y_c_307_n 0.0137835f $X=2.395 $Y=0.51 $X2=0 $Y2=0
cc_160 N_A_40_93#_c_183_n N_Y_c_307_n 0.0176473f $X=2.497 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_40_93#_c_193_n N_VGND_M1001_d 0.00902465f $X=1.2 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_162 N_A_40_93#_c_193_n N_VGND_c_355_n 0.0235676f $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A_40_93#_c_184_n N_VGND_c_355_n 0.00139179f $X=0.47 $Y=0.635 $X2=0
+ $Y2=0
cc_164 N_A_40_93#_c_199_n N_VGND_c_355_n 0.004476f $X=1.285 $Y=0.51 $X2=0 $Y2=0
cc_165 N_A_40_93#_c_180_n N_VGND_c_356_n 0.00436118f $X=2.56 $Y=0.995 $X2=0
+ $Y2=0
cc_166 N_A_40_93#_c_193_n N_VGND_c_356_n 0.00230621f $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A_40_93#_c_203_n N_VGND_c_356_n 0.0333809f $X=2.395 $Y=0.51 $X2=0 $Y2=0
cc_168 N_A_40_93#_c_199_n N_VGND_c_356_n 0.00448622f $X=1.285 $Y=0.51 $X2=0
+ $Y2=0
cc_169 N_A_40_93#_c_180_n N_VGND_c_357_n 0.00799415f $X=2.56 $Y=0.995 $X2=0
+ $Y2=0
cc_170 N_A_40_93#_c_193_n N_VGND_c_357_n 0.011166f $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A_40_93#_c_203_n N_VGND_c_357_n 0.0391223f $X=2.395 $Y=0.51 $X2=0 $Y2=0
cc_172 N_A_40_93#_c_184_n N_VGND_c_357_n 0.0129566f $X=0.47 $Y=0.635 $X2=0 $Y2=0
cc_173 N_A_40_93#_c_199_n N_VGND_c_357_n 0.00548271f $X=1.285 $Y=0.51 $X2=0
+ $Y2=0
cc_174 N_A_40_93#_c_193_n N_VGND_c_358_n 0.00274635f $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A_40_93#_c_184_n N_VGND_c_358_n 0.0118851f $X=0.47 $Y=0.635 $X2=0 $Y2=0
cc_176 N_A_40_93#_c_203_n A_251_47# 0.00515702f $X=2.395 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_177 N_A_40_93#_c_199_n A_251_47# 0.00465616f $X=1.285 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_178 N_A_40_93#_c_203_n A_334_47# 0.00912908f $X=2.395 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_179 N_A_40_93#_c_203_n A_431_47# 0.00816035f $X=2.395 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_180 N_A_40_93#_c_183_n A_431_47# 0.00313788f $X=2.497 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_181 N_VPWR_c_261_n N_Y_M1008_d 0.00231261f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_182 N_VPWR_c_261_n N_Y_M1000_d 0.00239291f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_183 N_VPWR_c_262_n N_Y_c_310_n 0.0137304f $X=0.92 $Y=1.66 $X2=0 $Y2=0
cc_184 N_VPWR_c_262_n N_Y_c_312_n 0.0614133f $X=0.92 $Y=1.66 $X2=0 $Y2=0
cc_185 N_VPWR_c_268_n N_Y_c_312_n 0.0223557f $X=1.725 $Y=2.72 $X2=0 $Y2=0
cc_186 N_VPWR_c_261_n N_Y_c_312_n 0.0140101f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_187 N_VPWR_M1006_d N_Y_c_316_n 0.00782613f $X=1.715 $Y=1.485 $X2=0 $Y2=0
cc_188 N_VPWR_c_263_n N_Y_c_316_n 0.0151327f $X=1.86 $Y=2 $X2=0 $Y2=0
cc_189 N_VPWR_c_265_n N_Y_c_318_n 0.0260218f $X=2.96 $Y=2 $X2=0 $Y2=0
cc_190 N_VPWR_c_270_n N_Y_c_318_n 0.0189681f $X=2.875 $Y=2.72 $X2=0 $Y2=0
cc_191 N_VPWR_c_261_n N_Y_c_318_n 0.0123589f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_192 N_VPWR_M1003_d N_Y_c_308_n 0.0128821f $X=2.675 $Y=1.485 $X2=0 $Y2=0
cc_193 N_VPWR_c_265_n N_Y_c_308_n 0.0192186f $X=2.96 $Y=2 $X2=0 $Y2=0
cc_194 N_VPWR_M1003_d N_Y_c_305_n 2.11855e-19 $X=2.675 $Y=1.485 $X2=0 $Y2=0
cc_195 N_Y_c_307_n N_VGND_c_356_n 0.0251617f $X=2.94 $Y=0.405 $X2=0 $Y2=0
cc_196 N_Y_M1005_d N_VGND_c_357_n 0.00855375f $X=2.635 $Y=0.235 $X2=0 $Y2=0
cc_197 N_Y_c_307_n N_VGND_c_357_n 0.0137714f $X=2.94 $Y=0.405 $X2=0 $Y2=0
cc_198 N_VGND_c_357_n A_251_47# 0.00237957f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_199 N_VGND_c_357_n A_334_47# 0.00302096f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_200 N_VGND_c_357_n A_431_47# 0.00297499f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
