* File: sky130_fd_sc_hdll__a21bo_4.spice
* Created: Thu Aug 27 18:52:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a21bo_4.pex.spice"
.subckt sky130_fd_sc_hdll__a21bo_4  VNB VPB B1_N A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_B1_N_M1013_g N_A_36_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.28275 PD=0.93 PS=2.17 NRD=0 NRS=23.988 M=1 R=4.33333 SA=75000.4
+ SB=75005.5 A=0.0975 P=1.6 MULT=1
MM1001 N_X_M1001_d N_A_209_21#_M1001_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.091 PD=0.98 PS=0.93 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.8
+ SB=75005 A=0.0975 P=1.6 MULT=1
MM1004 N_X_M1001_d N_A_209_21#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75001.3
+ SB=75004.6 A=0.0975 P=1.6 MULT=1
MM1007 N_X_M1007_d N_A_209_21#_M1007_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1007_d N_A_209_21#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.29575 PD=0.98 PS=1.56 NRD=0 NRS=29.532 M=1 R=4.33333
+ SA=75002.2 SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1009_s N_A_36_47#_M1010_g N_A_209_21#_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.29575 AS=0.104 PD=1.56 PS=0.97 NRD=11.988 NRS=0 M=1 R=4.33333
+ SA=75003.3 SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1016_d N_A_36_47#_M1016_g N_A_209_21#_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.117 AS=0.104 PD=1.01 PS=0.97 NRD=6.456 NRS=8.304 M=1 R=4.33333
+ SA=75003.8 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1015 A_1115_47# N_A2_M1015_g N_VGND_M1016_d VNB NSHORT L=0.15 W=0.65
+ AD=0.07475 AS=0.117 PD=0.88 PS=1.01 NRD=11.076 NRS=8.304 M=1 R=4.33333
+ SA=75004.3 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1011 N_A_209_21#_M1011_d N_A1_M1011_g A_1115_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.07475 PD=1.02 PS=0.88 NRD=8.304 NRS=11.076 M=1 R=4.33333
+ SA=75004.6 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1021 N_A_209_21#_M1011_d N_A1_M1021_g A_935_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=14.76 M=1 R=4.33333
+ SA=75005.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1017 A_935_47# N_A2_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.2015 PD=0.92 PS=1.92 NRD=14.76 NRS=8.304 M=1 R=4.33333 SA=75005.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_B1_N_M1003_g N_A_36_47#_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90002.1 A=0.18 P=2.36 MULT=1
MM1000 N_X_M1000_d N_A_209_21#_M1000_g N_VPWR_M1003_d VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1006 N_X_M1000_d N_A_209_21#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.1
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1012 N_X_M1012_d N_A_209_21#_M1012_g N_VPWR_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.6
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1018 N_X_M1012_d N_A_209_21#_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.29 PD=1.3 PS=2.58 NRD=1.9503 NRS=0.9653 M=1 R=5.55556 SA=90002.1
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1005 N_A_647_297#_M1005_d N_A_36_47#_M1005_g N_A_209_21#_M1005_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.2 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1019 N_A_647_297#_M1019_d N_A_36_47#_M1019_g N_A_209_21#_M1005_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A2_M1002_g N_A_647_297#_M1019_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1014 N_VPWR_M1002_d N_A1_M1014_g N_A_647_297#_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1020 N_VPWR_M1020_d N_A1_M1020_g N_A_647_297#_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1020_d N_A2_M1008_g N_A_647_297#_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90000.2 A=0.18 P=2.36 MULT=1
DX22_noxref VNB VPB NWDIODE A=10.9461 P=16.85
pX23_noxref noxref_14 A2 A2 PROBETYPE=1
c_42 VNB 0 1.1034e-19 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hdll__a21bo_4.pxi.spice"
*
.ends
*
*
