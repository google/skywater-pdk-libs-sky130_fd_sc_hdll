* File: sky130_fd_sc_hdll__nor2_8.pxi.spice
* Created: Thu Aug 27 19:15:43 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR2_8%A N_A_c_113_n N_A_M1004_g N_A_c_123_n N_A_M1001_g
+ N_A_c_114_n N_A_M1010_g N_A_c_124_n N_A_M1002_g N_A_c_115_n N_A_M1012_g
+ N_A_c_125_n N_A_M1008_g N_A_c_116_n N_A_M1016_g N_A_c_126_n N_A_M1013_g
+ N_A_c_117_n N_A_M1022_g N_A_c_127_n N_A_M1018_g N_A_c_118_n N_A_M1025_g
+ N_A_c_128_n N_A_M1021_g N_A_c_119_n N_A_M1027_g N_A_c_129_n N_A_M1026_g
+ N_A_c_130_n N_A_M1030_g N_A_c_120_n N_A_M1028_g A N_A_c_121_n N_A_c_122_n A
+ PM_SKY130_FD_SC_HDLL__NOR2_8%A
x_PM_SKY130_FD_SC_HDLL__NOR2_8%B N_B_c_253_n N_B_M1000_g N_B_c_262_n N_B_M1003_g
+ N_B_c_254_n N_B_M1005_g N_B_c_263_n N_B_M1006_g N_B_c_255_n N_B_M1007_g
+ N_B_c_264_n N_B_M1009_g N_B_c_256_n N_B_M1014_g N_B_c_265_n N_B_M1011_g
+ N_B_c_257_n N_B_M1017_g N_B_c_266_n N_B_M1015_g N_B_c_258_n N_B_M1020_g
+ N_B_c_267_n N_B_M1019_g N_B_c_259_n N_B_M1023_g N_B_c_268_n N_B_M1024_g
+ N_B_c_269_n N_B_M1029_g N_B_c_260_n N_B_M1031_g B N_B_c_273_n N_B_c_261_n B
+ PM_SKY130_FD_SC_HDLL__NOR2_8%B
x_PM_SKY130_FD_SC_HDLL__NOR2_8%A_27_297# N_A_27_297#_M1001_s N_A_27_297#_M1002_s
+ N_A_27_297#_M1013_s N_A_27_297#_M1021_s N_A_27_297#_M1030_s
+ N_A_27_297#_M1006_s N_A_27_297#_M1011_s N_A_27_297#_M1019_s
+ N_A_27_297#_M1029_s N_A_27_297#_c_392_n N_A_27_297#_c_393_n
+ N_A_27_297#_c_394_n N_A_27_297#_c_440_p N_A_27_297#_c_395_n
+ N_A_27_297#_c_442_p N_A_27_297#_c_396_n N_A_27_297#_c_444_p
+ N_A_27_297#_c_397_n N_A_27_297#_c_398_n N_A_27_297#_c_446_p
+ N_A_27_297#_c_427_n N_A_27_297#_c_483_p N_A_27_297#_c_429_n
+ N_A_27_297#_c_487_p N_A_27_297#_c_431_n N_A_27_297#_c_490_p
+ N_A_27_297#_c_433_n N_A_27_297#_c_493_p N_A_27_297#_c_399_n
+ N_A_27_297#_c_400_n N_A_27_297#_c_401_n N_A_27_297#_c_451_p
+ N_A_27_297#_c_452_p N_A_27_297#_c_453_p PM_SKY130_FD_SC_HDLL__NOR2_8%A_27_297#
x_PM_SKY130_FD_SC_HDLL__NOR2_8%VPWR N_VPWR_M1001_d N_VPWR_M1008_d N_VPWR_M1018_d
+ N_VPWR_M1026_d N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n
+ N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_502_n VPWR N_VPWR_c_503_n
+ N_VPWR_c_495_n N_VPWR_c_505_n N_VPWR_c_506_n N_VPWR_c_507_n N_VPWR_c_508_n
+ PM_SKY130_FD_SC_HDLL__NOR2_8%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR2_8%Y N_Y_M1004_s N_Y_M1012_s N_Y_M1022_s N_Y_M1027_s
+ N_Y_M1000_d N_Y_M1007_d N_Y_M1017_d N_Y_M1023_d N_Y_M1003_d N_Y_M1009_d
+ N_Y_M1015_d N_Y_M1024_d N_Y_c_617_n N_Y_c_594_n N_Y_c_595_n N_Y_c_628_n
+ N_Y_c_596_n N_Y_c_636_n N_Y_c_597_n N_Y_c_644_n N_Y_c_598_n N_Y_c_648_n
+ N_Y_c_731_n N_Y_c_610_n N_Y_c_611_n N_Y_c_599_n N_Y_c_676_n N_Y_c_735_n
+ N_Y_c_612_n N_Y_c_600_n N_Y_c_688_n N_Y_c_738_n N_Y_c_613_n N_Y_c_601_n
+ N_Y_c_741_n N_Y_c_602_n N_Y_c_603_n N_Y_c_604_n N_Y_c_605_n N_Y_c_606_n
+ N_Y_c_614_n N_Y_c_607_n N_Y_c_615_n N_Y_c_608_n Y
+ PM_SKY130_FD_SC_HDLL__NOR2_8%Y
x_PM_SKY130_FD_SC_HDLL__NOR2_8%VGND N_VGND_M1004_d N_VGND_M1010_d N_VGND_M1016_d
+ N_VGND_M1025_d N_VGND_M1028_d N_VGND_M1005_s N_VGND_M1014_s N_VGND_M1020_s
+ N_VGND_M1031_s N_VGND_c_817_n N_VGND_c_818_n N_VGND_c_819_n N_VGND_c_820_n
+ N_VGND_c_821_n N_VGND_c_822_n N_VGND_c_823_n N_VGND_c_824_n N_VGND_c_825_n
+ N_VGND_c_826_n N_VGND_c_827_n N_VGND_c_828_n N_VGND_c_829_n N_VGND_c_830_n
+ N_VGND_c_831_n N_VGND_c_832_n N_VGND_c_833_n N_VGND_c_834_n N_VGND_c_835_n
+ N_VGND_c_836_n N_VGND_c_837_n N_VGND_c_838_n N_VGND_c_839_n N_VGND_c_840_n
+ N_VGND_c_841_n N_VGND_c_842_n VGND N_VGND_c_843_n N_VGND_c_844_n
+ PM_SKY130_FD_SC_HDLL__NOR2_8%VGND
cc_1 VNB N_A_c_113_n 0.0218461f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_114_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_3 VNB N_A_c_115_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_4 VNB N_A_c_116_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=0.995
cc_5 VNB N_A_c_117_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=2.37 $Y2=0.995
cc_6 VNB N_A_c_118_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=2.84 $Y2=0.995
cc_7 VNB N_A_c_119_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=3.31 $Y2=0.995
cc_8 VNB N_A_c_120_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=3.83 $Y2=0.995
cc_9 VNB N_A_c_121_n 0.0124434f $X=-0.19 $Y=-0.24 $X2=3.67 $Y2=1.16
cc_10 VNB N_A_c_122_n 0.155395f $X=-0.19 $Y=-0.24 $X2=3.805 $Y2=1.202
cc_11 VNB N_B_c_253_n 0.0164943f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_12 VNB N_B_c_254_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_13 VNB N_B_c_255_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_14 VNB N_B_c_256_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=0.995
cc_15 VNB N_B_c_257_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=2.37 $Y2=0.995
cc_16 VNB N_B_c_258_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=2.84 $Y2=0.995
cc_17 VNB N_B_c_259_n 0.0171931f $X=-0.19 $Y=-0.24 $X2=3.31 $Y2=0.995
cc_18 VNB N_B_c_260_n 0.0203186f $X=-0.19 $Y=-0.24 $X2=3.83 $Y2=0.995
cc_19 VNB N_B_c_261_n 0.153702f $X=-0.19 $Y=-0.24 $X2=3.805 $Y2=1.202
cc_20 VNB N_VPWR_c_495_n 0.345644f $X=-0.19 $Y=-0.24 $X2=3.805 $Y2=1.985
cc_21 VNB N_Y_c_594_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=3.335 $Y2=1.985
cc_22 VNB N_Y_c_595_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=3.335 $Y2=1.985
cc_23 VNB N_Y_c_596_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=3.83 $Y2=0.56
cc_24 VNB N_Y_c_597_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.202
cc_25 VNB N_Y_c_598_n 0.0043236f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.202
cc_26 VNB N_Y_c_599_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=3.805 $Y2=1.202
cc_27 VNB N_Y_c_600_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_Y_c_601_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_Y_c_602_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_Y_c_603_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_Y_c_604_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_605_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_Y_c_606_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_Y_c_607_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_Y_c_608_n 0.0117165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB Y 0.0190689f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_817_n 0.0103581f $X=-0.19 $Y=-0.24 $X2=2.395 $Y2=1.41
cc_38 VNB N_VGND_c_818_n 0.0351736f $X=-0.19 $Y=-0.24 $X2=2.395 $Y2=1.985
cc_39 VNB N_VGND_c_819_n 0.0198149f $X=-0.19 $Y=-0.24 $X2=2.84 $Y2=0.56
cc_40 VNB N_VGND_c_820_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=2.865 $Y2=1.985
cc_41 VNB N_VGND_c_821_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=3.335 $Y2=1.41
cc_42 VNB N_VGND_c_822_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=3.805 $Y2=1.985
cc_43 VNB N_VGND_c_823_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=3.83 $Y2=0.56
cc_44 VNB N_VGND_c_824_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_45 VNB N_VGND_c_825_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=1.202
cc_46 VNB N_VGND_c_826_n 0.00467908f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=1.202
cc_47 VNB N_VGND_c_827_n 0.0187002f $X=-0.19 $Y=-0.24 $X2=2.84 $Y2=1.202
cc_48 VNB N_VGND_c_828_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=3.335 $Y2=1.202
cc_49 VNB N_VGND_c_829_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=3.67 $Y2=1.202
cc_50 VNB N_VGND_c_830_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=3.67 $Y2=1.16
cc_51 VNB N_VGND_c_831_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=3.805 $Y2=1.202
cc_52 VNB N_VGND_c_832_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.175
cc_53 VNB N_VGND_c_833_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_834_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.19
cc_55 VNB N_VGND_c_835_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0.74 $Y2=1.175
cc_56 VNB N_VGND_c_836_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_837_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_838_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_839_n 0.00323927f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_840_n 0.0108236f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_841_n 0.0192963f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_842_n 0.00555039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_843_n 0.396068f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_844_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VPB N_A_c_123_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_66 VPB N_A_c_124_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_67 VPB N_A_c_125_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_68 VPB N_A_c_126_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_69 VPB N_A_c_127_n 0.0159747f $X=-0.19 $Y=1.305 $X2=2.395 $Y2=1.41
cc_70 VPB N_A_c_128_n 0.0159747f $X=-0.19 $Y=1.305 $X2=2.865 $Y2=1.41
cc_71 VPB N_A_c_129_n 0.0159747f $X=-0.19 $Y=1.305 $X2=3.335 $Y2=1.41
cc_72 VPB N_A_c_130_n 0.0161059f $X=-0.19 $Y=1.305 $X2=3.805 $Y2=1.41
cc_73 VPB N_A_c_122_n 0.0997653f $X=-0.19 $Y=1.305 $X2=3.805 $Y2=1.202
cc_74 VPB N_B_c_262_n 0.0164196f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_75 VPB N_B_c_263_n 0.0158911f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_76 VPB N_B_c_264_n 0.0158911f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_77 VPB N_B_c_265_n 0.0158911f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_78 VPB N_B_c_266_n 0.0158911f $X=-0.19 $Y=1.305 $X2=2.395 $Y2=1.41
cc_79 VPB N_B_c_267_n 0.0158911f $X=-0.19 $Y=1.305 $X2=2.865 $Y2=1.41
cc_80 VPB N_B_c_268_n 0.0158911f $X=-0.19 $Y=1.305 $X2=3.335 $Y2=1.41
cc_81 VPB N_B_c_269_n 0.0192434f $X=-0.19 $Y=1.305 $X2=3.805 $Y2=1.41
cc_82 VPB N_B_c_261_n 0.0978077f $X=-0.19 $Y=1.305 $X2=3.805 $Y2=1.202
cc_83 VPB N_A_27_297#_c_392_n 0.013626f $X=-0.19 $Y=1.305 $X2=2.395 $Y2=1.41
cc_84 VPB N_A_27_297#_c_393_n 0.0312291f $X=-0.19 $Y=1.305 $X2=2.395 $Y2=1.985
cc_85 VPB N_A_27_297#_c_394_n 0.00200404f $X=-0.19 $Y=1.305 $X2=2.84 $Y2=0.56
cc_86 VPB N_A_27_297#_c_395_n 0.00197374f $X=-0.19 $Y=1.305 $X2=3.31 $Y2=0.56
cc_87 VPB N_A_27_297#_c_396_n 0.00197374f $X=-0.19 $Y=1.305 $X2=3.805 $Y2=1.985
cc_88 VPB N_A_27_297#_c_397_n 0.00200404f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_27_297#_c_398_n 0.00410774f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_90 VPB N_A_27_297#_c_399_n 0.0015364f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_27_297#_c_400_n 0.0015364f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_27_297#_c_401_n 0.0015364f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_496_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.985
cc_94 VPB N_VPWR_c_497_n 0.0195604f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=0.995
cc_95 VPB N_VPWR_c_498_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.985
cc_96 VPB N_VPWR_c_499_n 0.0195604f $X=-0.19 $Y=1.305 $X2=2.37 $Y2=0.995
cc_97 VPB N_VPWR_c_500_n 0.00516582f $X=-0.19 $Y=1.305 $X2=2.395 $Y2=1.985
cc_98 VPB N_VPWR_c_501_n 0.0195604f $X=-0.19 $Y=1.305 $X2=2.84 $Y2=0.995
cc_99 VPB N_VPWR_c_502_n 0.00516582f $X=-0.19 $Y=1.305 $X2=2.865 $Y2=1.985
cc_100 VPB N_VPWR_c_503_n 0.10924f $X=-0.19 $Y=1.305 $X2=3.805 $Y2=1.985
cc_101 VPB N_VPWR_c_495_n 0.0548233f $X=-0.19 $Y=1.305 $X2=3.805 $Y2=1.985
cc_102 VPB N_VPWR_c_505_n 0.0238702f $X=-0.19 $Y=1.305 $X2=3.83 $Y2=0.56
cc_103 VPB N_VPWR_c_506_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.202
cc_104 VPB N_VPWR_c_507_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_105 VPB N_VPWR_c_508_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_106 VPB N_Y_c_610_n 0.00192677f $X=-0.19 $Y=1.305 $X2=3.67 $Y2=1.16
cc_107 VPB N_Y_c_611_n 0.00188018f $X=-0.19 $Y=1.305 $X2=3.67 $Y2=1.16
cc_108 VPB N_Y_c_612_n 0.00192677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_Y_c_613_n 0.00192677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_Y_c_614_n 0.0014926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_Y_c_615_n 0.0014926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB Y 0.0204115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 N_A_c_120_n N_B_c_253_n 0.0245267f $X=3.83 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_114 N_A_c_130_n N_B_c_262_n 0.00966468f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A_c_121_n N_B_c_273_n 0.0124677f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_c_122_n N_B_c_273_n 2.30564e-19 $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_117 N_A_c_121_n N_B_c_261_n 0.00158796f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_c_122_n N_B_c_261_n 0.0245267f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_119 N_A_c_121_n N_A_27_297#_c_392_n 0.0036906f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A_c_123_n N_A_27_297#_c_394_n 0.0173206f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_c_124_n N_A_27_297#_c_394_n 0.0170871f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A_c_121_n N_A_27_297#_c_394_n 0.0472209f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A_c_122_n N_A_27_297#_c_394_n 0.00845817f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_124 N_A_c_125_n N_A_27_297#_c_395_n 0.0170871f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A_c_126_n N_A_27_297#_c_395_n 0.0170871f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A_c_121_n N_A_27_297#_c_395_n 0.047182f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A_c_122_n N_A_27_297#_c_395_n 0.00873423f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_128 N_A_c_127_n N_A_27_297#_c_396_n 0.0170871f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_c_128_n N_A_27_297#_c_396_n 0.0170871f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_c_121_n N_A_27_297#_c_396_n 0.047182f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_c_122_n N_A_27_297#_c_396_n 0.00873423f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_132 N_A_c_129_n N_A_27_297#_c_397_n 0.0170871f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A_c_130_n N_A_27_297#_c_397_n 0.0170264f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_c_121_n N_A_27_297#_c_397_n 0.0472209f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_c_122_n N_A_27_297#_c_397_n 0.00825244f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_136 N_A_c_121_n N_A_27_297#_c_398_n 0.0012302f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_c_121_n N_A_27_297#_c_399_n 0.019528f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_c_122_n N_A_27_297#_c_399_n 0.00661013f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_139 N_A_c_121_n N_A_27_297#_c_400_n 0.019528f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A_c_122_n N_A_27_297#_c_400_n 0.00661013f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_141 N_A_c_121_n N_A_27_297#_c_401_n 0.019528f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_c_122_n N_A_27_297#_c_401_n 0.00661013f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_143 N_A_c_123_n N_VPWR_c_496_n 0.00300743f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_124_n N_VPWR_c_496_n 0.00300743f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_c_124_n N_VPWR_c_497_n 0.00702461f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_c_125_n N_VPWR_c_497_n 0.00702461f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_c_125_n N_VPWR_c_498_n 0.00300743f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_c_126_n N_VPWR_c_498_n 0.00300743f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_c_126_n N_VPWR_c_499_n 0.00702461f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_c_127_n N_VPWR_c_499_n 0.00702461f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_c_127_n N_VPWR_c_500_n 0.00300743f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_c_128_n N_VPWR_c_500_n 0.00300743f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_c_128_n N_VPWR_c_501_n 0.00702461f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_c_129_n N_VPWR_c_501_n 0.00702461f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_c_129_n N_VPWR_c_502_n 0.00300743f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_c_130_n N_VPWR_c_502_n 0.00300743f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_c_130_n N_VPWR_c_503_n 0.00702461f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_c_123_n N_VPWR_c_495_n 0.0133387f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_c_124_n N_VPWR_c_495_n 0.0124092f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A_c_125_n N_VPWR_c_495_n 0.0124092f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A_c_126_n N_VPWR_c_495_n 0.0124092f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_c_127_n N_VPWR_c_495_n 0.0124092f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A_c_128_n N_VPWR_c_495_n 0.0124092f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_c_129_n N_VPWR_c_495_n 0.0124092f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A_c_130_n N_VPWR_c_495_n 0.0124344f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_c_123_n N_VPWR_c_505_n 0.00702461f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_c_113_n N_Y_c_617_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_c_114_n N_Y_c_617_n 0.00686626f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_c_115_n N_Y_c_617_n 5.45498e-19 $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_c_114_n N_Y_c_594_n 0.00901745f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A_c_115_n N_Y_c_594_n 0.00901745f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_c_121_n N_Y_c_594_n 0.0397461f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_c_122_n N_Y_c_594_n 0.00345541f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_174 N_A_c_113_n N_Y_c_595_n 0.00266157f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A_c_114_n N_Y_c_595_n 0.00116636f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_c_121_n N_Y_c_595_n 0.0306016f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_c_122_n N_Y_c_595_n 0.00358305f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_178 N_A_c_114_n N_Y_c_628_n 5.24597e-19 $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_c_115_n N_Y_c_628_n 0.00651696f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_c_116_n N_Y_c_628_n 0.00686626f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_c_117_n N_Y_c_628_n 5.45498e-19 $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_c_116_n N_Y_c_596_n 0.00901745f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_c_117_n N_Y_c_596_n 0.00901745f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_c_121_n N_Y_c_596_n 0.0397461f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_c_122_n N_Y_c_596_n 0.00345541f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_186 N_A_c_116_n N_Y_c_636_n 5.24597e-19 $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_c_117_n N_Y_c_636_n 0.00651696f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_c_118_n N_Y_c_636_n 0.00686626f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_c_119_n N_Y_c_636_n 5.45498e-19 $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_c_118_n N_Y_c_597_n 0.00901745f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_c_119_n N_Y_c_597_n 0.00901745f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_c_121_n N_Y_c_597_n 0.0397461f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_c_122_n N_Y_c_597_n 0.00345541f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_194 N_A_c_118_n N_Y_c_644_n 5.24597e-19 $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_c_119_n N_Y_c_644_n 0.00651696f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_c_120_n N_Y_c_598_n 0.0106151f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_c_121_n N_Y_c_598_n 0.0136715f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A_c_120_n N_Y_c_648_n 5.32212e-19 $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_c_115_n N_Y_c_602_n 0.00116636f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_c_116_n N_Y_c_602_n 0.00116636f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_c_121_n N_Y_c_602_n 0.0306016f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_202 N_A_c_122_n N_Y_c_602_n 0.00358305f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_203 N_A_c_117_n N_Y_c_603_n 0.00116636f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A_c_118_n N_Y_c_603_n 0.00116636f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A_c_121_n N_Y_c_603_n 0.0306016f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A_c_122_n N_Y_c_603_n 0.00358305f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_207 N_A_c_119_n N_Y_c_604_n 0.00119564f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A_c_121_n N_Y_c_604_n 0.0307352f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A_c_122_n N_Y_c_604_n 0.00486271f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_210 N_A_c_113_n N_VGND_c_818_n 0.00496762f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A_c_113_n N_VGND_c_819_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A_c_114_n N_VGND_c_819_n 0.00423334f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A_c_114_n N_VGND_c_820_n 0.00379224f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A_c_115_n N_VGND_c_820_n 0.00276126f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A_c_116_n N_VGND_c_821_n 0.00379224f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A_c_117_n N_VGND_c_821_n 0.00276126f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A_c_118_n N_VGND_c_822_n 0.00379224f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A_c_119_n N_VGND_c_822_n 0.00276126f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A_c_120_n N_VGND_c_823_n 0.00268723f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_c_115_n N_VGND_c_828_n 0.00423334f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A_c_116_n N_VGND_c_828_n 0.00423334f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A_c_117_n N_VGND_c_830_n 0.00423334f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A_c_118_n N_VGND_c_830_n 0.00423334f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A_c_119_n N_VGND_c_832_n 0.00423334f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A_c_120_n N_VGND_c_832_n 0.00437852f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A_c_113_n N_VGND_c_843_n 0.0106014f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A_c_114_n N_VGND_c_843_n 0.006093f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A_c_115_n N_VGND_c_843_n 0.00597024f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A_c_116_n N_VGND_c_843_n 0.006093f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A_c_117_n N_VGND_c_843_n 0.00597024f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A_c_118_n N_VGND_c_843_n 0.006093f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_c_119_n N_VGND_c_843_n 0.00608558f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_c_120_n N_VGND_c_843_n 0.00615622f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_234 N_B_c_262_n N_A_27_297#_c_398_n 2.98195e-19 $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_235 N_B_c_262_n N_A_27_297#_c_427_n 0.0143578f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_236 N_B_c_263_n N_A_27_297#_c_427_n 0.0143578f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_237 N_B_c_264_n N_A_27_297#_c_429_n 0.0143578f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_238 N_B_c_265_n N_A_27_297#_c_429_n 0.0143578f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_239 N_B_c_266_n N_A_27_297#_c_431_n 0.0143578f $X=6.155 $Y=1.41 $X2=0 $Y2=0
cc_240 N_B_c_267_n N_A_27_297#_c_431_n 0.0143578f $X=6.625 $Y=1.41 $X2=0 $Y2=0
cc_241 N_B_c_268_n N_A_27_297#_c_433_n 0.0143578f $X=7.095 $Y=1.41 $X2=0 $Y2=0
cc_242 N_B_c_269_n N_A_27_297#_c_433_n 0.0143578f $X=7.565 $Y=1.41 $X2=0 $Y2=0
cc_243 N_B_c_262_n N_VPWR_c_503_n 0.00429453f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_244 N_B_c_263_n N_VPWR_c_503_n 0.00429453f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_245 N_B_c_264_n N_VPWR_c_503_n 0.00429453f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_246 N_B_c_265_n N_VPWR_c_503_n 0.00429453f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_247 N_B_c_266_n N_VPWR_c_503_n 0.00429453f $X=6.155 $Y=1.41 $X2=0 $Y2=0
cc_248 N_B_c_267_n N_VPWR_c_503_n 0.00429453f $X=6.625 $Y=1.41 $X2=0 $Y2=0
cc_249 N_B_c_268_n N_VPWR_c_503_n 0.00429453f $X=7.095 $Y=1.41 $X2=0 $Y2=0
cc_250 N_B_c_269_n N_VPWR_c_503_n 0.00429453f $X=7.565 $Y=1.41 $X2=0 $Y2=0
cc_251 N_B_c_262_n N_VPWR_c_495_n 0.00609021f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_252 N_B_c_263_n N_VPWR_c_495_n 0.00606499f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_253 N_B_c_264_n N_VPWR_c_495_n 0.00606499f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_254 N_B_c_265_n N_VPWR_c_495_n 0.00606499f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_255 N_B_c_266_n N_VPWR_c_495_n 0.00606499f $X=6.155 $Y=1.41 $X2=0 $Y2=0
cc_256 N_B_c_267_n N_VPWR_c_495_n 0.00606499f $X=6.625 $Y=1.41 $X2=0 $Y2=0
cc_257 N_B_c_268_n N_VPWR_c_495_n 0.00606499f $X=7.095 $Y=1.41 $X2=0 $Y2=0
cc_258 N_B_c_269_n N_VPWR_c_495_n 0.00712629f $X=7.565 $Y=1.41 $X2=0 $Y2=0
cc_259 N_B_c_253_n N_Y_c_598_n 0.00940242f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_260 N_B_c_273_n N_Y_c_598_n 0.00651491f $X=7.055 $Y=1.16 $X2=0 $Y2=0
cc_261 N_B_c_253_n N_Y_c_648_n 0.00644736f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_262 N_B_c_254_n N_Y_c_648_n 0.00686626f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_263 N_B_c_255_n N_Y_c_648_n 5.45498e-19 $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_264 N_B_c_263_n N_Y_c_610_n 0.015669f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_265 N_B_c_264_n N_Y_c_610_n 0.0157513f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_266 N_B_c_273_n N_Y_c_610_n 0.0485189f $X=7.055 $Y=1.16 $X2=0 $Y2=0
cc_267 N_B_c_261_n N_Y_c_610_n 0.00875187f $X=7.565 $Y=1.202 $X2=0 $Y2=0
cc_268 N_B_c_262_n N_Y_c_611_n 6.32035e-19 $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_269 N_B_c_273_n N_Y_c_611_n 0.020385f $X=7.055 $Y=1.16 $X2=0 $Y2=0
cc_270 N_B_c_261_n N_Y_c_611_n 0.00663436f $X=7.565 $Y=1.202 $X2=0 $Y2=0
cc_271 N_B_c_254_n N_Y_c_599_n 0.00901745f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_272 N_B_c_255_n N_Y_c_599_n 0.00901745f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_273 N_B_c_273_n N_Y_c_599_n 0.0397461f $X=7.055 $Y=1.16 $X2=0 $Y2=0
cc_274 N_B_c_261_n N_Y_c_599_n 0.00345541f $X=7.565 $Y=1.202 $X2=0 $Y2=0
cc_275 N_B_c_254_n N_Y_c_676_n 5.24597e-19 $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_276 N_B_c_255_n N_Y_c_676_n 0.00651696f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_277 N_B_c_256_n N_Y_c_676_n 0.00686626f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_278 N_B_c_257_n N_Y_c_676_n 5.45498e-19 $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_279 N_B_c_265_n N_Y_c_612_n 0.0157513f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_280 N_B_c_266_n N_Y_c_612_n 0.0157513f $X=6.155 $Y=1.41 $X2=0 $Y2=0
cc_281 N_B_c_273_n N_Y_c_612_n 0.0485189f $X=7.055 $Y=1.16 $X2=0 $Y2=0
cc_282 N_B_c_261_n N_Y_c_612_n 0.00875187f $X=7.565 $Y=1.202 $X2=0 $Y2=0
cc_283 N_B_c_256_n N_Y_c_600_n 0.00901745f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_284 N_B_c_257_n N_Y_c_600_n 0.00901745f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_285 N_B_c_273_n N_Y_c_600_n 0.0397461f $X=7.055 $Y=1.16 $X2=0 $Y2=0
cc_286 N_B_c_261_n N_Y_c_600_n 0.00345541f $X=7.565 $Y=1.202 $X2=0 $Y2=0
cc_287 N_B_c_256_n N_Y_c_688_n 5.24597e-19 $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_288 N_B_c_257_n N_Y_c_688_n 0.00651696f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_289 N_B_c_258_n N_Y_c_688_n 0.00686352f $X=6.6 $Y=0.995 $X2=0 $Y2=0
cc_290 N_B_c_259_n N_Y_c_688_n 5.45311e-19 $X=7.07 $Y=0.995 $X2=0 $Y2=0
cc_291 N_B_c_267_n N_Y_c_613_n 0.0157513f $X=6.625 $Y=1.41 $X2=0 $Y2=0
cc_292 N_B_c_268_n N_Y_c_613_n 0.0157513f $X=7.095 $Y=1.41 $X2=0 $Y2=0
cc_293 N_B_c_273_n N_Y_c_613_n 0.0485189f $X=7.055 $Y=1.16 $X2=0 $Y2=0
cc_294 N_B_c_261_n N_Y_c_613_n 0.00875187f $X=7.565 $Y=1.202 $X2=0 $Y2=0
cc_295 N_B_c_258_n N_Y_c_601_n 0.00901745f $X=6.6 $Y=0.995 $X2=0 $Y2=0
cc_296 N_B_c_259_n N_Y_c_601_n 0.00901745f $X=7.07 $Y=0.995 $X2=0 $Y2=0
cc_297 N_B_c_273_n N_Y_c_601_n 0.0397461f $X=7.055 $Y=1.16 $X2=0 $Y2=0
cc_298 N_B_c_261_n N_Y_c_601_n 0.00345541f $X=7.565 $Y=1.202 $X2=0 $Y2=0
cc_299 N_B_c_253_n N_Y_c_605_n 0.00116636f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_300 N_B_c_254_n N_Y_c_605_n 0.00116636f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_301 N_B_c_273_n N_Y_c_605_n 0.0306016f $X=7.055 $Y=1.16 $X2=0 $Y2=0
cc_302 N_B_c_261_n N_Y_c_605_n 0.00358305f $X=7.565 $Y=1.202 $X2=0 $Y2=0
cc_303 N_B_c_255_n N_Y_c_606_n 0.00116636f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_304 N_B_c_256_n N_Y_c_606_n 0.00116636f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_305 N_B_c_273_n N_Y_c_606_n 0.0306016f $X=7.055 $Y=1.16 $X2=0 $Y2=0
cc_306 N_B_c_261_n N_Y_c_606_n 0.00358305f $X=7.565 $Y=1.202 $X2=0 $Y2=0
cc_307 N_B_c_273_n N_Y_c_614_n 0.020385f $X=7.055 $Y=1.16 $X2=0 $Y2=0
cc_308 N_B_c_261_n N_Y_c_614_n 0.00663436f $X=7.565 $Y=1.202 $X2=0 $Y2=0
cc_309 N_B_c_257_n N_Y_c_607_n 0.00116636f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_310 N_B_c_258_n N_Y_c_607_n 0.00116636f $X=6.6 $Y=0.995 $X2=0 $Y2=0
cc_311 N_B_c_273_n N_Y_c_607_n 0.0306016f $X=7.055 $Y=1.16 $X2=0 $Y2=0
cc_312 N_B_c_261_n N_Y_c_607_n 0.00358305f $X=7.565 $Y=1.202 $X2=0 $Y2=0
cc_313 N_B_c_273_n N_Y_c_615_n 0.020385f $X=7.055 $Y=1.16 $X2=0 $Y2=0
cc_314 N_B_c_261_n N_Y_c_615_n 0.00663436f $X=7.565 $Y=1.202 $X2=0 $Y2=0
cc_315 N_B_c_258_n N_Y_c_608_n 5.25778e-19 $X=6.6 $Y=0.995 $X2=0 $Y2=0
cc_316 N_B_c_259_n N_Y_c_608_n 0.00777632f $X=7.07 $Y=0.995 $X2=0 $Y2=0
cc_317 N_B_c_260_n N_Y_c_608_n 0.0103608f $X=7.59 $Y=0.995 $X2=0 $Y2=0
cc_318 N_B_c_273_n N_Y_c_608_n 0.0140822f $X=7.055 $Y=1.16 $X2=0 $Y2=0
cc_319 N_B_c_261_n N_Y_c_608_n 0.0056758f $X=7.565 $Y=1.202 $X2=0 $Y2=0
cc_320 N_B_c_259_n Y 9.09931e-19 $X=7.07 $Y=0.995 $X2=0 $Y2=0
cc_321 N_B_c_269_n Y 0.0178942f $X=7.565 $Y=1.41 $X2=0 $Y2=0
cc_322 N_B_c_260_n Y 0.00407608f $X=7.59 $Y=0.995 $X2=0 $Y2=0
cc_323 N_B_c_273_n Y 0.0233758f $X=7.055 $Y=1.16 $X2=0 $Y2=0
cc_324 N_B_c_261_n Y 0.0361146f $X=7.565 $Y=1.202 $X2=0 $Y2=0
cc_325 N_B_c_253_n N_VGND_c_823_n 0.00268723f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_326 N_B_c_254_n N_VGND_c_824_n 0.00379224f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_327 N_B_c_255_n N_VGND_c_824_n 0.00276126f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_328 N_B_c_256_n N_VGND_c_825_n 0.00379224f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_329 N_B_c_257_n N_VGND_c_825_n 0.00276126f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_330 N_B_c_258_n N_VGND_c_826_n 0.00379224f $X=6.6 $Y=0.995 $X2=0 $Y2=0
cc_331 N_B_c_259_n N_VGND_c_826_n 0.00276126f $X=7.07 $Y=0.995 $X2=0 $Y2=0
cc_332 N_B_c_260_n N_VGND_c_827_n 0.0045387f $X=7.59 $Y=0.995 $X2=0 $Y2=0
cc_333 N_B_c_253_n N_VGND_c_834_n 0.00423334f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_334 N_B_c_254_n N_VGND_c_834_n 0.00423334f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_335 N_B_c_255_n N_VGND_c_836_n 0.00423334f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_336 N_B_c_256_n N_VGND_c_836_n 0.00423334f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_337 N_B_c_257_n N_VGND_c_838_n 0.00423334f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_338 N_B_c_258_n N_VGND_c_838_n 0.00423334f $X=6.6 $Y=0.995 $X2=0 $Y2=0
cc_339 N_B_c_259_n N_VGND_c_841_n 0.00421816f $X=7.07 $Y=0.995 $X2=0 $Y2=0
cc_340 N_B_c_260_n N_VGND_c_841_n 0.00437716f $X=7.59 $Y=0.995 $X2=0 $Y2=0
cc_341 N_B_c_253_n N_VGND_c_843_n 0.00587047f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_342 N_B_c_254_n N_VGND_c_843_n 0.006093f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_343 N_B_c_255_n N_VGND_c_843_n 0.00597024f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_344 N_B_c_256_n N_VGND_c_843_n 0.006093f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_345 N_B_c_257_n N_VGND_c_843_n 0.00597024f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_346 N_B_c_258_n N_VGND_c_843_n 0.006093f $X=6.6 $Y=0.995 $X2=0 $Y2=0
cc_347 N_B_c_259_n N_VGND_c_843_n 0.00609466f $X=7.07 $Y=0.995 $X2=0 $Y2=0
cc_348 N_B_c_260_n N_VGND_c_843_n 0.00723526f $X=7.59 $Y=0.995 $X2=0 $Y2=0
cc_349 N_A_27_297#_c_394_n N_VPWR_M1001_d 0.00188315f $X=1.095 $Y=1.56 $X2=-0.19
+ $Y2=1.305
cc_350 N_A_27_297#_c_395_n N_VPWR_M1008_d 0.00188315f $X=2.035 $Y=1.56 $X2=0
+ $Y2=0
cc_351 N_A_27_297#_c_396_n N_VPWR_M1018_d 0.00188315f $X=2.975 $Y=1.56 $X2=0
+ $Y2=0
cc_352 N_A_27_297#_c_397_n N_VPWR_M1026_d 0.00188315f $X=3.915 $Y=1.56 $X2=0
+ $Y2=0
cc_353 N_A_27_297#_c_394_n N_VPWR_c_496_n 0.0145257f $X=1.095 $Y=1.56 $X2=0
+ $Y2=0
cc_354 N_A_27_297#_c_440_p N_VPWR_c_497_n 0.0149311f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_355 N_A_27_297#_c_395_n N_VPWR_c_498_n 0.0145257f $X=2.035 $Y=1.56 $X2=0
+ $Y2=0
cc_356 N_A_27_297#_c_442_p N_VPWR_c_499_n 0.0149311f $X=2.16 $Y=2.3 $X2=0 $Y2=0
cc_357 N_A_27_297#_c_396_n N_VPWR_c_500_n 0.0145257f $X=2.975 $Y=1.56 $X2=0
+ $Y2=0
cc_358 N_A_27_297#_c_444_p N_VPWR_c_501_n 0.0149311f $X=3.1 $Y=2.3 $X2=0 $Y2=0
cc_359 N_A_27_297#_c_397_n N_VPWR_c_502_n 0.0145257f $X=3.915 $Y=1.56 $X2=0
+ $Y2=0
cc_360 N_A_27_297#_c_446_p N_VPWR_c_503_n 0.015002f $X=4.04 $Y=2.295 $X2=0 $Y2=0
cc_361 N_A_27_297#_c_427_n N_VPWR_c_503_n 0.0386815f $X=4.855 $Y=2.38 $X2=0
+ $Y2=0
cc_362 N_A_27_297#_c_429_n N_VPWR_c_503_n 0.0386815f $X=5.795 $Y=2.38 $X2=0
+ $Y2=0
cc_363 N_A_27_297#_c_431_n N_VPWR_c_503_n 0.0386815f $X=6.735 $Y=2.38 $X2=0
+ $Y2=0
cc_364 N_A_27_297#_c_433_n N_VPWR_c_503_n 0.0549726f $X=7.675 $Y=2.38 $X2=0
+ $Y2=0
cc_365 N_A_27_297#_c_451_p N_VPWR_c_503_n 0.015002f $X=4.98 $Y=2.38 $X2=0 $Y2=0
cc_366 N_A_27_297#_c_452_p N_VPWR_c_503_n 0.015002f $X=5.92 $Y=2.38 $X2=0 $Y2=0
cc_367 N_A_27_297#_c_453_p N_VPWR_c_503_n 0.015002f $X=6.86 $Y=2.38 $X2=0 $Y2=0
cc_368 N_A_27_297#_M1001_s N_VPWR_c_495_n 0.00303344f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_369 N_A_27_297#_M1002_s N_VPWR_c_495_n 0.00370124f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_370 N_A_27_297#_M1013_s N_VPWR_c_495_n 0.00370124f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_371 N_A_27_297#_M1021_s N_VPWR_c_495_n 0.00370124f $X=2.955 $Y=1.485 $X2=0
+ $Y2=0
cc_372 N_A_27_297#_M1030_s N_VPWR_c_495_n 0.00297222f $X=3.895 $Y=1.485 $X2=0
+ $Y2=0
cc_373 N_A_27_297#_M1006_s N_VPWR_c_495_n 0.00231264f $X=4.835 $Y=1.485 $X2=0
+ $Y2=0
cc_374 N_A_27_297#_M1011_s N_VPWR_c_495_n 0.00231264f $X=5.775 $Y=1.485 $X2=0
+ $Y2=0
cc_375 N_A_27_297#_M1019_s N_VPWR_c_495_n 0.00231264f $X=6.715 $Y=1.485 $X2=0
+ $Y2=0
cc_376 N_A_27_297#_M1029_s N_VPWR_c_495_n 0.00260432f $X=7.655 $Y=1.485 $X2=0
+ $Y2=0
cc_377 N_A_27_297#_c_393_n N_VPWR_c_495_n 0.0120542f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_378 N_A_27_297#_c_440_p N_VPWR_c_495_n 0.00955092f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_379 N_A_27_297#_c_442_p N_VPWR_c_495_n 0.00955092f $X=2.16 $Y=2.3 $X2=0 $Y2=0
cc_380 N_A_27_297#_c_444_p N_VPWR_c_495_n 0.00955092f $X=3.1 $Y=2.3 $X2=0 $Y2=0
cc_381 N_A_27_297#_c_446_p N_VPWR_c_495_n 0.00962794f $X=4.04 $Y=2.295 $X2=0
+ $Y2=0
cc_382 N_A_27_297#_c_427_n N_VPWR_c_495_n 0.0239144f $X=4.855 $Y=2.38 $X2=0
+ $Y2=0
cc_383 N_A_27_297#_c_429_n N_VPWR_c_495_n 0.0239144f $X=5.795 $Y=2.38 $X2=0
+ $Y2=0
cc_384 N_A_27_297#_c_431_n N_VPWR_c_495_n 0.0239144f $X=6.735 $Y=2.38 $X2=0
+ $Y2=0
cc_385 N_A_27_297#_c_433_n N_VPWR_c_495_n 0.0335424f $X=7.675 $Y=2.38 $X2=0
+ $Y2=0
cc_386 N_A_27_297#_c_451_p N_VPWR_c_495_n 0.00962794f $X=4.98 $Y=2.38 $X2=0
+ $Y2=0
cc_387 N_A_27_297#_c_452_p N_VPWR_c_495_n 0.00962794f $X=5.92 $Y=2.38 $X2=0
+ $Y2=0
cc_388 N_A_27_297#_c_453_p N_VPWR_c_495_n 0.00962794f $X=6.86 $Y=2.38 $X2=0
+ $Y2=0
cc_389 N_A_27_297#_c_393_n N_VPWR_c_505_n 0.0208166f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_390 N_A_27_297#_c_427_n N_Y_M1003_d 0.00352392f $X=4.855 $Y=2.38 $X2=0 $Y2=0
cc_391 N_A_27_297#_c_429_n N_Y_M1009_d 0.00352392f $X=5.795 $Y=2.38 $X2=0 $Y2=0
cc_392 N_A_27_297#_c_431_n N_Y_M1015_d 0.00352392f $X=6.735 $Y=2.38 $X2=0 $Y2=0
cc_393 N_A_27_297#_c_433_n N_Y_M1024_d 0.00352392f $X=7.675 $Y=2.38 $X2=0 $Y2=0
cc_394 N_A_27_297#_c_398_n N_Y_c_598_n 0.0088033f $X=4.04 $Y=1.665 $X2=0 $Y2=0
cc_395 N_A_27_297#_c_427_n N_Y_c_731_n 0.0134104f $X=4.855 $Y=2.38 $X2=0 $Y2=0
cc_396 N_A_27_297#_M1006_s N_Y_c_610_n 0.00187091f $X=4.835 $Y=1.485 $X2=0 $Y2=0
cc_397 N_A_27_297#_c_483_p N_Y_c_610_n 0.0143191f $X=4.98 $Y=1.96 $X2=0 $Y2=0
cc_398 N_A_27_297#_c_398_n N_Y_c_611_n 0.00226124f $X=4.04 $Y=1.665 $X2=0 $Y2=0
cc_399 N_A_27_297#_c_429_n N_Y_c_735_n 0.0134104f $X=5.795 $Y=2.38 $X2=0 $Y2=0
cc_400 N_A_27_297#_M1011_s N_Y_c_612_n 0.00187091f $X=5.775 $Y=1.485 $X2=0 $Y2=0
cc_401 N_A_27_297#_c_487_p N_Y_c_612_n 0.0143191f $X=5.92 $Y=1.96 $X2=0 $Y2=0
cc_402 N_A_27_297#_c_431_n N_Y_c_738_n 0.0134104f $X=6.735 $Y=2.38 $X2=0 $Y2=0
cc_403 N_A_27_297#_M1019_s N_Y_c_613_n 0.00187091f $X=6.715 $Y=1.485 $X2=0 $Y2=0
cc_404 N_A_27_297#_c_490_p N_Y_c_613_n 0.0143191f $X=6.86 $Y=1.96 $X2=0 $Y2=0
cc_405 N_A_27_297#_c_433_n N_Y_c_741_n 0.0134104f $X=7.675 $Y=2.38 $X2=0 $Y2=0
cc_406 N_A_27_297#_M1029_s Y 0.0035037f $X=7.655 $Y=1.485 $X2=0 $Y2=0
cc_407 N_A_27_297#_c_493_p Y 0.0191143f $X=7.8 $Y=1.96 $X2=0 $Y2=0
cc_408 N_A_27_297#_c_392_n N_VGND_c_818_n 0.0111859f $X=0.247 $Y=1.665 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_495_n N_Y_M1003_d 0.00232895f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_410 N_VPWR_c_495_n N_Y_M1009_d 0.00232895f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_411 N_VPWR_c_495_n N_Y_M1015_d 0.00232895f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_412 N_VPWR_c_495_n N_Y_M1024_d 0.00232895f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_413 N_Y_c_594_n N_VGND_M1010_d 0.00251047f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_414 N_Y_c_596_n N_VGND_M1016_d 0.00251047f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_415 N_Y_c_597_n N_VGND_M1025_d 0.00251047f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_416 N_Y_c_598_n N_VGND_M1028_d 0.00162089f $X=4.295 $Y=0.815 $X2=0 $Y2=0
cc_417 N_Y_c_599_n N_VGND_M1005_s 0.00251047f $X=5.235 $Y=0.815 $X2=0 $Y2=0
cc_418 N_Y_c_600_n N_VGND_M1014_s 0.00251047f $X=6.175 $Y=0.815 $X2=0 $Y2=0
cc_419 N_Y_c_601_n N_VGND_M1020_s 0.00251047f $X=7.115 $Y=0.815 $X2=0 $Y2=0
cc_420 N_Y_c_608_n N_VGND_M1031_s 0.00290026f $X=7.33 $Y=0.39 $X2=0 $Y2=0
cc_421 N_Y_c_595_n N_VGND_c_818_n 0.00835456f $X=0.915 $Y=0.815 $X2=0 $Y2=0
cc_422 N_Y_c_617_n N_VGND_c_819_n 0.0223596f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_423 N_Y_c_594_n N_VGND_c_819_n 0.00266636f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_424 N_Y_c_617_n N_VGND_c_820_n 0.0183628f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_425 N_Y_c_594_n N_VGND_c_820_n 0.0127273f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_426 N_Y_c_628_n N_VGND_c_821_n 0.0183628f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_427 N_Y_c_596_n N_VGND_c_821_n 0.0127273f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_428 N_Y_c_636_n N_VGND_c_822_n 0.0183628f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_429 N_Y_c_597_n N_VGND_c_822_n 0.0127273f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_430 N_Y_c_598_n N_VGND_c_823_n 0.0122559f $X=4.295 $Y=0.815 $X2=0 $Y2=0
cc_431 N_Y_c_648_n N_VGND_c_824_n 0.0183628f $X=4.51 $Y=0.39 $X2=0 $Y2=0
cc_432 N_Y_c_599_n N_VGND_c_824_n 0.0127273f $X=5.235 $Y=0.815 $X2=0 $Y2=0
cc_433 N_Y_c_676_n N_VGND_c_825_n 0.0183628f $X=5.45 $Y=0.39 $X2=0 $Y2=0
cc_434 N_Y_c_600_n N_VGND_c_825_n 0.0127273f $X=6.175 $Y=0.815 $X2=0 $Y2=0
cc_435 N_Y_c_688_n N_VGND_c_826_n 0.0183628f $X=6.39 $Y=0.39 $X2=0 $Y2=0
cc_436 N_Y_c_601_n N_VGND_c_826_n 0.0127273f $X=7.115 $Y=0.815 $X2=0 $Y2=0
cc_437 N_Y_c_608_n N_VGND_c_827_n 0.0246547f $X=7.33 $Y=0.39 $X2=0 $Y2=0
cc_438 N_Y_c_594_n N_VGND_c_828_n 0.00198695f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_439 N_Y_c_628_n N_VGND_c_828_n 0.0223596f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_440 N_Y_c_596_n N_VGND_c_828_n 0.00266636f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_441 N_Y_c_596_n N_VGND_c_830_n 0.00198695f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_442 N_Y_c_636_n N_VGND_c_830_n 0.0223596f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_443 N_Y_c_597_n N_VGND_c_830_n 0.00266636f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_444 N_Y_c_597_n N_VGND_c_832_n 0.00198695f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_445 N_Y_c_644_n N_VGND_c_832_n 0.0231806f $X=3.57 $Y=0.39 $X2=0 $Y2=0
cc_446 N_Y_c_598_n N_VGND_c_832_n 0.00254521f $X=4.295 $Y=0.815 $X2=0 $Y2=0
cc_447 N_Y_c_598_n N_VGND_c_834_n 0.00198695f $X=4.295 $Y=0.815 $X2=0 $Y2=0
cc_448 N_Y_c_648_n N_VGND_c_834_n 0.0223596f $X=4.51 $Y=0.39 $X2=0 $Y2=0
cc_449 N_Y_c_599_n N_VGND_c_834_n 0.00266636f $X=5.235 $Y=0.815 $X2=0 $Y2=0
cc_450 N_Y_c_599_n N_VGND_c_836_n 0.00198695f $X=5.235 $Y=0.815 $X2=0 $Y2=0
cc_451 N_Y_c_676_n N_VGND_c_836_n 0.0223596f $X=5.45 $Y=0.39 $X2=0 $Y2=0
cc_452 N_Y_c_600_n N_VGND_c_836_n 0.00266636f $X=6.175 $Y=0.815 $X2=0 $Y2=0
cc_453 N_Y_c_600_n N_VGND_c_838_n 0.00198695f $X=6.175 $Y=0.815 $X2=0 $Y2=0
cc_454 N_Y_c_688_n N_VGND_c_838_n 0.0223596f $X=6.39 $Y=0.39 $X2=0 $Y2=0
cc_455 N_Y_c_601_n N_VGND_c_838_n 0.00266636f $X=7.115 $Y=0.815 $X2=0 $Y2=0
cc_456 N_Y_c_608_n N_VGND_c_840_n 3.327e-19 $X=7.33 $Y=0.39 $X2=0 $Y2=0
cc_457 N_Y_c_601_n N_VGND_c_841_n 0.00198695f $X=7.115 $Y=0.815 $X2=0 $Y2=0
cc_458 N_Y_c_608_n N_VGND_c_841_n 0.0260268f $X=7.33 $Y=0.39 $X2=0 $Y2=0
cc_459 N_Y_M1004_s N_VGND_c_843_n 0.0025535f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_460 N_Y_M1012_s N_VGND_c_843_n 0.0025535f $X=1.505 $Y=0.235 $X2=0 $Y2=0
cc_461 N_Y_M1022_s N_VGND_c_843_n 0.0025535f $X=2.445 $Y=0.235 $X2=0 $Y2=0
cc_462 N_Y_M1027_s N_VGND_c_843_n 0.00304143f $X=3.385 $Y=0.235 $X2=0 $Y2=0
cc_463 N_Y_M1000_d N_VGND_c_843_n 0.0025535f $X=4.325 $Y=0.235 $X2=0 $Y2=0
cc_464 N_Y_M1007_d N_VGND_c_843_n 0.0025535f $X=5.265 $Y=0.235 $X2=0 $Y2=0
cc_465 N_Y_M1017_d N_VGND_c_843_n 0.0025535f $X=6.205 $Y=0.235 $X2=0 $Y2=0
cc_466 N_Y_M1023_d N_VGND_c_843_n 0.00304917f $X=7.145 $Y=0.235 $X2=0 $Y2=0
cc_467 N_Y_c_617_n N_VGND_c_843_n 0.0141302f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_468 N_Y_c_594_n N_VGND_c_843_n 0.00972452f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_469 N_Y_c_628_n N_VGND_c_843_n 0.0141302f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_470 N_Y_c_596_n N_VGND_c_843_n 0.00972452f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_471 N_Y_c_636_n N_VGND_c_843_n 0.0141302f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_472 N_Y_c_597_n N_VGND_c_843_n 0.00972452f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_473 N_Y_c_644_n N_VGND_c_843_n 0.0143352f $X=3.57 $Y=0.39 $X2=0 $Y2=0
cc_474 N_Y_c_598_n N_VGND_c_843_n 0.0094839f $X=4.295 $Y=0.815 $X2=0 $Y2=0
cc_475 N_Y_c_648_n N_VGND_c_843_n 0.0141302f $X=4.51 $Y=0.39 $X2=0 $Y2=0
cc_476 N_Y_c_599_n N_VGND_c_843_n 0.00972452f $X=5.235 $Y=0.815 $X2=0 $Y2=0
cc_477 N_Y_c_676_n N_VGND_c_843_n 0.0141302f $X=5.45 $Y=0.39 $X2=0 $Y2=0
cc_478 N_Y_c_600_n N_VGND_c_843_n 0.00972452f $X=6.175 $Y=0.815 $X2=0 $Y2=0
cc_479 N_Y_c_688_n N_VGND_c_843_n 0.0141302f $X=6.39 $Y=0.39 $X2=0 $Y2=0
cc_480 N_Y_c_601_n N_VGND_c_843_n 0.00972452f $X=7.115 $Y=0.815 $X2=0 $Y2=0
cc_481 N_Y_c_608_n N_VGND_c_843_n 0.0215948f $X=7.33 $Y=0.39 $X2=0 $Y2=0
