* File: sky130_fd_sc_hdll__a211oi_1.spice
* Created: Wed Sep  2 08:16:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a211oi_1.pex.spice"
.subckt sky130_fd_sc_hdll__a211oi_1  VNB VPB A2 A1 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1002 A_123_47# N_A2_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.092625 AS=0.2145 PD=0.935 PS=1.96 NRD=16.152 NRS=11.988 M=1 R=4.33333
+ SA=75000.3 SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1006_d N_A1_M1006_g A_123_47# VNB NSHORT L=0.15 W=0.65 AD=0.125125
+ AS=0.092625 PD=1.035 PS=0.935 NRD=9.228 NRS=16.152 M=1 R=4.33333 SA=75000.7
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_B1_M1004_g N_Y_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.112125 AS=0.125125 PD=0.995 PS=1.035 NRD=7.38 NRS=10.152 M=1 R=4.33333
+ SA=75001.2 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1007 N_Y_M1007_d N_C1_M1007_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65 AD=0.26
+ AS=0.112125 PD=2.1 PS=0.995 NRD=24.912 NRS=4.608 M=1 R=4.33333 SA=75001.7
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A2_M1000_g N_A_27_297#_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1525 AS=0.29 PD=1.305 PS=2.58 NRD=2.9353 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1003 N_A_27_297#_M1003_d N_A1_M1003_g N_VPWR_M1000_d VPB PHIGHVT L=0.18 W=1
+ AD=0.1775 AS=0.1525 PD=1.355 PS=1.305 NRD=1.9503 NRS=1.9503 M=1 R=5.55556
+ SA=90000.7 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1005 A_325_297# N_B1_M1005_g N_A_27_297#_M1003_d VPB PHIGHVT L=0.18 W=1
+ AD=0.1575 AS=0.1775 PD=1.315 PS=1.355 NRD=20.1728 NRS=12.7853 M=1 R=5.55556
+ SA=90001.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1001 N_Y_M1001_d N_C1_M1001_g A_325_297# VPB PHIGHVT L=0.18 W=1 AD=0.36
+ AS=0.1575 PD=2.72 PS=1.315 NRD=18.715 NRS=20.1728 M=1 R=5.55556 SA=90001.7
+ SB=90000.3 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
pX9_noxref noxref_13 B1 B1 PROBETYPE=1
pX10_noxref noxref_14 B1 B1 PROBETYPE=1
pX11_noxref noxref_15 B1 B1 PROBETYPE=1
pX12_noxref noxref_16 B1 B1 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__a211oi_1.pxi.spice"
*
.ends
*
*
