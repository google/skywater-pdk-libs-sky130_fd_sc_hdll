* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nand3b_4 A_N B C VGND VNB VPB VPWR Y
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_683_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 a_683_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_27_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 a_225_47# B a_683_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 Y a_27_47# a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 a_225_47# B a_683_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND C a_683_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND C a_683_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 Y a_27_47# a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 a_27_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_225_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 a_683_47# B a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 a_225_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_683_47# B a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
