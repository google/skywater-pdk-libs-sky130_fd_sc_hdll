* File: sky130_fd_sc_hdll__nand3b_2.pxi.spice
* Created: Wed Sep  2 08:38:02 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND3B_2%A_N N_A_N_M1013_g N_A_N_c_75_n N_A_N_c_76_n
+ N_A_N_M1002_g A_N N_A_N_c_74_n A_N PM_SKY130_FD_SC_HDLL__NAND3B_2%A_N
x_PM_SKY130_FD_SC_HDLL__NAND3B_2%C N_C_M1000_g N_C_c_109_n N_C_M1006_g
+ N_C_c_110_n N_C_M1011_g N_C_M1007_g C C N_C_c_108_n C
+ PM_SKY130_FD_SC_HDLL__NAND3B_2%C
x_PM_SKY130_FD_SC_HDLL__NAND3B_2%B N_B_c_156_n N_B_M1003_g N_B_c_157_n
+ N_B_M1012_g N_B_M1004_g N_B_M1005_g N_B_c_153_n N_B_c_154_n B B B B
+ PM_SKY130_FD_SC_HDLL__NAND3B_2%B
x_PM_SKY130_FD_SC_HDLL__NAND3B_2%A_27_47# N_A_27_47#_M1013_s N_A_27_47#_M1002_s
+ N_A_27_47#_M1001_g N_A_27_47#_c_201_n N_A_27_47#_M1008_g N_A_27_47#_c_202_n
+ N_A_27_47#_M1009_g N_A_27_47#_M1010_g N_A_27_47#_c_198_n N_A_27_47#_c_204_n
+ N_A_27_47#_c_205_n N_A_27_47#_c_199_n N_A_27_47#_c_206_n N_A_27_47#_c_207_n
+ N_A_27_47#_c_208_n N_A_27_47#_c_200_n PM_SKY130_FD_SC_HDLL__NAND3B_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NAND3B_2%VPWR N_VPWR_M1002_d N_VPWR_M1011_d
+ N_VPWR_M1012_s N_VPWR_M1008_d N_VPWR_M1009_d N_VPWR_c_283_n N_VPWR_c_284_n
+ N_VPWR_c_285_n N_VPWR_c_286_n N_VPWR_c_287_n N_VPWR_c_288_n N_VPWR_c_289_n
+ N_VPWR_c_290_n N_VPWR_c_291_n N_VPWR_c_292_n N_VPWR_c_293_n N_VPWR_c_294_n
+ VPWR N_VPWR_c_295_n N_VPWR_c_296_n N_VPWR_c_282_n
+ PM_SKY130_FD_SC_HDLL__NAND3B_2%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND3B_2%Y N_Y_M1001_d N_Y_M1006_s N_Y_M1003_d
+ N_Y_M1008_s N_Y_c_366_n N_Y_c_362_n N_Y_c_360_n N_Y_c_363_n N_Y_c_365_n
+ N_Y_c_369_n N_Y_c_390_n Y Y PM_SKY130_FD_SC_HDLL__NAND3B_2%Y
x_PM_SKY130_FD_SC_HDLL__NAND3B_2%VGND N_VGND_M1013_d N_VGND_M1007_d
+ N_VGND_c_435_n N_VGND_c_436_n N_VGND_c_437_n N_VGND_c_438_n VGND
+ N_VGND_c_439_n N_VGND_c_440_n N_VGND_c_441_n VGND
+ PM_SKY130_FD_SC_HDLL__NAND3B_2%VGND
x_PM_SKY130_FD_SC_HDLL__NAND3B_2%A_228_47# N_A_228_47#_M1000_s
+ N_A_228_47#_M1004_s N_A_228_47#_c_495_n N_A_228_47#_c_491_n
+ N_A_228_47#_c_492_n N_A_228_47#_c_493_n N_A_228_47#_c_494_n
+ PM_SKY130_FD_SC_HDLL__NAND3B_2%A_228_47#
x_PM_SKY130_FD_SC_HDLL__NAND3B_2%A_448_47# N_A_448_47#_M1004_d
+ N_A_448_47#_M1005_d N_A_448_47#_M1010_s N_A_448_47#_c_522_n
+ N_A_448_47#_c_523_n N_A_448_47#_c_524_n N_A_448_47#_c_543_n
+ PM_SKY130_FD_SC_HDLL__NAND3B_2%A_448_47#
cc_1 VNB N_A_N_M1013_g 0.0351013f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB A_N 0.00224942f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_3 VNB N_A_N_c_74_n 0.0321034f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_4 VNB N_C_M1000_g 0.0201045f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_5 VNB N_C_M1007_g 0.0249344f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_6 VNB C 0.00593113f $X=-0.19 $Y=-0.24 $X2=0.587 $Y2=1.325
cc_7 VNB N_C_c_108_n 0.039763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_B_M1004_g 0.0244378f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_9 VNB N_B_M1005_g 0.0183135f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_10 VNB N_B_c_153_n 0.0527685f $X=-0.19 $Y=-0.24 $X2=0.587 $Y2=0.995
cc_11 VNB N_B_c_154_n 0.0323772f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.175
cc_12 VNB B 0.00625415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_M1001_g 0.0186958f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_14 VNB N_A_27_47#_M1010_g 0.0218952f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.175
cc_15 VNB N_A_27_47#_c_198_n 0.0308455f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_199_n 0.0188007f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_200_n 0.0434924f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_282_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_Y_c_360_n 0.0217723f $X=-0.19 $Y=-0.24 $X2=0.745 $Y2=1.175
cc_20 VNB Y 0.0207716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_435_n 0.0110084f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_436_n 0.00916027f $X=-0.19 $Y=-0.24 $X2=0.587 $Y2=0.995
cc_23 VNB N_VGND_c_437_n 0.019915f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_438_n 0.00478085f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.175
cc_25 VNB N_VGND_c_439_n 0.0633763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_440_n 0.242894f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_441_n 0.0250348f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_228_47#_c_491_n 0.00263458f $X=-0.19 $Y=-0.24 $X2=0.587 $Y2=1.16
cc_29 VNB N_A_228_47#_c_492_n 0.00280152f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_30 VNB N_A_228_47#_c_493_n 0.00375931f $X=-0.19 $Y=-0.24 $X2=0.587 $Y2=0.995
cc_31 VNB N_A_228_47#_c_494_n 0.0108006f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.175
cc_32 VNB N_A_448_47#_c_522_n 0.00263291f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_33 VNB N_A_448_47#_c_523_n 0.00186742f $X=-0.19 $Y=-0.24 $X2=0.587 $Y2=1.325
cc_34 VNB N_A_448_47#_c_524_n 0.0103948f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_35 VPB N_A_N_c_75_n 0.0379169f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_36 VPB N_A_N_c_76_n 0.0274831f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_37 VPB N_A_N_c_74_n 0.00599428f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_38 VPB N_C_c_109_n 0.0168631f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_39 VPB N_C_c_110_n 0.0160057f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_40 VPB N_C_c_108_n 0.0133458f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_B_c_156_n 0.0160057f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_42 VPB N_B_c_157_n 0.0201091f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_B_c_153_n 0.0160676f $X=-0.19 $Y=1.305 $X2=0.587 $Y2=0.995
cc_44 VPB N_A_27_47#_c_201_n 0.0200795f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_47#_c_202_n 0.0188554f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_46 VPB N_A_27_47#_c_198_n 0.00671796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_27_47#_c_204_n 0.0307013f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_27_47#_c_205_n 0.00136324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_27_47#_c_206_n 0.00770964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_47#_c_207_n 0.0168572f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_c_208_n 0.0214915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_47#_c_200_n 0.0161165f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_283_n 0.00786588f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.19
cc_54 VPB N_VPWR_c_284_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_285_n 0.00636464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_286_n 0.00764677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_287_n 0.0123745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_288_n 0.018317f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_289_n 0.0197985f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_290_n 0.00323937f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_291_n 0.0199879f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_292_n 0.00478085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_293_n 0.00598254f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_294_n 0.00573887f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_295_n 0.0203512f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_296_n 0.0249986f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_282_n 0.0470105f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_Y_c_362_n 0.00859173f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.175
cc_69 VPB N_Y_c_363_n 0.0111887f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB Y 0.0212803f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 N_A_N_M1013_g N_C_M1000_g 0.012851f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_72 N_A_N_c_74_n N_C_M1000_g 0.0230255f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_N_c_75_n N_C_c_109_n 0.01718f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_74 N_A_N_c_76_n N_C_c_109_n 0.0140826f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_75 A_N C 0.0132612f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_76 N_A_N_c_74_n C 2.0081e-19 $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_N_c_75_n N_C_c_108_n 0.00328354f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_78 A_N N_C_c_108_n 0.00145408f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_79 N_A_N_M1013_g N_A_27_47#_c_198_n 0.0231375f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_80 A_N N_A_27_47#_c_198_n 0.0151756f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_81 N_A_N_c_75_n N_A_27_47#_c_204_n 0.0213619f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_82 A_N N_A_27_47#_c_204_n 0.0285273f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_83 N_A_N_c_74_n N_A_27_47#_c_204_n 0.00439952f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_N_M1013_g N_A_27_47#_c_199_n 0.00595292f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_85 N_A_N_c_76_n N_A_27_47#_c_207_n 0.00515834f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_86 N_A_N_c_75_n N_A_27_47#_c_208_n 0.0116827f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_87 N_A_N_c_76_n N_A_27_47#_c_208_n 0.00168084f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_88 N_A_N_c_75_n N_VPWR_c_283_n 0.00201236f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_89 N_A_N_c_76_n N_VPWR_c_283_n 0.00668171f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_90 N_A_N_c_76_n N_VPWR_c_296_n 0.00717092f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_91 N_A_N_c_76_n N_VPWR_c_282_n 0.0138978f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_92 N_A_N_c_75_n N_Y_c_365_n 2.749e-19 $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_93 N_A_N_M1013_g N_VGND_c_435_n 0.0102192f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_94 A_N N_VGND_c_435_n 0.0164192f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_95 N_A_N_c_74_n N_VGND_c_435_n 0.00382571f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_N_M1013_g N_VGND_c_440_n 0.0115873f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A_N_M1013_g N_VGND_c_441_n 0.00564131f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_98 N_C_c_110_n N_B_c_156_n 0.0391101f $X=1.56 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_99 C N_B_c_153_n 0.00234736f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_100 N_C_c_108_n N_B_c_153_n 0.0204203f $X=1.56 $Y=1.217 $X2=0 $Y2=0
cc_101 C B 0.0128159f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_102 N_C_c_109_n N_A_27_47#_c_204_n 0.0177841f $X=1.09 $Y=1.41 $X2=0 $Y2=0
cc_103 N_C_c_110_n N_A_27_47#_c_204_n 0.0118662f $X=1.56 $Y=1.41 $X2=0 $Y2=0
cc_104 C N_A_27_47#_c_204_n 0.059498f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_105 N_C_c_108_n N_A_27_47#_c_204_n 0.00775184f $X=1.56 $Y=1.217 $X2=0 $Y2=0
cc_106 N_C_c_109_n N_VPWR_c_283_n 0.00932674f $X=1.09 $Y=1.41 $X2=0 $Y2=0
cc_107 N_C_c_110_n N_VPWR_c_284_n 0.00402622f $X=1.56 $Y=1.41 $X2=0 $Y2=0
cc_108 N_C_c_109_n N_VPWR_c_289_n 0.00597712f $X=1.09 $Y=1.41 $X2=0 $Y2=0
cc_109 N_C_c_110_n N_VPWR_c_289_n 0.00514793f $X=1.56 $Y=1.41 $X2=0 $Y2=0
cc_110 N_C_c_109_n N_VPWR_c_282_n 0.010376f $X=1.09 $Y=1.41 $X2=0 $Y2=0
cc_111 N_C_c_110_n N_VPWR_c_282_n 0.00680054f $X=1.56 $Y=1.41 $X2=0 $Y2=0
cc_112 N_C_c_110_n N_Y_c_366_n 0.012081f $X=1.56 $Y=1.41 $X2=0 $Y2=0
cc_113 N_C_c_109_n N_Y_c_365_n 0.0120228f $X=1.09 $Y=1.41 $X2=0 $Y2=0
cc_114 N_C_c_110_n N_Y_c_365_n 0.00757084f $X=1.56 $Y=1.41 $X2=0 $Y2=0
cc_115 N_C_c_110_n N_Y_c_369_n 5.5123e-19 $X=1.56 $Y=1.41 $X2=0 $Y2=0
cc_116 N_C_M1000_g N_VGND_c_435_n 0.00329166f $X=1.065 $Y=0.56 $X2=0 $Y2=0
cc_117 N_C_M1007_g N_VGND_c_436_n 0.0044954f $X=1.585 $Y=0.56 $X2=0 $Y2=0
cc_118 N_C_M1000_g N_VGND_c_437_n 0.00541359f $X=1.065 $Y=0.56 $X2=0 $Y2=0
cc_119 N_C_M1007_g N_VGND_c_437_n 0.00436487f $X=1.585 $Y=0.56 $X2=0 $Y2=0
cc_120 N_C_M1000_g N_VGND_c_440_n 0.0101418f $X=1.065 $Y=0.56 $X2=0 $Y2=0
cc_121 N_C_M1007_g N_VGND_c_440_n 0.00743054f $X=1.585 $Y=0.56 $X2=0 $Y2=0
cc_122 N_C_M1000_g N_A_228_47#_c_495_n 0.00514417f $X=1.065 $Y=0.56 $X2=0 $Y2=0
cc_123 N_C_M1000_g N_A_228_47#_c_491_n 0.00274259f $X=1.065 $Y=0.56 $X2=0 $Y2=0
cc_124 C N_A_228_47#_c_491_n 0.0307358f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_125 N_C_c_108_n N_A_228_47#_c_491_n 0.00450572f $X=1.56 $Y=1.217 $X2=0 $Y2=0
cc_126 N_C_M1007_g N_A_228_47#_c_492_n 0.00220648f $X=1.585 $Y=0.56 $X2=0 $Y2=0
cc_127 N_C_M1007_g N_A_228_47#_c_494_n 0.0132378f $X=1.585 $Y=0.56 $X2=0 $Y2=0
cc_128 C N_A_228_47#_c_494_n 0.0294895f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_129 N_B_M1005_g N_A_27_47#_M1001_g 0.0139634f $X=3.095 $Y=0.56 $X2=0 $Y2=0
cc_130 N_B_c_156_n N_A_27_47#_c_204_n 0.0134721f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_131 N_B_c_157_n N_A_27_47#_c_204_n 0.013909f $X=2.5 $Y=1.41 $X2=0 $Y2=0
cc_132 N_B_c_153_n N_A_27_47#_c_204_n 0.0218847f $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_133 B N_A_27_47#_c_204_n 0.0936703f $X=3.23 $Y=1.105 $X2=0 $Y2=0
cc_134 N_B_c_154_n N_A_27_47#_c_205_n 2.24692e-19 $X=3.02 $Y=1.16 $X2=0 $Y2=0
cc_135 B N_A_27_47#_c_205_n 0.0123975f $X=3.23 $Y=1.105 $X2=0 $Y2=0
cc_136 N_B_c_154_n N_A_27_47#_c_200_n 0.0139634f $X=3.02 $Y=1.16 $X2=0 $Y2=0
cc_137 B N_A_27_47#_c_200_n 0.00240847f $X=3.23 $Y=1.105 $X2=0 $Y2=0
cc_138 N_B_c_156_n N_VPWR_c_284_n 0.00381622f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_139 N_B_c_157_n N_VPWR_c_285_n 0.0059385f $X=2.5 $Y=1.41 $X2=0 $Y2=0
cc_140 N_B_c_156_n N_VPWR_c_291_n 0.0048852f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_141 N_B_c_157_n N_VPWR_c_291_n 0.00673617f $X=2.5 $Y=1.41 $X2=0 $Y2=0
cc_142 N_B_c_156_n N_VPWR_c_282_n 0.00653068f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_143 N_B_c_157_n N_VPWR_c_282_n 0.00818986f $X=2.5 $Y=1.41 $X2=0 $Y2=0
cc_144 N_B_c_156_n N_Y_c_366_n 0.009108f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_145 N_B_c_157_n N_Y_c_362_n 0.0122434f $X=2.5 $Y=1.41 $X2=0 $Y2=0
cc_146 N_B_c_156_n N_Y_c_365_n 5.16456e-19 $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_147 N_B_c_156_n N_Y_c_369_n 0.010999f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_148 N_B_c_157_n N_Y_c_369_n 0.0143512f $X=2.5 $Y=1.41 $X2=0 $Y2=0
cc_149 N_B_M1004_g N_VGND_c_436_n 0.00195249f $X=2.625 $Y=0.56 $X2=0 $Y2=0
cc_150 N_B_M1004_g N_VGND_c_439_n 0.00357877f $X=2.625 $Y=0.56 $X2=0 $Y2=0
cc_151 N_B_M1005_g N_VGND_c_439_n 0.00357877f $X=3.095 $Y=0.56 $X2=0 $Y2=0
cc_152 N_B_M1004_g N_VGND_c_440_n 0.00668309f $X=2.625 $Y=0.56 $X2=0 $Y2=0
cc_153 N_B_M1005_g N_VGND_c_440_n 0.00538422f $X=3.095 $Y=0.56 $X2=0 $Y2=0
cc_154 N_B_M1004_g N_A_228_47#_c_493_n 0.0143183f $X=2.625 $Y=0.56 $X2=0 $Y2=0
cc_155 N_B_c_154_n N_A_228_47#_c_493_n 0.00323379f $X=3.02 $Y=1.16 $X2=0 $Y2=0
cc_156 N_B_c_153_n N_A_228_47#_c_494_n 0.0168924f $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_157 B N_A_228_47#_c_494_n 0.063036f $X=3.23 $Y=1.105 $X2=0 $Y2=0
cc_158 N_B_M1004_g N_A_448_47#_c_522_n 0.00903374f $X=2.625 $Y=0.56 $X2=0 $Y2=0
cc_159 N_B_M1005_g N_A_448_47#_c_522_n 0.0111176f $X=3.095 $Y=0.56 $X2=0 $Y2=0
cc_160 B N_A_448_47#_c_522_n 0.00464179f $X=3.23 $Y=1.105 $X2=0 $Y2=0
cc_161 B N_A_448_47#_c_523_n 0.0142952f $X=3.23 $Y=1.105 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_204_n N_VPWR_M1002_d 0.0035219f $X=3.67 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_163 N_A_27_47#_c_204_n N_VPWR_M1011_d 0.00179023f $X=3.67 $Y=1.53 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_204_n N_VPWR_M1012_s 0.00286974f $X=3.67 $Y=1.53 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_204_n N_VPWR_M1008_d 0.00286974f $X=3.67 $Y=1.53 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_204_n N_VPWR_c_283_n 0.0208167f $X=3.67 $Y=1.53 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_208_n N_VPWR_c_283_n 0.0105094f $X=0.25 $Y=2.065 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_201_n N_VPWR_c_286_n 0.00581355f $X=3.54 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_202_n N_VPWR_c_288_n 0.00639018f $X=4.01 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_201_n N_VPWR_c_295_n 0.00597712f $X=3.54 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_202_n N_VPWR_c_295_n 0.00523784f $X=4.01 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_207_n N_VPWR_c_296_n 0.0201557f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_173 N_A_27_47#_M1002_s N_VPWR_c_282_n 0.00217517f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_c_201_n N_VPWR_c_282_n 0.00787843f $X=3.54 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_27_47#_c_202_n N_VPWR_c_282_n 0.00787547f $X=4.01 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A_27_47#_c_207_n N_VPWR_c_282_n 0.0120807f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_177 N_A_27_47#_c_204_n N_Y_M1006_s 0.00187091f $X=3.67 $Y=1.53 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_204_n N_Y_M1003_d 0.00187091f $X=3.67 $Y=1.53 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_204_n N_Y_M1008_s 0.00190105f $X=3.67 $Y=1.53 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_204_n N_Y_c_366_n 0.0316355f $X=3.67 $Y=1.53 $X2=0 $Y2=0
cc_181 N_A_27_47#_c_201_n N_Y_c_362_n 0.00967226f $X=3.54 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A_27_47#_c_204_n N_Y_c_362_n 0.0732708f $X=3.67 $Y=1.53 $X2=0 $Y2=0
cc_183 N_A_27_47#_M1001_g N_Y_c_360_n 0.00426831f $X=3.515 $Y=0.56 $X2=0 $Y2=0
cc_184 N_A_27_47#_M1010_g N_Y_c_360_n 0.0174772f $X=4.035 $Y=0.56 $X2=0 $Y2=0
cc_185 N_A_27_47#_c_204_n N_Y_c_360_n 0.00344548f $X=3.67 $Y=1.53 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_205_n N_Y_c_360_n 0.0264832f $X=3.835 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_27_47#_c_200_n N_Y_c_360_n 0.00438594f $X=4.01 $Y=1.217 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_202_n N_Y_c_363_n 0.0184579f $X=4.01 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A_27_47#_c_204_n N_Y_c_363_n 0.00614204f $X=3.67 $Y=1.53 $X2=0 $Y2=0
cc_190 N_A_27_47#_c_204_n N_Y_c_365_n 0.0211749f $X=3.67 $Y=1.53 $X2=0 $Y2=0
cc_191 N_A_27_47#_c_204_n N_Y_c_369_n 0.0211749f $X=3.67 $Y=1.53 $X2=0 $Y2=0
cc_192 N_A_27_47#_c_201_n N_Y_c_390_n 0.0173634f $X=3.54 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_204_n N_Y_c_390_n 0.020626f $X=3.67 $Y=1.53 $X2=0 $Y2=0
cc_194 N_A_27_47#_c_200_n N_Y_c_390_n 7.26953e-19 $X=4.01 $Y=1.217 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_202_n Y 0.0106918f $X=4.01 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A_27_47#_M1010_g Y 0.0153288f $X=4.035 $Y=0.56 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_204_n Y 0.0102207f $X=3.67 $Y=1.53 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_205_n Y 0.0213532f $X=3.835 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A_27_47#_c_198_n N_VGND_c_435_n 0.0114533f $X=0.175 $Y=1.445 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_204_n N_VGND_c_435_n 0.00412107f $X=3.67 $Y=1.53 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_199_n N_VGND_c_435_n 0.0252887f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_202 N_A_27_47#_M1001_g N_VGND_c_439_n 0.00357877f $X=3.515 $Y=0.56 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_M1010_g N_VGND_c_439_n 0.00357877f $X=4.035 $Y=0.56 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_M1013_s N_VGND_c_440_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_M1001_g N_VGND_c_440_n 0.005504f $X=3.515 $Y=0.56 $X2=0 $Y2=0
cc_206 N_A_27_47#_M1010_g N_VGND_c_440_n 0.00651046f $X=4.035 $Y=0.56 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_199_n N_VGND_c_440_n 0.012035f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_208 N_A_27_47#_c_199_n N_VGND_c_441_n 0.0201353f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_209 N_A_27_47#_c_204_n N_A_228_47#_c_494_n 0.00813711f $X=3.67 $Y=1.53 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_M1001_g N_A_448_47#_c_524_n 0.0131041f $X=3.515 $Y=0.56 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_M1010_g N_A_448_47#_c_524_n 0.00935436f $X=4.035 $Y=0.56 $X2=0
+ $Y2=0
cc_212 N_VPWR_c_282_n N_Y_M1006_s 0.00231261f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_213 N_VPWR_c_282_n N_Y_M1003_d 0.00231261f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_214 N_VPWR_c_282_n N_Y_M1008_s 0.00258911f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_215 N_VPWR_M1011_d N_Y_c_366_n 0.00364456f $X=1.65 $Y=1.485 $X2=0 $Y2=0
cc_216 N_VPWR_c_284_n N_Y_c_366_n 0.0133389f $X=1.795 $Y=2.34 $X2=0 $Y2=0
cc_217 N_VPWR_c_289_n N_Y_c_366_n 0.00271054f $X=1.71 $Y=2.72 $X2=0 $Y2=0
cc_218 N_VPWR_c_291_n N_Y_c_366_n 0.00201496f $X=2.65 $Y=2.72 $X2=0 $Y2=0
cc_219 N_VPWR_c_282_n N_Y_c_366_n 0.00979995f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_220 N_VPWR_M1012_s N_Y_c_362_n 0.00527719f $X=2.59 $Y=1.485 $X2=0 $Y2=0
cc_221 N_VPWR_M1008_d N_Y_c_362_n 0.00553617f $X=3.18 $Y=1.485 $X2=0 $Y2=0
cc_222 N_VPWR_c_285_n N_Y_c_362_n 0.0157895f $X=2.735 $Y=2.34 $X2=0 $Y2=0
cc_223 N_VPWR_c_286_n N_Y_c_362_n 0.0191028f $X=3.305 $Y=2.34 $X2=0 $Y2=0
cc_224 N_VPWR_c_282_n N_Y_c_362_n 0.0215419f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_225 N_VPWR_M1009_d N_Y_c_363_n 0.00691947f $X=4.1 $Y=1.485 $X2=0 $Y2=0
cc_226 N_VPWR_c_287_n N_Y_c_363_n 6.86176e-19 $X=4.305 $Y=2.635 $X2=0 $Y2=0
cc_227 N_VPWR_c_288_n N_Y_c_363_n 0.0244211f $X=4.245 $Y=2.34 $X2=0 $Y2=0
cc_228 N_VPWR_c_295_n N_Y_c_363_n 0.00346609f $X=4.16 $Y=2.72 $X2=0 $Y2=0
cc_229 N_VPWR_c_282_n N_Y_c_363_n 0.00949941f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_230 N_VPWR_c_283_n N_Y_c_365_n 0.0498192f $X=0.795 $Y=2 $X2=0 $Y2=0
cc_231 N_VPWR_c_284_n N_Y_c_365_n 0.0177504f $X=1.795 $Y=2.34 $X2=0 $Y2=0
cc_232 N_VPWR_c_289_n N_Y_c_365_n 0.0223557f $X=1.71 $Y=2.72 $X2=0 $Y2=0
cc_233 N_VPWR_c_282_n N_Y_c_365_n 0.0140101f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_234 N_VPWR_c_284_n N_Y_c_369_n 0.02165f $X=1.795 $Y=2.34 $X2=0 $Y2=0
cc_235 N_VPWR_c_285_n N_Y_c_369_n 0.0182679f $X=2.735 $Y=2.34 $X2=0 $Y2=0
cc_236 N_VPWR_c_291_n N_Y_c_369_n 0.0223557f $X=2.65 $Y=2.72 $X2=0 $Y2=0
cc_237 N_VPWR_c_282_n N_Y_c_369_n 0.0140101f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_238 N_VPWR_c_286_n N_Y_c_390_n 0.0221891f $X=3.305 $Y=2.34 $X2=0 $Y2=0
cc_239 N_VPWR_c_288_n N_Y_c_390_n 0.0150554f $X=4.245 $Y=2.34 $X2=0 $Y2=0
cc_240 N_VPWR_c_295_n N_Y_c_390_n 0.0187893f $X=4.16 $Y=2.72 $X2=0 $Y2=0
cc_241 N_VPWR_c_282_n N_Y_c_390_n 0.0110885f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_242 N_VPWR_M1009_d Y 0.0049632f $X=4.1 $Y=1.485 $X2=0 $Y2=0
cc_243 N_Y_c_360_n N_VGND_c_439_n 8.12174e-19 $X=4.25 $Y=0.77 $X2=0 $Y2=0
cc_244 N_Y_M1001_d N_VGND_c_440_n 0.00297142f $X=3.59 $Y=0.235 $X2=0 $Y2=0
cc_245 N_Y_c_360_n N_VGND_c_440_n 0.00171309f $X=4.25 $Y=0.77 $X2=0 $Y2=0
cc_246 N_Y_c_360_n N_A_448_47#_M1010_s 0.00324009f $X=4.25 $Y=0.77 $X2=0 $Y2=0
cc_247 N_Y_c_360_n N_A_448_47#_c_523_n 0.0119693f $X=4.25 $Y=0.77 $X2=0 $Y2=0
cc_248 N_Y_M1001_d N_A_448_47#_c_524_n 0.00508685f $X=3.59 $Y=0.235 $X2=0 $Y2=0
cc_249 N_Y_c_360_n N_A_448_47#_c_524_n 0.0524427f $X=4.25 $Y=0.77 $X2=0 $Y2=0
cc_250 N_VGND_c_440_n N_A_228_47#_M1000_s 0.0030386f $X=4.37 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_251 N_VGND_c_440_n N_A_228_47#_M1004_s 0.00256987f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_252 N_VGND_c_437_n N_A_228_47#_c_495_n 0.0231806f $X=1.71 $Y=0 $X2=0 $Y2=0
cc_253 N_VGND_c_440_n N_A_228_47#_c_495_n 0.0143352f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_254 N_VGND_c_435_n N_A_228_47#_c_491_n 0.00878993f $X=0.795 $Y=0.38 $X2=0
+ $Y2=0
cc_255 N_VGND_M1007_d N_A_228_47#_c_494_n 0.00285834f $X=1.66 $Y=0.235 $X2=0
+ $Y2=0
cc_256 N_VGND_c_436_n N_A_228_47#_c_494_n 0.0191473f $X=1.795 $Y=0.38 $X2=0
+ $Y2=0
cc_257 N_VGND_c_437_n N_A_228_47#_c_494_n 0.00260993f $X=1.71 $Y=0 $X2=0 $Y2=0
cc_258 N_VGND_c_439_n N_A_228_47#_c_494_n 0.00374451f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_259 N_VGND_c_440_n N_A_228_47#_c_494_n 0.0124612f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_260 N_VGND_c_440_n N_A_448_47#_M1004_d 0.00250339f $X=4.37 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_261 N_VGND_c_440_n N_A_448_47#_M1005_d 0.0021521f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_262 N_VGND_c_440_n N_A_448_47#_M1010_s 0.00209344f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_263 N_VGND_c_436_n N_A_448_47#_c_522_n 0.0141662f $X=1.795 $Y=0.38 $X2=0
+ $Y2=0
cc_264 N_VGND_c_439_n N_A_448_47#_c_522_n 0.0585829f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_265 N_VGND_c_440_n N_A_448_47#_c_522_n 0.0366524f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_266 N_VGND_c_439_n N_A_448_47#_c_524_n 0.061198f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_267 N_VGND_c_440_n N_A_448_47#_c_524_n 0.038149f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_268 N_VGND_c_439_n N_A_448_47#_c_543_n 0.0114305f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_269 N_VGND_c_440_n N_A_448_47#_c_543_n 0.00653933f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_270 N_A_228_47#_c_492_n N_A_448_47#_M1004_d 0.00229711f $X=2.335 $Y=0.77
+ $X2=-0.19 $Y2=-0.24
cc_271 N_A_228_47#_c_493_n N_A_448_47#_M1004_d 0.00210106f $X=2.835 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_272 N_A_228_47#_M1004_s N_A_448_47#_c_522_n 0.00401386f $X=2.7 $Y=0.235 $X2=0
+ $Y2=0
cc_273 N_A_228_47#_c_492_n N_A_448_47#_c_522_n 0.0463045f $X=2.335 $Y=0.77 $X2=0
+ $Y2=0
cc_274 N_A_228_47#_c_493_n N_A_448_47#_c_523_n 0.00126647f $X=2.835 $Y=0.72
+ $X2=0 $Y2=0
