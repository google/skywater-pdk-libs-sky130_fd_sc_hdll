* File: sky130_fd_sc_hdll__o211a_4.pxi.spice
* Created: Thu Aug 27 19:18:24 2020
* 
x_PM_SKY130_FD_SC_HDLL__O211A_4%A_80_21# N_A_80_21#_M1023_d N_A_80_21#_M1001_d
+ N_A_80_21#_M1014_s N_A_80_21#_M1006_s N_A_80_21#_c_96_n N_A_80_21#_M1009_g
+ N_A_80_21#_c_105_n N_A_80_21#_M1005_g N_A_80_21#_c_97_n N_A_80_21#_M1013_g
+ N_A_80_21#_c_106_n N_A_80_21#_M1010_g N_A_80_21#_c_98_n N_A_80_21#_M1021_g
+ N_A_80_21#_c_99_n N_A_80_21#_M1022_g N_A_80_21#_c_107_n N_A_80_21#_M1012_g
+ N_A_80_21#_c_108_n N_A_80_21#_M1017_g N_A_80_21#_c_204_p N_A_80_21#_c_100_n
+ N_A_80_21#_c_101_n N_A_80_21#_c_102_n N_A_80_21#_c_103_n N_A_80_21#_c_115_p
+ N_A_80_21#_c_116_p N_A_80_21#_c_160_p N_A_80_21#_c_141_p N_A_80_21#_c_136_p
+ N_A_80_21#_c_120_p N_A_80_21#_c_121_p N_A_80_21#_c_104_n N_A_80_21#_c_132_p
+ N_A_80_21#_c_122_p N_A_80_21#_c_149_p PM_SKY130_FD_SC_HDLL__O211A_4%A_80_21#
x_PM_SKY130_FD_SC_HDLL__O211A_4%B1 N_B1_c_257_n N_B1_M1001_g N_B1_c_258_n
+ N_B1_M1008_g N_B1_c_259_n N_B1_M1015_g N_B1_c_260_n N_B1_M1002_g N_B1_c_261_n
+ N_B1_c_285_n B1 N_B1_c_262_n PM_SKY130_FD_SC_HDLL__O211A_4%B1
x_PM_SKY130_FD_SC_HDLL__O211A_4%C1 N_C1_c_341_n N_C1_M1023_g N_C1_c_345_n
+ N_C1_M1004_g N_C1_c_346_n N_C1_M1014_g N_C1_c_342_n N_C1_M1019_g C1
+ N_C1_c_343_n N_C1_c_344_n C1 PM_SKY130_FD_SC_HDLL__O211A_4%C1
x_PM_SKY130_FD_SC_HDLL__O211A_4%A1 N_A1_c_388_n N_A1_M1007_g N_A1_c_389_n
+ N_A1_M1018_g N_A1_c_390_n N_A1_M1016_g N_A1_c_391_n N_A1_M1011_g N_A1_c_392_n
+ N_A1_c_402_n N_A1_c_405_n A1 N_A1_c_393_n PM_SKY130_FD_SC_HDLL__O211A_4%A1
x_PM_SKY130_FD_SC_HDLL__O211A_4%A2 N_A2_c_461_n N_A2_M1000_g N_A2_c_465_n
+ N_A2_M1006_g N_A2_c_462_n N_A2_M1003_g N_A2_c_466_n N_A2_M1020_g A2
+ N_A2_c_463_n N_A2_c_464_n A2 PM_SKY130_FD_SC_HDLL__O211A_4%A2
x_PM_SKY130_FD_SC_HDLL__O211A_4%VPWR N_VPWR_M1005_d N_VPWR_M1010_d
+ N_VPWR_M1017_d N_VPWR_M1004_d N_VPWR_M1002_s N_VPWR_M1011_d N_VPWR_c_515_n
+ N_VPWR_c_516_n N_VPWR_c_517_n N_VPWR_c_518_n N_VPWR_c_519_n N_VPWR_c_520_n
+ N_VPWR_c_521_n N_VPWR_c_522_n N_VPWR_c_523_n VPWR N_VPWR_c_524_n
+ N_VPWR_c_525_n N_VPWR_c_526_n N_VPWR_c_527_n N_VPWR_c_528_n N_VPWR_c_529_n
+ N_VPWR_c_530_n N_VPWR_c_531_n N_VPWR_c_532_n N_VPWR_c_514_n
+ PM_SKY130_FD_SC_HDLL__O211A_4%VPWR
x_PM_SKY130_FD_SC_HDLL__O211A_4%X N_X_M1009_d N_X_M1021_d N_X_M1005_s
+ N_X_M1012_s N_X_c_629_n N_X_c_624_n N_X_c_625_n N_X_c_674_p N_X_c_634_n
+ N_X_c_638_n N_X_c_626_n N_X_c_677_p N_X_c_645_n N_X_c_648_n N_X_c_627_n X
+ N_X_c_622_n X PM_SKY130_FD_SC_HDLL__O211A_4%X
x_PM_SKY130_FD_SC_HDLL__O211A_4%VGND N_VGND_M1009_s N_VGND_M1013_s
+ N_VGND_M1022_s N_VGND_M1007_s N_VGND_M1003_s N_VGND_c_697_n N_VGND_c_698_n
+ N_VGND_c_699_n N_VGND_c_700_n N_VGND_c_701_n N_VGND_c_702_n N_VGND_c_703_n
+ N_VGND_c_704_n N_VGND_c_705_n VGND N_VGND_c_706_n N_VGND_c_707_n
+ N_VGND_c_708_n N_VGND_c_709_n N_VGND_c_710_n
+ PM_SKY130_FD_SC_HDLL__O211A_4%VGND
x_PM_SKY130_FD_SC_HDLL__O211A_4%A_524_47# N_A_524_47#_M1008_s
+ N_A_524_47#_M1015_s N_A_524_47#_M1000_d N_A_524_47#_M1016_d
+ N_A_524_47#_c_797_n N_A_524_47#_c_815_n N_A_524_47#_c_804_n
+ N_A_524_47#_c_817_n N_A_524_47#_c_805_n N_A_524_47#_c_821_n
+ N_A_524_47#_c_798_n N_A_524_47#_c_799_n N_A_524_47#_c_837_n
+ PM_SKY130_FD_SC_HDLL__O211A_4%A_524_47#
cc_1 VNB N_A_80_21#_c_96_n 0.0187769f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_2 VNB N_A_80_21#_c_97_n 0.0169667f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=0.995
cc_3 VNB N_A_80_21#_c_98_n 0.0167707f $X=-0.19 $Y=-0.24 $X2=1.415 $Y2=0.995
cc_4 VNB N_A_80_21#_c_99_n 0.0193579f $X=-0.19 $Y=-0.24 $X2=1.885 $Y2=0.995
cc_5 VNB N_A_80_21#_c_100_n 0.107986f $X=-0.19 $Y=-0.24 $X2=2.26 $Y2=1.16
cc_6 VNB N_A_80_21#_c_101_n 0.00456197f $X=-0.19 $Y=-0.24 $X2=2.51 $Y2=1.065
cc_7 VNB N_A_80_21#_c_102_n 2.30681e-19 $X=-0.19 $Y=-0.24 $X2=2.51 $Y2=1.855
cc_8 VNB N_A_80_21#_c_103_n 0.00634842f $X=-0.19 $Y=-0.24 $X2=2.62 $Y2=0.725
cc_9 VNB N_A_80_21#_c_104_n 0.00120371f $X=-0.19 $Y=-0.24 $X2=2.51 $Y2=1.165
cc_10 VNB N_B1_c_257_n 0.0225703f $X=-0.19 $Y=-0.24 $X2=3.395 $Y2=0.235
cc_11 VNB N_B1_c_258_n 0.0190789f $X=-0.19 $Y=-0.24 $X2=5.53 $Y2=1.485
cc_12 VNB N_B1_c_259_n 0.0166507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_B1_c_260_n 0.0198564f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_B1_c_261_n 0.00353893f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.56
cc_15 VNB N_B1_c_262_n 0.00421326f $X=-0.19 $Y=-0.24 $X2=1.415 $Y2=0.56
cc_16 VNB N_C1_c_341_n 0.0178645f $X=-0.19 $Y=-0.24 $X2=3.395 $Y2=0.235
cc_17 VNB N_C1_c_342_n 0.0181228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_C1_c_343_n 0.00151558f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=0.995
cc_19 VNB N_C1_c_344_n 0.0460125f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=0.56
cc_20 VNB N_A1_c_388_n 0.0180289f $X=-0.19 $Y=-0.24 $X2=3.395 $Y2=0.235
cc_21 VNB N_A1_c_389_n 0.0239403f $X=-0.19 $Y=-0.24 $X2=5.53 $Y2=1.485
cc_22 VNB N_A1_c_390_n 0.0227688f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A1_c_391_n 0.0369999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A1_c_392_n 0.00191122f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.56
cc_25 VNB N_A1_c_393_n 0.0115052f $X=-0.19 $Y=-0.24 $X2=1.415 $Y2=0.995
cc_26 VNB N_A2_c_461_n 0.0178602f $X=-0.19 $Y=-0.24 $X2=3.395 $Y2=0.235
cc_27 VNB N_A2_c_462_n 0.0173683f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A2_c_463_n 0.038012f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.985
cc_29 VNB N_A2_c_464_n 0.00366605f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=0.995
cc_30 VNB N_VPWR_c_514_n 0.288713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_X_c_622_n 0.0076991f $X=-0.19 $Y=-0.24 $X2=2.26 $Y2=1.16
cc_32 VNB X 0.0253296f $X=-0.19 $Y=-0.24 $X2=2.51 $Y2=0.815
cc_33 VNB N_VGND_c_697_n 0.010288f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.41
cc_34 VNB N_VGND_c_698_n 0.011915f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.985
cc_35 VNB N_VGND_c_699_n 0.00214953f $X=-0.19 $Y=-0.24 $X2=1.42 $Y2=1.41
cc_36 VNB N_VGND_c_700_n 0.00546668f $X=-0.19 $Y=-0.24 $X2=1.415 $Y2=0.56
cc_37 VNB N_VGND_c_701_n 0.00479809f $X=-0.19 $Y=-0.24 $X2=1.885 $Y2=0.56
cc_38 VNB N_VGND_c_702_n 0.0609626f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=1.985
cc_39 VNB N_VGND_c_703_n 0.00602438f $X=-0.19 $Y=-0.24 $X2=2.38 $Y2=1.41
cc_40 VNB N_VGND_c_704_n 0.0190856f $X=-0.19 $Y=-0.24 $X2=2.38 $Y2=1.985
cc_41 VNB N_VGND_c_705_n 0.00362328f $X=-0.19 $Y=-0.24 $X2=2.4 $Y2=1.165
cc_42 VNB N_VGND_c_706_n 0.0147094f $X=-0.19 $Y=-0.24 $X2=0.75 $Y2=1.16
cc_43 VNB N_VGND_c_707_n 0.0258086f $X=-0.19 $Y=-0.24 $X2=2.51 $Y2=0.815
cc_44 VNB N_VGND_c_708_n 0.0183091f $X=-0.19 $Y=-0.24 $X2=4.25 $Y2=2.025
cc_45 VNB N_VGND_c_709_n 0.33776f $X=-0.19 $Y=-0.24 $X2=4.25 $Y2=2.3
cc_46 VNB N_VGND_c_710_n 0.00510002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_524_47#_c_797_n 0.00276851f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_48 VNB N_A_524_47#_c_798_n 0.00752521f $X=-0.19 $Y=-0.24 $X2=1.415 $Y2=0.995
cc_49 VNB N_A_524_47#_c_799_n 0.0175626f $X=-0.19 $Y=-0.24 $X2=1.885 $Y2=0.56
cc_50 VPB N_A_80_21#_c_105_n 0.0186521f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.41
cc_51 VPB N_A_80_21#_c_106_n 0.0155203f $X=-0.19 $Y=1.305 $X2=1.42 $Y2=1.41
cc_52 VPB N_A_80_21#_c_107_n 0.0158533f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=1.41
cc_53 VPB N_A_80_21#_c_108_n 0.0155987f $X=-0.19 $Y=1.305 $X2=2.38 $Y2=1.41
cc_54 VPB N_A_80_21#_c_100_n 0.0596483f $X=-0.19 $Y=1.305 $X2=2.26 $Y2=1.16
cc_55 VPB N_A_80_21#_c_102_n 0.00107122f $X=-0.19 $Y=1.305 $X2=2.51 $Y2=1.855
cc_56 VPB N_B1_c_257_n 0.0267566f $X=-0.19 $Y=1.305 $X2=3.395 $Y2=0.235
cc_57 VPB N_B1_c_260_n 0.0240364f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_B1_c_261_n 0.00159688f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_59 VPB B1 0.0122338f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=0.995
cc_60 VPB N_B1_c_262_n 0.00242379f $X=-0.19 $Y=1.305 $X2=1.415 $Y2=0.56
cc_61 VPB N_C1_c_345_n 0.0168366f $X=-0.19 $Y=1.305 $X2=5.53 $Y2=1.485
cc_62 VPB N_C1_c_346_n 0.0161061f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_C1_c_344_n 0.0247051f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=0.56
cc_64 VPB N_A1_c_389_n 0.0255352f $X=-0.19 $Y=1.305 $X2=5.53 $Y2=1.485
cc_65 VPB N_A1_c_391_n 0.0337389f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A1_c_392_n 0.00290466f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_67 VPB N_A1_c_393_n 0.0169895f $X=-0.19 $Y=1.305 $X2=1.415 $Y2=0.995
cc_68 VPB N_A2_c_465_n 0.0165852f $X=-0.19 $Y=1.305 $X2=5.53 $Y2=1.485
cc_69 VPB N_A2_c_466_n 0.0165913f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A2_c_463_n 0.0215172f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.985
cc_71 VPB N_A2_c_464_n 4.74361e-19 $X=-0.19 $Y=1.305 $X2=0.945 $Y2=0.995
cc_72 VPB N_VPWR_c_515_n 0.0274981f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=0.56
cc_73 VPB N_VPWR_c_516_n 3.26289e-19 $X=-0.19 $Y=1.305 $X2=1.415 $Y2=0.995
cc_74 VPB N_VPWR_c_517_n 4.07994e-19 $X=-0.19 $Y=1.305 $X2=1.885 $Y2=0.56
cc_75 VPB N_VPWR_c_518_n 4.89699e-19 $X=-0.19 $Y=1.305 $X2=1.9 $Y2=1.985
cc_76 VPB N_VPWR_c_519_n 0.00524989f $X=-0.19 $Y=1.305 $X2=2.4 $Y2=1.165
cc_77 VPB N_VPWR_c_520_n 0.0110648f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_78 VPB N_VPWR_c_521_n 0.0256219f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_522_n 0.0169255f $X=-0.19 $Y=1.305 $X2=2.26 $Y2=1.16
cc_80 VPB N_VPWR_c_523_n 0.00503031f $X=-0.19 $Y=1.305 $X2=2.51 $Y2=0.815
cc_81 VPB N_VPWR_c_524_n 0.0174178f $X=-0.19 $Y=1.305 $X2=2.51 $Y2=1.855
cc_82 VPB N_VPWR_c_525_n 0.014625f $X=-0.19 $Y=1.305 $X2=3 $Y2=1.94
cc_83 VPB N_VPWR_c_526_n 0.0145309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_527_n 0.0159194f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_528_n 0.0424952f $X=-0.19 $Y=1.305 $X2=4.25 $Y2=1.94
cc_86 VPB N_VPWR_c_529_n 0.00615892f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=1.202
cc_87 VPB N_VPWR_c_530_n 0.00503453f $X=-0.19 $Y=1.305 $X2=1.885 $Y2=1.202
cc_88 VPB N_VPWR_c_531_n 0.00502999f $X=-0.19 $Y=1.305 $X2=2.38 $Y2=1.202
cc_89 VPB N_VPWR_c_532_n 0.00502957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_514_n 0.0596295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_X_c_624_n 0.0100031f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_92 VPB N_X_c_625_n 0.0248561f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.41
cc_93 VPB N_X_c_626_n 0.00398104f $X=-0.19 $Y=1.305 $X2=1.415 $Y2=0.56
cc_94 VPB N_X_c_627_n 0.00107973f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.16
cc_95 VPB X 0.00764395f $X=-0.19 $Y=1.305 $X2=2.51 $Y2=0.815
cc_96 N_A_80_21#_c_108_n N_B1_c_257_n 0.0337282f $X=2.38 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_97 N_A_80_21#_c_100_n N_B1_c_257_n 0.0190762f $X=2.26 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_98 N_A_80_21#_c_101_n N_B1_c_257_n 4.59577e-19 $X=2.51 $Y=1.065 $X2=-0.19
+ $Y2=-0.24
cc_99 N_A_80_21#_c_102_n N_B1_c_257_n 0.00649141f $X=2.51 $Y=1.855 $X2=-0.19
+ $Y2=-0.24
cc_100 N_A_80_21#_c_115_p N_B1_c_257_n 0.00253744f $X=3.605 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_101 N_A_80_21#_c_116_p N_B1_c_257_n 0.0152274f $X=3 $Y=1.94 $X2=-0.19
+ $Y2=-0.24
cc_102 N_A_80_21#_c_104_n N_B1_c_257_n 0.00148116f $X=2.51 $Y=1.165 $X2=-0.19
+ $Y2=-0.24
cc_103 N_A_80_21#_c_101_n N_B1_c_258_n 0.00570677f $X=2.51 $Y=1.065 $X2=0 $Y2=0
cc_104 N_A_80_21#_c_115_p N_B1_c_258_n 0.0122418f $X=3.605 $Y=0.73 $X2=0 $Y2=0
cc_105 N_A_80_21#_c_120_p N_B1_c_260_n 0.0071253f $X=4.25 $Y=2.3 $X2=0 $Y2=0
cc_106 N_A_80_21#_c_121_p N_B1_c_260_n 0.0106439f $X=5.465 $Y=1.94 $X2=0 $Y2=0
cc_107 N_A_80_21#_c_122_p N_B1_c_260_n 0.00302271f $X=4.25 $Y=1.94 $X2=0 $Y2=0
cc_108 N_A_80_21#_c_100_n N_B1_c_261_n 3.86288e-19 $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_80_21#_c_101_n N_B1_c_261_n 0.00528199f $X=2.51 $Y=1.065 $X2=0 $Y2=0
cc_110 N_A_80_21#_c_102_n N_B1_c_261_n 0.0135702f $X=2.51 $Y=1.855 $X2=0 $Y2=0
cc_111 N_A_80_21#_c_115_p N_B1_c_261_n 0.0182618f $X=3.605 $Y=0.73 $X2=0 $Y2=0
cc_112 N_A_80_21#_c_104_n N_B1_c_261_n 0.0167371f $X=2.51 $Y=1.165 $X2=0 $Y2=0
cc_113 N_A_80_21#_M1001_d N_B1_c_285_n 9.07836e-19 $X=2.945 $Y=1.485 $X2=0 $Y2=0
cc_114 N_A_80_21#_c_108_n N_B1_c_285_n 2.29829e-19 $X=2.38 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A_80_21#_c_102_n N_B1_c_285_n 0.0192641f $X=2.51 $Y=1.855 $X2=0 $Y2=0
cc_116 N_A_80_21#_c_116_p N_B1_c_285_n 0.0117795f $X=3 $Y=1.94 $X2=0 $Y2=0
cc_117 N_A_80_21#_c_132_p N_B1_c_285_n 0.00743164f $X=3.18 $Y=1.94 $X2=0 $Y2=0
cc_118 N_A_80_21#_M1001_d B1 0.0040638f $X=2.945 $Y=1.485 $X2=0 $Y2=0
cc_119 N_A_80_21#_M1014_s B1 0.0021586f $X=4.08 $Y=1.485 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_115_p B1 0.00412163f $X=3.605 $Y=0.73 $X2=0 $Y2=0
cc_121 N_A_80_21#_c_136_p B1 0.0390477f $X=4.085 $Y=1.94 $X2=0 $Y2=0
cc_122 N_A_80_21#_c_121_p B1 0.0121079f $X=5.465 $Y=1.94 $X2=0 $Y2=0
cc_123 N_A_80_21#_c_132_p B1 0.0226705f $X=3.18 $Y=1.94 $X2=0 $Y2=0
cc_124 N_A_80_21#_c_122_p B1 0.01868f $X=4.25 $Y=1.94 $X2=0 $Y2=0
cc_125 N_A_80_21#_c_115_p N_C1_c_341_n 0.011593f $X=3.605 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_126 N_A_80_21#_c_141_p N_C1_c_345_n 0.00782047f $X=3.195 $Y=2.3 $X2=0 $Y2=0
cc_127 N_A_80_21#_c_136_p N_C1_c_345_n 0.0140035f $X=4.085 $Y=1.94 $X2=0 $Y2=0
cc_128 N_A_80_21#_c_136_p N_C1_c_346_n 0.013845f $X=4.085 $Y=1.94 $X2=0 $Y2=0
cc_129 N_A_80_21#_c_115_p N_C1_c_342_n 0.00305762f $X=3.605 $Y=0.73 $X2=0 $Y2=0
cc_130 N_A_80_21#_c_115_p N_C1_c_343_n 0.0314639f $X=3.605 $Y=0.73 $X2=0 $Y2=0
cc_131 N_A_80_21#_c_115_p N_C1_c_344_n 0.0080867f $X=3.605 $Y=0.73 $X2=0 $Y2=0
cc_132 N_A_80_21#_c_120_p N_A1_c_389_n 7.91317e-19 $X=4.25 $Y=2.3 $X2=0 $Y2=0
cc_133 N_A_80_21#_c_121_p N_A1_c_389_n 0.0146234f $X=5.465 $Y=1.94 $X2=0 $Y2=0
cc_134 N_A_80_21#_c_149_p N_A1_c_389_n 0.00171453f $X=5.68 $Y=2.02 $X2=0 $Y2=0
cc_135 N_A_80_21#_c_149_p N_A1_c_391_n 0.00185764f $X=5.68 $Y=2.02 $X2=0 $Y2=0
cc_136 N_A_80_21#_M1006_s N_A1_c_402_n 0.00354602f $X=5.53 $Y=1.485 $X2=0 $Y2=0
cc_137 N_A_80_21#_c_121_p N_A1_c_402_n 0.0178989f $X=5.465 $Y=1.94 $X2=0 $Y2=0
cc_138 N_A_80_21#_c_149_p N_A1_c_402_n 0.0211177f $X=5.68 $Y=2.02 $X2=0 $Y2=0
cc_139 N_A_80_21#_c_121_p N_A1_c_405_n 0.0175059f $X=5.465 $Y=1.94 $X2=0 $Y2=0
cc_140 N_A_80_21#_c_121_p N_A2_c_465_n 0.00824561f $X=5.465 $Y=1.94 $X2=0 $Y2=0
cc_141 N_A_80_21#_c_149_p N_A2_c_465_n 0.0122625f $X=5.68 $Y=2.02 $X2=0 $Y2=0
cc_142 N_A_80_21#_c_149_p N_A2_c_466_n 0.0116285f $X=5.68 $Y=2.02 $X2=0 $Y2=0
cc_143 N_A_80_21#_c_102_n N_VPWR_M1017_d 0.00366084f $X=2.51 $Y=1.855 $X2=0
+ $Y2=0
cc_144 N_A_80_21#_c_116_p N_VPWR_M1017_d 0.00422875f $X=3 $Y=1.94 $X2=0 $Y2=0
cc_145 N_A_80_21#_c_160_p N_VPWR_M1017_d 0.00100096f $X=2.62 $Y=1.94 $X2=0 $Y2=0
cc_146 N_A_80_21#_c_136_p N_VPWR_M1004_d 0.00369907f $X=4.085 $Y=1.94 $X2=0
+ $Y2=0
cc_147 N_A_80_21#_c_121_p N_VPWR_M1002_s 0.00848532f $X=5.465 $Y=1.94 $X2=0
+ $Y2=0
cc_148 N_A_80_21#_c_105_n N_VPWR_c_515_n 0.0116301f $X=0.94 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_80_21#_c_106_n N_VPWR_c_515_n 5.93577e-19 $X=1.42 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_80_21#_c_105_n N_VPWR_c_516_n 6.53476e-19 $X=0.94 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_80_21#_c_106_n N_VPWR_c_516_n 0.0150594f $X=1.42 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_80_21#_c_107_n N_VPWR_c_516_n 0.0105403f $X=1.9 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_80_21#_c_108_n N_VPWR_c_516_n 5.93577e-19 $X=2.38 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_80_21#_c_107_n N_VPWR_c_517_n 5.52618e-19 $X=1.9 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_80_21#_c_108_n N_VPWR_c_517_n 0.0102575f $X=2.38 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_80_21#_c_116_p N_VPWR_c_517_n 0.00758095f $X=3 $Y=1.94 $X2=0 $Y2=0
cc_157 N_A_80_21#_c_160_p N_VPWR_c_517_n 0.0131021f $X=2.62 $Y=1.94 $X2=0 $Y2=0
cc_158 N_A_80_21#_c_141_p N_VPWR_c_518_n 0.020849f $X=3.195 $Y=2.3 $X2=0 $Y2=0
cc_159 N_A_80_21#_c_136_p N_VPWR_c_518_n 0.0200311f $X=4.085 $Y=1.94 $X2=0 $Y2=0
cc_160 N_A_80_21#_c_121_p N_VPWR_c_519_n 0.0140554f $X=5.465 $Y=1.94 $X2=0 $Y2=0
cc_161 N_A_80_21#_c_149_p N_VPWR_c_521_n 0.0154573f $X=5.68 $Y=2.02 $X2=0 $Y2=0
cc_162 N_A_80_21#_c_116_p N_VPWR_c_522_n 0.00280993f $X=3 $Y=1.94 $X2=0 $Y2=0
cc_163 N_A_80_21#_c_141_p N_VPWR_c_522_n 0.0249412f $X=3.195 $Y=2.3 $X2=0 $Y2=0
cc_164 N_A_80_21#_c_136_p N_VPWR_c_522_n 0.00213732f $X=4.085 $Y=1.94 $X2=0
+ $Y2=0
cc_165 N_A_80_21#_c_105_n N_VPWR_c_525_n 0.00661659f $X=0.94 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_80_21#_c_106_n N_VPWR_c_525_n 0.00427505f $X=1.42 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_80_21#_c_107_n N_VPWR_c_526_n 0.00661659f $X=1.9 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A_80_21#_c_108_n N_VPWR_c_526_n 0.00427505f $X=2.38 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_80_21#_c_136_p N_VPWR_c_527_n 0.00239127f $X=4.085 $Y=1.94 $X2=0
+ $Y2=0
cc_170 N_A_80_21#_c_120_p N_VPWR_c_527_n 0.0191076f $X=4.25 $Y=2.3 $X2=0 $Y2=0
cc_171 N_A_80_21#_c_121_p N_VPWR_c_527_n 0.0024395f $X=5.465 $Y=1.94 $X2=0 $Y2=0
cc_172 N_A_80_21#_c_121_p N_VPWR_c_528_n 0.00810298f $X=5.465 $Y=1.94 $X2=0
+ $Y2=0
cc_173 N_A_80_21#_c_149_p N_VPWR_c_528_n 0.0222328f $X=5.68 $Y=2.02 $X2=0 $Y2=0
cc_174 N_A_80_21#_M1001_d N_VPWR_c_514_n 0.00433794f $X=2.945 $Y=1.485 $X2=0
+ $Y2=0
cc_175 N_A_80_21#_M1014_s N_VPWR_c_514_n 0.00247321f $X=4.08 $Y=1.485 $X2=0
+ $Y2=0
cc_176 N_A_80_21#_M1006_s N_VPWR_c_514_n 0.00239291f $X=5.53 $Y=1.485 $X2=0
+ $Y2=0
cc_177 N_A_80_21#_c_105_n N_VPWR_c_514_n 0.0110408f $X=0.94 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A_80_21#_c_106_n N_VPWR_c_514_n 0.00735516f $X=1.42 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_80_21#_c_107_n N_VPWR_c_514_n 0.0110408f $X=1.9 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_80_21#_c_108_n N_VPWR_c_514_n 0.00735516f $X=2.38 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_80_21#_c_116_p N_VPWR_c_514_n 0.00578962f $X=3 $Y=1.94 $X2=0 $Y2=0
cc_182 N_A_80_21#_c_160_p N_VPWR_c_514_n 9.77785e-19 $X=2.62 $Y=1.94 $X2=0 $Y2=0
cc_183 N_A_80_21#_c_141_p N_VPWR_c_514_n 0.013743f $X=3.195 $Y=2.3 $X2=0 $Y2=0
cc_184 N_A_80_21#_c_136_p N_VPWR_c_514_n 0.00941998f $X=4.085 $Y=1.94 $X2=0
+ $Y2=0
cc_185 N_A_80_21#_c_120_p N_VPWR_c_514_n 0.0124369f $X=4.25 $Y=2.3 $X2=0 $Y2=0
cc_186 N_A_80_21#_c_121_p N_VPWR_c_514_n 0.019917f $X=5.465 $Y=1.94 $X2=0 $Y2=0
cc_187 N_A_80_21#_c_149_p N_VPWR_c_514_n 0.0140151f $X=5.68 $Y=2.02 $X2=0 $Y2=0
cc_188 N_A_80_21#_c_96_n N_X_c_629_n 0.0148988f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_80_21#_c_204_p N_X_c_629_n 0.00406679f $X=2.4 $Y=1.165 $X2=0 $Y2=0
cc_190 N_A_80_21#_c_105_n N_X_c_624_n 0.0240816f $X=0.94 $Y=1.41 $X2=0 $Y2=0
cc_191 N_A_80_21#_c_204_p N_X_c_624_n 0.04012f $X=2.4 $Y=1.165 $X2=0 $Y2=0
cc_192 N_A_80_21#_c_100_n N_X_c_624_n 0.0145033f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_80_21#_c_97_n N_X_c_634_n 0.0135395f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_80_21#_c_98_n N_X_c_634_n 0.0128738f $X=1.415 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_80_21#_c_204_p N_X_c_634_n 0.0425368f $X=2.4 $Y=1.165 $X2=0 $Y2=0
cc_196 N_A_80_21#_c_100_n N_X_c_634_n 0.00655314f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A_80_21#_c_106_n N_X_c_638_n 0.00531491f $X=1.42 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_80_21#_c_106_n N_X_c_626_n 0.0190848f $X=1.42 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A_80_21#_c_107_n N_X_c_626_n 0.0204373f $X=1.9 $Y=1.41 $X2=0 $Y2=0
cc_200 N_A_80_21#_c_108_n N_X_c_626_n 0.00200601f $X=2.38 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A_80_21#_c_204_p N_X_c_626_n 0.0724824f $X=2.4 $Y=1.165 $X2=0 $Y2=0
cc_202 N_A_80_21#_c_100_n N_X_c_626_n 0.0160724f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A_80_21#_c_102_n N_X_c_626_n 0.0213684f $X=2.51 $Y=1.855 $X2=0 $Y2=0
cc_204 N_A_80_21#_c_108_n N_X_c_645_n 0.0054687f $X=2.38 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A_80_21#_c_102_n N_X_c_645_n 0.0111166f $X=2.51 $Y=1.855 $X2=0 $Y2=0
cc_206 N_A_80_21#_c_160_p N_X_c_645_n 0.013466f $X=2.62 $Y=1.94 $X2=0 $Y2=0
cc_207 N_A_80_21#_c_96_n N_X_c_648_n 6.12342e-19 $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A_80_21#_c_204_p N_X_c_648_n 0.0095549f $X=2.4 $Y=1.165 $X2=0 $Y2=0
cc_209 N_A_80_21#_c_100_n N_X_c_648_n 0.00322408f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_210 N_A_80_21#_c_204_p N_X_c_627_n 0.014677f $X=2.4 $Y=1.165 $X2=0 $Y2=0
cc_211 N_A_80_21#_c_100_n N_X_c_627_n 0.0046779f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_80_21#_c_96_n X 0.0190162f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A_80_21#_c_105_n X 6.39036e-19 $X=0.94 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A_80_21#_c_204_p X 0.0164096f $X=2.4 $Y=1.165 $X2=0 $Y2=0
cc_215 N_A_80_21#_c_100_n X 0.00231286f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A_80_21#_c_121_p A_1010_297# 0.00540949f $X=5.465 $Y=1.94 $X2=-0.19
+ $Y2=-0.24
cc_217 N_A_80_21#_c_96_n N_VGND_c_698_n 0.00796324f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_218 N_A_80_21#_c_97_n N_VGND_c_698_n 5.21831e-19 $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_219 N_A_80_21#_c_97_n N_VGND_c_699_n 0.00170235f $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_220 N_A_80_21#_c_98_n N_VGND_c_699_n 0.0064878f $X=1.415 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A_80_21#_c_99_n N_VGND_c_699_n 4.97619e-19 $X=1.885 $Y=0.995 $X2=0
+ $Y2=0
cc_222 N_A_80_21#_c_103_n N_VGND_c_702_n 0.00365478f $X=2.62 $Y=0.725 $X2=0
+ $Y2=0
cc_223 N_A_80_21#_c_96_n N_VGND_c_706_n 0.00353537f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_224 N_A_80_21#_c_97_n N_VGND_c_706_n 0.00422112f $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_225 N_A_80_21#_c_98_n N_VGND_c_707_n 0.00401717f $X=1.415 $Y=0.995 $X2=0
+ $Y2=0
cc_226 N_A_80_21#_c_99_n N_VGND_c_707_n 0.0132813f $X=1.885 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A_80_21#_c_204_p N_VGND_c_707_n 0.0110453f $X=2.4 $Y=1.165 $X2=0 $Y2=0
cc_228 N_A_80_21#_c_100_n N_VGND_c_707_n 0.00698009f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A_80_21#_M1023_d N_VGND_c_709_n 0.00440791f $X=3.395 $Y=0.235 $X2=0
+ $Y2=0
cc_230 N_A_80_21#_c_96_n N_VGND_c_709_n 0.00421368f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_231 N_A_80_21#_c_97_n N_VGND_c_709_n 0.00578703f $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_232 N_A_80_21#_c_98_n N_VGND_c_709_n 0.0041737f $X=1.415 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_80_21#_c_99_n N_VGND_c_709_n 0.00771167f $X=1.885 $Y=0.995 $X2=0
+ $Y2=0
cc_234 N_A_80_21#_c_103_n N_VGND_c_709_n 0.00551779f $X=2.62 $Y=0.725 $X2=0
+ $Y2=0
cc_235 N_A_80_21#_c_115_p N_A_524_47#_M1008_s 0.00844235f $X=3.605 $Y=0.73
+ $X2=-0.19 $Y2=-0.24
cc_236 N_A_80_21#_M1023_d N_A_524_47#_c_797_n 0.0109193f $X=3.395 $Y=0.235 $X2=0
+ $Y2=0
cc_237 N_A_80_21#_c_103_n N_A_524_47#_c_797_n 0.00323932f $X=2.62 $Y=0.725 $X2=0
+ $Y2=0
cc_238 N_A_80_21#_c_115_p N_A_524_47#_c_797_n 0.0669402f $X=3.605 $Y=0.73 $X2=0
+ $Y2=0
cc_239 N_A_80_21#_c_115_p N_A_524_47#_c_804_n 0.00187101f $X=3.605 $Y=0.73 $X2=0
+ $Y2=0
cc_240 N_A_80_21#_c_115_p N_A_524_47#_c_805_n 0.00406359f $X=3.605 $Y=0.73 $X2=0
+ $Y2=0
cc_241 N_A_80_21#_c_115_p A_818_47# 0.00295109f $X=3.605 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_242 N_B1_c_258_n N_C1_c_341_n 0.0399482f $X=2.96 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_243 N_B1_c_257_n N_C1_c_345_n 0.0258892f $X=2.855 $Y=1.41 $X2=0 $Y2=0
cc_244 N_B1_c_261_n N_C1_c_345_n 6.99636e-19 $X=2.875 $Y=1.16 $X2=0 $Y2=0
cc_245 B1 N_C1_c_345_n 0.0161206f $X=4.27 $Y=1.445 $X2=0 $Y2=0
cc_246 N_B1_c_260_n N_C1_c_346_n 0.0336169f $X=4.485 $Y=1.41 $X2=0 $Y2=0
cc_247 B1 N_C1_c_346_n 0.0151154f $X=4.27 $Y=1.445 $X2=0 $Y2=0
cc_248 N_B1_c_262_n N_C1_c_346_n 7.98535e-19 $X=4.435 $Y=1.16 $X2=0 $Y2=0
cc_249 N_B1_c_259_n N_C1_c_342_n 0.0498851f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_250 N_B1_c_257_n N_C1_c_343_n 2.62802e-19 $X=2.855 $Y=1.41 $X2=0 $Y2=0
cc_251 N_B1_c_260_n N_C1_c_343_n 2.79707e-19 $X=4.485 $Y=1.41 $X2=0 $Y2=0
cc_252 N_B1_c_261_n N_C1_c_343_n 0.0198042f $X=2.875 $Y=1.16 $X2=0 $Y2=0
cc_253 B1 N_C1_c_343_n 0.0615379f $X=4.27 $Y=1.445 $X2=0 $Y2=0
cc_254 N_B1_c_262_n N_C1_c_343_n 0.0191246f $X=4.435 $Y=1.16 $X2=0 $Y2=0
cc_255 N_B1_c_257_n N_C1_c_344_n 0.041767f $X=2.855 $Y=1.41 $X2=0 $Y2=0
cc_256 N_B1_c_260_n N_C1_c_344_n 0.0253684f $X=4.485 $Y=1.41 $X2=0 $Y2=0
cc_257 N_B1_c_261_n N_C1_c_344_n 0.00543635f $X=2.875 $Y=1.16 $X2=0 $Y2=0
cc_258 B1 N_C1_c_344_n 0.0127918f $X=4.27 $Y=1.445 $X2=0 $Y2=0
cc_259 N_B1_c_262_n N_C1_c_344_n 0.00400401f $X=4.435 $Y=1.16 $X2=0 $Y2=0
cc_260 N_B1_c_259_n N_A1_c_388_n 0.0103831f $X=4.4 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_261 N_B1_c_260_n N_A1_c_389_n 0.0641616f $X=4.485 $Y=1.41 $X2=0 $Y2=0
cc_262 B1 N_A1_c_389_n 2.98987e-19 $X=4.27 $Y=1.445 $X2=0 $Y2=0
cc_263 N_B1_c_262_n N_A1_c_389_n 0.00217398f $X=4.435 $Y=1.16 $X2=0 $Y2=0
cc_264 N_B1_c_260_n N_A1_c_392_n 9.2565e-19 $X=4.485 $Y=1.41 $X2=0 $Y2=0
cc_265 B1 N_A1_c_392_n 0.00283176f $X=4.27 $Y=1.445 $X2=0 $Y2=0
cc_266 N_B1_c_262_n N_A1_c_392_n 0.026792f $X=4.435 $Y=1.16 $X2=0 $Y2=0
cc_267 B1 N_VPWR_M1004_d 0.00200322f $X=4.27 $Y=1.445 $X2=0 $Y2=0
cc_268 N_B1_c_257_n N_VPWR_c_517_n 0.00829753f $X=2.855 $Y=1.41 $X2=0 $Y2=0
cc_269 N_B1_c_257_n N_VPWR_c_518_n 9.42083e-19 $X=2.855 $Y=1.41 $X2=0 $Y2=0
cc_270 N_B1_c_260_n N_VPWR_c_518_n 9.62811e-19 $X=4.485 $Y=1.41 $X2=0 $Y2=0
cc_271 N_B1_c_260_n N_VPWR_c_519_n 0.00303345f $X=4.485 $Y=1.41 $X2=0 $Y2=0
cc_272 N_B1_c_257_n N_VPWR_c_522_n 0.00476322f $X=2.855 $Y=1.41 $X2=0 $Y2=0
cc_273 N_B1_c_260_n N_VPWR_c_527_n 0.00511838f $X=4.485 $Y=1.41 $X2=0 $Y2=0
cc_274 N_B1_c_257_n N_VPWR_c_514_n 0.00590401f $X=2.855 $Y=1.41 $X2=0 $Y2=0
cc_275 N_B1_c_260_n N_VPWR_c_514_n 0.00674312f $X=4.485 $Y=1.41 $X2=0 $Y2=0
cc_276 N_B1_c_258_n N_VGND_c_702_n 0.00357877f $X=2.96 $Y=0.995 $X2=0 $Y2=0
cc_277 N_B1_c_259_n N_VGND_c_702_n 0.00357877f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_278 N_B1_c_258_n N_VGND_c_707_n 0.0021963f $X=2.96 $Y=0.995 $X2=0 $Y2=0
cc_279 N_B1_c_258_n N_VGND_c_709_n 0.00641668f $X=2.96 $Y=0.995 $X2=0 $Y2=0
cc_280 N_B1_c_259_n N_VGND_c_709_n 0.00531727f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_281 N_B1_c_258_n N_A_524_47#_c_797_n 0.00812316f $X=2.96 $Y=0.995 $X2=0 $Y2=0
cc_282 N_B1_c_259_n N_A_524_47#_c_797_n 0.0102718f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_283 N_B1_c_262_n N_A_524_47#_c_797_n 0.00520326f $X=4.435 $Y=1.16 $X2=0 $Y2=0
cc_284 N_B1_c_260_n N_A_524_47#_c_805_n 0.00291696f $X=4.485 $Y=1.41 $X2=0 $Y2=0
cc_285 N_B1_c_262_n N_A_524_47#_c_805_n 0.00824741f $X=4.435 $Y=1.16 $X2=0 $Y2=0
cc_286 N_C1_c_345_n N_VPWR_c_517_n 8.67235e-19 $X=3.51 $Y=1.41 $X2=0 $Y2=0
cc_287 N_C1_c_345_n N_VPWR_c_518_n 0.0112559f $X=3.51 $Y=1.41 $X2=0 $Y2=0
cc_288 N_C1_c_346_n N_VPWR_c_518_n 0.00798483f $X=3.99 $Y=1.41 $X2=0 $Y2=0
cc_289 N_C1_c_345_n N_VPWR_c_522_n 0.0033175f $X=3.51 $Y=1.41 $X2=0 $Y2=0
cc_290 N_C1_c_346_n N_VPWR_c_527_n 0.00476322f $X=3.99 $Y=1.41 $X2=0 $Y2=0
cc_291 N_C1_c_345_n N_VPWR_c_514_n 0.00442855f $X=3.51 $Y=1.41 $X2=0 $Y2=0
cc_292 N_C1_c_346_n N_VPWR_c_514_n 0.0055254f $X=3.99 $Y=1.41 $X2=0 $Y2=0
cc_293 N_C1_c_341_n N_VGND_c_702_n 0.00357877f $X=3.32 $Y=0.995 $X2=0 $Y2=0
cc_294 N_C1_c_342_n N_VGND_c_702_n 0.00357877f $X=4.015 $Y=0.995 $X2=0 $Y2=0
cc_295 N_C1_c_341_n N_VGND_c_709_n 0.00572034f $X=3.32 $Y=0.995 $X2=0 $Y2=0
cc_296 N_C1_c_342_n N_VGND_c_709_n 0.00579034f $X=4.015 $Y=0.995 $X2=0 $Y2=0
cc_297 N_C1_c_341_n N_A_524_47#_c_797_n 0.0120961f $X=3.32 $Y=0.995 $X2=0 $Y2=0
cc_298 N_C1_c_342_n N_A_524_47#_c_797_n 0.0142615f $X=4.015 $Y=0.995 $X2=0 $Y2=0
cc_299 N_C1_c_343_n N_A_524_47#_c_797_n 0.00646074f $X=3.875 $Y=1.16 $X2=0 $Y2=0
cc_300 N_C1_c_344_n N_A_524_47#_c_797_n 9.21206e-19 $X=3.99 $Y=1.202 $X2=0 $Y2=0
cc_301 N_A1_c_388_n N_A2_c_461_n 0.0216271f $X=4.875 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_302 N_A1_c_389_n N_A2_c_465_n 0.0512846f $X=4.96 $Y=1.41 $X2=0 $Y2=0
cc_303 N_A1_c_392_n N_A2_c_465_n 0.00194785f $X=4.99 $Y=1.16 $X2=0 $Y2=0
cc_304 N_A1_c_402_n N_A2_c_465_n 0.0128446f $X=6.3 $Y=1.59 $X2=0 $Y2=0
cc_305 N_A1_c_390_n N_A2_c_462_n 0.0219536f $X=6.375 $Y=0.995 $X2=0 $Y2=0
cc_306 N_A1_c_391_n N_A2_c_466_n 0.0502727f $X=6.4 $Y=1.41 $X2=0 $Y2=0
cc_307 N_A1_c_402_n N_A2_c_466_n 0.0176526f $X=6.3 $Y=1.59 $X2=0 $Y2=0
cc_308 N_A1_c_393_n N_A2_c_466_n 0.00170661f $X=6.495 $Y=1.16 $X2=0 $Y2=0
cc_309 N_A1_c_389_n N_A2_c_463_n 0.025595f $X=4.96 $Y=1.41 $X2=0 $Y2=0
cc_310 N_A1_c_391_n N_A2_c_463_n 0.0258696f $X=6.4 $Y=1.41 $X2=0 $Y2=0
cc_311 N_A1_c_392_n N_A2_c_463_n 0.00297212f $X=4.99 $Y=1.16 $X2=0 $Y2=0
cc_312 N_A1_c_402_n N_A2_c_463_n 0.00806196f $X=6.3 $Y=1.59 $X2=0 $Y2=0
cc_313 N_A1_c_393_n N_A2_c_463_n 8.83304e-19 $X=6.495 $Y=1.16 $X2=0 $Y2=0
cc_314 N_A1_c_389_n N_A2_c_464_n 3.41803e-19 $X=4.96 $Y=1.41 $X2=0 $Y2=0
cc_315 N_A1_c_391_n N_A2_c_464_n 0.00184721f $X=6.4 $Y=1.41 $X2=0 $Y2=0
cc_316 N_A1_c_392_n N_A2_c_464_n 0.0226678f $X=4.99 $Y=1.16 $X2=0 $Y2=0
cc_317 N_A1_c_402_n N_A2_c_464_n 0.0496628f $X=6.3 $Y=1.59 $X2=0 $Y2=0
cc_318 N_A1_c_393_n N_A2_c_464_n 0.0235053f $X=6.495 $Y=1.16 $X2=0 $Y2=0
cc_319 N_A1_c_393_n N_VPWR_M1011_d 0.00365535f $X=6.495 $Y=1.16 $X2=0 $Y2=0
cc_320 N_A1_c_389_n N_VPWR_c_519_n 0.00309306f $X=4.96 $Y=1.41 $X2=0 $Y2=0
cc_321 N_A1_c_391_n N_VPWR_c_521_n 0.0214786f $X=6.4 $Y=1.41 $X2=0 $Y2=0
cc_322 N_A1_c_393_n N_VPWR_c_521_n 0.0227717f $X=6.495 $Y=1.16 $X2=0 $Y2=0
cc_323 N_A1_c_389_n N_VPWR_c_528_n 0.0052046f $X=4.96 $Y=1.41 $X2=0 $Y2=0
cc_324 N_A1_c_391_n N_VPWR_c_528_n 0.00447018f $X=6.4 $Y=1.41 $X2=0 $Y2=0
cc_325 N_A1_c_389_n N_VPWR_c_514_n 0.00683647f $X=4.96 $Y=1.41 $X2=0 $Y2=0
cc_326 N_A1_c_391_n N_VPWR_c_514_n 0.00776557f $X=6.4 $Y=1.41 $X2=0 $Y2=0
cc_327 N_A1_c_402_n A_1010_297# 0.00427495f $X=6.3 $Y=1.59 $X2=-0.19 $Y2=-0.24
cc_328 N_A1_c_405_n A_1010_297# 5.20676e-19 $X=5.155 $Y=1.59 $X2=-0.19 $Y2=-0.24
cc_329 N_A1_c_402_n A_1202_297# 0.0104842f $X=6.3 $Y=1.59 $X2=-0.19 $Y2=-0.24
cc_330 N_A1_c_388_n N_VGND_c_700_n 0.00315768f $X=4.875 $Y=0.995 $X2=0 $Y2=0
cc_331 N_A1_c_390_n N_VGND_c_701_n 0.00283414f $X=6.375 $Y=0.995 $X2=0 $Y2=0
cc_332 N_A1_c_388_n N_VGND_c_702_n 0.00431182f $X=4.875 $Y=0.995 $X2=0 $Y2=0
cc_333 N_A1_c_390_n N_VGND_c_708_n 0.0042256f $X=6.375 $Y=0.995 $X2=0 $Y2=0
cc_334 N_A1_c_388_n N_VGND_c_709_n 0.00615698f $X=4.875 $Y=0.995 $X2=0 $Y2=0
cc_335 N_A1_c_390_n N_VGND_c_709_n 0.00684075f $X=6.375 $Y=0.995 $X2=0 $Y2=0
cc_336 N_A1_c_388_n N_A_524_47#_c_815_n 0.00190274f $X=4.875 $Y=0.995 $X2=0
+ $Y2=0
cc_337 N_A1_c_388_n N_A_524_47#_c_804_n 0.00369077f $X=4.875 $Y=0.995 $X2=0
+ $Y2=0
cc_338 N_A1_c_388_n N_A_524_47#_c_817_n 0.0108633f $X=4.875 $Y=0.995 $X2=0 $Y2=0
cc_339 N_A1_c_389_n N_A_524_47#_c_817_n 0.00451584f $X=4.96 $Y=1.41 $X2=0 $Y2=0
cc_340 N_A1_c_392_n N_A_524_47#_c_817_n 0.0234144f $X=4.99 $Y=1.16 $X2=0 $Y2=0
cc_341 N_A1_c_402_n N_A_524_47#_c_817_n 0.00363505f $X=6.3 $Y=1.59 $X2=0 $Y2=0
cc_342 N_A1_c_388_n N_A_524_47#_c_821_n 5.15987e-19 $X=4.875 $Y=0.995 $X2=0
+ $Y2=0
cc_343 N_A1_c_390_n N_A_524_47#_c_821_n 5.3197e-19 $X=6.375 $Y=0.995 $X2=0 $Y2=0
cc_344 N_A1_c_390_n N_A_524_47#_c_798_n 0.00963893f $X=6.375 $Y=0.995 $X2=0
+ $Y2=0
cc_345 N_A1_c_391_n N_A_524_47#_c_798_n 0.00728853f $X=6.4 $Y=1.41 $X2=0 $Y2=0
cc_346 N_A1_c_402_n N_A_524_47#_c_798_n 0.00364888f $X=6.3 $Y=1.59 $X2=0 $Y2=0
cc_347 N_A1_c_393_n N_A_524_47#_c_798_n 0.0398854f $X=6.495 $Y=1.16 $X2=0 $Y2=0
cc_348 N_A1_c_390_n N_A_524_47#_c_799_n 0.00607657f $X=6.375 $Y=0.995 $X2=0
+ $Y2=0
cc_349 N_A2_c_466_n N_VPWR_c_521_n 0.00287102f $X=5.92 $Y=1.41 $X2=0 $Y2=0
cc_350 N_A2_c_465_n N_VPWR_c_528_n 0.00489024f $X=5.44 $Y=1.41 $X2=0 $Y2=0
cc_351 N_A2_c_466_n N_VPWR_c_528_n 0.00681208f $X=5.92 $Y=1.41 $X2=0 $Y2=0
cc_352 N_A2_c_465_n N_VPWR_c_514_n 0.00671454f $X=5.44 $Y=1.41 $X2=0 $Y2=0
cc_353 N_A2_c_466_n N_VPWR_c_514_n 0.0122805f $X=5.92 $Y=1.41 $X2=0 $Y2=0
cc_354 N_A2_c_461_n N_VGND_c_700_n 0.00471866f $X=5.415 $Y=0.995 $X2=0 $Y2=0
cc_355 N_A2_c_462_n N_VGND_c_701_n 0.00380362f $X=5.895 $Y=0.995 $X2=0 $Y2=0
cc_356 N_A2_c_461_n N_VGND_c_704_n 0.0042256f $X=5.415 $Y=0.995 $X2=0 $Y2=0
cc_357 N_A2_c_462_n N_VGND_c_704_n 0.0042256f $X=5.895 $Y=0.995 $X2=0 $Y2=0
cc_358 N_A2_c_461_n N_VGND_c_709_n 0.00616982f $X=5.415 $Y=0.995 $X2=0 $Y2=0
cc_359 N_A2_c_462_n N_VGND_c_709_n 0.00611417f $X=5.895 $Y=0.995 $X2=0 $Y2=0
cc_360 N_A2_c_461_n N_A_524_47#_c_804_n 5.24878e-19 $X=5.415 $Y=0.995 $X2=0
+ $Y2=0
cc_361 N_A2_c_461_n N_A_524_47#_c_817_n 0.00923148f $X=5.415 $Y=0.995 $X2=0
+ $Y2=0
cc_362 N_A2_c_464_n N_A_524_47#_c_817_n 0.00880077f $X=5.895 $Y=1.16 $X2=0 $Y2=0
cc_363 N_A2_c_461_n N_A_524_47#_c_821_n 0.00636077f $X=5.415 $Y=0.995 $X2=0
+ $Y2=0
cc_364 N_A2_c_462_n N_A_524_47#_c_821_n 0.00639223f $X=5.895 $Y=0.995 $X2=0
+ $Y2=0
cc_365 N_A2_c_462_n N_A_524_47#_c_798_n 0.00894266f $X=5.895 $Y=0.995 $X2=0
+ $Y2=0
cc_366 N_A2_c_463_n N_A_524_47#_c_798_n 0.0028605f $X=5.895 $Y=1.16 $X2=0 $Y2=0
cc_367 N_A2_c_464_n N_A_524_47#_c_798_n 0.0174317f $X=5.895 $Y=1.16 $X2=0 $Y2=0
cc_368 N_A2_c_462_n N_A_524_47#_c_799_n 5.13858e-19 $X=5.895 $Y=0.995 $X2=0
+ $Y2=0
cc_369 N_A2_c_461_n N_A_524_47#_c_837_n 7.16038e-19 $X=5.415 $Y=0.995 $X2=0
+ $Y2=0
cc_370 N_A2_c_462_n N_A_524_47#_c_837_n 7.16038e-19 $X=5.895 $Y=0.995 $X2=0
+ $Y2=0
cc_371 N_A2_c_463_n N_A_524_47#_c_837_n 0.00364896f $X=5.895 $Y=1.16 $X2=0 $Y2=0
cc_372 N_A2_c_464_n N_A_524_47#_c_837_n 0.0255748f $X=5.895 $Y=1.16 $X2=0 $Y2=0
cc_373 N_VPWR_c_514_n N_X_M1005_s 0.00655879f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_374 N_VPWR_c_514_n N_X_M1012_s 0.00621163f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_375 N_VPWR_M1005_d N_X_c_624_n 0.00471874f $X=0.52 $Y=1.485 $X2=0 $Y2=0
cc_376 N_VPWR_c_515_n N_X_c_624_n 0.0269571f $X=0.695 $Y=1.955 $X2=0 $Y2=0
cc_377 N_VPWR_c_516_n N_X_c_638_n 0.0426768f $X=1.655 $Y=1.955 $X2=0 $Y2=0
cc_378 N_VPWR_c_525_n N_X_c_638_n 0.012308f $X=1.44 $Y=2.72 $X2=0 $Y2=0
cc_379 N_VPWR_c_514_n N_X_c_638_n 0.00685509f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_380 N_VPWR_M1010_d N_X_c_626_n 0.00200444f $X=1.51 $Y=1.485 $X2=0 $Y2=0
cc_381 N_VPWR_c_516_n N_X_c_626_n 0.0216439f $X=1.655 $Y=1.955 $X2=0 $Y2=0
cc_382 N_VPWR_c_517_n N_X_c_645_n 0.0199455f $X=2.615 $Y=2.32 $X2=0 $Y2=0
cc_383 N_VPWR_c_526_n N_X_c_645_n 0.0130112f $X=2.4 $Y=2.72 $X2=0 $Y2=0
cc_384 N_VPWR_c_514_n N_X_c_645_n 0.00724021f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_385 N_VPWR_c_514_n A_1010_297# 0.00376671f $X=6.67 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_386 N_VPWR_c_514_n A_1202_297# 0.0128237f $X=6.67 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_387 N_X_c_622_n N_VGND_M1009_s 0.00301407f $X=0.225 $Y=0.805 $X2=-0.19
+ $Y2=-0.24
cc_388 X N_VGND_M1009_s 3.71677e-19 $X=0.23 $Y=0.85 $X2=-0.19 $Y2=-0.24
cc_389 N_X_c_634_n N_VGND_M1013_s 0.00432468f $X=1.585 $Y=0.71 $X2=0 $Y2=0
cc_390 N_X_c_622_n N_VGND_c_697_n 2.03606e-19 $X=0.225 $Y=0.805 $X2=0 $Y2=0
cc_391 N_X_c_629_n N_VGND_c_698_n 0.00167305f $X=0.645 $Y=0.72 $X2=0 $Y2=0
cc_392 N_X_c_674_p N_VGND_c_698_n 0.012714f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_393 N_X_c_622_n N_VGND_c_698_n 0.0209438f $X=0.225 $Y=0.805 $X2=0 $Y2=0
cc_394 N_X_c_634_n N_VGND_c_699_n 0.017404f $X=1.585 $Y=0.71 $X2=0 $Y2=0
cc_395 N_X_c_677_p N_VGND_c_699_n 0.0115031f $X=1.67 $Y=0.42 $X2=0 $Y2=0
cc_396 N_X_c_629_n N_VGND_c_706_n 0.00325081f $X=0.645 $Y=0.72 $X2=0 $Y2=0
cc_397 N_X_c_674_p N_VGND_c_706_n 0.0115988f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_398 N_X_c_634_n N_VGND_c_706_n 0.00330209f $X=1.585 $Y=0.71 $X2=0 $Y2=0
cc_399 N_X_c_634_n N_VGND_c_707_n 0.00342879f $X=1.585 $Y=0.71 $X2=0 $Y2=0
cc_400 N_X_c_677_p N_VGND_c_707_n 0.0115988f $X=1.67 $Y=0.42 $X2=0 $Y2=0
cc_401 N_X_M1009_d N_VGND_c_709_n 0.00306192f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_402 N_X_M1021_d N_VGND_c_709_n 0.00477085f $X=1.49 $Y=0.235 $X2=0 $Y2=0
cc_403 N_X_c_629_n N_VGND_c_709_n 0.00584642f $X=0.645 $Y=0.72 $X2=0 $Y2=0
cc_404 N_X_c_674_p N_VGND_c_709_n 0.00642947f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_405 N_X_c_634_n N_VGND_c_709_n 0.0127472f $X=1.585 $Y=0.71 $X2=0 $Y2=0
cc_406 N_X_c_677_p N_VGND_c_709_n 0.00642947f $X=1.67 $Y=0.42 $X2=0 $Y2=0
cc_407 N_X_c_622_n N_VGND_c_709_n 0.00170408f $X=0.225 $Y=0.805 $X2=0 $Y2=0
cc_408 N_VGND_c_709_n N_A_524_47#_M1008_s 0.00213443f $X=6.67 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_409 N_VGND_c_709_n N_A_524_47#_M1015_s 0.00259365f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_410 N_VGND_c_709_n N_A_524_47#_M1000_d 0.0026338f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_411 N_VGND_c_709_n N_A_524_47#_M1016_d 0.00254408f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_412 N_VGND_c_702_n N_A_524_47#_c_797_n 0.109102f $X=4.98 $Y=0 $X2=0 $Y2=0
cc_413 N_VGND_c_707_n N_A_524_47#_c_797_n 0.014688f $X=1.925 $Y=0 $X2=0 $Y2=0
cc_414 N_VGND_c_709_n N_A_524_47#_c_797_n 0.0680659f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_415 N_VGND_c_702_n N_A_524_47#_c_815_n 0.0190711f $X=4.98 $Y=0 $X2=0 $Y2=0
cc_416 N_VGND_c_709_n N_A_524_47#_c_815_n 0.0125393f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_417 N_VGND_M1007_s N_A_524_47#_c_817_n 0.00699963f $X=4.95 $Y=0.235 $X2=0
+ $Y2=0
cc_418 N_VGND_c_700_n N_A_524_47#_c_817_n 0.0214325f $X=5.13 $Y=0.36 $X2=0 $Y2=0
cc_419 N_VGND_c_702_n N_A_524_47#_c_817_n 0.00230889f $X=4.98 $Y=0 $X2=0 $Y2=0
cc_420 N_VGND_c_704_n N_A_524_47#_c_817_n 0.0021487f $X=6.065 $Y=0 $X2=0 $Y2=0
cc_421 N_VGND_c_709_n N_A_524_47#_c_817_n 0.00917919f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_422 N_VGND_c_701_n N_A_524_47#_c_821_n 0.0166628f $X=6.16 $Y=0.36 $X2=0 $Y2=0
cc_423 N_VGND_c_704_n N_A_524_47#_c_821_n 0.0222964f $X=6.065 $Y=0 $X2=0 $Y2=0
cc_424 N_VGND_c_709_n N_A_524_47#_c_821_n 0.0141522f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_425 N_VGND_M1003_s N_A_524_47#_c_798_n 0.00593833f $X=5.97 $Y=0.235 $X2=0
+ $Y2=0
cc_426 N_VGND_c_701_n N_A_524_47#_c_798_n 0.0137448f $X=6.16 $Y=0.36 $X2=0 $Y2=0
cc_427 N_VGND_c_704_n N_A_524_47#_c_798_n 0.00283421f $X=6.065 $Y=0 $X2=0 $Y2=0
cc_428 N_VGND_c_708_n N_A_524_47#_c_798_n 0.0021487f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_429 N_VGND_c_709_n N_A_524_47#_c_798_n 0.0100001f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_430 N_VGND_c_708_n N_A_524_47#_c_799_n 0.024386f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_431 N_VGND_c_709_n N_A_524_47#_c_799_n 0.0143342f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_432 N_VGND_c_709_n A_818_47# 0.00168648f $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24
cc_433 N_VGND_c_709_n A_607_47# 0.00188725f $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24
cc_434 N_A_524_47#_c_797_n A_818_47# 0.00193721f $X=4.475 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_435 N_A_524_47#_c_797_n A_607_47# 0.00588031f $X=4.475 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
