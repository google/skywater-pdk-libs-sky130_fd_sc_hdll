* File: sky130_fd_sc_hdll__mux2_12.pex.spice
* Created: Wed Sep  2 08:34:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUX2_12%A1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39
r88 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.88 $Y=1.202
+ $X2=1.905 $Y2=1.202
r89 37 39 16.8441 $w=3.72e-07 $l=1.3e-07 $layer=POLY_cond $X=1.75 $Y=1.202
+ $X2=1.88 $Y2=1.202
r90 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.75
+ $Y=1.16 $X2=1.75 $Y2=1.16
r91 35 37 37.5753 $w=3.72e-07 $l=2.9e-07 $layer=POLY_cond $X=1.46 $Y=1.202
+ $X2=1.75 $Y2=1.202
r92 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.46 $Y2=1.202
r93 33 34 60.8979 $w=3.72e-07 $l=4.7e-07 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=1.435 $Y2=1.202
r94 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.202
+ $X2=0.965 $Y2=1.202
r95 30 32 27.2097 $w=3.72e-07 $l=2.1e-07 $layer=POLY_cond $X=0.73 $Y=1.202
+ $X2=0.94 $Y2=1.202
r96 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.73
+ $Y=1.16 $X2=0.73 $Y2=1.16
r97 28 30 27.2097 $w=3.72e-07 $l=2.1e-07 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.73 $Y2=1.202
r98 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r99 25 38 27.6586 $w=2.48e-07 $l=6e-07 $layer=LI1_cond $X=1.15 $Y=1.2 $X2=1.75
+ $Y2=1.2
r100 25 31 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=1.15 $Y=1.2 $X2=0.73
+ $Y2=1.2
r101 22 40 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r102 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r103 19 39 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.88 $Y=0.995
+ $X2=1.88 $Y2=1.202
r104 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.88 $Y=0.995
+ $X2=1.88 $Y2=0.56
r105 16 35 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=1.202
r106 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=0.56
r107 13 34 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r108 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r109 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r110 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r111 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=1.202
r112 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=0.56
r113 4 28 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r114 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=0.56
r115 1 27 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r116 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_12%S 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 43 55
r124 55 56 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.22 $Y=1.202
+ $X2=5.245 $Y2=1.202
r125 54 55 54.7135 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.8 $Y=1.202
+ $X2=5.22 $Y2=1.202
r126 53 54 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=4.775 $Y=1.202
+ $X2=4.8 $Y2=1.202
r127 52 53 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=4.305 $Y=1.202
+ $X2=4.775 $Y2=1.202
r128 51 52 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=4.28 $Y=1.202
+ $X2=4.305 $Y2=1.202
r129 49 51 22.1459 $w=3.7e-07 $l=1.7e-07 $layer=POLY_cond $X=4.11 $Y=1.202
+ $X2=4.28 $Y2=1.202
r130 47 49 32.5676 $w=3.7e-07 $l=2.5e-07 $layer=POLY_cond $X=3.86 $Y=1.202
+ $X2=4.11 $Y2=1.202
r131 46 47 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=3.835 $Y=1.202
+ $X2=3.86 $Y2=1.202
r132 45 46 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=3.365 $Y=1.202
+ $X2=3.835 $Y2=1.202
r133 44 45 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=3.34 $Y=1.202
+ $X2=3.365 $Y2=1.202
r134 43 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.11
+ $Y=1.16 $X2=4.11 $Y2=1.16
r135 42 44 32.5676 $w=3.7e-07 $l=2.5e-07 $layer=POLY_cond $X=3.09 $Y=1.202
+ $X2=3.34 $Y2=1.202
r136 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.09
+ $Y=1.16 $X2=3.09 $Y2=1.16
r137 40 42 22.1459 $w=3.7e-07 $l=1.7e-07 $layer=POLY_cond $X=2.92 $Y=1.202
+ $X2=3.09 $Y2=1.202
r138 39 40 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=2.895 $Y=1.202
+ $X2=2.92 $Y2=1.202
r139 37 43 0.271111 $w=1.348e-06 $l=3e-08 $layer=LI1_cond $X=3.6 $Y=1.19 $X2=3.6
+ $Y2=1.16
r140 34 56 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.202
r141 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.985
r142 31 55 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.22 $Y=0.995
+ $X2=5.22 $Y2=1.202
r143 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.22 $Y=0.995
+ $X2=5.22 $Y2=0.56
r144 28 54 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.8 $Y=0.995
+ $X2=4.8 $Y2=1.202
r145 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.8 $Y=0.995
+ $X2=4.8 $Y2=0.56
r146 25 53 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.202
r147 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
r148 22 52 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.202
r149 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.985
r150 19 51 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.28 $Y=0.995
+ $X2=4.28 $Y2=1.202
r151 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.28 $Y=0.995
+ $X2=4.28 $Y2=0.56
r152 16 47 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.86 $Y=0.995
+ $X2=3.86 $Y2=1.202
r153 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.86 $Y=0.995
+ $X2=3.86 $Y2=0.56
r154 13 46 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.202
r155 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.985
r156 10 45 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.202
r157 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.985
r158 7 44 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.34 $Y=0.995
+ $X2=3.34 $Y2=1.202
r159 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.34 $Y=0.995
+ $X2=3.34 $Y2=0.56
r160 4 40 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.92 $Y=0.995
+ $X2=2.92 $Y2=1.202
r161 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.92 $Y=0.995
+ $X2=2.92 $Y2=0.56
r162 1 39 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.202
r163 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_12%A_973_297# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 33 37 46 49 58
r122 58 59 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.1 $Y=1.202
+ $X2=7.125 $Y2=1.202
r123 55 56 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.655 $Y=1.202
+ $X2=6.68 $Y2=1.202
r124 54 55 60.8979 $w=3.72e-07 $l=4.7e-07 $layer=POLY_cond $X=6.185 $Y=1.202
+ $X2=6.655 $Y2=1.202
r125 53 54 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.16 $Y=1.202
+ $X2=6.185 $Y2=1.202
r126 50 51 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.715 $Y=1.202
+ $X2=5.74 $Y2=1.202
r127 47 58 22.0269 $w=3.72e-07 $l=1.7e-07 $layer=POLY_cond $X=6.93 $Y=1.202
+ $X2=7.1 $Y2=1.202
r128 47 56 32.3925 $w=3.72e-07 $l=2.5e-07 $layer=POLY_cond $X=6.93 $Y=1.202
+ $X2=6.68 $Y2=1.202
r129 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.93
+ $Y=1.16 $X2=6.93 $Y2=1.16
r130 44 53 32.3925 $w=3.72e-07 $l=2.5e-07 $layer=POLY_cond $X=5.91 $Y=1.202
+ $X2=6.16 $Y2=1.202
r131 44 51 22.0269 $w=3.72e-07 $l=1.7e-07 $layer=POLY_cond $X=5.91 $Y=1.202
+ $X2=5.74 $Y2=1.202
r132 43 46 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=5.91 $Y=1.2
+ $X2=6.93 $Y2=1.2
r133 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.91
+ $Y=1.16 $X2=5.91 $Y2=1.16
r134 41 49 2.3589 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.175 $Y=1.2
+ $X2=5.01 $Y2=1.2
r135 41 43 33.8818 $w=2.48e-07 $l=7.35e-07 $layer=LI1_cond $X=5.175 $Y=1.2
+ $X2=5.91 $Y2=1.2
r136 37 39 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.01 $Y=1.66
+ $X2=5.01 $Y2=2.34
r137 35 49 4.07664 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=5.01 $Y=1.325
+ $X2=5.01 $Y2=1.2
r138 35 37 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.01 $Y=1.325
+ $X2=5.01 $Y2=1.66
r139 31 49 4.07664 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=5.01 $Y=1.075
+ $X2=5.01 $Y2=1.2
r140 31 33 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=5.01 $Y=1.075
+ $X2=5.01 $Y2=0.42
r141 28 59 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.202
r142 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.985
r143 25 58 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.1 $Y=0.995
+ $X2=7.1 $Y2=1.202
r144 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.1 $Y=0.995
+ $X2=7.1 $Y2=0.56
r145 22 56 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.68 $Y=0.995
+ $X2=6.68 $Y2=1.202
r146 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.68 $Y=0.995
+ $X2=6.68 $Y2=0.56
r147 19 55 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.202
r148 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.985
r149 16 54 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.202
r150 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.985
r151 13 53 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=1.202
r152 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=0.56
r153 10 51 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.74 $Y=0.995
+ $X2=5.74 $Y2=1.202
r154 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.74 $Y=0.995
+ $X2=5.74 $Y2=0.56
r155 7 50 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.202
r156 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.985
r157 2 39 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=2.34
r158 2 37 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=1.66
r159 1 33 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=4.875
+ $Y=0.235 $X2=5.01 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_12%A0 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39
r92 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=9.5 $Y=1.202
+ $X2=9.525 $Y2=1.202
r93 37 39 27.2097 $w=3.72e-07 $l=2.1e-07 $layer=POLY_cond $X=9.29 $Y=1.202
+ $X2=9.5 $Y2=1.202
r94 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.29
+ $Y=1.16 $X2=9.29 $Y2=1.16
r95 35 37 27.2097 $w=3.72e-07 $l=2.1e-07 $layer=POLY_cond $X=9.08 $Y=1.202
+ $X2=9.29 $Y2=1.202
r96 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=9.055 $Y=1.202
+ $X2=9.08 $Y2=1.202
r97 33 34 60.8979 $w=3.72e-07 $l=4.7e-07 $layer=POLY_cond $X=8.585 $Y=1.202
+ $X2=9.055 $Y2=1.202
r98 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.56 $Y=1.202
+ $X2=8.585 $Y2=1.202
r99 30 32 37.5753 $w=3.72e-07 $l=2.9e-07 $layer=POLY_cond $X=8.27 $Y=1.202
+ $X2=8.56 $Y2=1.202
r100 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.27
+ $Y=1.16 $X2=8.27 $Y2=1.16
r101 28 30 16.8441 $w=3.72e-07 $l=1.3e-07 $layer=POLY_cond $X=8.14 $Y=1.202
+ $X2=8.27 $Y2=1.202
r102 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.115 $Y=1.202
+ $X2=8.14 $Y2=1.202
r103 25 38 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=8.97 $Y=1.2
+ $X2=9.29 $Y2=1.2
r104 25 31 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=8.97 $Y=1.2 $X2=8.27
+ $Y2=1.2
r105 22 40 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.525 $Y=1.41
+ $X2=9.525 $Y2=1.202
r106 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.525 $Y=1.41
+ $X2=9.525 $Y2=1.985
r107 19 39 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.5 $Y=0.995
+ $X2=9.5 $Y2=1.202
r108 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.5 $Y=0.995
+ $X2=9.5 $Y2=0.56
r109 16 35 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.08 $Y=0.995
+ $X2=9.08 $Y2=1.202
r110 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.08 $Y=0.995
+ $X2=9.08 $Y2=0.56
r111 13 34 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.055 $Y=1.41
+ $X2=9.055 $Y2=1.202
r112 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.055 $Y=1.41
+ $X2=9.055 $Y2=1.985
r113 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.585 $Y=1.41
+ $X2=8.585 $Y2=1.202
r114 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.585 $Y=1.41
+ $X2=8.585 $Y2=1.985
r115 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.56 $Y=0.995
+ $X2=8.56 $Y2=1.202
r116 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.56 $Y=0.995
+ $X2=8.56 $Y2=0.56
r117 4 28 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.14 $Y=0.995
+ $X2=8.14 $Y2=1.202
r118 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.14 $Y=0.995
+ $X2=8.14 $Y2=0.56
r119 1 27 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.115 $Y=1.41
+ $X2=8.115 $Y2=1.202
r120 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.115 $Y=1.41
+ $X2=8.115 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_12%A_27_47# 1 2 3 4 5 6 7 8 9 10 11 12 37 39
+ 40 42 43 45 46 48 49 51 52 54 55 57 58 60 61 63 64 66 67 69 70 72 73 75 76 78
+ 79 81 82 84 85 87 88 90 91 93 94 96 97 99 100 102 103 105 106 108 111 115 119
+ 121 123 125 127 131 135 137 139 142 144 150 153 156 161 162 163 165 166 173
+ 178 179 180 181 185 188 189 192 195 196 222
c480 195 0 1.96891e-19 $X=9.76 $Y=0.51
c481 189 0 1.96891e-19 $X=0.405 $Y=0.51
r482 222 223 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=15.66 $Y=1.202
+ $X2=15.685 $Y2=1.202
r483 221 222 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=15.24 $Y=1.202
+ $X2=15.66 $Y2=1.202
r484 220 221 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=15.215 $Y=1.202
+ $X2=15.24 $Y2=1.202
r485 219 220 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=14.745 $Y=1.202
+ $X2=15.215 $Y2=1.202
r486 218 219 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=14.72 $Y=1.202
+ $X2=14.745 $Y2=1.202
r487 215 216 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=14.275 $Y=1.202
+ $X2=14.3 $Y2=1.202
r488 214 215 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=13.805 $Y=1.202
+ $X2=14.275 $Y2=1.202
r489 213 214 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=13.78 $Y=1.202
+ $X2=13.805 $Y2=1.202
r490 212 213 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=13.36 $Y=1.202
+ $X2=13.78 $Y2=1.202
r491 211 212 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=13.335 $Y=1.202
+ $X2=13.36 $Y2=1.202
r492 210 211 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=12.865 $Y=1.202
+ $X2=13.335 $Y2=1.202
r493 209 210 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=12.84 $Y=1.202
+ $X2=12.865 $Y2=1.202
r494 208 209 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=12.42 $Y=1.202
+ $X2=12.84 $Y2=1.202
r495 207 208 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=12.395 $Y=1.202
+ $X2=12.42 $Y2=1.202
r496 206 207 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=11.925 $Y=1.202
+ $X2=12.395 $Y2=1.202
r497 205 206 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=11.9 $Y=1.202
+ $X2=11.925 $Y2=1.202
r498 204 205 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=11.48 $Y=1.202
+ $X2=11.9 $Y2=1.202
r499 203 204 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=11.455 $Y=1.202
+ $X2=11.48 $Y2=1.202
r500 202 203 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=10.985 $Y=1.202
+ $X2=11.455 $Y2=1.202
r501 201 202 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=10.96 $Y=1.202
+ $X2=10.985 $Y2=1.202
r502 198 199 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=10.515 $Y=1.202
+ $X2=10.54 $Y2=1.202
r503 195 196 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.76 $Y=0.51
+ $X2=9.76 $Y2=0.51
r504 192 226 44.177 $w=2.98e-07 $l=1.15e-06 $layer=LI1_cond $X=0.245 $Y=0.51
+ $X2=0.245 $Y2=1.66
r505 191 192 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=0.51
+ $X2=0.26 $Y2=0.51
r506 189 191 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.405 $Y=0.51
+ $X2=0.26 $Y2=0.51
r507 188 195 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.615 $Y=0.51
+ $X2=9.76 $Y2=0.51
r508 188 189 11.3985 $w=1.4e-07 $l=9.21e-06 $layer=MET1_cond $X=9.615 $Y=0.51
+ $X2=0.405 $Y2=0.51
r509 184 196 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=9.775 $Y=1.075
+ $X2=9.775 $Y2=0.51
r510 184 185 4.4274 $w=3e-07 $l=1.25e-07 $layer=LI1_cond $X=9.775 $Y=1.075
+ $X2=9.775 $Y2=1.2
r511 181 196 3.26526 $w=2.98e-07 $l=8.5e-08 $layer=LI1_cond $X=9.775 $Y=0.425
+ $X2=9.775 $Y2=0.51
r512 181 183 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.775 $Y=0.425
+ $X2=9.775 $Y2=0.34
r513 177 179 7.32169 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=8.82 $Y=0.4
+ $X2=8.955 $Y2=0.4
r514 177 178 7.32169 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=8.82 $Y=0.4
+ $X2=8.685 $Y2=0.4
r515 173 178 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.015 $Y=0.34
+ $X2=8.685 $Y2=0.34
r516 171 173 7.32568 $w=2.93e-07 $l=1.35e-07 $layer=LI1_cond $X=7.88 $Y=0.402
+ $X2=8.015 $Y2=0.402
r517 165 166 7.32568 $w=2.93e-07 $l=1.35e-07 $layer=LI1_cond $X=2.14 $Y=0.402
+ $X2=2.005 $Y2=0.402
r518 162 166 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.335 $Y=0.34
+ $X2=2.005 $Y2=0.34
r519 160 162 7.32169 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.2 $Y=0.4
+ $X2=1.335 $Y2=0.4
r520 160 161 7.32169 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.2 $Y=0.4
+ $X2=1.065 $Y2=0.4
r521 156 226 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=0.245 $Y=2.295
+ $X2=0.245 $Y2=1.66
r522 156 158 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=2.295
+ $X2=0.245 $Y2=2.38
r523 153 192 3.26526 $w=2.98e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=0.425
+ $X2=0.245 $Y2=0.51
r524 153 155 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=0.425
+ $X2=0.245 $Y2=0.34
r525 151 218 7.88011 $w=3.67e-07 $l=6e-08 $layer=POLY_cond $X=14.66 $Y=1.202
+ $X2=14.72 $Y2=1.202
r526 151 216 47.2807 $w=3.67e-07 $l=3.6e-07 $layer=POLY_cond $X=14.66 $Y=1.202
+ $X2=14.3 $Y2=1.202
r527 150 151 22.3508 $w=1.7e-07 $l=1.105e-06 $layer=licon1_POLY $count=6
+ $X=14.66 $Y=1.16 $X2=14.66 $Y2=1.16
r528 148 201 49.9074 $w=3.67e-07 $l=3.8e-07 $layer=POLY_cond $X=10.58 $Y=1.202
+ $X2=10.96 $Y2=1.202
r529 148 199 5.25341 $w=3.67e-07 $l=4e-08 $layer=POLY_cond $X=10.58 $Y=1.202
+ $X2=10.54 $Y2=1.202
r530 147 150 188.079 $w=2.48e-07 $l=4.08e-06 $layer=LI1_cond $X=10.58 $Y=1.2
+ $X2=14.66 $Y2=1.2
r531 147 148 22.3508 $w=1.7e-07 $l=1.105e-06 $layer=licon1_POLY $count=6
+ $X=10.58 $Y=1.16 $X2=10.58 $Y2=1.16
r532 145 185 2.0066 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=9.925 $Y=1.2
+ $X2=9.775 $Y2=1.2
r533 145 147 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=9.925 $Y=1.2
+ $X2=10.58 $Y2=1.2
r534 142 187 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.775 $Y=2.295
+ $X2=9.775 $Y2=2.38
r535 142 144 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=9.775 $Y=2.295
+ $X2=9.775 $Y2=1.66
r536 141 185 4.4274 $w=3e-07 $l=1.25e-07 $layer=LI1_cond $X=9.775 $Y=1.325
+ $X2=9.775 $Y2=1.2
r537 141 144 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=9.775 $Y=1.325
+ $X2=9.775 $Y2=1.66
r538 140 180 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.955 $Y=2.38
+ $X2=8.82 $Y2=2.38
r539 139 187 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=9.625 $Y=2.38
+ $X2=9.775 $Y2=2.38
r540 139 140 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.625 $Y=2.38
+ $X2=8.955 $Y2=2.38
r541 137 183 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=9.625 $Y=0.34
+ $X2=9.775 $Y2=0.34
r542 137 179 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.625 $Y=0.34
+ $X2=8.955 $Y2=0.34
r543 133 180 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.82 $Y=2.295
+ $X2=8.82 $Y2=2.38
r544 133 135 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.82 $Y=2.295
+ $X2=8.82 $Y2=2
r545 132 175 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=8.015 $Y=2.38
+ $X2=7.865 $Y2=2.38
r546 131 180 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.685 $Y=2.38
+ $X2=8.82 $Y2=2.38
r547 131 132 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.685 $Y=2.38
+ $X2=8.015 $Y2=2.38
r548 125 175 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.865 $Y=2.295
+ $X2=7.865 $Y2=2.38
r549 125 127 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=7.865 $Y=2.295
+ $X2=7.865 $Y2=1.66
r550 121 169 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=2.295
+ $X2=2.155 $Y2=2.38
r551 121 123 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=2.155 $Y=2.295
+ $X2=2.155 $Y2=1.66
r552 120 163 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=2.38
+ $X2=1.2 $Y2=2.38
r553 119 169 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.005 $Y=2.38
+ $X2=2.155 $Y2=2.38
r554 119 120 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=2.38
+ $X2=1.335 $Y2=2.38
r555 113 163 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.295
+ $X2=1.2 $Y2=2.38
r556 113 115 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=2.295
+ $X2=1.2 $Y2=2
r557 112 158 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.395 $Y=2.38
+ $X2=0.245 $Y2=2.38
r558 111 163 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=2.38
+ $X2=1.2 $Y2=2.38
r559 111 112 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.065 $Y=2.38
+ $X2=0.395 $Y2=2.38
r560 110 155 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.395 $Y=0.34
+ $X2=0.245 $Y2=0.34
r561 110 161 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.395 $Y=0.34
+ $X2=1.065 $Y2=0.34
r562 106 223 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=15.685 $Y=1.41
+ $X2=15.685 $Y2=1.202
r563 106 108 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.685 $Y=1.41
+ $X2=15.685 $Y2=1.985
r564 103 222 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=15.66 $Y=0.995
+ $X2=15.66 $Y2=1.202
r565 103 105 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=15.66 $Y=0.995
+ $X2=15.66 $Y2=0.56
r566 100 221 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=15.24 $Y=0.995
+ $X2=15.24 $Y2=1.202
r567 100 102 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=15.24 $Y=0.995
+ $X2=15.24 $Y2=0.56
r568 97 220 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=15.215 $Y=1.41
+ $X2=15.215 $Y2=1.202
r569 97 99 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.215 $Y=1.41
+ $X2=15.215 $Y2=1.985
r570 94 219 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=14.745 $Y=1.41
+ $X2=14.745 $Y2=1.202
r571 94 96 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=14.745 $Y=1.41
+ $X2=14.745 $Y2=1.985
r572 91 218 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=14.72 $Y=0.995
+ $X2=14.72 $Y2=1.202
r573 91 93 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=14.72 $Y=0.995
+ $X2=14.72 $Y2=0.56
r574 88 216 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=14.3 $Y=0.995
+ $X2=14.3 $Y2=1.202
r575 88 90 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=14.3 $Y=0.995
+ $X2=14.3 $Y2=0.56
r576 85 215 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=14.275 $Y=1.41
+ $X2=14.275 $Y2=1.202
r577 85 87 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=14.275 $Y=1.41
+ $X2=14.275 $Y2=1.985
r578 82 214 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=13.805 $Y=1.41
+ $X2=13.805 $Y2=1.202
r579 82 84 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=13.805 $Y=1.41
+ $X2=13.805 $Y2=1.985
r580 79 213 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=13.78 $Y=0.995
+ $X2=13.78 $Y2=1.202
r581 79 81 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.78 $Y=0.995
+ $X2=13.78 $Y2=0.56
r582 76 212 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=13.36 $Y=0.995
+ $X2=13.36 $Y2=1.202
r583 76 78 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.36 $Y=0.995
+ $X2=13.36 $Y2=0.56
r584 73 211 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=13.335 $Y=1.41
+ $X2=13.335 $Y2=1.202
r585 73 75 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=13.335 $Y=1.41
+ $X2=13.335 $Y2=1.985
r586 70 210 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=12.865 $Y=1.41
+ $X2=12.865 $Y2=1.202
r587 70 72 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.865 $Y=1.41
+ $X2=12.865 $Y2=1.985
r588 67 209 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=12.84 $Y=0.995
+ $X2=12.84 $Y2=1.202
r589 67 69 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.84 $Y=0.995
+ $X2=12.84 $Y2=0.56
r590 64 208 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=12.42 $Y=0.995
+ $X2=12.42 $Y2=1.202
r591 64 66 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.42 $Y=0.995
+ $X2=12.42 $Y2=0.56
r592 61 207 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=12.395 $Y=1.41
+ $X2=12.395 $Y2=1.202
r593 61 63 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.395 $Y=1.41
+ $X2=12.395 $Y2=1.985
r594 58 206 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=11.925 $Y=1.41
+ $X2=11.925 $Y2=1.202
r595 58 60 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.925 $Y=1.41
+ $X2=11.925 $Y2=1.985
r596 55 205 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.9 $Y=0.995
+ $X2=11.9 $Y2=1.202
r597 55 57 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.9 $Y=0.995
+ $X2=11.9 $Y2=0.56
r598 52 204 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.48 $Y=0.995
+ $X2=11.48 $Y2=1.202
r599 52 54 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.48 $Y=0.995
+ $X2=11.48 $Y2=0.56
r600 49 203 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=11.455 $Y=1.41
+ $X2=11.455 $Y2=1.202
r601 49 51 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.455 $Y=1.41
+ $X2=11.455 $Y2=1.985
r602 46 202 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.985 $Y=1.41
+ $X2=10.985 $Y2=1.202
r603 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.985 $Y=1.41
+ $X2=10.985 $Y2=1.985
r604 43 201 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.96 $Y=0.995
+ $X2=10.96 $Y2=1.202
r605 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.96 $Y=0.995
+ $X2=10.96 $Y2=0.56
r606 40 199 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.54 $Y=0.995
+ $X2=10.54 $Y2=1.202
r607 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.54 $Y=0.995
+ $X2=10.54 $Y2=0.56
r608 37 198 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.515 $Y=1.41
+ $X2=10.515 $Y2=1.202
r609 37 39 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.515 $Y=1.41
+ $X2=10.515 $Y2=1.985
r610 12 187 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=9.615
+ $Y=1.485 $X2=9.76 $Y2=2.34
r611 12 144 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=9.615
+ $Y=1.485 $X2=9.76 $Y2=1.66
r612 11 135 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=8.675
+ $Y=1.485 $X2=8.82 $Y2=2
r613 10 175 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=7.755
+ $Y=1.485 $X2=7.88 $Y2=2.34
r614 10 127 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=7.755
+ $Y=1.485 $X2=7.88 $Y2=1.66
r615 9 169 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2.34
r616 9 123 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.66
r617 8 115 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r618 7 226 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r619 7 158 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r620 6 183 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=9.575
+ $Y=0.235 $X2=9.76 $Y2=0.4
r621 5 177 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=8.635
+ $Y=0.235 $X2=8.82 $Y2=0.38
r622 4 171 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=7.755
+ $Y=0.235 $X2=7.88 $Y2=0.385
r623 3 165 182 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.235 $X2=2.14 $Y2=0.385
r624 2 160 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.38
r625 1 155 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_12%A_117_297# 1 2 3 4 13 15 17 20 23 26 29 30
+ 31 32 33 34 37 41 44 46 47
r131 47 59 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=6.89 $Y=1.87
+ $X2=6.89 $Y2=2.34
r132 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.89 $Y=1.87
+ $X2=6.89 $Y2=1.87
r133 44 55 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=5.95 $Y=1.87
+ $X2=5.95 $Y2=2.34
r134 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.95 $Y=1.87
+ $X2=5.95 $Y2=1.87
r135 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.67 $Y=1.87
+ $X2=1.67 $Y2=1.87
r136 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.73 $Y=1.87
+ $X2=0.73 $Y2=1.87
r137 34 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.095 $Y=1.87
+ $X2=5.95 $Y2=1.87
r138 33 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.745 $Y=1.87
+ $X2=6.89 $Y2=1.87
r139 33 34 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=6.745 $Y=1.87
+ $X2=6.095 $Y2=1.87
r140 32 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.815 $Y=1.87
+ $X2=1.67 $Y2=1.87
r141 31 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.805 $Y=1.87
+ $X2=5.95 $Y2=1.87
r142 31 32 4.93811 $w=1.4e-07 $l=3.99e-06 $layer=MET1_cond $X=5.805 $Y=1.87
+ $X2=1.815 $Y2=1.87
r143 30 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.875 $Y=1.87
+ $X2=0.73 $Y2=1.87
r144 29 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.525 $Y=1.87
+ $X2=1.67 $Y2=1.87
r145 29 30 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=1.525 $Y=1.87
+ $X2=0.875 $Y2=1.87
r146 26 47 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=6.89 $Y=1.665
+ $X2=6.89 $Y2=1.87
r147 26 28 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=1.665
+ $X2=6.89 $Y2=1.58
r148 23 44 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=5.95 $Y=1.665
+ $X2=5.95 $Y2=1.87
r149 23 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=1.665
+ $X2=5.95 $Y2=1.58
r150 20 41 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=1.87
r151 20 22 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=1.58
r152 17 37 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=1.87
r153 17 19 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=1.58
r154 16 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.115 $Y=1.58
+ $X2=5.95 $Y2=1.58
r155 15 28 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.725 $Y=1.58
+ $X2=6.89 $Y2=1.58
r156 15 16 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.725 $Y=1.58
+ $X2=6.115 $Y2=1.58
r157 14 19 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.73 $Y2=1.58
r158 13 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=1.67 $Y2=1.58
r159 13 14 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=0.895 $Y2=1.58
r160 4 59 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=2.34
r161 4 28 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=1.66
r162 3 55 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=2.34
r163 3 25 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=1.66
r164 2 22 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r165 1 19 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_12%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 42 48
+ 52 58 64 68 74 80 84 88 92 96 100 105 106 108 109 111 112 114 115 117 118 120
+ 121 122 124 151 155 160 165 170 175 182 183 186 189 192 195 198 201 204 208
c273 108 0 1.97192e-19 $X=4.405 $Y=2.72
c274 105 0 1.97192e-19 $X=3.465 $Y=2.72
c275 5 0 1.91318e-19 $X=6.275 $Y=1.485
c276 2 0 1.91318e-19 $X=3.455 $Y=1.485
r277 204 205 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.87 $Y=2.72
+ $X2=15.87 $Y2=2.72
r278 201 202 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.95 $Y=2.72
+ $X2=14.95 $Y2=2.72
r279 198 199 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=2.72
+ $X2=14.03 $Y2=2.72
r280 195 196 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r281 192 193 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r282 189 190 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r283 186 187 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r284 183 205 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=16.33 $Y=2.72
+ $X2=15.87 $Y2=2.72
r285 182 183 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.33 $Y=2.72
+ $X2=16.33 $Y2=2.72
r286 180 204 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=16.055 $Y=2.72
+ $X2=15.92 $Y2=2.72
r287 180 182 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=16.055 $Y=2.72
+ $X2=16.33 $Y2=2.72
r288 179 205 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.41 $Y=2.72
+ $X2=15.87 $Y2=2.72
r289 179 202 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.41 $Y=2.72
+ $X2=14.95 $Y2=2.72
r290 178 179 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.41 $Y=2.72
+ $X2=15.41 $Y2=2.72
r291 176 201 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=15.115 $Y=2.72
+ $X2=14.98 $Y2=2.72
r292 176 178 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=15.115 $Y=2.72
+ $X2=15.41 $Y2=2.72
r293 175 204 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=15.785 $Y=2.72
+ $X2=15.92 $Y2=2.72
r294 175 178 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=15.785 $Y=2.72
+ $X2=15.41 $Y2=2.72
r295 174 202 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=2.72
+ $X2=14.95 $Y2=2.72
r296 174 199 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=2.72
+ $X2=14.03 $Y2=2.72
r297 173 174 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.49 $Y=2.72
+ $X2=14.49 $Y2=2.72
r298 171 198 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.175 $Y=2.72
+ $X2=14.04 $Y2=2.72
r299 171 173 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=14.175 $Y=2.72
+ $X2=14.49 $Y2=2.72
r300 170 201 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.845 $Y=2.72
+ $X2=14.98 $Y2=2.72
r301 170 173 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=14.845 $Y=2.72
+ $X2=14.49 $Y2=2.72
r302 169 199 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=2.72
+ $X2=14.03 $Y2=2.72
r303 169 196 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=2.72
+ $X2=13.11 $Y2=2.72
r304 168 169 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=2.72
+ $X2=13.57 $Y2=2.72
r305 166 195 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.235 $Y=2.72
+ $X2=13.1 $Y2=2.72
r306 166 168 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.235 $Y=2.72
+ $X2=13.57 $Y2=2.72
r307 165 198 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.905 $Y=2.72
+ $X2=14.04 $Y2=2.72
r308 165 168 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.905 $Y=2.72
+ $X2=13.57 $Y2=2.72
r309 164 196 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=13.11 $Y2=2.72
r310 164 193 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=12.19 $Y2=2.72
r311 163 164 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r312 161 192 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.295 $Y=2.72
+ $X2=12.16 $Y2=2.72
r313 161 163 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=12.295 $Y=2.72
+ $X2=12.65 $Y2=2.72
r314 160 195 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.965 $Y=2.72
+ $X2=13.1 $Y2=2.72
r315 160 163 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.965 $Y=2.72
+ $X2=12.65 $Y2=2.72
r316 159 193 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=12.19 $Y2=2.72
r317 159 190 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=11.27 $Y2=2.72
r318 158 159 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r319 156 189 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.355 $Y=2.72
+ $X2=11.22 $Y2=2.72
r320 156 158 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.355 $Y=2.72
+ $X2=11.73 $Y2=2.72
r321 155 192 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.025 $Y=2.72
+ $X2=12.16 $Y2=2.72
r322 155 158 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.025 $Y=2.72
+ $X2=11.73 $Y2=2.72
r323 154 190 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.27 $Y2=2.72
r324 153 154 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r325 151 189 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.085 $Y=2.72
+ $X2=11.22 $Y2=2.72
r326 151 153 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.085 $Y=2.72
+ $X2=10.81 $Y2=2.72
r327 150 154 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.81 $Y2=2.72
r328 149 150 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r329 147 150 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=9.89 $Y2=2.72
r330 146 149 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=7.59 $Y=2.72
+ $X2=9.89 $Y2=2.72
r331 146 147 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r332 144 147 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r333 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r334 141 144 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r335 140 141 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r336 138 141 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r337 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r338 135 138 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r339 134 135 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r340 132 135 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r341 132 187 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r342 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r343 129 186 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=2.66 $Y2=2.72
r344 129 131 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=3.45 $Y2=2.72
r345 126 208 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r346 124 186 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.66 $Y2=2.72
r347 124 126 149.727 $w=1.68e-07 $l=2.295e-06 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=0.23 $Y2=2.72
r348 122 187 0.653023 $w=4.8e-07 $l=2.295e-06 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=2.53 $Y2=2.72
r349 122 208 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r350 120 149 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=10.145 $Y=2.72
+ $X2=9.89 $Y2=2.72
r351 120 121 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.145 $Y=2.72
+ $X2=10.28 $Y2=2.72
r352 119 153 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.415 $Y=2.72
+ $X2=10.81 $Y2=2.72
r353 119 121 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.415 $Y=2.72
+ $X2=10.28 $Y2=2.72
r354 117 143 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.225 $Y=2.72
+ $X2=7.13 $Y2=2.72
r355 117 118 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.225 $Y=2.72
+ $X2=7.36 $Y2=2.72
r356 116 146 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.495 $Y=2.72
+ $X2=7.59 $Y2=2.72
r357 116 118 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.495 $Y=2.72
+ $X2=7.36 $Y2=2.72
r358 114 140 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.285 $Y=2.72
+ $X2=6.21 $Y2=2.72
r359 114 115 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.285 $Y=2.72
+ $X2=6.42 $Y2=2.72
r360 113 143 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.555 $Y=2.72
+ $X2=7.13 $Y2=2.72
r361 113 115 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.555 $Y=2.72
+ $X2=6.42 $Y2=2.72
r362 111 137 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=5.345 $Y=2.72
+ $X2=5.29 $Y2=2.72
r363 111 112 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.345 $Y=2.72
+ $X2=5.48 $Y2=2.72
r364 110 140 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.615 $Y=2.72
+ $X2=6.21 $Y2=2.72
r365 110 112 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.615 $Y=2.72
+ $X2=5.48 $Y2=2.72
r366 108 134 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.405 $Y=2.72
+ $X2=4.37 $Y2=2.72
r367 108 109 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.405 $Y=2.72
+ $X2=4.54 $Y2=2.72
r368 107 137 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.675 $Y=2.72
+ $X2=5.29 $Y2=2.72
r369 107 109 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.675 $Y=2.72
+ $X2=4.54 $Y2=2.72
r370 105 131 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.465 $Y=2.72
+ $X2=3.45 $Y2=2.72
r371 105 106 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.465 $Y=2.72
+ $X2=3.6 $Y2=2.72
r372 104 134 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.735 $Y=2.72
+ $X2=4.37 $Y2=2.72
r373 104 106 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.735 $Y=2.72
+ $X2=3.6 $Y2=2.72
r374 100 103 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=15.92 $Y=1.66
+ $X2=15.92 $Y2=2.34
r375 98 204 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.92 $Y=2.635
+ $X2=15.92 $Y2=2.72
r376 98 103 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=15.92 $Y=2.635
+ $X2=15.92 $Y2=2.34
r377 94 201 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.98 $Y=2.635
+ $X2=14.98 $Y2=2.72
r378 94 96 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=14.98 $Y=2.635
+ $X2=14.98 $Y2=2
r379 90 198 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.04 $Y=2.635
+ $X2=14.04 $Y2=2.72
r380 90 92 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=14.04 $Y=2.635
+ $X2=14.04 $Y2=2
r381 86 195 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.1 $Y=2.635
+ $X2=13.1 $Y2=2.72
r382 86 88 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=13.1 $Y=2.635
+ $X2=13.1 $Y2=2
r383 82 192 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.16 $Y=2.635
+ $X2=12.16 $Y2=2.72
r384 82 84 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=12.16 $Y=2.635
+ $X2=12.16 $Y2=2
r385 78 189 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.22 $Y=2.635
+ $X2=11.22 $Y2=2.72
r386 78 80 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=11.22 $Y=2.635
+ $X2=11.22 $Y2=2
r387 74 77 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=10.28 $Y=1.66
+ $X2=10.28 $Y2=2.34
r388 72 121 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.28 $Y=2.635
+ $X2=10.28 $Y2=2.72
r389 72 77 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.28 $Y=2.635
+ $X2=10.28 $Y2=2.34
r390 68 71 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.36 $Y=1.66
+ $X2=7.36 $Y2=2.34
r391 66 118 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=2.635
+ $X2=7.36 $Y2=2.72
r392 66 71 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.36 $Y=2.635
+ $X2=7.36 $Y2=2.34
r393 62 115 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=2.72
r394 62 64 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=2
r395 58 61 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.48 $Y=1.66
+ $X2=5.48 $Y2=2.34
r396 56 112 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2.72
r397 56 61 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2.34
r398 52 55 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.54 $Y=1.66
+ $X2=4.54 $Y2=2.34
r399 50 109 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=2.635
+ $X2=4.54 $Y2=2.72
r400 50 55 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.54 $Y=2.635
+ $X2=4.54 $Y2=2.34
r401 46 106 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=2.635
+ $X2=3.6 $Y2=2.72
r402 46 48 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.6 $Y=2.635
+ $X2=3.6 $Y2=2
r403 42 45 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.66 $Y=1.66
+ $X2=2.66 $Y2=2.34
r404 40 186 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=2.635
+ $X2=2.66 $Y2=2.72
r405 40 45 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.66 $Y=2.635
+ $X2=2.66 $Y2=2.34
r406 13 103 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=15.775
+ $Y=1.485 $X2=15.92 $Y2=2.34
r407 13 100 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=15.775
+ $Y=1.485 $X2=15.92 $Y2=1.66
r408 12 96 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=14.835
+ $Y=1.485 $X2=14.98 $Y2=2
r409 11 92 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=13.895
+ $Y=1.485 $X2=14.04 $Y2=2
r410 10 88 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=12.955
+ $Y=1.485 $X2=13.1 $Y2=2
r411 9 84 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=12.015
+ $Y=1.485 $X2=12.16 $Y2=2
r412 8 80 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=11.075
+ $Y=1.485 $X2=11.22 $Y2=2
r413 7 77 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=10.155
+ $Y=1.485 $X2=10.28 $Y2=2.34
r414 7 74 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=10.155
+ $Y=1.485 $X2=10.28 $Y2=1.66
r415 6 71 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.215
+ $Y=1.485 $X2=7.36 $Y2=2.34
r416 6 68 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=7.215
+ $Y=1.485 $X2=7.36 $Y2=1.66
r417 5 64 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.275
+ $Y=1.485 $X2=6.42 $Y2=2
r418 4 61 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=2.34
r419 4 58 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=1.66
r420 3 55 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.485 $X2=4.54 $Y2=2.34
r421 3 52 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.485 $X2=4.54 $Y2=1.66
r422 2 48 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.455
+ $Y=1.485 $X2=3.6 $Y2=2
r423 1 45 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.535
+ $Y=1.485 $X2=2.66 $Y2=2.34
r424 1 42 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=2.535
+ $Y=1.485 $X2=2.66 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_12%A_597_297# 1 2 3 4 13 15 17 20 23 26 29 30
+ 31 32 34 35 36 37 38 41 45 48 50 51
c138 32 0 1.97192e-19 $X=4.215 $Y=2.21
c139 31 0 1.91318e-19 $X=7.52 $Y=2.21
c140 30 0 1.97192e-19 $X=3.275 $Y=2.21
c141 29 0 1.91318e-19 $X=3.925 $Y=2.21
r142 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.29 $Y=1.87
+ $X2=9.29 $Y2=1.87
r143 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.35 $Y=1.87
+ $X2=8.35 $Y2=1.87
r144 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.07 $Y=2.21
+ $X2=4.07 $Y2=2.21
r145 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.13 $Y=2.21
+ $X2=3.13 $Y2=2.21
r146 38 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.495 $Y=1.87
+ $X2=8.35 $Y2=1.87
r147 37 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.145 $Y=1.87
+ $X2=9.29 $Y2=1.87
r148 37 38 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=9.145 $Y=1.87
+ $X2=8.495 $Y2=1.87
r149 35 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.205 $Y=1.87
+ $X2=8.35 $Y2=1.87
r150 35 36 0.674504 $w=1.4e-07 $l=5.45e-07 $layer=MET1_cond $X=8.205 $Y=1.87
+ $X2=7.66 $Y2=1.87
r151 33 36 0.0698411 $w=1.4e-07 $l=9.89949e-08 $layer=MET1_cond $X=7.59 $Y=1.94
+ $X2=7.66 $Y2=1.87
r152 33 34 0.247524 $w=1.4e-07 $l=2e-07 $layer=MET1_cond $X=7.59 $Y=1.94
+ $X2=7.59 $Y2=2.14
r153 32 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.215 $Y=2.21
+ $X2=4.07 $Y2=2.21
r154 31 34 0.0698411 $w=1.4e-07 $l=9.89949e-08 $layer=MET1_cond $X=7.52 $Y=2.21
+ $X2=7.59 $Y2=2.14
r155 31 32 4.09034 $w=1.4e-07 $l=3.305e-06 $layer=MET1_cond $X=7.52 $Y=2.21
+ $X2=4.215 $Y2=2.21
r156 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.275 $Y=2.21
+ $X2=3.13 $Y2=2.21
r157 29 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.925 $Y=2.21
+ $X2=4.07 $Y2=2.21
r158 29 30 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=3.925 $Y=2.21
+ $X2=3.275 $Y2=2.21
r159 26 51 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=9.29 $Y=1.665
+ $X2=9.29 $Y2=1.87
r160 26 28 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.29 $Y=1.665
+ $X2=9.29 $Y2=1.58
r161 23 48 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=8.35 $Y=1.665
+ $X2=8.35 $Y2=1.87
r162 23 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.35 $Y=1.665
+ $X2=8.35 $Y2=1.58
r163 20 45 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=4.07 $Y=1.665
+ $X2=4.07 $Y2=2.21
r164 20 22 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=1.665
+ $X2=4.07 $Y2=1.58
r165 17 41 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=3.13 $Y=1.665
+ $X2=3.13 $Y2=2.21
r166 17 19 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=1.665
+ $X2=3.13 $Y2=1.58
r167 16 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.515 $Y=1.58
+ $X2=8.35 $Y2=1.58
r168 15 28 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.125 $Y=1.58
+ $X2=9.29 $Y2=1.58
r169 15 16 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=9.125 $Y=1.58
+ $X2=8.515 $Y2=1.58
r170 14 19 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=1.58
+ $X2=3.13 $Y2=1.58
r171 13 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.905 $Y=1.58
+ $X2=4.07 $Y2=1.58
r172 13 14 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.905 $Y=1.58
+ $X2=3.295 $Y2=1.58
r173 4 28 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=9.145
+ $Y=1.485 $X2=9.29 $Y2=1.66
r174 3 25 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=8.205
+ $Y=1.485 $X2=8.35 $Y2=1.66
r175 2 45 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=2.34
r176 2 22 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=1.66
r177 1 41 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.985
+ $Y=1.485 $X2=3.13 $Y2=2.34
r178 1 19 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.985
+ $Y=1.485 $X2=3.13 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_12%X 1 2 3 4 5 6 7 8 9 10 11 12 39 41 43 45
+ 46 47 51 55 57 59 63 67 69 71 75 79 81 83 87 91 93 95 99 103 107 109 110 112
+ 113 115 116 118 120 123 124
r219 121 124 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=15.45 $Y=1.495
+ $X2=15.45 $Y2=1.19
r220 121 123 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.45 $Y=1.495
+ $X2=15.45 $Y2=1.58
r221 119 124 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=15.45 $Y=0.905
+ $X2=15.45 $Y2=1.19
r222 119 120 3.0419 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=15.45 $Y=0.905
+ $X2=15.45 $Y2=0.815
r223 101 123 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.45 $Y=1.665
+ $X2=15.45 $Y2=1.58
r224 101 103 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=15.45 $Y=1.665
+ $X2=15.45 $Y2=2.34
r225 97 120 3.0419 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=15.45 $Y=0.725
+ $X2=15.45 $Y2=0.815
r226 97 99 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=15.45 $Y=0.725
+ $X2=15.45 $Y2=0.42
r227 96 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.675 $Y=1.58
+ $X2=14.51 $Y2=1.58
r228 95 123 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.285 $Y=1.58
+ $X2=15.45 $Y2=1.58
r229 95 96 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=15.285 $Y=1.58
+ $X2=14.675 $Y2=1.58
r230 94 116 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=14.675 $Y=0.815
+ $X2=14.51 $Y2=0.815
r231 93 120 3.59259 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=15.285 $Y=0.815
+ $X2=15.45 $Y2=0.815
r232 93 94 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=15.285 $Y=0.815
+ $X2=14.675 $Y2=0.815
r233 89 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.51 $Y=1.665
+ $X2=14.51 $Y2=1.58
r234 89 91 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=14.51 $Y=1.665
+ $X2=14.51 $Y2=2.34
r235 85 116 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=14.51 $Y=0.725
+ $X2=14.51 $Y2=0.815
r236 85 87 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=14.51 $Y=0.725
+ $X2=14.51 $Y2=0.42
r237 84 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.735 $Y=1.58
+ $X2=13.57 $Y2=1.58
r238 83 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.345 $Y=1.58
+ $X2=14.51 $Y2=1.58
r239 83 84 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=14.345 $Y=1.58
+ $X2=13.735 $Y2=1.58
r240 82 113 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=13.735 $Y=0.815
+ $X2=13.57 $Y2=0.815
r241 81 116 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=14.345 $Y=0.815
+ $X2=14.51 $Y2=0.815
r242 81 82 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=14.345 $Y=0.815
+ $X2=13.735 $Y2=0.815
r243 77 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.57 $Y=1.665
+ $X2=13.57 $Y2=1.58
r244 77 79 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=13.57 $Y=1.665
+ $X2=13.57 $Y2=2.34
r245 73 113 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=13.57 $Y=0.725
+ $X2=13.57 $Y2=0.815
r246 73 75 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=13.57 $Y=0.725
+ $X2=13.57 $Y2=0.42
r247 72 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.795 $Y=1.58
+ $X2=12.63 $Y2=1.58
r248 71 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.405 $Y=1.58
+ $X2=13.57 $Y2=1.58
r249 71 72 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=13.405 $Y=1.58
+ $X2=12.795 $Y2=1.58
r250 70 110 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=12.795 $Y=0.815
+ $X2=12.63 $Y2=0.815
r251 69 113 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=13.405 $Y=0.815
+ $X2=13.57 $Y2=0.815
r252 69 70 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=13.405 $Y=0.815
+ $X2=12.795 $Y2=0.815
r253 65 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.63 $Y=1.665
+ $X2=12.63 $Y2=1.58
r254 65 67 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=12.63 $Y=1.665
+ $X2=12.63 $Y2=2.34
r255 61 110 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=12.63 $Y=0.725
+ $X2=12.63 $Y2=0.815
r256 61 63 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=12.63 $Y=0.725
+ $X2=12.63 $Y2=0.42
r257 60 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.855 $Y=1.58
+ $X2=11.69 $Y2=1.58
r258 59 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.465 $Y=1.58
+ $X2=12.63 $Y2=1.58
r259 59 60 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=12.465 $Y=1.58
+ $X2=11.855 $Y2=1.58
r260 58 107 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=11.855 $Y=0.815
+ $X2=11.69 $Y2=0.815
r261 57 110 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=12.465 $Y=0.815
+ $X2=12.63 $Y2=0.815
r262 57 58 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=12.465 $Y=0.815
+ $X2=11.855 $Y2=0.815
r263 53 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.69 $Y=1.665
+ $X2=11.69 $Y2=1.58
r264 53 55 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=11.69 $Y=1.665
+ $X2=11.69 $Y2=2.34
r265 49 107 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=11.69 $Y=0.725
+ $X2=11.69 $Y2=0.815
r266 49 51 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=11.69 $Y=0.725
+ $X2=11.69 $Y2=0.42
r267 48 106 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.915 $Y=1.58
+ $X2=10.75 $Y2=1.58
r268 47 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.525 $Y=1.58
+ $X2=11.69 $Y2=1.58
r269 47 48 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=11.525 $Y=1.58
+ $X2=10.915 $Y2=1.58
r270 45 107 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=11.525 $Y=0.815
+ $X2=11.69 $Y2=0.815
r271 45 46 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=11.525 $Y=0.815
+ $X2=10.915 $Y2=0.815
r272 41 106 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.75 $Y=1.665
+ $X2=10.75 $Y2=1.58
r273 41 43 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=10.75 $Y=1.665
+ $X2=10.75 $Y2=2.34
r274 37 46 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=10.75 $Y=0.725
+ $X2=10.915 $Y2=0.815
r275 37 39 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=10.75 $Y=0.725
+ $X2=10.75 $Y2=0.42
r276 12 123 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=15.305
+ $Y=1.485 $X2=15.45 $Y2=1.66
r277 12 103 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=15.305
+ $Y=1.485 $X2=15.45 $Y2=2.34
r278 11 118 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=14.365
+ $Y=1.485 $X2=14.51 $Y2=1.66
r279 11 91 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=14.365
+ $Y=1.485 $X2=14.51 $Y2=2.34
r280 10 115 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=13.425
+ $Y=1.485 $X2=13.57 $Y2=1.66
r281 10 79 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=13.425
+ $Y=1.485 $X2=13.57 $Y2=2.34
r282 9 112 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=12.485
+ $Y=1.485 $X2=12.63 $Y2=1.66
r283 9 67 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=12.485
+ $Y=1.485 $X2=12.63 $Y2=2.34
r284 8 109 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=11.545
+ $Y=1.485 $X2=11.69 $Y2=1.66
r285 8 55 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=11.545
+ $Y=1.485 $X2=11.69 $Y2=2.34
r286 7 106 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=10.605
+ $Y=1.485 $X2=10.75 $Y2=1.66
r287 7 43 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.605
+ $Y=1.485 $X2=10.75 $Y2=2.34
r288 6 99 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=15.315
+ $Y=0.235 $X2=15.45 $Y2=0.42
r289 5 87 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=14.375
+ $Y=0.235 $X2=14.51 $Y2=0.42
r290 4 75 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=13.435
+ $Y=0.235 $X2=13.57 $Y2=0.42
r291 3 63 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=12.495
+ $Y=0.235 $X2=12.63 $Y2=0.42
r292 2 51 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=11.555
+ $Y=0.235 $X2=11.69 $Y2=0.42
r293 1 39 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=10.615
+ $Y=0.235 $X2=10.75 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_12%A_119_47# 1 2 3 4 15 19 21 25 30 33 34 35
r83 32 34 8.14364 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.67 $Y=0.75
+ $X2=1.835 $Y2=0.75
r84 32 33 8.14364 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.67 $Y=0.75
+ $X2=1.505 $Y2=0.75
r85 30 33 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=0.895 $Y=0.815
+ $X2=1.505 $Y2=0.815
r86 28 30 8.14364 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=0.75
+ $X2=0.895 $Y2=0.75
r87 23 25 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.07 $Y=0.725
+ $X2=4.07 $Y2=0.42
r88 22 35 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=0.815
+ $X2=3.13 $Y2=0.815
r89 21 23 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=3.905 $Y=0.815
+ $X2=4.07 $Y2=0.725
r90 21 22 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=3.905 $Y=0.815
+ $X2=3.295 $Y2=0.815
r91 17 35 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.13 $Y=0.725 $X2=3.13
+ $Y2=0.815
r92 17 19 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=3.13 $Y=0.725
+ $X2=3.13 $Y2=0.42
r93 15 35 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=0.815
+ $X2=3.13 $Y2=0.815
r94 15 34 69.6263 $w=1.78e-07 $l=1.13e-06 $layer=LI1_cond $X=2.965 $Y=0.815
+ $X2=1.835 $Y2=0.815
r95 4 25 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=3.935
+ $Y=0.235 $X2=4.07 $Y2=0.42
r96 3 19 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=2.995
+ $Y=0.235 $X2=3.13 $Y2=0.42
r97 2 32 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.76
r98 1 28 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_12%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 42 46
+ 50 54 58 62 66 70 74 78 82 86 90 93 94 96 97 99 100 102 103 105 106 108 109
+ 110 112 139 143 148 153 158 163 170 171 174 177 180 183 186 189 192 196
c264 112 0 1.96891e-19 $X=2.525 $Y=0
c265 108 0 1.96891e-19 $X=10.145 $Y=0
r266 192 193 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.87 $Y=0
+ $X2=15.87 $Y2=0
r267 189 190 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.95 $Y=0
+ $X2=14.95 $Y2=0
r268 186 187 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=0
+ $X2=14.03 $Y2=0
r269 183 184 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r270 180 181 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r271 177 178 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r272 174 175 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r273 171 193 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=16.33 $Y=0
+ $X2=15.87 $Y2=0
r274 170 171 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.33 $Y=0
+ $X2=16.33 $Y2=0
r275 168 192 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=16.055 $Y=0
+ $X2=15.92 $Y2=0
r276 168 170 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=16.055 $Y=0
+ $X2=16.33 $Y2=0
r277 167 193 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.41 $Y=0
+ $X2=15.87 $Y2=0
r278 167 190 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.41 $Y=0
+ $X2=14.95 $Y2=0
r279 166 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.41 $Y=0
+ $X2=15.41 $Y2=0
r280 164 189 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=15.115 $Y=0
+ $X2=14.98 $Y2=0
r281 164 166 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=15.115 $Y=0
+ $X2=15.41 $Y2=0
r282 163 192 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=15.785 $Y=0
+ $X2=15.92 $Y2=0
r283 163 166 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=15.785 $Y=0
+ $X2=15.41 $Y2=0
r284 162 190 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=0
+ $X2=14.95 $Y2=0
r285 162 187 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=0
+ $X2=14.03 $Y2=0
r286 161 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.49 $Y=0
+ $X2=14.49 $Y2=0
r287 159 186 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.175 $Y=0
+ $X2=14.04 $Y2=0
r288 159 161 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=14.175 $Y=0
+ $X2=14.49 $Y2=0
r289 158 189 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.845 $Y=0
+ $X2=14.98 $Y2=0
r290 158 161 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=14.845 $Y=0
+ $X2=14.49 $Y2=0
r291 157 187 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=14.03 $Y2=0
r292 157 184 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=13.11 $Y2=0
r293 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r294 154 183 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.235 $Y=0
+ $X2=13.1 $Y2=0
r295 154 156 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.235 $Y=0
+ $X2=13.57 $Y2=0
r296 153 186 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.905 $Y=0
+ $X2=14.04 $Y2=0
r297 153 156 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.905 $Y=0
+ $X2=13.57 $Y2=0
r298 152 184 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.11 $Y2=0
r299 152 181 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=12.19 $Y2=0
r300 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r301 149 180 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.295 $Y=0
+ $X2=12.16 $Y2=0
r302 149 151 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=12.295 $Y=0
+ $X2=12.65 $Y2=0
r303 148 183 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.965 $Y=0
+ $X2=13.1 $Y2=0
r304 148 151 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.965 $Y=0
+ $X2=12.65 $Y2=0
r305 147 181 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.19 $Y2=0
r306 147 178 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=11.27 $Y2=0
r307 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r308 144 177 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.355 $Y=0
+ $X2=11.22 $Y2=0
r309 144 146 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.355 $Y=0
+ $X2=11.73 $Y2=0
r310 143 180 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.025 $Y=0
+ $X2=12.16 $Y2=0
r311 143 146 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.025 $Y=0
+ $X2=11.73 $Y2=0
r312 142 178 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.27 $Y2=0
r313 141 142 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r314 139 177 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.085 $Y=0
+ $X2=11.22 $Y2=0
r315 139 141 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.085 $Y=0
+ $X2=10.81 $Y2=0
r316 138 142 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.81 $Y2=0
r317 137 138 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r318 135 138 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=9.89 $Y2=0
r319 134 137 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=7.59 $Y=0
+ $X2=9.89 $Y2=0
r320 134 135 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r321 132 135 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=7.59 $Y2=0
r322 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r323 129 132 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.13 $Y2=0
r324 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r325 126 129 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.21 $Y2=0
r326 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r327 123 126 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.29 $Y2=0
r328 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r329 120 123 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.37 $Y2=0
r330 120 175 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=2.53 $Y2=0
r331 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r332 117 174 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.795 $Y=0
+ $X2=2.66 $Y2=0
r333 117 119 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.795 $Y=0
+ $X2=3.45 $Y2=0
r334 114 196 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r335 112 174 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.525 $Y=0
+ $X2=2.66 $Y2=0
r336 112 114 149.727 $w=1.68e-07 $l=2.295e-06 $layer=LI1_cond $X=2.525 $Y=0
+ $X2=0.23 $Y2=0
r337 110 175 0.653023 $w=4.8e-07 $l=2.295e-06 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=2.53 $Y2=0
r338 110 196 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r339 108 137 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=10.145 $Y=0
+ $X2=9.89 $Y2=0
r340 108 109 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.145 $Y=0
+ $X2=10.28 $Y2=0
r341 107 141 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.415 $Y=0
+ $X2=10.81 $Y2=0
r342 107 109 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.415 $Y=0
+ $X2=10.28 $Y2=0
r343 105 131 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.225 $Y=0
+ $X2=7.13 $Y2=0
r344 105 106 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.225 $Y=0
+ $X2=7.36 $Y2=0
r345 104 134 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.495 $Y=0
+ $X2=7.59 $Y2=0
r346 104 106 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.495 $Y=0
+ $X2=7.36 $Y2=0
r347 102 128 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.285 $Y=0
+ $X2=6.21 $Y2=0
r348 102 103 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.285 $Y=0
+ $X2=6.42 $Y2=0
r349 101 131 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.555 $Y=0
+ $X2=7.13 $Y2=0
r350 101 103 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.555 $Y=0
+ $X2=6.42 $Y2=0
r351 99 125 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=5.345 $Y=0
+ $X2=5.29 $Y2=0
r352 99 100 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.345 $Y=0
+ $X2=5.48 $Y2=0
r353 98 128 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.615 $Y=0
+ $X2=6.21 $Y2=0
r354 98 100 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.615 $Y=0
+ $X2=5.48 $Y2=0
r355 96 122 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.405 $Y=0
+ $X2=4.37 $Y2=0
r356 96 97 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.405 $Y=0 $X2=4.54
+ $Y2=0
r357 95 125 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.675 $Y=0
+ $X2=5.29 $Y2=0
r358 95 97 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.675 $Y=0 $X2=4.54
+ $Y2=0
r359 93 119 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.465 $Y=0
+ $X2=3.45 $Y2=0
r360 93 94 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.465 $Y=0 $X2=3.6
+ $Y2=0
r361 92 122 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.735 $Y=0
+ $X2=4.37 $Y2=0
r362 92 94 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.735 $Y=0 $X2=3.6
+ $Y2=0
r363 88 192 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.92 $Y=0.085
+ $X2=15.92 $Y2=0
r364 88 90 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=15.92 $Y=0.085
+ $X2=15.92 $Y2=0.38
r365 84 189 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.98 $Y=0.085
+ $X2=14.98 $Y2=0
r366 84 86 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=14.98 $Y=0.085
+ $X2=14.98 $Y2=0.38
r367 80 186 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.04 $Y=0.085
+ $X2=14.04 $Y2=0
r368 80 82 12.8049 $w=2.68e-07 $l=3e-07 $layer=LI1_cond $X=14.04 $Y=0.085
+ $X2=14.04 $Y2=0.385
r369 76 183 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.1 $Y=0.085
+ $X2=13.1 $Y2=0
r370 76 78 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.1 $Y=0.085
+ $X2=13.1 $Y2=0.38
r371 72 180 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.16 $Y=0.085
+ $X2=12.16 $Y2=0
r372 72 74 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.16 $Y=0.085
+ $X2=12.16 $Y2=0.38
r373 68 177 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.22 $Y=0.085
+ $X2=11.22 $Y2=0
r374 68 70 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=11.22 $Y=0.085
+ $X2=11.22 $Y2=0.38
r375 64 109 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.28 $Y=0.085
+ $X2=10.28 $Y2=0
r376 64 66 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.28 $Y=0.085
+ $X2=10.28 $Y2=0.38
r377 60 106 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0
r378 60 62 12.8049 $w=2.68e-07 $l=3e-07 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0.385
r379 56 103 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0
r380 56 58 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0.38
r381 52 100 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0
r382 52 54 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.38
r383 48 97 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0
r384 48 50 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0.38
r385 44 94 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=0.085
+ $X2=3.6 $Y2=0
r386 44 46 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.6 $Y=0.085
+ $X2=3.6 $Y2=0.38
r387 40 174 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=0.085
+ $X2=2.66 $Y2=0
r388 40 42 12.8049 $w=2.68e-07 $l=3e-07 $layer=LI1_cond $X=2.66 $Y=0.085
+ $X2=2.66 $Y2=0.385
r389 13 90 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=15.735
+ $Y=0.235 $X2=15.92 $Y2=0.38
r390 12 86 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=14.795
+ $Y=0.235 $X2=14.98 $Y2=0.38
r391 11 82 182 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_NDIFF $count=1 $X=13.855
+ $Y=0.235 $X2=14.04 $Y2=0.385
r392 10 78 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=12.915
+ $Y=0.235 $X2=13.1 $Y2=0.38
r393 9 74 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=11.975
+ $Y=0.235 $X2=12.16 $Y2=0.38
r394 8 70 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=11.035
+ $Y=0.235 $X2=11.22 $Y2=0.38
r395 7 66 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=10.155
+ $Y=0.235 $X2=10.28 $Y2=0.38
r396 6 62 182 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_NDIFF $count=1 $X=7.175
+ $Y=0.235 $X2=7.36 $Y2=0.385
r397 5 58 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=6.235
+ $Y=0.235 $X2=6.42 $Y2=0.38
r398 4 54 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=5.295
+ $Y=0.235 $X2=5.48 $Y2=0.38
r399 3 50 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=4.355
+ $Y=0.235 $X2=4.54 $Y2=0.38
r400 2 46 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.235 $X2=3.6 $Y2=0.38
r401 1 42 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.235 $X2=2.66 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_12%A_1163_47# 1 2 3 4 15 17 18 21 27 30 31 33
+ 34
r87 33 34 8.14364 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=9.29 $Y=0.75
+ $X2=9.125 $Y2=0.75
r88 31 34 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=8.515 $Y=0.815
+ $X2=9.125 $Y2=0.815
r89 29 31 8.14364 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=8.35 $Y=0.75
+ $X2=8.515 $Y2=0.75
r90 29 30 8.14364 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=8.35 $Y=0.75
+ $X2=8.185 $Y2=0.75
r91 24 27 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.055 $Y=0.815
+ $X2=6.89 $Y2=0.815
r92 24 30 69.6263 $w=1.78e-07 $l=1.13e-06 $layer=LI1_cond $X=7.055 $Y=0.815
+ $X2=8.185 $Y2=0.815
r93 19 27 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=6.89 $Y=0.725 $X2=6.89
+ $Y2=0.815
r94 19 21 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.89 $Y=0.725
+ $X2=6.89 $Y2=0.42
r95 17 27 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.725 $Y=0.815
+ $X2=6.89 $Y2=0.815
r96 17 18 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=6.725 $Y=0.815
+ $X2=6.115 $Y2=0.815
r97 13 18 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=5.95 $Y=0.725
+ $X2=6.115 $Y2=0.815
r98 13 15 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=5.95 $Y=0.725
+ $X2=5.95 $Y2=0.42
r99 4 33 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=9.155
+ $Y=0.235 $X2=9.29 $Y2=0.76
r100 3 29 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=8.215
+ $Y=0.235 $X2=8.35 $Y2=0.76
r101 2 21 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=6.755
+ $Y=0.235 $X2=6.89 $Y2=0.42
r102 1 15 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=5.815
+ $Y=0.235 $X2=5.95 $Y2=0.42
.ends

