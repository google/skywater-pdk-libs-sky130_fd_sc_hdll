* File: sky130_fd_sc_hdll__nand2_4.pex.spice
* Created: Thu Aug 27 19:12:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND2_4%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 27 28 45 50 53 56 59
r84 45 46 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=1.93 $Y2=1.202
r85 43 45 31.0329 $w=3.65e-07 $l=2.35e-07 $layer=POLY_cond $X=1.67 $Y=1.202
+ $X2=1.905 $Y2=1.202
r86 43 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.67
+ $Y=1.16 $X2=1.67 $Y2=1.16
r87 41 43 27.7315 $w=3.65e-07 $l=2.1e-07 $layer=POLY_cond $X=1.46 $Y=1.202
+ $X2=1.67 $Y2=1.202
r88 40 41 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.46 $Y2=1.202
r89 39 40 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=0.99 $Y=1.202
+ $X2=1.435 $Y2=1.202
r90 38 39 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r91 37 38 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.965 $Y2=1.202
r92 36 37 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r93 34 36 29.0521 $w=3.65e-07 $l=2.2e-07 $layer=POLY_cond $X=0.275 $Y=1.202
+ $X2=0.495 $Y2=1.202
r94 34 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r95 28 59 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.61 $Y=1.2 $X2=1.615
+ $Y2=1.2
r96 28 56 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=1.61 $Y=1.2
+ $X2=1.155 $Y2=1.2
r97 27 56 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.15 $Y=1.2 $X2=1.155
+ $Y2=1.2
r98 27 53 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=1.15 $Y=1.2
+ $X2=0.695 $Y2=1.2
r99 26 53 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.69 $Y=1.2 $X2=0.695
+ $Y2=1.2
r100 26 50 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=0.69 $Y=1.2
+ $X2=0.235 $Y2=1.2
r101 25 50 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.23 $Y=1.2
+ $X2=0.235 $Y2=1.2
r102 22 46 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r103 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r104 19 45 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r105 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r106 16 41 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=1.202
r107 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=0.56
r108 13 40 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r109 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r110 10 39 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r111 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r112 7 38 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r113 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r114 4 37 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r115 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=0.56
r116 1 36 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r117 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 37 38 43 46
c74 1 0 1.56657e-19 $X=2.35 $Y=0.995
r75 38 39 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.785 $Y=1.202
+ $X2=3.81 $Y2=1.202
r76 37 46 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=3.55 $Y=1.2
+ $X2=3.455 $Y2=1.2
r77 36 38 30.4489 $w=3.72e-07 $l=2.35e-07 $layer=POLY_cond $X=3.55 $Y=1.202
+ $X2=3.785 $Y2=1.202
r78 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.55
+ $Y=1.16 $X2=3.55 $Y2=1.16
r79 34 36 30.4489 $w=3.72e-07 $l=2.35e-07 $layer=POLY_cond $X=3.315 $Y=1.202
+ $X2=3.55 $Y2=1.202
r80 33 34 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.202
+ $X2=3.315 $Y2=1.202
r81 32 33 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=3.29 $Y2=1.202
r82 31 32 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.845 $Y2=1.202
r83 30 31 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.82 $Y2=1.202
r84 29 30 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.202
+ $X2=2.375 $Y2=1.202
r85 26 46 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=3.45 $Y=1.2 $X2=3.455
+ $Y2=1.2
r86 26 43 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=3.45 $Y=1.2
+ $X2=2.995 $Y2=1.2
r87 25 43 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=2.99 $Y=1.2 $X2=2.995
+ $Y2=1.2
r88 22 39 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=1.202
r89 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=0.56
r90 19 38 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.202
r91 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r92 16 34 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.202
r93 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r94 13 33 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=1.202
r95 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=0.56
r96 10 32 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r97 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r98 7 31 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=1.202
r99 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.82 $Y=0.995 $X2=2.82
+ $Y2=0.56
r100 4 30 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r101 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r102 1 29 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.202
r103 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_4%VPWR 1 2 3 4 5 16 18 22 26 28 32 36 40 43
+ 44 46 47 48 58 59 65 68
r72 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r73 66 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r74 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r75 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r76 56 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r77 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r78 53 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r79 53 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r80 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r81 50 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.14 $Y2=2.72
r82 50 52 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.99 $Y2=2.72
r83 48 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r84 48 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r85 46 55 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.935 $Y=2.72
+ $X2=3.91 $Y2=2.72
r86 46 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.935 $Y=2.72
+ $X2=4.06 $Y2=2.72
r87 45 58 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.185 $Y=2.72
+ $X2=4.37 $Y2=2.72
r88 45 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.185 $Y=2.72
+ $X2=4.06 $Y2=2.72
r89 43 52 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.995 $Y=2.72
+ $X2=2.99 $Y2=2.72
r90 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=2.72
+ $X2=3.08 $Y2=2.72
r91 42 55 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3.165 $Y=2.72
+ $X2=3.91 $Y2=2.72
r92 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=2.72
+ $X2=3.08 $Y2=2.72
r93 38 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.06 $Y=2.635
+ $X2=4.06 $Y2=2.72
r94 38 40 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=4.06 $Y=2.635
+ $X2=4.06 $Y2=2
r95 34 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2.72
r96 34 36 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2
r97 30 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.72
r98 30 32 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2
r99 29 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.72 $X2=1.2
+ $Y2=2.72
r100 28 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=2.14 $Y2=2.72
r101 28 29 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=1.285 $Y2=2.72
r102 24 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.72
r103 24 26 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r104 23 62 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r105 22 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=1.2 $Y2=2.72
r106 22 23 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=0.345 $Y2=2.72
r107 18 21 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.34
r108 16 62 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r109 16 21 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.34
r110 5 40 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=2
r111 4 36 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2
r112 3 32 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r113 2 26 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r114 1 21 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r115 1 18 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_4%Y 1 2 3 4 5 6 19 21 23 27 29 33 37 39 41
+ 43 48 49 54 55
r93 55 59 1.23714 $w=3e-07 $l=1.03078e-07 $layer=LI1_cond $X=2.585 $Y=1.58
+ $X2=2.545 $Y2=1.495
r94 55 59 0.960369 $w=2.98e-07 $l=2.5e-08 $layer=LI1_cond $X=2.545 $Y=1.47
+ $X2=2.545 $Y2=1.495
r95 54 55 10.7561 $w=2.98e-07 $l=2.8e-07 $layer=LI1_cond $X=2.545 $Y=1.19
+ $X2=2.545 $Y2=1.47
r96 49 54 14.7897 $w=2.98e-07 $l=3.85e-07 $layer=LI1_cond $X=2.545 $Y=0.805
+ $X2=2.545 $Y2=1.19
r97 49 51 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=0.805
+ $X2=2.545 $Y2=0.72
r98 41 53 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=1.665
+ $X2=3.525 $Y2=1.58
r99 41 43 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=3.525 $Y=1.665
+ $X2=3.525 $Y2=2.34
r100 40 55 5.3802 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=1.58
+ $X2=2.585 $Y2=1.58
r101 39 53 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.335 $Y=1.58
+ $X2=3.525 $Y2=1.58
r102 39 40 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.335 $Y=1.58
+ $X2=2.775 $Y2=1.58
r103 35 51 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.695 $Y=0.72
+ $X2=2.545 $Y2=0.72
r104 35 37 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=2.695 $Y=0.72
+ $X2=3.55 $Y2=0.72
r105 31 55 1.23714 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=1.665
+ $X2=2.585 $Y2=1.58
r106 31 33 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=2.585 $Y=1.665
+ $X2=2.585 $Y2=2.34
r107 30 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=1.58
+ $X2=1.645 $Y2=1.58
r108 29 55 5.3802 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=1.58
+ $X2=2.585 $Y2=1.58
r109 29 30 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.395 $Y=1.58
+ $X2=1.835 $Y2=1.58
r110 25 48 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.645 $Y2=1.58
r111 25 27 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.645 $Y2=2.34
r112 24 46 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.705 $Y2=1.58
r113 23 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=1.58
+ $X2=1.645 $Y2=1.58
r114 23 24 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.455 $Y=1.58
+ $X2=0.895 $Y2=1.58
r115 19 46 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=1.58
r116 19 21 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=2.34
r117 6 53 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.66
r118 6 43 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2.34
r119 5 55 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.66
r120 5 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.34
r121 4 48 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r122 4 27 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
r123 3 46 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r124 3 21 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r125 2 37 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.72
r126 1 51 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_4%A_27_47# 1 2 3 4 5 18 20 21 24 26 28 29 30
+ 34 36 38
c70 29 0 1.56657e-19 $X=2.075 $Y=0.715
r71 34 44 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=4.06 $Y=0.465
+ $X2=4.06 $Y2=0.36
r72 34 36 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.06 $Y=0.465
+ $X2=4.06 $Y2=0.72
r73 31 40 4.17428 $w=2.1e-07 $l=1.5e-07 $layer=LI1_cond $X=2.225 $Y=0.36
+ $X2=2.075 $Y2=0.36
r74 31 33 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=2.225 $Y=0.36
+ $X2=3.08 $Y2=0.36
r75 30 44 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=3.935 $Y=0.36
+ $X2=4.06 $Y2=0.36
r76 30 33 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=3.935 $Y=0.36
+ $X2=3.08 $Y2=0.36
r77 29 42 2.82016 $w=3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.075 $Y=0.715
+ $X2=2.075 $Y2=0.81
r78 28 40 2.92199 $w=3e-07 $l=1.05e-07 $layer=LI1_cond $X=2.075 $Y=0.465
+ $X2=2.075 $Y2=0.36
r79 28 29 9.60369 $w=2.98e-07 $l=2.5e-07 $layer=LI1_cond $X=2.075 $Y=0.465
+ $X2=2.075 $Y2=0.715
r80 27 38 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=1.365 $Y=0.81
+ $X2=1.175 $Y2=0.81
r81 26 42 4.45288 $w=1.9e-07 $l=1.5e-07 $layer=LI1_cond $X=1.925 $Y=0.81
+ $X2=2.075 $Y2=0.81
r82 26 27 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=1.925 $Y=0.81
+ $X2=1.365 $Y2=0.81
r83 22 38 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=1.175 $Y=0.715
+ $X2=1.175 $Y2=0.81
r84 22 24 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.175 $Y=0.715
+ $X2=1.175 $Y2=0.38
r85 20 38 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=0.985 $Y=0.81
+ $X2=1.175 $Y2=0.81
r86 20 21 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=0.985 $Y=0.81
+ $X2=0.425 $Y2=0.81
r87 16 21 7.51555 $w=1.9e-07 $l=2.102e-07 $layer=LI1_cond $X=0.257 $Y=0.715
+ $X2=0.425 $Y2=0.81
r88 16 18 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=0.257 $Y=0.715
+ $X2=0.257 $Y2=0.38
r89 5 44 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.235 $X2=4.02 $Y2=0.38
r90 5 36 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.235 $X2=4.02 $Y2=0.72
r91 4 33 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.38
r92 3 42 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.72
r93 3 40 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.38
r94 2 24 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.38
r95 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_4%VGND 1 2 11 13 17 19 26 27 30 33
r57 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r58 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r59 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r60 26 27 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r61 24 27 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=4.37
+ $Y2=0
r62 24 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r63 23 26 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=4.37
+ $Y2=0
r64 23 24 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r65 21 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=0 $X2=1.67
+ $Y2=0
r66 21 23 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.755 $Y=0 $X2=2.07
+ $Y2=0
r67 19 31 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r68 15 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0
r69 15 17 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0.38
r70 14 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.73
+ $Y2=0
r71 13 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=0 $X2=1.67
+ $Y2=0
r72 13 14 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.585 $Y=0 $X2=0.815
+ $Y2=0
r73 9 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085 $X2=0.73
+ $Y2=0
r74 9 11 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.38
r75 2 17 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.38
r76 1 11 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

