* File: sky130_fd_sc_hdll__a221oi_4.pex.spice
* Created: Thu Aug 27 18:53:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A221OI_4%C1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 36 39
r76 39 40 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.925 $Y=1.202
+ $X2=1.95 $Y2=1.202
r77 38 39 57.9703 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=1.48 $Y=1.202
+ $X2=1.925 $Y2=1.202
r78 37 38 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.48 $Y2=1.202
r79 35 37 24.1 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=1.27 $Y=1.202
+ $X2=1.455 $Y2=1.202
r80 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.27
+ $Y=1.16 $X2=1.27 $Y2=1.16
r81 33 35 33.8703 $w=3.7e-07 $l=2.6e-07 $layer=POLY_cond $X=1.01 $Y=1.202
+ $X2=1.27 $Y2=1.202
r82 32 33 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.01 $Y2=1.202
r83 31 32 57.9703 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=0.54 $Y=1.202
+ $X2=0.985 $Y2=1.202
r84 30 31 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.54 $Y2=1.202
r85 28 30 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.49 $Y=1.202
+ $X2=0.515 $Y2=1.202
r86 28 29 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.49
+ $Y=1.16 $X2=0.49 $Y2=1.16
r87 25 36 6.37727 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=1.27 $Y2=1.175
r88 25 29 36.8773 $w=1.98e-07 $l=6.65e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=0.49 $Y2=1.175
r89 22 40 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=1.202
r90 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=0.56
r91 19 39 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r92 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r93 16 38 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.48 $Y=0.995
+ $X2=1.48 $Y2=1.202
r94 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.48 $Y=0.995
+ $X2=1.48 $Y2=0.56
r95 13 37 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r96 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r97 10 33 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=1.202
r98 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=0.56
r99 7 32 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r100 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r101 4 31 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.54 $Y2=1.202
r102 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.54 $Y2=0.56
r103 1 30 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r104 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_4%B2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 27 31 32 35 36 47
c121 10 0 1.43003e-19 $X=3.38 $Y=0.995
c122 4 0 1.71792e-19 $X=2.91 $Y=0.995
r123 41 42 7.36389 $w=3.6e-07 $l=5.5e-08 $layer=POLY_cond $X=3.38 $Y=1.202
+ $X2=3.435 $Y2=1.202
r124 40 41 55.5639 $w=3.6e-07 $l=4.15e-07 $layer=POLY_cond $X=2.965 $Y=1.202
+ $X2=3.38 $Y2=1.202
r125 39 40 7.36389 $w=3.6e-07 $l=5.5e-08 $layer=POLY_cond $X=2.91 $Y=1.202
+ $X2=2.965 $Y2=1.202
r126 38 39 62.9278 $w=3.6e-07 $l=4.7e-07 $layer=POLY_cond $X=2.44 $Y=1.202
+ $X2=2.91 $Y2=1.202
r127 36 47 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.335 $Y=1.53
+ $X2=4.29 $Y2=1.53
r128 35 36 112.866 $w=1.68e-07 $l=1.73e-06 $layer=LI1_cond $X=6.065 $Y=1.53
+ $X2=4.335 $Y2=1.53
r129 34 47 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.165 $Y=1.53
+ $X2=4.29 $Y2=1.53
r130 33 34 4.34843 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=3.965 $Y=1.53
+ $X2=4.165 $Y2=1.53
r131 32 44 7.36389 $w=3.6e-07 $l=5.5e-08 $layer=POLY_cond $X=3.85 $Y=1.202
+ $X2=3.905 $Y2=1.202
r132 32 42 55.5639 $w=3.6e-07 $l=4.15e-07 $layer=POLY_cond $X=3.85 $Y=1.202
+ $X2=3.435 $Y2=1.202
r133 31 33 14.3302 $w=3.15e-07 $l=3.7e-07 $layer=LI1_cond $X=3.965 $Y=1.16
+ $X2=3.965 $Y2=1.53
r134 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.85
+ $Y=1.16 $X2=3.85 $Y2=1.16
r135 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.23
+ $Y=1.16 $X2=6.23 $Y2=1.16
r136 25 35 7.89393 $w=1.7e-07 $l=2.10247e-07 $layer=LI1_cond $X=6.237 $Y=1.445
+ $X2=6.065 $Y2=1.53
r137 25 27 9.52018 $w=3.43e-07 $l=2.85e-07 $layer=LI1_cond $X=6.237 $Y=1.445
+ $X2=6.237 $Y2=1.16
r138 22 28 38.6443 $w=2.87e-07 $l=1.79374e-07 $layer=POLY_cond $X=6.28 $Y=0.995
+ $X2=6.25 $Y2=1.16
r139 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.28 $Y=0.995
+ $X2=6.28 $Y2=0.56
r140 19 28 48.651 $w=2.87e-07 $l=2.52488e-07 $layer=POLY_cond $X=6.255 $Y=1.41
+ $X2=6.25 $Y2=1.16
r141 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.255 $Y=1.41
+ $X2=6.255 $Y2=1.985
r142 16 44 18.9685 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.905 $Y=1.41
+ $X2=3.905 $Y2=1.202
r143 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.905 $Y=1.41
+ $X2=3.905 $Y2=1.985
r144 13 42 18.9685 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.435 $Y=1.41
+ $X2=3.435 $Y2=1.202
r145 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.435 $Y=1.41
+ $X2=3.435 $Y2=1.985
r146 10 41 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.38 $Y=0.995
+ $X2=3.38 $Y2=1.202
r147 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.38 $Y=0.995
+ $X2=3.38 $Y2=0.56
r148 7 40 18.9685 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.965 $Y=1.41
+ $X2=2.965 $Y2=1.202
r149 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.965 $Y=1.41
+ $X2=2.965 $Y2=1.985
r150 4 39 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.91 $Y=0.995
+ $X2=2.91 $Y2=1.202
r151 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.91 $Y=0.995
+ $X2=2.91 $Y2=0.56
r152 1 38 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.44 $Y=0.995
+ $X2=2.44 $Y2=1.202
r153 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.44 $Y=0.995
+ $X2=2.44 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_4%B1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39 45
r66 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.785 $Y=1.202
+ $X2=5.81 $Y2=1.202
r67 38 45 33.1327 $w=2.78e-07 $l=8.05e-07 $layer=LI1_cond $X=5.67 $Y=1.135
+ $X2=4.865 $Y2=1.135
r68 37 39 14.9005 $w=3.72e-07 $l=1.15e-07 $layer=POLY_cond $X=5.67 $Y=1.202
+ $X2=5.785 $Y2=1.202
r69 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.67
+ $Y=1.16 $X2=5.67 $Y2=1.16
r70 35 37 45.9973 $w=3.72e-07 $l=3.55e-07 $layer=POLY_cond $X=5.315 $Y=1.202
+ $X2=5.67 $Y2=1.202
r71 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.29 $Y=1.202
+ $X2=5.315 $Y2=1.202
r72 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=4.845 $Y=1.202
+ $X2=5.29 $Y2=1.202
r73 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.82 $Y=1.202
+ $X2=4.845 $Y2=1.202
r74 30 32 41.4624 $w=3.72e-07 $l=3.2e-07 $layer=POLY_cond $X=4.5 $Y=1.202
+ $X2=4.82 $Y2=1.202
r75 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.5 $Y=1.16
+ $X2=4.5 $Y2=1.16
r76 28 30 16.1962 $w=3.72e-07 $l=1.25e-07 $layer=POLY_cond $X=4.375 $Y=1.202
+ $X2=4.5 $Y2=1.202
r77 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.35 $Y=1.202
+ $X2=4.375 $Y2=1.202
r78 25 45 0.823174 $w=2.78e-07 $l=2e-08 $layer=LI1_cond $X=4.845 $Y=1.135
+ $X2=4.865 $Y2=1.135
r79 25 31 14.1997 $w=2.78e-07 $l=3.45e-07 $layer=LI1_cond $X=4.845 $Y=1.135
+ $X2=4.5 $Y2=1.135
r80 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.81 $Y=0.995
+ $X2=5.81 $Y2=1.202
r81 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.81 $Y=0.995
+ $X2=5.81 $Y2=0.56
r82 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.785 $Y=1.41
+ $X2=5.785 $Y2=1.202
r83 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.785 $Y=1.41
+ $X2=5.785 $Y2=1.985
r84 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.315 $Y=1.41
+ $X2=5.315 $Y2=1.202
r85 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.315 $Y=1.41
+ $X2=5.315 $Y2=1.985
r86 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.29 $Y=0.995
+ $X2=5.29 $Y2=1.202
r87 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.29 $Y=0.995
+ $X2=5.29 $Y2=0.56
r88 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.845 $Y=1.41
+ $X2=4.845 $Y2=1.202
r89 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.845 $Y=1.41
+ $X2=4.845 $Y2=1.985
r90 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.82 $Y=0.995
+ $X2=4.82 $Y2=1.202
r91 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.82 $Y=0.995 $X2=4.82
+ $Y2=0.56
r92 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.375 $Y=1.41
+ $X2=4.375 $Y2=1.202
r93 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.375 $Y=1.41
+ $X2=4.375 $Y2=1.985
r94 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=1.202
r95 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.35 $Y=0.995 $X2=4.35
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_4%A2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 28 30 35 36 48 49 53
c122 1 0 1.20734e-19 $X=6.775 $Y=1.41
r123 49 50 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=10.04 $Y=1.202
+ $X2=10.065 $Y2=1.202
r124 47 49 9.04558 $w=3.73e-07 $l=7e-08 $layer=POLY_cond $X=9.97 $Y=1.202
+ $X2=10.04 $Y2=1.202
r125 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9.97
+ $Y=1.16 $X2=9.97 $Y2=1.16
r126 45 47 48.4584 $w=3.73e-07 $l=3.75e-07 $layer=POLY_cond $X=9.595 $Y=1.202
+ $X2=9.97 $Y2=1.202
r127 44 45 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=9.57 $Y=1.202
+ $X2=9.595 $Y2=1.202
r128 43 53 6.1 $w=1.98e-07 $l=1.1e-07 $layer=LI1_cond $X=9.19 $Y=1.175 $X2=9.3
+ $Y2=1.175
r129 42 44 49.1046 $w=3.73e-07 $l=3.8e-07 $layer=POLY_cond $X=9.19 $Y=1.202
+ $X2=9.57 $Y2=1.202
r130 42 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9.19
+ $Y=1.16 $X2=9.19 $Y2=1.16
r131 40 42 8.39946 $w=3.73e-07 $l=6.5e-08 $layer=POLY_cond $X=9.125 $Y=1.202
+ $X2=9.19 $Y2=1.202
r132 39 40 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=9.1 $Y=1.202
+ $X2=9.125 $Y2=1.202
r133 36 48 28.5591 $w=1.98e-07 $l=5.15e-07 $layer=LI1_cond $X=9.455 $Y=1.175
+ $X2=9.97 $Y2=1.175
r134 36 53 8.59545 $w=1.98e-07 $l=1.55e-07 $layer=LI1_cond $X=9.455 $Y=1.175
+ $X2=9.3 $Y2=1.175
r135 35 43 3.05 $w=1.98e-07 $l=5.5e-08 $layer=LI1_cond $X=9.135 $Y=1.175
+ $X2=9.19 $Y2=1.175
r136 30 33 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=6.775 $Y=1.16
+ $X2=6.775 $Y2=1.53
r137 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.75
+ $Y=1.16 $X2=6.75 $Y2=1.16
r138 27 35 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=9.05 $Y=1.275
+ $X2=9.135 $Y2=1.175
r139 27 28 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.05 $Y=1.275
+ $X2=9.05 $Y2=1.445
r140 26 33 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.965 $Y=1.53
+ $X2=6.775 $Y2=1.53
r141 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.965 $Y=1.53
+ $X2=9.05 $Y2=1.445
r142 25 26 130.481 $w=1.68e-07 $l=2e-06 $layer=LI1_cond $X=8.965 $Y=1.53
+ $X2=6.965 $Y2=1.53
r143 22 50 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.065 $Y=1.41
+ $X2=10.065 $Y2=1.202
r144 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.065 $Y=1.41
+ $X2=10.065 $Y2=1.985
r145 19 49 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.04 $Y=0.995
+ $X2=10.04 $Y2=1.202
r146 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.04 $Y=0.995
+ $X2=10.04 $Y2=0.56
r147 16 45 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.595 $Y=1.41
+ $X2=9.595 $Y2=1.202
r148 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.595 $Y=1.41
+ $X2=9.595 $Y2=1.985
r149 13 44 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.57 $Y=0.995
+ $X2=9.57 $Y2=1.202
r150 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.57 $Y=0.995
+ $X2=9.57 $Y2=0.56
r151 10 40 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.125 $Y=1.41
+ $X2=9.125 $Y2=1.202
r152 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.125 $Y=1.41
+ $X2=9.125 $Y2=1.985
r153 7 39 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.1 $Y=0.995 $X2=9.1
+ $Y2=1.202
r154 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.1 $Y=0.995 $X2=9.1
+ $Y2=0.56
r155 4 31 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=6.8 $Y=0.995
+ $X2=6.775 $Y2=1.16
r156 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.8 $Y=0.995 $X2=6.8
+ $Y2=0.56
r157 1 31 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=6.775 $Y=1.41
+ $X2=6.775 $Y2=1.16
r158 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.775 $Y=1.41
+ $X2=6.775 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_4%A1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 36 39 44
r60 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.655 $Y=1.202
+ $X2=8.68 $Y2=1.202
r61 38 39 60.8979 $w=3.72e-07 $l=4.7e-07 $layer=POLY_cond $X=8.185 $Y=1.202
+ $X2=8.655 $Y2=1.202
r62 37 38 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.16 $Y=1.202
+ $X2=8.185 $Y2=1.202
r63 35 37 9.06989 $w=3.72e-07 $l=7e-08 $layer=POLY_cond $X=8.09 $Y=1.202
+ $X2=8.16 $Y2=1.202
r64 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.09
+ $Y=1.16 $X2=8.09 $Y2=1.16
r65 33 35 48.5887 $w=3.72e-07 $l=3.75e-07 $layer=POLY_cond $X=7.715 $Y=1.202
+ $X2=8.09 $Y2=1.202
r66 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.69 $Y=1.202
+ $X2=7.715 $Y2=1.202
r67 31 44 11.9227 $w=1.98e-07 $l=2.15e-07 $layer=LI1_cond $X=7.31 $Y=1.175
+ $X2=7.525 $Y2=1.175
r68 30 32 49.2366 $w=3.72e-07 $l=3.8e-07 $layer=POLY_cond $X=7.31 $Y=1.202
+ $X2=7.69 $Y2=1.202
r69 30 31 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.31
+ $Y=1.16 $X2=7.31 $Y2=1.16
r70 28 30 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=7.245 $Y=1.202
+ $X2=7.31 $Y2=1.202
r71 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.22 $Y=1.202
+ $X2=7.245 $Y2=1.202
r72 25 36 27.45 $w=1.98e-07 $l=4.95e-07 $layer=LI1_cond $X=7.595 $Y=1.175
+ $X2=8.09 $Y2=1.175
r73 25 44 3.88182 $w=1.98e-07 $l=7e-08 $layer=LI1_cond $X=7.595 $Y=1.175
+ $X2=7.525 $Y2=1.175
r74 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.68 $Y=0.995
+ $X2=8.68 $Y2=1.202
r75 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.68 $Y=0.995
+ $X2=8.68 $Y2=0.56
r76 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.655 $Y=1.41
+ $X2=8.655 $Y2=1.202
r77 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.655 $Y=1.41
+ $X2=8.655 $Y2=1.985
r78 16 38 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.185 $Y=1.41
+ $X2=8.185 $Y2=1.202
r79 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.185 $Y=1.41
+ $X2=8.185 $Y2=1.985
r80 13 37 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.16 $Y=0.995
+ $X2=8.16 $Y2=1.202
r81 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.16 $Y=0.995
+ $X2=8.16 $Y2=0.56
r82 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.715 $Y=1.41
+ $X2=7.715 $Y2=1.202
r83 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.715 $Y=1.41
+ $X2=7.715 $Y2=1.985
r84 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.69 $Y=0.995
+ $X2=7.69 $Y2=1.202
r85 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.69 $Y=0.995 $X2=7.69
+ $Y2=0.56
r86 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.245 $Y=1.41
+ $X2=7.245 $Y2=1.202
r87 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.245 $Y=1.41
+ $X2=7.245 $Y2=1.985
r88 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.22 $Y=0.995
+ $X2=7.22 $Y2=1.202
r89 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.22 $Y=0.995 $X2=7.22
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_4%A_27_297# 1 2 3 4 5 6 7 22 24 26 30 32 35
+ 37 38 39 41 43 50 54
r81 48 50 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=5.08 $Y=1.94 $X2=6.02
+ $Y2=1.94
r82 46 48 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=4.14 $Y=1.94 $X2=5.08
+ $Y2=1.94
r83 44 58 4.13622 $w=2.1e-07 $l=1.48e-07 $layer=LI1_cond $X=3.33 $Y=1.94
+ $X2=3.182 $Y2=1.94
r84 44 46 42.7792 $w=2.08e-07 $l=8.1e-07 $layer=LI1_cond $X=3.33 $Y=1.94
+ $X2=4.14 $Y2=1.94
r85 41 58 2.93448 $w=2.95e-07 $l=1.05e-07 $layer=LI1_cond $X=3.182 $Y=1.835
+ $X2=3.182 $Y2=1.94
r86 41 43 8.39916 $w=2.93e-07 $l=2.15e-07 $layer=LI1_cond $X=3.182 $Y=1.835
+ $X2=3.182 $Y2=1.62
r87 40 43 0.195329 $w=2.93e-07 $l=5e-09 $layer=LI1_cond $X=3.182 $Y=1.615
+ $X2=3.182 $Y2=1.62
r88 38 40 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=3.035 $Y=1.53
+ $X2=3.182 $Y2=1.615
r89 38 39 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.035 $Y=1.53
+ $X2=2.325 $Y2=1.53
r90 35 56 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=2.295 $X2=2.2
+ $Y2=2.38
r91 35 37 30.655 $w=2.48e-07 $l=6.65e-07 $layer=LI1_cond $X=2.2 $Y=2.295 $X2=2.2
+ $Y2=1.63
r92 34 39 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.2 $Y=1.615
+ $X2=2.325 $Y2=1.53
r93 34 37 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=2.2 $Y=1.615
+ $X2=2.2 $Y2=1.63
r94 33 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=2.38
+ $X2=1.22 $Y2=2.38
r95 32 56 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.075 $Y=2.38
+ $X2=2.2 $Y2=2.38
r96 32 33 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.075 $Y=2.38
+ $X2=1.345 $Y2=2.38
r97 28 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=2.295
+ $X2=1.22 $Y2=2.38
r98 28 30 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.22 $Y=2.295
+ $X2=1.22 $Y2=1.96
r99 27 53 4.96789 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=0.405 $Y=2.38
+ $X2=0.247 $Y2=2.38
r100 26 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=2.38
+ $X2=1.22 $Y2=2.38
r101 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=2.38
+ $X2=0.405 $Y2=2.38
r102 22 53 2.6726 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.247 $Y=2.295
+ $X2=0.247 $Y2=2.38
r103 22 24 24.6952 $w=3.13e-07 $l=6.75e-07 $layer=LI1_cond $X=0.247 $Y=2.295
+ $X2=0.247 $Y2=1.62
r104 7 50 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=5.875
+ $Y=1.485 $X2=6.02 $Y2=1.96
r105 6 48 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=4.935
+ $Y=1.485 $X2=5.08 $Y2=1.96
r106 5 46 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=3.995
+ $Y=1.485 $X2=4.14 $Y2=1.96
r107 4 58 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=3.055
+ $Y=1.485 $X2=3.2 $Y2=1.96
r108 4 43 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.055
+ $Y=1.485 $X2=3.2 $Y2=1.62
r109 3 56 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=2.31
r110 3 37 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=1.63
r111 2 30 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.96
r112 1 53 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r113 1 24 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_4%Y 1 2 3 4 5 6 7 8 27 31 33 34 35 36 39 43
+ 46 47 50 52 63 65 66 67 68 69 70 71 72
r147 70 71 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=6.96 $Y=0.775
+ $X2=7.13 $Y2=0.775
r148 69 70 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.28 $Y=0.82
+ $X2=6.96 $Y2=0.82
r149 68 69 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=6.11 $Y=0.775
+ $X2=6.28 $Y2=0.775
r150 66 72 6.57889 $w=3.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.755 $Y=1.445
+ $X2=1.755 $Y2=1.275
r151 66 67 4.06715 $w=2.25e-07 $l=1.05119e-07 $layer=LI1_cond $X=1.755 $Y=1.445
+ $X2=1.71 $Y2=1.53
r152 61 63 59.574 $w=1.73e-07 $l=9.4e-07 $layer=LI1_cond $X=7.48 $Y=0.732
+ $X2=8.42 $Y2=0.732
r153 61 71 22.1818 $w=1.73e-07 $l=3.5e-07 $layer=LI1_cond $X=7.48 $Y=0.732
+ $X2=7.13 $Y2=0.732
r154 56 68 35.4909 $w=1.73e-07 $l=5.6e-07 $layer=LI1_cond $X=5.55 $Y=0.732
+ $X2=6.11 $Y2=0.732
r155 54 56 59.574 $w=1.73e-07 $l=9.4e-07 $layer=LI1_cond $X=4.61 $Y=0.732
+ $X2=5.55 $Y2=0.732
r156 52 54 64.3273 $w=1.73e-07 $l=1.015e-06 $layer=LI1_cond $X=3.595 $Y=0.732
+ $X2=4.61 $Y2=0.732
r157 49 52 6.93219 $w=1.75e-07 $l=1.4758e-07 $layer=LI1_cond $X=3.485 $Y=0.82
+ $X2=3.595 $Y2=0.732
r158 49 50 14.4055 $w=2.18e-07 $l=2.75e-07 $layer=LI1_cond $X=3.485 $Y=0.82
+ $X2=3.485 $Y2=1.095
r159 48 72 1.72457 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=1.855 $Y=1.185
+ $X2=1.755 $Y2=1.185
r160 47 50 6.90553 $w=1.8e-07 $l=1.48324e-07 $layer=LI1_cond $X=3.375 $Y=1.185
+ $X2=3.485 $Y2=1.095
r161 47 48 93.6566 $w=1.78e-07 $l=1.52e-06 $layer=LI1_cond $X=3.375 $Y=1.185
+ $X2=1.855 $Y2=1.185
r162 46 72 4.72821 $w=2e-07 $l=9e-08 $layer=LI1_cond $X=1.755 $Y=1.095 $X2=1.755
+ $Y2=1.185
r163 45 65 3.41797 $w=2.9e-07 $l=1.27279e-07 $layer=LI1_cond $X=1.755 $Y=0.905
+ $X2=1.665 $Y2=0.815
r164 45 46 10.5364 $w=1.98e-07 $l=1.9e-07 $layer=LI1_cond $X=1.755 $Y=0.905
+ $X2=1.755 $Y2=1.095
r165 41 67 4.06715 $w=2.25e-07 $l=9.44722e-08 $layer=LI1_cond $X=1.69 $Y=1.615
+ $X2=1.71 $Y2=1.53
r166 41 43 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.69 $Y=1.615
+ $X2=1.69 $Y2=1.62
r167 37 65 3.41797 $w=2.9e-07 $l=9e-08 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.815
r168 37 39 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.39
r169 35 65 3.10432 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=1.665 $Y2=0.815
r170 35 36 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=0.915 $Y2=0.815
r171 33 67 2.36881 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.565 $Y=1.53
+ $X2=1.71 $Y2=1.53
r172 33 34 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.565 $Y=1.53
+ $X2=0.875 $Y2=1.53
r173 29 34 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.75 $Y=1.615
+ $X2=0.875 $Y2=1.53
r174 29 31 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.75 $Y=1.615
+ $X2=0.75 $Y2=1.62
r175 25 36 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.915 $Y2=0.815
r176 25 27 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.725 $Y2=0.39
r177 8 43 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=1.62
r178 7 31 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=1.62
r179 6 63 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=8.235
+ $Y=0.235 $X2=8.42 $Y2=0.73
r180 5 61 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=7.295
+ $Y=0.235 $X2=7.48 $Y2=0.73
r181 4 56 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=5.365
+ $Y=0.235 $X2=5.55 $Y2=0.73
r182 3 54 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.61 $Y2=0.73
r183 2 39 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.555
+ $Y=0.235 $X2=1.69 $Y2=0.39
r184 1 27 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.615
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_4%A_511_297# 1 2 3 4 5 6 7 8 9 28 30 32 40
+ 41 42 50 53 54 55 58 67
c94 40 0 1.20734e-19 $X=6.53 $Y=2.045
r95 56 58 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=10.3 $Y=1.615
+ $X2=10.3 $Y2=1.82
r96 54 56 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.175 $Y=1.53
+ $X2=10.3 $Y2=1.615
r97 54 55 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=10.175 $Y=1.53
+ $X2=9.525 $Y2=1.53
r98 53 67 7.24004 $w=1.7e-07 $l=1.48661e-07 $layer=LI1_cond $X=9.44 $Y=1.785
+ $X2=9.4 $Y2=1.915
r99 52 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.44 $Y=1.615
+ $X2=9.525 $Y2=1.53
r100 52 53 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.44 $Y=1.615
+ $X2=9.44 $Y2=1.785
r101 48 67 7.24004 $w=1.7e-07 $l=1.48661e-07 $layer=LI1_cond $X=9.36 $Y=2.045
+ $X2=9.4 $Y2=1.915
r102 48 50 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=9.36 $Y=2.045
+ $X2=9.36 $Y2=2.3
r103 45 47 41.6652 $w=2.58e-07 $l=9.4e-07 $layer=LI1_cond $X=7.48 $Y=1.915
+ $X2=8.42 $Y2=1.915
r104 43 63 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=6.655 $Y=1.915
+ $X2=6.53 $Y2=1.915
r105 43 45 36.5679 $w=2.58e-07 $l=8.25e-07 $layer=LI1_cond $X=6.655 $Y=1.915
+ $X2=7.48 $Y2=1.915
r106 42 67 0.132371 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=9.275 $Y=1.915
+ $X2=9.4 $Y2=1.915
r107 42 47 37.8976 $w=2.58e-07 $l=8.55e-07 $layer=LI1_cond $X=9.275 $Y=1.915
+ $X2=8.42 $Y2=1.915
r108 41 65 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.53 $Y=2.215
+ $X2=6.53 $Y2=2.34
r109 40 63 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=6.53 $Y=2.045
+ $X2=6.53 $Y2=1.915
r110 40 41 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=6.53 $Y=2.045
+ $X2=6.53 $Y2=2.215
r111 37 39 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=4.61 $Y=2.34
+ $X2=5.55 $Y2=2.34
r112 35 37 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=3.67 $Y=2.34
+ $X2=4.61 $Y2=2.34
r113 33 61 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=2.815 $Y=2.34
+ $X2=2.69 $Y2=2.34
r114 33 35 39.4136 $w=2.48e-07 $l=8.55e-07 $layer=LI1_cond $X=2.815 $Y=2.34
+ $X2=3.67 $Y2=2.34
r115 32 65 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.405 $Y=2.34
+ $X2=6.53 $Y2=2.34
r116 32 39 39.4136 $w=2.48e-07 $l=8.55e-07 $layer=LI1_cond $X=6.405 $Y=2.34
+ $X2=5.55 $Y2=2.34
r117 28 61 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=2.69 $Y=2.215
+ $X2=2.69 $Y2=2.34
r118 28 30 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=2.69 $Y=2.215
+ $X2=2.69 $Y2=1.96
r119 9 58 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=10.155
+ $Y=1.485 $X2=10.3 $Y2=1.82
r120 8 67 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=9.215
+ $Y=1.485 $X2=9.36 $Y2=1.96
r121 8 50 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=9.215
+ $Y=1.485 $X2=9.36 $Y2=2.3
r122 7 47 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=8.275
+ $Y=1.485 $X2=8.42 $Y2=1.96
r123 6 45 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=7.335
+ $Y=1.485 $X2=7.48 $Y2=1.96
r124 5 65 600 $w=1.7e-07 $l=9.02773e-07 $layer=licon1_PDIFF $count=1 $X=6.345
+ $Y=1.485 $X2=6.53 $Y2=2.3
r125 5 63 600 $w=1.7e-07 $l=5.59911e-07 $layer=licon1_PDIFF $count=1 $X=6.345
+ $Y=1.485 $X2=6.53 $Y2=1.96
r126 4 39 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.405
+ $Y=1.485 $X2=5.55 $Y2=2.3
r127 3 37 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.465
+ $Y=1.485 $X2=4.61 $Y2=2.3
r128 2 35 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.525
+ $Y=1.485 $X2=3.67 $Y2=2.3
r129 1 61 600 $w=1.7e-07 $l=8.98248e-07 $layer=licon1_PDIFF $count=1 $X=2.555
+ $Y=1.485 $X2=2.73 $Y2=2.3
r130 1 30 600 $w=1.7e-07 $l=5.55653e-07 $layer=licon1_PDIFF $count=1 $X=2.555
+ $Y=1.485 $X2=2.73 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_4%VPWR 1 2 3 4 15 17 21 23 24 25 34 45 46
+ 53
r108 51 53 9.0773 $w=5.88e-07 $l=1.15e-07 $layer=LI1_cond $X=8.97 $Y=2.51
+ $X2=9.085 $Y2=2.51
r109 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r110 49 51 1.6218 $w=5.88e-07 $l=8e-08 $layer=LI1_cond $X=8.89 $Y=2.51 $X2=8.97
+ $Y2=2.51
r111 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r112 43 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=10.35 $Y2=2.72
r113 43 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=8.97 $Y2=2.72
r114 42 53 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.43 $Y=2.72
+ $X2=9.085 $Y2=2.72
r115 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r116 37 52 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.97 $Y2=2.72
r117 36 39 16.6235 $w=5.88e-07 $l=8.2e-07 $layer=LI1_cond $X=7.13 $Y=2.51
+ $X2=7.95 $Y2=2.51
r118 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r119 34 49 2.02725 $w=5.88e-07 $l=1e-07 $layer=LI1_cond $X=8.79 $Y=2.51 $X2=8.89
+ $Y2=2.51
r120 34 39 17.0289 $w=5.88e-07 $l=8.4e-07 $layer=LI1_cond $X=8.79 $Y=2.51
+ $X2=7.95 $Y2=2.51
r121 33 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r122 32 33 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r123 28 32 420.15 $w=1.68e-07 $l=6.44e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=6.67 $Y2=2.72
r124 25 33 1.83245 $w=4.8e-07 $l=6.44e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=6.67 $Y2=2.72
r125 25 28 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r126 23 42 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.745 $Y=2.72
+ $X2=9.43 $Y2=2.72
r127 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.745 $Y=2.72
+ $X2=9.83 $Y2=2.72
r128 22 45 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=9.915 $Y=2.72
+ $X2=10.35 $Y2=2.72
r129 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.915 $Y=2.72
+ $X2=9.83 $Y2=2.72
r130 21 32 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=6.825 $Y=2.72
+ $X2=6.67 $Y2=2.72
r131 20 21 10.4964 $w=5.88e-07 $l=1.85e-07 $layer=LI1_cond $X=7.01 $Y=2.51
+ $X2=6.825 $Y2=2.51
r132 17 36 0.202725 $w=5.88e-07 $l=1e-08 $layer=LI1_cond $X=7.12 $Y=2.51
+ $X2=7.13 $Y2=2.51
r133 17 20 2.22998 $w=5.88e-07 $l=1.1e-07 $layer=LI1_cond $X=7.12 $Y=2.51
+ $X2=7.01 $Y2=2.51
r134 13 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.83 $Y=2.635
+ $X2=9.83 $Y2=2.72
r135 13 15 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=9.83 $Y=2.635
+ $X2=9.83 $Y2=1.96
r136 4 15 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=9.685
+ $Y=1.485 $X2=9.83 $Y2=1.96
r137 3 49 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=8.745
+ $Y=1.485 $X2=8.89 $Y2=2.3
r138 2 39 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=7.805
+ $Y=1.485 $X2=7.95 $Y2=2.3
r139 1 20 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=6.865
+ $Y=1.485 $X2=7.01 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_4%VGND 1 2 3 4 5 6 7 22 24 26 30 35 37 40
+ 44 46 48 51 52 54 55 58 59 61 62 63 81 89 93
r143 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r144 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r145 84 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.35 $Y2=0
r146 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r147 81 92 3.40825 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=10.165 $Y=0
+ $X2=10.372 $Y2=0
r148 81 83 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.165 $Y=0
+ $X2=9.89 $Y2=0
r149 80 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=9.89
+ $Y2=0
r150 79 80 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r151 77 80 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=6.67 $Y=0 $X2=8.97
+ $Y2=0
r152 76 79 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=6.67 $Y=0 $X2=8.97
+ $Y2=0
r153 76 77 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r154 74 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r155 73 74 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r156 71 74 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=2.53 $Y=0 $X2=6.21
+ $Y2=0
r157 70 73 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=6.21
+ $Y2=0
r158 70 71 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r159 68 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r160 68 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r161 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r162 65 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.22
+ $Y2=0
r163 65 67 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.305 $Y=0
+ $X2=2.07 $Y2=0
r164 63 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r165 63 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r166 61 79 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.275 $Y=0
+ $X2=8.97 $Y2=0
r167 61 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.275 $Y=0 $X2=9.36
+ $Y2=0
r168 60 83 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=9.445 $Y=0
+ $X2=9.89 $Y2=0
r169 60 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.445 $Y=0 $X2=9.36
+ $Y2=0
r170 58 73 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.455 $Y=0 $X2=6.21
+ $Y2=0
r171 58 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.455 $Y=0 $X2=6.54
+ $Y2=0
r172 57 76 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=6.625 $Y=0 $X2=6.67
+ $Y2=0
r173 57 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.625 $Y=0 $X2=6.54
+ $Y2=0
r174 54 55 3.26614 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=0.76
+ $X2=3.035 $Y2=0.76
r175 51 67 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.07
+ $Y2=0
r176 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.16
+ $Y2=0
r177 50 70 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.245 $Y=0
+ $X2=2.53 $Y2=0
r178 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.16
+ $Y2=0
r179 46 92 3.40825 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=10.25 $Y=0.085
+ $X2=10.372 $Y2=0
r180 46 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.25 $Y=0.085
+ $X2=10.25 $Y2=0.39
r181 42 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.36 $Y=0.085
+ $X2=9.36 $Y2=0
r182 42 44 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.36 $Y=0.085
+ $X2=9.36 $Y2=0.39
r183 38 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.54 $Y=0.085
+ $X2=6.54 $Y2=0
r184 38 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.54 $Y=0.085
+ $X2=6.54 $Y2=0.39
r185 37 55 32.5154 $w=2.78e-07 $l=7.9e-07 $layer=LI1_cond $X=2.245 $Y=0.785
+ $X2=3.035 $Y2=0.785
r186 33 37 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.16 $Y=0.645
+ $X2=2.245 $Y2=0.785
r187 33 35 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.16 $Y=0.645
+ $X2=2.16 $Y2=0.39
r188 32 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0
r189 32 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0.39
r190 28 89 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r191 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.39
r192 27 86 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r193 26 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.22
+ $Y2=0
r194 26 27 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=0
+ $X2=0.365 $Y2=0
r195 22 86 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r196 22 24 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.39
r197 7 48 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=10.115
+ $Y=0.235 $X2=10.25 $Y2=0.39
r198 6 44 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=9.175
+ $Y=0.235 $X2=9.36 $Y2=0.39
r199 5 40 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=6.355
+ $Y=0.235 $X2=6.54 $Y2=0.39
r200 4 54 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=2.985
+ $Y=0.235 $X2=3.12 $Y2=0.76
r201 3 35 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.16 $Y2=0.39
r202 2 30 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.235 $X2=1.22 $Y2=0.39
r203 1 24 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_4%A_503_47# 1 2 3 4 13 19 25 27 28
c36 27 0 1.43003e-19 $X=2.86 $Y=0.365
c37 19 0 1.71792e-19 $X=3.555 $Y=0.365
r38 27 28 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.86 $Y=0.34
+ $X2=3.335 $Y2=0.34
r39 23 25 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=5.08 $Y=0.365
+ $X2=6.02 $Y2=0.365
r40 21 23 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=4.14 $Y=0.365
+ $X2=5.08 $Y2=0.365
r41 19 28 12.1497 $w=2.18e-07 $l=2.2e-07 $layer=LI1_cond $X=3.555 $Y=0.365
+ $X2=3.335 $Y2=0.365
r42 19 21 30.6445 $w=2.18e-07 $l=5.85e-07 $layer=LI1_cond $X=3.555 $Y=0.365
+ $X2=4.14 $Y2=0.365
r43 13 27 6.3875 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=2.75 $Y=0.365
+ $X2=2.86 $Y2=0.365
r44 13 15 5.23838 $w=2.18e-07 $l=1e-07 $layer=LI1_cond $X=2.75 $Y=0.365 $X2=2.65
+ $Y2=0.365
r45 4 25 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.885
+ $Y=0.235 $X2=6.02 $Y2=0.39
r46 3 23 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.895
+ $Y=0.235 $X2=5.08 $Y2=0.39
r47 2 21 91 $w=1.7e-07 $l=7.58551e-07 $layer=licon1_NDIFF $count=2 $X=3.455
+ $Y=0.235 $X2=4.14 $Y2=0.39
r48 1 15 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.515
+ $Y=0.235 $X2=2.65 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A221OI_4%A_1375_47# 1 2 3 4 13 19 20 21 25
r49 23 25 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=9.805 $Y=0.725
+ $X2=9.805 $Y2=0.39
r50 22 30 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=9.055 $Y=0.815
+ $X2=8.93 $Y2=0.815
r51 21 23 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=9.615 $Y=0.815
+ $X2=9.805 $Y2=0.725
r52 21 22 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=9.615 $Y=0.815
+ $X2=9.055 $Y2=0.815
r53 20 30 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=8.93 $Y=0.725 $X2=8.93
+ $Y2=0.815
r54 19 28 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=8.93 $Y=0.475
+ $X2=8.93 $Y2=0.365
r55 19 20 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=8.93 $Y=0.475
+ $X2=8.93 $Y2=0.725
r56 15 18 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=7.01 $Y=0.365
+ $X2=7.95 $Y2=0.365
r57 13 28 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=8.805 $Y=0.365
+ $X2=8.93 $Y2=0.365
r58 13 18 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=8.805 $Y=0.365
+ $X2=7.95 $Y2=0.365
r59 4 25 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=9.645
+ $Y=0.235 $X2=9.83 $Y2=0.39
r60 3 30 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=8.755
+ $Y=0.235 $X2=8.89 $Y2=0.73
r61 3 28 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=8.755
+ $Y=0.235 $X2=8.89 $Y2=0.39
r62 2 18 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=7.765
+ $Y=0.235 $X2=7.95 $Y2=0.39
r63 1 15 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.875
+ $Y=0.235 $X2=7.01 $Y2=0.39
.ends

