* File: sky130_fd_sc_hdll__muxb4to1_2.pex.spice
* Created: Wed Sep  2 08:35:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%D[0] 3 7 11 15 17 27 29
r47 28 29 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.16
+ $X2=0.965 $Y2=1.16
r48 26 28 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=0.75 $Y=1.16 $X2=0.94
+ $Y2=1.16
r49 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.16 $X2=0.75 $Y2=1.16
r50 24 26 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=0.52 $Y=1.16 $X2=0.75
+ $Y2=1.16
r51 23 24 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r52 21 27 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.41 $Y=1.19
+ $X2=0.75 $Y2=1.19
r53 20 23 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=0.41 $Y=1.16
+ $X2=0.495 $Y2=1.16
r54 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r55 17 21 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.23 $Y=1.19
+ $X2=0.41 $Y2=1.19
r56 13 29 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=0.965 $Y=1.295
+ $X2=0.965 $Y2=1.16
r57 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.965 $Y=1.295
+ $X2=0.965 $Y2=1.985
r58 9 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.94 $Y=1.025
+ $X2=0.94 $Y2=1.16
r59 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.94 $Y=1.025
+ $X2=0.94 $Y2=0.56
r60 5 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=1.16
r61 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=0.56
r62 1 23 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=1.16
r63 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_278_265# 1 2 9 11 12 15 17 18 21 28
+ 32
c77 9 0 1.30521e-19 $X=1.49 $Y=2.075
r78 26 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=2.43 $Y=1.42
+ $X2=2.715 $Y2=1.63
r79 25 32 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=2.265 $Y=1.34
+ $X2=1.96 $Y2=1.34
r80 24 26 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=1.42
+ $X2=2.43 $Y2=1.42
r81 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.265
+ $Y=1.34 $X2=2.265 $Y2=1.34
r82 21 28 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.715 $Y=2.31
+ $X2=2.715 $Y2=1.635
r83 18 26 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.43 $Y=1.205
+ $X2=2.43 $Y2=1.42
r84 17 31 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=2.43 $Y=0.755
+ $X2=2.8 $Y2=0.457
r85 17 18 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.43 $Y=0.755
+ $X2=2.43 $Y2=1.205
r86 13 32 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=1.96 $Y=1.475
+ $X2=1.96 $Y2=1.34
r87 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=1.96 $Y=1.475 $X2=1.96
+ $Y2=2.075
r88 11 32 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=1.87 $Y=1.4
+ $X2=1.96 $Y2=1.34
r89 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.87 $Y=1.4 $X2=1.58
+ $Y2=1.4
r90 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.49 $Y=1.475
+ $X2=1.58 $Y2=1.4
r91 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=1.49 $Y=1.475 $X2=1.49
+ $Y2=2.075
r92 2 28 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.59
+ $Y=1.485 $X2=2.715 $Y2=1.63
r93 2 21 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=2.59
+ $Y=1.485 $X2=2.715 $Y2=2.31
r94 1 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=2.675
+ $Y=0.235 $X2=2.8 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%S[0] 1 3 4 5 6 8 9 12 13 14 15 17 18 20
+ 21 22
r65 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=2.955 $Y=0.92
+ $X2=2.955 $Y2=1.16
r66 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.955
+ $Y=1.16 $X2=2.955 $Y2=1.16
r67 18 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=3.01 $Y=0.845
+ $X2=2.955 $Y2=0.92
r68 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.01 $Y=0.845
+ $X2=3.01 $Y2=0.495
r69 15 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=2.95 $Y=1.41
+ $X2=2.955 $Y2=1.16
r70 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.95 $Y=1.41
+ $X2=2.95 $Y2=1.985
r71 13 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.82 $Y=0.92
+ $X2=2.955 $Y2=0.92
r72 13 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.82 $Y=0.92
+ $X2=2.44 $Y2=0.92
r73 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.365 $Y=0.845
+ $X2=2.44 $Y2=0.92
r74 11 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.365 $Y=0.255
+ $X2=2.365 $Y2=0.845
r75 10 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.955 $Y=0.18
+ $X2=1.88 $Y2=0.18
r76 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.29 $Y=0.18
+ $X2=2.365 $Y2=0.255
r77 9 10 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.29 $Y=0.18
+ $X2=1.955 $Y2=0.18
r78 6 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.88 $Y=0.255
+ $X2=1.88 $Y2=0.18
r79 6 8 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.88 $Y=0.255 $X2=1.88
+ $Y2=0.605
r80 4 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.805 $Y=0.18
+ $X2=1.88 $Y2=0.18
r81 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.805 $Y=0.18
+ $X2=1.535 $Y2=0.18
r82 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.46 $Y=0.255
+ $X2=1.535 $Y2=0.18
r83 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.46 $Y=0.255 $X2=1.46
+ $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%S[1] 1 3 4 6 7 10 11 12 13 15 16 18 20
+ 21 22
r62 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=3.485 $Y=0.92
+ $X2=3.485 $Y2=1.16
r63 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.485
+ $Y=1.16 $X2=3.485 $Y2=1.16
r64 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.98 $Y=0.255
+ $X2=4.98 $Y2=0.605
r65 17 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.635 $Y=0.18
+ $X2=4.56 $Y2=0.18
r66 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.905 $Y=0.18
+ $X2=4.98 $Y2=0.255
r67 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.905 $Y=0.18
+ $X2=4.635 $Y2=0.18
r68 13 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.56 $Y=0.255
+ $X2=4.56 $Y2=0.18
r69 13 15 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.56 $Y=0.255
+ $X2=4.56 $Y2=0.605
r70 11 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.485 $Y=0.18
+ $X2=4.56 $Y2=0.18
r71 11 12 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=4.485 $Y=0.18
+ $X2=4.15 $Y2=0.18
r72 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.075 $Y=0.255
+ $X2=4.15 $Y2=0.18
r73 9 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=4.075 $Y=0.255
+ $X2=4.075 $Y2=0.845
r74 8 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.62 $Y=0.92
+ $X2=3.485 $Y2=0.92
r75 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4 $Y=0.92
+ $X2=4.075 $Y2=0.845
r76 7 8 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=4 $Y=0.92 $X2=3.62
+ $Y2=0.92
r77 4 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=3.49 $Y=1.41
+ $X2=3.485 $Y2=1.16
r78 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.49 $Y=1.41 $X2=3.49
+ $Y2=1.985
r79 1 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=3.43 $Y=0.845
+ $X2=3.485 $Y2=0.92
r80 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.43 $Y=0.845 $X2=3.43
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_701_47# 1 2 9 11 12 15 19 22 24 28
c74 15 0 1.69024e-19 $X=4.95 $Y=2.075
c75 11 0 1.93373e-19 $X=4.86 $Y=1.4
r76 31 33 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=4.175 $Y=1.34
+ $X2=4.48 $Y2=1.34
r77 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.175
+ $Y=1.34 $X2=4.175 $Y2=1.34
r78 28 30 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.01 $Y=1.42
+ $X2=4.175 $Y2=1.42
r79 27 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=3.725 $Y=1.63
+ $X2=4.01 $Y2=1.42
r80 22 28 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=4.01 $Y=1.205
+ $X2=4.01 $Y2=1.42
r81 21 24 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=4.01 $Y=0.755
+ $X2=3.64 $Y2=0.457
r82 21 22 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.01 $Y=0.755
+ $X2=4.01 $Y2=1.205
r83 19 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.725 $Y=2.31
+ $X2=3.725 $Y2=1.635
r84 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=4.95 $Y=1.475 $X2=4.95
+ $Y2=2.075
r85 12 33 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=4.57 $Y=1.4
+ $X2=4.48 $Y2=1.34
r86 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.86 $Y=1.4
+ $X2=4.95 $Y2=1.475
r87 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.86 $Y=1.4 $X2=4.57
+ $Y2=1.4
r88 7 33 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=4.48 $Y=1.475
+ $X2=4.48 $Y2=1.34
r89 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=4.48 $Y=1.475 $X2=4.48
+ $Y2=2.075
r90 2 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=1.485 $X2=3.725 $Y2=1.63
r91 2 19 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=1.485 $X2=3.725 $Y2=2.31
r92 1 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=3.505
+ $Y=0.235 $X2=3.64 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%D[1] 3 7 11 15 17 28
c53 17 0 1.17966e-19 $X=6.21 $Y=1.19
c54 15 0 1.17966e-19 $X=5.945 $Y=1.985
r55 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.03
+ $Y=1.16 $X2=6.03 $Y2=1.16
r56 26 28 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=5.945 $Y=1.16
+ $X2=6.03 $Y2=1.16
r57 25 26 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.92 $Y=1.16
+ $X2=5.945 $Y2=1.16
r58 24 29 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.69 $Y=1.19
+ $X2=6.03 $Y2=1.19
r59 23 25 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=5.69 $Y=1.16 $X2=5.92
+ $Y2=1.16
r60 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.69
+ $Y=1.16 $X2=5.69 $Y2=1.16
r61 21 23 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=5.5 $Y=1.16 $X2=5.69
+ $Y2=1.16
r62 19 21 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.475 $Y=1.16
+ $X2=5.5 $Y2=1.16
r63 17 29 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.21 $Y=1.19
+ $X2=6.03 $Y2=1.19
r64 13 26 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.945 $Y=1.295
+ $X2=5.945 $Y2=1.16
r65 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=5.945 $Y=1.295
+ $X2=5.945 $Y2=1.985
r66 9 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.92 $Y=1.025
+ $X2=5.92 $Y2=1.16
r67 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.92 $Y=1.025
+ $X2=5.92 $Y2=0.56
r68 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.5 $Y=1.025 $X2=5.5
+ $Y2=1.16
r69 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.5 $Y=1.025 $X2=5.5
+ $Y2=0.56
r70 1 19 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.475 $Y=1.295
+ $X2=5.475 $Y2=1.16
r71 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=5.475 $Y=1.295
+ $X2=5.475 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%D[2] 3 7 11 15 17 27 29
c54 27 0 1.17966e-19 $X=7.19 $Y=1.16
c55 3 0 1.17966e-19 $X=6.935 $Y=1.985
r56 28 29 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=7.38 $Y=1.16
+ $X2=7.405 $Y2=1.16
r57 26 28 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=7.19 $Y=1.16 $X2=7.38
+ $Y2=1.16
r58 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.19
+ $Y=1.16 $X2=7.19 $Y2=1.16
r59 24 26 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=6.96 $Y=1.16 $X2=7.19
+ $Y2=1.16
r60 23 24 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=6.935 $Y=1.16
+ $X2=6.96 $Y2=1.16
r61 21 27 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.85 $Y=1.19
+ $X2=7.19 $Y2=1.19
r62 20 23 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=6.85 $Y=1.16
+ $X2=6.935 $Y2=1.16
r63 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.85
+ $Y=1.16 $X2=6.85 $Y2=1.16
r64 17 21 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.67 $Y=1.19
+ $X2=6.85 $Y2=1.19
r65 13 29 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=7.405 $Y=1.295
+ $X2=7.405 $Y2=1.16
r66 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=7.405 $Y=1.295
+ $X2=7.405 $Y2=1.985
r67 9 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.38 $Y=1.025
+ $X2=7.38 $Y2=1.16
r68 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.38 $Y=1.025
+ $X2=7.38 $Y2=0.56
r69 5 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.96 $Y=1.025
+ $X2=6.96 $Y2=1.16
r70 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.96 $Y=1.025
+ $X2=6.96 $Y2=0.56
r71 1 23 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=6.935 $Y=1.295
+ $X2=6.935 $Y2=1.16
r72 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=6.935 $Y=1.295
+ $X2=6.935 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_1566_265# 1 2 9 11 12 15 17 18 21 28
+ 32
c78 12 0 1.93373e-19 $X=8.02 $Y=1.4
c79 9 0 1.69024e-19 $X=7.93 $Y=2.075
r80 26 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=8.87 $Y=1.42
+ $X2=9.155 $Y2=1.63
r81 25 32 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=8.705 $Y=1.34
+ $X2=8.4 $Y2=1.34
r82 24 26 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=8.705 $Y=1.42
+ $X2=8.87 $Y2=1.42
r83 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.705
+ $Y=1.34 $X2=8.705 $Y2=1.34
r84 21 28 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=9.155 $Y=2.31
+ $X2=9.155 $Y2=1.635
r85 18 26 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=8.87 $Y=1.205
+ $X2=8.87 $Y2=1.42
r86 17 31 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=8.87 $Y=0.755
+ $X2=9.24 $Y2=0.457
r87 17 18 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.87 $Y=0.755
+ $X2=8.87 $Y2=1.205
r88 13 32 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=8.4 $Y=1.475
+ $X2=8.4 $Y2=1.34
r89 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=8.4 $Y=1.475 $X2=8.4
+ $Y2=2.075
r90 11 32 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=8.31 $Y=1.4
+ $X2=8.4 $Y2=1.34
r91 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.31 $Y=1.4 $X2=8.02
+ $Y2=1.4
r92 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=7.93 $Y=1.475
+ $X2=8.02 $Y2=1.4
r93 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=7.93 $Y=1.475 $X2=7.93
+ $Y2=2.075
r94 2 28 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=9.03
+ $Y=1.485 $X2=9.155 $Y2=1.63
r95 2 21 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=9.03
+ $Y=1.485 $X2=9.155 $Y2=2.31
r96 1 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=9.115
+ $Y=0.235 $X2=9.24 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%S[2] 1 3 4 5 6 8 9 12 13 14 15 17 18 20
+ 21 22
r65 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=9.395 $Y=0.92
+ $X2=9.395 $Y2=1.16
r66 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.395
+ $Y=1.16 $X2=9.395 $Y2=1.16
r67 18 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=9.45 $Y=0.845
+ $X2=9.395 $Y2=0.92
r68 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.45 $Y=0.845
+ $X2=9.45 $Y2=0.495
r69 15 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=9.39 $Y=1.41
+ $X2=9.395 $Y2=1.16
r70 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.39 $Y=1.41
+ $X2=9.39 $Y2=1.985
r71 13 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.26 $Y=0.92
+ $X2=9.395 $Y2=0.92
r72 13 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=9.26 $Y=0.92
+ $X2=8.88 $Y2=0.92
r73 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.805 $Y=0.845
+ $X2=8.88 $Y2=0.92
r74 11 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=8.805 $Y=0.255
+ $X2=8.805 $Y2=0.845
r75 10 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.395 $Y=0.18
+ $X2=8.32 $Y2=0.18
r76 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.73 $Y=0.18
+ $X2=8.805 $Y2=0.255
r77 9 10 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=8.73 $Y=0.18
+ $X2=8.395 $Y2=0.18
r78 6 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.32 $Y=0.255
+ $X2=8.32 $Y2=0.18
r79 6 8 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=8.32 $Y=0.255 $X2=8.32
+ $Y2=0.605
r80 4 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.245 $Y=0.18
+ $X2=8.32 $Y2=0.18
r81 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.245 $Y=0.18
+ $X2=7.975 $Y2=0.18
r82 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.9 $Y=0.255
+ $X2=7.975 $Y2=0.18
r83 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=7.9 $Y=0.255 $X2=7.9
+ $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%S[3] 1 3 4 6 7 10 11 12 13 15 16 18 20
+ 21 22
r62 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=9.925 $Y=0.92
+ $X2=9.925 $Y2=1.16
r63 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.925
+ $Y=1.16 $X2=9.925 $Y2=1.16
r64 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=11.42 $Y=0.255
+ $X2=11.42 $Y2=0.605
r65 17 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.075 $Y=0.18
+ $X2=11 $Y2=0.18
r66 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.345 $Y=0.18
+ $X2=11.42 $Y2=0.255
r67 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=11.345 $Y=0.18
+ $X2=11.075 $Y2=0.18
r68 13 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11 $Y=0.255 $X2=11
+ $Y2=0.18
r69 13 15 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=11 $Y=0.255 $X2=11
+ $Y2=0.605
r70 11 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.925 $Y=0.18
+ $X2=11 $Y2=0.18
r71 11 12 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.925 $Y=0.18
+ $X2=10.59 $Y2=0.18
r72 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.515 $Y=0.255
+ $X2=10.59 $Y2=0.18
r73 9 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=10.515 $Y=0.255
+ $X2=10.515 $Y2=0.845
r74 8 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.06 $Y=0.92
+ $X2=9.925 $Y2=0.92
r75 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.44 $Y=0.92
+ $X2=10.515 $Y2=0.845
r76 7 8 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=10.44 $Y=0.92
+ $X2=10.06 $Y2=0.92
r77 4 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=9.93 $Y=1.41
+ $X2=9.925 $Y2=1.16
r78 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.93 $Y=1.41 $X2=9.93
+ $Y2=1.985
r79 1 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=9.87 $Y=0.845
+ $X2=9.925 $Y2=0.92
r80 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.87 $Y=0.845 $X2=9.87
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_1989_47# 1 2 9 11 12 15 19 22 24 28
c73 15 0 1.30521e-19 $X=11.39 $Y=2.075
r74 31 33 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=10.615 $Y=1.34
+ $X2=10.92 $Y2=1.34
r75 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.615
+ $Y=1.34 $X2=10.615 $Y2=1.34
r76 28 30 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=10.45 $Y=1.42
+ $X2=10.615 $Y2=1.42
r77 27 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=10.165 $Y=1.63
+ $X2=10.45 $Y2=1.42
r78 22 28 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=10.45 $Y=1.205
+ $X2=10.45 $Y2=1.42
r79 21 24 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=10.45 $Y=0.755
+ $X2=10.08 $Y2=0.457
r80 21 22 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=10.45 $Y=0.755
+ $X2=10.45 $Y2=1.205
r81 19 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=10.165 $Y=2.31
+ $X2=10.165 $Y2=1.635
r82 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=11.39 $Y=1.475
+ $X2=11.39 $Y2=2.075
r83 12 33 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=11.01 $Y=1.4
+ $X2=10.92 $Y2=1.34
r84 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=11.3 $Y=1.4
+ $X2=11.39 $Y2=1.475
r85 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=11.3 $Y=1.4
+ $X2=11.01 $Y2=1.4
r86 7 33 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=10.92 $Y=1.475
+ $X2=10.92 $Y2=1.34
r87 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=10.92 $Y=1.475 $X2=10.92
+ $Y2=2.075
r88 2 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.02
+ $Y=1.485 $X2=10.165 $Y2=1.63
r89 2 19 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=10.02
+ $Y=1.485 $X2=10.165 $Y2=2.31
r90 1 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=9.945
+ $Y=0.235 $X2=10.08 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%D[3] 3 7 11 15 17 28
r46 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.47
+ $Y=1.16 $X2=12.47 $Y2=1.16
r47 26 28 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=12.385 $Y=1.16
+ $X2=12.47 $Y2=1.16
r48 25 26 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=12.36 $Y=1.16
+ $X2=12.385 $Y2=1.16
r49 24 29 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=12.13 $Y=1.19
+ $X2=12.47 $Y2=1.19
r50 23 25 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=12.13 $Y=1.16 $X2=12.36
+ $Y2=1.16
r51 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.13
+ $Y=1.16 $X2=12.13 $Y2=1.16
r52 21 23 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=11.94 $Y=1.16
+ $X2=12.13 $Y2=1.16
r53 19 21 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=11.915 $Y=1.16
+ $X2=11.94 $Y2=1.16
r54 17 29 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=12.65 $Y=1.19
+ $X2=12.47 $Y2=1.19
r55 13 26 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=12.385 $Y=1.295
+ $X2=12.385 $Y2=1.16
r56 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=12.385 $Y=1.295
+ $X2=12.385 $Y2=1.985
r57 9 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=12.36 $Y=1.025
+ $X2=12.36 $Y2=1.16
r58 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=12.36 $Y=1.025
+ $X2=12.36 $Y2=0.56
r59 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.94 $Y=1.025
+ $X2=11.94 $Y2=1.16
r60 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.94 $Y=1.025
+ $X2=11.94 $Y2=0.56
r61 1 19 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=11.915 $Y=1.295
+ $X2=11.915 $Y2=1.16
r62 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=11.915 $Y=1.295
+ $X2=11.915 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_27_297# 1 2 3 10 12 17 18 19 22 27 28
r47 27 28 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.26 $Y=2.34
+ $X2=0.26 $Y2=2.21
r48 20 22 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.195 $Y=2.295
+ $X2=2.195 $Y2=1.81
r49 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.11 $Y=2.38
+ $X2=2.195 $Y2=2.295
r50 18 19 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=2.11 $Y=2.38
+ $X2=1.285 $Y2=2.38
r51 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.2 $Y=2.295
+ $X2=1.285 $Y2=2.38
r52 15 17 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=1.2 $Y=2.295
+ $X2=1.2 $Y2=1.78
r53 14 17 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.665
+ $X2=1.2 $Y2=1.78
r54 13 25 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.395 $Y=1.58
+ $X2=0.245 $Y2=1.58
r55 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.115 $Y=1.58
+ $X2=1.2 $Y2=1.665
r56 12 13 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.115 $Y=1.58
+ $X2=0.395 $Y2=1.58
r57 10 25 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=1.665
+ $X2=0.245 $Y2=1.58
r58 10 28 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=0.245 $Y=1.665
+ $X2=0.245 $Y2=2.21
r59 3 22 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=2.05
+ $Y=1.665 $X2=2.195 $Y2=1.81
r60 2 17 300 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.78
r61 1 27 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r62 1 25 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%VPWR 1 2 3 4 5 6 22 25 32 36 39 46 48
+ 52 53 55 59 63 64 66 69 70 71 72 77 89 96 108 117 121 124 127 130
c182 66 0 1.30521e-19 $X=12.15 $Y=1.94
c183 59 0 1.69024e-19 $X=7.17 $Y=1.94
c184 55 0 1.69024e-19 $X=5.71 $Y=1.94
c185 48 0 1.30521e-19 $X=0.73 $Y=1.94
r186 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r187 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r188 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r189 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r190 115 130 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=12.285 $Y=2.72
+ $X2=12.135 $Y2=2.72
r191 115 117 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=12.285 $Y=2.72
+ $X2=12.65 $Y2=2.72
r192 114 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=12.19 $Y2=2.72
r193 113 114 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r194 111 114 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=11.73 $Y2=2.72
r195 110 113 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=9.89 $Y=2.72
+ $X2=11.73 $Y2=2.72
r196 110 111 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r197 108 130 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=11.985 $Y=2.72
+ $X2=12.135 $Y2=2.72
r198 108 113 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.985 $Y=2.72
+ $X2=11.73 $Y2=2.72
r199 107 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=9.89 $Y2=2.72
r200 106 107 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r201 104 107 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=9.43 $Y2=2.72
r202 104 128 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r203 103 106 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=7.59 $Y=2.72
+ $X2=9.43 $Y2=2.72
r204 103 104 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r205 101 127 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=7.335 $Y=2.72
+ $X2=7.185 $Y2=2.72
r206 101 103 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.335 $Y=2.72
+ $X2=7.59 $Y2=2.72
r207 97 124 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.845 $Y=2.72
+ $X2=5.695 $Y2=2.72
r208 97 99 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=5.845 $Y=2.72
+ $X2=6.67 $Y2=2.72
r209 96 127 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=7.035 $Y=2.72
+ $X2=7.185 $Y2=2.72
r210 96 99 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.035 $Y=2.72
+ $X2=6.67 $Y2=2.72
r211 95 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r212 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r213 92 95 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=5.29 $Y2=2.72
r214 91 94 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=5.29 $Y2=2.72
r215 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r216 89 124 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.545 $Y=2.72
+ $X2=5.695 $Y2=2.72
r217 89 94 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.545 $Y=2.72
+ $X2=5.29 $Y2=2.72
r218 88 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r219 87 88 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r220 85 88 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r221 85 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r222 84 87 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r223 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r224 82 121 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.745 $Y2=2.72
r225 82 84 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r226 77 121 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.745 $Y2=2.72
r227 77 79 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r228 72 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=12.19 $Y2=2.72
r229 72 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r230 71 128 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r231 71 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r232 70 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r233 70 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r234 69 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r235 69 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r236 66 68 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.15 $Y=1.94
+ $X2=12.15 $Y2=2.105
r237 63 106 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=9.495 $Y=2.72
+ $X2=9.43 $Y2=2.72
r238 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.495 $Y=2.72
+ $X2=9.66 $Y2=2.72
r239 62 110 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=9.825 $Y=2.72
+ $X2=9.89 $Y2=2.72
r240 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.825 $Y=2.72
+ $X2=9.66 $Y2=2.72
r241 59 61 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.17 $Y=1.94
+ $X2=7.17 $Y2=2.105
r242 55 57 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.71 $Y=1.94
+ $X2=5.71 $Y2=2.105
r243 52 87 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.055 $Y=2.72
+ $X2=2.99 $Y2=2.72
r244 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.055 $Y=2.72
+ $X2=3.22 $Y2=2.72
r245 51 91 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.385 $Y=2.72
+ $X2=3.45 $Y2=2.72
r246 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=2.72
+ $X2=3.22 $Y2=2.72
r247 48 50 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=1.94
+ $X2=0.73 $Y2=2.105
r248 46 68 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=12.135 $Y=2.34
+ $X2=12.135 $Y2=2.105
r249 44 130 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.135 $Y=2.635
+ $X2=12.135 $Y2=2.72
r250 44 46 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=12.135 $Y=2.635
+ $X2=12.135 $Y2=2.34
r251 39 42 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.66 $Y=1.63
+ $X2=9.66 $Y2=2.31
r252 37 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.66 $Y=2.635
+ $X2=9.66 $Y2=2.72
r253 37 42 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=9.66 $Y=2.635
+ $X2=9.66 $Y2=2.31
r254 36 61 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=7.185 $Y=2.34
+ $X2=7.185 $Y2=2.105
r255 34 127 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.185 $Y=2.635
+ $X2=7.185 $Y2=2.72
r256 34 36 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=7.185 $Y=2.635
+ $X2=7.185 $Y2=2.34
r257 32 57 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=5.695 $Y=2.34
+ $X2=5.695 $Y2=2.105
r258 30 124 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.695 $Y=2.635
+ $X2=5.695 $Y2=2.72
r259 30 32 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=5.695 $Y=2.635
+ $X2=5.695 $Y2=2.34
r260 25 28 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.22 $Y=1.63
+ $X2=3.22 $Y2=2.31
r261 23 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=2.635
+ $X2=3.22 $Y2=2.72
r262 23 28 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.22 $Y=2.635
+ $X2=3.22 $Y2=2.31
r263 22 50 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=0.745 $Y=2.34
+ $X2=0.745 $Y2=2.105
r264 20 121 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=2.635
+ $X2=0.745 $Y2=2.72
r265 20 22 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.745 $Y=2.635
+ $X2=0.745 $Y2=2.34
r266 6 66 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=12.005
+ $Y=1.485 $X2=12.15 $Y2=1.94
r267 6 46 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=12.005
+ $Y=1.485 $X2=12.15 $Y2=2.34
r268 5 42 400 $w=1.7e-07 $l=9.10563e-07 $layer=licon1_PDIFF $count=1 $X=9.48
+ $Y=1.485 $X2=9.66 $Y2=2.31
r269 5 39 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=9.48
+ $Y=1.485 $X2=9.66 $Y2=1.63
r270 4 59 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=7.025
+ $Y=1.485 $X2=7.17 $Y2=1.94
r271 4 36 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.025
+ $Y=1.485 $X2=7.17 $Y2=2.34
r272 3 55 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=1.485 $X2=5.71 $Y2=1.94
r273 3 32 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=1.485 $X2=5.71 $Y2=2.34
r274 2 28 400 $w=1.7e-07 $l=9.10563e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=1.485 $X2=3.22 $Y2=2.31
r275 2 25 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=1.485 $X2=3.22 $Y2=1.63
r276 1 48 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.94
r277 1 22 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%Z 1 2 3 4 5 6 7 8 34 37 40 43 45 46 47
+ 48 49 50 51 52 53 54 60 62 66 68 72 74 78 80
c228 47 0 6.32252e-19 $X=7.905 $Y=1.87
r229 78 80 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=11.2 $Y=1.87
+ $X2=11.2 $Y2=1.755
r230 72 74 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=8.12 $Y=1.87
+ $X2=8.12 $Y2=1.755
r231 66 68 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.76 $Y=1.87
+ $X2=4.76 $Y2=1.755
r232 60 62 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.87
+ $X2=1.68 $Y2=1.755
r233 54 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=1.87
+ $X2=11.27 $Y2=1.87
r234 53 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=1.87
+ $X2=8.05 $Y2=1.87
r235 52 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=1.87
+ $X2=4.83 $Y2=1.87
r236 51 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=1.87
+ $X2=1.61 $Y2=1.87
r237 50 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.195 $Y=1.87
+ $X2=8.05 $Y2=1.87
r238 49 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.125 $Y=1.87
+ $X2=11.27 $Y2=1.87
r239 49 50 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=11.125 $Y=1.87
+ $X2=8.195 $Y2=1.87
r240 48 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.975 $Y=1.87
+ $X2=4.83 $Y2=1.87
r241 47 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.905 $Y=1.87
+ $X2=8.05 $Y2=1.87
r242 47 48 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=7.905 $Y=1.87
+ $X2=4.975 $Y2=1.87
r243 46 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.755 $Y=1.87
+ $X2=1.61 $Y2=1.87
r244 45 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.685 $Y=1.87
+ $X2=4.83 $Y2=1.87
r245 45 46 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=4.685 $Y=1.87
+ $X2=1.755 $Y2=1.87
r246 31 43 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=11.21 $Y=0.885
+ $X2=11.21 $Y2=0.68
r247 31 80 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=11.21 $Y=0.885
+ $X2=11.21 $Y2=1.755
r248 29 40 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=8.11 $Y=0.885
+ $X2=8.11 $Y2=0.68
r249 29 74 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=8.11 $Y=0.885
+ $X2=8.11 $Y2=1.755
r250 27 37 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=4.77 $Y=0.885
+ $X2=4.77 $Y2=0.68
r251 27 68 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=4.77 $Y=0.885
+ $X2=4.77 $Y2=1.755
r252 25 34 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.67 $Y=0.885
+ $X2=1.67 $Y2=0.68
r253 25 62 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=1.67 $Y=0.885
+ $X2=1.67 $Y2=1.755
r254 8 78 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=11.01
+ $Y=1.665 $X2=11.155 $Y2=2.02
r255 7 72 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=8.02
+ $Y=1.665 $X2=8.165 $Y2=2.02
r256 6 66 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=4.57
+ $Y=1.665 $X2=4.715 $Y2=2.02
r257 5 60 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.665 $X2=1.725 $Y2=2.02
r258 4 43 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=11.075
+ $Y=0.345 $X2=11.21 $Y2=0.68
r259 3 40 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=7.975
+ $Y=0.345 $X2=8.11 $Y2=0.68
r260 2 37 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=4.635
+ $Y=0.345 $X2=4.77 $Y2=0.68
r261 1 34 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.345 $X2=1.67 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_824_333# 1 2 3 12 14 15 19 20 21 22
+ 25 26
c59 3 0 1.22753e-19 $X=6.035 $Y=1.485
r60 25 26 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=6.18 $Y=2.34
+ $X2=6.18 $Y2=2.21
r61 22 29 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.195 $Y=1.665
+ $X2=6.195 $Y2=1.58
r62 22 26 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=6.195 $Y=1.665
+ $X2=6.195 $Y2=2.21
r63 20 29 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.045 $Y=1.58
+ $X2=6.195 $Y2=1.58
r64 20 21 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.045 $Y=1.58
+ $X2=5.325 $Y2=1.58
r65 17 19 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=5.24 $Y=2.295
+ $X2=5.24 $Y2=1.78
r66 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.24 $Y=1.665
+ $X2=5.325 $Y2=1.58
r67 16 19 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=5.24 $Y=1.665
+ $X2=5.24 $Y2=1.78
r68 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.155 $Y=2.38
+ $X2=5.24 $Y2=2.295
r69 14 15 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=5.155 $Y=2.38
+ $X2=4.33 $Y2=2.38
r70 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.245 $Y=2.295
+ $X2=4.33 $Y2=2.38
r71 10 12 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.245 $Y=2.295
+ $X2=4.245 $Y2=1.81
r72 3 29 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=6.035
+ $Y=1.485 $X2=6.18 $Y2=1.66
r73 3 25 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.035
+ $Y=1.485 $X2=6.18 $Y2=2.34
r74 2 19 300 $w=1.7e-07 $l=2.50998e-07 $layer=licon1_PDIFF $count=2 $X=5.04
+ $Y=1.665 $X2=5.24 $Y2=1.78
r75 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=4.12
+ $Y=1.665 $X2=4.245 $Y2=1.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_1315_297# 1 2 3 10 12 17 18 19 22 27
+ 28
c57 1 0 1.22753e-19 $X=6.575 $Y=1.485
r58 27 28 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=6.7 $Y=2.34 $X2=6.7
+ $Y2=2.21
r59 20 22 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=8.635 $Y=2.295
+ $X2=8.635 $Y2=1.81
r60 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.55 $Y=2.38
+ $X2=8.635 $Y2=2.295
r61 18 19 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=8.55 $Y=2.38
+ $X2=7.725 $Y2=2.38
r62 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.64 $Y=2.295
+ $X2=7.725 $Y2=2.38
r63 15 17 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=7.64 $Y=2.295
+ $X2=7.64 $Y2=1.78
r64 14 17 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.64 $Y=1.665
+ $X2=7.64 $Y2=1.78
r65 13 25 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.835 $Y=1.58
+ $X2=6.685 $Y2=1.58
r66 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.555 $Y=1.58
+ $X2=7.64 $Y2=1.665
r67 12 13 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=7.555 $Y=1.58
+ $X2=6.835 $Y2=1.58
r68 10 25 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.685 $Y=1.665
+ $X2=6.685 $Y2=1.58
r69 10 28 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=6.685 $Y=1.665
+ $X2=6.685 $Y2=2.21
r70 3 22 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=8.49
+ $Y=1.665 $X2=8.635 $Y2=1.81
r71 2 17 300 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=2 $X=7.495
+ $Y=1.485 $X2=7.64 $Y2=1.78
r72 1 27 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=6.575
+ $Y=1.485 $X2=6.7 $Y2=2.34
r73 1 25 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=6.575
+ $Y=1.485 $X2=6.7 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_2112_333# 1 2 3 12 14 15 19 20 21 22
+ 25 26
r49 25 26 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=12.62 $Y=2.34
+ $X2=12.62 $Y2=2.21
r50 22 29 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.635 $Y=1.665
+ $X2=12.635 $Y2=1.58
r51 22 26 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=12.635 $Y=1.665
+ $X2=12.635 $Y2=2.21
r52 20 29 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=12.485 $Y=1.58
+ $X2=12.635 $Y2=1.58
r53 20 21 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=12.485 $Y=1.58
+ $X2=11.765 $Y2=1.58
r54 17 19 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=11.68 $Y=2.295
+ $X2=11.68 $Y2=1.78
r55 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.68 $Y=1.665
+ $X2=11.765 $Y2=1.58
r56 16 19 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=11.68 $Y=1.665
+ $X2=11.68 $Y2=1.78
r57 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.595 $Y=2.38
+ $X2=11.68 $Y2=2.295
r58 14 15 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=11.595 $Y=2.38
+ $X2=10.77 $Y2=2.38
r59 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.685 $Y=2.295
+ $X2=10.77 $Y2=2.38
r60 10 12 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=10.685 $Y=2.295
+ $X2=10.685 $Y2=1.81
r61 3 29 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=12.475
+ $Y=1.485 $X2=12.62 $Y2=1.66
r62 3 25 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=12.475
+ $Y=1.485 $X2=12.62 $Y2=2.34
r63 2 19 300 $w=1.7e-07 $l=2.50998e-07 $layer=licon1_PDIFF $count=2 $X=11.48
+ $Y=1.665 $X2=11.68 $Y2=1.78
r64 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=10.56
+ $Y=1.665 $X2=10.685 $Y2=1.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_27_47# 1 2 3 12 14 15 16 18 22
c42 16 0 1.81988e-19 $X=1.182 $Y=0.425
r43 20 22 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.09 $Y=0.425
+ $X2=2.09 $Y2=0.605
r44 19 25 4.85887 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.335 $Y=0.34
+ $X2=1.182 $Y2=0.34
r45 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.005 $Y=0.34
+ $X2=2.09 $Y2=0.425
r46 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=0.34
+ $X2=1.335 $Y2=0.34
r47 16 25 2.69937 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.182 $Y=0.425
+ $X2=1.182 $Y2=0.34
r48 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=1.182 $Y=0.425
+ $X2=1.182 $Y2=0.715
r49 14 17 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=1.03 $Y=0.8
+ $X2=1.182 $Y2=0.715
r50 14 15 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.03 $Y=0.8
+ $X2=0.475 $Y2=0.8
r51 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.31 $Y=0.715
+ $X2=0.475 $Y2=0.8
r52 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.31 $Y=0.715
+ $X2=0.31 $Y2=0.38
r53 3 22 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.345 $X2=2.09 $Y2=0.605
r54 2 25 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.235 $X2=1.175 $Y2=0.42
r55 1 12 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.31 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%VGND 1 2 3 4 5 6 23 27 31 33 37 41 45
+ 48 49 51 52 54 55 56 57 58 59 71 92 96 99 102
r143 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r144 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r145 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r146 89 90 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r147 87 90 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=11.73 $Y2=0
r148 86 89 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=9.89 $Y=0
+ $X2=11.73 $Y2=0
r149 86 87 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r150 84 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0 $X2=9.89
+ $Y2=0
r151 83 84 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r152 81 84 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=9.43 $Y2=0
r153 81 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=7.13 $Y2=0
r154 80 83 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=7.59 $Y=0 $X2=9.43
+ $Y2=0
r155 80 81 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r156 78 102 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=7.3 $Y=0 $X2=7.192
+ $Y2=0
r157 78 80 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.3 $Y=0 $X2=7.59
+ $Y2=0
r158 77 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=5.75 $Y2=0
r159 76 77 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r160 74 77 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=5.29 $Y2=0
r161 73 76 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=3.45 $Y=0 $X2=5.29
+ $Y2=0
r162 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r163 71 99 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=5.58 $Y=0 $X2=5.687
+ $Y2=0
r164 71 76 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.58 $Y=0 $X2=5.29
+ $Y2=0
r165 70 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r166 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r167 67 70 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.99 $Y2=0
r168 67 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r169 66 69 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r170 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r171 64 96 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=0.86 $Y=0 $X2=0.752
+ $Y2=0
r172 64 66 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.86 $Y=0 $X2=1.15
+ $Y2=0
r173 59 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=11.73 $Y2=0
r174 59 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r175 58 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r176 57 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r177 57 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=5.75 $Y2=0
r178 56 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r179 54 89 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=12.02 $Y=0
+ $X2=11.73 $Y2=0
r180 54 55 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=12.02 $Y=0
+ $X2=12.127 $Y2=0
r181 53 92 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=12.235 $Y=0
+ $X2=12.65 $Y2=0
r182 53 55 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=12.235 $Y=0
+ $X2=12.127 $Y2=0
r183 51 83 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=9.535 $Y=0
+ $X2=9.43 $Y2=0
r184 51 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.535 $Y=0 $X2=9.66
+ $Y2=0
r185 50 86 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=9.785 $Y=0
+ $X2=9.89 $Y2=0
r186 50 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.785 $Y=0 $X2=9.66
+ $Y2=0
r187 48 69 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.095 $Y=0
+ $X2=2.99 $Y2=0
r188 48 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.095 $Y=0 $X2=3.22
+ $Y2=0
r189 47 73 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.345 $Y=0
+ $X2=3.45 $Y2=0
r190 47 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.345 $Y=0 $X2=3.22
+ $Y2=0
r191 43 55 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=12.127 $Y=0.085
+ $X2=12.127 $Y2=0
r192 43 45 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=12.127 $Y=0.085
+ $X2=12.127 $Y2=0.38
r193 39 52 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.66 $Y=0.085
+ $X2=9.66 $Y2=0
r194 39 41 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=9.66 $Y=0.085
+ $X2=9.66 $Y2=0.495
r195 35 102 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=7.192 $Y=0.085
+ $X2=7.192 $Y2=0
r196 35 37 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=7.192 $Y=0.085
+ $X2=7.192 $Y2=0.38
r197 34 99 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=5.795 $Y=0
+ $X2=5.687 $Y2=0
r198 33 102 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=7.085 $Y=0
+ $X2=7.192 $Y2=0
r199 33 34 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=7.085 $Y=0
+ $X2=5.795 $Y2=0
r200 29 99 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.687 $Y=0.085
+ $X2=5.687 $Y2=0
r201 29 31 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=5.687 $Y=0.085
+ $X2=5.687 $Y2=0.38
r202 25 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=0.085
+ $X2=3.22 $Y2=0
r203 25 27 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=3.22 $Y=0.085
+ $X2=3.22 $Y2=0.495
r204 21 96 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.752 $Y=0.085
+ $X2=0.752 $Y2=0
r205 21 23 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=0.752 $Y=0.085
+ $X2=0.752 $Y2=0.38
r206 6 45 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=12.015
+ $Y=0.235 $X2=12.15 $Y2=0.38
r207 5 41 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=9.525
+ $Y=0.235 $X2=9.66 $Y2=0.495
r208 4 37 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.035
+ $Y=0.235 $X2=7.17 $Y2=0.38
r209 3 31 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.575
+ $Y=0.235 $X2=5.71 $Y2=0.38
r210 2 27 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=3.085
+ $Y=0.235 $X2=3.22 $Y2=0.495
r211 1 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_845_69# 1 2 3 12 14 15 16 18 19 22
c48 16 0 1.81988e-19 $X=5.257 $Y=0.425
r49 20 22 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.13 $Y=0.715
+ $X2=6.13 $Y2=0.38
r50 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.965 $Y=0.8
+ $X2=6.13 $Y2=0.715
r51 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=5.965 $Y=0.8
+ $X2=5.41 $Y2=0.8
r52 17 19 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=5.257 $Y=0.715
+ $X2=5.41 $Y2=0.8
r53 16 25 2.71076 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.257 $Y=0.425
+ $X2=5.257 $Y2=0.34
r54 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=5.257 $Y=0.425
+ $X2=5.257 $Y2=0.715
r55 14 25 4.84748 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.105 $Y=0.34
+ $X2=5.257 $Y2=0.34
r56 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.105 $Y=0.34
+ $X2=4.435 $Y2=0.34
r57 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.35 $Y=0.425
+ $X2=4.435 $Y2=0.34
r58 10 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.35 $Y=0.425
+ $X2=4.35 $Y2=0.605
r59 3 22 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.995
+ $Y=0.235 $X2=6.13 $Y2=0.38
r60 2 25 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=5.055
+ $Y=0.345 $X2=5.265 $Y2=0.42
r61 1 12 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=4.225
+ $Y=0.345 $X2=4.35 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_1315_47# 1 2 3 12 14 15 16 18 22
c44 16 0 1.81988e-19 $X=7.622 $Y=0.425
r45 20 22 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.53 $Y=0.425
+ $X2=8.53 $Y2=0.605
r46 19 25 4.85887 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.775 $Y=0.34
+ $X2=7.622 $Y2=0.34
r47 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.445 $Y=0.34
+ $X2=8.53 $Y2=0.425
r48 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.445 $Y=0.34
+ $X2=7.775 $Y2=0.34
r49 16 25 2.69937 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.622 $Y=0.425
+ $X2=7.622 $Y2=0.34
r50 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=7.622 $Y=0.425
+ $X2=7.622 $Y2=0.715
r51 14 17 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=7.47 $Y=0.8
+ $X2=7.622 $Y2=0.715
r52 14 15 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=7.47 $Y=0.8
+ $X2=6.915 $Y2=0.8
r53 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.75 $Y=0.715
+ $X2=6.915 $Y2=0.8
r54 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.75 $Y=0.715
+ $X2=6.75 $Y2=0.38
r55 3 22 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=8.395
+ $Y=0.345 $X2=8.53 $Y2=0.605
r56 2 25 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=7.455
+ $Y=0.235 $X2=7.615 $Y2=0.42
r57 1 12 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=6.575
+ $Y=0.235 $X2=6.75 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_2%A_2133_69# 1 2 3 12 14 15 16 18 19 22
c46 16 0 1.81988e-19 $X=11.697 $Y=0.425
r47 20 22 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=12.57 $Y=0.715
+ $X2=12.57 $Y2=0.38
r48 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.405 $Y=0.8
+ $X2=12.57 $Y2=0.715
r49 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=12.405 $Y=0.8
+ $X2=11.85 $Y2=0.8
r50 17 19 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=11.697 $Y=0.715
+ $X2=11.85 $Y2=0.8
r51 16 25 2.71076 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=11.697 $Y=0.425
+ $X2=11.697 $Y2=0.34
r52 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=11.697 $Y=0.425
+ $X2=11.697 $Y2=0.715
r53 14 25 4.84748 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=11.545 $Y=0.34
+ $X2=11.697 $Y2=0.34
r54 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.545 $Y=0.34
+ $X2=10.875 $Y2=0.34
r55 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.79 $Y=0.425
+ $X2=10.875 $Y2=0.34
r56 10 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=10.79 $Y=0.425
+ $X2=10.79 $Y2=0.605
r57 3 22 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=12.435
+ $Y=0.235 $X2=12.57 $Y2=0.38
r58 2 25 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=11.495
+ $Y=0.345 $X2=11.705 $Y2=0.42
r59 1 12 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=10.665
+ $Y=0.345 $X2=10.79 $Y2=0.605
.ends

