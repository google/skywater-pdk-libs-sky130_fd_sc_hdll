* File: sky130_fd_sc_hdll__a31oi_1.pex.spice
* Created: Thu Aug 27 18:55:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A31OI_1%A3 1 3 4 6 7 11
r20 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.35
+ $Y=1.16 $X2=0.35 $Y2=1.16
r21 7 11 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.23 $Y=1.16 $X2=0.35
+ $Y2=1.16
r22 4 10 38.7084 $w=3.43e-07 $l=2.14942e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.405 $Y2=1.16
r23 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r24 1 10 45.964 $w=3.43e-07 $l=2.91548e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.405 $Y2=1.16
r25 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_1%A2 1 3 4 6 7 8 9
r32 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.16
+ $X2=1 $Y2=1.16
r33 9 15 0.640756 $w=5.58e-07 $l=3e-08 $layer=LI1_cond $X=0.885 $Y=1.19
+ $X2=0.885 $Y2=1.16
r34 8 15 6.62115 $w=5.58e-07 $l=3.1e-07 $layer=LI1_cond $X=0.885 $Y=0.85
+ $X2=0.885 $Y2=1.16
r35 7 8 7.2619 $w=5.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.885 $Y=0.51 $X2=0.885
+ $Y2=0.85
r36 4 14 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=1 $Y2=1.16
r37 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r38 1 14 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=1 $Y2=1.16
r39 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995 $X2=0.94
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_1%A1 1 3 4 6 9 12 13 19
r38 13 19 7.33373 $w=2.18e-07 $l=1.4e-07 $layer=LI1_cond $X=1.15 $Y=1.555
+ $X2=1.29 $Y2=1.555
r39 12 19 4.1907 $w=2.18e-07 $l=8e-08 $layer=LI1_cond $X=1.37 $Y=1.555 $X2=1.29
+ $Y2=1.555
r40 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.505
+ $Y=1.16 $X2=1.505 $Y2=1.16
r41 7 12 7.15082 $w=2.2e-07 $l=2.09914e-07 $layer=LI1_cond $X=1.532 $Y=1.445
+ $X2=1.37 $Y2=1.555
r42 7 9 10.106 $w=3.23e-07 $l=2.85e-07 $layer=LI1_cond $X=1.532 $Y=1.445
+ $X2=1.532 $Y2=1.16
r43 4 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.47 $Y=1.41
+ $X2=1.505 $Y2=1.16
r44 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.47 $Y=1.41 $X2=1.47
+ $Y2=1.985
r45 1 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.445 $Y=0.995
+ $X2=1.505 $Y2=1.16
r46 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.445 $Y=0.995
+ $X2=1.445 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_1%B1 1 3 4 6 8 9 12 18
r34 13 18 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.41 $Y=1.16
+ $X2=2.505 $Y2=1.16
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.41
+ $Y=1.16 $X2=2.41 $Y2=1.16
r36 9 18 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=2.55 $Y=1.16
+ $X2=2.505 $Y2=1.16
r37 7 12 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=2.095 $Y=1.16
+ $X2=2.41 $Y2=1.16
r38 7 8 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=2.095 $Y=1.16
+ $X2=1.995 $Y2=1.202
r39 4 8 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=1.995 $Y=1.41
+ $X2=1.995 $Y2=1.202
r40 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.995 $Y=1.41
+ $X2=1.995 $Y2=1.985
r41 1 8 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=1.97 $Y=0.995
+ $X2=1.995 $Y2=1.202
r42 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.97 $Y=0.995 $X2=1.97
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_1%VPWR 1 2 7 9 15 17 19 29 30 36
r38 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r39 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r40 27 30 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r41 27 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r42 26 29 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r43 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r44 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.2 $Y2=2.72
r45 24 26 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.61 $Y2=2.72
r46 23 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r47 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 20 33 4.79676 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=0.42 $Y=2.72 $X2=0.21
+ $Y2=2.72
r49 20 22 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.42 $Y=2.72 $X2=0.69
+ $Y2=2.72
r50 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=1.2 $Y2=2.72
r51 19 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 17 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r53 17 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r54 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.72
r55 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.34
r56 9 12 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.255 $Y=1.66
+ $X2=0.255 $Y2=2.34
r57 7 33 2.96942 $w=3.3e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.255 $Y=2.635
+ $X2=0.21 $Y2=2.72
r58 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.255 $Y=2.635
+ $X2=0.255 $Y2=2.34
r59 2 15 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.34
r60 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r61 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_1%A_117_297# 1 2 9 11 12 15
r24 13 15 13.9347 $w=1.93e-07 $l=2.45e-07 $layer=LI1_cond $X=1.717 $Y=2.005
+ $X2=1.717 $Y2=2.25
r25 11 13 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=1.62 $Y=1.92
+ $X2=1.717 $Y2=2.005
r26 11 12 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.62 $Y=1.92
+ $X2=0.815 $Y2=1.92
r27 7 12 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.727 $Y=2.005
+ $X2=0.815 $Y2=1.92
r28 7 9 15.5273 $w=1.73e-07 $l=2.45e-07 $layer=LI1_cond $X=0.727 $Y=2.005
+ $X2=0.727 $Y2=2.25
r29 2 15 600 $w=1.7e-07 $l=8.34356e-07 $layer=licon1_PDIFF $count=1 $X=1.56
+ $Y=1.485 $X2=1.705 $Y2=2.25
r30 1 9 600 $w=1.7e-07 $l=8.34356e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.25
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_1%Y 1 2 12 16 17 18 19
r37 19 27 3.52512 $w=4.23e-07 $l=1.3e-07 $layer=LI1_cond $X=2.197 $Y=2.21
+ $X2=2.197 $Y2=2.34
r38 18 19 9.21954 $w=4.23e-07 $l=3.4e-07 $layer=LI1_cond $X=2.197 $Y=1.87
+ $X2=2.197 $Y2=2.21
r39 16 17 8.76046 $w=4.23e-07 $l=1.65e-07 $layer=LI1_cond $X=2.197 $Y=1.66
+ $X2=2.197 $Y2=1.495
r40 14 18 4.41996 $w=4.23e-07 $l=1.63e-07 $layer=LI1_cond $X=2.197 $Y=1.707
+ $X2=2.197 $Y2=1.87
r41 14 16 1.27447 $w=4.23e-07 $l=4.7e-08 $layer=LI1_cond $X=2.197 $Y=1.707
+ $X2=2.197 $Y2=1.66
r42 10 12 8.23714 $w=5.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=0.56
+ $X2=2.07 $Y2=0.56
r43 7 12 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=2.07 $Y=0.825
+ $X2=2.07 $Y2=0.56
r44 7 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.07 $Y=0.825
+ $X2=2.07 $Y2=1.495
r45 2 27 400 $w=1.7e-07 $l=9.29274e-07 $layer=licon1_PDIFF $count=1 $X=2.085
+ $Y=1.485 $X2=2.24 $Y2=2.34
r46 2 16 400 $w=1.7e-07 $l=2.40312e-07 $layer=licon1_PDIFF $count=1 $X=2.085
+ $Y=1.485 $X2=2.24 $Y2=1.66
r47 1 10 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=1.52
+ $Y=0.235 $X2=1.705 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_1%VGND 1 2 7 9 11 13 15 17 30
r30 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r31 24 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r32 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r33 21 24 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r34 20 23 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r35 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r36 18 26 4.89275 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.215
+ $Y2=0
r37 18 20 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.69
+ $Y2=0
r38 17 29 4.02327 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=2.542
+ $Y2=0
r39 17 23 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=2.07
+ $Y2=0
r40 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r41 15 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r42 11 29 3.18895 $w=2.6e-07 $l=1.22327e-07 $layer=LI1_cond $X=2.455 $Y=0.085
+ $X2=2.542 $Y2=0
r43 11 13 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=2.455 $Y=0.085
+ $X2=2.455 $Y2=0.4
r44 7 26 2.95841 $w=3.4e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.215 $Y2=0
r45 7 9 10.3381 $w=3.38e-07 $l=3.05e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.39
r46 2 13 182 $w=1.7e-07 $l=4.39829e-07 $layer=licon1_NDIFF $count=1 $X=2.045
+ $Y=0.235 $X2=2.41 $Y2=0.4
r47 1 9 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

