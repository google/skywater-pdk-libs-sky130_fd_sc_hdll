* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nor3_2 A B C VGND VNB VPB VPWR Y
X0 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 Y C a_309_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 a_309_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 a_309_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_297# B a_309_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
