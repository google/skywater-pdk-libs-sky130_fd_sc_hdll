* File: sky130_fd_sc_hdll__decap_6.pxi.spice
* Created: Wed Sep  2 08:27:46 2020
* 
x_PM_SKY130_FD_SC_HDLL__DECAP_6%VGND N_VGND_M1001_s N_VGND_c_16_n VGND
+ N_VGND_c_17_n N_VGND_M1000_g N_VGND_c_18_n N_VGND_c_19_n N_VGND_c_20_n
+ PM_SKY130_FD_SC_HDLL__DECAP_6%VGND
x_PM_SKY130_FD_SC_HDLL__DECAP_6%VPWR N_VPWR_M1000_s N_VPWR_M1001_g N_VPWR_c_42_n
+ N_VPWR_c_43_n VPWR N_VPWR_c_38_n N_VPWR_c_39_n N_VPWR_c_40_n N_VPWR_c_41_n
+ PM_SKY130_FD_SC_HDLL__DECAP_6%VPWR
cc_1 VNB N_VGND_c_16_n 0.0120582f $X=-0.19 $Y=-0.24 $X2=2.205 $Y2=0.385
cc_2 VNB N_VGND_c_17_n 0.0332598f $X=-0.19 $Y=-0.24 $X2=1.11 $Y2=1.29
cc_3 VNB N_VGND_c_18_n 0.0745114f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=0.475
cc_4 VNB N_VGND_c_19_n 0.0439751f $X=-0.19 $Y=-0.24 $X2=2.5 $Y2=0.475
cc_5 VNB N_VGND_c_20_n 0.159975f $X=-0.19 $Y=-0.24 $X2=2.53 $Y2=0
cc_6 VNB N_VPWR_c_38_n 0.121206f $X=-0.19 $Y=-0.24 $X2=1.38 $Y2=2.05
cc_7 VNB N_VPWR_c_39_n 0.0831799f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=0
cc_8 VNB N_VPWR_c_40_n 0.0178259f $X=-0.19 $Y=-0.24 $X2=2.5 $Y2=0.475
cc_9 VNB N_VPWR_c_41_n 0.117919f $X=-0.19 $Y=-0.24 $X2=2.53 $Y2=0
cc_10 VPB N_VGND_c_17_n 0.17121f $X=-0.19 $Y=1.305 $X2=1.11 $Y2=1.29
cc_11 VPB N_VGND_c_18_n 0.0068688f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=0.475
cc_12 VPB N_VPWR_c_42_n 0.00993338f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_13 VPB N_VPWR_c_43_n 0.0597303f $X=-0.19 $Y=1.305 $X2=1.11 $Y2=1.29
cc_14 VPB N_VPWR_c_40_n 0.0771788f $X=-0.19 $Y=1.305 $X2=2.5 $Y2=0.475
cc_15 VPB N_VPWR_c_41_n 0.0420516f $X=-0.19 $Y=1.305 $X2=2.53 $Y2=0
cc_16 N_VGND_c_17_n N_VPWR_c_42_n 0.100391f $X=1.11 $Y=1.29 $X2=0 $Y2=0
cc_17 N_VGND_c_18_n N_VPWR_c_42_n 0.0489119f $X=0.26 $Y=0.475 $X2=0 $Y2=0
cc_18 N_VGND_c_17_n N_VPWR_c_43_n 0.0493583f $X=1.11 $Y=1.29 $X2=0 $Y2=0
cc_19 N_VGND_c_18_n N_VPWR_c_43_n 0.0561345f $X=0.26 $Y=0.475 $X2=0 $Y2=0
cc_20 N_VGND_c_16_n N_VPWR_c_38_n 0.0738934f $X=2.205 $Y=0.385 $X2=0 $Y2=0
cc_21 N_VGND_c_17_n N_VPWR_c_38_n 0.0673714f $X=1.11 $Y=1.29 $X2=0 $Y2=0
cc_22 N_VGND_c_18_n N_VPWR_c_38_n 0.00648593f $X=0.26 $Y=0.475 $X2=0 $Y2=0
cc_23 N_VGND_c_19_n N_VPWR_c_38_n 0.0237188f $X=2.5 $Y=0.475 $X2=0 $Y2=0
cc_24 N_VGND_c_16_n N_VPWR_c_39_n 0.0203068f $X=2.205 $Y=0.385 $X2=0 $Y2=0
cc_25 N_VGND_c_17_n N_VPWR_c_39_n 0.0617788f $X=1.11 $Y=1.29 $X2=0 $Y2=0
cc_26 N_VGND_c_18_n N_VPWR_c_39_n 0.105038f $X=0.26 $Y=0.475 $X2=0 $Y2=0
cc_27 N_VGND_c_16_n N_VPWR_c_40_n 0.0623495f $X=2.205 $Y=0.385 $X2=0 $Y2=0
cc_28 N_VGND_c_17_n N_VPWR_c_40_n 0.138185f $X=1.11 $Y=1.29 $X2=0 $Y2=0
cc_29 N_VGND_c_18_n N_VPWR_c_40_n 0.0327855f $X=0.26 $Y=0.475 $X2=0 $Y2=0
cc_30 N_VGND_c_19_n N_VPWR_c_40_n 0.0425904f $X=2.5 $Y=0.475 $X2=0 $Y2=0
