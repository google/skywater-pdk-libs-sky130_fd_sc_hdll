* NGSPICE file created from sky130_fd_sc_hdll__o211a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=1.12e+12p pd=8.24e+06u as=3e+11p ps=2.6e+06u
M1001 a_120_47# C1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=2.0475e+11p ps=1.93e+06u
M1002 VPWR C1 a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.055e+12p ps=6.11e+06u
M1003 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_206_47# B1 a_120_47# VNB nshort w=650000u l=150000u
+  ad=3.7375e+11p pd=3.75e+06u as=0p ps=0u
M1005 a_206_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.4425e+11p ps=6.19e+06u
M1006 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=2.34e+11p pd=2.02e+06u as=0p ps=0u
M1007 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_47# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A1 a_206_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_406_297# A2 a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=2.3e+11p pd=2.46e+06u as=0p ps=0u
M1011 VPWR A1 a_406_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

