* File: sky130_fd_sc_hdll__sdfxbp_2.pxi.spice
* Created: Wed Sep  2 08:52:13 2020
* 
x_PM_SKY130_FD_SC_HDLL__SDFXBP_2%CLK N_CLK_c_241_n N_CLK_c_245_n N_CLK_c_246_n
+ N_CLK_M1010_g N_CLK_c_242_n N_CLK_M1029_g CLK
+ PM_SKY130_FD_SC_HDLL__SDFXBP_2%CLK
x_PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_27_47# N_A_27_47#_M1029_s N_A_27_47#_M1010_s
+ N_A_27_47#_c_294_n N_A_27_47#_c_295_n N_A_27_47#_M1033_g N_A_27_47#_M1001_g
+ N_A_27_47#_M1009_g N_A_27_47#_c_283_n N_A_27_47#_c_284_n N_A_27_47#_c_298_n
+ N_A_27_47#_c_299_n N_A_27_47#_M1023_g N_A_27_47#_c_300_n N_A_27_47#_c_301_n
+ N_A_27_47#_M1008_g N_A_27_47#_c_285_n N_A_27_47#_M1038_g N_A_27_47#_c_511_p
+ N_A_27_47#_c_287_n N_A_27_47#_c_288_n N_A_27_47#_c_303_n N_A_27_47#_c_289_n
+ N_A_27_47#_c_400_p N_A_27_47#_c_304_n N_A_27_47#_c_305_n N_A_27_47#_c_290_n
+ N_A_27_47#_c_306_n N_A_27_47#_c_307_n N_A_27_47#_c_308_n N_A_27_47#_c_309_n
+ N_A_27_47#_c_310_n N_A_27_47#_c_311_n N_A_27_47#_c_291_n N_A_27_47#_c_292_n
+ N_A_27_47#_c_293_n PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_319_47# N_A_319_47#_M1021_s
+ N_A_319_47#_M1022_s N_A_319_47#_M1031_g N_A_319_47#_c_532_n
+ N_A_319_47#_M1011_g N_A_319_47#_c_526_n N_A_319_47#_c_534_n
+ N_A_319_47#_c_541_n N_A_319_47#_c_527_n N_A_319_47#_c_528_n
+ N_A_319_47#_c_529_n N_A_319_47#_c_543_n N_A_319_47#_c_536_n
+ N_A_319_47#_c_530_n N_A_319_47#_c_537_n N_A_319_47#_c_547_n
+ N_A_319_47#_c_538_n N_A_319_47#_c_531_n
+ PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_319_47#
x_PM_SKY130_FD_SC_HDLL__SDFXBP_2%SCE N_SCE_c_652_n N_SCE_M1022_g N_SCE_M1021_g
+ N_SCE_c_654_n N_SCE_c_655_n N_SCE_M1016_g N_SCE_M1019_g N_SCE_c_656_n
+ N_SCE_c_647_n N_SCE_c_648_n N_SCE_c_649_n SCE N_SCE_c_650_n N_SCE_c_716_p SCE
+ PM_SKY130_FD_SC_HDLL__SDFXBP_2%SCE
x_PM_SKY130_FD_SC_HDLL__SDFXBP_2%D N_D_c_749_n N_D_M1020_g N_D_M1014_g D
+ PM_SKY130_FD_SC_HDLL__SDFXBP_2%D
x_PM_SKY130_FD_SC_HDLL__SDFXBP_2%SCD N_SCD_M1037_g N_SCD_c_788_n N_SCD_c_789_n
+ N_SCD_M1007_g SCD N_SCD_c_787_n PM_SKY130_FD_SC_HDLL__SDFXBP_2%SCD
x_PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_211_363# N_A_211_363#_M1001_d
+ N_A_211_363#_M1033_d N_A_211_363#_c_848_n N_A_211_363#_M1028_g
+ N_A_211_363#_c_835_n N_A_211_363#_M1034_g N_A_211_363#_c_836_n
+ N_A_211_363#_M1030_g N_A_211_363#_c_849_n N_A_211_363#_M1036_g
+ N_A_211_363#_c_837_n N_A_211_363#_c_838_n N_A_211_363#_c_839_n
+ N_A_211_363#_c_852_n N_A_211_363#_c_840_n N_A_211_363#_c_841_n
+ N_A_211_363#_c_842_n N_A_211_363#_c_843_n N_A_211_363#_c_957_p
+ N_A_211_363#_c_844_n N_A_211_363#_c_845_n N_A_211_363#_c_901_n
+ N_A_211_363#_c_846_n N_A_211_363#_c_847_n
+ PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_211_363#
x_PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_1179_183# N_A_1179_183#_M1002_d
+ N_A_1179_183#_M1025_d N_A_1179_183#_c_1040_n N_A_1179_183#_c_1048_n
+ N_A_1179_183#_M1000_g N_A_1179_183#_M1017_g N_A_1179_183#_c_1042_n
+ N_A_1179_183#_c_1072_n N_A_1179_183#_c_1092_p N_A_1179_183#_c_1073_n
+ N_A_1179_183#_c_1043_n N_A_1179_183#_c_1044_n N_A_1179_183#_c_1059_n
+ N_A_1179_183#_c_1045_n N_A_1179_183#_c_1046_n
+ PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_1179_183#
x_PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_1001_47# N_A_1001_47#_M1009_d
+ N_A_1001_47#_M1028_d N_A_1001_47#_c_1140_n N_A_1001_47#_c_1147_n
+ N_A_1001_47#_M1025_g N_A_1001_47#_M1002_g N_A_1001_47#_c_1141_n
+ N_A_1001_47#_c_1142_n N_A_1001_47#_c_1143_n N_A_1001_47#_c_1144_n
+ N_A_1001_47#_c_1162_n N_A_1001_47#_c_1167_n N_A_1001_47#_c_1145_n
+ N_A_1001_47#_c_1150_n N_A_1001_47#_c_1146_n
+ PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_1001_47#
x_PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_1653_315# N_A_1653_315#_M1039_s
+ N_A_1653_315#_M1015_s N_A_1653_315#_c_1266_n N_A_1653_315#_M1032_g
+ N_A_1653_315#_M1024_g N_A_1653_315#_c_1268_n N_A_1653_315#_M1003_g
+ N_A_1653_315#_c_1257_n N_A_1653_315#_M1013_g N_A_1653_315#_c_1269_n
+ N_A_1653_315#_M1026_g N_A_1653_315#_c_1258_n N_A_1653_315#_M1035_g
+ N_A_1653_315#_c_1259_n N_A_1653_315#_c_1260_n N_A_1653_315#_c_1272_n
+ N_A_1653_315#_c_1273_n N_A_1653_315#_M1018_g N_A_1653_315#_M1027_g
+ N_A_1653_315#_c_1262_n N_A_1653_315#_c_1275_n N_A_1653_315#_c_1276_n
+ N_A_1653_315#_c_1263_n N_A_1653_315#_c_1277_n N_A_1653_315#_c_1264_n
+ N_A_1653_315#_c_1265_n N_A_1653_315#_c_1279_n N_A_1653_315#_c_1293_p
+ PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_1653_315#
x_PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_1464_413# N_A_1464_413#_M1030_d
+ N_A_1464_413#_M1008_d N_A_1464_413#_c_1378_n N_A_1464_413#_M1015_g
+ N_A_1464_413#_c_1372_n N_A_1464_413#_M1039_g N_A_1464_413#_c_1373_n
+ N_A_1464_413#_c_1374_n N_A_1464_413#_c_1384_n N_A_1464_413#_c_1388_n
+ N_A_1464_413#_c_1381_n N_A_1464_413#_c_1375_n N_A_1464_413#_c_1376_n
+ N_A_1464_413#_c_1377_n PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_1464_413#
x_PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_2234_47# N_A_2234_47#_M1027_s
+ N_A_2234_47#_M1018_s N_A_2234_47#_c_1461_n N_A_2234_47#_M1005_g
+ N_A_2234_47#_c_1455_n N_A_2234_47#_M1004_g N_A_2234_47#_c_1462_n
+ N_A_2234_47#_M1012_g N_A_2234_47#_c_1456_n N_A_2234_47#_M1006_g
+ N_A_2234_47#_c_1457_n N_A_2234_47#_c_1463_n N_A_2234_47#_c_1458_n
+ N_A_2234_47#_c_1459_n N_A_2234_47#_c_1460_n
+ PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_2234_47#
x_PM_SKY130_FD_SC_HDLL__SDFXBP_2%VPWR N_VPWR_M1010_d N_VPWR_M1022_d
+ N_VPWR_M1007_d N_VPWR_M1000_d N_VPWR_M1032_d N_VPWR_M1015_d N_VPWR_M1026_d
+ N_VPWR_M1018_d N_VPWR_M1012_d N_VPWR_c_1518_n N_VPWR_c_1519_n N_VPWR_c_1520_n
+ N_VPWR_c_1521_n N_VPWR_c_1522_n N_VPWR_c_1523_n N_VPWR_c_1524_n
+ N_VPWR_c_1525_n N_VPWR_c_1526_n N_VPWR_c_1527_n N_VPWR_c_1528_n
+ N_VPWR_c_1529_n N_VPWR_c_1530_n N_VPWR_c_1531_n N_VPWR_c_1532_n
+ N_VPWR_c_1533_n N_VPWR_c_1534_n VPWR N_VPWR_c_1535_n N_VPWR_c_1536_n
+ N_VPWR_c_1537_n N_VPWR_c_1538_n N_VPWR_c_1539_n N_VPWR_c_1540_n
+ N_VPWR_c_1541_n N_VPWR_c_1542_n N_VPWR_c_1543_n N_VPWR_c_1544_n
+ N_VPWR_c_1517_n PM_SKY130_FD_SC_HDLL__SDFXBP_2%VPWR
x_PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_604_369# N_A_604_369#_M1014_d
+ N_A_604_369#_M1009_s N_A_604_369#_M1020_d N_A_604_369#_M1028_s
+ N_A_604_369#_c_1727_n N_A_604_369#_c_1740_n N_A_604_369#_c_1741_n
+ N_A_604_369#_c_1716_n N_A_604_369#_c_1723_n N_A_604_369#_c_1724_n
+ N_A_604_369#_c_1717_n N_A_604_369#_c_1718_n N_A_604_369#_c_1719_n
+ N_A_604_369#_c_1720_n N_A_604_369#_c_1721_n N_A_604_369#_c_1722_n
+ N_A_604_369#_c_1726_n PM_SKY130_FD_SC_HDLL__SDFXBP_2%A_604_369#
x_PM_SKY130_FD_SC_HDLL__SDFXBP_2%Q N_Q_M1013_d N_Q_M1003_s Q N_Q_c_1844_n
+ PM_SKY130_FD_SC_HDLL__SDFXBP_2%Q
x_PM_SKY130_FD_SC_HDLL__SDFXBP_2%Q_N N_Q_N_M1004_s N_Q_N_M1005_s Q_N
+ N_Q_N_c_1863_n PM_SKY130_FD_SC_HDLL__SDFXBP_2%Q_N
x_PM_SKY130_FD_SC_HDLL__SDFXBP_2%VGND N_VGND_M1029_d N_VGND_M1021_d
+ N_VGND_M1037_d N_VGND_M1017_d N_VGND_M1024_d N_VGND_M1039_d N_VGND_M1035_s
+ N_VGND_M1027_d N_VGND_M1006_d N_VGND_c_1880_n N_VGND_c_1881_n N_VGND_c_1882_n
+ N_VGND_c_1883_n N_VGND_c_1884_n N_VGND_c_1885_n N_VGND_c_1886_n
+ N_VGND_c_1887_n N_VGND_c_1888_n N_VGND_c_1889_n N_VGND_c_1890_n
+ N_VGND_c_1891_n N_VGND_c_1892_n N_VGND_c_1893_n VGND N_VGND_c_1894_n
+ N_VGND_c_1895_n N_VGND_c_1896_n N_VGND_c_1897_n N_VGND_c_1898_n
+ N_VGND_c_1899_n N_VGND_c_1900_n N_VGND_c_1901_n N_VGND_c_1902_n
+ N_VGND_c_1903_n N_VGND_c_1904_n N_VGND_c_1905_n N_VGND_c_1906_n
+ PM_SKY130_FD_SC_HDLL__SDFXBP_2%VGND
cc_1 VNB N_CLK_c_241_n 0.0607903f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.325
cc_2 VNB N_CLK_c_242_n 0.0173562f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_3 VNB CLK 0.0188452f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_27_47#_M1001_g 0.0398894f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_27_47#_M1009_g 0.0541072f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_c_283_n 0.0165761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_284_n 0.00284949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_285_n 0.0212345f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1038_g 0.0472025f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_287_n 0.00339765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_288_n 0.00647711f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_289_n 0.00204906f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_290_n 0.00522807f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_291_n 0.0260131f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_292_n 0.0106395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_293_n 0.00177482f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_319_47#_M1031_g 0.0244273f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_18 VNB N_A_319_47#_c_526_n 0.0147622f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_19 VNB N_A_319_47#_c_527_n 0.00282526f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_319_47#_c_528_n 0.00166871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_319_47#_c_529_n 0.00382184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_319_47#_c_530_n 0.00277255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_319_47#_c_531_n 0.0296191f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_SCE_M1021_g 0.0562132f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_25 VNB N_SCE_M1019_g 0.0173732f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_26 VNB N_SCE_c_647_n 0.00476782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_SCE_c_648_n 0.0171124f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_SCE_c_649_n 0.00121137f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_SCE_c_650_n 0.0320765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB SCE 0.00162963f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_D_M1014_g 0.0503241f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_32 VNB N_SCD_M1037_g 0.046913f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.74
cc_33 VNB SCD 0.00538176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_SCD_c_787_n 0.0173777f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_35 VNB N_A_211_363#_c_835_n 0.0184077f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_211_363#_c_836_n 0.0191164f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_37 VNB N_A_211_363#_c_837_n 0.00361085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_211_363#_c_838_n 0.00443734f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_211_363#_c_839_n 0.00672004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_211_363#_c_840_n 0.00954394f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_211_363#_c_841_n 0.0015014f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_211_363#_c_842_n 0.00211521f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_211_363#_c_843_n 0.0110991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_211_363#_c_844_n 0.0136749f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_211_363#_c_845_n 0.00640764f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_211_363#_c_846_n 0.0312456f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_211_363#_c_847_n 0.0341862f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_1179_183#_c_1040_n 0.0161342f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_49 VNB N_A_1179_183#_M1017_g 0.0216963f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_1179_183#_c_1042_n 0.00354578f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_51 VNB N_A_1179_183#_c_1043_n 0.0043246f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_1179_183#_c_1044_n 0.00133147f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_1179_183#_c_1045_n 0.00316561f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1179_183#_c_1046_n 0.0370936f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_1001_47#_c_1140_n 0.0127944f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_56 VNB N_A_1001_47#_c_1141_n 0.0162173f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_57 VNB N_A_1001_47#_c_1142_n 0.017433f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_58 VNB N_A_1001_47#_c_1143_n 0.00914068f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_59 VNB N_A_1001_47#_c_1144_n 0.00101096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_1001_47#_c_1145_n 0.0131749f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_1001_47#_c_1146_n 0.00182328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_1653_315#_M1024_g 0.0483572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1653_315#_c_1257_n 0.018089f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_64 VNB N_A_1653_315#_c_1258_n 0.0199361f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_1653_315#_c_1259_n 0.0499109f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1653_315#_c_1260_n 0.0418231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1653_315#_M1027_g 0.0377787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1653_315#_c_1262_n 0.0127355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_1653_315#_c_1263_n 0.00257179f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_1653_315#_c_1264_n 0.00241353f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_1653_315#_c_1265_n 0.00808857f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_1464_413#_c_1372_n 0.0207831f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1464_413#_c_1373_n 0.0410096f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.105
cc_74 VNB N_A_1464_413#_c_1374_n 0.0116501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1464_413#_c_1375_n 0.00860132f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_1464_413#_c_1376_n 0.00584669f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1464_413#_c_1377_n 0.00364926f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_2234_47#_c_1455_n 0.0195452f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_2234_47#_c_1456_n 0.0205912f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_80 VNB N_A_2234_47#_c_1457_n 0.0114678f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_2234_47#_c_1458_n 0.00720247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_2234_47#_c_1459_n 4.07275e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_2234_47#_c_1460_n 0.0595632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VPWR_c_1517_n 0.554392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_604_369#_c_1716_n 3.46824e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_604_369#_c_1717_n 0.0166845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_604_369#_c_1718_n 0.00543757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_604_369#_c_1719_n 0.00314477f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_604_369#_c_1720_n 0.00896062f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_604_369#_c_1721_n 0.00188916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_604_369#_c_1722_n 0.00194402f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_Q_c_1844_n 0.00105123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_Q_N_c_1863_n 0.0018494f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1880_n 0.00562936f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1881_n 0.00491179f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1882_n 0.00586751f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1883_n 0.00404537f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1884_n 0.00611774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1885_n 0.00967872f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1886_n 0.0220055f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1887_n 0.00892965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1888_n 0.0113721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1889_n 0.0103365f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1890_n 0.033696f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1891_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1892_n 0.0405525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1893_n 0.0038195f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1894_n 0.0154125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1895_n 0.0494436f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1896_n 0.0477763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1897_n 0.0213119f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1898_n 0.0191557f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1899_n 0.0194083f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1900_n 0.0085923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1901_n 0.00709041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1902_n 0.00580517f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1903_n 0.0080786f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1904_n 0.00442399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1905_n 0.0121179f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1906_n 0.626053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VPB N_CLK_c_241_n 0.00482568f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_122 VPB N_CLK_c_245_n 0.0148284f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.59
cc_123 VPB N_CLK_c_246_n 0.0462588f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.74
cc_124 VPB CLK 0.0178738f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_125 VPB N_A_27_47#_c_294_n 0.0193314f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_126 VPB N_A_27_47#_c_295_n 0.0253151f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_127 VPB N_A_27_47#_c_283_n 0.0157793f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_27_47#_c_284_n 0.00578676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_27_47#_c_298_n 0.0117214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_27_47#_c_299_n 0.0505757f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_27_47#_c_300_n 0.015896f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_27_47#_c_301_n 0.022678f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_27_47#_c_285_n 0.0244074f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_27_47#_c_303_n 0.00217719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_27_47#_c_304_n 0.00381244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_27_47#_c_305_n 0.0035907f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_27_47#_c_306_n 0.0588483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_27_47#_c_307_n 0.0013034f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_27_47#_c_308_n 0.00246423f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_27_47#_c_309_n 9.17012e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_27_47#_c_310_n 0.0087556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_27_47#_c_311_n 0.00434106f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_27_47#_c_291_n 0.0119092f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_27_47#_c_292_n 0.0223895f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_27_47#_c_293_n 0.00461343f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_319_47#_c_532_n 0.0520644f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.665
cc_147 VPB N_A_319_47#_c_526_n 0.0109024f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.16
cc_148 VPB N_A_319_47#_c_534_n 0.00448421f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_319_47#_c_527_n 0.00468231f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_319_47#_c_536_n 0.00160776f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_319_47#_c_537_n 0.00202192f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_319_47#_c_538_n 0.00186942f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_SCE_c_652_n 0.0621217f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_154 VPB N_SCE_M1021_g 0.0054864f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_155 VPB N_SCE_c_654_n 0.0129207f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_156 VPB N_SCE_c_655_n 0.0159667f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_SCE_c_656_n 0.0162338f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_158 VPB N_SCE_c_647_n 7.34924e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_D_c_749_n 0.0504862f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_160 VPB N_D_M1014_g 0.0044562f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_161 VPB D 0.00614535f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_162 VPB N_SCD_c_788_n 0.00981036f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_163 VPB N_SCD_c_789_n 0.02746f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_164 VPB SCD 0.00583016f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_SCD_c_787_n 0.0217377f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_166 VPB N_A_211_363#_c_848_n 0.0628983f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_167 VPB N_A_211_363#_c_849_n 0.0544959f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_168 VPB N_A_211_363#_c_837_n 0.00470057f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_211_363#_c_838_n 0.00380616f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_211_363#_c_852_n 0.00625509f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_211_363#_c_844_n 0.0118281f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_1179_183#_c_1040_n 0.0313232f $X=-0.19 $Y=1.305 $X2=0.52
+ $Y2=0.445
cc_173 VPB N_A_1179_183#_c_1048_n 0.0245924f $X=-0.19 $Y=1.305 $X2=0.31
+ $Y2=1.665
cc_174 VPB N_A_1179_183#_c_1045_n 0.00256319f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_1001_47#_c_1147_n 0.018063f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_176 VPB N_A_1001_47#_c_1143_n 0.0189969f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_177 VPB N_A_1001_47#_c_1144_n 0.0158981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_1001_47#_c_1150_n 0.00162511f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_1001_47#_c_1146_n 0.00893798f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_1653_315#_c_1266_n 0.0705156f $X=-0.19 $Y=1.305 $X2=0.52
+ $Y2=0.445
cc_181 VPB N_A_1653_315#_M1024_g 0.0179547f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_1653_315#_c_1268_n 0.0170437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_1653_315#_c_1269_n 0.0193533f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_A_1653_315#_c_1259_n 0.0318469f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_1653_315#_c_1260_n 0.0280345f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_1653_315#_c_1272_n 0.0272315f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_1653_315#_c_1273_n 0.0305021f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_1653_315#_c_1262_n 8.03011e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_1653_315#_c_1275_n 0.0110649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_A_1653_315#_c_1276_n 0.00737531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_A_1653_315#_c_1277_n 0.00231467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_A_1653_315#_c_1264_n 0.00241353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_A_1653_315#_c_1279_n 9.71818e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_A_1464_413#_c_1378_n 0.0206604f $X=-0.19 $Y=1.305 $X2=0.52
+ $Y2=0.445
cc_195 VPB N_A_1464_413#_c_1373_n 0.0157025f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_196 VPB N_A_1464_413#_c_1374_n 0.00763995f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_A_1464_413#_c_1381_n 0.00777195f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_A_1464_413#_c_1375_n 0.00382552f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_A_1464_413#_c_1376_n 0.0071082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_A_2234_47#_c_1461_n 0.0182155f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_201 VPB N_A_2234_47#_c_1462_n 0.0188164f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_202 VPB N_A_2234_47#_c_1463_n 0.0130405f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_A_2234_47#_c_1458_n 0.00634334f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_A_2234_47#_c_1460_n 0.0298458f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1518_n 0.00126291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1519_n 4.89699e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1520_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1521_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1522_n 0.00550337f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1523_n 0.00331524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1524_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1525_n 0.023495f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1526_n 0.00699073f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1527_n 0.0113462f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1528_n 0.0112895f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1529_n 0.0425429f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1530_n 0.00324297f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1531_n 0.0547273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1532_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1533_n 0.0513405f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1534_n 0.00584025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1535_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1536_n 0.0274845f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1537_n 0.0207768f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1538_n 0.0186002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1539_n 0.0189301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1540_n 0.0054556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1541_n 0.00502699f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1542_n 0.00686913f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1543_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1544_n 0.0104276f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1517_n 0.0736121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_A_604_369#_c_1723_n 0.00779562f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_A_604_369#_c_1724_n 0.00158613f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_A_604_369#_c_1720_n 0.0110413f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_A_604_369#_c_1726_n 0.00897532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_Q_c_1844_n 0.00154493f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_Q_N_c_1863_n 0.00153806f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 N_CLK_c_245_n N_A_27_47#_c_294_n 0.00267643f $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_240 N_CLK_c_246_n N_A_27_47#_c_294_n 0.0066814f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_241 CLK N_A_27_47#_c_294_n 8.10055e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_242 N_CLK_c_246_n N_A_27_47#_c_295_n 0.0193458f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_243 N_CLK_c_241_n N_A_27_47#_M1001_g 0.00195891f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_244 N_CLK_c_242_n N_A_27_47#_M1001_g 0.01543f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_245 N_CLK_c_241_n N_A_27_47#_c_287_n 0.0107312f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_246 N_CLK_c_242_n N_A_27_47#_c_287_n 0.00638787f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_247 CLK N_A_27_47#_c_287_n 0.00774265f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_248 N_CLK_c_241_n N_A_27_47#_c_288_n 0.00622672f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_249 CLK N_A_27_47#_c_288_n 0.0144574f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_250 N_CLK_c_246_n N_A_27_47#_c_303_n 0.0170291f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_251 CLK N_A_27_47#_c_303_n 0.00769886f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_252 N_CLK_c_241_n N_A_27_47#_c_289_n 5.45607e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_253 CLK N_A_27_47#_c_289_n 0.0429117f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_254 N_CLK_c_241_n N_A_27_47#_c_304_n 3.04005e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_255 N_CLK_c_245_n N_A_27_47#_c_304_n 4.49617e-19 $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_256 N_CLK_c_246_n N_A_27_47#_c_304_n 0.00442243f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_257 N_CLK_c_241_n N_A_27_47#_c_305_n 2.46885e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_258 N_CLK_c_246_n N_A_27_47#_c_305_n 0.00784199f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_259 CLK N_A_27_47#_c_305_n 0.0153591f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_260 N_CLK_c_241_n N_A_27_47#_c_290_n 0.00189681f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_261 N_CLK_c_246_n N_A_27_47#_c_307_n 0.00101717f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_262 N_CLK_c_241_n N_A_27_47#_c_291_n 0.0130772f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_263 CLK N_A_27_47#_c_291_n 0.00184152f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_264 N_CLK_c_242_n N_A_211_363#_c_841_n 5.8539e-19 $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_265 N_CLK_c_246_n N_VPWR_c_1518_n 0.0125197f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_266 N_CLK_c_246_n N_VPWR_c_1535_n 0.00304525f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_267 N_CLK_c_246_n N_VPWR_c_1517_n 0.00454898f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_268 N_CLK_c_241_n N_VGND_c_1894_n 6.28829e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_269 N_CLK_c_242_n N_VGND_c_1894_n 0.00198377f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_270 N_CLK_c_242_n N_VGND_c_1900_n 0.0142867f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_271 N_CLK_c_242_n N_VGND_c_1906_n 0.00367064f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_272 N_A_27_47#_c_306_n N_A_319_47#_c_532_n 0.00327847f $X=5.555 $Y=1.87 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_306_n N_A_319_47#_c_526_n 0.0122495f $X=5.555 $Y=1.87 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_306_n N_A_319_47#_c_541_n 0.0180318f $X=5.555 $Y=1.87 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_306_n N_A_319_47#_c_527_n 0.0087525f $X=5.555 $Y=1.87 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_306_n N_A_319_47#_c_543_n 0.0423833f $X=5.555 $Y=1.87 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_306_n N_A_319_47#_c_536_n 0.012446f $X=5.555 $Y=1.87 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_M1001_g N_A_319_47#_c_530_n 0.00138585f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_306_n N_A_319_47#_c_537_n 0.0137859f $X=5.555 $Y=1.87 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_306_n N_A_319_47#_c_547_n 0.0046091f $X=5.555 $Y=1.87 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_306_n N_A_319_47#_c_538_n 7.81108e-19 $X=5.555 $Y=1.87 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_306_n N_A_319_47#_c_531_n 0.00297526f $X=5.555 $Y=1.87 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_294_n N_SCE_c_652_n 0.00238227f $X=0.965 $Y=1.64 $X2=-0.19
+ $Y2=-0.24
cc_284 N_A_27_47#_c_306_n N_SCE_c_652_n 0.0101204f $X=5.555 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_285 N_A_27_47#_c_306_n N_SCE_c_655_n 0.0021692f $X=5.555 $Y=1.87 $X2=0 $Y2=0
cc_286 N_A_27_47#_c_306_n N_SCE_c_656_n 2.52518e-19 $X=5.555 $Y=1.87 $X2=0 $Y2=0
cc_287 N_A_27_47#_c_306_n N_SCE_c_647_n 0.00399737f $X=5.555 $Y=1.87 $X2=0 $Y2=0
cc_288 N_A_27_47#_c_306_n N_D_c_749_n 0.00594499f $X=5.555 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_289 N_A_27_47#_c_306_n D 0.00929306f $X=5.555 $Y=1.87 $X2=0 $Y2=0
cc_290 N_A_27_47#_c_306_n N_SCD_c_789_n 0.00274884f $X=5.555 $Y=1.87 $X2=0 $Y2=0
cc_291 N_A_27_47#_c_306_n SCD 0.0133868f $X=5.555 $Y=1.87 $X2=0 $Y2=0
cc_292 N_A_27_47#_M1009_g N_SCD_c_787_n 0.00191568f $X=4.93 $Y=0.415 $X2=0 $Y2=0
cc_293 N_A_27_47#_c_306_n N_A_211_363#_M1033_d 0.00143359f $X=5.555 $Y=1.87
+ $X2=0 $Y2=0
cc_294 N_A_27_47#_c_284_n N_A_211_363#_c_848_n 0.0194945f $X=5.005 $Y=1.32 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_299_n N_A_211_363#_c_848_n 0.0316622f $X=5.465 $Y=1.99 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_306_n N_A_211_363#_c_848_n 0.0095879f $X=5.555 $Y=1.87 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_310_n N_A_211_363#_c_848_n 0.00224123f $X=5.7 $Y=1.87 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_M1009_g N_A_211_363#_c_835_n 0.0125566f $X=4.93 $Y=0.415 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_M1038_g N_A_211_363#_c_836_n 0.0136788f $X=8 $Y=0.415 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_300_n N_A_211_363#_c_849_n 0.0184225f $X=7.23 $Y=1.89 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_301_n N_A_211_363#_c_849_n 0.0117705f $X=7.23 $Y=1.99 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_285_n N_A_211_363#_c_849_n 0.0237682f $X=7.925 $Y=1.32 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_311_n N_A_211_363#_c_849_n 0.00137325f $X=7.26 $Y=1.87 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_293_n N_A_211_363#_c_849_n 0.00168213f $X=7.2 $Y=1.41 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_M1009_g N_A_211_363#_c_837_n 0.00797646f $X=4.93 $Y=0.415
+ $X2=0 $Y2=0
cc_306 N_A_27_47#_c_283_n N_A_211_363#_c_837_n 0.00920069f $X=5.365 $Y=1.32
+ $X2=0 $Y2=0
cc_307 N_A_27_47#_c_284_n N_A_211_363#_c_837_n 0.00418731f $X=5.005 $Y=1.32
+ $X2=0 $Y2=0
cc_308 N_A_27_47#_c_298_n N_A_211_363#_c_837_n 0.00641846f $X=5.465 $Y=1.575
+ $X2=0 $Y2=0
cc_309 N_A_27_47#_c_299_n N_A_211_363#_c_837_n 7.35344e-19 $X=5.465 $Y=1.99
+ $X2=0 $Y2=0
cc_310 N_A_27_47#_c_306_n N_A_211_363#_c_837_n 0.0161657f $X=5.555 $Y=1.87 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_310_n N_A_211_363#_c_837_n 0.0171769f $X=5.7 $Y=1.87 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_285_n N_A_211_363#_c_838_n 0.0121391f $X=7.925 $Y=1.32 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_M1038_g N_A_211_363#_c_838_n 0.00393345f $X=8 $Y=0.415 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_292_n N_A_211_363#_c_838_n 0.00416507f $X=7.225 $Y=1.32
+ $X2=0 $Y2=0
cc_315 N_A_27_47#_c_293_n N_A_211_363#_c_838_n 0.023853f $X=7.2 $Y=1.41 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_M1038_g N_A_211_363#_c_839_n 0.0022503f $X=8 $Y=0.415 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_292_n N_A_211_363#_c_839_n 0.00228363f $X=7.225 $Y=1.32
+ $X2=0 $Y2=0
cc_318 N_A_27_47#_c_293_n N_A_211_363#_c_839_n 0.0149393f $X=7.2 $Y=1.41 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_300_n N_A_211_363#_c_852_n 0.0011999f $X=7.23 $Y=1.89 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_285_n N_A_211_363#_c_852_n 0.00449357f $X=7.925 $Y=1.32
+ $X2=0 $Y2=0
cc_321 N_A_27_47#_c_311_n N_A_211_363#_c_852_n 0.00509777f $X=7.26 $Y=1.87 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_293_n N_A_211_363#_c_852_n 0.0251353f $X=7.2 $Y=1.41 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_M1009_g N_A_211_363#_c_840_n 0.00298f $X=4.93 $Y=0.415 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_M1001_g N_A_211_363#_c_841_n 0.006485f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_M1009_g N_A_211_363#_c_842_n 0.00182155f $X=4.93 $Y=0.415
+ $X2=0 $Y2=0
cc_326 N_A_27_47#_c_283_n N_A_211_363#_c_843_n 4.20893e-19 $X=5.365 $Y=1.32
+ $X2=0 $Y2=0
cc_327 N_A_27_47#_c_292_n N_A_211_363#_c_843_n 0.00111403f $X=7.225 $Y=1.32
+ $X2=0 $Y2=0
cc_328 N_A_27_47#_c_295_n N_A_211_363#_c_844_n 0.00679553f $X=0.965 $Y=1.74
+ $X2=0 $Y2=0
cc_329 N_A_27_47#_M1001_g N_A_211_363#_c_844_n 0.0252255f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_287_n N_A_211_363#_c_844_n 0.00946411f $X=0.665 $Y=0.72
+ $X2=0 $Y2=0
cc_331 N_A_27_47#_c_289_n N_A_211_363#_c_844_n 0.0495956f $X=0.78 $Y=1.085 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_400_p N_A_211_363#_c_844_n 0.00860964f $X=0.78 $Y=1.795
+ $X2=0 $Y2=0
cc_333 N_A_27_47#_c_290_n N_A_211_363#_c_844_n 0.00939236f $X=0.78 $Y=0.97 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_306_n N_A_211_363#_c_844_n 0.0198063f $X=5.555 $Y=1.87 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_307_n N_A_211_363#_c_844_n 0.00261995f $X=0.925 $Y=1.87
+ $X2=0 $Y2=0
cc_336 N_A_27_47#_M1009_g N_A_211_363#_c_845_n 0.0119703f $X=4.93 $Y=0.415 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_283_n N_A_211_363#_c_845_n 0.00609027f $X=5.365 $Y=1.32
+ $X2=0 $Y2=0
cc_338 N_A_27_47#_c_310_n N_A_211_363#_c_845_n 0.00398178f $X=5.7 $Y=1.87 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_293_n N_A_211_363#_c_901_n 0.00152544f $X=7.2 $Y=1.41 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_M1009_g N_A_211_363#_c_846_n 0.0163791f $X=4.93 $Y=0.415 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_c_283_n N_A_211_363#_c_846_n 0.0211553f $X=5.365 $Y=1.32 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_299_n N_A_211_363#_c_846_n 5.43883e-19 $X=5.465 $Y=1.99
+ $X2=0 $Y2=0
cc_343 N_A_27_47#_c_310_n N_A_211_363#_c_846_n 6.38247e-19 $X=5.7 $Y=1.87 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_M1038_g N_A_211_363#_c_847_n 0.0118259f $X=8 $Y=0.415 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_292_n N_A_211_363#_c_847_n 0.0234243f $X=7.225 $Y=1.32 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_293_n N_A_211_363#_c_847_n 3.7895e-19 $X=7.2 $Y=1.41 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_308_n N_A_1179_183#_M1025_d 0.00523078f $X=7.115 $Y=1.87
+ $X2=0 $Y2=0
cc_348 N_A_27_47#_c_283_n N_A_1179_183#_c_1040_n 0.0116665f $X=5.365 $Y=1.32
+ $X2=0 $Y2=0
cc_349 N_A_27_47#_c_299_n N_A_1179_183#_c_1040_n 0.0209627f $X=5.465 $Y=1.99
+ $X2=0 $Y2=0
cc_350 N_A_27_47#_c_308_n N_A_1179_183#_c_1040_n 0.00150072f $X=7.115 $Y=1.87
+ $X2=0 $Y2=0
cc_351 N_A_27_47#_c_309_n N_A_1179_183#_c_1040_n 7.30561e-19 $X=5.845 $Y=1.87
+ $X2=0 $Y2=0
cc_352 N_A_27_47#_c_310_n N_A_1179_183#_c_1040_n 0.00212256f $X=5.7 $Y=1.87
+ $X2=0 $Y2=0
cc_353 N_A_27_47#_c_299_n N_A_1179_183#_c_1048_n 0.0264165f $X=5.465 $Y=1.99
+ $X2=0 $Y2=0
cc_354 N_A_27_47#_c_308_n N_A_1179_183#_c_1048_n 0.00126931f $X=7.115 $Y=1.87
+ $X2=0 $Y2=0
cc_355 N_A_27_47#_c_309_n N_A_1179_183#_c_1048_n 7.78138e-19 $X=5.845 $Y=1.87
+ $X2=0 $Y2=0
cc_356 N_A_27_47#_c_301_n N_A_1179_183#_c_1059_n 0.00554009f $X=7.23 $Y=1.99
+ $X2=0 $Y2=0
cc_357 N_A_27_47#_c_308_n N_A_1179_183#_c_1059_n 0.00261642f $X=7.115 $Y=1.87
+ $X2=0 $Y2=0
cc_358 N_A_27_47#_c_300_n N_A_1179_183#_c_1045_n 0.00121845f $X=7.23 $Y=1.89
+ $X2=0 $Y2=0
cc_359 N_A_27_47#_c_301_n N_A_1179_183#_c_1045_n 0.00368889f $X=7.23 $Y=1.99
+ $X2=0 $Y2=0
cc_360 N_A_27_47#_c_308_n N_A_1179_183#_c_1045_n 0.0240109f $X=7.115 $Y=1.87
+ $X2=0 $Y2=0
cc_361 N_A_27_47#_c_311_n N_A_1179_183#_c_1045_n 0.00301429f $X=7.26 $Y=1.87
+ $X2=0 $Y2=0
cc_362 N_A_27_47#_c_292_n N_A_1179_183#_c_1045_n 0.00232864f $X=7.225 $Y=1.32
+ $X2=0 $Y2=0
cc_363 N_A_27_47#_c_293_n N_A_1179_183#_c_1045_n 0.0533394f $X=7.2 $Y=1.41 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_292_n N_A_1001_47#_c_1140_n 0.0159377f $X=7.225 $Y=1.32
+ $X2=0 $Y2=0
cc_365 N_A_27_47#_c_293_n N_A_1001_47#_c_1140_n 3.02222e-19 $X=7.2 $Y=1.41 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_300_n N_A_1001_47#_c_1147_n 0.0117884f $X=7.23 $Y=1.89 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_301_n N_A_1001_47#_c_1147_n 0.0139731f $X=7.23 $Y=1.99 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_308_n N_A_1001_47#_c_1147_n 0.00642704f $X=7.115 $Y=1.87
+ $X2=0 $Y2=0
cc_369 N_A_27_47#_c_293_n N_A_1001_47#_c_1147_n 6.30062e-19 $X=7.2 $Y=1.41 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_c_308_n N_A_1001_47#_c_1143_n 0.00109659f $X=7.115 $Y=1.87
+ $X2=0 $Y2=0
cc_371 N_A_27_47#_c_300_n N_A_1001_47#_c_1144_n 0.00314415f $X=7.23 $Y=1.89
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_c_308_n N_A_1001_47#_c_1144_n 2.82791e-19 $X=7.115 $Y=1.87
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_293_n N_A_1001_47#_c_1144_n 2.11637e-19 $X=7.2 $Y=1.41 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_c_299_n N_A_1001_47#_c_1162_n 0.0105456f $X=5.465 $Y=1.99
+ $X2=0 $Y2=0
cc_375 N_A_27_47#_c_306_n N_A_1001_47#_c_1162_n 0.00761843f $X=5.555 $Y=1.87
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_c_308_n N_A_1001_47#_c_1162_n 0.00373305f $X=7.115 $Y=1.87
+ $X2=0 $Y2=0
cc_377 N_A_27_47#_c_309_n N_A_1001_47#_c_1162_n 0.00172919f $X=5.845 $Y=1.87
+ $X2=0 $Y2=0
cc_378 N_A_27_47#_c_310_n N_A_1001_47#_c_1162_n 0.0280962f $X=5.7 $Y=1.87 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_M1009_g N_A_1001_47#_c_1167_n 0.00154152f $X=4.93 $Y=0.415
+ $X2=0 $Y2=0
cc_380 N_A_27_47#_c_283_n N_A_1001_47#_c_1145_n 8.60771e-19 $X=5.365 $Y=1.32
+ $X2=0 $Y2=0
cc_381 N_A_27_47#_c_299_n N_A_1001_47#_c_1150_n 0.00172804f $X=5.465 $Y=1.99
+ $X2=0 $Y2=0
cc_382 N_A_27_47#_c_308_n N_A_1001_47#_c_1150_n 0.0228785f $X=7.115 $Y=1.87
+ $X2=0 $Y2=0
cc_383 N_A_27_47#_c_309_n N_A_1001_47#_c_1150_n 0.00260208f $X=5.845 $Y=1.87
+ $X2=0 $Y2=0
cc_384 N_A_27_47#_c_310_n N_A_1001_47#_c_1150_n 0.0253723f $X=5.7 $Y=1.87 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_283_n N_A_1001_47#_c_1146_n 0.00241105f $X=5.365 $Y=1.32
+ $X2=0 $Y2=0
cc_386 N_A_27_47#_c_298_n N_A_1001_47#_c_1146_n 4.58825e-19 $X=5.465 $Y=1.575
+ $X2=0 $Y2=0
cc_387 N_A_27_47#_c_308_n N_A_1001_47#_c_1146_n 0.0173913f $X=7.115 $Y=1.87
+ $X2=0 $Y2=0
cc_388 N_A_27_47#_c_309_n N_A_1001_47#_c_1146_n 0.00179088f $X=5.845 $Y=1.87
+ $X2=0 $Y2=0
cc_389 N_A_27_47#_c_310_n N_A_1001_47#_c_1146_n 0.00980238f $X=5.7 $Y=1.87 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_M1038_g N_A_1653_315#_M1024_g 0.0411339f $X=8 $Y=0.415 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_c_301_n N_A_1464_413#_c_1384_n 0.00454762f $X=7.23 $Y=1.99
+ $X2=0 $Y2=0
cc_392 N_A_27_47#_c_311_n N_A_1464_413#_c_1384_n 0.00257575f $X=7.26 $Y=1.87
+ $X2=0 $Y2=0
cc_393 N_A_27_47#_c_292_n N_A_1464_413#_c_1384_n 4.94934e-19 $X=7.225 $Y=1.32
+ $X2=0 $Y2=0
cc_394 N_A_27_47#_c_293_n N_A_1464_413#_c_1384_n 0.0045378f $X=7.2 $Y=1.41 $X2=0
+ $Y2=0
cc_395 N_A_27_47#_M1038_g N_A_1464_413#_c_1388_n 0.00871365f $X=8 $Y=0.415 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_M1038_g N_A_1464_413#_c_1375_n 3.40832e-19 $X=8 $Y=0.415 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_c_285_n N_A_1464_413#_c_1376_n 0.00740284f $X=7.925 $Y=1.32
+ $X2=0 $Y2=0
cc_398 N_A_27_47#_M1038_g N_A_1464_413#_c_1376_n 0.00740571f $X=8 $Y=0.415 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_M1038_g N_A_1464_413#_c_1377_n 0.0136883f $X=8 $Y=0.415 $X2=0
+ $Y2=0
cc_400 N_A_27_47#_c_400_p N_VPWR_M1010_d 7.14517e-19 $X=0.78 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_401 N_A_27_47#_c_307_n N_VPWR_M1010_d 0.001801f $X=0.925 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_402 N_A_27_47#_c_308_n N_VPWR_M1000_d 0.00711371f $X=7.115 $Y=1.87 $X2=0
+ $Y2=0
cc_403 N_A_27_47#_c_295_n N_VPWR_c_1518_n 0.00966647f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_404 N_A_27_47#_c_303_n N_VPWR_c_1518_n 0.00676847f $X=0.665 $Y=1.88 $X2=0
+ $Y2=0
cc_405 N_A_27_47#_c_400_p N_VPWR_c_1518_n 0.0133392f $X=0.78 $Y=1.795 $X2=0
+ $Y2=0
cc_406 N_A_27_47#_c_305_n N_VPWR_c_1518_n 0.0246493f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_407 N_A_27_47#_c_307_n N_VPWR_c_1518_n 0.00311184f $X=0.925 $Y=1.87 $X2=0
+ $Y2=0
cc_408 N_A_27_47#_c_306_n N_VPWR_c_1519_n 0.00142334f $X=5.555 $Y=1.87 $X2=0
+ $Y2=0
cc_409 N_A_27_47#_c_306_n N_VPWR_c_1520_n 8.00522e-19 $X=5.555 $Y=1.87 $X2=0
+ $Y2=0
cc_410 N_A_27_47#_c_308_n N_VPWR_c_1521_n 0.00944753f $X=7.115 $Y=1.87 $X2=0
+ $Y2=0
cc_411 N_A_27_47#_c_299_n N_VPWR_c_1531_n 0.00454633f $X=5.465 $Y=1.99 $X2=0
+ $Y2=0
cc_412 N_A_27_47#_c_301_n N_VPWR_c_1533_n 0.00519523f $X=7.23 $Y=1.99 $X2=0
+ $Y2=0
cc_413 N_A_27_47#_c_293_n N_VPWR_c_1533_n 0.00157744f $X=7.2 $Y=1.41 $X2=0 $Y2=0
cc_414 N_A_27_47#_c_303_n N_VPWR_c_1535_n 0.00180073f $X=0.665 $Y=1.88 $X2=0
+ $Y2=0
cc_415 N_A_27_47#_c_305_n N_VPWR_c_1535_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_416 N_A_27_47#_c_295_n N_VPWR_c_1536_n 0.00590576f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_417 N_A_27_47#_c_295_n N_VPWR_c_1517_n 0.00664518f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_c_299_n N_VPWR_c_1517_n 0.00640619f $X=5.465 $Y=1.99 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_c_301_n N_VPWR_c_1517_n 0.00675888f $X=7.23 $Y=1.99 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_c_303_n N_VPWR_c_1517_n 0.00427626f $X=0.665 $Y=1.88 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_c_305_n N_VPWR_c_1517_n 0.00646745f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_c_306_n N_VPWR_c_1517_n 0.215775f $X=5.555 $Y=1.87 $X2=0 $Y2=0
cc_423 N_A_27_47#_c_307_n N_VPWR_c_1517_n 0.0146104f $X=0.925 $Y=1.87 $X2=0
+ $Y2=0
cc_424 N_A_27_47#_c_308_n N_VPWR_c_1517_n 0.0602887f $X=7.115 $Y=1.87 $X2=0
+ $Y2=0
cc_425 N_A_27_47#_c_309_n N_VPWR_c_1517_n 0.014713f $X=5.845 $Y=1.87 $X2=0 $Y2=0
cc_426 N_A_27_47#_c_311_n N_VPWR_c_1517_n 0.0158133f $X=7.26 $Y=1.87 $X2=0 $Y2=0
cc_427 N_A_27_47#_c_293_n N_VPWR_c_1517_n 0.0010813f $X=7.2 $Y=1.41 $X2=0 $Y2=0
cc_428 N_A_27_47#_c_306_n N_A_604_369#_c_1727_n 0.00614591f $X=5.555 $Y=1.87
+ $X2=0 $Y2=0
cc_429 N_A_27_47#_c_306_n N_A_604_369#_c_1723_n 0.0232744f $X=5.555 $Y=1.87
+ $X2=0 $Y2=0
cc_430 N_A_27_47#_c_306_n N_A_604_369#_c_1724_n 0.0102316f $X=5.555 $Y=1.87
+ $X2=0 $Y2=0
cc_431 N_A_27_47#_M1009_g N_A_604_369#_c_1719_n 0.00473651f $X=4.93 $Y=0.415
+ $X2=0 $Y2=0
cc_432 N_A_27_47#_M1009_g N_A_604_369#_c_1720_n 0.00646253f $X=4.93 $Y=0.415
+ $X2=0 $Y2=0
cc_433 N_A_27_47#_c_306_n N_A_604_369#_c_1720_n 0.0104876f $X=5.555 $Y=1.87
+ $X2=0 $Y2=0
cc_434 N_A_27_47#_M1009_g N_A_604_369#_c_1721_n 0.00160472f $X=4.93 $Y=0.415
+ $X2=0 $Y2=0
cc_435 N_A_27_47#_M1009_g N_A_604_369#_c_1722_n 0.00136206f $X=4.93 $Y=0.415
+ $X2=0 $Y2=0
cc_436 N_A_27_47#_c_306_n N_A_604_369#_c_1726_n 0.0128459f $X=5.555 $Y=1.87
+ $X2=0 $Y2=0
cc_437 N_A_27_47#_c_310_n N_A_604_369#_c_1726_n 0.00293569f $X=5.7 $Y=1.87 $X2=0
+ $Y2=0
cc_438 N_A_27_47#_c_306_n A_698_369# 0.00134881f $X=5.555 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_439 N_A_27_47#_c_287_n N_VGND_M1029_d 0.00226918f $X=0.665 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_440 N_A_27_47#_M1009_g N_VGND_c_1881_n 0.00353857f $X=4.93 $Y=0.415 $X2=0
+ $Y2=0
cc_441 N_A_27_47#_M1038_g N_VGND_c_1883_n 0.00230088f $X=8 $Y=0.415 $X2=0 $Y2=0
cc_442 N_A_27_47#_M1001_g N_VGND_c_1890_n 0.00585385f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_443 N_A_27_47#_c_511_p N_VGND_c_1894_n 0.00725596f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_444 N_A_27_47#_c_287_n N_VGND_c_1894_n 0.00244154f $X=0.665 $Y=0.72 $X2=0
+ $Y2=0
cc_445 N_A_27_47#_M1009_g N_VGND_c_1895_n 0.00431421f $X=4.93 $Y=0.415 $X2=0
+ $Y2=0
cc_446 N_A_27_47#_M1038_g N_VGND_c_1896_n 0.00379633f $X=8 $Y=0.415 $X2=0 $Y2=0
cc_447 N_A_27_47#_M1001_g N_VGND_c_1900_n 0.00317372f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_448 N_A_27_47#_c_511_p N_VGND_c_1900_n 0.00895866f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_449 N_A_27_47#_c_287_n N_VGND_c_1900_n 0.0228245f $X=0.665 $Y=0.72 $X2=0
+ $Y2=0
cc_450 N_A_27_47#_c_291_n N_VGND_c_1900_n 6.84019e-19 $X=0.99 $Y=1.235 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_M1029_s N_VGND_c_1906_n 0.00437169f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_452 N_A_27_47#_M1001_g N_VGND_c_1906_n 0.0098507f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_453 N_A_27_47#_M1009_g N_VGND_c_1906_n 0.00680361f $X=4.93 $Y=0.415 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_M1038_g N_VGND_c_1906_n 0.00610845f $X=8 $Y=0.415 $X2=0 $Y2=0
cc_455 N_A_27_47#_c_511_p N_VGND_c_1906_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_c_287_n N_VGND_c_1906_n 0.00609319f $X=0.665 $Y=0.72 $X2=0
+ $Y2=0
cc_457 N_A_319_47#_c_526_n N_SCE_c_652_n 0.0082304f $X=1.605 $Y=1.86 $X2=-0.19
+ $Y2=-0.24
cc_458 N_A_319_47#_c_534_n N_SCE_c_652_n 0.00582986f $X=1.72 $Y=2.175 $X2=-0.19
+ $Y2=-0.24
cc_459 N_A_319_47#_c_541_n N_SCE_c_652_n 0.0213633f $X=2.25 $Y=1.967 $X2=-0.19
+ $Y2=-0.24
cc_460 N_A_319_47#_c_527_n N_SCE_c_652_n 0.0031289f $X=2.335 $Y=1.86 $X2=-0.19
+ $Y2=-0.24
cc_461 N_A_319_47#_c_537_n N_SCE_c_652_n 8.40582e-19 $X=1.662 $Y=1.967 $X2=-0.19
+ $Y2=-0.24
cc_462 N_A_319_47#_M1031_g N_SCE_M1021_g 0.016781f $X=2.57 $Y=0.445 $X2=0 $Y2=0
cc_463 N_A_319_47#_c_526_n N_SCE_M1021_g 0.00802403f $X=1.605 $Y=1.86 $X2=0
+ $Y2=0
cc_464 N_A_319_47#_c_527_n N_SCE_M1021_g 0.00399271f $X=2.335 $Y=1.86 $X2=0
+ $Y2=0
cc_465 N_A_319_47#_c_528_n N_SCE_M1021_g 0.00106798f $X=2.42 $Y=1.04 $X2=0 $Y2=0
cc_466 N_A_319_47#_c_531_n N_SCE_M1021_g 0.0124737f $X=2.57 $Y=1.04 $X2=0 $Y2=0
cc_467 N_A_319_47#_c_527_n N_SCE_c_654_n 0.00655628f $X=2.335 $Y=1.86 $X2=0
+ $Y2=0
cc_468 N_A_319_47#_c_531_n N_SCE_c_654_n 0.0081608f $X=2.57 $Y=1.04 $X2=0 $Y2=0
cc_469 N_A_319_47#_c_527_n N_SCE_c_655_n 0.00275035f $X=2.335 $Y=1.86 $X2=0
+ $Y2=0
cc_470 N_A_319_47#_c_543_n N_SCE_c_655_n 0.00894721f $X=3.335 $Y=1.967 $X2=0
+ $Y2=0
cc_471 N_A_319_47#_c_547_n N_SCE_c_655_n 0.00611955f $X=2.335 $Y=1.967 $X2=0
+ $Y2=0
cc_472 N_A_319_47#_c_527_n N_SCE_c_656_n 0.00763267f $X=2.335 $Y=1.86 $X2=0
+ $Y2=0
cc_473 N_A_319_47#_c_529_n N_SCE_c_656_n 6.87639e-19 $X=2.48 $Y=1.04 $X2=0 $Y2=0
cc_474 N_A_319_47#_c_543_n N_SCE_c_656_n 2.9076e-19 $X=3.335 $Y=1.967 $X2=0
+ $Y2=0
cc_475 N_A_319_47#_M1031_g N_SCE_c_647_n 6.40825e-19 $X=2.57 $Y=0.445 $X2=0
+ $Y2=0
cc_476 N_A_319_47#_c_526_n N_SCE_c_647_n 0.066591f $X=1.605 $Y=1.86 $X2=0 $Y2=0
cc_477 N_A_319_47#_c_541_n N_SCE_c_647_n 0.0106871f $X=2.25 $Y=1.967 $X2=0 $Y2=0
cc_478 N_A_319_47#_c_527_n N_SCE_c_647_n 0.0323992f $X=2.335 $Y=1.86 $X2=0 $Y2=0
cc_479 N_A_319_47#_c_528_n N_SCE_c_647_n 0.0109125f $X=2.42 $Y=1.04 $X2=0 $Y2=0
cc_480 N_A_319_47#_c_531_n N_SCE_c_647_n 5.75109e-19 $X=2.57 $Y=1.04 $X2=0 $Y2=0
cc_481 N_A_319_47#_M1031_g N_SCE_c_648_n 0.0120677f $X=2.57 $Y=0.445 $X2=0 $Y2=0
cc_482 N_A_319_47#_c_528_n N_SCE_c_648_n 0.0130764f $X=2.42 $Y=1.04 $X2=0 $Y2=0
cc_483 N_A_319_47#_c_529_n N_SCE_c_648_n 0.0182303f $X=2.48 $Y=1.04 $X2=0 $Y2=0
cc_484 N_A_319_47#_c_531_n N_SCE_c_648_n 0.00410724f $X=2.57 $Y=1.04 $X2=0 $Y2=0
cc_485 N_A_319_47#_c_526_n N_SCE_c_649_n 0.0123907f $X=1.605 $Y=1.86 $X2=0 $Y2=0
cc_486 N_A_319_47#_c_532_n N_SCE_c_650_n 0.0173476f $X=3.4 $Y=1.77 $X2=0 $Y2=0
cc_487 N_A_319_47#_c_538_n N_SCE_c_650_n 4.0176e-19 $X=3.42 $Y=1.52 $X2=0 $Y2=0
cc_488 N_A_319_47#_c_532_n SCE 4.01315e-19 $X=3.4 $Y=1.77 $X2=0 $Y2=0
cc_489 N_A_319_47#_c_529_n SCE 0.00470053f $X=2.48 $Y=1.04 $X2=0 $Y2=0
cc_490 N_A_319_47#_c_538_n SCE 0.0124391f $X=3.42 $Y=1.52 $X2=0 $Y2=0
cc_491 N_A_319_47#_c_532_n N_D_c_749_n 0.0473597f $X=3.4 $Y=1.77 $X2=-0.19
+ $Y2=-0.24
cc_492 N_A_319_47#_c_527_n N_D_c_749_n 0.00182775f $X=2.335 $Y=1.86 $X2=-0.19
+ $Y2=-0.24
cc_493 N_A_319_47#_c_543_n N_D_c_749_n 0.0163489f $X=3.335 $Y=1.967 $X2=-0.19
+ $Y2=-0.24
cc_494 N_A_319_47#_c_536_n N_D_c_749_n 0.00121919f $X=3.432 $Y=1.86 $X2=-0.19
+ $Y2=-0.24
cc_495 N_A_319_47#_c_538_n N_D_c_749_n 3.48252e-19 $X=3.42 $Y=1.52 $X2=-0.19
+ $Y2=-0.24
cc_496 N_A_319_47#_M1031_g N_D_M1014_g 0.0537503f $X=2.57 $Y=0.445 $X2=0 $Y2=0
cc_497 N_A_319_47#_c_527_n N_D_M1014_g 0.00461931f $X=2.335 $Y=1.86 $X2=0 $Y2=0
cc_498 N_A_319_47#_c_529_n N_D_M1014_g 0.00191253f $X=2.48 $Y=1.04 $X2=0 $Y2=0
cc_499 N_A_319_47#_c_532_n D 0.00208935f $X=3.4 $Y=1.77 $X2=0 $Y2=0
cc_500 N_A_319_47#_c_527_n D 0.0143404f $X=2.335 $Y=1.86 $X2=0 $Y2=0
cc_501 N_A_319_47#_c_543_n D 0.0209635f $X=3.335 $Y=1.967 $X2=0 $Y2=0
cc_502 N_A_319_47#_c_538_n D 0.021827f $X=3.42 $Y=1.52 $X2=0 $Y2=0
cc_503 N_A_319_47#_c_532_n N_SCD_c_789_n 0.0337266f $X=3.4 $Y=1.77 $X2=0 $Y2=0
cc_504 N_A_319_47#_c_543_n N_SCD_c_789_n 2.18774e-19 $X=3.335 $Y=1.967 $X2=0
+ $Y2=0
cc_505 N_A_319_47#_c_536_n N_SCD_c_789_n 0.00255837f $X=3.432 $Y=1.86 $X2=0
+ $Y2=0
cc_506 N_A_319_47#_c_532_n SCD 0.00107609f $X=3.4 $Y=1.77 $X2=0 $Y2=0
cc_507 N_A_319_47#_c_538_n SCD 0.0161232f $X=3.42 $Y=1.52 $X2=0 $Y2=0
cc_508 N_A_319_47#_c_532_n N_SCD_c_787_n 0.0199907f $X=3.4 $Y=1.77 $X2=0 $Y2=0
cc_509 N_A_319_47#_c_538_n N_SCD_c_787_n 0.00110894f $X=3.42 $Y=1.52 $X2=0 $Y2=0
cc_510 N_A_319_47#_M1021_s N_A_211_363#_c_840_n 0.00682674f $X=1.595 $Y=0.235
+ $X2=0 $Y2=0
cc_511 N_A_319_47#_M1031_g N_A_211_363#_c_840_n 0.00386001f $X=2.57 $Y=0.445
+ $X2=0 $Y2=0
cc_512 N_A_319_47#_c_526_n N_A_211_363#_c_840_n 0.0174641f $X=1.605 $Y=1.86
+ $X2=0 $Y2=0
cc_513 N_A_319_47#_c_530_n N_A_211_363#_c_840_n 0.00905429f $X=1.74 $Y=0.36
+ $X2=0 $Y2=0
cc_514 N_A_319_47#_c_526_n N_A_211_363#_c_841_n 0.00136191f $X=1.605 $Y=1.86
+ $X2=0 $Y2=0
cc_515 N_A_319_47#_c_530_n N_A_211_363#_c_841_n 0.00139336f $X=1.74 $Y=0.36
+ $X2=0 $Y2=0
cc_516 N_A_319_47#_c_526_n N_A_211_363#_c_844_n 0.0822487f $X=1.605 $Y=1.86
+ $X2=0 $Y2=0
cc_517 N_A_319_47#_c_534_n N_A_211_363#_c_844_n 0.022567f $X=1.72 $Y=2.175 $X2=0
+ $Y2=0
cc_518 N_A_319_47#_c_530_n N_A_211_363#_c_844_n 0.00554179f $X=1.74 $Y=0.36
+ $X2=0 $Y2=0
cc_519 N_A_319_47#_c_537_n N_A_211_363#_c_844_n 0.0128392f $X=1.662 $Y=1.967
+ $X2=0 $Y2=0
cc_520 N_A_319_47#_c_541_n N_VPWR_M1022_d 0.00402367f $X=2.25 $Y=1.967 $X2=0
+ $Y2=0
cc_521 N_A_319_47#_c_547_n N_VPWR_M1022_d 2.87958e-19 $X=2.335 $Y=1.967 $X2=0
+ $Y2=0
cc_522 N_A_319_47#_c_534_n N_VPWR_c_1519_n 0.015515f $X=1.72 $Y=2.175 $X2=0
+ $Y2=0
cc_523 N_A_319_47#_c_541_n N_VPWR_c_1519_n 0.0152093f $X=2.25 $Y=1.967 $X2=0
+ $Y2=0
cc_524 N_A_319_47#_c_547_n N_VPWR_c_1519_n 0.00353227f $X=2.335 $Y=1.967 $X2=0
+ $Y2=0
cc_525 N_A_319_47#_c_532_n N_VPWR_c_1529_n 0.00441747f $X=3.4 $Y=1.77 $X2=0
+ $Y2=0
cc_526 N_A_319_47#_c_543_n N_VPWR_c_1529_n 0.00685978f $X=3.335 $Y=1.967 $X2=0
+ $Y2=0
cc_527 N_A_319_47#_c_547_n N_VPWR_c_1529_n 0.00112385f $X=2.335 $Y=1.967 $X2=0
+ $Y2=0
cc_528 N_A_319_47#_c_534_n N_VPWR_c_1536_n 0.0176557f $X=1.72 $Y=2.175 $X2=0
+ $Y2=0
cc_529 N_A_319_47#_c_541_n N_VPWR_c_1536_n 0.00234063f $X=2.25 $Y=1.967 $X2=0
+ $Y2=0
cc_530 N_A_319_47#_M1022_s N_VPWR_c_1517_n 0.0019314f $X=1.595 $Y=1.845 $X2=0
+ $Y2=0
cc_531 N_A_319_47#_c_532_n N_VPWR_c_1517_n 0.00617905f $X=3.4 $Y=1.77 $X2=0
+ $Y2=0
cc_532 N_A_319_47#_c_534_n N_VPWR_c_1517_n 0.00512382f $X=1.72 $Y=2.175 $X2=0
+ $Y2=0
cc_533 N_A_319_47#_c_541_n N_VPWR_c_1517_n 0.00257024f $X=2.25 $Y=1.967 $X2=0
+ $Y2=0
cc_534 N_A_319_47#_c_543_n N_VPWR_c_1517_n 0.0062042f $X=3.335 $Y=1.967 $X2=0
+ $Y2=0
cc_535 N_A_319_47#_c_547_n N_VPWR_c_1517_n 0.00109221f $X=2.335 $Y=1.967 $X2=0
+ $Y2=0
cc_536 N_A_319_47#_c_543_n A_503_369# 0.00701041f $X=3.335 $Y=1.967 $X2=-0.19
+ $Y2=-0.24
cc_537 N_A_319_47#_c_543_n N_A_604_369#_M1020_d 0.00423765f $X=3.335 $Y=1.967
+ $X2=0 $Y2=0
cc_538 N_A_319_47#_c_532_n N_A_604_369#_c_1727_n 0.0107746f $X=3.4 $Y=1.77 $X2=0
+ $Y2=0
cc_539 N_A_319_47#_c_543_n N_A_604_369#_c_1727_n 0.0322478f $X=3.335 $Y=1.967
+ $X2=0 $Y2=0
cc_540 N_A_319_47#_M1031_g N_A_604_369#_c_1740_n 4.80357e-19 $X=2.57 $Y=0.445
+ $X2=0 $Y2=0
cc_541 N_A_319_47#_c_532_n N_A_604_369#_c_1741_n 0.00368652f $X=3.4 $Y=1.77
+ $X2=0 $Y2=0
cc_542 N_A_319_47#_c_532_n N_A_604_369#_c_1724_n 5.35252e-19 $X=3.4 $Y=1.77
+ $X2=0 $Y2=0
cc_543 N_A_319_47#_c_543_n N_A_604_369#_c_1724_n 0.00683184f $X=3.335 $Y=1.967
+ $X2=0 $Y2=0
cc_544 N_A_319_47#_c_536_n N_A_604_369#_c_1724_n 0.00221871f $X=3.432 $Y=1.86
+ $X2=0 $Y2=0
cc_545 N_A_319_47#_M1031_g N_VGND_c_1880_n 0.00333207f $X=2.57 $Y=0.445 $X2=0
+ $Y2=0
cc_546 N_A_319_47#_c_530_n N_VGND_c_1880_n 0.0121274f $X=1.74 $Y=0.36 $X2=0
+ $Y2=0
cc_547 N_A_319_47#_c_530_n N_VGND_c_1890_n 0.0230378f $X=1.74 $Y=0.36 $X2=0
+ $Y2=0
cc_548 N_A_319_47#_M1031_g N_VGND_c_1892_n 0.00422112f $X=2.57 $Y=0.445 $X2=0
+ $Y2=0
cc_549 N_A_319_47#_M1021_s N_VGND_c_1906_n 0.0014225f $X=1.595 $Y=0.235 $X2=0
+ $Y2=0
cc_550 N_A_319_47#_M1031_g N_VGND_c_1906_n 0.00514507f $X=2.57 $Y=0.445 $X2=0
+ $Y2=0
cc_551 N_A_319_47#_c_530_n N_VGND_c_1906_n 0.00372846f $X=1.74 $Y=0.36 $X2=0
+ $Y2=0
cc_552 N_SCE_c_652_n N_D_c_749_n 0.0015819f $X=1.955 $Y=1.77 $X2=-0.19 $Y2=-0.24
cc_553 N_SCE_M1021_g N_D_c_749_n 2.78202e-19 $X=1.98 $Y=0.445 $X2=-0.19
+ $Y2=-0.24
cc_554 N_SCE_c_655_n N_D_c_749_n 0.0337703f $X=2.425 $Y=1.77 $X2=-0.19 $Y2=-0.24
cc_555 N_SCE_c_656_n N_D_c_749_n 0.0142795f $X=2.425 $Y=1.58 $X2=-0.19 $Y2=-0.24
cc_556 N_SCE_c_648_n N_D_c_749_n 0.00298034f $X=3.315 $Y=0.7 $X2=-0.19 $Y2=-0.24
cc_557 N_SCE_M1019_g N_D_M1014_g 0.0117825f $X=3.51 $Y=0.445 $X2=0 $Y2=0
cc_558 N_SCE_c_648_n N_D_M1014_g 0.0137087f $X=3.315 $Y=0.7 $X2=0 $Y2=0
cc_559 N_SCE_c_650_n N_D_M1014_g 0.0208345f $X=3.51 $Y=0.95 $X2=0 $Y2=0
cc_560 SCE N_D_M1014_g 0.00157285f $X=3.45 $Y=0.85 $X2=0 $Y2=0
cc_561 N_SCE_c_656_n D 7.72287e-19 $X=2.425 $Y=1.58 $X2=0 $Y2=0
cc_562 N_SCE_c_648_n D 0.010785f $X=3.315 $Y=0.7 $X2=0 $Y2=0
cc_563 N_SCE_M1019_g N_SCD_M1037_g 0.057552f $X=3.51 $Y=0.445 $X2=0 $Y2=0
cc_564 SCE N_SCD_M1037_g 0.00126634f $X=3.45 $Y=0.85 $X2=0 $Y2=0
cc_565 N_SCE_c_650_n SCD 2.22853e-19 $X=3.51 $Y=0.95 $X2=0 $Y2=0
cc_566 SCE SCD 0.0030443f $X=3.45 $Y=0.85 $X2=0 $Y2=0
cc_567 N_SCE_M1021_g N_A_211_363#_c_840_n 0.00434342f $X=1.98 $Y=0.445 $X2=0
+ $Y2=0
cc_568 N_SCE_M1019_g N_A_211_363#_c_840_n 0.00376966f $X=3.51 $Y=0.445 $X2=0
+ $Y2=0
cc_569 N_SCE_c_648_n N_A_211_363#_c_840_n 0.0405406f $X=3.315 $Y=0.7 $X2=0 $Y2=0
cc_570 N_SCE_c_649_n N_A_211_363#_c_840_n 0.00558867f $X=2.03 $Y=0.7 $X2=0 $Y2=0
cc_571 N_SCE_c_716_p N_A_211_363#_c_840_n 0.00624733f $X=3.425 $Y=0.785 $X2=0
+ $Y2=0
cc_572 N_SCE_c_652_n N_A_211_363#_c_844_n 0.00157278f $X=1.955 $Y=1.77 $X2=0
+ $Y2=0
cc_573 N_SCE_c_652_n N_VPWR_c_1519_n 0.0118271f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_574 N_SCE_c_654_n N_VPWR_c_1519_n 3.93315e-19 $X=2.325 $Y=1.58 $X2=0 $Y2=0
cc_575 N_SCE_c_655_n N_VPWR_c_1519_n 0.00940281f $X=2.425 $Y=1.77 $X2=0 $Y2=0
cc_576 N_SCE_c_655_n N_VPWR_c_1529_n 0.00454221f $X=2.425 $Y=1.77 $X2=0 $Y2=0
cc_577 N_SCE_c_652_n N_VPWR_c_1536_n 0.00312096f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_578 N_SCE_c_652_n N_VPWR_c_1517_n 0.00489637f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_579 N_SCE_c_655_n N_VPWR_c_1517_n 0.0050148f $X=2.425 $Y=1.77 $X2=0 $Y2=0
cc_580 N_SCE_c_648_n N_A_604_369#_M1014_d 0.00189963f $X=3.315 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_581 N_SCE_c_716_p N_A_604_369#_M1014_d 6.01405e-19 $X=3.425 $Y=0.785
+ $X2=-0.19 $Y2=-0.24
cc_582 N_SCE_c_655_n N_A_604_369#_c_1727_n 6.13327e-19 $X=2.425 $Y=1.77 $X2=0
+ $Y2=0
cc_583 N_SCE_M1019_g N_A_604_369#_c_1740_n 0.00733119f $X=3.51 $Y=0.445 $X2=0
+ $Y2=0
cc_584 N_SCE_c_648_n N_A_604_369#_c_1740_n 0.014004f $X=3.315 $Y=0.7 $X2=0 $Y2=0
cc_585 N_SCE_c_650_n N_A_604_369#_c_1740_n 4.69407e-19 $X=3.51 $Y=0.95 $X2=0
+ $Y2=0
cc_586 N_SCE_c_716_p N_A_604_369#_c_1740_n 0.0117118f $X=3.425 $Y=0.785 $X2=0
+ $Y2=0
cc_587 N_SCE_M1019_g N_A_604_369#_c_1716_n 0.00363713f $X=3.51 $Y=0.445 $X2=0
+ $Y2=0
cc_588 N_SCE_c_716_p N_A_604_369#_c_1716_n 0.00790081f $X=3.425 $Y=0.785 $X2=0
+ $Y2=0
cc_589 N_SCE_M1019_g N_A_604_369#_c_1718_n 0.0011534f $X=3.51 $Y=0.445 $X2=0
+ $Y2=0
cc_590 N_SCE_c_716_p N_A_604_369#_c_1718_n 0.00619806f $X=3.425 $Y=0.785 $X2=0
+ $Y2=0
cc_591 SCE N_A_604_369#_c_1718_n 0.00817005f $X=3.45 $Y=0.85 $X2=0 $Y2=0
cc_592 N_SCE_c_648_n N_VGND_M1021_d 0.0034102f $X=3.315 $Y=0.7 $X2=0 $Y2=0
cc_593 N_SCE_M1021_g N_VGND_c_1880_n 0.00527118f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_594 N_SCE_c_648_n N_VGND_c_1880_n 0.0192779f $X=3.315 $Y=0.7 $X2=0 $Y2=0
cc_595 N_SCE_M1021_g N_VGND_c_1890_n 0.00421987f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_596 N_SCE_c_648_n N_VGND_c_1890_n 0.00149634f $X=3.315 $Y=0.7 $X2=0 $Y2=0
cc_597 N_SCE_c_649_n N_VGND_c_1890_n 0.00208705f $X=2.03 $Y=0.7 $X2=0 $Y2=0
cc_598 N_SCE_M1019_g N_VGND_c_1892_n 0.00362032f $X=3.51 $Y=0.445 $X2=0 $Y2=0
cc_599 N_SCE_c_648_n N_VGND_c_1892_n 0.00830546f $X=3.315 $Y=0.7 $X2=0 $Y2=0
cc_600 N_SCE_M1021_g N_VGND_c_1906_n 0.00665851f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_601 N_SCE_M1019_g N_VGND_c_1906_n 0.00492794f $X=3.51 $Y=0.445 $X2=0 $Y2=0
cc_602 N_SCE_c_648_n A_529_47# 0.00220129f $X=3.315 $Y=0.7 $X2=-0.19 $Y2=-0.24
cc_603 N_D_M1014_g N_A_211_363#_c_840_n 0.00371598f $X=2.98 $Y=0.445 $X2=0 $Y2=0
cc_604 N_D_c_749_n N_VPWR_c_1519_n 0.0017204f $X=2.93 $Y=1.77 $X2=0 $Y2=0
cc_605 N_D_c_749_n N_VPWR_c_1529_n 0.00455384f $X=2.93 $Y=1.77 $X2=0 $Y2=0
cc_606 N_D_c_749_n N_VPWR_c_1517_n 0.00624738f $X=2.93 $Y=1.77 $X2=0 $Y2=0
cc_607 N_D_c_749_n N_A_604_369#_c_1727_n 0.00790861f $X=2.93 $Y=1.77 $X2=0 $Y2=0
cc_608 N_D_M1014_g N_A_604_369#_c_1740_n 0.00274813f $X=2.98 $Y=0.445 $X2=0
+ $Y2=0
cc_609 N_D_M1014_g N_VGND_c_1892_n 0.0042011f $X=2.98 $Y=0.445 $X2=0 $Y2=0
cc_610 N_D_M1014_g N_VGND_c_1906_n 0.00519902f $X=2.98 $Y=0.445 $X2=0 $Y2=0
cc_611 N_SCD_M1037_g N_A_211_363#_c_840_n 0.00364748f $X=3.89 $Y=0.445 $X2=0
+ $Y2=0
cc_612 SCD N_A_211_363#_c_840_n 0.00124159f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_613 N_SCD_c_789_n N_VPWR_c_1520_n 0.00627598f $X=3.915 $Y=1.77 $X2=0 $Y2=0
cc_614 N_SCD_c_789_n N_VPWR_c_1529_n 0.00504444f $X=3.915 $Y=1.77 $X2=0 $Y2=0
cc_615 N_SCD_c_789_n N_VPWR_c_1517_n 0.00784388f $X=3.915 $Y=1.77 $X2=0 $Y2=0
cc_616 N_SCD_c_789_n N_A_604_369#_c_1727_n 0.00520197f $X=3.915 $Y=1.77 $X2=0
+ $Y2=0
cc_617 N_SCD_M1037_g N_A_604_369#_c_1740_n 0.00466603f $X=3.89 $Y=0.445 $X2=0
+ $Y2=0
cc_618 N_SCD_c_789_n N_A_604_369#_c_1741_n 0.00716226f $X=3.915 $Y=1.77 $X2=0
+ $Y2=0
cc_619 N_SCD_M1037_g N_A_604_369#_c_1716_n 0.00621204f $X=3.89 $Y=0.445 $X2=0
+ $Y2=0
cc_620 N_SCD_c_789_n N_A_604_369#_c_1723_n 0.0107892f $X=3.915 $Y=1.77 $X2=0
+ $Y2=0
cc_621 SCD N_A_604_369#_c_1723_n 0.0333186f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_622 N_SCD_c_787_n N_A_604_369#_c_1723_n 5.47062e-19 $X=3.95 $Y=1.355 $X2=0
+ $Y2=0
cc_623 N_SCD_c_789_n N_A_604_369#_c_1724_n 0.00273267f $X=3.915 $Y=1.77 $X2=0
+ $Y2=0
cc_624 SCD N_A_604_369#_c_1724_n 0.00363458f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_625 N_SCD_M1037_g N_A_604_369#_c_1717_n 0.00869578f $X=3.89 $Y=0.445 $X2=0
+ $Y2=0
cc_626 SCD N_A_604_369#_c_1717_n 0.0368172f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_627 N_SCD_c_787_n N_A_604_369#_c_1717_n 8.52981e-19 $X=3.95 $Y=1.355 $X2=0
+ $Y2=0
cc_628 N_SCD_M1037_g N_A_604_369#_c_1718_n 0.00268499f $X=3.89 $Y=0.445 $X2=0
+ $Y2=0
cc_629 SCD N_A_604_369#_c_1718_n 0.00472161f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_630 N_SCD_M1037_g N_A_604_369#_c_1719_n 0.00234067f $X=3.89 $Y=0.445 $X2=0
+ $Y2=0
cc_631 N_SCD_M1037_g N_A_604_369#_c_1720_n 0.00433743f $X=3.89 $Y=0.445 $X2=0
+ $Y2=0
cc_632 N_SCD_c_788_n N_A_604_369#_c_1720_n 0.00333631f $X=3.915 $Y=1.67 $X2=0
+ $Y2=0
cc_633 N_SCD_c_789_n N_A_604_369#_c_1720_n 0.00109095f $X=3.915 $Y=1.77 $X2=0
+ $Y2=0
cc_634 SCD N_A_604_369#_c_1720_n 0.0494238f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_635 N_SCD_c_787_n N_A_604_369#_c_1720_n 0.00106267f $X=3.95 $Y=1.355 $X2=0
+ $Y2=0
cc_636 N_SCD_c_789_n N_A_604_369#_c_1726_n 0.00296158f $X=3.915 $Y=1.77 $X2=0
+ $Y2=0
cc_637 N_SCD_M1037_g N_VGND_c_1881_n 0.0104431f $X=3.89 $Y=0.445 $X2=0 $Y2=0
cc_638 N_SCD_M1037_g N_VGND_c_1892_n 0.00406622f $X=3.89 $Y=0.445 $X2=0 $Y2=0
cc_639 N_SCD_M1037_g N_VGND_c_1906_n 0.00624566f $X=3.89 $Y=0.445 $X2=0 $Y2=0
cc_640 N_A_211_363#_c_839_n N_A_1179_183#_M1002_d 0.00152085f $X=7.525 $Y=0.87
+ $X2=-0.19 $Y2=-0.24
cc_641 N_A_211_363#_c_843_n N_A_1179_183#_M1002_d 0.00127469f $X=7.125 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_642 N_A_211_363#_c_835_n N_A_1179_183#_M1017_g 0.0138322f $X=5.51 $Y=0.705
+ $X2=0 $Y2=0
cc_643 N_A_211_363#_c_843_n N_A_1179_183#_M1017_g 0.00275613f $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_644 N_A_211_363#_c_843_n N_A_1179_183#_c_1042_n 0.021665f $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_645 N_A_211_363#_c_901_n N_A_1179_183#_c_1072_n 2.22072e-19 $X=7.27 $Y=0.85
+ $X2=0 $Y2=0
cc_646 N_A_211_363#_c_839_n N_A_1179_183#_c_1073_n 0.00717359f $X=7.525 $Y=0.87
+ $X2=0 $Y2=0
cc_647 N_A_211_363#_c_843_n N_A_1179_183#_c_1073_n 0.0048041f $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_648 N_A_211_363#_c_901_n N_A_1179_183#_c_1073_n 4.51578e-19 $X=7.27 $Y=0.85
+ $X2=0 $Y2=0
cc_649 N_A_211_363#_c_843_n N_A_1179_183#_c_1043_n 0.00936146f $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_650 N_A_211_363#_c_838_n N_A_1179_183#_c_1044_n 0.00106902f $X=7.62 $Y=1.575
+ $X2=0 $Y2=0
cc_651 N_A_211_363#_c_839_n N_A_1179_183#_c_1044_n 0.0193507f $X=7.525 $Y=0.87
+ $X2=0 $Y2=0
cc_652 N_A_211_363#_c_843_n N_A_1179_183#_c_1044_n 0.0215929f $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_653 N_A_211_363#_c_901_n N_A_1179_183#_c_1044_n 4.94929e-19 $X=7.27 $Y=0.85
+ $X2=0 $Y2=0
cc_654 N_A_211_363#_c_847_n N_A_1179_183#_c_1044_n 5.8166e-19 $X=7.48 $Y=0.87
+ $X2=0 $Y2=0
cc_655 N_A_211_363#_c_838_n N_A_1179_183#_c_1045_n 0.00592824f $X=7.62 $Y=1.575
+ $X2=0 $Y2=0
cc_656 N_A_211_363#_c_843_n N_A_1179_183#_c_1046_n 0.00386411f $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_657 N_A_211_363#_c_846_n N_A_1179_183#_c_1046_n 0.0180796f $X=5.51 $Y=0.87
+ $X2=0 $Y2=0
cc_658 N_A_211_363#_c_840_n N_A_1001_47#_M1009_d 0.00163744f $X=5.085 $Y=0.51
+ $X2=-0.19 $Y2=-0.24
cc_659 N_A_211_363#_c_842_n N_A_1001_47#_M1009_d 3.07407e-19 $X=5.155 $Y=0.735
+ $X2=-0.19 $Y2=-0.24
cc_660 N_A_211_363#_c_836_n N_A_1001_47#_c_1141_n 0.00960751f $X=7.335 $Y=0.705
+ $X2=0 $Y2=0
cc_661 N_A_211_363#_c_839_n N_A_1001_47#_c_1141_n 0.0010974f $X=7.525 $Y=0.87
+ $X2=0 $Y2=0
cc_662 N_A_211_363#_c_838_n N_A_1001_47#_c_1142_n 3.2664e-19 $X=7.62 $Y=1.575
+ $X2=0 $Y2=0
cc_663 N_A_211_363#_c_847_n N_A_1001_47#_c_1142_n 0.00960751f $X=7.48 $Y=0.87
+ $X2=0 $Y2=0
cc_664 N_A_211_363#_c_848_n N_A_1001_47#_c_1162_n 0.00432343f $X=4.95 $Y=1.99
+ $X2=0 $Y2=0
cc_665 N_A_211_363#_c_837_n N_A_1001_47#_c_1162_n 0.00454699f $X=4.94 $Y=1.74
+ $X2=0 $Y2=0
cc_666 N_A_211_363#_c_835_n N_A_1001_47#_c_1167_n 0.00854005f $X=5.51 $Y=0.705
+ $X2=0 $Y2=0
cc_667 N_A_211_363#_c_840_n N_A_1001_47#_c_1167_n 0.007819f $X=5.085 $Y=0.51
+ $X2=0 $Y2=0
cc_668 N_A_211_363#_c_843_n N_A_1001_47#_c_1167_n 0.00608741f $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_669 N_A_211_363#_c_957_p N_A_1001_47#_c_1167_n 6.15789e-19 $X=5.375 $Y=0.85
+ $X2=0 $Y2=0
cc_670 N_A_211_363#_c_845_n N_A_1001_47#_c_1167_n 0.0249559f $X=5.23 $Y=0.85
+ $X2=0 $Y2=0
cc_671 N_A_211_363#_c_846_n N_A_1001_47#_c_1167_n 0.00368644f $X=5.51 $Y=0.87
+ $X2=0 $Y2=0
cc_672 N_A_211_363#_c_835_n N_A_1001_47#_c_1145_n 0.00628549f $X=5.51 $Y=0.705
+ $X2=0 $Y2=0
cc_673 N_A_211_363#_c_837_n N_A_1001_47#_c_1145_n 0.00929804f $X=4.94 $Y=1.74
+ $X2=0 $Y2=0
cc_674 N_A_211_363#_c_840_n N_A_1001_47#_c_1145_n 0.00600133f $X=5.085 $Y=0.51
+ $X2=0 $Y2=0
cc_675 N_A_211_363#_c_843_n N_A_1001_47#_c_1145_n 0.0194801f $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_676 N_A_211_363#_c_957_p N_A_1001_47#_c_1145_n 5.14709e-19 $X=5.375 $Y=0.85
+ $X2=0 $Y2=0
cc_677 N_A_211_363#_c_845_n N_A_1001_47#_c_1145_n 0.0189145f $X=5.23 $Y=0.85
+ $X2=0 $Y2=0
cc_678 N_A_211_363#_c_837_n N_A_1001_47#_c_1146_n 0.00612128f $X=4.94 $Y=1.74
+ $X2=0 $Y2=0
cc_679 N_A_211_363#_c_843_n N_A_1001_47#_c_1146_n 0.00977661f $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_680 N_A_211_363#_c_849_n N_A_1653_315#_c_1266_n 0.0285138f $X=7.7 $Y=1.99
+ $X2=0 $Y2=0
cc_681 N_A_211_363#_c_852_n N_A_1653_315#_c_1266_n 4.80585e-19 $X=7.76 $Y=1.74
+ $X2=0 $Y2=0
cc_682 N_A_211_363#_c_849_n N_A_1464_413#_c_1384_n 0.0143918f $X=7.7 $Y=1.99
+ $X2=0 $Y2=0
cc_683 N_A_211_363#_c_852_n N_A_1464_413#_c_1384_n 0.0153945f $X=7.76 $Y=1.74
+ $X2=0 $Y2=0
cc_684 N_A_211_363#_c_836_n N_A_1464_413#_c_1388_n 0.00196231f $X=7.335 $Y=0.705
+ $X2=0 $Y2=0
cc_685 N_A_211_363#_c_839_n N_A_1464_413#_c_1388_n 0.0153898f $X=7.525 $Y=0.87
+ $X2=0 $Y2=0
cc_686 N_A_211_363#_c_847_n N_A_1464_413#_c_1388_n 8.58658e-19 $X=7.48 $Y=0.87
+ $X2=0 $Y2=0
cc_687 N_A_211_363#_c_849_n N_A_1464_413#_c_1381_n 0.00703212f $X=7.7 $Y=1.99
+ $X2=0 $Y2=0
cc_688 N_A_211_363#_c_838_n N_A_1464_413#_c_1381_n 0.00712801f $X=7.62 $Y=1.575
+ $X2=0 $Y2=0
cc_689 N_A_211_363#_c_852_n N_A_1464_413#_c_1381_n 0.020822f $X=7.76 $Y=1.74
+ $X2=0 $Y2=0
cc_690 N_A_211_363#_c_849_n N_A_1464_413#_c_1376_n 0.00102186f $X=7.7 $Y=1.99
+ $X2=0 $Y2=0
cc_691 N_A_211_363#_c_838_n N_A_1464_413#_c_1376_n 0.0226171f $X=7.62 $Y=1.575
+ $X2=0 $Y2=0
cc_692 N_A_211_363#_c_836_n N_A_1464_413#_c_1377_n 8.84292e-19 $X=7.335 $Y=0.705
+ $X2=0 $Y2=0
cc_693 N_A_211_363#_c_839_n N_A_1464_413#_c_1377_n 0.0213581f $X=7.525 $Y=0.87
+ $X2=0 $Y2=0
cc_694 N_A_211_363#_c_901_n N_A_1464_413#_c_1377_n 8.51213e-19 $X=7.27 $Y=0.85
+ $X2=0 $Y2=0
cc_695 N_A_211_363#_c_847_n N_A_1464_413#_c_1377_n 3.55894e-19 $X=7.48 $Y=0.87
+ $X2=0 $Y2=0
cc_696 N_A_211_363#_c_844_n N_VPWR_c_1518_n 0.0202126f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_697 N_A_211_363#_c_848_n N_VPWR_c_1520_n 0.00269426f $X=4.95 $Y=1.99 $X2=0
+ $Y2=0
cc_698 N_A_211_363#_c_848_n N_VPWR_c_1531_n 0.00659238f $X=4.95 $Y=1.99 $X2=0
+ $Y2=0
cc_699 N_A_211_363#_c_849_n N_VPWR_c_1533_n 0.00460277f $X=7.7 $Y=1.99 $X2=0
+ $Y2=0
cc_700 N_A_211_363#_c_844_n N_VPWR_c_1536_n 0.0120448f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_701 N_A_211_363#_c_848_n N_VPWR_c_1517_n 0.00850916f $X=4.95 $Y=1.99 $X2=0
+ $Y2=0
cc_702 N_A_211_363#_c_849_n N_VPWR_c_1517_n 0.006692f $X=7.7 $Y=1.99 $X2=0 $Y2=0
cc_703 N_A_211_363#_c_837_n N_VPWR_c_1517_n 0.00196481f $X=4.94 $Y=1.74 $X2=0
+ $Y2=0
cc_704 N_A_211_363#_c_844_n N_VPWR_c_1517_n 0.00308197f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_705 N_A_211_363#_c_840_n N_A_604_369#_M1014_d 0.00275032f $X=5.085 $Y=0.51
+ $X2=-0.19 $Y2=-0.24
cc_706 N_A_211_363#_c_840_n N_A_604_369#_M1009_s 0.00646594f $X=5.085 $Y=0.51
+ $X2=0 $Y2=0
cc_707 N_A_211_363#_c_840_n N_A_604_369#_c_1740_n 0.0162091f $X=5.085 $Y=0.51
+ $X2=0 $Y2=0
cc_708 N_A_211_363#_c_840_n N_A_604_369#_c_1716_n 0.0147466f $X=5.085 $Y=0.51
+ $X2=0 $Y2=0
cc_709 N_A_211_363#_c_840_n N_A_604_369#_c_1717_n 0.0192039f $X=5.085 $Y=0.51
+ $X2=0 $Y2=0
cc_710 N_A_211_363#_c_840_n N_A_604_369#_c_1719_n 0.0121812f $X=5.085 $Y=0.51
+ $X2=0 $Y2=0
cc_711 N_A_211_363#_c_842_n N_A_604_369#_c_1719_n 0.00459717f $X=5.155 $Y=0.735
+ $X2=0 $Y2=0
cc_712 N_A_211_363#_c_845_n N_A_604_369#_c_1719_n 6.47147e-19 $X=5.23 $Y=0.85
+ $X2=0 $Y2=0
cc_713 N_A_211_363#_c_848_n N_A_604_369#_c_1720_n 0.00543259f $X=4.95 $Y=1.99
+ $X2=0 $Y2=0
cc_714 N_A_211_363#_c_837_n N_A_604_369#_c_1720_n 0.0594075f $X=4.94 $Y=1.74
+ $X2=0 $Y2=0
cc_715 N_A_211_363#_c_957_p N_A_604_369#_c_1720_n 3.52067e-19 $X=5.375 $Y=0.85
+ $X2=0 $Y2=0
cc_716 N_A_211_363#_c_845_n N_A_604_369#_c_1720_n 0.0115017f $X=5.23 $Y=0.85
+ $X2=0 $Y2=0
cc_717 N_A_211_363#_c_840_n N_A_604_369#_c_1721_n 0.0120713f $X=5.085 $Y=0.51
+ $X2=0 $Y2=0
cc_718 N_A_211_363#_c_845_n N_A_604_369#_c_1721_n 6.25683e-19 $X=5.23 $Y=0.85
+ $X2=0 $Y2=0
cc_719 N_A_211_363#_c_842_n N_A_604_369#_c_1722_n 8.48865e-19 $X=5.155 $Y=0.735
+ $X2=0 $Y2=0
cc_720 N_A_211_363#_c_845_n N_A_604_369#_c_1722_n 0.0142932f $X=5.23 $Y=0.85
+ $X2=0 $Y2=0
cc_721 N_A_211_363#_c_848_n N_A_604_369#_c_1726_n 0.0122886f $X=4.95 $Y=1.99
+ $X2=0 $Y2=0
cc_722 N_A_211_363#_c_837_n N_A_604_369#_c_1726_n 0.00558961f $X=4.94 $Y=1.74
+ $X2=0 $Y2=0
cc_723 N_A_211_363#_c_840_n N_VGND_M1021_d 0.00386578f $X=5.085 $Y=0.51 $X2=0
+ $Y2=0
cc_724 N_A_211_363#_c_840_n N_VGND_M1037_d 0.00349104f $X=5.085 $Y=0.51 $X2=0
+ $Y2=0
cc_725 N_A_211_363#_c_840_n N_VGND_c_1880_n 0.00746988f $X=5.085 $Y=0.51 $X2=0
+ $Y2=0
cc_726 N_A_211_363#_c_840_n N_VGND_c_1881_n 0.00839237f $X=5.085 $Y=0.51 $X2=0
+ $Y2=0
cc_727 N_A_211_363#_c_843_n N_VGND_c_1882_n 0.00197288f $X=7.125 $Y=0.85 $X2=0
+ $Y2=0
cc_728 N_A_211_363#_c_840_n N_VGND_c_1890_n 0.00187533f $X=5.085 $Y=0.51 $X2=0
+ $Y2=0
cc_729 N_A_211_363#_c_841_n N_VGND_c_1890_n 0.00104058f $X=1.345 $Y=0.51 $X2=0
+ $Y2=0
cc_730 N_A_211_363#_c_844_n N_VGND_c_1890_n 0.00732874f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_731 N_A_211_363#_c_840_n N_VGND_c_1892_n 0.00298108f $X=5.085 $Y=0.51 $X2=0
+ $Y2=0
cc_732 N_A_211_363#_c_835_n N_VGND_c_1895_n 0.0037981f $X=5.51 $Y=0.705 $X2=0
+ $Y2=0
cc_733 N_A_211_363#_c_840_n N_VGND_c_1895_n 0.00181568f $X=5.085 $Y=0.51 $X2=0
+ $Y2=0
cc_734 N_A_211_363#_c_845_n N_VGND_c_1895_n 0.00291348f $X=5.23 $Y=0.85 $X2=0
+ $Y2=0
cc_735 N_A_211_363#_c_836_n N_VGND_c_1896_n 0.00435108f $X=7.335 $Y=0.705 $X2=0
+ $Y2=0
cc_736 N_A_211_363#_c_839_n N_VGND_c_1896_n 0.00414043f $X=7.525 $Y=0.87 $X2=0
+ $Y2=0
cc_737 N_A_211_363#_c_847_n N_VGND_c_1896_n 0.00152809f $X=7.48 $Y=0.87 $X2=0
+ $Y2=0
cc_738 N_A_211_363#_c_841_n N_VGND_c_1900_n 0.0021356f $X=1.345 $Y=0.51 $X2=0
+ $Y2=0
cc_739 N_A_211_363#_M1001_d N_VGND_c_1906_n 0.00151052f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_740 N_A_211_363#_c_835_n N_VGND_c_1906_n 0.00584986f $X=5.51 $Y=0.705 $X2=0
+ $Y2=0
cc_741 N_A_211_363#_c_836_n N_VGND_c_1906_n 0.0063925f $X=7.335 $Y=0.705 $X2=0
+ $Y2=0
cc_742 N_A_211_363#_c_839_n N_VGND_c_1906_n 0.00468679f $X=7.525 $Y=0.87 $X2=0
+ $Y2=0
cc_743 N_A_211_363#_c_840_n N_VGND_c_1906_n 0.332687f $X=5.085 $Y=0.51 $X2=0
+ $Y2=0
cc_744 N_A_211_363#_c_841_n N_VGND_c_1906_n 0.0338686f $X=1.345 $Y=0.51 $X2=0
+ $Y2=0
cc_745 N_A_211_363#_c_843_n N_VGND_c_1906_n 0.0810653f $X=7.125 $Y=0.85 $X2=0
+ $Y2=0
cc_746 N_A_211_363#_c_957_p N_VGND_c_1906_n 0.00755712f $X=5.375 $Y=0.85 $X2=0
+ $Y2=0
cc_747 N_A_211_363#_c_844_n N_VGND_c_1906_n 0.00169577f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_748 N_A_211_363#_c_901_n N_VGND_c_1906_n 0.0145657f $X=7.27 $Y=0.85 $X2=0
+ $Y2=0
cc_749 N_A_211_363#_c_847_n N_VGND_c_1906_n 0.00251234f $X=7.48 $Y=0.87 $X2=0
+ $Y2=0
cc_750 N_A_211_363#_c_840_n A_529_47# 0.0033455f $X=5.085 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_751 N_A_211_363#_c_840_n A_717_47# 0.00460223f $X=5.085 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_752 N_A_1179_183#_c_1045_n N_A_1001_47#_c_1140_n 0.00685148f $X=6.875
+ $Y=2.135 $X2=0 $Y2=0
cc_753 N_A_1179_183#_c_1040_n N_A_1001_47#_c_1147_n 0.00419555f $X=5.995 $Y=1.89
+ $X2=0 $Y2=0
cc_754 N_A_1179_183#_c_1048_n N_A_1001_47#_c_1147_n 0.00719967f $X=5.995 $Y=1.99
+ $X2=0 $Y2=0
cc_755 N_A_1179_183#_c_1059_n N_A_1001_47#_c_1147_n 0.00529276f $X=6.94 $Y=2.3
+ $X2=0 $Y2=0
cc_756 N_A_1179_183#_c_1045_n N_A_1001_47#_c_1147_n 0.0113977f $X=6.875 $Y=2.135
+ $X2=0 $Y2=0
cc_757 N_A_1179_183#_M1017_g N_A_1001_47#_c_1141_n 0.00774331f $X=6 $Y=0.445
+ $X2=0 $Y2=0
cc_758 N_A_1179_183#_c_1072_n N_A_1001_47#_c_1141_n 0.00627039f $X=6.835
+ $Y=0.765 $X2=0 $Y2=0
cc_759 N_A_1179_183#_c_1092_p N_A_1001_47#_c_1141_n 0.00614274f $X=6.945 $Y=0.45
+ $X2=0 $Y2=0
cc_760 N_A_1179_183#_c_1044_n N_A_1001_47#_c_1141_n 0.00666077f $X=6.835
+ $Y=0.915 $X2=0 $Y2=0
cc_761 N_A_1179_183#_c_1046_n N_A_1001_47#_c_1141_n 0.00413835f $X=6 $Y=0.93
+ $X2=0 $Y2=0
cc_762 N_A_1179_183#_c_1040_n N_A_1001_47#_c_1142_n 0.00485524f $X=5.995 $Y=1.89
+ $X2=0 $Y2=0
cc_763 N_A_1179_183#_c_1042_n N_A_1001_47#_c_1142_n 0.0102886f $X=6.725 $Y=0.915
+ $X2=0 $Y2=0
cc_764 N_A_1179_183#_c_1043_n N_A_1001_47#_c_1142_n 2.52267e-19 $X=6.265 $Y=0.93
+ $X2=0 $Y2=0
cc_765 N_A_1179_183#_c_1044_n N_A_1001_47#_c_1142_n 0.00358011f $X=6.835
+ $Y=0.915 $X2=0 $Y2=0
cc_766 N_A_1179_183#_c_1045_n N_A_1001_47#_c_1142_n 0.00411223f $X=6.875
+ $Y=2.135 $X2=0 $Y2=0
cc_767 N_A_1179_183#_c_1046_n N_A_1001_47#_c_1142_n 0.00574663f $X=6 $Y=0.93
+ $X2=0 $Y2=0
cc_768 N_A_1179_183#_c_1040_n N_A_1001_47#_c_1143_n 0.017484f $X=5.995 $Y=1.89
+ $X2=0 $Y2=0
cc_769 N_A_1179_183#_c_1042_n N_A_1001_47#_c_1143_n 0.00400764f $X=6.725
+ $Y=0.915 $X2=0 $Y2=0
cc_770 N_A_1179_183#_c_1046_n N_A_1001_47#_c_1143_n 0.00238133f $X=6 $Y=0.93
+ $X2=0 $Y2=0
cc_771 N_A_1179_183#_c_1040_n N_A_1001_47#_c_1144_n 0.00203945f $X=5.995 $Y=1.89
+ $X2=0 $Y2=0
cc_772 N_A_1179_183#_c_1045_n N_A_1001_47#_c_1144_n 0.011008f $X=6.875 $Y=2.135
+ $X2=0 $Y2=0
cc_773 N_A_1179_183#_c_1048_n N_A_1001_47#_c_1162_n 0.0109992f $X=5.995 $Y=1.99
+ $X2=0 $Y2=0
cc_774 N_A_1179_183#_M1017_g N_A_1001_47#_c_1145_n 0.00451615f $X=6 $Y=0.445
+ $X2=0 $Y2=0
cc_775 N_A_1179_183#_c_1043_n N_A_1001_47#_c_1145_n 0.0195837f $X=6.265 $Y=0.93
+ $X2=0 $Y2=0
cc_776 N_A_1179_183#_c_1046_n N_A_1001_47#_c_1145_n 0.010005f $X=6 $Y=0.93 $X2=0
+ $Y2=0
cc_777 N_A_1179_183#_c_1040_n N_A_1001_47#_c_1150_n 0.00884796f $X=5.995 $Y=1.89
+ $X2=0 $Y2=0
cc_778 N_A_1179_183#_c_1048_n N_A_1001_47#_c_1150_n 0.00967444f $X=5.995 $Y=1.99
+ $X2=0 $Y2=0
cc_779 N_A_1179_183#_c_1045_n N_A_1001_47#_c_1150_n 0.00780656f $X=6.875
+ $Y=2.135 $X2=0 $Y2=0
cc_780 N_A_1179_183#_c_1040_n N_A_1001_47#_c_1146_n 0.0162689f $X=5.995 $Y=1.89
+ $X2=0 $Y2=0
cc_781 N_A_1179_183#_c_1042_n N_A_1001_47#_c_1146_n 0.0186614f $X=6.725 $Y=0.915
+ $X2=0 $Y2=0
cc_782 N_A_1179_183#_c_1043_n N_A_1001_47#_c_1146_n 0.0112018f $X=6.265 $Y=0.93
+ $X2=0 $Y2=0
cc_783 N_A_1179_183#_c_1045_n N_A_1001_47#_c_1146_n 0.0251292f $X=6.875 $Y=2.135
+ $X2=0 $Y2=0
cc_784 N_A_1179_183#_c_1046_n N_A_1001_47#_c_1146_n 0.0021403f $X=6 $Y=0.93
+ $X2=0 $Y2=0
cc_785 N_A_1179_183#_c_1059_n N_A_1464_413#_c_1384_n 0.0110665f $X=6.94 $Y=2.3
+ $X2=0 $Y2=0
cc_786 N_A_1179_183#_c_1040_n N_VPWR_c_1521_n 3.85242e-19 $X=5.995 $Y=1.89 $X2=0
+ $Y2=0
cc_787 N_A_1179_183#_c_1048_n N_VPWR_c_1521_n 0.00532796f $X=5.995 $Y=1.99 $X2=0
+ $Y2=0
cc_788 N_A_1179_183#_c_1045_n N_VPWR_c_1521_n 0.0450469f $X=6.875 $Y=2.135 $X2=0
+ $Y2=0
cc_789 N_A_1179_183#_c_1048_n N_VPWR_c_1531_n 0.00457093f $X=5.995 $Y=1.99 $X2=0
+ $Y2=0
cc_790 N_A_1179_183#_c_1059_n N_VPWR_c_1533_n 0.0185094f $X=6.94 $Y=2.3 $X2=0
+ $Y2=0
cc_791 N_A_1179_183#_M1025_d N_VPWR_c_1517_n 0.0030383f $X=6.795 $Y=1.735 $X2=0
+ $Y2=0
cc_792 N_A_1179_183#_c_1048_n N_VPWR_c_1517_n 0.00678138f $X=5.995 $Y=1.99 $X2=0
+ $Y2=0
cc_793 N_A_1179_183#_c_1059_n N_VPWR_c_1517_n 0.00522915f $X=6.94 $Y=2.3 $X2=0
+ $Y2=0
cc_794 N_A_1179_183#_c_1042_n N_VGND_M1017_d 0.00408144f $X=6.725 $Y=0.915 $X2=0
+ $Y2=0
cc_795 N_A_1179_183#_M1017_g N_VGND_c_1882_n 0.00984181f $X=6 $Y=0.445 $X2=0
+ $Y2=0
cc_796 N_A_1179_183#_c_1043_n N_VGND_c_1882_n 0.0260635f $X=6.265 $Y=0.93 $X2=0
+ $Y2=0
cc_797 N_A_1179_183#_c_1046_n N_VGND_c_1882_n 0.00123827f $X=6 $Y=0.93 $X2=0
+ $Y2=0
cc_798 N_A_1179_183#_M1017_g N_VGND_c_1895_n 0.00585385f $X=6 $Y=0.445 $X2=0
+ $Y2=0
cc_799 N_A_1179_183#_c_1092_p N_VGND_c_1896_n 0.00738334f $X=6.945 $Y=0.45 $X2=0
+ $Y2=0
cc_800 N_A_1179_183#_c_1073_n N_VGND_c_1896_n 0.0100275f $X=7.07 $Y=0.45 $X2=0
+ $Y2=0
cc_801 N_A_1179_183#_M1002_d N_VGND_c_1906_n 0.00247799f $X=6.905 $Y=0.235 $X2=0
+ $Y2=0
cc_802 N_A_1179_183#_M1017_g N_VGND_c_1906_n 0.00740521f $X=6 $Y=0.445 $X2=0
+ $Y2=0
cc_803 N_A_1179_183#_c_1042_n N_VGND_c_1906_n 0.00430476f $X=6.725 $Y=0.915
+ $X2=0 $Y2=0
cc_804 N_A_1179_183#_c_1092_p N_VGND_c_1906_n 0.00343551f $X=6.945 $Y=0.45 $X2=0
+ $Y2=0
cc_805 N_A_1179_183#_c_1073_n N_VGND_c_1906_n 0.00445429f $X=7.07 $Y=0.45 $X2=0
+ $Y2=0
cc_806 N_A_1179_183#_c_1043_n N_VGND_c_1906_n 0.00284313f $X=6.265 $Y=0.93 $X2=0
+ $Y2=0
cc_807 N_A_1001_47#_c_1162_n N_VPWR_M1000_d 0.00249014f $X=5.995 $Y=2.275 $X2=0
+ $Y2=0
cc_808 N_A_1001_47#_c_1150_n N_VPWR_M1000_d 0.00416039f $X=6.105 $Y=2.19 $X2=0
+ $Y2=0
cc_809 N_A_1001_47#_c_1147_n N_VPWR_c_1521_n 0.00502749f $X=6.705 $Y=1.66 $X2=0
+ $Y2=0
cc_810 N_A_1001_47#_c_1143_n N_VPWR_c_1521_n 9.59975e-19 $X=6.605 $Y=1.41 $X2=0
+ $Y2=0
cc_811 N_A_1001_47#_c_1162_n N_VPWR_c_1521_n 0.0138309f $X=5.995 $Y=2.275 $X2=0
+ $Y2=0
cc_812 N_A_1001_47#_c_1150_n N_VPWR_c_1521_n 0.0256293f $X=6.105 $Y=2.19 $X2=0
+ $Y2=0
cc_813 N_A_1001_47#_c_1146_n N_VPWR_c_1521_n 0.00748119f $X=6.105 $Y=1.41 $X2=0
+ $Y2=0
cc_814 N_A_1001_47#_c_1162_n N_VPWR_c_1531_n 0.0416565f $X=5.995 $Y=2.275 $X2=0
+ $Y2=0
cc_815 N_A_1001_47#_c_1147_n N_VPWR_c_1533_n 0.00597712f $X=6.705 $Y=1.66 $X2=0
+ $Y2=0
cc_816 N_A_1001_47#_M1028_d N_VPWR_c_1517_n 0.00230779f $X=5.04 $Y=2.065 $X2=0
+ $Y2=0
cc_817 N_A_1001_47#_c_1147_n N_VPWR_c_1517_n 0.00740372f $X=6.705 $Y=1.66 $X2=0
+ $Y2=0
cc_818 N_A_1001_47#_c_1162_n N_VPWR_c_1517_n 0.0183713f $X=5.995 $Y=2.275 $X2=0
+ $Y2=0
cc_819 N_A_1001_47#_c_1167_n N_A_604_369#_c_1721_n 0.00994528f $X=5.705 $Y=0.45
+ $X2=0 $Y2=0
cc_820 N_A_1001_47#_c_1162_n N_A_604_369#_c_1726_n 0.0123679f $X=5.995 $Y=2.275
+ $X2=0 $Y2=0
cc_821 N_A_1001_47#_c_1162_n A_1111_413# 0.0050022f $X=5.995 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_822 N_A_1001_47#_c_1141_n N_VGND_c_1882_n 0.00681995f $X=6.755 $Y=0.95 $X2=0
+ $Y2=0
cc_823 N_A_1001_47#_c_1167_n N_VGND_c_1895_n 0.027869f $X=5.705 $Y=0.45 $X2=0
+ $Y2=0
cc_824 N_A_1001_47#_c_1141_n N_VGND_c_1896_n 0.0037962f $X=6.755 $Y=0.95 $X2=0
+ $Y2=0
cc_825 N_A_1001_47#_M1009_d N_VGND_c_1906_n 0.00259162f $X=5.005 $Y=0.235 $X2=0
+ $Y2=0
cc_826 N_A_1001_47#_c_1141_n N_VGND_c_1906_n 0.006268f $X=6.755 $Y=0.95 $X2=0
+ $Y2=0
cc_827 N_A_1001_47#_c_1167_n N_VGND_c_1906_n 0.0113167f $X=5.705 $Y=0.45 $X2=0
+ $Y2=0
cc_828 N_A_1001_47#_c_1167_n A_1117_47# 0.00455507f $X=5.705 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_829 N_A_1001_47#_c_1145_n A_1117_47# 0.00131375f $X=5.79 $Y=1.315 $X2=-0.19
+ $Y2=-0.24
cc_830 N_A_1653_315#_c_1268_n N_A_1464_413#_c_1378_n 0.0299413f $X=10.06 $Y=1.41
+ $X2=0 $Y2=0
cc_831 N_A_1653_315#_c_1276_n N_A_1464_413#_c_1378_n 0.00603579f $X=9.235
+ $Y=2.34 $X2=0 $Y2=0
cc_832 N_A_1653_315#_c_1277_n N_A_1464_413#_c_1378_n 0.00443259f $X=9.307
+ $Y=1.575 $X2=0 $Y2=0
cc_833 N_A_1653_315#_c_1279_n N_A_1464_413#_c_1378_n 0.00411833f $X=9.235
+ $Y=1.66 $X2=0 $Y2=0
cc_834 N_A_1653_315#_c_1257_n N_A_1464_413#_c_1372_n 0.0158017f $X=10.085
+ $Y=0.995 $X2=0 $Y2=0
cc_835 N_A_1653_315#_c_1263_n N_A_1464_413#_c_1372_n 0.0044201f $X=9.307
+ $Y=0.995 $X2=0 $Y2=0
cc_836 N_A_1653_315#_M1024_g N_A_1464_413#_c_1373_n 0.017717f $X=8.505 $Y=0.445
+ $X2=0 $Y2=0
cc_837 N_A_1653_315#_c_1275_n N_A_1464_413#_c_1373_n 0.00567751f $X=9.07 $Y=1.74
+ $X2=0 $Y2=0
cc_838 N_A_1653_315#_c_1265_n N_A_1464_413#_c_1373_n 0.00747686f $X=9.235
+ $Y=0.385 $X2=0 $Y2=0
cc_839 N_A_1653_315#_c_1279_n N_A_1464_413#_c_1373_n 0.00591375f $X=9.235
+ $Y=1.66 $X2=0 $Y2=0
cc_840 N_A_1653_315#_c_1293_p N_A_1464_413#_c_1373_n 0.0168182f $X=9.307 $Y=1.16
+ $X2=0 $Y2=0
cc_841 N_A_1653_315#_c_1260_n N_A_1464_413#_c_1374_n 0.0241585f $X=10.63 $Y=1.16
+ $X2=0 $Y2=0
cc_842 N_A_1653_315#_c_1277_n N_A_1464_413#_c_1374_n 0.0034091f $X=9.307
+ $Y=1.575 $X2=0 $Y2=0
cc_843 N_A_1653_315#_c_1264_n N_A_1464_413#_c_1374_n 0.0241415f $X=9.915 $Y=1.16
+ $X2=0 $Y2=0
cc_844 N_A_1653_315#_c_1293_p N_A_1464_413#_c_1374_n 0.00162165f $X=9.307
+ $Y=1.16 $X2=0 $Y2=0
cc_845 N_A_1653_315#_c_1266_n N_A_1464_413#_c_1384_n 0.00511661f $X=8.365
+ $Y=1.99 $X2=0 $Y2=0
cc_846 N_A_1653_315#_M1024_g N_A_1464_413#_c_1388_n 6.7345e-19 $X=8.505 $Y=0.445
+ $X2=0 $Y2=0
cc_847 N_A_1653_315#_c_1266_n N_A_1464_413#_c_1381_n 0.0214064f $X=8.365 $Y=1.99
+ $X2=0 $Y2=0
cc_848 N_A_1653_315#_c_1275_n N_A_1464_413#_c_1381_n 0.0219216f $X=9.07 $Y=1.74
+ $X2=0 $Y2=0
cc_849 N_A_1653_315#_c_1266_n N_A_1464_413#_c_1375_n 0.00861313f $X=8.365
+ $Y=1.99 $X2=0 $Y2=0
cc_850 N_A_1653_315#_M1024_g N_A_1464_413#_c_1375_n 0.0184544f $X=8.505 $Y=0.445
+ $X2=0 $Y2=0
cc_851 N_A_1653_315#_c_1275_n N_A_1464_413#_c_1375_n 0.033362f $X=9.07 $Y=1.74
+ $X2=0 $Y2=0
cc_852 N_A_1653_315#_c_1265_n N_A_1464_413#_c_1375_n 7.42989e-19 $X=9.235
+ $Y=0.385 $X2=0 $Y2=0
cc_853 N_A_1653_315#_c_1293_p N_A_1464_413#_c_1375_n 0.0277655f $X=9.307 $Y=1.16
+ $X2=0 $Y2=0
cc_854 N_A_1653_315#_M1024_g N_A_1464_413#_c_1376_n 0.00857838f $X=8.505
+ $Y=0.445 $X2=0 $Y2=0
cc_855 N_A_1653_315#_M1024_g N_A_1464_413#_c_1377_n 0.00777602f $X=8.505
+ $Y=0.445 $X2=0 $Y2=0
cc_856 N_A_1653_315#_c_1272_n N_A_2234_47#_c_1461_n 0.00499537f $X=11.53 $Y=1.67
+ $X2=0 $Y2=0
cc_857 N_A_1653_315#_c_1273_n N_A_2234_47#_c_1461_n 0.00920897f $X=11.53 $Y=1.77
+ $X2=0 $Y2=0
cc_858 N_A_1653_315#_M1027_g N_A_2234_47#_c_1455_n 0.0110006f $X=11.555 $Y=0.445
+ $X2=0 $Y2=0
cc_859 N_A_1653_315#_c_1258_n N_A_2234_47#_c_1457_n 0.00514121f $X=10.555
+ $Y=0.995 $X2=0 $Y2=0
cc_860 N_A_1653_315#_M1027_g N_A_2234_47#_c_1457_n 0.0120696f $X=11.555 $Y=0.445
+ $X2=0 $Y2=0
cc_861 N_A_1653_315#_c_1269_n N_A_2234_47#_c_1463_n 0.00476119f $X=10.53 $Y=1.41
+ $X2=0 $Y2=0
cc_862 N_A_1653_315#_c_1260_n N_A_2234_47#_c_1463_n 0.00146603f $X=10.63 $Y=1.16
+ $X2=0 $Y2=0
cc_863 N_A_1653_315#_c_1272_n N_A_2234_47#_c_1463_n 0.0168274f $X=11.53 $Y=1.67
+ $X2=0 $Y2=0
cc_864 N_A_1653_315#_c_1273_n N_A_2234_47#_c_1463_n 0.0135486f $X=11.53 $Y=1.77
+ $X2=0 $Y2=0
cc_865 N_A_1653_315#_c_1262_n N_A_2234_47#_c_1458_n 0.0271722f $X=11.53 $Y=1.16
+ $X2=0 $Y2=0
cc_866 N_A_1653_315#_c_1259_n N_A_2234_47#_c_1459_n 0.0346091f $X=11.43 $Y=1.16
+ $X2=0 $Y2=0
cc_867 N_A_1653_315#_c_1262_n N_A_2234_47#_c_1459_n 0.00248969f $X=11.53 $Y=1.16
+ $X2=0 $Y2=0
cc_868 N_A_1653_315#_c_1272_n N_A_2234_47#_c_1460_n 0.00210665f $X=11.53 $Y=1.67
+ $X2=0 $Y2=0
cc_869 N_A_1653_315#_c_1262_n N_A_2234_47#_c_1460_n 0.00671506f $X=11.53 $Y=1.16
+ $X2=0 $Y2=0
cc_870 N_A_1653_315#_c_1266_n N_VPWR_c_1522_n 0.0200676f $X=8.365 $Y=1.99 $X2=0
+ $Y2=0
cc_871 N_A_1653_315#_c_1275_n N_VPWR_c_1522_n 0.0192158f $X=9.07 $Y=1.74 $X2=0
+ $Y2=0
cc_872 N_A_1653_315#_c_1276_n N_VPWR_c_1522_n 0.0197296f $X=9.235 $Y=2.34 $X2=0
+ $Y2=0
cc_873 N_A_1653_315#_c_1268_n N_VPWR_c_1523_n 0.0282178f $X=10.06 $Y=1.41 $X2=0
+ $Y2=0
cc_874 N_A_1653_315#_c_1269_n N_VPWR_c_1523_n 0.00103735f $X=10.53 $Y=1.41 $X2=0
+ $Y2=0
cc_875 N_A_1653_315#_c_1260_n N_VPWR_c_1523_n 0.00370295f $X=10.63 $Y=1.16 $X2=0
+ $Y2=0
cc_876 N_A_1653_315#_c_1264_n N_VPWR_c_1523_n 0.0201149f $X=9.915 $Y=1.16 $X2=0
+ $Y2=0
cc_877 N_A_1653_315#_c_1269_n N_VPWR_c_1524_n 0.0107752f $X=10.53 $Y=1.41 $X2=0
+ $Y2=0
cc_878 N_A_1653_315#_c_1259_n N_VPWR_c_1524_n 0.00666742f $X=11.43 $Y=1.16 $X2=0
+ $Y2=0
cc_879 N_A_1653_315#_c_1272_n N_VPWR_c_1524_n 5.68274e-19 $X=11.53 $Y=1.67 $X2=0
+ $Y2=0
cc_880 N_A_1653_315#_c_1273_n N_VPWR_c_1524_n 0.00358544f $X=11.53 $Y=1.77 $X2=0
+ $Y2=0
cc_881 N_A_1653_315#_c_1273_n N_VPWR_c_1525_n 0.00674661f $X=11.53 $Y=1.77 $X2=0
+ $Y2=0
cc_882 N_A_1653_315#_c_1272_n N_VPWR_c_1526_n 0.00374694f $X=11.53 $Y=1.67 $X2=0
+ $Y2=0
cc_883 N_A_1653_315#_c_1273_n N_VPWR_c_1526_n 0.0141193f $X=11.53 $Y=1.77 $X2=0
+ $Y2=0
cc_884 N_A_1653_315#_c_1266_n N_VPWR_c_1533_n 0.00712364f $X=8.365 $Y=1.99 $X2=0
+ $Y2=0
cc_885 N_A_1653_315#_c_1276_n N_VPWR_c_1537_n 0.0197996f $X=9.235 $Y=2.34 $X2=0
+ $Y2=0
cc_886 N_A_1653_315#_c_1268_n N_VPWR_c_1538_n 0.00622633f $X=10.06 $Y=1.41 $X2=0
+ $Y2=0
cc_887 N_A_1653_315#_c_1269_n N_VPWR_c_1538_n 0.00628756f $X=10.53 $Y=1.41 $X2=0
+ $Y2=0
cc_888 N_A_1653_315#_M1015_s N_VPWR_c_1517_n 0.00217852f $X=9.11 $Y=1.485 $X2=0
+ $Y2=0
cc_889 N_A_1653_315#_c_1266_n N_VPWR_c_1517_n 0.015655f $X=8.365 $Y=1.99 $X2=0
+ $Y2=0
cc_890 N_A_1653_315#_c_1268_n N_VPWR_c_1517_n 0.0104011f $X=10.06 $Y=1.41 $X2=0
+ $Y2=0
cc_891 N_A_1653_315#_c_1269_n N_VPWR_c_1517_n 0.0120424f $X=10.53 $Y=1.41 $X2=0
+ $Y2=0
cc_892 N_A_1653_315#_c_1273_n N_VPWR_c_1517_n 0.0139192f $X=11.53 $Y=1.77 $X2=0
+ $Y2=0
cc_893 N_A_1653_315#_c_1275_n N_VPWR_c_1517_n 0.0115245f $X=9.07 $Y=1.74 $X2=0
+ $Y2=0
cc_894 N_A_1653_315#_c_1276_n N_VPWR_c_1517_n 0.0124126f $X=9.235 $Y=2.34 $X2=0
+ $Y2=0
cc_895 N_A_1653_315#_c_1268_n N_Q_c_1844_n 0.00828013f $X=10.06 $Y=1.41 $X2=0
+ $Y2=0
cc_896 N_A_1653_315#_c_1257_n N_Q_c_1844_n 0.00293751f $X=10.085 $Y=0.995 $X2=0
+ $Y2=0
cc_897 N_A_1653_315#_c_1269_n N_Q_c_1844_n 0.0177553f $X=10.53 $Y=1.41 $X2=0
+ $Y2=0
cc_898 N_A_1653_315#_c_1258_n N_Q_c_1844_n 0.0119447f $X=10.555 $Y=0.995 $X2=0
+ $Y2=0
cc_899 N_A_1653_315#_c_1260_n N_Q_c_1844_n 0.037412f $X=10.63 $Y=1.16 $X2=0
+ $Y2=0
cc_900 N_A_1653_315#_c_1264_n N_Q_c_1844_n 0.0218309f $X=9.915 $Y=1.16 $X2=0
+ $Y2=0
cc_901 N_A_1653_315#_M1024_g N_VGND_c_1883_n 0.0192246f $X=8.505 $Y=0.445 $X2=0
+ $Y2=0
cc_902 N_A_1653_315#_c_1265_n N_VGND_c_1883_n 0.0209343f $X=9.235 $Y=0.385 $X2=0
+ $Y2=0
cc_903 N_A_1653_315#_c_1257_n N_VGND_c_1884_n 0.00643251f $X=10.085 $Y=0.995
+ $X2=0 $Y2=0
cc_904 N_A_1653_315#_c_1260_n N_VGND_c_1884_n 0.00444835f $X=10.63 $Y=1.16 $X2=0
+ $Y2=0
cc_905 N_A_1653_315#_c_1264_n N_VGND_c_1884_n 0.0204927f $X=9.915 $Y=1.16 $X2=0
+ $Y2=0
cc_906 N_A_1653_315#_c_1258_n N_VGND_c_1885_n 0.00628799f $X=10.555 $Y=0.995
+ $X2=0 $Y2=0
cc_907 N_A_1653_315#_c_1259_n N_VGND_c_1885_n 0.0072715f $X=11.43 $Y=1.16 $X2=0
+ $Y2=0
cc_908 N_A_1653_315#_M1027_g N_VGND_c_1885_n 0.0044645f $X=11.555 $Y=0.445 $X2=0
+ $Y2=0
cc_909 N_A_1653_315#_M1027_g N_VGND_c_1886_n 0.00585385f $X=11.555 $Y=0.445
+ $X2=0 $Y2=0
cc_910 N_A_1653_315#_M1027_g N_VGND_c_1887_n 0.00979412f $X=11.555 $Y=0.445
+ $X2=0 $Y2=0
cc_911 N_A_1653_315#_c_1265_n N_VGND_c_1897_n 0.0187449f $X=9.235 $Y=0.385 $X2=0
+ $Y2=0
cc_912 N_A_1653_315#_c_1257_n N_VGND_c_1898_n 0.00585385f $X=10.085 $Y=0.995
+ $X2=0 $Y2=0
cc_913 N_A_1653_315#_c_1258_n N_VGND_c_1898_n 0.00571722f $X=10.555 $Y=0.995
+ $X2=0 $Y2=0
cc_914 N_A_1653_315#_M1039_s N_VGND_c_1906_n 0.00322755f $X=9.11 $Y=0.235 $X2=0
+ $Y2=0
cc_915 N_A_1653_315#_c_1257_n N_VGND_c_1906_n 0.0110683f $X=10.085 $Y=0.995
+ $X2=0 $Y2=0
cc_916 N_A_1653_315#_c_1258_n N_VGND_c_1906_n 0.0118209f $X=10.555 $Y=0.995
+ $X2=0 $Y2=0
cc_917 N_A_1653_315#_M1027_g N_VGND_c_1906_n 0.0128045f $X=11.555 $Y=0.445 $X2=0
+ $Y2=0
cc_918 N_A_1653_315#_c_1265_n N_VGND_c_1906_n 0.0136152f $X=9.235 $Y=0.385 $X2=0
+ $Y2=0
cc_919 N_A_1464_413#_c_1378_n N_VPWR_c_1522_n 0.00222629f $X=9.47 $Y=1.41 $X2=0
+ $Y2=0
cc_920 N_A_1464_413#_c_1384_n N_VPWR_c_1522_n 0.0110234f $X=8.115 $Y=2.25 $X2=0
+ $Y2=0
cc_921 N_A_1464_413#_c_1381_n N_VPWR_c_1522_n 0.00172289f $X=8.2 $Y=2.165 $X2=0
+ $Y2=0
cc_922 N_A_1464_413#_c_1378_n N_VPWR_c_1523_n 0.00915264f $X=9.47 $Y=1.41 $X2=0
+ $Y2=0
cc_923 N_A_1464_413#_c_1384_n N_VPWR_c_1533_n 0.0324354f $X=8.115 $Y=2.25 $X2=0
+ $Y2=0
cc_924 N_A_1464_413#_c_1378_n N_VPWR_c_1537_n 0.00673882f $X=9.47 $Y=1.41 $X2=0
+ $Y2=0
cc_925 N_A_1464_413#_M1008_d N_VPWR_c_1517_n 0.00234902f $X=7.32 $Y=2.065 $X2=0
+ $Y2=0
cc_926 N_A_1464_413#_c_1378_n N_VPWR_c_1517_n 0.0133725f $X=9.47 $Y=1.41 $X2=0
+ $Y2=0
cc_927 N_A_1464_413#_c_1384_n N_VPWR_c_1517_n 0.0315385f $X=8.115 $Y=2.25 $X2=0
+ $Y2=0
cc_928 N_A_1464_413#_c_1384_n A_1558_413# 0.0125149f $X=8.115 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_929 N_A_1464_413#_c_1381_n A_1558_413# 0.00130185f $X=8.2 $Y=2.165 $X2=-0.19
+ $Y2=-0.24
cc_930 N_A_1464_413#_c_1372_n N_VGND_c_1883_n 0.00303997f $X=9.495 $Y=0.995
+ $X2=0 $Y2=0
cc_931 N_A_1464_413#_c_1375_n N_VGND_c_1883_n 0.0166909f $X=8.96 $Y=1.16 $X2=0
+ $Y2=0
cc_932 N_A_1464_413#_c_1372_n N_VGND_c_1884_n 0.00420747f $X=9.495 $Y=0.995
+ $X2=0 $Y2=0
cc_933 N_A_1464_413#_c_1388_n N_VGND_c_1896_n 0.0223802f $X=7.935 $Y=0.45 $X2=0
+ $Y2=0
cc_934 N_A_1464_413#_c_1372_n N_VGND_c_1897_n 0.00583607f $X=9.495 $Y=0.995
+ $X2=0 $Y2=0
cc_935 N_A_1464_413#_M1030_d N_VGND_c_1906_n 0.00482596f $X=7.41 $Y=0.235 $X2=0
+ $Y2=0
cc_936 N_A_1464_413#_c_1372_n N_VGND_c_1906_n 0.0122173f $X=9.495 $Y=0.995 $X2=0
+ $Y2=0
cc_937 N_A_1464_413#_c_1388_n N_VGND_c_1906_n 0.0218104f $X=7.935 $Y=0.45 $X2=0
+ $Y2=0
cc_938 N_A_1464_413#_c_1388_n A_1615_47# 0.00198116f $X=7.935 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_939 N_A_1464_413#_c_1377_n A_1615_47# 0.00129418f $X=8.11 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_940 N_A_2234_47#_c_1463_n N_VPWR_c_1524_n 0.0453754f $X=11.295 $Y=2 $X2=0
+ $Y2=0
cc_941 N_A_2234_47#_c_1463_n N_VPWR_c_1525_n 0.0167768f $X=11.295 $Y=2 $X2=0
+ $Y2=0
cc_942 N_A_2234_47#_c_1461_n N_VPWR_c_1526_n 0.0382543f $X=12.365 $Y=1.41 $X2=0
+ $Y2=0
cc_943 N_A_2234_47#_c_1462_n N_VPWR_c_1526_n 0.0019742f $X=12.835 $Y=1.41 $X2=0
+ $Y2=0
cc_944 N_A_2234_47#_c_1463_n N_VPWR_c_1526_n 0.0606213f $X=11.295 $Y=2 $X2=0
+ $Y2=0
cc_945 N_A_2234_47#_c_1458_n N_VPWR_c_1526_n 0.0489737f $X=12.255 $Y=1.16 $X2=0
+ $Y2=0
cc_946 N_A_2234_47#_c_1460_n N_VPWR_c_1526_n 0.00323466f $X=12.835 $Y=1.202
+ $X2=0 $Y2=0
cc_947 N_A_2234_47#_c_1462_n N_VPWR_c_1528_n 0.0118238f $X=12.835 $Y=1.41 $X2=0
+ $Y2=0
cc_948 N_A_2234_47#_c_1460_n N_VPWR_c_1528_n 3.5734e-19 $X=12.835 $Y=1.202 $X2=0
+ $Y2=0
cc_949 N_A_2234_47#_c_1461_n N_VPWR_c_1539_n 0.00622633f $X=12.365 $Y=1.41 $X2=0
+ $Y2=0
cc_950 N_A_2234_47#_c_1462_n N_VPWR_c_1539_n 0.00650422f $X=12.835 $Y=1.41 $X2=0
+ $Y2=0
cc_951 N_A_2234_47#_M1018_s N_VPWR_c_1517_n 0.00219849f $X=11.17 $Y=1.845 $X2=0
+ $Y2=0
cc_952 N_A_2234_47#_c_1461_n N_VPWR_c_1517_n 0.010479f $X=12.365 $Y=1.41 $X2=0
+ $Y2=0
cc_953 N_A_2234_47#_c_1462_n N_VPWR_c_1517_n 0.0120963f $X=12.835 $Y=1.41 $X2=0
+ $Y2=0
cc_954 N_A_2234_47#_c_1463_n N_VPWR_c_1517_n 0.0122224f $X=11.295 $Y=2 $X2=0
+ $Y2=0
cc_955 N_A_2234_47#_c_1457_n N_Q_c_1844_n 0.00849653f $X=11.295 $Y=0.51 $X2=0
+ $Y2=0
cc_956 N_A_2234_47#_c_1463_n N_Q_c_1844_n 0.00827397f $X=11.295 $Y=2 $X2=0 $Y2=0
cc_957 N_A_2234_47#_c_1459_n N_Q_c_1844_n 0.00861103f $X=11.295 $Y=1.16 $X2=0
+ $Y2=0
cc_958 N_A_2234_47#_c_1461_n N_Q_N_c_1863_n 0.00601391f $X=12.365 $Y=1.41 $X2=0
+ $Y2=0
cc_959 N_A_2234_47#_c_1455_n N_Q_N_c_1863_n 0.00401633f $X=12.39 $Y=0.995 $X2=0
+ $Y2=0
cc_960 N_A_2234_47#_c_1462_n N_Q_N_c_1863_n 0.0146652f $X=12.835 $Y=1.41 $X2=0
+ $Y2=0
cc_961 N_A_2234_47#_c_1456_n N_Q_N_c_1863_n 0.00300534f $X=12.86 $Y=0.995 $X2=0
+ $Y2=0
cc_962 N_A_2234_47#_c_1458_n N_Q_N_c_1863_n 0.0252112f $X=12.255 $Y=1.16 $X2=0
+ $Y2=0
cc_963 N_A_2234_47#_c_1460_n N_Q_N_c_1863_n 0.0418304f $X=12.835 $Y=1.202 $X2=0
+ $Y2=0
cc_964 N_A_2234_47#_c_1457_n N_VGND_c_1885_n 0.0228545f $X=11.295 $Y=0.51 $X2=0
+ $Y2=0
cc_965 N_A_2234_47#_c_1457_n N_VGND_c_1886_n 0.011052f $X=11.295 $Y=0.51 $X2=0
+ $Y2=0
cc_966 N_A_2234_47#_c_1455_n N_VGND_c_1887_n 0.00913159f $X=12.39 $Y=0.995 $X2=0
+ $Y2=0
cc_967 N_A_2234_47#_c_1457_n N_VGND_c_1887_n 0.0170933f $X=11.295 $Y=0.51 $X2=0
+ $Y2=0
cc_968 N_A_2234_47#_c_1458_n N_VGND_c_1887_n 0.0480657f $X=12.255 $Y=1.16 $X2=0
+ $Y2=0
cc_969 N_A_2234_47#_c_1460_n N_VGND_c_1887_n 0.00398003f $X=12.835 $Y=1.202
+ $X2=0 $Y2=0
cc_970 N_A_2234_47#_c_1456_n N_VGND_c_1889_n 0.00595917f $X=12.86 $Y=0.995 $X2=0
+ $Y2=0
cc_971 N_A_2234_47#_c_1455_n N_VGND_c_1899_n 0.00585385f $X=12.39 $Y=0.995 $X2=0
+ $Y2=0
cc_972 N_A_2234_47#_c_1456_n N_VGND_c_1899_n 0.00585385f $X=12.86 $Y=0.995 $X2=0
+ $Y2=0
cc_973 N_A_2234_47#_M1027_s N_VGND_c_1906_n 0.0060859f $X=11.17 $Y=0.235 $X2=0
+ $Y2=0
cc_974 N_A_2234_47#_c_1455_n N_VGND_c_1906_n 0.0115217f $X=12.39 $Y=0.995 $X2=0
+ $Y2=0
cc_975 N_A_2234_47#_c_1456_n N_VGND_c_1906_n 0.0117085f $X=12.86 $Y=0.995 $X2=0
+ $Y2=0
cc_976 N_A_2234_47#_c_1457_n N_VGND_c_1906_n 0.00910216f $X=11.295 $Y=0.51 $X2=0
+ $Y2=0
cc_977 N_VPWR_c_1517_n A_503_369# 0.00287867f $X=13.11 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_978 N_VPWR_c_1517_n N_A_604_369#_M1020_d 0.00192656f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_979 N_VPWR_c_1517_n N_A_604_369#_M1028_s 0.00209341f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_980 N_VPWR_c_1519_n N_A_604_369#_c_1727_n 0.00541311f $X=2.19 $Y=2.33 $X2=0
+ $Y2=0
cc_981 N_VPWR_c_1520_n N_A_604_369#_c_1727_n 0.0109395f $X=4.175 $Y=2.33 $X2=0
+ $Y2=0
cc_982 N_VPWR_c_1529_n N_A_604_369#_c_1727_n 0.0429697f $X=4.09 $Y=2.72 $X2=0
+ $Y2=0
cc_983 N_VPWR_c_1517_n N_A_604_369#_c_1727_n 0.0157065f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_984 N_VPWR_c_1520_n N_A_604_369#_c_1741_n 0.00457937f $X=4.175 $Y=2.33 $X2=0
+ $Y2=0
cc_985 N_VPWR_M1007_d N_A_604_369#_c_1723_n 0.00399644f $X=4.005 $Y=1.845 $X2=0
+ $Y2=0
cc_986 N_VPWR_c_1520_n N_A_604_369#_c_1723_n 0.0119067f $X=4.175 $Y=2.33 $X2=0
+ $Y2=0
cc_987 N_VPWR_c_1529_n N_A_604_369#_c_1723_n 0.00264158f $X=4.09 $Y=2.72 $X2=0
+ $Y2=0
cc_988 N_VPWR_c_1531_n N_A_604_369#_c_1723_n 0.00384075f $X=6.385 $Y=2.72 $X2=0
+ $Y2=0
cc_989 N_VPWR_c_1517_n N_A_604_369#_c_1723_n 0.00546859f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_990 N_VPWR_c_1520_n N_A_604_369#_c_1726_n 0.0159048f $X=4.175 $Y=2.33 $X2=0
+ $Y2=0
cc_991 N_VPWR_c_1531_n N_A_604_369#_c_1726_n 0.017039f $X=6.385 $Y=2.72 $X2=0
+ $Y2=0
cc_992 N_VPWR_c_1517_n N_A_604_369#_c_1726_n 0.0050874f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_993 N_VPWR_c_1517_n A_698_369# 0.00224063f $X=13.11 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_994 N_VPWR_c_1517_n A_1111_413# 0.00234053f $X=13.11 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_995 N_VPWR_c_1517_n A_1558_413# 0.00421708f $X=13.11 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_996 N_VPWR_c_1517_n N_Q_M1003_s 0.00439839f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_997 N_VPWR_c_1523_n N_Q_c_1844_n 0.0531342f $X=9.765 $Y=1.79 $X2=0 $Y2=0
cc_998 N_VPWR_c_1524_n N_Q_c_1844_n 0.0540272f $X=10.775 $Y=1.78 $X2=0 $Y2=0
cc_999 N_VPWR_c_1538_n N_Q_c_1844_n 0.0163795f $X=10.69 $Y=2.72 $X2=0 $Y2=0
cc_1000 N_VPWR_c_1517_n N_Q_c_1844_n 0.010358f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_1001 N_VPWR_c_1517_n N_Q_N_M1005_s 0.0046067f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_1002 N_VPWR_c_1526_n N_Q_N_c_1863_n 0.0544967f $X=11.985 $Y=1.66 $X2=0 $Y2=0
cc_1003 N_VPWR_c_1528_n N_Q_N_c_1863_n 0.0597406f $X=13.07 $Y=1.66 $X2=0 $Y2=0
cc_1004 N_VPWR_c_1539_n N_Q_N_c_1863_n 0.00877801f $X=12.985 $Y=2.72 $X2=0 $Y2=0
cc_1005 N_VPWR_c_1517_n N_Q_N_c_1863_n 0.00933345f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_1006 N_VPWR_c_1528_n N_VGND_c_1889_n 0.00811802f $X=13.07 $Y=1.66 $X2=0 $Y2=0
cc_1007 N_A_604_369#_c_1727_n A_698_369# 0.00415924f $X=3.7 $Y=2.33 $X2=-0.19
+ $Y2=-0.24
cc_1008 N_A_604_369#_c_1741_n A_698_369# 0.00267751f $X=3.785 $Y=2.245 $X2=-0.19
+ $Y2=-0.24
cc_1009 N_A_604_369#_c_1724_n A_698_369# 9.2722e-19 $X=3.87 $Y=1.91 $X2=-0.19
+ $Y2=-0.24
cc_1010 N_A_604_369#_c_1740_n N_VGND_c_1880_n 0.00256403f $X=3.705 $Y=0.36 $X2=0
+ $Y2=0
cc_1011 N_A_604_369#_c_1740_n N_VGND_c_1881_n 0.0109973f $X=3.705 $Y=0.36 $X2=0
+ $Y2=0
cc_1012 N_A_604_369#_c_1716_n N_VGND_c_1881_n 0.00505946f $X=3.79 $Y=0.715 $X2=0
+ $Y2=0
cc_1013 N_A_604_369#_c_1717_n N_VGND_c_1881_n 0.0130184f $X=4.515 $Y=0.8 $X2=0
+ $Y2=0
cc_1014 N_A_604_369#_c_1719_n N_VGND_c_1881_n 5.38578e-19 $X=4.6 $Y=0.715 $X2=0
+ $Y2=0
cc_1015 N_A_604_369#_c_1721_n N_VGND_c_1881_n 0.0100351f $X=4.7 $Y=0.45 $X2=0
+ $Y2=0
cc_1016 N_A_604_369#_c_1740_n N_VGND_c_1892_n 0.0409578f $X=3.705 $Y=0.36 $X2=0
+ $Y2=0
cc_1017 N_A_604_369#_c_1717_n N_VGND_c_1892_n 0.00279549f $X=4.515 $Y=0.8 $X2=0
+ $Y2=0
cc_1018 N_A_604_369#_c_1717_n N_VGND_c_1895_n 0.00291197f $X=4.515 $Y=0.8 $X2=0
+ $Y2=0
cc_1019 N_A_604_369#_c_1721_n N_VGND_c_1895_n 0.012161f $X=4.7 $Y=0.45 $X2=0
+ $Y2=0
cc_1020 N_A_604_369#_M1014_d N_VGND_c_1906_n 0.00171875f $X=3.055 $Y=0.235 $X2=0
+ $Y2=0
cc_1021 N_A_604_369#_M1009_s N_VGND_c_1906_n 0.00134242f $X=4.575 $Y=0.235 $X2=0
+ $Y2=0
cc_1022 N_A_604_369#_c_1740_n N_VGND_c_1906_n 0.00783828f $X=3.705 $Y=0.36 $X2=0
+ $Y2=0
cc_1023 N_A_604_369#_c_1721_n N_VGND_c_1906_n 0.00330494f $X=4.7 $Y=0.45 $X2=0
+ $Y2=0
cc_1024 N_A_604_369#_c_1740_n A_717_47# 0.00220454f $X=3.705 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_1025 N_A_604_369#_c_1716_n A_717_47# 0.00299808f $X=3.79 $Y=0.715 $X2=-0.19
+ $Y2=-0.24
cc_1026 N_Q_c_1844_n N_VGND_c_1898_n 0.0173023f $X=10.295 $Y=0.42 $X2=0 $Y2=0
cc_1027 N_Q_M1013_d N_VGND_c_1906_n 0.00428929f $X=10.16 $Y=0.235 $X2=0 $Y2=0
cc_1028 N_Q_c_1844_n N_VGND_c_1906_n 0.0105927f $X=10.295 $Y=0.42 $X2=0 $Y2=0
cc_1029 N_Q_N_c_1863_n N_VGND_c_1889_n 0.0188376f $X=12.6 $Y=0.63 $X2=0 $Y2=0
cc_1030 N_Q_N_c_1863_n N_VGND_c_1899_n 0.0156894f $X=12.6 $Y=0.63 $X2=0 $Y2=0
cc_1031 N_Q_N_M1004_s N_VGND_c_1906_n 0.00433537f $X=12.465 $Y=0.235 $X2=0 $Y2=0
cc_1032 N_Q_N_c_1863_n N_VGND_c_1906_n 0.0102724f $X=12.6 $Y=0.63 $X2=0 $Y2=0
cc_1033 N_VGND_c_1906_n A_529_47# 0.00151964f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1034 N_VGND_c_1906_n A_717_47# 0.00104569f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1035 N_VGND_c_1906_n A_1117_47# 0.00272292f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1036 N_VGND_c_1906_n A_1615_47# 0.0102544f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
