* File: sky130_fd_sc_hdll__xnor2_1.spice
* Created: Thu Aug 27 19:29:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__xnor2_1.pex.spice"
.subckt sky130_fd_sc_hdll__xnor2_1  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1002 A_139_47# N_B_M1002_g N_A_47_47#_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.2015 PD=0.86 PS=1.92 NRD=9.228 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g A_139_47# VNB NSHORT L=0.15 W=0.65 AD=0.12025
+ AS=0.06825 PD=1.02 PS=0.86 NRD=8.304 NRS=9.228 M=1 R=4.33333 SA=75000.6
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1004 N_A_315_47#_M1004_d N_A_M1004_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_A_315_47#_M1006_d N_B_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.2015 PD=0.97 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1005 N_Y_M1005_d N_A_47_47#_M1005_g N_A_315_47#_M1006_d VNB NSHORT L=0.15
+ W=0.65 AD=0.195 AS=0.104 PD=1.9 PS=0.97 NRD=6.456 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_A_47_47#_M1008_d N_B_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.31 PD=1.29 PS=2.62 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.7 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_47_47#_M1008_d VPB PHIGHVT L=0.18 W=1
+ AD=0.4 AS=0.145 PD=1.8 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.7
+ SB=90002.2 A=0.18 P=2.36 MULT=1
MM1001 A_415_297# N_A_M1001_g N_VPWR_M1003_d VPB PHIGHVT L=0.18 W=1 AD=0.115
+ AS=0.4 PD=1.23 PS=1.8 NRD=11.8003 NRS=0.9653 M=1 R=5.55556 SA=90001.7
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1000 N_Y_M1000_d N_B_M1000_g A_415_297# VPB PHIGHVT L=0.18 W=1 AD=0.175
+ AS=0.115 PD=1.35 PS=1.23 NRD=12.7853 NRS=11.8003 M=1 R=5.55556 SA=90002.1
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A_47_47#_M1009_g N_Y_M1000_d VPB PHIGHVT L=0.18 W=1
+ AD=0.37 AS=0.175 PD=2.74 PS=1.35 NRD=8.8453 NRS=0.9653 M=1 R=5.55556
+ SA=90002.6 SB=90000.3 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
pX11_noxref noxref_12 Y Y PROBETYPE=1
*
.include "sky130_fd_sc_hdll__xnor2_1.pxi.spice"
*
.ends
*
*
