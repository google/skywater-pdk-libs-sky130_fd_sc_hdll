# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a211o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a211o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.535000 1.020000 5.930000 1.330000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.945000 1.020000 5.325000 1.510000 ;
        RECT 4.945000 1.510000 6.445000 1.700000 ;
        RECT 6.125000 1.020000 6.875000 1.320000 ;
        RECT 6.125000 1.320000 6.445000 1.510000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 0.985000 3.105000 1.325000 ;
        RECT 2.875000 1.325000 3.105000 1.445000 ;
        RECT 2.875000 1.445000 4.625000 1.700000 ;
        RECT 4.245000 0.985000 4.625000 1.445000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.275000 0.985000 4.045000 1.275000 ;
    END
  END C1
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN X
    ANTENNADIFFAREA  1.071250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.635000 2.225000 0.875000 ;
        RECT 0.085000 0.875000 0.340000 1.495000 ;
        RECT 0.085000 1.495000 1.790000 1.705000 ;
        RECT 0.645000 1.705000 0.830000 2.465000 ;
        RECT 1.085000 0.255000 1.275000 0.615000 ;
        RECT 1.085000 0.615000 2.225000 0.635000 ;
        RECT 1.600000 1.705000 1.790000 2.465000 ;
        RECT 2.045000 0.255000 2.225000 0.615000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.090000  1.875000 0.425000 2.635000 ;
      RECT 0.485000  0.085000 0.865000 0.465000 ;
      RECT 0.525000  1.045000 2.620000 1.325000 ;
      RECT 1.050000  1.875000 1.380000 2.635000 ;
      RECT 1.445000  0.085000 1.825000 0.445000 ;
      RECT 2.010000  1.835000 2.260000 2.635000 ;
      RECT 2.385000  1.325000 2.620000 1.505000 ;
      RECT 2.385000  1.505000 2.705000 1.675000 ;
      RECT 2.395000  0.615000 6.040000 0.805000 ;
      RECT 2.395000  0.805000 2.620000 1.045000 ;
      RECT 2.420000  0.085000 2.805000 0.445000 ;
      RECT 2.530000  1.675000 2.705000 1.870000 ;
      RECT 2.530000  1.870000 3.860000 2.040000 ;
      RECT 2.570000  2.210000 4.900000 2.465000 ;
      RECT 3.025000  0.255000 3.270000 0.615000 ;
      RECT 3.440000  0.085000 3.820000 0.445000 ;
      RECT 4.040000  0.255000 4.420000 0.615000 ;
      RECT 4.570000  1.880000 6.995000 2.105000 ;
      RECT 4.570000  2.105000 4.900000 2.210000 ;
      RECT 4.640000  0.085000 5.010000 0.445000 ;
      RECT 5.070000  2.275000 5.450000 2.635000 ;
      RECT 5.660000  0.275000 6.040000 0.615000 ;
      RECT 5.660000  2.105000 5.970000 2.465000 ;
      RECT 6.140000  2.275000 6.520000 2.635000 ;
      RECT 6.615000  0.085000 6.995000 0.805000 ;
      RECT 6.615000  1.535000 6.995000 1.880000 ;
      RECT 6.740000  2.105000 6.995000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a211o_4
END LIBRARY
