* NGSPICE file created from sky130_fd_sc_hdll__a22o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 a_1008_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=3.835e+11p pd=3.78e+06u as=1.3975e+12p ps=1.08e+07u
M1001 X a_96_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=1.43e+12p ps=1.286e+07u
M1002 VPWR A2 a_524_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.515e+12p ps=1.303e+07u
M1003 a_96_21# B1 a_524_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1004 VGND A2 a_1008_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_96_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_524_297# B1 a_96_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_96_21# VGND VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=0p ps=0u
M1008 VGND a_96_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_616_47# B1 a_96_21# VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=4.81e+11p ps=4.08e+06u
M1010 a_524_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1008_47# A1 a_96_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_96_21# B2 a_524_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_96_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND B2 a_616_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_96_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_96_21# B1 a_616_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A1 a_524_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_96_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_616_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_96_21# A1 a_1008_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_524_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_96_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_524_297# B2 a_96_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

