* File: sky130_fd_sc_hdll__a32oi_2.pxi.spice
* Created: Thu Aug 27 18:56:31 2020
* 
x_PM_SKY130_FD_SC_HDLL__A32OI_2%B2 N_B2_c_78_n N_B2_M1001_g N_B2_c_73_n
+ N_B2_M1002_g N_B2_c_79_n N_B2_M1007_g N_B2_c_74_n N_B2_M1014_g B2 B2 B2
+ N_B2_c_76_n N_B2_c_77_n PM_SKY130_FD_SC_HDLL__A32OI_2%B2
x_PM_SKY130_FD_SC_HDLL__A32OI_2%B1 N_B1_c_122_n N_B1_M1004_g N_B1_c_126_n
+ N_B1_M1013_g N_B1_c_127_n N_B1_M1018_g N_B1_c_123_n N_B1_M1015_g B1 B1
+ N_B1_c_125_n B1 PM_SKY130_FD_SC_HDLL__A32OI_2%B1
x_PM_SKY130_FD_SC_HDLL__A32OI_2%A1 N_A1_c_180_n N_A1_M1003_g N_A1_c_175_n
+ N_A1_c_176_n N_A1_M1011_g N_A1_c_182_n N_A1_M1010_g N_A1_M1012_g A1 A1
+ N_A1_c_186_n N_A1_c_179_n A1 A1 PM_SKY130_FD_SC_HDLL__A32OI_2%A1
x_PM_SKY130_FD_SC_HDLL__A32OI_2%A2 N_A2_M1008_g N_A2_c_229_n N_A2_M1000_g
+ N_A2_M1016_g N_A2_c_230_n N_A2_M1017_g A2 A2 N_A2_c_228_n A2 A2
+ PM_SKY130_FD_SC_HDLL__A32OI_2%A2
x_PM_SKY130_FD_SC_HDLL__A32OI_2%A3 N_A3_c_276_n N_A3_M1005_g N_A3_M1006_g
+ N_A3_c_277_n N_A3_M1009_g N_A3_M1019_g N_A3_c_272_n A3 A3 A3 A3 A3
+ N_A3_c_274_n N_A3_c_275_n A3 PM_SKY130_FD_SC_HDLL__A32OI_2%A3
x_PM_SKY130_FD_SC_HDLL__A32OI_2%A_27_297# N_A_27_297#_M1001_d
+ N_A_27_297#_M1007_d N_A_27_297#_M1018_d N_A_27_297#_M1010_d
+ N_A_27_297#_M1017_s N_A_27_297#_M1009_d N_A_27_297#_c_319_n
+ N_A_27_297#_c_322_n N_A_27_297#_c_370_p N_A_27_297#_c_345_p
+ N_A_27_297#_c_324_n N_A_27_297#_c_352_p N_A_27_297#_c_353_p
+ N_A_27_297#_c_326_n N_A_27_297#_c_330_n N_A_27_297#_c_335_n
+ N_A_27_297#_c_375_p N_A_27_297#_c_376_p N_A_27_297#_c_377_p
+ N_A_27_297#_c_339_n PM_SKY130_FD_SC_HDLL__A32OI_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A32OI_2%Y N_Y_M1004_d N_Y_M1011_s N_Y_M1001_s
+ N_Y_M1013_s N_Y_c_404_n N_Y_c_399_n N_Y_c_400_n N_Y_c_417_n N_Y_c_421_n
+ N_Y_c_401_n N_Y_c_397_n N_Y_c_402_n Y Y Y N_Y_c_429_n Y
+ PM_SKY130_FD_SC_HDLL__A32OI_2%Y
x_PM_SKY130_FD_SC_HDLL__A32OI_2%VPWR N_VPWR_M1003_s N_VPWR_M1000_d
+ N_VPWR_M1005_s VPWR N_VPWR_c_485_n N_VPWR_c_484_n N_VPWR_c_487_n
+ N_VPWR_c_488_n N_VPWR_c_489_n N_VPWR_c_490_n N_VPWR_c_491_n N_VPWR_c_492_n
+ PM_SKY130_FD_SC_HDLL__A32OI_2%VPWR
x_PM_SKY130_FD_SC_HDLL__A32OI_2%A_27_47# N_A_27_47#_M1002_d N_A_27_47#_M1014_d
+ N_A_27_47#_M1015_s N_A_27_47#_c_566_n N_A_27_47#_c_570_n N_A_27_47#_c_567_n
+ N_A_27_47#_c_577_n N_A_27_47#_c_568_n N_A_27_47#_c_569_n
+ PM_SKY130_FD_SC_HDLL__A32OI_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__A32OI_2%VGND N_VGND_M1002_s N_VGND_M1006_d
+ N_VGND_M1019_d N_VGND_c_610_n N_VGND_c_611_n N_VGND_c_612_n N_VGND_c_613_n
+ VGND N_VGND_c_614_n N_VGND_c_615_n N_VGND_c_616_n
+ PM_SKY130_FD_SC_HDLL__A32OI_2%VGND
x_PM_SKY130_FD_SC_HDLL__A32OI_2%A_507_47# N_A_507_47#_M1011_d
+ N_A_507_47#_M1012_d N_A_507_47#_M1016_d N_A_507_47#_c_677_n
+ PM_SKY130_FD_SC_HDLL__A32OI_2%A_507_47#
x_PM_SKY130_FD_SC_HDLL__A32OI_2%A_757_47# N_A_757_47#_M1008_s
+ N_A_757_47#_M1006_s N_A_757_47#_c_696_n N_A_757_47#_c_705_n
+ PM_SKY130_FD_SC_HDLL__A32OI_2%A_757_47#
cc_1 VNB N_B2_c_73_n 0.0223829f $X=-0.195 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB N_B2_c_74_n 0.0166793f $X=-0.195 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB B2 6.57328e-19 $X=-0.195 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_4 VNB N_B2_c_76_n 0.0557501f $X=-0.195 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_5 VNB N_B2_c_77_n 0.00864012f $X=-0.195 $Y=-0.24 $X2=0.235 $Y2=1.285
cc_6 VNB N_B1_c_122_n 0.016055f $X=-0.195 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_7 VNB N_B1_c_123_n 0.0195547f $X=-0.195 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_8 VNB B1 0.00606283f $X=-0.195 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_9 VNB N_B1_c_125_n 0.0447809f $X=-0.195 $Y=-0.24 $X2=0.71 $Y2=1.16
cc_10 VNB N_A1_c_175_n 0.0258737f $X=-0.195 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_11 VNB N_A1_c_176_n 0.0168792f $X=-0.195 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_12 VNB N_A1_M1011_g 0.0220338f $X=-0.195 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_13 VNB N_A1_M1012_g 0.017802f $X=-0.195 $Y=-0.24 $X2=0.625 $Y2=1.105
cc_14 VNB N_A1_c_179_n 0.0349865f $X=-0.195 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A2_M1008_g 0.0183466f $X=-0.195 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_16 VNB N_A2_M1016_g 0.0249276f $X=-0.195 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_17 VNB N_A2_c_228_n 0.0717265f $X=-0.195 $Y=-0.24 $X2=0.235 $Y2=1.53
cc_18 VNB N_A3_M1006_g 0.0258898f $X=-0.195 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_19 VNB N_A3_M1019_g 0.0250322f $X=-0.195 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_20 VNB N_A3_c_272_n 0.0420443f $X=-0.195 $Y=-0.24 $X2=0.625 $Y2=1.105
cc_21 VNB A3 0.00932659f $X=-0.195 $Y=-0.24 $X2=0.71 $Y2=1.16
cc_22 VNB N_A3_c_274_n 0.0270733f $X=-0.195 $Y=-0.24 $X2=0.325 $Y2=1.18
cc_23 VNB N_A3_c_275_n 0.0342242f $X=-0.195 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_Y_c_397_n 0.00730405f $X=-0.195 $Y=-0.24 $X2=0.695 $Y2=1.18
cc_25 VNB Y 0.00401828f $X=-0.195 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_484_n 0.269736f $X=-0.195 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_566_n 0.0165239f $X=-0.195 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_28 VNB N_A_27_47#_c_567_n 0.0106747f $X=-0.195 $Y=-0.24 $X2=0.625 $Y2=1.105
cc_29 VNB N_A_27_47#_c_568_n 0.00151873f $X=-0.195 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_27_47#_c_569_n 0.00214428f $X=-0.195 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_31 VNB N_VGND_c_610_n 0.00472845f $X=-0.195 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_32 VNB N_VGND_c_611_n 0.0110531f $X=-0.195 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_612_n 0.00574094f $X=-0.195 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_613_n 0.113238f $X=-0.195 $Y=-0.24 $X2=0.71 $Y2=1.202
cc_35 VNB N_VGND_c_614_n 0.0226698f $X=-0.195 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_615_n 0.0222151f $X=-0.195 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_616_n 0.322575f $X=-0.195 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_507_47#_c_677_n 0.00588558f $X=-0.195 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_757_47#_c_696_n 0.0171405f $X=-0.195 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_40 VPB N_B2_c_78_n 0.0190112f $X=-0.195 $Y=1.305 $X2=0.495 $Y2=1.41
cc_41 VPB N_B2_c_79_n 0.0161009f $X=-0.195 $Y=1.305 $X2=0.965 $Y2=1.41
cc_42 VPB B2 0.00761758f $X=-0.195 $Y=1.305 $X2=0.15 $Y2=1.445
cc_43 VPB N_B2_c_76_n 0.0288252f $X=-0.195 $Y=1.305 $X2=0.965 $Y2=1.202
cc_44 VPB N_B1_c_126_n 0.0160857f $X=-0.195 $Y=1.305 $X2=0.52 $Y2=0.995
cc_45 VPB N_B1_c_127_n 0.0158275f $X=-0.195 $Y=1.305 $X2=0.965 $Y2=1.41
cc_46 VPB N_B1_c_125_n 0.012412f $X=-0.195 $Y=1.305 $X2=0.71 $Y2=1.16
cc_47 VPB N_A1_c_180_n 0.0180073f $X=-0.195 $Y=1.305 $X2=0.495 $Y2=1.41
cc_48 VPB N_A1_c_176_n 0.00723915f $X=-0.195 $Y=1.305 $X2=0.52 $Y2=0.56
cc_49 VPB N_A1_c_182_n 0.0183492f $X=-0.195 $Y=1.305 $X2=0.99 $Y2=0.995
cc_50 VPB N_A1_c_179_n 0.00727992f $X=-0.195 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A2_c_229_n 0.0175941f $X=-0.195 $Y=1.305 $X2=0.52 $Y2=0.56
cc_52 VPB N_A2_c_230_n 0.0175864f $X=-0.195 $Y=1.305 $X2=0.99 $Y2=0.56
cc_53 VPB N_A2_c_228_n 0.0143264f $X=-0.195 $Y=1.305 $X2=0.235 $Y2=1.53
cc_54 VPB N_A3_c_276_n 0.0198686f $X=-0.195 $Y=1.305 $X2=0.495 $Y2=1.41
cc_55 VPB N_A3_c_277_n 0.0229729f $X=-0.195 $Y=1.305 $X2=0.965 $Y2=1.985
cc_56 VPB N_A3_c_272_n 0.00734255f $X=-0.195 $Y=1.305 $X2=0.625 $Y2=1.105
cc_57 VPB A3 0.0137974f $X=-0.195 $Y=1.305 $X2=0.71 $Y2=1.16
cc_58 VPB N_A3_c_275_n 0.0161937f $X=-0.195 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_Y_c_399_n 0.00297822f $X=-0.195 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_Y_c_400_n 0.00174853f $X=-0.195 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_Y_c_401_n 4.02974e-19 $X=-0.195 $Y=1.305 $X2=0.235 $Y2=1.53
cc_62 VPB N_Y_c_402_n 0.00102672f $X=-0.195 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB Y 9.35342e-19 $X=-0.195 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_485_n 0.0186134f $X=-0.195 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_484_n 0.0473008f $X=-0.195 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_487_n 0.0582958f $X=-0.195 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_488_n 0.0170733f $X=-0.195 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_489_n 0.0141177f $X=-0.195 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_490_n 0.0134558f $X=-0.195 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_491_n 0.0139761f $X=-0.195 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_492_n 0.0210296f $X=-0.195 $Y=1.305 $X2=0 $Y2=0
cc_72 N_B2_c_74_n N_B1_c_122_n 0.0175843f $X=0.99 $Y=0.995 $X2=-0.195 $Y2=-0.24
cc_73 N_B2_c_79_n N_B1_c_126_n 0.02168f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_74 B2 B1 0.0160896f $X=0.625 $Y=1.105 $X2=0 $Y2=0
cc_75 N_B2_c_76_n B1 0.00235992f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_76 N_B2_c_76_n N_B1_c_125_n 0.0175843f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_77 B2 N_A_27_297#_M1001_d 0.0108175f $X=0.15 $Y=1.445 $X2=-0.195 $Y2=-0.24
cc_78 B2 N_A_27_297#_c_319_n 0.0131226f $X=0.15 $Y=1.445 $X2=0 $Y2=0
cc_79 B2 N_A_27_297#_c_319_n 6.33088e-19 $X=0.625 $Y=1.105 $X2=0 $Y2=0
cc_80 N_B2_c_76_n N_A_27_297#_c_319_n 0.00100981f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_81 N_B2_c_78_n N_A_27_297#_c_322_n 0.0137768f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_82 N_B2_c_79_n N_A_27_297#_c_322_n 0.0112487f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_83 N_B2_c_78_n N_Y_c_404_n 0.0116496f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_84 N_B2_c_79_n N_Y_c_404_n 0.00726135f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_85 N_B2_c_79_n N_Y_c_399_n 0.0133552f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_86 N_B2_c_76_n N_Y_c_399_n 3.5658e-19 $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_87 N_B2_c_78_n N_Y_c_400_n 0.00308953f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_88 N_B2_c_79_n N_Y_c_400_n 0.00146147f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_89 B2 N_Y_c_400_n 0.0103134f $X=0.15 $Y=1.445 $X2=0 $Y2=0
cc_90 B2 N_Y_c_400_n 0.0252371f $X=0.625 $Y=1.105 $X2=0 $Y2=0
cc_91 N_B2_c_76_n N_Y_c_400_n 0.00775434f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_92 N_B2_c_78_n N_VPWR_c_484_n 0.00697643f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_93 N_B2_c_79_n N_VPWR_c_484_n 0.00609021f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_94 N_B2_c_78_n N_VPWR_c_487_n 0.00429453f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_95 N_B2_c_79_n N_VPWR_c_487_n 0.00429453f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_96 N_B2_c_73_n N_A_27_47#_c_570_n 0.0104412f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_97 N_B2_c_74_n N_A_27_47#_c_570_n 0.0102701f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_98 B2 N_A_27_47#_c_570_n 0.0259185f $X=0.625 $Y=1.105 $X2=0 $Y2=0
cc_99 N_B2_c_76_n N_A_27_47#_c_570_n 0.00340637f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_100 B2 N_A_27_47#_c_567_n 0.00573168f $X=0.625 $Y=1.105 $X2=0 $Y2=0
cc_101 N_B2_c_76_n N_A_27_47#_c_567_n 0.00677682f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_102 N_B2_c_77_n N_A_27_47#_c_567_n 0.0140961f $X=0.235 $Y=1.285 $X2=0 $Y2=0
cc_103 N_B2_c_74_n N_A_27_47#_c_577_n 0.00229336f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_104 N_B2_c_73_n N_A_27_47#_c_568_n 4.8427e-19 $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_105 N_B2_c_74_n N_A_27_47#_c_568_n 0.00542267f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_106 N_B2_c_73_n N_VGND_c_610_n 0.00276126f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_107 N_B2_c_74_n N_VGND_c_610_n 0.00437853f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_108 N_B2_c_74_n N_VGND_c_613_n 0.00422371f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_109 N_B2_c_73_n N_VGND_c_615_n 0.00436487f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_110 N_B2_c_73_n N_VGND_c_616_n 0.00698799f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_111 N_B2_c_74_n N_VGND_c_616_n 0.0059854f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_112 N_B1_c_127_n N_A1_c_180_n 0.0211043f $X=1.905 $Y=1.41 $X2=-0.195
+ $Y2=-0.24
cc_113 N_B1_c_125_n N_A1_c_176_n 0.0177293f $X=1.905 $Y=1.192 $X2=0 $Y2=0
cc_114 N_B1_c_125_n N_A1_c_186_n 2.6501e-19 $X=1.905 $Y=1.192 $X2=0 $Y2=0
cc_115 N_B1_c_126_n N_A_27_297#_c_324_n 0.0115669f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_116 N_B1_c_127_n N_A_27_297#_c_324_n 0.0115805f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_117 N_B1_c_126_n N_Y_c_404_n 8.27825e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_118 N_B1_c_126_n N_Y_c_399_n 0.0145582f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_119 B1 N_Y_c_399_n 0.0381122f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_120 N_B1_c_125_n N_Y_c_399_n 0.00190063f $X=1.905 $Y=1.192 $X2=0 $Y2=0
cc_121 N_B1_c_122_n N_Y_c_417_n 0.00266083f $X=1.41 $Y=0.975 $X2=0 $Y2=0
cc_122 N_B1_c_123_n N_Y_c_417_n 0.00622332f $X=1.93 $Y=0.975 $X2=0 $Y2=0
cc_123 B1 N_Y_c_417_n 0.0163828f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_124 N_B1_c_125_n N_Y_c_417_n 0.00451586f $X=1.905 $Y=1.192 $X2=0 $Y2=0
cc_125 N_B1_c_126_n N_Y_c_421_n 0.00543807f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_126 N_B1_c_127_n N_Y_c_421_n 0.00543583f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_127 N_B1_c_127_n N_Y_c_401_n 0.0128196f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_128 B1 N_Y_c_401_n 0.00286809f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_129 N_B1_c_125_n N_Y_c_401_n 0.00169959f $X=1.905 $Y=1.192 $X2=0 $Y2=0
cc_130 B1 N_Y_c_402_n 0.0138898f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_131 N_B1_c_125_n N_Y_c_402_n 0.00397531f $X=1.905 $Y=1.192 $X2=0 $Y2=0
cc_132 N_B1_c_123_n Y 0.00534332f $X=1.93 $Y=0.975 $X2=0 $Y2=0
cc_133 N_B1_c_127_n N_Y_c_429_n 0.00285969f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_134 N_B1_c_122_n Y 5.69995e-19 $X=1.41 $Y=0.975 $X2=0 $Y2=0
cc_135 N_B1_c_126_n Y 2.06485e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_136 N_B1_c_127_n Y 0.00118503f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_137 N_B1_c_123_n Y 0.00566227f $X=1.93 $Y=0.975 $X2=0 $Y2=0
cc_138 B1 Y 0.0161814f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_139 N_B1_c_125_n Y 0.0160029f $X=1.905 $Y=1.192 $X2=0 $Y2=0
cc_140 N_B1_c_126_n N_VPWR_c_484_n 0.00609021f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_141 N_B1_c_127_n N_VPWR_c_484_n 0.00609021f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_142 N_B1_c_126_n N_VPWR_c_487_n 0.00429453f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_143 N_B1_c_127_n N_VPWR_c_487_n 0.00429453f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_144 N_B1_c_127_n N_VPWR_c_488_n 0.00105559f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_145 B1 N_A_27_47#_c_568_n 0.0142485f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_146 N_B1_c_122_n N_A_27_47#_c_569_n 0.010118f $X=1.41 $Y=0.975 $X2=0 $Y2=0
cc_147 N_B1_c_123_n N_A_27_47#_c_569_n 0.00856614f $X=1.93 $Y=0.975 $X2=0 $Y2=0
cc_148 B1 N_A_27_47#_c_569_n 0.00365692f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_149 N_B1_c_122_n N_VGND_c_613_n 0.00366111f $X=1.41 $Y=0.975 $X2=0 $Y2=0
cc_150 N_B1_c_123_n N_VGND_c_613_n 0.00366111f $X=1.93 $Y=0.975 $X2=0 $Y2=0
cc_151 N_B1_c_122_n N_VGND_c_616_n 0.00551892f $X=1.41 $Y=0.975 $X2=0 $Y2=0
cc_152 N_B1_c_123_n N_VGND_c_616_n 0.00681779f $X=1.93 $Y=0.975 $X2=0 $Y2=0
cc_153 N_A1_M1012_g N_A2_M1008_g 0.0242938f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_154 N_A1_c_182_n N_A2_c_229_n 0.0217955f $X=3.265 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A1_c_186_n N_A2_c_229_n 6.61778e-19 $X=3 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A1_c_186_n N_A2_c_228_n 0.0011995f $X=3 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A1_c_179_n N_A2_c_228_n 0.0242938f $X=3.265 $Y=1.217 $X2=0 $Y2=0
cc_158 N_A1_c_182_n A2 6.95708e-19 $X=3.265 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A1_c_186_n A2 0.0203366f $X=3 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A1_c_179_n A2 0.00126078f $X=3.265 $Y=1.217 $X2=0 $Y2=0
cc_161 N_A1_c_180_n N_A_27_297#_c_326_n 0.0160889f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A1_c_175_n N_A_27_297#_c_326_n 0.00227113f $X=2.795 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A1_c_182_n N_A_27_297#_c_326_n 0.0163779f $X=3.265 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A1_c_186_n N_A_27_297#_c_326_n 0.0600964f $X=3 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A1_c_176_n N_Y_c_397_n 0.0133122f $X=2.475 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A1_M1011_g N_Y_c_397_n 0.0110467f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_167 N_A1_M1012_g N_Y_c_397_n 0.0038838f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_168 N_A1_c_186_n N_Y_c_397_n 0.0447212f $X=3 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A1_c_179_n N_Y_c_397_n 0.00194825f $X=3.265 $Y=1.217 $X2=0 $Y2=0
cc_170 N_A1_c_180_n N_Y_c_429_n 0.00137947f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A1_c_186_n N_Y_c_429_n 0.014179f $X=3 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A1_c_180_n Y 3.13013e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A1_c_176_n Y 0.00400549f $X=2.475 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A1_M1011_g Y 0.00451941f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_175 N_A1_c_186_n Y 0.0295633f $X=3 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A1_c_186_n N_VPWR_M1003_s 0.00916097f $X=3 $Y=1.16 $X2=-0.195 $Y2=-0.24
cc_177 N_A1_c_180_n N_VPWR_c_484_n 0.00546112f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A1_c_182_n N_VPWR_c_484_n 0.00764137f $X=3.265 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A1_c_180_n N_VPWR_c_487_n 0.00470513f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A1_c_180_n N_VPWR_c_488_n 0.00907217f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A1_c_182_n N_VPWR_c_488_n 0.00238515f $X=3.265 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A1_c_182_n N_VPWR_c_489_n 0.00412417f $X=3.265 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A1_c_182_n N_VPWR_c_490_n 5.54128e-19 $X=3.265 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A1_M1011_g N_VGND_c_613_n 0.00366111f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_185 N_A1_M1012_g N_VGND_c_613_n 0.00366111f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_186 N_A1_M1011_g N_VGND_c_616_n 0.00656615f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_187 N_A1_M1012_g N_VGND_c_616_n 0.00526729f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_188 N_A1_M1011_g N_A_507_47#_c_677_n 0.00801257f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_189 N_A1_M1012_g N_A_507_47#_c_677_n 0.0113833f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_190 N_A1_c_186_n N_A_507_47#_c_677_n 2.58419e-19 $X=3 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A1_M1012_g N_A_757_47#_c_696_n 5.30585e-19 $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_192 N_A2_c_230_n N_A3_c_276_n 0.0209655f $X=4.545 $Y=1.41 $X2=-0.195
+ $Y2=-0.24
cc_193 A2 N_A3_c_276_n 7.14961e-19 $X=4.365 $Y=1.19 $X2=-0.195 $Y2=-0.24
cc_194 N_A2_c_228_n N_A3_c_272_n 0.0190496f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_195 A2 N_A3_c_272_n 0.0013001f $X=4.365 $Y=1.19 $X2=0 $Y2=0
cc_196 N_A2_c_230_n A3 6.73468e-19 $X=4.545 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A2_c_228_n A3 0.00122491f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_198 A2 A3 0.0209182f $X=4.365 $Y=1.19 $X2=0 $Y2=0
cc_199 N_A2_c_229_n N_A_27_297#_c_330_n 0.0149571f $X=3.735 $Y=1.41 $X2=0 $Y2=0
cc_200 N_A2_c_230_n N_A_27_297#_c_330_n 0.014379f $X=4.545 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A2_c_228_n N_A_27_297#_c_330_n 0.00199706f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_202 A2 N_A_27_297#_c_330_n 0.0578242f $X=4.365 $Y=1.19 $X2=0 $Y2=0
cc_203 N_A2_M1008_g N_Y_c_397_n 5.30585e-19 $X=3.71 $Y=0.56 $X2=0 $Y2=0
cc_204 A2 N_VPWR_M1000_d 0.00766166f $X=4.365 $Y=1.19 $X2=0 $Y2=0
cc_205 N_A2_c_229_n N_VPWR_c_484_n 0.00439345f $X=3.735 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A2_c_230_n N_VPWR_c_484_n 0.00395957f $X=4.545 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A2_c_229_n N_VPWR_c_489_n 0.00220938f $X=3.735 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A2_c_229_n N_VPWR_c_490_n 0.0100685f $X=3.735 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A2_c_230_n N_VPWR_c_490_n 0.0109248f $X=4.545 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A2_c_230_n N_VPWR_c_491_n 0.0017675f $X=4.545 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A2_M1008_g N_VGND_c_613_n 0.00366111f $X=3.71 $Y=0.56 $X2=0 $Y2=0
cc_212 N_A2_M1016_g N_VGND_c_613_n 0.00614817f $X=4.18 $Y=0.56 $X2=0 $Y2=0
cc_213 N_A2_M1008_g N_VGND_c_616_n 0.00539914f $X=3.71 $Y=0.56 $X2=0 $Y2=0
cc_214 N_A2_M1016_g N_VGND_c_616_n 0.00669801f $X=4.18 $Y=0.56 $X2=0 $Y2=0
cc_215 N_A2_M1008_g N_A_507_47#_c_677_n 0.0112375f $X=3.71 $Y=0.56 $X2=0 $Y2=0
cc_216 N_A2_M1016_g N_A_507_47#_c_677_n 0.00818766f $X=4.18 $Y=0.56 $X2=0 $Y2=0
cc_217 A2 N_A_507_47#_c_677_n 9.04466e-19 $X=4.365 $Y=1.19 $X2=0 $Y2=0
cc_218 N_A2_M1008_g N_A_757_47#_c_696_n 0.00388163f $X=3.71 $Y=0.56 $X2=0 $Y2=0
cc_219 N_A2_M1016_g N_A_757_47#_c_696_n 0.0110355f $X=4.18 $Y=0.56 $X2=0 $Y2=0
cc_220 N_A2_c_228_n N_A_757_47#_c_696_n 0.0129334f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_221 A2 N_A_757_47#_c_696_n 0.0393572f $X=4.365 $Y=1.19 $X2=0 $Y2=0
cc_222 A3 N_A_27_297#_M1009_d 0.00426621f $X=6.11 $Y=1.105 $X2=0 $Y2=0
cc_223 N_A3_c_276_n N_A_27_297#_c_335_n 0.0165615f $X=5.025 $Y=1.41 $X2=0 $Y2=0
cc_224 N_A3_c_277_n N_A_27_297#_c_335_n 0.0140197f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A3_c_272_n N_A_27_297#_c_335_n 0.00237574f $X=5.475 $Y=1.16 $X2=0 $Y2=0
cc_226 A3 N_A_27_297#_c_335_n 0.0700262f $X=6.11 $Y=1.105 $X2=0 $Y2=0
cc_227 A3 N_A_27_297#_c_339_n 0.0150029f $X=6.11 $Y=1.105 $X2=0 $Y2=0
cc_228 N_A3_c_275_n N_A_27_297#_c_339_n 6.78074e-19 $X=5.97 $Y=1.212 $X2=0 $Y2=0
cc_229 A3 N_VPWR_M1005_s 0.00972321f $X=6.11 $Y=1.105 $X2=0 $Y2=0
cc_230 N_A3_c_277_n N_VPWR_c_485_n 0.0053025f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_231 N_A3_c_276_n N_VPWR_c_484_n 0.00820862f $X=5.025 $Y=1.41 $X2=0 $Y2=0
cc_232 N_A3_c_277_n N_VPWR_c_484_n 0.00907115f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_233 N_A3_c_276_n N_VPWR_c_490_n 5.60508e-19 $X=5.025 $Y=1.41 $X2=0 $Y2=0
cc_234 N_A3_c_276_n N_VPWR_c_491_n 0.00412417f $X=5.025 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A3_c_276_n N_VPWR_c_492_n 0.00360215f $X=5.025 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A3_c_277_n N_VPWR_c_492_n 0.00523602f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_237 N_A3_M1019_g N_VGND_c_612_n 0.00438629f $X=5.97 $Y=0.56 $X2=0 $Y2=0
cc_238 A3 N_VGND_c_612_n 0.0129521f $X=6.11 $Y=1.105 $X2=0 $Y2=0
cc_239 N_A3_c_275_n N_VGND_c_612_n 0.00404225f $X=5.97 $Y=1.212 $X2=0 $Y2=0
cc_240 N_A3_M1006_g N_VGND_c_613_n 0.0101966f $X=5.4 $Y=0.56 $X2=0 $Y2=0
cc_241 N_A3_M1006_g N_VGND_c_614_n 0.00403386f $X=5.4 $Y=0.56 $X2=0 $Y2=0
cc_242 N_A3_M1019_g N_VGND_c_614_n 0.00585385f $X=5.97 $Y=0.56 $X2=0 $Y2=0
cc_243 N_A3_M1006_g N_VGND_c_616_n 0.00727001f $X=5.4 $Y=0.56 $X2=0 $Y2=0
cc_244 N_A3_M1019_g N_VGND_c_616_n 0.0119276f $X=5.97 $Y=0.56 $X2=0 $Y2=0
cc_245 N_A3_M1006_g N_A_757_47#_c_696_n 0.0103949f $X=5.4 $Y=0.56 $X2=0 $Y2=0
cc_246 N_A3_c_272_n N_A_757_47#_c_696_n 0.010561f $X=5.475 $Y=1.16 $X2=0 $Y2=0
cc_247 A3 N_A_757_47#_c_696_n 0.0195748f $X=6.11 $Y=1.105 $X2=0 $Y2=0
cc_248 N_A3_M1006_g N_A_757_47#_c_705_n 0.0132038f $X=5.4 $Y=0.56 $X2=0 $Y2=0
cc_249 N_A3_M1019_g N_A_757_47#_c_705_n 0.00558621f $X=5.97 $Y=0.56 $X2=0 $Y2=0
cc_250 A3 N_A_757_47#_c_705_n 0.0202833f $X=6.11 $Y=1.105 $X2=0 $Y2=0
cc_251 N_A3_c_274_n N_A_757_47#_c_705_n 0.00520972f $X=5.845 $Y=1.16 $X2=0 $Y2=0
cc_252 N_A_27_297#_c_322_n N_Y_M1001_s 0.00352392f $X=1.115 $Y=2.38 $X2=0.495
+ $Y2=1.985
cc_253 N_A_27_297#_c_324_n N_Y_M1013_s 0.00343888f $X=2.055 $Y=2.38 $X2=0.52
+ $Y2=0.995
cc_254 N_A_27_297#_c_319_n N_Y_c_404_n 0.0199789f $X=0.26 $Y=1.96 $X2=0.625
+ $Y2=1.105
cc_255 N_A_27_297#_c_322_n N_Y_c_404_n 0.016028f $X=1.115 $Y=2.38 $X2=0.625
+ $Y2=1.105
cc_256 N_A_27_297#_c_345_p N_Y_c_404_n 0.0199789f $X=1.2 $Y=1.96 $X2=0.625
+ $Y2=1.105
cc_257 N_A_27_297#_M1007_d N_Y_c_399_n 0.00178587f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_258 N_A_27_297#_c_322_n N_Y_c_399_n 0.00346334f $X=1.115 $Y=2.38 $X2=0 $Y2=0
cc_259 N_A_27_297#_c_345_p N_Y_c_399_n 0.0136517f $X=1.2 $Y=1.96 $X2=0 $Y2=0
cc_260 N_A_27_297#_c_324_n N_Y_c_399_n 0.00394364f $X=2.055 $Y=2.38 $X2=0 $Y2=0
cc_261 N_A_27_297#_c_345_p N_Y_c_421_n 0.0157757f $X=1.2 $Y=1.96 $X2=0.99
+ $Y2=1.202
cc_262 N_A_27_297#_c_324_n N_Y_c_421_n 0.0127862f $X=2.055 $Y=2.38 $X2=0.99
+ $Y2=1.202
cc_263 N_A_27_297#_c_352_p N_Y_c_421_n 0.00908546f $X=2.14 $Y=1.965 $X2=0.99
+ $Y2=1.202
cc_264 N_A_27_297#_c_353_p N_Y_c_421_n 0.00762492f $X=2.14 $Y=2.295 $X2=0.99
+ $Y2=1.202
cc_265 N_A_27_297#_c_324_n N_Y_c_401_n 0.00325872f $X=2.055 $Y=2.38 $X2=0.235
+ $Y2=1.53
cc_266 N_A_27_297#_M1018_d N_Y_c_429_n 0.00284406f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_267 N_A_27_297#_c_324_n N_Y_c_429_n 7.47417e-19 $X=2.055 $Y=2.38 $X2=0 $Y2=0
cc_268 N_A_27_297#_c_352_p N_Y_c_429_n 0.0126088f $X=2.14 $Y=1.965 $X2=0 $Y2=0
cc_269 N_A_27_297#_c_326_n N_VPWR_M1003_s 0.0167687f $X=3.415 $Y=1.88 $X2=0.495
+ $Y2=1.41
cc_270 N_A_27_297#_c_330_n N_VPWR_M1000_d 0.0142108f $X=4.695 $Y=1.88 $X2=0.495
+ $Y2=1.985
cc_271 N_A_27_297#_c_335_n N_VPWR_M1005_s 0.0177279f $X=6.095 $Y=1.88 $X2=0.495
+ $Y2=1.985
cc_272 N_A_27_297#_c_335_n N_VPWR_c_485_n 0.0027521f $X=6.095 $Y=1.88 $X2=0
+ $Y2=0
cc_273 N_A_27_297#_c_339_n N_VPWR_c_485_n 0.011801f $X=6.18 $Y=1.96 $X2=0 $Y2=0
cc_274 N_A_27_297#_M1001_d N_VPWR_c_484_n 0.00356385f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_275 N_A_27_297#_M1007_d N_VPWR_c_484_n 0.00231272f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_276 N_A_27_297#_M1018_d N_VPWR_c_484_n 0.00263241f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_277 N_A_27_297#_M1010_d N_VPWR_c_484_n 0.00293603f $X=3.355 $Y=1.485 $X2=0
+ $Y2=0
cc_278 N_A_27_297#_M1017_s N_VPWR_c_484_n 0.00307053f $X=4.635 $Y=1.485 $X2=0
+ $Y2=0
cc_279 N_A_27_297#_M1009_d N_VPWR_c_484_n 0.00391023f $X=6.035 $Y=1.485 $X2=0
+ $Y2=0
cc_280 N_A_27_297#_c_322_n N_VPWR_c_484_n 0.0268781f $X=1.115 $Y=2.38 $X2=0
+ $Y2=0
cc_281 N_A_27_297#_c_370_p N_VPWR_c_484_n 0.00654447f $X=0.345 $Y=2.38 $X2=0
+ $Y2=0
cc_282 N_A_27_297#_c_324_n N_VPWR_c_484_n 0.0334225f $X=2.055 $Y=2.38 $X2=0
+ $Y2=0
cc_283 N_A_27_297#_c_326_n N_VPWR_c_484_n 0.0140711f $X=3.415 $Y=1.88 $X2=0
+ $Y2=0
cc_284 N_A_27_297#_c_330_n N_VPWR_c_484_n 0.0122072f $X=4.695 $Y=1.88 $X2=0
+ $Y2=0
cc_285 N_A_27_297#_c_335_n N_VPWR_c_484_n 0.0149689f $X=6.095 $Y=1.88 $X2=0
+ $Y2=0
cc_286 N_A_27_297#_c_375_p N_VPWR_c_484_n 0.00654447f $X=1.2 $Y=2.38 $X2=0 $Y2=0
cc_287 N_A_27_297#_c_376_p N_VPWR_c_484_n 0.00646745f $X=3.5 $Y=1.96 $X2=0 $Y2=0
cc_288 N_A_27_297#_c_377_p N_VPWR_c_484_n 0.00646745f $X=4.78 $Y=1.96 $X2=0
+ $Y2=0
cc_289 N_A_27_297#_c_339_n N_VPWR_c_484_n 0.00646745f $X=6.18 $Y=1.96 $X2=0
+ $Y2=0
cc_290 N_A_27_297#_c_322_n N_VPWR_c_487_n 0.0415032f $X=1.115 $Y=2.38 $X2=0
+ $Y2=0
cc_291 N_A_27_297#_c_370_p N_VPWR_c_487_n 0.0119417f $X=0.345 $Y=2.38 $X2=0
+ $Y2=0
cc_292 N_A_27_297#_c_324_n N_VPWR_c_487_n 0.0534447f $X=2.055 $Y=2.38 $X2=0
+ $Y2=0
cc_293 N_A_27_297#_c_326_n N_VPWR_c_487_n 0.00242894f $X=3.415 $Y=1.88 $X2=0
+ $Y2=0
cc_294 N_A_27_297#_c_375_p N_VPWR_c_487_n 0.0119417f $X=1.2 $Y=2.38 $X2=0 $Y2=0
cc_295 N_A_27_297#_c_324_n N_VPWR_c_488_n 0.0122124f $X=2.055 $Y=2.38 $X2=0
+ $Y2=0
cc_296 N_A_27_297#_c_353_p N_VPWR_c_488_n 0.00249118f $X=2.14 $Y=2.295 $X2=0
+ $Y2=0
cc_297 N_A_27_297#_c_326_n N_VPWR_c_488_n 0.0299101f $X=3.415 $Y=1.88 $X2=0
+ $Y2=0
cc_298 N_A_27_297#_c_326_n N_VPWR_c_489_n 0.00218485f $X=3.415 $Y=1.88 $X2=0
+ $Y2=0
cc_299 N_A_27_297#_c_330_n N_VPWR_c_489_n 0.00136817f $X=4.695 $Y=1.88 $X2=0
+ $Y2=0
cc_300 N_A_27_297#_c_376_p N_VPWR_c_489_n 0.011801f $X=3.5 $Y=1.96 $X2=0 $Y2=0
cc_301 N_A_27_297#_c_330_n N_VPWR_c_490_n 0.0306127f $X=4.695 $Y=1.88 $X2=0
+ $Y2=0
cc_302 N_A_27_297#_c_376_p N_VPWR_c_490_n 0.0153798f $X=3.5 $Y=1.96 $X2=0 $Y2=0
cc_303 N_A_27_297#_c_377_p N_VPWR_c_490_n 0.016427f $X=4.78 $Y=1.96 $X2=0 $Y2=0
cc_304 N_A_27_297#_c_330_n N_VPWR_c_491_n 0.00117971f $X=4.695 $Y=1.88 $X2=0
+ $Y2=0
cc_305 N_A_27_297#_c_335_n N_VPWR_c_491_n 0.00233417f $X=6.095 $Y=1.88 $X2=0
+ $Y2=0
cc_306 N_A_27_297#_c_377_p N_VPWR_c_491_n 0.011801f $X=4.78 $Y=1.96 $X2=0 $Y2=0
cc_307 N_A_27_297#_c_335_n N_VPWR_c_492_n 0.0305174f $X=6.095 $Y=1.88 $X2=0
+ $Y2=0
cc_308 N_Y_M1001_s N_VPWR_c_484_n 0.00232895f $X=0.585 $Y=1.485 $X2=0 $Y2=0
cc_309 N_Y_M1013_s N_VPWR_c_484_n 0.00232895f $X=1.525 $Y=1.485 $X2=0 $Y2=0
cc_310 N_Y_c_397_n N_A_27_47#_M1015_s 0.00401694f $X=3.08 $Y=0.74 $X2=0 $Y2=0
cc_311 Y N_A_27_47#_M1015_s 0.00158476f $X=2.005 $Y=0.765 $X2=0 $Y2=0
cc_312 Y N_A_27_47#_M1015_s 0.00105541f $X=2.095 $Y=0.85 $X2=0 $Y2=0
cc_313 N_Y_c_399_n N_A_27_47#_c_570_n 0.00322894f $X=1.585 $Y=1.54 $X2=0 $Y2=0
cc_314 N_Y_c_399_n N_A_27_47#_c_568_n 8.51236e-19 $X=1.585 $Y=1.54 $X2=0 $Y2=0
cc_315 N_Y_M1004_d N_A_27_47#_c_569_n 0.00530193f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_316 N_Y_c_417_n N_A_27_47#_c_569_n 0.0241477f $X=1.965 $Y=0.74 $X2=0 $Y2=0
cc_317 N_Y_c_397_n N_A_27_47#_c_569_n 0.00698264f $X=3.08 $Y=0.74 $X2=0 $Y2=0
cc_318 Y N_A_27_47#_c_569_n 0.0118629f $X=2.005 $Y=0.765 $X2=0 $Y2=0
cc_319 N_Y_c_397_n N_VGND_c_613_n 0.00332968f $X=3.08 $Y=0.74 $X2=0 $Y2=0
cc_320 N_Y_M1004_d N_VGND_c_616_n 0.00300439f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_321 N_Y_M1011_s N_VGND_c_616_n 0.00219239f $X=2.945 $Y=0.235 $X2=0 $Y2=0
cc_322 N_Y_c_397_n N_VGND_c_616_n 0.0070144f $X=3.08 $Y=0.74 $X2=0 $Y2=0
cc_323 N_Y_c_397_n N_A_507_47#_M1011_d 0.00493096f $X=3.08 $Y=0.74 $X2=-0.195
+ $Y2=-0.24
cc_324 N_Y_M1011_s N_A_507_47#_c_677_n 0.00324009f $X=2.945 $Y=0.235 $X2=0 $Y2=0
cc_325 N_Y_c_397_n N_A_507_47#_c_677_n 0.0355575f $X=3.08 $Y=0.74 $X2=0 $Y2=0
cc_326 N_Y_c_397_n N_A_757_47#_c_696_n 0.00507639f $X=3.08 $Y=0.74 $X2=0 $Y2=0
cc_327 N_A_27_47#_c_570_n N_VGND_M1002_s 0.00443346f $X=1.035 $Y=0.8 $X2=-0.195
+ $Y2=-0.24
cc_328 N_A_27_47#_c_570_n N_VGND_c_610_n 0.0126475f $X=1.035 $Y=0.8 $X2=0 $Y2=0
cc_329 N_A_27_47#_c_577_n N_VGND_c_610_n 0.0109395f $X=1.16 $Y=0.465 $X2=0 $Y2=0
cc_330 N_A_27_47#_c_568_n N_VGND_c_610_n 0.00471242f $X=1.16 $Y=0.715 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_570_n N_VGND_c_613_n 0.00271675f $X=1.035 $Y=0.8 $X2=0 $Y2=0
cc_332 N_A_27_47#_c_577_n N_VGND_c_613_n 0.0120504f $X=1.16 $Y=0.465 $X2=0 $Y2=0
cc_333 N_A_27_47#_c_569_n N_VGND_c_613_n 0.0462122f $X=2.14 $Y=0.38 $X2=0 $Y2=0
cc_334 N_A_27_47#_c_566_n N_VGND_c_615_n 0.0172428f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_335 N_A_27_47#_c_570_n N_VGND_c_615_n 0.00259521f $X=1.035 $Y=0.8 $X2=0 $Y2=0
cc_336 N_A_27_47#_M1002_d N_VGND_c_616_n 0.00261174f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_M1014_d N_VGND_c_616_n 0.00217541f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_M1015_s N_VGND_c_616_n 0.00211652f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_566_n N_VGND_c_616_n 0.0123301f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_340 N_A_27_47#_c_570_n N_VGND_c_616_n 0.0109206f $X=1.035 $Y=0.8 $X2=0 $Y2=0
cc_341 N_A_27_47#_c_577_n N_VGND_c_616_n 0.00918694f $X=1.16 $Y=0.465 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_569_n N_VGND_c_616_n 0.035531f $X=2.14 $Y=0.38 $X2=0 $Y2=0
cc_343 N_A_27_47#_c_569_n N_A_507_47#_c_677_n 0.0145425f $X=2.14 $Y=0.38 $X2=0
+ $Y2=0
cc_344 N_VGND_c_616_n N_A_507_47#_M1011_d 0.00211652f $X=6.21 $Y=0 $X2=-0.195
+ $Y2=-0.24
cc_345 N_VGND_c_616_n N_A_507_47#_M1012_d 0.00217615f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_346 N_VGND_c_616_n N_A_507_47#_M1016_d 0.00211652f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_347 N_VGND_c_613_n N_A_507_47#_c_677_n 0.10687f $X=4.865 $Y=0 $X2=0 $Y2=0
cc_348 N_VGND_c_616_n N_A_507_47#_c_677_n 0.0736146f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_349 N_VGND_c_616_n N_A_757_47#_M1008_s 0.00259839f $X=6.21 $Y=0 $X2=-0.195
+ $Y2=-0.24
cc_350 N_VGND_c_616_n N_A_757_47#_M1006_s 0.00671736f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_351 N_VGND_M1006_d N_A_757_47#_c_696_n 0.0102367f $X=4.91 $Y=0.235 $X2=0
+ $Y2=0
cc_352 N_VGND_c_613_n N_A_757_47#_c_696_n 0.0341008f $X=4.865 $Y=0 $X2=0 $Y2=0
cc_353 N_VGND_c_614_n N_A_757_47#_c_696_n 0.00242734f $X=6.095 $Y=0 $X2=0 $Y2=0
cc_354 N_VGND_c_616_n N_A_757_47#_c_696_n 0.0150728f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_355 N_VGND_c_613_n N_A_757_47#_c_705_n 0.0150815f $X=4.865 $Y=0 $X2=0 $Y2=0
cc_356 N_VGND_c_614_n N_A_757_47#_c_705_n 0.0213183f $X=6.095 $Y=0 $X2=0 $Y2=0
cc_357 N_VGND_c_616_n N_A_757_47#_c_705_n 0.0139973f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_358 N_A_507_47#_c_677_n N_A_757_47#_M1008_s 0.00416045f $X=4.39 $Y=0.38
+ $X2=-0.195 $Y2=-0.24
cc_359 N_A_507_47#_M1016_d N_A_757_47#_c_696_n 0.0049097f $X=4.255 $Y=0.235
+ $X2=0 $Y2=0
cc_360 N_A_507_47#_c_677_n N_A_757_47#_c_696_n 0.0461069f $X=4.39 $Y=0.38 $X2=0
+ $Y2=0
