* File: sky130_fd_sc_hdll__or4b_2.pxi.spice
* Created: Wed Sep  2 08:49:42 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR4B_2%D_N N_D_N_c_75_n N_D_N_M1004_g N_D_N_M1010_g D_N
+ N_D_N_c_74_n PM_SKY130_FD_SC_HDLL__OR4B_2%D_N
x_PM_SKY130_FD_SC_HDLL__OR4B_2%A_186_21# N_A_186_21#_M1009_d N_A_186_21#_M1011_d
+ N_A_186_21#_M1003_d N_A_186_21#_c_100_n N_A_186_21#_M1001_g
+ N_A_186_21#_c_109_n N_A_186_21#_M1005_g N_A_186_21#_c_101_n
+ N_A_186_21#_M1013_g N_A_186_21#_c_110_n N_A_186_21#_M1012_g
+ N_A_186_21#_c_102_n N_A_186_21#_c_103_n N_A_186_21#_c_104_n
+ N_A_186_21#_c_105_n N_A_186_21#_c_106_n N_A_186_21#_c_107_n
+ N_A_186_21#_c_108_n N_A_186_21#_c_113_n N_A_186_21#_c_114_n
+ PM_SKY130_FD_SC_HDLL__OR4B_2%A_186_21#
x_PM_SKY130_FD_SC_HDLL__OR4B_2%A N_A_M1009_g N_A_c_219_n N_A_M1000_g A A
+ PM_SKY130_FD_SC_HDLL__OR4B_2%A
x_PM_SKY130_FD_SC_HDLL__OR4B_2%B N_B_M1007_g N_B_c_255_n N_B_M1008_g N_B_c_257_n
+ B B PM_SKY130_FD_SC_HDLL__OR4B_2%B
x_PM_SKY130_FD_SC_HDLL__OR4B_2%C N_C_M1011_g N_C_c_296_n N_C_M1006_g C C C
+ PM_SKY130_FD_SC_HDLL__OR4B_2%C
x_PM_SKY130_FD_SC_HDLL__OR4B_2%A_27_47# N_A_27_47#_M1010_s N_A_27_47#_M1004_s
+ N_A_27_47#_M1002_g N_A_27_47#_c_333_n N_A_27_47#_M1003_g N_A_27_47#_c_335_n
+ N_A_27_47#_c_328_n N_A_27_47#_c_336_n N_A_27_47#_c_329_n N_A_27_47#_c_330_n
+ N_A_27_47#_c_362_n N_A_27_47#_c_337_n N_A_27_47#_c_338_n N_A_27_47#_c_339_n
+ N_A_27_47#_c_340_n N_A_27_47#_c_331_n N_A_27_47#_c_342_n
+ PM_SKY130_FD_SC_HDLL__OR4B_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__OR4B_2%VPWR N_VPWR_M1004_d N_VPWR_M1012_d N_VPWR_c_440_n
+ N_VPWR_c_441_n VPWR N_VPWR_c_442_n N_VPWR_c_443_n N_VPWR_c_439_n
+ N_VPWR_c_445_n PM_SKY130_FD_SC_HDLL__OR4B_2%VPWR
x_PM_SKY130_FD_SC_HDLL__OR4B_2%X N_X_M1001_d N_X_M1005_s N_X_c_490_n N_X_c_499_n
+ N_X_c_501_n X PM_SKY130_FD_SC_HDLL__OR4B_2%X
x_PM_SKY130_FD_SC_HDLL__OR4B_2%VGND N_VGND_M1010_d N_VGND_M1013_s N_VGND_M1007_d
+ N_VGND_M1002_d N_VGND_c_523_n N_VGND_c_524_n N_VGND_c_525_n N_VGND_c_526_n
+ N_VGND_c_527_n N_VGND_c_528_n N_VGND_c_529_n VGND N_VGND_c_530_n
+ N_VGND_c_531_n N_VGND_c_532_n N_VGND_c_533_n VGND
+ PM_SKY130_FD_SC_HDLL__OR4B_2%VGND
cc_1 VNB N_D_N_M1010_g 0.0359501f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB D_N 0.00896472f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_D_N_c_74_n 0.040435f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_A_186_21#_c_100_n 0.0167914f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.202
cc_5 VNB N_A_186_21#_c_101_n 0.0172537f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_186_21#_c_102_n 0.0035936f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_186_21#_c_103_n 8.46298e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_186_21#_c_104_n 0.0143026f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_186_21#_c_105_n 9.56716e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_186_21#_c_106_n 0.0039387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_186_21#_c_107_n 0.0416341f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_186_21#_c_108_n 0.00155697f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_M1009_g 0.030306f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.695
cc_14 VNB N_A_c_219_n 0.0232575f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_15 VNB A 0.00582735f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_16 VNB N_B_M1007_g 0.0429934f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.695
cc_17 VNB N_C_M1011_g 0.0282187f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.695
cc_18 VNB N_C_c_296_n 0.0209354f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_19 VNB C 0.0276101f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_M1002_g 0.0621061f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_328_n 0.0171283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_329_n 0.00489827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_330_n 0.00968315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_331_n 0.00708948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_439_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_X_c_490_n 7.75412e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_27 VNB N_VGND_c_523_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_524_n 0.0175973f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_525_n 3.37329e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_526_n 0.0157371f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_527_n 0.0171871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_528_n 0.0142853f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_529_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_530_n 0.0148517f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_531_n 0.0236557f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_532_n 0.00642776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_533_n 0.224139f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VPB N_D_N_c_75_n 0.0227508f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_39 VPB D_N 0.00782582f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_40 VPB N_D_N_c_74_n 0.0162789f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_41 VPB N_A_186_21#_c_109_n 0.0187975f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_42 VPB N_A_186_21#_c_110_n 0.0186905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_186_21#_c_106_n 9.29639e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_186_21#_c_107_n 0.0221617f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_186_21#_c_113_n 0.0186879f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_186_21#_c_114_n 0.0110764f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_c_219_n 0.0279852f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_48 VPB N_B_M1007_g 9.70307e-19 $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.695
cc_49 VPB N_B_c_255_n 0.0480812f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_50 VPB N_B_M1008_g 0.0107369f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_51 VPB N_B_c_257_n 0.00653992f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.202
cc_52 VPB B 0.0148678f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_C_c_296_n 0.0253125f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_54 VPB N_A_27_47#_M1002_g 0.00153908f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_27_47#_c_333_n 0.0510487f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_56 VPB N_A_27_47#_M1003_g 0.0168697f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_57 VPB N_A_27_47#_c_335_n 0.00885218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_47#_c_336_n 0.0188451f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_47#_c_337_n 0.00810067f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_27_47#_c_338_n 0.0045818f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_27_47#_c_339_n 0.00228849f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_27_47#_c_340_n 0.00860011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_27_47#_c_331_n 0.00324685f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_27_47#_c_342_n 0.00264403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_440_n 0.0142662f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_66 VPB N_VPWR_c_441_n 0.0195535f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_67 VPB N_VPWR_c_442_n 0.0185074f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_443_n 0.0608312f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_439_n 0.0803247f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_445_n 0.018077f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_X_c_490_n 0.00114407f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_72 N_D_N_M1010_g N_A_186_21#_c_100_n 0.0155847f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_73 N_D_N_c_75_n N_A_186_21#_c_109_n 0.0177394f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_74 N_D_N_c_74_n N_A_186_21#_c_107_n 0.0155847f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_75 N_D_N_M1010_g N_A_27_47#_c_328_n 0.00422527f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_76 N_D_N_c_75_n N_A_27_47#_c_336_n 0.029625f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_77 D_N N_A_27_47#_c_336_n 0.0253129f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_78 N_D_N_c_74_n N_A_27_47#_c_336_n 0.00140343f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_79 N_D_N_M1010_g N_A_27_47#_c_329_n 0.0180619f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_80 D_N N_A_27_47#_c_329_n 0.00558788f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_81 N_D_N_c_74_n N_A_27_47#_c_329_n 0.00286467f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_82 D_N N_A_27_47#_c_330_n 0.0223758f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_83 N_D_N_c_74_n N_A_27_47#_c_330_n 0.00573424f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_84 N_D_N_c_75_n N_A_27_47#_c_331_n 0.00442551f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_85 N_D_N_M1010_g N_A_27_47#_c_331_n 0.00755038f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_86 D_N N_A_27_47#_c_331_n 0.0223143f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_87 N_D_N_c_75_n N_VPWR_c_442_n 0.00231735f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_88 N_D_N_c_75_n N_VPWR_c_439_n 0.00295025f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_89 N_D_N_c_75_n N_VPWR_c_445_n 3.77688e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_90 N_D_N_M1010_g X 5.80526e-19 $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_91 N_D_N_M1010_g N_VGND_c_523_n 0.00539494f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_92 N_D_N_M1010_g N_VGND_c_531_n 0.00439206f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_93 N_D_N_M1010_g N_VGND_c_533_n 0.00725985f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_94 N_A_186_21#_c_101_n N_A_M1009_g 0.019762f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_186_21#_c_102_n N_A_M1009_g 0.0128181f $X=2.185 $Y=0.785 $X2=0 $Y2=0
cc_96 N_A_186_21#_c_103_n N_A_M1009_g 0.00494164f $X=2.27 $Y=0.47 $X2=0 $Y2=0
cc_97 N_A_186_21#_c_106_n N_A_M1009_g 0.00357737f $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_186_21#_c_110_n N_A_c_219_n 0.021222f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A_186_21#_c_102_n N_A_c_219_n 0.00258294f $X=2.185 $Y=0.785 $X2=0 $Y2=0
cc_100 N_A_186_21#_c_106_n N_A_c_219_n 0.00337086f $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_186_21#_c_107_n N_A_c_219_n 0.0179781f $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A_186_21#_c_108_n N_A_c_219_n 0.00175462f $X=2.27 $Y=0.785 $X2=0 $Y2=0
cc_103 N_A_186_21#_c_114_n N_A_c_219_n 0.0159306f $X=3.525 $Y=1.612 $X2=0 $Y2=0
cc_104 N_A_186_21#_c_102_n A 0.0171267f $X=2.185 $Y=0.785 $X2=0 $Y2=0
cc_105 N_A_186_21#_c_104_n A 0.0105717f $X=3.135 $Y=0.785 $X2=0 $Y2=0
cc_106 N_A_186_21#_c_106_n A 0.0174525f $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_186_21#_c_107_n A 6.38059e-19 $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A_186_21#_c_108_n A 0.0123175f $X=2.27 $Y=0.785 $X2=0 $Y2=0
cc_109 N_A_186_21#_c_114_n A 0.0445983f $X=3.525 $Y=1.612 $X2=0 $Y2=0
cc_110 N_A_186_21#_c_103_n N_B_M1007_g 0.00490687f $X=2.27 $Y=0.47 $X2=0 $Y2=0
cc_111 N_A_186_21#_c_104_n N_B_M1007_g 0.0134671f $X=3.135 $Y=0.785 $X2=0 $Y2=0
cc_112 N_A_186_21#_c_114_n N_B_M1008_g 0.0131893f $X=3.525 $Y=1.612 $X2=0 $Y2=0
cc_113 N_A_186_21#_c_104_n N_B_c_257_n 8.69515e-19 $X=3.135 $Y=0.785 $X2=0 $Y2=0
cc_114 N_A_186_21#_c_110_n B 0.00489105f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A_186_21#_c_104_n N_C_M1011_g 0.0119333f $X=3.135 $Y=0.785 $X2=0 $Y2=0
cc_116 N_A_186_21#_c_105_n N_C_M1011_g 0.00493603f $X=3.22 $Y=0.47 $X2=0 $Y2=0
cc_117 N_A_186_21#_c_104_n N_C_c_296_n 0.00308437f $X=3.135 $Y=0.785 $X2=0 $Y2=0
cc_118 N_A_186_21#_c_113_n N_C_c_296_n 8.16039e-19 $X=3.74 $Y=1.655 $X2=0 $Y2=0
cc_119 N_A_186_21#_c_114_n N_C_c_296_n 0.0140358f $X=3.525 $Y=1.612 $X2=0 $Y2=0
cc_120 N_A_186_21#_c_104_n C 0.0333197f $X=3.135 $Y=0.785 $X2=0 $Y2=0
cc_121 N_A_186_21#_c_114_n C 0.082366f $X=3.525 $Y=1.612 $X2=0 $Y2=0
cc_122 N_A_186_21#_c_104_n N_A_27_47#_M1002_g 0.00527111f $X=3.135 $Y=0.785
+ $X2=0 $Y2=0
cc_123 N_A_186_21#_c_105_n N_A_27_47#_M1002_g 0.00338478f $X=3.22 $Y=0.47 $X2=0
+ $Y2=0
cc_124 N_A_186_21#_c_114_n N_A_27_47#_c_333_n 0.00127261f $X=3.525 $Y=1.612
+ $X2=0 $Y2=0
cc_125 N_A_186_21#_c_113_n N_A_27_47#_M1003_g 0.00811418f $X=3.74 $Y=1.655 $X2=0
+ $Y2=0
cc_126 N_A_186_21#_c_114_n N_A_27_47#_M1003_g 0.00848704f $X=3.525 $Y=1.612
+ $X2=0 $Y2=0
cc_127 N_A_186_21#_c_109_n N_A_27_47#_c_336_n 8.18622e-19 $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_128 N_A_186_21#_c_100_n N_A_27_47#_c_329_n 0.00143019f $X=1.005 $Y=0.995
+ $X2=0 $Y2=0
cc_129 N_A_186_21#_c_109_n N_A_27_47#_c_362_n 0.0159769f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_130 N_A_186_21#_c_110_n N_A_27_47#_c_362_n 0.0108558f $X=1.5 $Y=1.41 $X2=0
+ $Y2=0
cc_131 N_A_186_21#_c_106_n N_A_27_47#_c_362_n 0.00337526f $X=1.49 $Y=1.16 $X2=0
+ $Y2=0
cc_132 N_A_186_21#_c_107_n N_A_27_47#_c_362_n 8.57262e-19 $X=1.49 $Y=1.16 $X2=0
+ $Y2=0
cc_133 N_A_186_21#_c_114_n N_A_27_47#_c_337_n 0.0802533f $X=3.525 $Y=1.612 $X2=0
+ $Y2=0
cc_134 N_A_186_21#_c_113_n N_A_27_47#_c_340_n 0.00511705f $X=3.74 $Y=1.655 $X2=0
+ $Y2=0
cc_135 N_A_186_21#_c_114_n N_A_27_47#_c_340_n 0.00401454f $X=3.525 $Y=1.612
+ $X2=0 $Y2=0
cc_136 N_A_186_21#_c_100_n N_A_27_47#_c_331_n 0.00430733f $X=1.005 $Y=0.995
+ $X2=0 $Y2=0
cc_137 N_A_186_21#_c_109_n N_A_27_47#_c_331_n 0.00760096f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_138 N_A_186_21#_c_109_n N_A_27_47#_c_342_n 8.48942e-19 $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_139 N_A_186_21#_c_110_n N_A_27_47#_c_342_n 0.0125424f $X=1.5 $Y=1.41 $X2=0
+ $Y2=0
cc_140 N_A_186_21#_c_106_n N_A_27_47#_c_342_n 0.0115726f $X=1.49 $Y=1.16 $X2=0
+ $Y2=0
cc_141 N_A_186_21#_c_114_n N_A_27_47#_c_342_n 0.00998003f $X=3.525 $Y=1.612
+ $X2=0 $Y2=0
cc_142 N_A_186_21#_c_106_n N_VPWR_M1012_d 9.73829e-19 $X=1.49 $Y=1.16 $X2=0
+ $Y2=0
cc_143 N_A_186_21#_c_114_n N_VPWR_M1012_d 0.00160576f $X=3.525 $Y=1.612 $X2=0
+ $Y2=0
cc_144 N_A_186_21#_c_110_n N_VPWR_c_440_n 0.00774299f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_186_21#_c_109_n N_VPWR_c_441_n 0.00495396f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_146 N_A_186_21#_c_110_n N_VPWR_c_441_n 0.00496495f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_186_21#_c_109_n N_VPWR_c_439_n 0.00781284f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_148 N_A_186_21#_c_110_n N_VPWR_c_439_n 0.00778764f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_186_21#_c_109_n N_VPWR_c_445_n 0.00772305f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_150 N_A_186_21#_c_100_n N_X_c_490_n 0.00443195f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_186_21#_c_109_n N_X_c_490_n 0.00222567f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_186_21#_c_101_n N_X_c_490_n 0.00157178f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_186_21#_c_110_n N_X_c_490_n 5.7361e-19 $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_186_21#_c_106_n N_X_c_490_n 0.0417298f $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_186_21#_c_107_n N_X_c_490_n 0.0200289f $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_186_21#_c_100_n N_X_c_499_n 0.00404212f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A_186_21#_c_107_n N_X_c_499_n 0.00309179f $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A_186_21#_c_109_n N_X_c_501_n 0.00723721f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_186_21#_c_106_n N_X_c_501_n 0.0098555f $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_186_21#_c_107_n N_X_c_501_n 0.0053503f $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A_186_21#_c_100_n X 0.00631372f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_186_21#_c_114_n A_425_297# 0.0023755f $X=3.525 $Y=1.612 $X2=-0.19
+ $Y2=-0.24
cc_163 N_A_186_21#_c_114_n A_531_297# 0.00134267f $X=3.525 $Y=1.612 $X2=-0.19
+ $Y2=-0.24
cc_164 N_A_186_21#_c_114_n A_615_297# 0.00250556f $X=3.525 $Y=1.612 $X2=-0.19
+ $Y2=-0.24
cc_165 N_A_186_21#_c_102_n N_VGND_M1013_s 0.00379245f $X=2.185 $Y=0.785 $X2=0
+ $Y2=0
cc_166 N_A_186_21#_c_106_n N_VGND_M1013_s 0.0020976f $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_186_21#_c_100_n N_VGND_c_523_n 0.00385938f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_168 N_A_186_21#_c_100_n N_VGND_c_524_n 0.00496228f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_169 N_A_186_21#_c_101_n N_VGND_c_524_n 0.00526846f $X=1.475 $Y=0.995 $X2=0
+ $Y2=0
cc_170 N_A_186_21#_c_103_n N_VGND_c_525_n 0.0125809f $X=2.27 $Y=0.47 $X2=0 $Y2=0
cc_171 N_A_186_21#_c_104_n N_VGND_c_525_n 0.0165174f $X=3.135 $Y=0.785 $X2=0
+ $Y2=0
cc_172 N_A_186_21#_c_105_n N_VGND_c_525_n 0.0130167f $X=3.22 $Y=0.47 $X2=0 $Y2=0
cc_173 N_A_186_21#_c_105_n N_VGND_c_527_n 0.0192809f $X=3.22 $Y=0.47 $X2=0 $Y2=0
cc_174 N_A_186_21#_c_102_n N_VGND_c_528_n 0.00328839f $X=2.185 $Y=0.785 $X2=0
+ $Y2=0
cc_175 N_A_186_21#_c_103_n N_VGND_c_528_n 0.010678f $X=2.27 $Y=0.47 $X2=0 $Y2=0
cc_176 N_A_186_21#_c_104_n N_VGND_c_528_n 0.00344013f $X=3.135 $Y=0.785 $X2=0
+ $Y2=0
cc_177 N_A_186_21#_c_104_n N_VGND_c_530_n 0.00328013f $X=3.135 $Y=0.785 $X2=0
+ $Y2=0
cc_178 N_A_186_21#_c_105_n N_VGND_c_530_n 0.010678f $X=3.22 $Y=0.47 $X2=0 $Y2=0
cc_179 N_A_186_21#_c_100_n N_VGND_c_532_n 0.00116825f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_180 N_A_186_21#_c_101_n N_VGND_c_532_n 0.0116888f $X=1.475 $Y=0.995 $X2=0
+ $Y2=0
cc_181 N_A_186_21#_c_102_n N_VGND_c_532_n 0.0122657f $X=2.185 $Y=0.785 $X2=0
+ $Y2=0
cc_182 N_A_186_21#_c_103_n N_VGND_c_532_n 0.013288f $X=2.27 $Y=0.47 $X2=0 $Y2=0
cc_183 N_A_186_21#_c_106_n N_VGND_c_532_n 0.00974716f $X=1.49 $Y=1.16 $X2=0
+ $Y2=0
cc_184 N_A_186_21#_c_107_n N_VGND_c_532_n 3.46465e-19 $X=1.49 $Y=1.16 $X2=0
+ $Y2=0
cc_185 N_A_186_21#_M1009_d N_VGND_c_533_n 0.00400479f $X=2.085 $Y=0.235 $X2=0
+ $Y2=0
cc_186 N_A_186_21#_M1011_d N_VGND_c_533_n 0.00693283f $X=3.035 $Y=0.235 $X2=0
+ $Y2=0
cc_187 N_A_186_21#_c_100_n N_VGND_c_533_n 0.0088172f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_188 N_A_186_21#_c_101_n N_VGND_c_533_n 0.00902097f $X=1.475 $Y=0.995 $X2=0
+ $Y2=0
cc_189 N_A_186_21#_c_102_n N_VGND_c_533_n 0.00634556f $X=2.185 $Y=0.785 $X2=0
+ $Y2=0
cc_190 N_A_186_21#_c_103_n N_VGND_c_533_n 0.00640162f $X=2.27 $Y=0.47 $X2=0
+ $Y2=0
cc_191 N_A_186_21#_c_104_n N_VGND_c_533_n 0.0123938f $X=3.135 $Y=0.785 $X2=0
+ $Y2=0
cc_192 N_A_186_21#_c_105_n N_VGND_c_533_n 0.00640162f $X=3.22 $Y=0.47 $X2=0
+ $Y2=0
cc_193 N_A_186_21#_c_106_n N_VGND_c_533_n 8.61174e-19 $X=1.49 $Y=1.16 $X2=0
+ $Y2=0
cc_194 N_A_M1009_g N_B_M1007_g 0.0166634f $X=2.01 $Y=0.445 $X2=0 $Y2=0
cc_195 N_A_c_219_n N_B_M1007_g 0.0219951f $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_196 A N_B_M1007_g 0.00623202f $X=2.185 $Y=1.105 $X2=0 $Y2=0
cc_197 N_A_c_219_n N_B_M1008_g 0.0232186f $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_c_219_n N_B_c_257_n 0.0038729f $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_199 A C 0.0120461f $X=2.185 $Y=1.105 $X2=0 $Y2=0
cc_200 N_A_c_219_n N_A_27_47#_c_337_n 0.0121855f $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A_c_219_n N_A_27_47#_c_342_n 0.00254462f $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A_c_219_n N_VPWR_c_440_n 4.84843e-19 $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A_c_219_n N_VPWR_c_443_n 0.00349789f $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A_c_219_n N_VPWR_c_439_n 0.00448105f $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A_M1009_g N_VGND_c_525_n 5.82695e-19 $X=2.01 $Y=0.445 $X2=0 $Y2=0
cc_206 N_A_M1009_g N_VGND_c_528_n 0.00347531f $X=2.01 $Y=0.445 $X2=0 $Y2=0
cc_207 N_A_M1009_g N_VGND_c_532_n 0.00802887f $X=2.01 $Y=0.445 $X2=0 $Y2=0
cc_208 N_A_M1009_g N_VGND_c_533_n 0.00439991f $X=2.01 $Y=0.445 $X2=0 $Y2=0
cc_209 N_B_M1007_g N_C_M1011_g 0.0410744f $X=2.54 $Y=0.445 $X2=0 $Y2=0
cc_210 N_B_M1008_g N_C_c_296_n 0.0353329f $X=2.565 $Y=1.695 $X2=0 $Y2=0
cc_211 N_B_c_257_n N_C_c_296_n 0.00536912f $X=2.56 $Y=1.41 $X2=0 $Y2=0
cc_212 B N_C_c_296_n 7.32077e-19 $X=2.785 $Y=2.305 $X2=0 $Y2=0
cc_213 N_B_M1007_g C 0.00154316f $X=2.54 $Y=0.445 $X2=0 $Y2=0
cc_214 N_B_c_255_n N_A_27_47#_c_333_n 0.00395002f $X=2.565 $Y=2.035 $X2=0 $Y2=0
cc_215 B N_A_27_47#_c_333_n 0.0016216f $X=2.785 $Y=2.305 $X2=0 $Y2=0
cc_216 N_B_c_255_n N_A_27_47#_c_337_n 0.00133343f $X=2.565 $Y=2.035 $X2=0 $Y2=0
cc_217 N_B_M1008_g N_A_27_47#_c_337_n 0.0118247f $X=2.565 $Y=1.695 $X2=0 $Y2=0
cc_218 B N_A_27_47#_c_337_n 0.054362f $X=2.785 $Y=2.305 $X2=0 $Y2=0
cc_219 N_B_c_255_n N_A_27_47#_c_338_n 0.00256058f $X=2.565 $Y=2.035 $X2=0 $Y2=0
cc_220 B N_A_27_47#_c_338_n 0.00587192f $X=2.785 $Y=2.305 $X2=0 $Y2=0
cc_221 N_B_c_255_n N_A_27_47#_c_339_n 4.83868e-19 $X=2.565 $Y=2.035 $X2=0 $Y2=0
cc_222 B N_A_27_47#_c_339_n 0.0122703f $X=2.785 $Y=2.305 $X2=0 $Y2=0
cc_223 N_B_c_255_n N_A_27_47#_c_342_n 0.00238089f $X=2.565 $Y=2.035 $X2=0 $Y2=0
cc_224 B N_A_27_47#_c_342_n 0.00221937f $X=2.785 $Y=2.305 $X2=0 $Y2=0
cc_225 N_B_c_255_n N_VPWR_c_440_n 0.00112818f $X=2.565 $Y=2.035 $X2=0 $Y2=0
cc_226 B N_VPWR_c_440_n 0.00583495f $X=2.785 $Y=2.305 $X2=0 $Y2=0
cc_227 N_B_c_255_n N_VPWR_c_443_n 0.00813358f $X=2.565 $Y=2.035 $X2=0 $Y2=0
cc_228 B N_VPWR_c_443_n 0.0364283f $X=2.785 $Y=2.305 $X2=0 $Y2=0
cc_229 N_B_c_255_n N_VPWR_c_439_n 0.0115323f $X=2.565 $Y=2.035 $X2=0 $Y2=0
cc_230 B N_VPWR_c_439_n 0.0266655f $X=2.785 $Y=2.305 $X2=0 $Y2=0
cc_231 N_B_M1007_g N_VGND_c_525_n 0.00761566f $X=2.54 $Y=0.445 $X2=0 $Y2=0
cc_232 N_B_M1007_g N_VGND_c_528_n 0.0034676f $X=2.54 $Y=0.445 $X2=0 $Y2=0
cc_233 N_B_M1007_g N_VGND_c_532_n 5.85038e-19 $X=2.54 $Y=0.445 $X2=0 $Y2=0
cc_234 N_B_M1007_g N_VGND_c_533_n 0.00439987f $X=2.54 $Y=0.445 $X2=0 $Y2=0
cc_235 N_C_M1011_g N_A_27_47#_M1002_g 0.0165487f $X=2.96 $Y=0.445 $X2=0 $Y2=0
cc_236 N_C_c_296_n N_A_27_47#_M1002_g 0.0180491f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_237 C N_A_27_47#_M1002_g 0.0171899f $X=3.715 $Y=1.105 $X2=0 $Y2=0
cc_238 N_C_c_296_n N_A_27_47#_M1003_g 0.021451f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_239 N_C_c_296_n N_A_27_47#_c_335_n 0.00398214f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_240 C N_A_27_47#_c_335_n 0.00121851f $X=3.715 $Y=1.105 $X2=0 $Y2=0
cc_241 N_C_c_296_n N_A_27_47#_c_337_n 0.0120264f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_242 N_C_c_296_n N_A_27_47#_c_338_n 0.00189355f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_243 N_C_c_296_n N_VPWR_c_443_n 0.00340707f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_244 N_C_c_296_n N_VPWR_c_439_n 0.00431405f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_245 N_C_M1011_g N_VGND_c_525_n 0.00753553f $X=2.96 $Y=0.445 $X2=0 $Y2=0
cc_246 N_C_M1011_g N_VGND_c_527_n 6.1514e-19 $X=2.96 $Y=0.445 $X2=0 $Y2=0
cc_247 C N_VGND_c_527_n 0.0132765f $X=3.715 $Y=1.105 $X2=0 $Y2=0
cc_248 N_C_M1011_g N_VGND_c_530_n 0.0034676f $X=2.96 $Y=0.445 $X2=0 $Y2=0
cc_249 N_C_M1011_g N_VGND_c_533_n 0.00437864f $X=2.96 $Y=0.445 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_336_n N_VPWR_M1004_d 0.00653872f $X=0.51 $Y=1.747 $X2=-0.19
+ $Y2=-0.24
cc_251 N_A_27_47#_c_362_n N_VPWR_M1004_d 0.00375559f $X=1.54 $Y=2.08 $X2=-0.19
+ $Y2=-0.24
cc_252 N_A_27_47#_c_331_n N_VPWR_M1004_d 0.00267665f $X=0.662 $Y=1.605 $X2=-0.19
+ $Y2=-0.24
cc_253 N_A_27_47#_c_337_n N_VPWR_M1012_d 5.43066e-19 $X=3.16 $Y=1.87 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_342_n N_VPWR_M1012_d 0.00497025f $X=1.702 $Y=1.87 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_337_n N_VPWR_c_440_n 0.00383286f $X=3.16 $Y=1.87 $X2=0 $Y2=0
cc_256 N_A_27_47#_c_342_n N_VPWR_c_440_n 0.0170862f $X=1.702 $Y=1.87 $X2=0 $Y2=0
cc_257 N_A_27_47#_c_362_n N_VPWR_c_441_n 0.011801f $X=1.54 $Y=2.08 $X2=0 $Y2=0
cc_258 N_A_27_47#_c_342_n N_VPWR_c_441_n 0.00151337f $X=1.702 $Y=1.87 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_333_n N_VPWR_c_443_n 0.00790512f $X=3.505 $Y=2.035 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_339_n N_VPWR_c_443_n 0.00780423f $X=3.33 $Y=2.3 $X2=0 $Y2=0
cc_261 N_A_27_47#_c_340_n N_VPWR_c_443_n 0.0149599f $X=3.44 $Y=2.3 $X2=0 $Y2=0
cc_262 N_A_27_47#_c_333_n N_VPWR_c_439_n 0.0110773f $X=3.505 $Y=2.035 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_c_336_n N_VPWR_c_439_n 0.0169864f $X=0.51 $Y=1.747 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_362_n N_VPWR_c_439_n 0.0182974f $X=1.54 $Y=2.08 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_337_n N_VPWR_c_439_n 0.0174073f $X=3.16 $Y=1.87 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_339_n N_VPWR_c_439_n 0.0061985f $X=3.33 $Y=2.3 $X2=0 $Y2=0
cc_267 N_A_27_47#_c_340_n N_VPWR_c_439_n 0.0127153f $X=3.44 $Y=2.3 $X2=0 $Y2=0
cc_268 N_A_27_47#_c_342_n N_VPWR_c_439_n 0.00381682f $X=1.702 $Y=1.87 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_336_n N_VPWR_c_445_n 0.0245412f $X=0.51 $Y=1.747 $X2=0 $Y2=0
cc_270 N_A_27_47#_c_362_n N_VPWR_c_445_n 0.00504782f $X=1.54 $Y=2.08 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_362_n N_X_M1005_s 0.00449183f $X=1.54 $Y=2.08 $X2=0 $Y2=0
cc_272 N_A_27_47#_c_331_n N_X_c_490_n 0.0372026f $X=0.662 $Y=1.605 $X2=0 $Y2=0
cc_273 N_A_27_47#_c_329_n N_X_c_499_n 0.0119177f $X=0.645 $Y=0.82 $X2=0 $Y2=0
cc_274 N_A_27_47#_c_362_n N_X_c_501_n 0.0202872f $X=1.54 $Y=2.08 $X2=0 $Y2=0
cc_275 N_A_27_47#_c_331_n N_X_c_501_n 0.0216559f $X=0.662 $Y=1.605 $X2=0 $Y2=0
cc_276 N_A_27_47#_c_342_n N_X_c_501_n 0.00278809f $X=1.702 $Y=1.87 $X2=0 $Y2=0
cc_277 N_A_27_47#_c_328_n X 0.00443712f $X=0.26 $Y=0.5 $X2=0 $Y2=0
cc_278 N_A_27_47#_c_337_n A_425_297# 0.00241926f $X=3.16 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_279 N_A_27_47#_c_337_n A_531_297# 0.00134267f $X=3.16 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_280 N_A_27_47#_c_337_n A_615_297# 0.00412715f $X=3.16 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_281 N_A_27_47#_c_329_n N_VGND_M1010_d 0.00336683f $X=0.645 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_282 N_A_27_47#_c_328_n N_VGND_c_523_n 0.0110639f $X=0.26 $Y=0.5 $X2=0 $Y2=0
cc_283 N_A_27_47#_c_329_n N_VGND_c_523_n 0.0116177f $X=0.645 $Y=0.82 $X2=0 $Y2=0
cc_284 N_A_27_47#_M1002_g N_VGND_c_525_n 5.83747e-19 $X=3.48 $Y=0.445 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_M1002_g N_VGND_c_527_n 0.0117016f $X=3.48 $Y=0.445 $X2=0 $Y2=0
cc_286 N_A_27_47#_M1002_g N_VGND_c_530_n 0.0046653f $X=3.48 $Y=0.445 $X2=0 $Y2=0
cc_287 N_A_27_47#_c_328_n N_VGND_c_531_n 0.0126415f $X=0.26 $Y=0.5 $X2=0 $Y2=0
cc_288 N_A_27_47#_c_329_n N_VGND_c_531_n 0.00468693f $X=0.645 $Y=0.82 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_M1010_s N_VGND_c_533_n 0.00303542f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_M1002_g N_VGND_c_533_n 0.00823078f $X=3.48 $Y=0.445 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_328_n N_VGND_c_533_n 0.00971608f $X=0.26 $Y=0.5 $X2=0 $Y2=0
cc_292 N_A_27_47#_c_329_n N_VGND_c_533_n 0.00853072f $X=0.645 $Y=0.82 $X2=0
+ $Y2=0
cc_293 N_VPWR_c_439_n N_X_M1005_s 0.00306279f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_294 X N_VGND_c_523_n 0.0225201f $X=1.17 $Y=0.425 $X2=0 $Y2=0
cc_295 X N_VGND_c_524_n 0.0199697f $X=1.17 $Y=0.425 $X2=0 $Y2=0
cc_296 N_X_M1001_d N_VGND_c_533_n 0.00434153f $X=1.08 $Y=0.235 $X2=0 $Y2=0
cc_297 X N_VGND_c_533_n 0.0123029f $X=1.17 $Y=0.425 $X2=0 $Y2=0
