* File: sky130_fd_sc_hdll__a21oi_4.spice
* Created: Thu Aug 27 18:53:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a21oi_4.pex.spice"
.subckt sky130_fd_sc_hdll__a21oi_4  VNB VPB B1 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_B1_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.1235 PD=1.83 PS=1.03 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75000.2
+ SB=75005.6 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_B1_M1003_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.1235 PD=0.98 PS=1.03 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75000.7
+ SB=75005 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1003_d N_B1_M1010_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_B1_M1013_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.10725 PD=0.97 PS=0.98 NRD=7.38 NRS=9.228 M=1 R=4.33333 SA=75001.7
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1005 N_A_502_47#_M1005_d N_A2_M1005_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.104 PD=0.98 PS=0.97 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1015 N_Y_M1015_d N_A1_M1015_g N_A_502_47#_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75002.6
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1016 N_Y_M1015_d N_A1_M1016_g N_A_502_47#_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75003.1
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1019 N_Y_M1019_d N_A1_M1019_g N_A_502_47#_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.10725 PD=1.03 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75003.6
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1023 N_Y_M1019_d N_A1_M1023_g N_A_502_47#_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.091 PD=1.03 PS=0.93 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75004.1
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1008 N_A_502_47#_M1023_s N_A2_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.10725 PD=0.93 PS=0.98 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75004.5
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1011 N_A_502_47#_M1011_d N_A2_M1011_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75005
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1014 N_A_502_47#_M1011_d N_A2_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.20475 PD=0.98 PS=1.93 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75005.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1006_d N_B1_M1006_g N_A_28_297#_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.27 PD=1.3 PS=2.54 NRD=1.9503 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90005.5 A=0.18 P=2.36 MULT=1
MM1009 N_Y_M1006_d N_B1_M1009_g N_A_28_297#_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90005 A=0.18 P=2.36 MULT=1
MM1017 N_Y_M1017_d N_B1_M1017_g N_A_28_297#_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.1
+ SB=90004.5 A=0.18 P=2.36 MULT=1
MM1020 N_Y_M1017_d N_B1_M1020_g N_A_28_297#_M1020_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.165 PD=1.3 PS=1.33 NRD=1.9503 NRS=7.8603 M=1 R=5.55556 SA=90001.6
+ SB=90004.1 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A2_M1002_g N_A_28_297#_M1020_s VPB PHIGHVT L=0.18 W=1
+ AD=0.155 AS=0.165 PD=1.31 PS=1.33 NRD=3.9203 NRS=1.9503 M=1 R=5.55556
+ SA=90002.1 SB=90003.6 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1002_d N_A1_M1000_g N_A_28_297#_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.155 AS=0.15 PD=1.31 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.6
+ SB=90003.1 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g N_A_28_297#_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90003.1
+ SB=90002.6 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1004_d N_A1_M1007_g N_A_28_297#_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90003.6
+ SB=90002.1 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_A1_M1012_g N_A_28_297#_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90004.1
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1012_d N_A2_M1018_g N_A_28_297#_M1018_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90004.5
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1021 N_VPWR_M1021_d N_A2_M1021_g N_A_28_297#_M1018_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90005
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1022 N_VPWR_M1021_d N_A2_M1022_g N_A_28_297#_M1022_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90005.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX24_noxref VNB VPB NWDIODE A=10.9461 P=16.85
pX25_noxref noxref_11 A2 A2 PROBETYPE=1
c_43 VNB 0 1.1531e-19 $X=0.15 $Y=-0.085
c_79 VPB 0 3.14505e-20 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__a21oi_4.pxi.spice"
*
.ends
*
*
