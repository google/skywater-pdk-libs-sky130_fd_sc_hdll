* NGSPICE file created from sky130_fd_sc_hdll__o21ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 a_29_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=8.7425e+11p pd=7.89e+06u as=5.005e+11p ps=4.14e+06u
M1001 Y B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6e+11p pd=5.2e+06u as=9.95e+11p ps=7.99e+06u
M1002 a_120_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6.7e+11p pd=5.34e+06u as=0p ps=0u
M1003 a_120_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y B1 a_29_47# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=0p ps=0u
M1005 VPWR A1 a_120_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_29_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A2 a_120_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A1 a_29_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_29_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A2 a_29_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

