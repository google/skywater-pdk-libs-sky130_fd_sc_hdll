* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__clkbuf_2 A VGND VNB VPB VPWR X
M1000 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=2.457e+11p pd=2.85e+06u as=1.323e+11p ps=1.47e+06u
M1001 VGND a_27_47# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.554e+11p ps=1.58e+06u
M1002 VPWR A a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=6.15e+11p pd=5.23e+06u as=2.75e+11p ps=2.55e+06u
M1003 X a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1005 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
