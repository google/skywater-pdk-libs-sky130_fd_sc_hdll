* File: sky130_fd_sc_hdll__sdfstp_4.spice
* Created: Wed Sep  2 08:51:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__sdfstp_4.pex.spice"
.subckt sky130_fd_sc_hdll__sdfstp_4  VNB VPB SCD SCE D CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* SCE	SCE
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1027 A_119_47# N_SCD_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.42 AD=0.0546
+ AS=0.1302 PD=0.68 PS=1.46 NRD=21.42 NRS=12.852 M=1 R=2.8 SA=75000.2 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1037 N_A_201_47#_M1037_d N_SCE_M1037_g A_119_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0546 PD=0.74 PS=0.68 NRD=0 NRS=21.42 M=1 R=2.8 SA=75000.6
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1035 A_295_47# N_D_M1035_g N_A_201_47#_M1037_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0672 PD=0.69 PS=0.74 NRD=22.848 NRS=12.852 M=1 R=2.8 SA=75001.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_349_21#_M1001_g A_295_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1428 AS=0.0567 PD=1.52 PS=0.69 NRD=21.42 NRS=22.848 M=1 R=2.8 SA=75001.5
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_SCE_M1007_g N_A_349_21#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1302 PD=1.36 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_CLK_M1021_g N_A_693_369#_M1021_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1018 N_A_877_369#_M1018_d N_A_693_369#_M1018_g N_VGND_M1021_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1092 AS=0.0672 PD=1.36 PS=0.74 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1033 N_A_1075_413#_M1033_d N_A_693_369#_M1033_g N_A_201_47#_M1033_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1028 A_1177_47# N_A_877_369#_M1028_g N_A_1075_413#_M1033_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0546 AS=0.0672 PD=0.68 PS=0.74 NRD=21.42 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_1229_21#_M1019_g A_1177_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0546 PD=1.36 PS=0.68 NRD=0 NRS=21.42 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1024 A_1467_47# N_A_1075_413#_M1024_g N_A_1229_21#_M1024_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0546 AS=0.1512 PD=0.68 PS=1.56 NRD=21.42 NRS=27.132 M=1 R=2.8
+ SA=75000.3 SB=75004.6 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_SET_B_M1017_g A_1467_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0885566 AS=0.0546 PD=0.80434 PS=0.68 NRD=1.428 NRS=21.42 M=1 R=2.8
+ SA=75000.7 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1023 A_1654_47# N_A_1075_413#_M1023_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.64
+ AD=0.2544 AS=0.134943 PD=1.435 PS=1.22566 NRD=64.212 NRS=16.872 M=1 R=4.26667
+ SA=75000.9 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1045 N_A_1745_329#_M1045_d N_A_877_369#_M1045_g A_1654_47# VNB NSHORT L=0.15
+ W=0.64 AD=0.201177 AS=0.2544 PD=1.50943 PS=1.435 NRD=14.052 NRS=64.212 M=1
+ R=4.26667 SA=75001.8 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1005 A_1995_47# N_A_693_369#_M1005_g N_A_1745_329#_M1045_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.132023 PD=0.63 PS=0.990566 NRD=14.28 NRS=72.852 M=1
+ R=2.8 SA=75002.9 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1002 A_2067_47# N_A_1951_295#_M1002_g A_1995_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1008 AS=0.0441 PD=0.9 PS=0.63 NRD=52.848 NRS=14.28 M=1 R=2.8 SA=75003.3
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_SET_B_M1015_g A_2067_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0987 AS=0.1008 PD=0.89 PS=0.9 NRD=41.424 NRS=52.848 M=1 R=2.8 SA=75003.9
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1022 N_A_1951_295#_M1022_d N_A_1745_329#_M1022_g N_VGND_M1015_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1596 AS=0.0987 PD=1.6 PS=0.89 NRD=32.856 NRS=12.852 M=1
+ R=2.8 SA=75004.5 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1030 N_VGND_M1030_d N_A_1745_329#_M1030_g N_A_2447_47#_M1030_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.121875 AS=0.2015 PD=1.025 PS=1.92 NRD=3.684 NRS=8.304 M=1
+ R=4.33333 SA=75000.2 SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1030_d N_A_2447_47#_M1009_g N_Q_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.121875 AS=0.104 PD=1.025 PS=0.97 NRD=13.836 NRS=0 M=1 R=4.33333
+ SA=75000.8 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_A_2447_47#_M1013_g N_Q_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=8.304 M=1 R=4.33333
+ SA=75001.2 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1036 N_VGND_M1013_d N_A_2447_47#_M1036_g N_Q_M1036_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1038 N_VGND_M1038_d N_A_2447_47#_M1038_g N_Q_M1036_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=8.304 M=1 R=4.33333
+ SA=75002.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_VPWR_M1010_d N_SCD_M1010_g N_A_27_369#_M1010_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90001.5 A=0.1152 P=1.64 MULT=1
MM1039 A_211_369# N_SCE_M1039_g N_VPWR_M1010_d VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0736 AS=0.0928 PD=0.87 PS=0.93 NRD=18.4589 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90001.1 A=0.1152 P=1.64 MULT=1
MM1041 N_A_201_47#_M1041_d N_D_M1041_g A_211_369# VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.0736 PD=0.93 PS=0.87 NRD=1.5366 NRS=18.4589 M=1 R=3.55556
+ SA=90001.1 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1026 N_A_27_369#_M1026_d N_A_349_21#_M1026_g N_A_201_47#_M1041_d VPB PHIGHVT
+ L=0.18 W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1
+ R=3.55556 SA=90001.5 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1014 N_VPWR_M1014_d N_SCE_M1014_g N_A_349_21#_M1014_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.1728 PD=1.82 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1044 N_VPWR_M1044_d N_CLK_M1044_g N_A_693_369#_M1044_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1031 N_A_877_369#_M1031_d N_A_693_369#_M1031_g N_VPWR_M1044_d VPB PHIGHVT
+ L=0.18 W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1
+ R=3.55556 SA=90000.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1008 N_A_1075_413#_M1008_d N_A_877_369#_M1008_g N_A_201_47#_M1008_s VPB
+ PHIGHVT L=0.18 W=0.42 AD=0.0609 AS=0.1134 PD=0.71 PS=1.38 NRD=2.3443
+ NRS=2.3443 M=1 R=2.33333 SA=90000.2 SB=90005.5 A=0.0756 P=1.2 MULT=1
MM1042 A_1169_413# N_A_693_369#_M1042_g N_A_1075_413#_M1008_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0798 AS=0.0609 PD=0.8 PS=0.71 NRD=63.3158 NRS=2.3443 M=1 R=2.33333
+ SA=90000.6 SB=90005 A=0.0756 P=1.2 MULT=1
MM1043 N_VPWR_M1043_d N_A_1229_21#_M1043_g A_1169_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.1071 AS=0.0798 PD=0.93 PS=0.8 NRD=30.4759 NRS=63.3158 M=1 R=2.33333
+ SA=90001.2 SB=90004.5 A=0.0756 P=1.2 MULT=1
MM1011 N_A_1229_21#_M1011_d N_A_1075_413#_M1011_g N_VPWR_M1043_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.0861 AS=0.1071 PD=0.83 PS=0.93 NRD=14.0658 NRS=77.3816 M=1
+ R=2.33333 SA=90001.9 SB=90003.8 A=0.0756 P=1.2 MULT=1
MM1000 N_VPWR_M1000_d N_SET_B_M1000_g N_A_1229_21#_M1011_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0994 AS=0.0861 PD=0.86 PS=0.83 NRD=23.443 NRS=46.886 M=1 R=2.33333
+ SA=90002.5 SB=90003.2 A=0.0756 P=1.2 MULT=1
MM1032 A_1663_329# N_A_1075_413#_M1032_g N_VPWR_M1000_d VPB PHIGHVT L=0.18
+ W=0.84 AD=0.0966 AS=0.1988 PD=1.07 PS=1.72 NRD=14.0658 NRS=28.1316 M=1
+ R=4.66667 SA=90001.6 SB=90001.6 A=0.1512 P=2.04 MULT=1
MM1034 N_A_1745_329#_M1034_d N_A_693_369#_M1034_g A_1663_329# VPB PHIGHVT L=0.18
+ W=0.84 AD=0.2268 AS=0.0966 PD=1.85333 PS=1.07 NRD=36.3465 NRS=14.0658 M=1
+ R=4.66667 SA=90002.1 SB=90001.2 A=0.1512 P=2.04 MULT=1
MM1006 A_1891_413# N_A_877_369#_M1006_g N_A_1745_329#_M1034_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0651 AS=0.1134 PD=0.73 PS=0.926667 NRD=46.886 NRS=53.9386 M=1
+ R=2.33333 SA=90004.3 SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1020 N_VPWR_M1020_d N_A_1951_295#_M1020_g A_1891_413# VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1113 AS=0.0651 PD=0.95 PS=0.73 NRD=65.6601 NRS=46.886 M=1
+ R=2.33333 SA=90004.7 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1003 N_A_1745_329#_M1003_d N_SET_B_M1003_g N_VPWR_M1020_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1344 AS=0.1113 PD=1.48 PS=0.95 NRD=2.3443 NRS=51.5943 M=1
+ R=2.33333 SA=90005.5 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1004 N_A_1951_295#_M1004_d N_A_1745_329#_M1004_g N_VPWR_M1004_s VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.1134 AS=0.1134 PD=1.38 PS=1.38 NRD=2.3443 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1040 N_VPWR_M1040_d N_A_1745_329#_M1040_g N_A_2447_47#_M1040_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.1725 AS=0.27 PD=1.345 PS=2.54 NRD=5.91 NRS=0.9653 M=1
+ R=5.55556 SA=90000.2 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1012 N_Q_M1012_d N_A_2447_47#_M1012_g N_VPWR_M1040_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.1725 PD=1.29 PS=1.345 NRD=0.9653 NRS=6.8753 M=1 R=5.55556
+ SA=90000.7 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1016 N_Q_M1012_d N_A_2447_47#_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.17 PD=1.29 PS=1.34 NRD=0.9653 NRS=10.8153 M=1 R=5.55556
+ SA=90001.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1025 N_Q_M1025_d N_A_2447_47#_M1025_g N_VPWR_M1016_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.17 PD=1.29 PS=1.34 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.7 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1029 N_Q_M1025_d N_A_2447_47#_M1029_g N_VPWR_M1029_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.32 PD=1.29 PS=2.64 NRD=0.9653 NRS=10.8153 M=1 R=5.55556
+ SA=90002.2 SB=90000.2 A=0.18 P=2.36 MULT=1
DX46_noxref VNB VPB NWDIODE A=24.9738 P=34.33
c_132 VNB 0 1.07953e-19 $X=0.145 $Y=-0.085
c_279 VPB 0 7.24997e-20 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__sdfstp_4.pxi.spice"
*
.ends
*
*
