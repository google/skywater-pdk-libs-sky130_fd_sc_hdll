* File: sky130_fd_sc_hdll__o21ba_1.pex.spice
* Created: Wed Sep  2 08:43:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O21BA_1%A_79_199# 1 2 7 9 10 12 14 16 19 23 29 32
+ 35
r76 33 35 0.268087 $w=5.78e-07 $l=1.3e-08 $layer=LI1_cond $X=2.432 $Y=1.745
+ $X2=2.445 $Y2=1.745
r77 31 33 9.42427 $w=5.78e-07 $l=4.57e-07 $layer=LI1_cond $X=1.975 $Y=1.745
+ $X2=2.432 $Y2=1.745
r78 31 32 8.37612 $w=5.78e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=1.745
+ $X2=1.89 $Y2=1.745
r79 26 29 5.48283 $w=3.28e-07 $l=1.57e-07 $layer=LI1_cond $X=0.595 $Y=1.16
+ $X2=0.752 $Y2=1.16
r80 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.595
+ $Y=1.16 $X2=0.595 $Y2=1.16
r81 21 33 4.51232 $w=3.05e-07 $l=2.9e-07 $layer=LI1_cond $X=2.432 $Y=2.035
+ $X2=2.432 $Y2=1.745
r82 21 23 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=2.432 $Y=2.035
+ $X2=2.432 $Y2=2.3
r83 17 31 8.09873 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=1.975 $Y=1.455
+ $X2=1.975 $Y2=1.745
r84 17 19 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=1.975 $Y=1.455
+ $X2=1.975 $Y2=0.57
r85 16 32 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.86 $Y=1.95
+ $X2=1.89 $Y2=1.95
r86 14 16 6.93832 $w=1.7e-07 $l=1.44375e-07 $layer=LI1_cond $X=0.752 $Y=1.865
+ $X2=0.86 $Y2=1.95
r87 13 29 3.26307 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=0.752 $Y=1.325
+ $X2=0.752 $Y2=1.16
r88 13 14 28.9451 $w=2.13e-07 $l=5.4e-07 $layer=LI1_cond $X=0.752 $Y=1.325
+ $X2=0.752 $Y2=1.865
r89 10 27 38.5336 $w=3.07e-07 $l=1.70895e-07 $layer=POLY_cond $X=0.55 $Y=0.995
+ $X2=0.562 $Y2=1.16
r90 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.55 $Y=0.995
+ $X2=0.55 $Y2=0.56
r91 7 27 47.4309 $w=3.07e-07 $l=2.81514e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.562 $Y2=1.16
r92 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r93 2 35 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.485 $X2=2.445 $Y2=1.62
r94 2 23 400 $w=1.7e-07 $l=8.89129e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.485 $X2=2.445 $Y2=2.3
r95 1 19 182 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_NDIFF $count=1 $X=1.85
+ $Y=0.235 $X2=1.975 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_1%B1_N 1 3 4 6 7 15
c29 4 0 2.13581e-19 $X=1.06 $Y=1.41
r30 7 15 2.30489 $w=3.48e-07 $l=7e-08 $layer=LI1_cond $X=1.205 $Y=1.16 $X2=1.205
+ $Y2=1.23
r31 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.135
+ $Y=1.16 $X2=1.135 $Y2=1.16
r32 4 10 48.651 $w=2.87e-07 $l=2.76134e-07 $layer=POLY_cond $X=1.06 $Y=1.41
+ $X2=1.115 $Y2=1.16
r33 4 6 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.06 $Y=1.41 $X2=1.06
+ $Y2=1.695
r34 1 10 38.6443 $w=2.87e-07 $l=2.0106e-07 $layer=POLY_cond $X=1.035 $Y=0.995
+ $X2=1.115 $Y2=1.16
r35 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.035 $Y=0.995
+ $X2=1.035 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_1%A_222_93# 1 2 7 9 10 12 13 14 15 22 25
r50 25 26 17.4286 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=1.295 $Y=0.655
+ $X2=1.635 $Y2=0.655
r51 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.635
+ $Y=1.16 $X2=1.635 $Y2=1.16
r52 20 22 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.635 $Y=1.525
+ $X2=1.635 $Y2=1.16
r53 19 26 2.70854 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.635 $Y=0.825
+ $X2=1.635 $Y2=0.655
r54 19 22 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.635 $Y=0.825
+ $X2=1.635 $Y2=1.16
r55 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.55 $Y=1.61
+ $X2=1.635 $Y2=1.525
r56 15 17 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.55 $Y=1.61
+ $X2=1.295 $Y2=1.61
r57 13 23 81.3105 $w=3.3e-07 $l=4.65e-07 $layer=POLY_cond $X=2.1 $Y=1.16
+ $X2=1.635 $Y2=1.16
r58 13 14 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=2.1 $Y=1.16
+ $X2=2.2 $Y2=1.202
r59 10 14 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=2.225 $Y=0.995
+ $X2=2.2 $Y2=1.202
r60 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.225 $Y=0.995
+ $X2=2.225 $Y2=0.56
r61 7 14 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=2.2 $Y=1.41 $X2=2.2
+ $Y2=1.202
r62 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.2 $Y=1.41 $X2=2.2
+ $Y2=1.985
r63 2 17 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.15
+ $Y=1.485 $X2=1.295 $Y2=1.61
r64 1 25 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=1.11
+ $Y=0.465 $X2=1.295 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_1%A2 1 3 4 6 7 13
r28 7 13 7.92208 $w=2.08e-07 $l=1.5e-07 $layer=LI1_cond $X=2.6 $Y=1.18 $X2=2.45
+ $Y2=1.18
r29 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.645
+ $Y=1.16 $X2=2.645 $Y2=1.16
r30 4 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.705 $Y=0.995
+ $X2=2.645 $Y2=1.16
r31 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.705 $Y=0.995
+ $X2=2.705 $Y2=0.56
r32 1 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.68 $Y=1.41
+ $X2=2.645 $Y2=1.16
r33 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.68 $Y=1.41 $X2=2.68
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_1%A1 1 3 4 6 7 15
r19 7 15 9.77056 $w=2.08e-07 $l=1.85e-07 $layer=LI1_cond $X=3.185 $Y=1.18
+ $X2=3.37 $Y2=1.18
r20 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.185
+ $Y=1.16 $X2=3.185 $Y2=1.16
r21 4 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.15 $Y=1.41
+ $X2=3.185 $Y2=1.16
r22 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.15 $Y=1.41 $X2=3.15
+ $Y2=1.985
r23 1 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.125 $Y=0.995
+ $X2=3.185 $Y2=1.16
r24 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.125 $Y=0.995
+ $X2=3.125 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_1%X 1 2 10 15 16 17
c20 17 0 1.1384e-19 $X=0.23 $Y=2.21
c21 15 0 9.97411e-20 $X=0.26 $Y=1.645
r22 17 22 3.89797 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=0.255 $Y=2.21
+ $X2=0.255 $Y2=2.325
r23 15 16 6.33887 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.255 $Y=1.645
+ $X2=0.255 $Y2=1.48
r24 13 17 18.9814 $w=3.38e-07 $l=5.6e-07 $layer=LI1_cond $X=0.255 $Y=1.65
+ $X2=0.255 $Y2=2.21
r25 13 15 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=0.255 $Y=1.65
+ $X2=0.255 $Y2=1.645
r26 12 16 29.602 $w=2.53e-07 $l=6.55e-07 $layer=LI1_cond $X=0.212 $Y=0.825
+ $X2=0.212 $Y2=1.48
r27 10 12 6.27783 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=0.66
+ $X2=0.265 $Y2=0.825
r28 2 22 400 $w=1.7e-07 $l=9.00333e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.325
r29 2 15 400 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.645
r30 1 10 182 $w=1.7e-07 $l=4.83477e-07 $layer=licon1_NDIFF $count=1 $X=0.215
+ $Y=0.235 $X2=0.34 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_1%VPWR 1 2 3 12 16 18 20 24 26 31 36 42 45
+ 49
r47 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r48 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r49 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 40 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r51 40 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r52 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 37 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.1 $Y=2.72
+ $X2=1.935 $Y2=2.72
r54 37 39 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=2.1 $Y=2.72 $X2=2.99
+ $Y2=2.72
r55 36 48 5.16088 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=3.17 $Y=2.72
+ $X2=3.425 $Y2=2.72
r56 36 39 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.17 $Y=2.72
+ $X2=2.99 $Y2=2.72
r57 35 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 35 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r59 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r60 32 42 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.005 $Y=2.72
+ $X2=0.8 $Y2=2.72
r61 32 34 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.005 $Y=2.72
+ $X2=1.61 $Y2=2.72
r62 31 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.77 $Y=2.72
+ $X2=1.935 $Y2=2.72
r63 31 34 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.77 $Y=2.72
+ $X2=1.61 $Y2=2.72
r64 26 42 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.8 $Y2=2.72
r65 26 28 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r66 24 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r67 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r68 20 23 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=3.36 $Y=1.62
+ $X2=3.36 $Y2=2.3
r69 18 48 3.03581 $w=3.8e-07 $l=1.12916e-07 $layer=LI1_cond $X=3.36 $Y=2.635
+ $X2=3.425 $Y2=2.72
r70 18 23 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.36 $Y=2.635
+ $X2=3.36 $Y2=2.3
r71 14 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.935 $Y=2.635
+ $X2=1.935 $Y2=2.72
r72 14 16 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.935 $Y=2.635
+ $X2=1.935 $Y2=2.3
r73 10 42 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=2.635 $X2=0.8
+ $Y2=2.72
r74 10 12 9.69739 $w=4.08e-07 $l=3.45e-07 $layer=LI1_cond $X=0.8 $Y=2.635
+ $X2=0.8 $Y2=2.29
r75 3 23 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.24
+ $Y=1.485 $X2=3.385 $Y2=2.3
r76 3 20 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.24
+ $Y=1.485 $X2=3.385 $Y2=1.62
r77 2 16 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=1.81
+ $Y=1.485 $X2=1.935 $Y2=2.3
r78 1 12 600 $w=1.7e-07 $l=8.882e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.76 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_1%VGND 1 2 11 15 18 19 20 30 31 34
r43 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r44 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r45 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r46 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r47 25 28 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r48 25 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r49 24 27 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r50 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r51 22 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.76
+ $Y2=0
r52 22 24 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r53 20 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r54 18 27 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.83 $Y=0 $X2=2.53
+ $Y2=0
r55 18 19 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.83 $Y=0 $X2=2.915
+ $Y2=0
r56 17 30 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3 $Y=0 $X2=3.45
+ $Y2=0
r57 17 19 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=0 $X2=2.915
+ $Y2=0
r58 13 19 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0
r59 13 15 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0.39
r60 9 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=0.085 $X2=0.76
+ $Y2=0
r61 9 11 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.76 $Y=0.085
+ $X2=0.76 $Y2=0.66
r62 2 15 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.78
+ $Y=0.235 $X2=2.915 $Y2=0.39
r63 1 11 182 $w=1.7e-07 $l=4.87852e-07 $layer=licon1_NDIFF $count=1 $X=0.625
+ $Y=0.235 $X2=0.76 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_1%A_460_47# 1 2 9 11 12 15
r26 13 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.4 $Y=0.735
+ $X2=3.4 $Y2=0.39
r27 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.235 $Y=0.82
+ $X2=3.4 $Y2=0.735
r28 11 12 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.235 $Y=0.82
+ $X2=2.61 $Y2=0.82
r29 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.445 $Y=0.735
+ $X2=2.61 $Y2=0.82
r30 7 9 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.445 $Y=0.735
+ $X2=2.445 $Y2=0.39
r31 2 15 91 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_NDIFF $count=2 $X=3.2
+ $Y=0.235 $X2=3.4 $Y2=0.39
r32 1 9 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=2.3
+ $Y=0.235 $X2=2.445 $Y2=0.39
.ends

