* File: sky130_fd_sc_hdll__o21a_1.spice
* Created: Wed Sep  2 08:43:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o21a_1.pex.spice"
.subckt sky130_fd_sc_hdll__o21a_1  VNB VPB B1 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_83_21#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.182 PD=1.82 PS=1.86 NRD=0 NRS=2.76 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_A_302_47#_M1003_d N_B1_M1003_g N_A_83_21#_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.17225 PD=0.92 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g N_A_302_47#_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.08775 PD=0.98 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1007 N_A_302_47#_M1007_d N_A1_M1007_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.10725 PD=1.82 PS=0.98 NRD=0 NRS=10.152 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_83_21#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.3225 AS=0.29 PD=1.645 PS=2.58 NRD=2.9353 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.4 A=0.18 P=2.36 MULT=1
MM1005 N_A_83_21#_M1005_d N_B1_M1005_g N_VPWR_M1000_d VPB PHIGHVT L=0.18 W=1
+ AD=0.18 AS=0.3225 PD=1.36 PS=1.645 NRD=14.775 NRS=1.9503 M=1 R=5.55556
+ SA=90001 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1001 A_394_297# N_A2_M1001_g N_A_83_21#_M1005_d VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.18 PD=1.3 PS=1.36 NRD=18.6953 NRS=0.9653 M=1 R=5.55556 SA=90001.6
+ SB=90001 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g A_394_297# VPB PHIGHVT L=0.18 W=1 AD=0.61
+ AS=0.15 PD=3.22 PS=1.3 NRD=0.9653 NRS=18.6953 M=1 R=5.55556 SA=90002
+ SB=90000.5 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.778 P=10.41
pX9_noxref noxref_12 N_B1_X9_noxref_CONDUCTOR B1 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o21a_1.pxi.spice"
*
.ends
*
*
