# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__dfrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dfrtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.50000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.615000 1.975000 1.665000 ;
        RECT 1.455000 1.665000 1.780000 2.450000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.475000 0.255000  9.855000 0.735000 ;
        RECT  9.475000 0.735000 11.405000 0.905000 ;
        RECT  9.565000 1.455000 11.405000 1.625000 ;
        RECT  9.565000 1.625000  9.855000 2.465000 ;
        RECT 10.415000 0.255000 10.795000 0.735000 ;
        RECT 10.505000 1.625000 10.755000 2.465000 ;
        RECT 10.995000 0.905000 11.405000 1.455000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.277200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175000 0.765000 4.945000 1.015000 ;
        RECT 7.805000 1.035000 8.395000 1.405000 ;
        RECT 8.155000 0.635000 8.395000 1.035000 ;
      LAYER mcon ;
        RECT 4.285000 0.765000 4.455000 0.935000 ;
        RECT 4.645000 0.765000 4.815000 0.935000 ;
        RECT 7.870000 1.080000 8.040000 1.250000 ;
        RECT 8.165000 0.765000 8.335000 0.935000 ;
      LAYER met1 ;
        RECT 4.175000 0.735000 4.925000 0.780000 ;
        RECT 4.175000 0.780000 8.395000 0.920000 ;
        RECT 4.175000 0.920000 4.925000 0.965000 ;
        RECT 7.810000 0.920000 8.395000 1.280000 ;
        RECT 8.105000 0.735000 8.395000 0.780000 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 11.500000 0.085000 ;
        RECT  0.515000  0.085000  0.895000 0.465000 ;
        RECT  1.645000  0.085000  1.975000 0.445000 ;
        RECT  4.825000  0.085000  5.155000 0.545000 ;
        RECT  7.355000  0.085000  7.595000 0.525000 ;
        RECT  9.135000  0.085000  9.305000 0.895000 ;
        RECT 10.075000  0.085000 10.245000 0.555000 ;
        RECT 11.015000  0.085000 11.185000 0.555000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
        RECT 10.725000 -0.085000 10.895000 0.085000 ;
        RECT 11.185000 -0.085000 11.355000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.500000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 11.500000 2.805000 ;
        RECT  0.515000 2.135000  0.895000 2.635000 ;
        RECT  1.950000 2.175000  2.200000 2.635000 ;
        RECT  4.290000 2.205000  4.620000 2.635000 ;
        RECT  5.305000 2.175000  5.725000 2.635000 ;
        RECT  7.640000 2.175000  7.890000 2.635000 ;
        RECT  8.460000 2.255000  8.840000 2.635000 ;
        RECT  9.135000 1.575000  9.305000 2.635000 ;
        RECT 10.075000 1.795000 10.245000 2.635000 ;
        RECT 11.015000 1.795000 11.185000 2.635000 ;
      LAYER mcon ;
        RECT  0.145000 2.635000  0.315000 2.805000 ;
        RECT  0.605000 2.635000  0.775000 2.805000 ;
        RECT  1.065000 2.635000  1.235000 2.805000 ;
        RECT  1.525000 2.635000  1.695000 2.805000 ;
        RECT  1.985000 2.635000  2.155000 2.805000 ;
        RECT  2.445000 2.635000  2.615000 2.805000 ;
        RECT  2.905000 2.635000  3.075000 2.805000 ;
        RECT  3.365000 2.635000  3.535000 2.805000 ;
        RECT  3.825000 2.635000  3.995000 2.805000 ;
        RECT  4.285000 2.635000  4.455000 2.805000 ;
        RECT  4.745000 2.635000  4.915000 2.805000 ;
        RECT  5.205000 2.635000  5.375000 2.805000 ;
        RECT  5.665000 2.635000  5.835000 2.805000 ;
        RECT  6.125000 2.635000  6.295000 2.805000 ;
        RECT  6.585000 2.635000  6.755000 2.805000 ;
        RECT  7.045000 2.635000  7.215000 2.805000 ;
        RECT  7.505000 2.635000  7.675000 2.805000 ;
        RECT  7.965000 2.635000  8.135000 2.805000 ;
        RECT  8.425000 2.635000  8.595000 2.805000 ;
        RECT  8.885000 2.635000  9.055000 2.805000 ;
        RECT  9.345000 2.635000  9.515000 2.805000 ;
        RECT  9.805000 2.635000  9.975000 2.805000 ;
        RECT 10.265000 2.635000 10.435000 2.805000 ;
        RECT 10.725000 2.635000 10.895000 2.805000 ;
        RECT 11.185000 2.635000 11.355000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 11.500000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 0.345000  0.345000 0.635000 ;
      RECT 0.090000 0.635000  0.890000 0.805000 ;
      RECT 0.090000 1.795000  0.890000 1.965000 ;
      RECT 0.090000 1.965000  0.345000 2.465000 ;
      RECT 0.660000 0.805000  0.890000 1.795000 ;
      RECT 1.115000 0.345000  1.285000 2.465000 ;
      RECT 2.145000 0.305000  2.690000 0.475000 ;
      RECT 2.145000 0.475000  2.315000 1.835000 ;
      RECT 2.145000 1.835000  2.590000 2.005000 ;
      RECT 2.420000 2.005000  2.590000 2.135000 ;
      RECT 2.420000 2.135000  2.670000 2.465000 ;
      RECT 2.535000 0.765000  2.935000 1.385000 ;
      RECT 2.760000 1.575000  3.275000 1.965000 ;
      RECT 2.935000 2.135000  3.665000 2.465000 ;
      RECT 2.945000 0.305000  3.850000 0.475000 ;
      RECT 3.105000 0.765000  3.510000 0.985000 ;
      RECT 3.105000 0.985000  3.275000 1.575000 ;
      RECT 3.495000 1.185000  5.285000 1.355000 ;
      RECT 3.495000 1.355000  3.665000 2.135000 ;
      RECT 3.680000 0.475000  3.850000 1.185000 ;
      RECT 3.835000 1.865000  5.010000 2.035000 ;
      RECT 3.835000 2.035000  4.005000 2.375000 ;
      RECT 4.025000 1.525000  5.675000 1.695000 ;
      RECT 4.840000 2.035000  5.010000 2.375000 ;
      RECT 5.115000 1.005000  5.285000 1.185000 ;
      RECT 5.365000 0.275000  5.765000 0.445000 ;
      RECT 5.365000 0.445000  5.675000 0.835000 ;
      RECT 5.505000 0.835000  5.675000 1.525000 ;
      RECT 5.505000 1.695000  5.675000 1.835000 ;
      RECT 5.505000 1.835000  6.115000 2.005000 ;
      RECT 5.915000 0.705000  6.125000 1.495000 ;
      RECT 5.915000 1.495000  6.690000 1.655000 ;
      RECT 5.915000 1.655000  7.030000 1.665000 ;
      RECT 5.945000 2.005000  6.115000 2.465000 ;
      RECT 6.035000 0.255000  7.135000 0.535000 ;
      RECT 6.295000 0.705000  6.745000 1.325000 ;
      RECT 6.350000 2.125000  7.470000 2.465000 ;
      RECT 6.470000 1.665000  7.030000 1.955000 ;
      RECT 6.965000 0.535000  7.135000 1.315000 ;
      RECT 6.965000 1.315000  7.470000 1.485000 ;
      RECT 7.250000 1.485000  7.470000 1.575000 ;
      RECT 7.250000 1.575000  8.620000 1.745000 ;
      RECT 7.250000 1.745000  7.470000 2.125000 ;
      RECT 7.355000 0.695000  7.935000 0.865000 ;
      RECT 7.355000 0.865000  7.625000 1.145000 ;
      RECT 7.765000 0.295000  8.935000 0.465000 ;
      RECT 7.765000 0.465000  7.935000 0.695000 ;
      RECT 8.110000 1.915000  8.960000 2.085000 ;
      RECT 8.110000 2.085000  8.280000 2.375000 ;
      RECT 8.615000 0.465000  8.935000 0.820000 ;
      RECT 8.615000 0.820000  8.940000 1.075000 ;
      RECT 8.615000 1.075000 10.795000 1.285000 ;
      RECT 8.615000 1.285000  8.960000 1.295000 ;
      RECT 8.790000 1.295000  8.960000 1.915000 ;
    LAYER mcon ;
      RECT 0.660000 1.105000 0.830000 1.275000 ;
      RECT 1.115000 1.785000 1.285000 1.955000 ;
      RECT 2.595000 1.105000 2.765000 1.275000 ;
      RECT 3.105000 1.785000 3.275000 1.955000 ;
      RECT 6.525000 1.105000 6.695000 1.275000 ;
      RECT 6.525000 1.785000 6.695000 1.955000 ;
    LAYER met1 ;
      RECT 0.600000 1.075000 0.890000 1.120000 ;
      RECT 0.600000 1.120000 6.805000 1.260000 ;
      RECT 0.600000 1.260000 0.890000 1.305000 ;
      RECT 1.005000 1.755000 1.345000 1.800000 ;
      RECT 1.005000 1.800000 6.805000 1.940000 ;
      RECT 1.005000 1.940000 1.345000 1.985000 ;
      RECT 2.535000 1.075000 2.825000 1.120000 ;
      RECT 2.535000 1.260000 2.825000 1.305000 ;
      RECT 3.045000 1.755000 3.335000 1.800000 ;
      RECT 3.045000 1.940000 3.335000 1.985000 ;
      RECT 6.465000 1.075000 6.805000 1.120000 ;
      RECT 6.465000 1.260000 6.805000 1.305000 ;
      RECT 6.465000 1.755000 6.805000 1.800000 ;
      RECT 6.465000 1.940000 6.805000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dfrtp_4
