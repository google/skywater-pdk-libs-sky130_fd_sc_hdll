* File: sky130_fd_sc_hdll__o221ai_2.pxi.spice
* Created: Wed Sep  2 08:44:59 2020
* 
x_PM_SKY130_FD_SC_HDLL__O221AI_2%C1 N_C1_c_87_n N_C1_M1006_g N_C1_c_83_n
+ N_C1_M1002_g N_C1_c_88_n N_C1_M1018_g N_C1_c_84_n N_C1_M1013_g C1 N_C1_c_86_n
+ PM_SKY130_FD_SC_HDLL__O221AI_2%C1
x_PM_SKY130_FD_SC_HDLL__O221AI_2%B1 N_B1_c_126_n N_B1_M1000_g N_B1_c_127_n
+ N_B1_M1003_g N_B1_c_128_n N_B1_M1010_g N_B1_c_129_n N_B1_M1014_g N_B1_c_135_n
+ N_B1_c_130_n N_B1_c_131_n N_B1_c_132_n B1 B1 PM_SKY130_FD_SC_HDLL__O221AI_2%B1
x_PM_SKY130_FD_SC_HDLL__O221AI_2%B2 N_B2_c_203_n N_B2_M1007_g N_B2_c_207_n
+ N_B2_M1004_g N_B2_c_208_n N_B2_M1008_g N_B2_c_204_n N_B2_M1015_g B2
+ N_B2_c_205_n N_B2_c_206_n B2 PM_SKY130_FD_SC_HDLL__O221AI_2%B2
x_PM_SKY130_FD_SC_HDLL__O221AI_2%A1 N_A1_c_246_n N_A1_M1005_g N_A1_c_247_n
+ N_A1_M1009_g N_A1_c_248_n N_A1_M1011_g N_A1_c_249_n N_A1_M1017_g N_A1_c_256_n
+ N_A1_c_250_n N_A1_c_251_n N_A1_c_252_n A1 A1 PM_SKY130_FD_SC_HDLL__O221AI_2%A1
x_PM_SKY130_FD_SC_HDLL__O221AI_2%A2 N_A2_c_319_n N_A2_M1001_g N_A2_c_323_n
+ N_A2_M1016_g N_A2_c_324_n N_A2_M1019_g N_A2_c_320_n N_A2_M1012_g A2
+ N_A2_c_322_n A2 PM_SKY130_FD_SC_HDLL__O221AI_2%A2
x_PM_SKY130_FD_SC_HDLL__O221AI_2%VPWR N_VPWR_M1006_s N_VPWR_M1018_s
+ N_VPWR_M1010_d N_VPWR_M1011_s N_VPWR_c_367_n N_VPWR_c_368_n N_VPWR_c_369_n
+ N_VPWR_c_370_n N_VPWR_c_371_n N_VPWR_c_372_n N_VPWR_c_373_n N_VPWR_c_374_n
+ VPWR N_VPWR_c_375_n N_VPWR_c_366_n N_VPWR_c_377_n N_VPWR_c_378_n
+ PM_SKY130_FD_SC_HDLL__O221AI_2%VPWR
x_PM_SKY130_FD_SC_HDLL__O221AI_2%Y N_Y_M1002_d N_Y_M1006_d N_Y_M1004_s
+ N_Y_M1016_s N_Y_c_440_n N_Y_c_445_n N_Y_c_476_n N_Y_c_457_n N_Y_c_446_n
+ N_Y_c_439_n N_Y_c_454_n N_Y_c_461_n N_Y_c_455_n N_Y_c_470_n Y Y
+ PM_SKY130_FD_SC_HDLL__O221AI_2%Y
x_PM_SKY130_FD_SC_HDLL__O221AI_2%A_410_297# N_A_410_297#_M1000_s
+ N_A_410_297#_M1008_d N_A_410_297#_c_508_n N_A_410_297#_c_514_n
+ N_A_410_297#_c_516_n PM_SKY130_FD_SC_HDLL__O221AI_2%A_410_297#
x_PM_SKY130_FD_SC_HDLL__O221AI_2%A_802_297# N_A_802_297#_M1005_d
+ N_A_802_297#_M1019_d N_A_802_297#_c_530_n N_A_802_297#_c_529_n
+ N_A_802_297#_c_536_n PM_SKY130_FD_SC_HDLL__O221AI_2%A_802_297#
x_PM_SKY130_FD_SC_HDLL__O221AI_2%A_28_47# N_A_28_47#_M1002_s N_A_28_47#_M1013_s
+ N_A_28_47#_M1003_d N_A_28_47#_M1015_s N_A_28_47#_c_543_n N_A_28_47#_c_544_n
+ N_A_28_47#_c_551_n N_A_28_47#_c_545_n N_A_28_47#_c_546_n N_A_28_47#_c_547_n
+ PM_SKY130_FD_SC_HDLL__O221AI_2%A_28_47#
x_PM_SKY130_FD_SC_HDLL__O221AI_2%A_320_47# N_A_320_47#_M1003_s
+ N_A_320_47#_M1007_d N_A_320_47#_M1014_s N_A_320_47#_M1001_s
+ N_A_320_47#_M1017_s N_A_320_47#_c_592_n N_A_320_47#_c_642_p
+ N_A_320_47#_c_593_n N_A_320_47#_c_594_n N_A_320_47#_c_613_n
+ N_A_320_47#_c_595_n N_A_320_47#_c_596_n N_A_320_47#_c_597_n
+ PM_SKY130_FD_SC_HDLL__O221AI_2%A_320_47#
x_PM_SKY130_FD_SC_HDLL__O221AI_2%VGND N_VGND_M1009_d N_VGND_M1012_d
+ N_VGND_c_660_n N_VGND_c_661_n N_VGND_c_662_n N_VGND_c_663_n N_VGND_c_664_n
+ N_VGND_c_665_n VGND N_VGND_c_666_n N_VGND_c_667_n
+ PM_SKY130_FD_SC_HDLL__O221AI_2%VGND
cc_1 VNB N_C1_c_83_n 0.0221646f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_2 VNB N_C1_c_84_n 0.0219018f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=0.995
cc_3 VNB C1 0.00869944f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_C1_c_86_n 0.0666947f $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=1.202
cc_5 VNB N_B1_c_126_n 0.0289223f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_6 VNB N_B1_c_127_n 0.0217065f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_7 VNB N_B1_c_128_n 0.0227592f $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=1.41
cc_8 VNB N_B1_c_129_n 0.0180397f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=0.995
cc_9 VNB N_B1_c_130_n 0.012072f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.202
cc_10 VNB N_B1_c_131_n 0.00215682f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.202
cc_11 VNB N_B1_c_132_n 0.00350331f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=1.202
cc_12 VNB N_B2_c_203_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_13 VNB N_B2_c_204_n 0.0173947f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=0.995
cc_14 VNB N_B2_c_205_n 0.00141641f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.202
cc_15 VNB N_B2_c_206_n 0.0356367f $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=1.202
cc_16 VNB N_A1_c_246_n 0.0222035f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_17 VNB N_A1_c_247_n 0.017338f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_18 VNB N_A1_c_248_n 0.0295756f $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=1.41
cc_19 VNB N_A1_c_249_n 0.0221445f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=0.995
cc_20 VNB N_A1_c_250_n 2.72331e-19 $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_21 VNB N_A1_c_251_n 0.00350331f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.202
cc_22 VNB N_A1_c_252_n 0.00200001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB A1 0.0221414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A2_c_319_n 0.0169338f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_25 VNB N_A2_c_320_n 0.0173947f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=0.995
cc_26 VNB A2 0.00141439f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_27 VNB N_A2_c_322_n 0.0356338f $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=1.202
cc_28 VNB N_VPWR_c_366_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_Y_c_439_n 0.00198262f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_28_47#_c_543_n 0.0095692f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_31 VNB N_A_28_47#_c_544_n 0.017326f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.202
cc_32 VNB N_A_28_47#_c_545_n 0.00229934f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.202
cc_33 VNB N_A_28_47#_c_546_n 0.00559164f $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=1.202
cc_34 VNB N_A_28_47#_c_547_n 0.0192549f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_320_47#_c_592_n 0.00262034f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_36 VNB N_A_320_47#_c_593_n 0.00337798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_320_47#_c_594_n 0.00828262f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_320_47#_c_595_n 0.0137528f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_320_47#_c_596_n 0.0187437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_320_47#_c_597_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_660_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=1.985
cc_42 VNB N_VGND_c_661_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_43 VNB N_VGND_c_662_n 0.0957397f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_44 VNB N_VGND_c_663_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_45 VNB N_VGND_c_664_n 0.0193035f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.202
cc_46 VNB N_VGND_c_665_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=1.202
cc_47 VNB N_VGND_c_666_n 0.023262f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_667_n 0.305295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VPB N_C1_c_87_n 0.0202702f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_50 VPB N_C1_c_88_n 0.0188045f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=1.41
cc_51 VPB N_C1_c_86_n 0.0335337f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=1.202
cc_52 VPB N_B1_c_126_n 0.030133f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_53 VPB N_B1_c_128_n 0.0256643f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=1.41
cc_54 VPB N_B1_c_135_n 0.00674463f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_55 VPB N_B1_c_130_n 0.00448438f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.202
cc_56 VPB N_B1_c_131_n 0.00156923f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.202
cc_57 VPB N_B1_c_132_n 0.00272944f $X=-0.19 $Y=1.305 $X2=0.995 $Y2=1.202
cc_58 VPB N_B2_c_207_n 0.0159754f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=0.995
cc_59 VPB N_B2_c_208_n 0.0159779f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=1.41
cc_60 VPB N_B2_c_206_n 0.0192421f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=1.202
cc_61 VPB N_A1_c_246_n 0.0256643f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_62 VPB N_A1_c_248_n 0.0345571f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=1.41
cc_63 VPB N_A1_c_256_n 0.00659403f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_64 VPB N_A1_c_250_n 0.00130718f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_65 VPB N_A1_c_251_n 0.00272944f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.202
cc_66 VPB N_A2_c_323_n 0.0159779f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=0.995
cc_67 VPB N_A2_c_324_n 0.0159751f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=1.41
cc_68 VPB N_A2_c_322_n 0.0192668f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=1.202
cc_69 VPB N_VPWR_c_367_n 0.0114496f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_70 VPB N_VPWR_c_368_n 0.00824103f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.202
cc_71 VPB N_VPWR_c_369_n 0.00561515f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_370_n 0.00835273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_371_n 0.0403375f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_372_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_373_n 0.0417635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_374_n 0.00391723f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_375_n 0.0113717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_366_n 0.0522956f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_377_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_378_n 0.0229095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_Y_c_440_n 6.37077e-19 $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_82 VPB N_Y_c_439_n 0.00113129f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 N_C1_c_88_n N_B1_c_130_n 0.00502141f $X=0.97 $Y=1.41 $X2=0 $Y2=0
cc_84 N_C1_c_86_n N_B1_c_130_n 0.0102649f $X=0.97 $Y=1.202 $X2=0 $Y2=0
cc_85 N_C1_c_87_n N_VPWR_c_368_n 0.0055335f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_86 C1 N_VPWR_c_368_n 0.0193718f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_87 N_C1_c_86_n N_VPWR_c_368_n 0.00610779f $X=0.97 $Y=1.202 $X2=0 $Y2=0
cc_88 N_C1_c_87_n N_VPWR_c_366_n 0.0133252f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_89 N_C1_c_88_n N_VPWR_c_366_n 0.00821414f $X=0.97 $Y=1.41 $X2=0 $Y2=0
cc_90 N_C1_c_87_n N_VPWR_c_377_n 0.00702461f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_91 N_C1_c_88_n N_VPWR_c_377_n 0.00702461f $X=0.97 $Y=1.41 $X2=0 $Y2=0
cc_92 N_C1_c_88_n N_VPWR_c_378_n 0.00514457f $X=0.97 $Y=1.41 $X2=0 $Y2=0
cc_93 N_C1_c_87_n N_Y_c_440_n 5.49698e-19 $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_94 N_C1_c_88_n N_Y_c_440_n 0.00218415f $X=0.97 $Y=1.41 $X2=0 $Y2=0
cc_95 N_C1_c_86_n N_Y_c_440_n 0.00155289f $X=0.97 $Y=1.202 $X2=0 $Y2=0
cc_96 N_C1_c_88_n N_Y_c_445_n 0.007541f $X=0.97 $Y=1.41 $X2=0 $Y2=0
cc_97 N_C1_c_83_n N_Y_c_446_n 0.00779402f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_98 N_C1_c_86_n N_Y_c_446_n 7.95032e-19 $X=0.97 $Y=1.202 $X2=0 $Y2=0
cc_99 N_C1_c_87_n N_Y_c_439_n 8.69791e-19 $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_100 N_C1_c_83_n N_Y_c_439_n 0.00269965f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_101 N_C1_c_88_n N_Y_c_439_n 7.15981e-19 $X=0.97 $Y=1.41 $X2=0 $Y2=0
cc_102 N_C1_c_84_n N_Y_c_439_n 0.00263234f $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_103 C1 N_Y_c_439_n 0.0119245f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_104 N_C1_c_86_n N_Y_c_439_n 0.0344199f $X=0.97 $Y=1.202 $X2=0 $Y2=0
cc_105 N_C1_c_88_n N_Y_c_454_n 7.63508e-19 $X=0.97 $Y=1.41 $X2=0 $Y2=0
cc_106 N_C1_c_88_n N_Y_c_455_n 0.0170995f $X=0.97 $Y=1.41 $X2=0 $Y2=0
cc_107 N_C1_c_83_n N_A_28_47#_c_544_n 0.00441832f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_108 C1 N_A_28_47#_c_544_n 0.0192857f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_109 N_C1_c_86_n N_A_28_47#_c_544_n 0.00621075f $X=0.97 $Y=1.202 $X2=0 $Y2=0
cc_110 N_C1_c_83_n N_A_28_47#_c_551_n 0.0115007f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_111 N_C1_c_84_n N_A_28_47#_c_551_n 0.0140389f $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_112 C1 N_A_28_47#_c_551_n 0.00165805f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_113 N_C1_c_86_n N_A_28_47#_c_551_n 0.00167844f $X=0.97 $Y=1.202 $X2=0 $Y2=0
cc_114 N_C1_c_84_n N_A_28_47#_c_546_n 4.79383e-19 $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_115 N_C1_c_83_n N_VGND_c_662_n 0.00357877f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_116 N_C1_c_84_n N_VGND_c_662_n 0.00357877f $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_117 N_C1_c_83_n N_VGND_c_667_n 0.00635999f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_118 N_C1_c_84_n N_VGND_c_667_n 0.00668309f $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_119 N_B1_c_127_n N_B2_c_203_n 0.0270078f $X=1.985 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_120 N_B1_c_126_n N_B2_c_207_n 0.0378374f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_121 N_B1_c_135_n N_B2_c_207_n 0.0120058f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_122 N_B1_c_131_n N_B2_c_207_n 9.86626e-19 $X=2.185 $Y=1.345 $X2=0 $Y2=0
cc_123 N_B1_c_128_n N_B2_c_208_n 0.0378352f $X=3.37 $Y=1.41 $X2=0 $Y2=0
cc_124 N_B1_c_135_n N_B2_c_208_n 0.0112841f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_125 N_B1_c_132_n N_B2_c_208_n 0.00101445f $X=3.345 $Y=1.16 $X2=0 $Y2=0
cc_126 N_B1_c_129_n N_B2_c_204_n 0.0219899f $X=3.395 $Y=0.995 $X2=0 $Y2=0
cc_127 N_B1_c_126_n N_B2_c_205_n 2.06438e-19 $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_128 N_B1_c_128_n N_B2_c_205_n 6.86695e-19 $X=3.37 $Y=1.41 $X2=0 $Y2=0
cc_129 N_B1_c_135_n N_B2_c_205_n 0.0461557f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_130 N_B1_c_131_n N_B2_c_205_n 0.0176043f $X=2.185 $Y=1.345 $X2=0 $Y2=0
cc_131 N_B1_c_132_n N_B2_c_205_n 0.0176354f $X=3.345 $Y=1.16 $X2=0 $Y2=0
cc_132 N_B1_c_126_n N_B2_c_206_n 0.0263716f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_133 N_B1_c_128_n N_B2_c_206_n 0.0263033f $X=3.37 $Y=1.41 $X2=0 $Y2=0
cc_134 N_B1_c_135_n N_B2_c_206_n 0.00803891f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_135 N_B1_c_131_n N_B2_c_206_n 0.00526937f $X=2.185 $Y=1.345 $X2=0 $Y2=0
cc_136 N_B1_c_132_n N_B2_c_206_n 0.00392336f $X=3.345 $Y=1.16 $X2=0 $Y2=0
cc_137 N_B1_c_128_n N_A1_c_246_n 0.056924f $X=3.37 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_138 N_B1_c_132_n N_A1_c_246_n 0.00168165f $X=3.345 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_139 N_B1_c_129_n N_A1_c_247_n 0.0154445f $X=3.395 $Y=0.995 $X2=0 $Y2=0
cc_140 N_B1_c_128_n N_A1_c_251_n 0.00168165f $X=3.37 $Y=1.41 $X2=0 $Y2=0
cc_141 N_B1_c_132_n N_A1_c_251_n 0.0455154f $X=3.345 $Y=1.16 $X2=0 $Y2=0
cc_142 N_B1_c_130_n N_VPWR_M1018_s 0.0127537f $X=1.915 $Y=1.345 $X2=0 $Y2=0
cc_143 N_B1_c_132_n N_VPWR_M1010_d 0.00161183f $X=3.345 $Y=1.16 $X2=0 $Y2=0
cc_144 N_B1_c_128_n N_VPWR_c_369_n 0.00322023f $X=3.37 $Y=1.41 $X2=0 $Y2=0
cc_145 N_B1_c_126_n N_VPWR_c_371_n 0.00702461f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_146 N_B1_c_128_n N_VPWR_c_371_n 0.00702461f $X=3.37 $Y=1.41 $X2=0 $Y2=0
cc_147 N_B1_c_126_n N_VPWR_c_366_n 0.00823967f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_148 N_B1_c_128_n N_VPWR_c_366_n 0.00716301f $X=3.37 $Y=1.41 $X2=0 $Y2=0
cc_149 N_B1_c_126_n N_VPWR_c_378_n 0.00514457f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_150 N_B1_c_135_n N_Y_M1004_s 0.00187091f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_151 N_B1_c_128_n N_Y_c_457_n 0.0140422f $X=3.37 $Y=1.41 $X2=0 $Y2=0
cc_152 N_B1_c_135_n N_Y_c_457_n 0.0218268f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_153 N_B1_c_132_n N_Y_c_457_n 0.0201576f $X=3.345 $Y=1.16 $X2=0 $Y2=0
cc_154 N_B1_c_130_n N_Y_c_439_n 0.0364668f $X=1.915 $Y=1.345 $X2=0 $Y2=0
cc_155 N_B1_c_135_n N_Y_c_461_n 0.0135474f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_156 N_B1_c_126_n N_Y_c_455_n 0.0156745f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_157 N_B1_c_130_n N_Y_c_455_n 0.0938664f $X=1.915 $Y=1.345 $X2=0 $Y2=0
cc_158 N_B1_c_135_n N_A_410_297#_M1000_s 0.00103364f $X=3.18 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_159 N_B1_c_131_n N_A_410_297#_M1000_s 8.61234e-19 $X=2.185 $Y=1.345 $X2=-0.19
+ $Y2=-0.24
cc_160 N_B1_c_135_n N_A_410_297#_M1008_d 0.00172342f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_161 N_B1_c_132_n N_A_410_297#_M1008_d 7.76441e-19 $X=3.345 $Y=1.16 $X2=0
+ $Y2=0
cc_162 N_B1_c_127_n N_A_28_47#_c_546_n 0.00285215f $X=1.985 $Y=0.995 $X2=0 $Y2=0
cc_163 N_B1_c_130_n N_A_28_47#_c_546_n 0.0228439f $X=1.915 $Y=1.345 $X2=0 $Y2=0
cc_164 N_B1_c_126_n N_A_28_47#_c_547_n 0.00441892f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_165 N_B1_c_127_n N_A_28_47#_c_547_n 0.0141874f $X=1.985 $Y=0.995 $X2=0 $Y2=0
cc_166 N_B1_c_128_n N_A_28_47#_c_547_n 0.00233856f $X=3.37 $Y=1.41 $X2=0 $Y2=0
cc_167 N_B1_c_135_n N_A_28_47#_c_547_n 0.0117006f $X=3.18 $Y=1.53 $X2=0 $Y2=0
cc_168 N_B1_c_130_n N_A_28_47#_c_547_n 0.0671947f $X=1.915 $Y=1.345 $X2=0 $Y2=0
cc_169 N_B1_c_132_n N_A_28_47#_c_547_n 0.00976394f $X=3.345 $Y=1.16 $X2=0 $Y2=0
cc_170 N_B1_c_127_n N_A_320_47#_c_592_n 0.00886996f $X=1.985 $Y=0.995 $X2=0
+ $Y2=0
cc_171 N_B1_c_128_n N_A_320_47#_c_592_n 3.99938e-19 $X=3.37 $Y=1.41 $X2=0 $Y2=0
cc_172 N_B1_c_129_n N_A_320_47#_c_592_n 0.0112894f $X=3.395 $Y=0.995 $X2=0 $Y2=0
cc_173 N_B1_c_132_n N_A_320_47#_c_592_n 0.00499729f $X=3.345 $Y=1.16 $X2=0 $Y2=0
cc_174 N_B1_c_128_n N_A_320_47#_c_594_n 2.55742e-19 $X=3.37 $Y=1.41 $X2=0 $Y2=0
cc_175 N_B1_c_129_n N_A_320_47#_c_594_n 2.31743e-19 $X=3.395 $Y=0.995 $X2=0
+ $Y2=0
cc_176 N_B1_c_132_n N_A_320_47#_c_594_n 0.00353546f $X=3.345 $Y=1.16 $X2=0 $Y2=0
cc_177 N_B1_c_127_n N_VGND_c_662_n 0.00357877f $X=1.985 $Y=0.995 $X2=0 $Y2=0
cc_178 N_B1_c_129_n N_VGND_c_662_n 0.00357877f $X=3.395 $Y=0.995 $X2=0 $Y2=0
cc_179 N_B1_c_127_n N_VGND_c_667_n 0.00657948f $X=1.985 $Y=0.995 $X2=0 $Y2=0
cc_180 N_B1_c_129_n N_VGND_c_667_n 0.00568976f $X=3.395 $Y=0.995 $X2=0 $Y2=0
cc_181 N_B2_c_207_n N_VPWR_c_371_n 0.00429453f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_182 N_B2_c_208_n N_VPWR_c_371_n 0.00429453f $X=2.9 $Y=1.41 $X2=0 $Y2=0
cc_183 N_B2_c_207_n N_VPWR_c_366_n 0.00609021f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_184 N_B2_c_208_n N_VPWR_c_366_n 0.00609021f $X=2.9 $Y=1.41 $X2=0 $Y2=0
cc_185 N_B2_c_208_n N_Y_c_457_n 0.0108425f $X=2.9 $Y=1.41 $X2=0 $Y2=0
cc_186 N_B2_c_207_n N_Y_c_455_n 0.0108425f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_187 N_B2_c_207_n N_A_410_297#_c_508_n 0.0099733f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_188 N_B2_c_208_n N_A_410_297#_c_508_n 0.0099733f $X=2.9 $Y=1.41 $X2=0 $Y2=0
cc_189 N_B2_c_203_n N_A_28_47#_c_547_n 0.0120916f $X=2.405 $Y=0.995 $X2=0 $Y2=0
cc_190 N_B2_c_204_n N_A_28_47#_c_547_n 0.0118103f $X=2.925 $Y=0.995 $X2=0 $Y2=0
cc_191 N_B2_c_205_n N_A_28_47#_c_547_n 0.0480026f $X=2.665 $Y=1.16 $X2=0 $Y2=0
cc_192 N_B2_c_206_n N_A_28_47#_c_547_n 0.0047334f $X=2.9 $Y=1.202 $X2=0 $Y2=0
cc_193 N_B2_c_203_n N_A_320_47#_c_592_n 0.00886996f $X=2.405 $Y=0.995 $X2=0
+ $Y2=0
cc_194 N_B2_c_204_n N_A_320_47#_c_592_n 0.00923997f $X=2.925 $Y=0.995 $X2=0
+ $Y2=0
cc_195 N_B2_c_203_n N_VGND_c_662_n 0.00357877f $X=2.405 $Y=0.995 $X2=0 $Y2=0
cc_196 N_B2_c_204_n N_VGND_c_662_n 0.00357877f $X=2.925 $Y=0.995 $X2=0 $Y2=0
cc_197 N_B2_c_203_n N_VGND_c_667_n 0.00549573f $X=2.405 $Y=0.995 $X2=0 $Y2=0
cc_198 N_B2_c_204_n N_VGND_c_667_n 0.00561849f $X=2.925 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A1_c_247_n N_A2_c_319_n 0.0258911f $X=3.945 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_200 N_A1_c_246_n N_A2_c_323_n 0.0378352f $X=3.92 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A1_c_256_n N_A2_c_323_n 0.0112841f $X=5.095 $Y=1.53 $X2=0 $Y2=0
cc_202 N_A1_c_251_n N_A2_c_323_n 0.00101445f $X=3.895 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A1_c_248_n N_A2_c_324_n 0.0219473f $X=5.33 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A1_c_256_n N_A2_c_324_n 0.0182308f $X=5.095 $Y=1.53 $X2=0 $Y2=0
cc_205 N_A1_c_250_n N_A2_c_324_n 7.34002e-19 $X=5.18 $Y=1.445 $X2=0 $Y2=0
cc_206 N_A1_c_249_n N_A2_c_320_n 0.0213001f $X=5.355 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A1_c_246_n A2 6.74634e-19 $X=3.92 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A1_c_256_n A2 0.0420374f $X=5.095 $Y=1.53 $X2=0 $Y2=0
cc_209 N_A1_c_251_n A2 0.0175037f $X=3.895 $Y=1.16 $X2=0 $Y2=0
cc_210 N_A1_c_252_n A2 0.0143894f $X=5.265 $Y=1.175 $X2=0 $Y2=0
cc_211 N_A1_c_246_n N_A2_c_322_n 0.0263033f $X=3.92 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A1_c_248_n N_A2_c_322_n 0.026336f $X=5.33 $Y=1.41 $X2=0 $Y2=0
cc_213 N_A1_c_256_n N_A2_c_322_n 0.00803891f $X=5.095 $Y=1.53 $X2=0 $Y2=0
cc_214 N_A1_c_250_n N_A2_c_322_n 0.0029218f $X=5.18 $Y=1.445 $X2=0 $Y2=0
cc_215 N_A1_c_251_n N_A2_c_322_n 0.00392336f $X=3.895 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A1_c_252_n N_A2_c_322_n 0.00164489f $X=5.265 $Y=1.175 $X2=0 $Y2=0
cc_217 N_A1_c_251_n N_VPWR_M1010_d 0.00161183f $X=3.895 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A1_c_246_n N_VPWR_c_369_n 0.00537492f $X=3.92 $Y=1.41 $X2=0 $Y2=0
cc_219 N_A1_c_248_n N_VPWR_c_370_n 0.0122183f $X=5.33 $Y=1.41 $X2=0 $Y2=0
cc_220 N_A1_c_256_n N_VPWR_c_370_n 0.0104762f $X=5.095 $Y=1.53 $X2=0 $Y2=0
cc_221 A1 N_VPWR_c_370_n 0.0166332f $X=5.62 $Y=1.105 $X2=0 $Y2=0
cc_222 N_A1_c_246_n N_VPWR_c_373_n 0.00702461f $X=3.92 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A1_c_248_n N_VPWR_c_373_n 0.00702461f $X=5.33 $Y=1.41 $X2=0 $Y2=0
cc_224 N_A1_c_246_n N_VPWR_c_366_n 0.00721773f $X=3.92 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A1_c_248_n N_VPWR_c_366_n 0.0135742f $X=5.33 $Y=1.41 $X2=0 $Y2=0
cc_226 N_A1_c_256_n N_Y_M1016_s 0.00187091f $X=5.095 $Y=1.53 $X2=0 $Y2=0
cc_227 N_A1_c_246_n N_Y_c_457_n 0.0140422f $X=3.92 $Y=1.41 $X2=0 $Y2=0
cc_228 N_A1_c_256_n N_Y_c_457_n 0.0218268f $X=5.095 $Y=1.53 $X2=0 $Y2=0
cc_229 N_A1_c_251_n N_Y_c_457_n 0.0201576f $X=3.895 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A1_c_256_n N_Y_c_470_n 0.0135474f $X=5.095 $Y=1.53 $X2=0 $Y2=0
cc_231 N_A1_c_256_n N_A_802_297#_M1005_d 0.00172342f $X=5.095 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_232 N_A1_c_251_n N_A_802_297#_M1005_d 7.76441e-19 $X=3.895 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_233 N_A1_c_256_n N_A_802_297#_M1019_d 0.00189183f $X=5.095 $Y=1.53 $X2=0
+ $Y2=0
cc_234 N_A1_c_256_n N_A_802_297#_c_529_n 0.014924f $X=5.095 $Y=1.53 $X2=0 $Y2=0
cc_235 N_A1_c_246_n N_A_320_47#_c_593_n 0.00205406f $X=3.92 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A1_c_247_n N_A_320_47#_c_593_n 0.0124528f $X=3.945 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A1_c_256_n N_A_320_47#_c_593_n 0.00574667f $X=5.095 $Y=1.53 $X2=0 $Y2=0
cc_238 N_A1_c_251_n N_A_320_47#_c_593_n 0.0198504f $X=3.895 $Y=1.16 $X2=0 $Y2=0
cc_239 N_A1_c_246_n N_A_320_47#_c_594_n 0.00239959f $X=3.92 $Y=1.41 $X2=0 $Y2=0
cc_240 N_A1_c_251_n N_A_320_47#_c_594_n 0.010525f $X=3.895 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A1_c_247_n N_A_320_47#_c_613_n 5.32212e-19 $X=3.945 $Y=0.995 $X2=0
+ $Y2=0
cc_242 N_A1_c_248_n N_A_320_47#_c_595_n 0.00443298f $X=5.33 $Y=1.41 $X2=0 $Y2=0
cc_243 N_A1_c_249_n N_A_320_47#_c_595_n 0.00903373f $X=5.355 $Y=0.995 $X2=0
+ $Y2=0
cc_244 N_A1_c_256_n N_A_320_47#_c_595_n 0.00684545f $X=5.095 $Y=1.53 $X2=0 $Y2=0
cc_245 N_A1_c_252_n N_A_320_47#_c_595_n 0.0137248f $X=5.265 $Y=1.175 $X2=0 $Y2=0
cc_246 A1 N_A_320_47#_c_595_n 0.0372828f $X=5.62 $Y=1.105 $X2=0 $Y2=0
cc_247 N_A1_c_249_n N_A_320_47#_c_596_n 0.00850899f $X=5.355 $Y=0.995 $X2=0
+ $Y2=0
cc_248 N_A1_c_247_n N_VGND_c_660_n 0.00268723f $X=3.945 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A1_c_249_n N_VGND_c_661_n 0.00359159f $X=5.355 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A1_c_247_n N_VGND_c_662_n 0.00439206f $X=3.945 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A1_c_249_n N_VGND_c_666_n 0.00396605f $X=5.355 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A1_c_247_n N_VGND_c_667_n 0.00630876f $X=3.945 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A1_c_249_n N_VGND_c_667_n 0.00677957f $X=5.355 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A2_c_323_n N_VPWR_c_373_n 0.00429453f $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_255 N_A2_c_324_n N_VPWR_c_373_n 0.00429453f $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_256 N_A2_c_323_n N_VPWR_c_366_n 0.00609021f $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_257 N_A2_c_324_n N_VPWR_c_366_n 0.00609021f $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_258 N_A2_c_323_n N_Y_c_457_n 0.0108425f $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A2_c_323_n N_A_802_297#_c_530_n 0.0100164f $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A2_c_324_n N_A_802_297#_c_530_n 0.0143148f $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A2_c_319_n N_A_320_47#_c_593_n 0.00845772f $X=4.365 $Y=0.995 $X2=0
+ $Y2=0
cc_262 A2 N_A_320_47#_c_593_n 0.00896514f $X=4.705 $Y=1.105 $X2=0 $Y2=0
cc_263 N_A2_c_319_n N_A_320_47#_c_613_n 0.00644736f $X=4.365 $Y=0.995 $X2=0
+ $Y2=0
cc_264 N_A2_c_320_n N_A_320_47#_c_595_n 0.011927f $X=4.885 $Y=0.995 $X2=0 $Y2=0
cc_265 A2 N_A_320_47#_c_595_n 0.00589753f $X=4.705 $Y=1.105 $X2=0 $Y2=0
cc_266 N_A2_c_320_n N_A_320_47#_c_596_n 5.82315e-19 $X=4.885 $Y=0.995 $X2=0
+ $Y2=0
cc_267 N_A2_c_319_n N_A_320_47#_c_597_n 0.00135102f $X=4.365 $Y=0.995 $X2=0
+ $Y2=0
cc_268 A2 N_A_320_47#_c_597_n 0.0307352f $X=4.705 $Y=1.105 $X2=0 $Y2=0
cc_269 N_A2_c_322_n N_A_320_47#_c_597_n 0.00486271f $X=4.86 $Y=1.202 $X2=0 $Y2=0
cc_270 N_A2_c_319_n N_VGND_c_660_n 0.00268723f $X=4.365 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A2_c_320_n N_VGND_c_661_n 0.00276126f $X=4.885 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A2_c_319_n N_VGND_c_664_n 0.00424416f $X=4.365 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A2_c_320_n N_VGND_c_664_n 0.00437852f $X=4.885 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A2_c_319_n N_VGND_c_667_n 0.00600559f $X=4.365 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A2_c_320_n N_VGND_c_667_n 0.00627444f $X=4.885 $Y=0.995 $X2=0 $Y2=0
cc_276 N_VPWR_c_366_n N_Y_M1006_d 0.00310442f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_277 N_VPWR_c_366_n N_Y_M1004_s 0.00231289f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_278 N_VPWR_c_366_n N_Y_M1016_s 0.00232092f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_279 N_VPWR_c_368_n N_Y_c_440_n 0.00195268f $X=0.265 $Y=1.65 $X2=0 $Y2=0
cc_280 N_VPWR_c_366_n N_Y_c_476_n 0.00955092f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_281 N_VPWR_c_377_n N_Y_c_476_n 0.0149311f $X=1.08 $Y=2.465 $X2=0 $Y2=0
cc_282 N_VPWR_M1010_d N_Y_c_457_n 0.0101824f $X=3.46 $Y=1.485 $X2=0 $Y2=0
cc_283 N_VPWR_c_369_n N_Y_c_457_n 0.020234f $X=3.605 $Y=2.3 $X2=0 $Y2=0
cc_284 N_VPWR_c_366_n N_Y_c_457_n 0.0165712f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_285 N_VPWR_c_366_n N_Y_c_454_n 0.00142525f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_286 N_VPWR_M1018_s N_Y_c_455_n 0.0187907f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_287 N_VPWR_c_366_n N_Y_c_455_n 0.01579f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_288 N_VPWR_c_378_n N_Y_c_455_n 0.0547305f $X=1.85 $Y=2.465 $X2=0 $Y2=0
cc_289 N_VPWR_c_366_n N_A_410_297#_M1000_s 0.00241598f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_290 N_VPWR_c_366_n N_A_410_297#_M1008_d 0.00241598f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_371_n N_A_410_297#_c_508_n 0.0386815f $X=3.48 $Y=2.72 $X2=0
+ $Y2=0
cc_292 N_VPWR_c_366_n N_A_410_297#_c_508_n 0.0239224f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_293 N_VPWR_c_371_n N_A_410_297#_c_514_n 0.014332f $X=3.48 $Y=2.72 $X2=0 $Y2=0
cc_294 N_VPWR_c_366_n N_A_410_297#_c_514_n 0.00938745f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_295 N_VPWR_c_371_n N_A_410_297#_c_516_n 0.0143006f $X=3.48 $Y=2.72 $X2=0
+ $Y2=0
cc_296 N_VPWR_c_366_n N_A_410_297#_c_516_n 0.00938288f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_297 N_VPWR_c_366_n N_A_802_297#_M1005_d 0.00241598f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_298 N_VPWR_c_366_n N_A_802_297#_M1019_d 0.00297222f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_299 N_VPWR_c_373_n N_A_802_297#_c_530_n 0.0536835f $X=5.485 $Y=2.72 $X2=0
+ $Y2=0
cc_300 N_VPWR_c_366_n N_A_802_297#_c_530_n 0.0335464f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_301 N_VPWR_c_373_n N_A_802_297#_c_536_n 0.0143006f $X=5.485 $Y=2.72 $X2=0
+ $Y2=0
cc_302 N_VPWR_c_366_n N_A_802_297#_c_536_n 0.00938288f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_303 N_Y_c_455_n N_A_410_297#_M1000_s 0.00369247f $X=2.54 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_304 N_Y_c_457_n N_A_410_297#_M1008_d 0.00367036f $X=4.5 $Y=1.87 $X2=0 $Y2=0
cc_305 N_Y_M1004_s N_A_410_297#_c_508_n 0.00352392f $X=2.52 $Y=1.485 $X2=0 $Y2=0
cc_306 N_Y_c_457_n N_A_410_297#_c_508_n 0.00608347f $X=4.5 $Y=1.87 $X2=0 $Y2=0
cc_307 N_Y_c_461_n N_A_410_297#_c_508_n 0.0127274f $X=2.665 $Y=1.87 $X2=0 $Y2=0
cc_308 N_Y_c_455_n N_A_410_297#_c_508_n 0.00608347f $X=2.54 $Y=1.87 $X2=0 $Y2=0
cc_309 N_Y_c_455_n N_A_410_297#_c_514_n 0.0131392f $X=2.54 $Y=1.87 $X2=0 $Y2=0
cc_310 N_Y_c_457_n N_A_410_297#_c_516_n 0.0130645f $X=4.5 $Y=1.87 $X2=0 $Y2=0
cc_311 N_Y_c_457_n N_A_802_297#_M1005_d 0.00367036f $X=4.5 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_312 N_Y_M1016_s N_A_802_297#_c_530_n 0.00352392f $X=4.48 $Y=1.485 $X2=0 $Y2=0
cc_313 N_Y_c_457_n N_A_802_297#_c_530_n 0.00608347f $X=4.5 $Y=1.87 $X2=0 $Y2=0
cc_314 N_Y_c_470_n N_A_802_297#_c_530_n 0.0127274f $X=4.625 $Y=1.87 $X2=0 $Y2=0
cc_315 N_Y_c_457_n N_A_802_297#_c_536_n 0.0130645f $X=4.5 $Y=1.87 $X2=0 $Y2=0
cc_316 N_Y_c_446_n N_A_28_47#_c_544_n 0.0168291f $X=0.777 $Y=0.755 $X2=0 $Y2=0
cc_317 N_Y_c_439_n N_A_28_47#_c_544_n 0.00100415f $X=0.755 $Y=1.445 $X2=0 $Y2=0
cc_318 N_Y_M1002_d N_A_28_47#_c_551_n 0.00400389f $X=0.6 $Y=0.235 $X2=0 $Y2=0
cc_319 N_Y_c_446_n N_A_28_47#_c_551_n 0.0201165f $X=0.777 $Y=0.755 $X2=0 $Y2=0
cc_320 N_Y_c_439_n N_A_28_47#_c_546_n 0.00137098f $X=0.755 $Y=1.445 $X2=0 $Y2=0
cc_321 N_Y_M1002_d N_VGND_c_667_n 0.00256987f $X=0.6 $Y=0.235 $X2=0 $Y2=0
cc_322 N_A_28_47#_c_547_n N_A_320_47#_M1003_s 0.00435219f $X=3.135 $Y=0.73
+ $X2=-0.19 $Y2=-0.24
cc_323 N_A_28_47#_c_547_n N_A_320_47#_M1007_d 0.00279596f $X=3.135 $Y=0.73 $X2=0
+ $Y2=0
cc_324 N_A_28_47#_M1003_d N_A_320_47#_c_592_n 0.00312026f $X=2.06 $Y=0.235 $X2=0
+ $Y2=0
cc_325 N_A_28_47#_M1015_s N_A_320_47#_c_592_n 0.0041027f $X=3 $Y=0.235 $X2=0
+ $Y2=0
cc_326 N_A_28_47#_c_545_n N_A_320_47#_c_592_n 0.0188708f $X=1.245 $Y=0.475 $X2=0
+ $Y2=0
cc_327 N_A_28_47#_c_547_n N_A_320_47#_c_592_n 0.0966135f $X=3.135 $Y=0.73 $X2=0
+ $Y2=0
cc_328 N_A_28_47#_c_547_n N_A_320_47#_c_594_n 0.00140356f $X=3.135 $Y=0.73 $X2=0
+ $Y2=0
cc_329 N_A_28_47#_c_543_n N_VGND_c_662_n 0.0175572f $X=0.225 $Y=0.475 $X2=0
+ $Y2=0
cc_330 N_A_28_47#_c_551_n N_VGND_c_662_n 0.0425444f $X=1.12 $Y=0.365 $X2=0 $Y2=0
cc_331 N_A_28_47#_c_545_n N_VGND_c_662_n 0.0173343f $X=1.245 $Y=0.475 $X2=0
+ $Y2=0
cc_332 N_A_28_47#_c_547_n N_VGND_c_662_n 0.00349681f $X=3.135 $Y=0.73 $X2=0
+ $Y2=0
cc_333 N_A_28_47#_M1002_s N_VGND_c_667_n 0.00250318f $X=0.14 $Y=0.235 $X2=0
+ $Y2=0
cc_334 N_A_28_47#_M1013_s N_VGND_c_667_n 0.00209324f $X=1.07 $Y=0.235 $X2=0
+ $Y2=0
cc_335 N_A_28_47#_M1003_d N_VGND_c_667_n 0.00216833f $X=2.06 $Y=0.235 $X2=0
+ $Y2=0
cc_336 N_A_28_47#_M1015_s N_VGND_c_667_n 0.00256987f $X=3 $Y=0.235 $X2=0 $Y2=0
cc_337 N_A_28_47#_c_543_n N_VGND_c_667_n 0.00961275f $X=0.225 $Y=0.475 $X2=0
+ $Y2=0
cc_338 N_A_28_47#_c_551_n N_VGND_c_667_n 0.0273233f $X=1.12 $Y=0.365 $X2=0 $Y2=0
cc_339 N_A_28_47#_c_545_n N_VGND_c_667_n 0.00961652f $X=1.245 $Y=0.475 $X2=0
+ $Y2=0
cc_340 N_A_28_47#_c_547_n N_VGND_c_667_n 0.00886559f $X=3.135 $Y=0.73 $X2=0
+ $Y2=0
cc_341 N_A_320_47#_c_593_n N_VGND_M1009_d 0.00165819f $X=4.41 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_342 N_A_320_47#_c_595_n N_VGND_M1012_d 0.00251047f $X=5.35 $Y=0.815 $X2=0
+ $Y2=0
cc_343 N_A_320_47#_c_593_n N_VGND_c_660_n 0.0116528f $X=4.41 $Y=0.82 $X2=0 $Y2=0
cc_344 N_A_320_47#_c_595_n N_VGND_c_661_n 0.0127273f $X=5.35 $Y=0.815 $X2=0
+ $Y2=0
cc_345 N_A_320_47#_c_596_n N_VGND_c_661_n 0.0223967f $X=5.565 $Y=0.39 $X2=0
+ $Y2=0
cc_346 N_A_320_47#_c_592_n N_VGND_c_662_n 0.112077f $X=3.52 $Y=0.365 $X2=0 $Y2=0
cc_347 N_A_320_47#_c_642_p N_VGND_c_662_n 0.0216064f $X=3.685 $Y=0.475 $X2=0
+ $Y2=0
cc_348 N_A_320_47#_c_593_n N_VGND_c_662_n 0.00248756f $X=4.41 $Y=0.82 $X2=0
+ $Y2=0
cc_349 N_A_320_47#_c_593_n N_VGND_c_664_n 0.00193763f $X=4.41 $Y=0.82 $X2=0
+ $Y2=0
cc_350 N_A_320_47#_c_613_n N_VGND_c_664_n 0.0231806f $X=4.625 $Y=0.39 $X2=0
+ $Y2=0
cc_351 N_A_320_47#_c_595_n N_VGND_c_664_n 0.00254521f $X=5.35 $Y=0.815 $X2=0
+ $Y2=0
cc_352 N_A_320_47#_c_595_n N_VGND_c_666_n 0.00199443f $X=5.35 $Y=0.815 $X2=0
+ $Y2=0
cc_353 N_A_320_47#_c_596_n N_VGND_c_666_n 0.024373f $X=5.565 $Y=0.39 $X2=0 $Y2=0
cc_354 N_A_320_47#_M1003_s N_VGND_c_667_n 0.00250339f $X=1.6 $Y=0.235 $X2=0
+ $Y2=0
cc_355 N_A_320_47#_M1007_d N_VGND_c_667_n 0.00295535f $X=2.48 $Y=0.235 $X2=0
+ $Y2=0
cc_356 N_A_320_47#_M1014_s N_VGND_c_667_n 0.00330638f $X=3.47 $Y=0.235 $X2=0
+ $Y2=0
cc_357 N_A_320_47#_M1001_s N_VGND_c_667_n 0.00304143f $X=4.44 $Y=0.235 $X2=0
+ $Y2=0
cc_358 N_A_320_47#_M1017_s N_VGND_c_667_n 0.00209319f $X=5.43 $Y=0.235 $X2=0
+ $Y2=0
cc_359 N_A_320_47#_c_592_n N_VGND_c_667_n 0.0703895f $X=3.52 $Y=0.365 $X2=0
+ $Y2=0
cc_360 N_A_320_47#_c_642_p N_VGND_c_667_n 0.0126938f $X=3.685 $Y=0.475 $X2=0
+ $Y2=0
cc_361 N_A_320_47#_c_593_n N_VGND_c_667_n 0.00943347f $X=4.41 $Y=0.82 $X2=0
+ $Y2=0
cc_362 N_A_320_47#_c_613_n N_VGND_c_667_n 0.0143352f $X=4.625 $Y=0.39 $X2=0
+ $Y2=0
cc_363 N_A_320_47#_c_595_n N_VGND_c_667_n 0.00977515f $X=5.35 $Y=0.815 $X2=0
+ $Y2=0
cc_364 N_A_320_47#_c_596_n N_VGND_c_667_n 0.0141066f $X=5.565 $Y=0.39 $X2=0
+ $Y2=0
