* NGSPICE file created from sky130_fd_sc_hdll__or3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__or3b_2 A B C_N VGND VNB VPB VPWR X
M1000 a_448_297# A VPWR VPB phighvt w=420000u l=180000u
+  ad=1.302e+11p pd=1.46e+06u as=6.164e+11p ps=5.43e+06u
M1001 X a_186_21# VGND VNB nshort w=650000u l=150000u
+  ad=3.4125e+11p pd=2.35e+06u as=5.5575e+11p ps=5.52e+06u
M1002 VGND B a_186_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.268e+11p ps=2.76e+06u
M1003 a_186_21# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_546_297# B a_448_297# VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1005 a_186_21# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR C_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1007 VPWR a_186_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=4e+11p ps=2.8e+06u
M1008 a_186_21# a_27_47# a_546_297# VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1009 VGND C_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1010 X a_186_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_186_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

