* File: sky130_fd_sc_hdll__nor2b_1.pex.spice
* Created: Wed Sep  2 08:39:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR2B_1%B_N 3 5 7 8 9 19
r26 9 19 1.70732 $w=2.68e-07 $l=4e-08 $layer=LI1_cond $X=0.65 $Y=1.58 $X2=0.65
+ $Y2=1.62
r27 8 9 17.9269 $w=2.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.65 $Y=1.16 $X2=0.65
+ $Y2=1.58
r28 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6 $Y=1.16
+ $X2=0.6 $Y2=1.16
r29 5 13 46.8073 $w=3.2e-07 $l=2.82843e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.565 $Y2=1.16
r30 5 7 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.695
r31 1 13 41.562 $w=3.2e-07 $l=2.27596e-07 $layer=POLY_cond $X=0.47 $Y=0.975
+ $X2=0.565 $Y2=1.16
r32 1 3 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.47 $Y=0.975 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2B_1%A 1 3 4 6 7
r32 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.16 $X2=1.12 $Y2=1.16
r33 4 10 49.9093 $w=2.71e-07 $l=2.7157e-07 $layer=POLY_cond $X=1.175 $Y=1.41
+ $X2=1.13 $Y2=1.16
r34 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.175 $Y=1.41
+ $X2=1.175 $Y2=1.985
r35 1 10 38.8824 $w=2.71e-07 $l=1.69926e-07 $layer=POLY_cond $X=1.14 $Y=0.995
+ $X2=1.13 $Y2=1.16
r36 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.14 $Y=0.995 $X2=1.14
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2B_1%A_27_47# 1 2 7 9 10 12 15 19 20 22 24 27
+ 30
r55 30 33 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=1.16
+ $X2=1.675 $Y2=1.325
r56 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.16 $X2=1.65 $Y2=1.16
r57 25 27 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.4 $Y=1.58 $X2=1.57
+ $Y2=1.58
r58 24 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=1.495
+ $X2=1.57 $Y2=1.58
r59 24 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.57 $Y=1.495
+ $X2=1.57 $Y2=1.325
r60 21 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.4 $Y=1.665 $X2=1.4
+ $Y2=1.58
r61 21 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.4 $Y=1.665 $X2=1.4
+ $Y2=1.915
r62 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.315 $Y=2
+ $X2=1.4 $Y2=1.915
r63 19 20 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.315 $Y=2 $X2=0.345
+ $Y2=2
r64 15 18 58.7746 $w=2.48e-07 $l=1.275e-06 $layer=LI1_cond $X=0.22 $Y=0.455
+ $X2=0.22 $Y2=1.73
r65 13 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.22 $Y=1.915
+ $X2=0.345 $Y2=2
r66 13 18 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=0.22 $Y=1.915
+ $X2=0.22 $Y2=1.73
r67 10 31 45.964 $w=3.43e-07 $l=2.91548e-07 $layer=POLY_cond $X=1.585 $Y=1.41
+ $X2=1.675 $Y2=1.16
r68 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.585 $Y=1.41
+ $X2=1.585 $Y2=1.985
r69 7 31 38.7084 $w=3.43e-07 $l=2.14942e-07 $layer=POLY_cond $X=1.56 $Y=0.995
+ $X2=1.675 $Y2=1.16
r70 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.56 $Y=0.995 $X2=1.56
+ $Y2=0.56
r71 2 18 600 $w=1.7e-07 $l=3.01081e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.73
r72 1 15 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2B_1%VPWR 1 6 9 10 11 21 22
r26 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r27 19 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r28 18 21 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r29 18 19 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r30 15 19 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r31 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r32 11 15 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r33 9 14 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=2.72
+ $X2=0.69 $Y2=2.72
r34 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.775 $Y=2.72
+ $X2=0.94 $Y2=2.72
r35 8 18 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.105 $Y=2.72
+ $X2=1.15 $Y2=2.72
r36 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.105 $Y=2.72
+ $X2=0.94 $Y2=2.72
r37 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.94 $Y=2.635 $X2=0.94
+ $Y2=2.72
r38 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.94 $Y=2.635
+ $X2=0.94 $Y2=2.34
r39 1 6 600 $w=1.7e-07 $l=1.01713e-06 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.94 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2B_1%Y 1 2 9 11 12 15 18 19
r40 18 19 9.16965 $w=5.58e-07 $l=1.5e-07 $layer=LI1_cond $X=1.935 $Y=2 $X2=1.935
+ $Y2=1.85
r41 15 18 4.48529 $w=5.58e-07 $l=2.1e-07 $layer=LI1_cond $X=1.935 $Y=2.21
+ $X2=1.935 $Y2=2
r42 13 19 58.8434 $w=1.78e-07 $l=9.55e-07 $layer=LI1_cond $X=2.125 $Y=0.895
+ $X2=2.125 $Y2=1.85
r43 11 13 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.035 $Y=0.81
+ $X2=2.125 $Y2=0.895
r44 11 12 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.035 $Y=0.81
+ $X2=1.515 $Y2=0.81
r45 7 12 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=1.325 $Y=0.725
+ $X2=1.515 $Y2=0.81
r46 7 9 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.325 $Y=0.725
+ $X2=1.325 $Y2=0.39
r47 2 18 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.675
+ $Y=1.485 $X2=1.82 $Y2=2
r48 1 9 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.215
+ $Y=0.235 $X2=1.35 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2B_1%VGND 1 2 11 13 15 17 19 25 29
r31 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r32 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r33 23 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r34 23 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r35 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r36 20 25 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=0.82
+ $Y2=0
r37 20 22 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=1.61
+ $Y2=0
r38 19 28 5.08477 $w=1.7e-07 $l=2.82e-07 $layer=LI1_cond $X=1.735 $Y=0 $X2=2.017
+ $Y2=0
r39 19 22 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.735 $Y=0 $X2=1.61
+ $Y2=0
r40 17 26 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r41 13 28 3.15544 $w=3.85e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.927 $Y=0.085
+ $X2=2.017 $Y2=0
r42 13 15 9.12974 $w=3.83e-07 $l=3.05e-07 $layer=LI1_cond $X=1.927 $Y=0.085
+ $X2=1.927 $Y2=0.39
r43 9 25 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=0.085
+ $X2=0.82 $Y2=0
r44 9 11 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=0.82 $Y=0.085
+ $X2=0.82 $Y2=0.39
r45 2 15 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.635
+ $Y=0.235 $X2=1.82 $Y2=0.39
r46 1 11 182 $w=1.7e-07 $l=4.05154e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.88 $Y2=0.39
.ends

