* File: sky130_fd_sc_hdll__nor2b_2.pex.spice
* Created: Thu Aug 27 19:15:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR2B_2%A 1 3 4 6 7 9 10 12 13 20 24
c37 10 0 1.19013e-19 $X=1.01 $Y=0.995
r38 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.01 $Y2=1.202
r39 18 20 43.1263 $w=3.8e-07 $l=3.4e-07 $layer=POLY_cond $X=0.645 $Y=1.202
+ $X2=0.985 $Y2=1.202
r40 18 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.645
+ $Y=1.16 $X2=0.645 $Y2=1.16
r41 16 18 16.4895 $w=3.8e-07 $l=1.3e-07 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.645 $Y2=1.202
r42 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.49 $Y=1.202
+ $X2=0.515 $Y2=1.202
r43 13 24 5.28139 $w=2.08e-07 $l=1e-07 $layer=LI1_cond $X=0.745 $Y=1.17
+ $X2=0.645 $Y2=1.17
r44 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=1.202
r45 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=0.56
r46 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r47 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r48 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r49 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r50 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.202
r51 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2B_2%A_271_21# 1 2 7 9 10 12 13 15 16 18 19 24
+ 27 31 35 37
c65 31 0 3.18361e-20 $X=2.68 $Y=0.68
r66 33 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=1.245
+ $X2=2.68 $Y2=1.16
r67 33 35 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=2.68 $Y=1.245
+ $X2=2.68 $Y2=2.28
r68 29 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=1.075
+ $X2=2.68 $Y2=1.16
r69 29 31 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.68 $Y=1.075
+ $X2=2.68 $Y2=0.68
r70 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.24
+ $Y=1.16 $X2=2.24 $Y2=1.16
r71 24 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=1.16
+ $X2=2.68 $Y2=1.16
r72 24 26 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.595 $Y=1.16
+ $X2=2.24 $Y2=1.16
r73 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.9 $Y=1.202
+ $X2=1.925 $Y2=1.202
r74 21 22 56.4447 $w=3.8e-07 $l=4.45e-07 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.9 $Y2=1.202
r75 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.43 $Y=1.202
+ $X2=1.455 $Y2=1.202
r76 19 27 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=2.025 $Y=1.16
+ $X2=2.24 $Y2=1.16
r77 19 23 13.6483 $w=3.8e-07 $l=1.19164e-07 $layer=POLY_cond $X=2.025 $Y=1.16
+ $X2=1.925 $Y2=1.202
r78 16 23 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r79 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r80 13 22 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.9 $Y=0.995
+ $X2=1.9 $Y2=1.202
r81 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.9 $Y=0.995 $X2=1.9
+ $Y2=0.56
r82 10 21 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r83 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r84 7 20 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=1.202
r85 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995 $X2=1.43
+ $Y2=0.56
r86 2 35 600 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=2.555
+ $Y=2.065 $X2=2.68 $Y2=2.28
r87 1 31 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=2.555
+ $Y=0.465 $X2=2.68 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2B_2%B_N 3 5 6 8 9 12 14 15 16 22
c32 12 0 3.18361e-20 $X=3.125 $Y=1.16
r33 15 16 14.7861 $w=2.63e-07 $l=3.4e-07 $layer=LI1_cond $X=3.402 $Y=1.53
+ $X2=3.402 $Y2=1.87
r34 14 15 8.50329 $w=4.33e-07 $l=2.55e-07 $layer=LI1_cond $X=3.402 $Y=1.275
+ $X2=3.402 $Y2=1.53
r35 12 23 37.7183 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=3.142 $Y=1.16
+ $X2=3.142 $Y2=1.325
r36 12 22 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=3.142 $Y=1.16
+ $X2=3.142 $Y2=0.995
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.125
+ $Y=1.16 $X2=3.125 $Y2=1.16
r38 9 14 3.86311 $w=2.1e-07 $l=1.32e-07 $layer=LI1_cond $X=3.27 $Y=1.17
+ $X2=3.402 $Y2=1.17
r39 9 11 7.65801 $w=2.08e-07 $l=1.45e-07 $layer=LI1_cond $X=3.27 $Y=1.17
+ $X2=3.125 $Y2=1.17
r40 6 8 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.075 $Y=1.99
+ $X2=3.075 $Y2=2.275
r41 5 6 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.075 $Y=1.89 $X2=3.075
+ $Y2=1.99
r42 5 23 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=3.075 $Y=1.89
+ $X2=3.075 $Y2=1.325
r43 3 22 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.05 $Y=0.675
+ $X2=3.05 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2B_2%A_27_297# 1 2 3 10 12 14 16 17 18 20 22
r39 20 31 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=2.295
+ $X2=2.18 $Y2=2.38
r40 20 22 26.4267 $w=2.88e-07 $l=6.65e-07 $layer=LI1_cond $X=2.18 $Y=2.295
+ $X2=2.18 $Y2=1.63
r41 19 29 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=2.38
+ $X2=1.22 $Y2=2.38
r42 18 31 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.035 $Y=2.38
+ $X2=2.18 $Y2=2.38
r43 18 19 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.035 $Y=2.38
+ $X2=1.345 $Y2=2.38
r44 17 29 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=2.295
+ $X2=1.22 $Y2=2.38
r45 16 27 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.22 $Y=1.655
+ $X2=1.22 $Y2=1.55
r46 16 17 29.5025 $w=2.48e-07 $l=6.4e-07 $layer=LI1_cond $X=1.22 $Y=1.655
+ $X2=1.22 $Y2=2.295
r47 15 25 4.35048 $w=2.1e-07 $l=1.6e-07 $layer=LI1_cond $X=0.405 $Y=1.55
+ $X2=0.245 $Y2=1.55
r48 14 27 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=1.55
+ $X2=1.22 $Y2=1.55
r49 14 15 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=1.55
+ $X2=0.405 $Y2=1.55
r50 10 25 2.855 $w=3.2e-07 $l=1.05e-07 $layer=LI1_cond $X=0.245 $Y=1.655
+ $X2=0.245 $Y2=1.55
r51 10 12 23.2289 $w=3.18e-07 $l=6.45e-07 $layer=LI1_cond $X=0.245 $Y=1.655
+ $X2=0.245 $Y2=2.3
r52 3 31 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=2.31
r53 3 22 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=1.63
r54 2 29 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.3
r55 2 27 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.62
r56 1 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r57 1 12 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2B_2%VPWR 1 2 11 13 15 17 19 28 32 34
r40 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r41 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r42 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r43 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r44 23 26 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 23 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r46 22 25 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r47 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r48 20 28 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=0.75 $Y2=2.72
r49 20 22 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=1.15 $Y2=2.72
r50 19 31 3.88626 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=3.185 $Y=2.72
+ $X2=3.432 $Y2=2.72
r51 19 25 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.185 $Y=2.72
+ $X2=2.99 $Y2=2.72
r52 17 29 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r53 17 34 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r54 13 31 3.2569 $w=2.5e-07 $l=1.58915e-07 $layer=LI1_cond $X=3.31 $Y=2.635
+ $X2=3.432 $Y2=2.72
r55 13 15 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=3.31 $Y=2.635
+ $X2=3.31 $Y2=2.31
r56 9 28 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r57 9 11 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2
r58 2 15 600 $w=1.7e-07 $l=3.09112e-07 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=2.065 $X2=3.31 $Y2=2.31
r59 1 11 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2B_2%Y 1 2 3 12 14 15 18 21 22 25
c45 15 0 1.19013e-19 $X=0.935 $Y=0.81
r46 22 25 3.63929 $w=3.78e-07 $l=1.2e-07 $layer=LI1_cond $X=1.665 $Y=0.51
+ $X2=1.665 $Y2=0.39
r47 20 22 6.5204 $w=3.78e-07 $l=2.15e-07 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.51
r48 20 21 3.01263 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.81
r49 16 21 3.01263 $w=3.15e-07 $l=9.66954e-08 $layer=LI1_cond $X=1.69 $Y=0.895
+ $X2=1.665 $Y2=0.81
r50 16 18 33.4208 $w=2.48e-07 $l=7.25e-07 $layer=LI1_cond $X=1.69 $Y=0.895
+ $X2=1.69 $Y2=1.62
r51 14 21 3.63293 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.475 $Y=0.81
+ $X2=1.665 $Y2=0.81
r52 14 15 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.475 $Y=0.81
+ $X2=0.935 $Y2=0.81
r53 10 15 8.37092 $w=1.7e-07 $l=2.38747e-07 $layer=LI1_cond $X=0.735 $Y=0.725
+ $X2=0.935 $Y2=0.81
r54 10 12 9.65171 $w=3.98e-07 $l=3.35e-07 $layer=LI1_cond $X=0.735 $Y=0.725
+ $X2=0.735 $Y2=0.39
r55 3 18 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=1.62
r56 2 25 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.505
+ $Y=0.235 $X2=1.69 $Y2=0.39
r57 1 12 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2B_2%VGND 1 2 3 4 13 15 17 21 25 27 29 32 33 34
+ 40 48 52
r51 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r52 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r53 43 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r54 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r55 40 51 3.92207 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=3.185 $Y=0 $X2=3.432
+ $Y2=0
r56 40 42 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.185 $Y=0 $X2=2.99
+ $Y2=0
r57 39 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r58 39 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r59 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r60 36 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.22
+ $Y2=0
r61 36 38 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=2.07
+ $Y2=0
r62 34 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r63 34 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r64 32 38 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.07
+ $Y2=0
r65 32 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.16
+ $Y2=0
r66 31 42 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.99
+ $Y2=0
r67 31 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.16
+ $Y2=0
r68 27 51 3.25516 $w=2.55e-07 $l=1.56844e-07 $layer=LI1_cond $X=3.312 $Y=0.085
+ $X2=3.432 $Y2=0
r69 27 29 26.8903 $w=2.53e-07 $l=5.95e-07 $layer=LI1_cond $X=3.312 $Y=0.085
+ $X2=3.312 $Y2=0.68
r70 23 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0
r71 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0.39
r72 19 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r73 19 21 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.39
r74 18 45 4.33083 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r75 17 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.22
+ $Y2=0
r76 17 18 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=0 $X2=0.365
+ $Y2=0
r77 13 45 3.02922 $w=2.8e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.182 $Y2=0
r78 13 15 12.5534 $w=2.78e-07 $l=3.05e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.225 $Y2=0.39
r79 4 29 182 $w=1.7e-07 $l=2.93258e-07 $layer=licon1_NDIFF $count=1 $X=3.125
+ $Y=0.465 $X2=3.31 $Y2=0.68
r80 3 25 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.975
+ $Y=0.235 $X2=2.16 $Y2=0.39
r81 2 21 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.235 $X2=1.22 $Y2=0.39
r82 1 15 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

