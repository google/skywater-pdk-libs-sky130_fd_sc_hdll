* File: sky130_fd_sc_hdll__nand4_1.pxi.spice
* Created: Wed Sep  2 08:38:17 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND4_1%D N_D_c_46_n N_D_M1004_g N_D_c_43_n N_D_M1006_g
+ D N_D_c_45_n PM_SKY130_FD_SC_HDLL__NAND4_1%D
x_PM_SKY130_FD_SC_HDLL__NAND4_1%C N_C_c_68_n N_C_M1000_g N_C_c_69_n N_C_M1001_g
+ C C C N_C_c_71_n C PM_SKY130_FD_SC_HDLL__NAND4_1%C
x_PM_SKY130_FD_SC_HDLL__NAND4_1%B N_B_c_104_n N_B_M1003_g N_B_c_105_n
+ N_B_M1007_g N_B_c_106_n N_B_c_107_n B PM_SKY130_FD_SC_HDLL__NAND4_1%B
x_PM_SKY130_FD_SC_HDLL__NAND4_1%A N_A_c_146_n N_A_M1002_g N_A_c_149_n
+ N_A_M1005_g A A N_A_c_147_n N_A_c_148_n PM_SKY130_FD_SC_HDLL__NAND4_1%A
x_PM_SKY130_FD_SC_HDLL__NAND4_1%VPWR N_VPWR_M1004_s N_VPWR_M1000_d
+ N_VPWR_M1005_d N_VPWR_c_175_n N_VPWR_c_176_n N_VPWR_c_177_n N_VPWR_c_178_n
+ N_VPWR_c_179_n N_VPWR_c_180_n N_VPWR_c_181_n VPWR N_VPWR_c_182_n
+ N_VPWR_c_174_n N_VPWR_c_184_n PM_SKY130_FD_SC_HDLL__NAND4_1%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND4_1%Y N_Y_M1002_d N_Y_M1004_d N_Y_M1007_d
+ N_Y_c_217_n N_Y_c_218_n N_Y_c_222_n N_Y_c_254_n N_Y_c_214_n N_Y_c_232_n Y
+ N_Y_c_215_n PM_SKY130_FD_SC_HDLL__NAND4_1%Y
x_PM_SKY130_FD_SC_HDLL__NAND4_1%VGND N_VGND_M1006_s N_VGND_c_260_n
+ N_VGND_c_261_n VGND N_VGND_c_262_n N_VGND_c_263_n
+ PM_SKY130_FD_SC_HDLL__NAND4_1%VGND
cc_1 VNB N_D_c_43_n 0.0226111f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB D 0.0139673f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_D_c_45_n 0.0370546f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_C_c_68_n 0.0248141f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_C_c_69_n 0.0168751f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB C 0.00259601f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_7 VNB N_C_c_71_n 9.39592e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_B_c_104_n 0.016758f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_9 VNB N_B_c_105_n 0.027656f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_10 VNB N_B_c_106_n 0.0011365f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B_c_107_n 0.0020905f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_12 VNB N_A_c_146_n 0.0225264f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_13 VNB N_A_c_147_n 0.0396652f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_14 VNB N_A_c_148_n 0.0241593f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VPWR_c_174_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_Y_c_214_n 0.00272979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_Y_c_215_n 0.0249461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_260_n 0.0115155f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_19 VNB N_VGND_c_261_n 0.0290471f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_20 VNB N_VGND_c_262_n 0.0637099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_263_n 0.171847f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VPB N_D_c_46_n 0.0212694f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_23 VPB D 0.00475375f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_24 VPB N_D_c_45_n 0.0177624f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_25 VPB N_C_c_68_n 0.026226f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_26 VPB N_C_c_71_n 0.00195866f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_B_c_105_n 0.026848f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_28 VPB N_B_c_107_n 9.4923e-19 $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_29 VPB N_A_c_149_n 0.0193513f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_30 VPB N_A_c_147_n 0.0183775f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_31 VPB N_A_c_148_n 0.0273723f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_175_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_33 VPB N_VPWR_c_176_n 0.0434419f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_34 VPB N_VPWR_c_177_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_178_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_179_n 0.0298966f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_180_n 0.0232629f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_181_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_182_n 0.0137583f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_174_n 0.0537295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_184_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_Y_c_214_n 0.00132922f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 N_D_c_46_n N_C_c_68_n 0.0100726f $X=0.495 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_44 D N_C_c_68_n 2.16942e-19 $X=0.15 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_45 N_D_c_45_n N_C_c_68_n 0.0261314f $X=0.495 $Y=1.202 $X2=-0.19 $Y2=-0.24
cc_46 N_D_c_43_n N_C_c_69_n 0.0281918f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_47 N_D_c_43_n C 0.00620227f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_48 D N_C_c_71_n 0.0221051f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_49 N_D_c_45_n N_C_c_71_n 0.00306671f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_50 N_D_c_46_n N_VPWR_c_176_n 0.00779021f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_51 D N_VPWR_c_176_n 0.0194376f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_52 N_D_c_45_n N_VPWR_c_176_n 0.00173333f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_53 N_D_c_46_n N_VPWR_c_177_n 0.00597712f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_54 N_D_c_46_n N_VPWR_c_174_n 0.0109312f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_55 N_D_c_46_n N_Y_c_217_n 0.00605425f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_56 N_D_c_46_n N_Y_c_218_n 0.0121679f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_57 N_D_c_43_n N_VGND_c_261_n 0.00483019f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_58 D N_VGND_c_261_n 0.0233168f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_59 N_D_c_45_n N_VGND_c_261_n 0.00211088f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_60 N_D_c_43_n N_VGND_c_262_n 0.00585385f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_61 N_D_c_43_n N_VGND_c_263_n 0.0116876f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_62 N_C_c_69_n N_B_c_104_n 0.0420218f $X=0.99 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_63 N_C_c_68_n N_B_c_105_n 0.0487615f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_64 N_C_c_71_n N_B_c_105_n 3.14501e-19 $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_65 N_C_c_69_n N_B_c_106_n 0.00129016f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_66 C N_B_c_106_n 0.00600179f $X=0.66 $Y=0.425 $X2=0 $Y2=0
cc_67 N_C_c_68_n N_B_c_107_n 0.00204979f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_68 N_C_c_71_n N_B_c_107_n 0.0271234f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_69 N_C_c_68_n B 0.00124263f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_70 N_C_c_69_n B 0.0125323f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_71 N_C_c_71_n B 0.00303576f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_72 N_C_c_68_n N_VPWR_c_177_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_73 N_C_c_68_n N_VPWR_c_178_n 0.0052072f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_74 N_C_c_68_n N_VPWR_c_174_n 0.0118942f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_75 N_C_c_68_n N_Y_c_217_n 0.0018341f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_76 N_C_c_71_n N_Y_c_217_n 0.0208725f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_77 N_C_c_68_n N_Y_c_218_n 0.0108293f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_78 N_C_c_68_n N_Y_c_222_n 0.0150546f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_79 N_C_c_71_n N_Y_c_222_n 0.0121426f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_80 N_C_c_69_n N_VGND_c_262_n 0.00535866f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_81 C N_VGND_c_262_n 0.012846f $X=0.66 $Y=0.425 $X2=0 $Y2=0
cc_82 N_C_c_69_n N_VGND_c_263_n 0.00973738f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_83 C N_VGND_c_263_n 0.00990262f $X=0.66 $Y=0.425 $X2=0 $Y2=0
cc_84 C A_119_47# 0.00790386f $X=0.66 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_85 N_B_c_104_n N_A_c_146_n 0.0254837f $X=1.41 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_86 B N_A_c_146_n 7.47222e-19 $X=1.17 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_87 N_B_c_105_n N_A_c_149_n 0.0075379f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_88 N_B_c_105_n N_A_c_147_n 0.0233591f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_89 N_B_c_107_n N_A_c_147_n 3.14127e-19 $X=1.47 $Y=1.16 $X2=0 $Y2=0
cc_90 N_B_c_105_n N_VPWR_c_178_n 0.00547142f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_91 N_B_c_105_n N_VPWR_c_180_n 0.00702461f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_92 N_B_c_105_n N_VPWR_c_174_n 0.0126959f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_93 N_B_c_105_n N_Y_c_218_n 6.38978e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_94 N_B_c_105_n N_Y_c_222_n 0.0152233f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_95 N_B_c_107_n N_Y_c_222_n 0.0188796f $X=1.47 $Y=1.16 $X2=0 $Y2=0
cc_96 B N_Y_c_222_n 0.00360423f $X=1.17 $Y=0.425 $X2=0 $Y2=0
cc_97 N_B_c_104_n N_Y_c_214_n 8.26784e-19 $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_98 N_B_c_105_n N_Y_c_214_n 0.0042985f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_99 N_B_c_106_n N_Y_c_214_n 0.00487915f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_100 N_B_c_107_n N_Y_c_214_n 0.0249362f $X=1.47 $Y=1.16 $X2=0 $Y2=0
cc_101 N_B_c_105_n N_Y_c_232_n 0.00370955f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_102 N_B_c_107_n N_Y_c_232_n 0.00367128f $X=1.47 $Y=1.16 $X2=0 $Y2=0
cc_103 N_B_c_104_n N_Y_c_215_n 0.0057426f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_104 B N_Y_c_215_n 0.0319866f $X=1.17 $Y=0.425 $X2=0 $Y2=0
cc_105 N_B_c_104_n N_VGND_c_262_n 0.00470326f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_106 B N_VGND_c_262_n 0.0174972f $X=1.17 $Y=0.425 $X2=0 $Y2=0
cc_107 N_B_c_104_n N_VGND_c_263_n 0.00821166f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_108 B N_VGND_c_263_n 0.0138313f $X=1.17 $Y=0.425 $X2=0 $Y2=0
cc_109 N_B_c_106_n A_213_47# 6.95655e-19 $X=1.33 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_110 B A_213_47# 0.00429481f $X=1.17 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_111 N_A_c_148_n N_VPWR_M1005_d 0.00546612f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_c_149_n N_VPWR_c_179_n 0.00763033f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_c_147_n N_VPWR_c_179_n 0.00270937f $X=1.965 $Y=1.202 $X2=0 $Y2=0
cc_114 N_A_c_148_n N_VPWR_c_179_n 0.0197361f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_c_149_n N_VPWR_c_180_n 0.00702461f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A_c_149_n N_VPWR_c_174_n 0.0137658f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A_c_146_n N_Y_c_214_n 0.0095216f $X=1.94 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A_c_149_n N_Y_c_214_n 0.00214305f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_c_147_n N_Y_c_214_n 0.0113334f $X=1.965 $Y=1.202 $X2=0 $Y2=0
cc_120 N_A_c_148_n N_Y_c_214_n 0.0298244f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_c_149_n N_Y_c_232_n 0.0062681f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A_c_148_n N_Y_c_232_n 0.0113746f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A_c_146_n N_Y_c_215_n 0.0187964f $X=1.94 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A_c_147_n N_Y_c_215_n 0.00751301f $X=1.965 $Y=1.202 $X2=0 $Y2=0
cc_125 N_A_c_148_n N_Y_c_215_n 0.0206713f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A_c_146_n N_VGND_c_262_n 0.00357668f $X=1.94 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_c_146_n N_VGND_c_263_n 0.00683541f $X=1.94 $Y=0.995 $X2=0 $Y2=0
cc_128 N_VPWR_c_174_n N_Y_M1004_d 0.00231261f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_129 N_VPWR_c_174_n N_Y_M1007_d 0.00348872f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_130 N_VPWR_c_176_n N_Y_c_217_n 0.013769f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_131 N_VPWR_c_176_n N_Y_c_218_n 0.0615942f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_132 N_VPWR_c_177_n N_Y_c_218_n 0.0223557f $X=1.115 $Y=2.72 $X2=0 $Y2=0
cc_133 N_VPWR_c_178_n N_Y_c_218_n 0.0385613f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_134 N_VPWR_c_174_n N_Y_c_218_n 0.0140101f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_135 N_VPWR_M1000_d N_Y_c_222_n 0.00495589f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_136 N_VPWR_c_178_n N_Y_c_222_n 0.0136682f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_137 N_VPWR_c_180_n N_Y_c_254_n 0.0198599f $X=2.115 $Y=2.72 $X2=0 $Y2=0
cc_138 N_VPWR_c_174_n N_Y_c_254_n 0.0126319f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_139 N_VPWR_c_176_n N_VGND_c_261_n 7.14544e-19 $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_140 N_Y_c_215_n N_VGND_c_262_n 0.0475266f $X=2.2 $Y=0.38 $X2=0 $Y2=0
cc_141 N_Y_M1002_d N_VGND_c_263_n 0.00283101f $X=2.015 $Y=0.235 $X2=0 $Y2=0
cc_142 N_Y_c_215_n N_VGND_c_263_n 0.0277553f $X=2.2 $Y=0.38 $X2=0 $Y2=0
cc_143 N_Y_c_215_n A_297_47# 0.00989808f $X=2.2 $Y=0.38 $X2=-0.19 $Y2=-0.24
cc_144 N_VGND_c_263_n A_119_47# 0.00453305f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24
cc_145 N_VGND_c_263_n A_213_47# 0.00219624f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24
cc_146 N_VGND_c_263_n A_297_47# 0.00950848f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24
