* File: sky130_fd_sc_hdll__nand4b_4.pex.spice
* Created: Wed Sep  2 08:38:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND4B_4%A_N 1 3 6 8 13
c30 8 0 1.24063e-19 $X=0.235 $Y=1.19
r31 13 14 3.61862 $w=3.33e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.212
+ $X2=0.52 $Y2=1.212
r32 11 13 31.8438 $w=3.33e-07 $l=2.2e-07 $layer=POLY_cond $X=0.275 $Y=1.212
+ $X2=0.495 $Y2=1.212
r33 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r34 4 14 21.4384 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=0.52 $Y=1.015
+ $X2=0.52 $Y2=1.212
r35 4 6 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.52 $Y=1.015
+ $X2=0.52 $Y2=0.56
r36 1 13 17.1428 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.212
r37 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_4%A_27_47# 1 2 9 11 14 16 18 21 23 25 28 30
+ 32 35 39 41 43 45 46 47 50 52 55 60 61 68
c130 61 0 1.24063e-19 $X=1.485 $Y=1.217
c131 16 0 1.81354e-19 $X=1.955 $Y=1.41
r132 68 69 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=2.895 $Y=1.217
+ $X2=2.92 $Y2=1.217
r133 67 68 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=2.45 $Y=1.217
+ $X2=2.895 $Y2=1.217
r134 66 67 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=2.425 $Y=1.217
+ $X2=2.45 $Y2=1.217
r135 65 66 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=1.98 $Y=1.217
+ $X2=2.425 $Y2=1.217
r136 64 65 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=1.955 $Y=1.217
+ $X2=1.98 $Y2=1.217
r137 61 62 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=1.485 $Y=1.217
+ $X2=1.51 $Y2=1.217
r138 56 64 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=1.72 $Y=1.217
+ $X2=1.955 $Y2=1.217
r139 56 62 30.9541 $w=3.27e-07 $l=2.1e-07 $layer=POLY_cond $X=1.72 $Y=1.217
+ $X2=1.51 $Y2=1.217
r140 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.72
+ $Y=1.16 $X2=1.72 $Y2=1.16
r141 53 60 1.25155 $w=2e-07 $l=9.8e-08 $layer=LI1_cond $X=0.855 $Y=1.175
+ $X2=0.757 $Y2=1.175
r142 53 55 47.9682 $w=1.98e-07 $l=8.65e-07 $layer=LI1_cond $X=0.855 $Y=1.175
+ $X2=1.72 $Y2=1.175
r143 51 60 5.27577 $w=1.95e-07 $l=1e-07 $layer=LI1_cond $X=0.757 $Y=1.275
+ $X2=0.757 $Y2=1.175
r144 51 52 12.5128 $w=1.93e-07 $l=2.2e-07 $layer=LI1_cond $X=0.757 $Y=1.275
+ $X2=0.757 $Y2=1.495
r145 50 60 5.27577 $w=1.95e-07 $l=1e-07 $layer=LI1_cond $X=0.757 $Y=1.075
+ $X2=0.757 $Y2=1.175
r146 49 50 9.669 $w=1.93e-07 $l=1.7e-07 $layer=LI1_cond $X=0.757 $Y=0.905
+ $X2=0.757 $Y2=1.075
r147 48 59 5.18513 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.425 $Y=1.58
+ $X2=0.257 $Y2=1.58
r148 47 52 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=0.66 $Y=1.58
+ $X2=0.757 $Y2=1.495
r149 47 48 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.66 $Y=1.58
+ $X2=0.425 $Y2=1.58
r150 45 49 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=0.66 $Y=0.82
+ $X2=0.757 $Y2=0.905
r151 45 46 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.66 $Y=0.82
+ $X2=0.425 $Y2=0.82
r152 41 59 2.62343 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.257 $Y=1.665
+ $X2=0.257 $Y2=1.58
r153 41 43 23.2209 $w=3.33e-07 $l=6.75e-07 $layer=LI1_cond $X=0.257 $Y=1.665
+ $X2=0.257 $Y2=2.34
r154 37 46 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.425 $Y2=0.82
r155 37 39 12.2125 $w=3.33e-07 $l=3.55e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.257 $Y2=0.38
r156 33 69 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.92 $Y=1.025
+ $X2=2.92 $Y2=1.217
r157 33 35 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.92 $Y=1.025
+ $X2=2.92 $Y2=0.56
r158 30 68 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.217
r159 30 32 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.985
r160 26 67 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.45 $Y=1.025
+ $X2=2.45 $Y2=1.217
r161 26 28 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.45 $Y=1.025
+ $X2=2.45 $Y2=0.56
r162 23 66 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.217
r163 23 25 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.985
r164 19 65 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.98 $Y=1.025
+ $X2=1.98 $Y2=1.217
r165 19 21 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.98 $Y=1.025
+ $X2=1.98 $Y2=0.56
r166 16 64 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.217
r167 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.985
r168 12 62 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.51 $Y=1.025
+ $X2=1.51 $Y2=1.217
r169 12 14 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.51 $Y=1.025
+ $X2=1.51 $Y2=0.56
r170 9 61 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.217
r171 9 11 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.985
r172 2 59 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r173 2 43 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r174 1 39 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_4%B 1 3 6 8 10 13 15 17 20 22 24 27 29 30
+ 31 32 47 55 58 61 64
c80 1 0 1.59082e-19 $X=3.365 $Y=1.41
r81 47 49 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=4.8 $Y=1.212
+ $X2=4.825 $Y2=1.212
r82 46 47 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=4.775 $Y=1.212
+ $X2=4.8 $Y2=1.212
r83 45 46 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=4.33 $Y=1.212
+ $X2=4.775 $Y2=1.212
r84 44 45 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=4.305 $Y=1.212
+ $X2=4.33 $Y2=1.212
r85 43 44 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=3.86 $Y=1.212
+ $X2=4.305 $Y2=1.212
r86 42 43 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=3.835 $Y=1.212
+ $X2=3.86 $Y2=1.212
r87 41 42 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=3.39 $Y=1.212
+ $X2=3.835 $Y2=1.212
r88 39 41 2.99379 $w=3.22e-07 $l=2e-08 $layer=POLY_cond $X=3.37 $Y=1.212
+ $X2=3.39 $Y2=1.212
r89 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.37
+ $Y=1.16 $X2=3.37 $Y2=1.16
r90 37 39 0.748447 $w=3.22e-07 $l=5e-09 $layer=POLY_cond $X=3.365 $Y=1.212
+ $X2=3.37 $Y2=1.212
r91 32 64 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=4.825 $Y=1.175
+ $X2=4.84 $Y2=1.175
r92 32 61 23.8455 $w=1.98e-07 $l=4.3e-07 $layer=LI1_cond $X=4.825 $Y=1.175
+ $X2=4.395 $Y2=1.175
r93 32 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.825
+ $Y=1.16 $X2=4.825 $Y2=1.16
r94 31 61 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=4.375 $Y=1.175
+ $X2=4.395 $Y2=1.175
r95 31 58 24.4 $w=1.98e-07 $l=4.4e-07 $layer=LI1_cond $X=4.375 $Y=1.175
+ $X2=3.935 $Y2=1.175
r96 30 58 1.66364 $w=1.98e-07 $l=3e-08 $layer=LI1_cond $X=3.905 $Y=1.175
+ $X2=3.935 $Y2=1.175
r97 30 55 23.8455 $w=1.98e-07 $l=4.3e-07 $layer=LI1_cond $X=3.905 $Y=1.175
+ $X2=3.475 $Y2=1.175
r98 29 55 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=3.47 $Y=1.175
+ $X2=3.475 $Y2=1.175
r99 29 40 5.54545 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=3.47 $Y=1.175 $X2=3.37
+ $Y2=1.175
r100 25 47 20.6399 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=4.8 $Y=1.015
+ $X2=4.8 $Y2=1.212
r101 25 27 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.8 $Y=1.015
+ $X2=4.8 $Y2=0.56
r102 22 46 16.3606 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.212
r103 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
r104 18 45 20.6399 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=4.33 $Y=1.025
+ $X2=4.33 $Y2=1.212
r105 18 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.33 $Y=1.025
+ $X2=4.33 $Y2=0.56
r106 15 44 16.3606 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.212
r107 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.985
r108 11 43 20.6399 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=3.86 $Y=1.025
+ $X2=3.86 $Y2=1.212
r109 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.86 $Y=1.025
+ $X2=3.86 $Y2=0.56
r110 8 42 16.3606 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.212
r111 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.985
r112 4 41 20.6399 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=3.39 $Y=1.025
+ $X2=3.39 $Y2=1.212
r113 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.39 $Y=1.025
+ $X2=3.39 $Y2=0.56
r114 1 37 16.3606 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.212
r115 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_4%C 1 3 6 8 10 13 15 17 20 22 24 27 29 30
+ 31 32 37 50 51 56 59 62 65
c80 27 0 3.89631e-19 $X=7.2 $Y=0.56
r81 51 52 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=7.175 $Y=1.217
+ $X2=7.2 $Y2=1.217
r82 49 51 33.9021 $w=3.27e-07 $l=2.3e-07 $layer=POLY_cond $X=6.945 $Y=1.217
+ $X2=7.175 $Y2=1.217
r83 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.945
+ $Y=1.16 $X2=6.945 $Y2=1.16
r84 47 49 31.6911 $w=3.27e-07 $l=2.15e-07 $layer=POLY_cond $X=6.73 $Y=1.217
+ $X2=6.945 $Y2=1.217
r85 46 47 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=6.705 $Y=1.217
+ $X2=6.73 $Y2=1.217
r86 45 46 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=6.26 $Y=1.217
+ $X2=6.705 $Y2=1.217
r87 44 45 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=6.235 $Y=1.217
+ $X2=6.26 $Y2=1.217
r88 43 44 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=5.79 $Y=1.217
+ $X2=6.235 $Y2=1.217
r89 42 43 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=5.765 $Y=1.217
+ $X2=5.79 $Y2=1.217
r90 40 59 19.9636 $w=1.98e-07 $l=3.6e-07 $layer=LI1_cond $X=5.435 $Y=1.175
+ $X2=5.795 $Y2=1.175
r91 40 56 5.54545 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=5.435 $Y=1.175
+ $X2=5.335 $Y2=1.175
r92 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.435
+ $Y=1.16 $X2=5.435 $Y2=1.16
r93 37 42 16.3472 $w=3.27e-07 $l=1.253e-07 $layer=POLY_cond $X=5.665 $Y=1.16
+ $X2=5.765 $Y2=1.217
r94 37 39 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=5.665 $Y=1.16 $X2=5.435
+ $Y2=1.16
r95 32 50 11.6455 $w=1.98e-07 $l=2.1e-07 $layer=LI1_cond $X=6.735 $Y=1.175
+ $X2=6.945 $Y2=1.175
r96 32 65 2.77273 $w=1.98e-07 $l=5e-08 $layer=LI1_cond $X=6.735 $Y=1.175
+ $X2=6.685 $Y2=1.175
r97 31 65 20.2409 $w=1.98e-07 $l=3.65e-07 $layer=LI1_cond $X=6.32 $Y=1.175
+ $X2=6.685 $Y2=1.175
r98 31 62 3.60455 $w=1.98e-07 $l=6.5e-08 $layer=LI1_cond $X=6.32 $Y=1.175
+ $X2=6.255 $Y2=1.175
r99 30 62 24.6773 $w=1.98e-07 $l=4.45e-07 $layer=LI1_cond $X=5.81 $Y=1.175
+ $X2=6.255 $Y2=1.175
r100 30 59 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=5.81 $Y=1.175
+ $X2=5.795 $Y2=1.175
r101 29 56 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=5.325 $Y=1.175
+ $X2=5.335 $Y2=1.175
r102 25 52 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.2 $Y=1.025
+ $X2=7.2 $Y2=1.217
r103 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.2 $Y=1.025
+ $X2=7.2 $Y2=0.56
r104 22 51 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.175 $Y=1.41
+ $X2=7.175 $Y2=1.217
r105 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.175 $Y=1.41
+ $X2=7.175 $Y2=1.985
r106 18 47 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.73 $Y=1.025
+ $X2=6.73 $Y2=1.217
r107 18 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.73 $Y=1.025
+ $X2=6.73 $Y2=0.56
r108 15 46 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.705 $Y=1.41
+ $X2=6.705 $Y2=1.217
r109 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.705 $Y=1.41
+ $X2=6.705 $Y2=1.985
r110 11 45 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.26 $Y=1.025
+ $X2=6.26 $Y2=1.217
r111 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.26 $Y=1.025
+ $X2=6.26 $Y2=0.56
r112 8 44 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.235 $Y=1.41
+ $X2=6.235 $Y2=1.217
r113 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.235 $Y=1.41
+ $X2=6.235 $Y2=1.985
r114 4 43 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.79 $Y=1.025
+ $X2=5.79 $Y2=1.217
r115 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.79 $Y=1.025
+ $X2=5.79 $Y2=0.56
r116 1 42 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.765 $Y=1.41
+ $X2=5.765 $Y2=1.217
r117 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.765 $Y=1.41
+ $X2=5.765 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_4%D 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 32 37 39 57 60 63 66
r88 51 52 3.67378 $w=3.28e-07 $l=2.5e-08 $layer=POLY_cond $X=9.03 $Y=1.212
+ $X2=9.055 $Y2=1.212
r89 50 51 65.3933 $w=3.28e-07 $l=4.45e-07 $layer=POLY_cond $X=8.585 $Y=1.212
+ $X2=9.03 $Y2=1.212
r90 49 50 3.67378 $w=3.28e-07 $l=2.5e-08 $layer=POLY_cond $X=8.56 $Y=1.212
+ $X2=8.585 $Y2=1.212
r91 48 49 65.3933 $w=3.28e-07 $l=4.45e-07 $layer=POLY_cond $X=8.115 $Y=1.212
+ $X2=8.56 $Y2=1.212
r92 47 48 3.67378 $w=3.28e-07 $l=2.5e-08 $layer=POLY_cond $X=8.09 $Y=1.212
+ $X2=8.115 $Y2=1.212
r93 45 47 30.8598 $w=3.28e-07 $l=2.1e-07 $layer=POLY_cond $X=7.88 $Y=1.212
+ $X2=8.09 $Y2=1.212
r94 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.88
+ $Y=1.16 $X2=7.88 $Y2=1.16
r95 43 45 34.5335 $w=3.28e-07 $l=2.35e-07 $layer=POLY_cond $X=7.645 $Y=1.212
+ $X2=7.88 $Y2=1.212
r96 42 43 3.67378 $w=3.28e-07 $l=2.5e-08 $layer=POLY_cond $X=7.62 $Y=1.212
+ $X2=7.645 $Y2=1.212
r97 37 52 15.4609 $w=3.28e-07 $l=1.23288e-07 $layer=POLY_cond $X=9.155 $Y=1.16
+ $X2=9.055 $Y2=1.212
r98 37 39 34.1305 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=9.155 $Y=1.16
+ $X2=9.32 $Y2=1.16
r99 32 66 3.88182 $w=1.98e-07 $l=7e-08 $layer=LI1_cond $X=9.32 $Y=1.175 $X2=9.39
+ $Y2=1.175
r100 32 63 23.0136 $w=1.98e-07 $l=4.15e-07 $layer=LI1_cond $X=9.32 $Y=1.175
+ $X2=8.905 $Y2=1.175
r101 32 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.32
+ $Y=1.16 $X2=9.32 $Y2=1.16
r102 31 63 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=8.895 $Y=1.175
+ $X2=8.905 $Y2=1.175
r103 31 60 21.35 $w=1.98e-07 $l=3.85e-07 $layer=LI1_cond $X=8.895 $Y=1.175
+ $X2=8.51 $Y2=1.175
r104 30 60 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=8.5 $Y=1.175
+ $X2=8.51 $Y2=1.175
r105 30 57 22.4591 $w=1.98e-07 $l=4.05e-07 $layer=LI1_cond $X=8.5 $Y=1.175
+ $X2=8.095 $Y2=1.175
r106 29 57 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=8.055 $Y=1.175
+ $X2=8.095 $Y2=1.175
r107 29 46 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=8.055 $Y=1.175
+ $X2=7.88 $Y2=1.175
r108 26 52 16.7902 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=9.055 $Y=1.41
+ $X2=9.055 $Y2=1.212
r109 26 28 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.055 $Y=1.41
+ $X2=9.055 $Y2=1.985
r110 22 51 21.0783 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=9.03 $Y=1.015
+ $X2=9.03 $Y2=1.212
r111 22 24 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=9.03 $Y=1.015
+ $X2=9.03 $Y2=0.56
r112 19 50 16.7902 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=8.585 $Y=1.41
+ $X2=8.585 $Y2=1.212
r113 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.585 $Y=1.41
+ $X2=8.585 $Y2=1.985
r114 15 49 21.0783 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=8.56 $Y=1.025
+ $X2=8.56 $Y2=1.212
r115 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.56 $Y=1.025
+ $X2=8.56 $Y2=0.56
r116 12 48 16.7902 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=8.115 $Y=1.41
+ $X2=8.115 $Y2=1.212
r117 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.115 $Y=1.41
+ $X2=8.115 $Y2=1.985
r118 8 47 21.0783 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=8.09 $Y=1.025
+ $X2=8.09 $Y2=1.212
r119 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.09 $Y=1.025
+ $X2=8.09 $Y2=0.56
r120 5 43 16.7902 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=7.645 $Y=1.41
+ $X2=7.645 $Y2=1.212
r121 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.645 $Y=1.41
+ $X2=7.645 $Y2=1.985
r122 1 42 21.0783 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=7.62 $Y=1.025
+ $X2=7.62 $Y2=1.212
r123 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.62 $Y=1.025
+ $X2=7.62 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_4%VPWR 1 2 3 4 5 6 7 8 9 10 36 39 43 47 51
+ 55 59 63 67 69 71 76 79 80 82 83 85 86 88 89 91 92 94 95 96 108 122 127 132
+ 136
r152 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r153 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r154 128 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r155 127 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r156 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r157 125 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.43 $Y2=2.72
r158 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r159 122 135 3.95444 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=9.205 $Y=2.72
+ $X2=9.432 $Y2=2.72
r160 122 124 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.205 $Y=2.72
+ $X2=8.97 $Y2=2.72
r161 121 125 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r162 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r163 118 121 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r164 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r165 115 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r166 115 133 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.29 $Y2=2.72
r167 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r168 112 132 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=5.615 $Y=2.72
+ $X2=5.27 $Y2=2.72
r169 112 114 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.615 $Y=2.72
+ $X2=6.21 $Y2=2.72
r170 111 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r171 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r172 108 132 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=4.925 $Y=2.72
+ $X2=5.27 $Y2=2.72
r173 108 110 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.925 $Y=2.72
+ $X2=4.83 $Y2=2.72
r174 107 111 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r175 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r176 104 107 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r177 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r178 101 104 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r179 101 128 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r180 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r181 98 127 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=0.99 $Y2=2.72
r182 98 100 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=2.07 $Y2=2.72
r183 96 130 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r184 94 120 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=8.265 $Y=2.72
+ $X2=8.05 $Y2=2.72
r185 94 95 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.265 $Y=2.72
+ $X2=8.35 $Y2=2.72
r186 93 124 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=8.435 $Y=2.72
+ $X2=8.97 $Y2=2.72
r187 93 95 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.435 $Y=2.72
+ $X2=8.35 $Y2=2.72
r188 91 117 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.325 $Y=2.72
+ $X2=7.13 $Y2=2.72
r189 91 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.325 $Y=2.72
+ $X2=7.41 $Y2=2.72
r190 90 120 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=7.495 $Y=2.72
+ $X2=8.05 $Y2=2.72
r191 90 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.495 $Y=2.72
+ $X2=7.41 $Y2=2.72
r192 88 114 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.385 $Y=2.72
+ $X2=6.21 $Y2=2.72
r193 88 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.385 $Y=2.72
+ $X2=6.47 $Y2=2.72
r194 87 117 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.555 $Y=2.72
+ $X2=7.13 $Y2=2.72
r195 87 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=2.72
+ $X2=6.47 $Y2=2.72
r196 85 106 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.985 $Y=2.72
+ $X2=3.91 $Y2=2.72
r197 85 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.985 $Y=2.72
+ $X2=4.07 $Y2=2.72
r198 84 110 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=4.155 $Y=2.72
+ $X2=4.83 $Y2=2.72
r199 84 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=2.72
+ $X2=4.07 $Y2=2.72
r200 82 103 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.045 $Y=2.72
+ $X2=2.99 $Y2=2.72
r201 82 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.045 $Y=2.72
+ $X2=3.13 $Y2=2.72
r202 81 106 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=3.91 $Y2=2.72
r203 81 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=3.13 $Y2=2.72
r204 79 100 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.07 $Y2=2.72
r205 79 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.19 $Y2=2.72
r206 78 103 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.99 $Y2=2.72
r207 78 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.19 $Y2=2.72
r208 76 77 6.97577 $w=6.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=2 $X2=0.99
+ $Y2=1.835
r209 71 74 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=9.332 $Y=1.66
+ $X2=9.332 $Y2=2.34
r210 69 135 3.22278 $w=2.55e-07 $l=1.36015e-07 $layer=LI1_cond $X=9.332 $Y=2.635
+ $X2=9.432 $Y2=2.72
r211 69 74 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=9.332 $Y=2.635
+ $X2=9.332 $Y2=2.34
r212 65 95 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.35 $Y=2.635
+ $X2=8.35 $Y2=2.72
r213 65 67 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.35 $Y=2.635
+ $X2=8.35 $Y2=2
r214 61 92 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.41 $Y=2.635
+ $X2=7.41 $Y2=2.72
r215 61 63 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.41 $Y=2.635
+ $X2=7.41 $Y2=2
r216 57 89 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=2.635
+ $X2=6.47 $Y2=2.72
r217 57 59 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.47 $Y=2.635
+ $X2=6.47 $Y2=2
r218 53 132 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.27 $Y=2.635
+ $X2=5.27 $Y2=2.72
r219 53 55 11.0074 $w=6.88e-07 $l=6.35e-07 $layer=LI1_cond $X=5.27 $Y=2.635
+ $X2=5.27 $Y2=2
r220 49 86 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=2.635
+ $X2=4.07 $Y2=2.72
r221 49 51 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.07 $Y=2.635
+ $X2=4.07 $Y2=2
r222 45 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=2.635
+ $X2=3.13 $Y2=2.72
r223 45 47 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.13 $Y=2.635
+ $X2=3.13 $Y2=2
r224 41 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2.72
r225 41 43 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2
r226 39 77 6.9544 $w=2.88e-07 $l=1.75e-07 $layer=LI1_cond $X=1.19 $Y=1.66
+ $X2=1.19 $Y2=1.835
r227 34 127 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.99 $Y=2.635
+ $X2=0.99 $Y2=2.72
r228 34 36 5.11367 $w=6.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.99 $Y=2.635
+ $X2=0.99 $Y2=2.34
r229 33 76 3.1202 $w=6.88e-07 $l=1.8e-07 $layer=LI1_cond $X=0.99 $Y=2.18
+ $X2=0.99 $Y2=2
r230 33 36 2.77352 $w=6.88e-07 $l=1.6e-07 $layer=LI1_cond $X=0.99 $Y=2.18
+ $X2=0.99 $Y2=2.34
r231 10 74 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=9.145
+ $Y=1.485 $X2=9.29 $Y2=2.34
r232 10 71 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=9.145
+ $Y=1.485 $X2=9.29 $Y2=1.66
r233 9 67 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=8.205
+ $Y=1.485 $X2=8.35 $Y2=2
r234 8 63 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=7.265
+ $Y=1.485 $X2=7.41 $Y2=2
r235 7 59 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.325
+ $Y=1.485 $X2=6.47 $Y2=2
r236 6 55 150 $w=1.7e-07 $l=8.02185e-07 $layer=licon1_PDIFF $count=4 $X=4.865
+ $Y=1.485 $X2=5.45 $Y2=2
r237 5 51 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=2
r238 4 47 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.985
+ $Y=1.485 $X2=3.13 $Y2=2
r239 3 43 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=1.485 $X2=2.19 $Y2=2
r240 2 39 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.25 $Y2=1.66
r241 2 36 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.25 $Y2=2.34
r242 1 76 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_4%Y 1 2 3 4 5 6 7 8 9 10 31 35 37 39 43 47
+ 49 53 55 59 61 65 67 71 73 75 77 81 83 85 87 89 91 94 95 96 103
c192 103 0 1.62009e-19 $X=2.625 $Y=0.905
c193 94 0 3.40437e-19 $X=2.745 $Y=0.85
r194 95 96 6.06193 $w=5.98e-07 $l=2.55e-07 $layer=LI1_cond $X=2.625 $Y=1.19
+ $X2=2.625 $Y2=1.445
r195 94 103 2.81193 $w=4.3e-07 $l=1.35e-07 $layer=LI1_cond $X=2.625 $Y=0.77
+ $X2=2.625 $Y2=0.905
r196 94 95 7.23627 $w=4.28e-07 $l=2.7e-07 $layer=LI1_cond $X=2.625 $Y=0.92
+ $X2=2.625 $Y2=1.19
r197 94 103 0.402015 $w=4.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.625 $Y=0.92
+ $X2=2.625 $Y2=0.905
r198 81 96 17.3778 $w=3.88e-07 $l=5.45e-07 $layer=LI1_cond $X=3.385 $Y=1.555
+ $X2=2.84 $Y2=1.555
r199 81 83 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=3.385 $Y=1.555
+ $X2=3.575 $Y2=1.555
r200 75 93 2.73777 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=8.795 $Y=1.665
+ $X2=8.795 $Y2=1.555
r201 75 77 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=8.795 $Y=1.665
+ $X2=8.795 $Y2=2.34
r202 74 91 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=8.045 $Y=1.555
+ $X2=7.855 $Y2=1.555
r203 73 93 4.72888 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=8.605 $Y=1.555
+ $X2=8.795 $Y2=1.555
r204 73 74 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=8.605 $Y=1.555
+ $X2=8.045 $Y2=1.555
r205 69 91 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=7.855 $Y=1.665
+ $X2=7.855 $Y2=1.555
r206 69 71 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=7.855 $Y=1.665
+ $X2=7.855 $Y2=2.34
r207 68 89 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=7.105 $Y=1.555
+ $X2=6.915 $Y2=1.555
r208 67 91 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=7.665 $Y=1.555
+ $X2=7.855 $Y2=1.555
r209 67 68 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=7.665 $Y=1.555
+ $X2=7.105 $Y2=1.555
r210 63 89 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=6.915 $Y=1.665
+ $X2=6.915 $Y2=1.555
r211 63 65 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=6.915 $Y=1.665
+ $X2=6.915 $Y2=2.34
r212 62 87 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=6.165 $Y=1.555
+ $X2=5.975 $Y2=1.555
r213 61 89 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=6.725 $Y=1.555
+ $X2=6.915 $Y2=1.555
r214 61 62 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=6.725 $Y=1.555
+ $X2=6.165 $Y2=1.555
r215 57 87 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=5.975 $Y=1.665
+ $X2=5.975 $Y2=1.555
r216 57 59 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=5.975 $Y=1.665
+ $X2=5.975 $Y2=2.34
r217 56 85 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=4.705 $Y=1.555
+ $X2=4.515 $Y2=1.555
r218 55 87 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=5.785 $Y=1.555
+ $X2=5.975 $Y2=1.555
r219 55 56 56.5745 $w=2.18e-07 $l=1.08e-06 $layer=LI1_cond $X=5.785 $Y=1.555
+ $X2=4.705 $Y2=1.555
r220 51 85 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=4.515 $Y=1.665
+ $X2=4.515 $Y2=1.555
r221 51 53 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=4.515 $Y=1.665
+ $X2=4.515 $Y2=2.34
r222 50 83 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=3.765 $Y=1.555
+ $X2=3.575 $Y2=1.555
r223 49 85 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=4.325 $Y=1.555
+ $X2=4.515 $Y2=1.555
r224 49 50 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=4.325 $Y=1.555
+ $X2=3.765 $Y2=1.555
r225 45 83 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=3.575 $Y=1.665
+ $X2=3.575 $Y2=1.555
r226 45 47 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=3.575 $Y=1.665
+ $X2=3.575 $Y2=2.34
r227 41 96 1.42006 $w=3.8e-07 $l=1.14891e-07 $layer=LI1_cond $X=2.635 $Y=1.665
+ $X2=2.625 $Y2=1.555
r228 41 43 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=2.635 $Y=1.665
+ $X2=2.635 $Y2=2.34
r229 40 80 4.72888 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.885 $Y=1.555
+ $X2=1.695 $Y2=1.555
r230 39 96 5.08349 $w=2.2e-07 $l=2.15e-07 $layer=LI1_cond $X=2.41 $Y=1.555
+ $X2=2.625 $Y2=1.555
r231 39 40 27.5015 $w=2.18e-07 $l=5.25e-07 $layer=LI1_cond $X=2.41 $Y=1.555
+ $X2=1.885 $Y2=1.555
r232 35 80 2.73777 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=1.555
r233 35 37 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=2.34
r234 31 94 4.47825 $w=2.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.41 $Y=0.77
+ $X2=2.625 $Y2=0.77
r235 31 33 29.4513 $w=2.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.41 $Y=0.77
+ $X2=1.72 $Y2=0.77
r236 10 93 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=8.675
+ $Y=1.485 $X2=8.82 $Y2=1.66
r237 10 77 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=8.675
+ $Y=1.485 $X2=8.82 $Y2=2.34
r238 9 91 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=7.735
+ $Y=1.485 $X2=7.88 $Y2=1.66
r239 9 71 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.735
+ $Y=1.485 $X2=7.88 $Y2=2.34
r240 8 89 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=6.795
+ $Y=1.485 $X2=6.94 $Y2=1.66
r241 8 65 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.795
+ $Y=1.485 $X2=6.94 $Y2=2.34
r242 7 87 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.855
+ $Y=1.485 $X2=6 $Y2=1.66
r243 7 59 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.855
+ $Y=1.485 $X2=6 $Y2=2.34
r244 6 85 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.485 $X2=4.54 $Y2=1.66
r245 6 53 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.485 $X2=4.54 $Y2=2.34
r246 5 83 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.455
+ $Y=1.485 $X2=3.6 $Y2=1.66
r247 5 47 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.455
+ $Y=1.485 $X2=3.6 $Y2=2.34
r248 4 96 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=1.485 $X2=2.66 $Y2=1.66
r249 4 43 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=1.485 $X2=2.66 $Y2=2.34
r250 3 80 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=1.485 $X2=1.72 $Y2=1.66
r251 3 37 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=1.485 $X2=1.72 $Y2=2.34
r252 2 94 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.525
+ $Y=0.235 $X2=2.66 $Y2=0.72
r253 1 33 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.235 $X2=1.72 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_4%VGND 1 2 3 14 18 22 25 26 28 29 30 43 44
+ 47
r103 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r104 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r105 41 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=9.43
+ $Y2=0
r106 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r107 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.51
+ $Y2=0
r108 37 38 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r109 35 38 1.83245 $w=4.8e-07 $l=6.44e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=7.59
+ $Y2=0
r110 35 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r111 34 37 420.15 $w=1.68e-07 $l=6.44e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=7.59
+ $Y2=0
r112 34 35 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r113 32 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.77
+ $Y2=0
r114 32 34 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r115 30 48 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r116 28 40 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=8.735 $Y=0
+ $X2=8.51 $Y2=0
r117 28 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.735 $Y=0 $X2=8.82
+ $Y2=0
r118 27 43 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=8.905 $Y=0
+ $X2=9.43 $Y2=0
r119 27 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.905 $Y=0 $X2=8.82
+ $Y2=0
r120 25 37 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.795 $Y=0
+ $X2=7.59 $Y2=0
r121 25 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.795 $Y=0 $X2=7.88
+ $Y2=0
r122 24 40 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=7.965 $Y=0
+ $X2=8.51 $Y2=0
r123 24 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.965 $Y=0 $X2=7.88
+ $Y2=0
r124 20 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.82 $Y=0.085
+ $X2=8.82 $Y2=0
r125 20 22 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.82 $Y=0.085
+ $X2=8.82 $Y2=0.38
r126 16 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.88 $Y=0.085
+ $X2=7.88 $Y2=0
r127 16 18 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.88 $Y=0.085
+ $X2=7.88 $Y2=0.38
r128 12 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=0.085
+ $X2=0.77 $Y2=0
r129 12 14 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.77 $Y=0.085
+ $X2=0.77 $Y2=0.38
r130 3 22 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=8.635
+ $Y=0.235 $X2=8.82 $Y2=0.38
r131 2 18 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=7.695
+ $Y=0.235 $X2=7.88 $Y2=0.38
r132 1 14 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_4%A_225_47# 1 2 3 4 5 16 18 28
r44 26 28 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=4.07 $Y=0.36 $X2=5.01
+ $Y2=0.36
r45 24 26 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=3.13 $Y=0.36 $X2=4.07
+ $Y2=0.36
r46 22 24 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=2.19 $Y=0.36 $X2=3.13
+ $Y2=0.36
r47 20 31 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.335 $Y=0.36
+ $X2=1.21 $Y2=0.36
r48 20 22 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=1.335 $Y=0.36
+ $X2=2.19 $Y2=0.36
r49 16 31 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.21 $Y=0.465
+ $X2=1.21 $Y2=0.36
r50 16 18 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=1.21 $Y=0.465
+ $X2=1.21 $Y2=0.72
r51 5 28 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.875
+ $Y=0.235 $X2=5.01 $Y2=0.38
r52 4 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.935
+ $Y=0.235 $X2=4.07 $Y2=0.38
r53 3 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.995
+ $Y=0.235 $X2=3.13 $Y2=0.38
r54 2 22 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.055
+ $Y=0.235 $X2=2.19 $Y2=0.38
r55 1 31 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.25 $Y2=0.38
r56 1 18 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.25 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_4%A_693_47# 1 2 3 4 21
c33 21 0 1.91072e-19 $X=6.94 $Y=0.72
r34 19 21 40.1221 $w=2.68e-07 $l=9.4e-07 $layer=LI1_cond $X=6 $Y=0.77 $X2=6.94
+ $Y2=0.77
r35 17 19 62.3173 $w=2.68e-07 $l=1.46e-06 $layer=LI1_cond $X=4.54 $Y=0.77 $X2=6
+ $Y2=0.77
r36 14 17 40.1221 $w=2.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.6 $Y=0.77 $X2=4.54
+ $Y2=0.77
r37 4 21 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=6.805
+ $Y=0.235 $X2=6.94 $Y2=0.72
r38 3 19 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=5.865
+ $Y=0.235 $X2=6 $Y2=0.72
r39 2 17 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=4.405
+ $Y=0.235 $X2=4.54 $Y2=0.72
r40 1 14 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.465
+ $Y=0.235 $X2=3.6 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4B_4%A_1081_47# 1 2 3 4 5 16 22 25 26 27 30 32
+ 36 40
c67 27 0 1.98558e-19 $X=7.575 $Y=0.82
r68 34 36 10.6264 $w=3.83e-07 $l=3.55e-07 $layer=LI1_cond $X=9.267 $Y=0.735
+ $X2=9.267 $Y2=0.38
r69 33 40 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.515 $Y=0.82
+ $X2=8.325 $Y2=0.82
r70 32 34 8.24022 $w=1.7e-07 $l=2.30617e-07 $layer=LI1_cond $X=9.075 $Y=0.82
+ $X2=9.267 $Y2=0.735
r71 32 33 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=9.075 $Y=0.82
+ $X2=8.515 $Y2=0.82
r72 28 40 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.325 $Y=0.735
+ $X2=8.325 $Y2=0.82
r73 28 30 10.7662 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=8.325 $Y=0.735
+ $X2=8.325 $Y2=0.38
r74 26 40 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.135 $Y=0.82
+ $X2=8.325 $Y2=0.82
r75 26 27 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.135 $Y=0.82
+ $X2=7.575 $Y2=0.82
r76 23 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.45 $Y=0.735
+ $X2=7.575 $Y2=0.82
r77 23 25 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=7.45 $Y=0.735
+ $X2=7.45 $Y2=0.72
r78 22 39 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=7.45 $Y=0.465
+ $X2=7.45 $Y2=0.36
r79 22 25 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=7.45 $Y=0.465
+ $X2=7.45 $Y2=0.72
r80 18 21 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=5.53 $Y=0.36 $X2=6.47
+ $Y2=0.36
r81 16 39 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=7.325 $Y=0.36
+ $X2=7.45 $Y2=0.36
r82 16 21 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=7.325 $Y=0.36
+ $X2=6.47 $Y2=0.36
r83 5 36 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=9.105
+ $Y=0.235 $X2=9.29 $Y2=0.38
r84 4 30 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=8.165
+ $Y=0.235 $X2=8.35 $Y2=0.38
r85 3 39 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.275
+ $Y=0.235 $X2=7.41 $Y2=0.38
r86 3 25 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=7.275
+ $Y=0.235 $X2=7.41 $Y2=0.72
r87 2 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.335
+ $Y=0.235 $X2=6.47 $Y2=0.38
r88 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.405
+ $Y=0.235 $X2=5.53 $Y2=0.38
.ends

