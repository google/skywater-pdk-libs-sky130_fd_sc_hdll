* File: sky130_fd_sc_hdll__nand2_16.pex.spice
* Created: Thu Aug 27 19:12:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND2_16%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 51 52 54 55 57 58 60 61
+ 63 64 66 67 69 70 72 73 75 76 78 79 81 82 84 85 87 88 90 91 93 94 96 97 134
+ 135
r328 135 136 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=7.545 $Y=1.202
+ $X2=7.57 $Y2=1.202
r329 133 135 24.297 $w=3.67e-07 $l=1.85e-07 $layer=POLY_cond $X=7.36 $Y=1.202
+ $X2=7.545 $Y2=1.202
r330 133 134 13.8362 $w=1.7e-07 $l=1.785e-06 $layer=licon1_POLY $count=10
+ $X=7.36 $Y=1.16 $X2=7.36 $Y2=1.16
r331 131 133 37.4305 $w=3.67e-07 $l=2.85e-07 $layer=POLY_cond $X=7.075 $Y=1.202
+ $X2=7.36 $Y2=1.202
r332 130 131 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=7.05 $Y=1.202
+ $X2=7.075 $Y2=1.202
r333 129 130 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=6.63 $Y=1.202
+ $X2=7.05 $Y2=1.202
r334 128 129 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=6.605 $Y=1.202
+ $X2=6.63 $Y2=1.202
r335 127 128 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=6.135 $Y=1.202
+ $X2=6.605 $Y2=1.202
r336 126 127 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=6.11 $Y=1.202
+ $X2=6.135 $Y2=1.202
r337 125 126 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=5.69 $Y=1.202
+ $X2=6.11 $Y2=1.202
r338 124 125 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=5.665 $Y=1.202
+ $X2=5.69 $Y2=1.202
r339 123 124 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=5.195 $Y=1.202
+ $X2=5.665 $Y2=1.202
r340 122 123 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=5.17 $Y=1.202
+ $X2=5.195 $Y2=1.202
r341 121 122 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=4.75 $Y=1.202
+ $X2=5.17 $Y2=1.202
r342 120 121 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=4.725 $Y=1.202
+ $X2=4.75 $Y2=1.202
r343 119 120 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=4.255 $Y=1.202
+ $X2=4.725 $Y2=1.202
r344 118 119 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=4.23 $Y=1.202
+ $X2=4.255 $Y2=1.202
r345 117 118 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=3.81 $Y=1.202
+ $X2=4.23 $Y2=1.202
r346 116 117 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=3.785 $Y=1.202
+ $X2=3.81 $Y2=1.202
r347 115 116 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=3.315 $Y=1.202
+ $X2=3.785 $Y2=1.202
r348 114 115 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.202
+ $X2=3.315 $Y2=1.202
r349 113 114 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=2.87 $Y=1.202
+ $X2=3.29 $Y2=1.202
r350 112 113 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=2.87 $Y2=1.202
r351 111 112 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.845 $Y2=1.202
r352 110 111 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.202
+ $X2=2.375 $Y2=1.202
r353 109 110 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=1.93 $Y=1.202
+ $X2=2.35 $Y2=1.202
r354 108 109 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=1.93 $Y2=1.202
r355 107 108 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.905 $Y2=1.202
r356 106 107 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.202
+ $X2=1.435 $Y2=1.202
r357 105 106 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=0.99 $Y=1.202
+ $X2=1.41 $Y2=1.202
r358 104 105 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r359 102 104 53.1907 $w=3.67e-07 $l=4.05e-07 $layer=POLY_cond $X=0.56 $Y=1.202
+ $X2=0.965 $Y2=1.202
r360 102 103 13.8362 $w=1.7e-07 $l=1.785e-06 $layer=licon1_POLY $count=10
+ $X=0.56 $Y=1.16 $X2=0.56 $Y2=1.16
r361 100 102 8.53679 $w=3.67e-07 $l=6.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.56 $Y2=1.202
r362 99 100 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r363 97 134 147.257 $w=2.68e-07 $l=3.45e-06 $layer=LI1_cond $X=3.91 $Y=1.19
+ $X2=7.36 $Y2=1.19
r364 97 103 142.988 $w=2.68e-07 $l=3.35e-06 $layer=LI1_cond $X=3.91 $Y=1.19
+ $X2=0.56 $Y2=1.19
r365 94 136 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.57 $Y=0.995
+ $X2=7.57 $Y2=1.202
r366 94 96 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.57 $Y=0.995
+ $X2=7.57 $Y2=0.56
r367 91 135 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.202
r368 91 93 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.985
r369 88 131 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.202
r370 88 90 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.985
r371 85 130 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.05 $Y=0.995
+ $X2=7.05 $Y2=1.202
r372 85 87 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.05 $Y=0.995
+ $X2=7.05 $Y2=0.56
r373 82 129 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=1.202
r374 82 84 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=0.56
r375 79 128 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.202
r376 79 81 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.985
r377 76 127 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.202
r378 76 78 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.985
r379 73 126 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.11 $Y=0.995
+ $X2=6.11 $Y2=1.202
r380 73 75 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.11 $Y=0.995
+ $X2=6.11 $Y2=0.56
r381 70 125 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=1.202
r382 70 72 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=0.56
r383 67 124 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.202
r384 67 69 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.985
r385 64 123 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.202
r386 64 66 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.985
r387 61 122 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.17 $Y=0.995
+ $X2=5.17 $Y2=1.202
r388 61 63 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.17 $Y=0.995
+ $X2=5.17 $Y2=0.56
r389 58 121 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.75 $Y=0.995
+ $X2=4.75 $Y2=1.202
r390 58 60 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.75 $Y=0.995
+ $X2=4.75 $Y2=0.56
r391 55 120 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.202
r392 55 57 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.985
r393 52 119 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.202
r394 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.985
r395 49 118 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.23 $Y=0.995
+ $X2=4.23 $Y2=1.202
r396 49 51 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.23 $Y=0.995
+ $X2=4.23 $Y2=0.56
r397 46 117 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=1.202
r398 46 48 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=0.56
r399 43 116 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.202
r400 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r401 40 115 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.202
r402 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r403 37 114 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=1.202
r404 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=0.56
r405 34 113 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.87 $Y=0.995
+ $X2=2.87 $Y2=1.202
r406 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.87 $Y=0.995
+ $X2=2.87 $Y2=0.56
r407 31 112 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r408 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r409 28 111 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r410 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r411 25 110 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.202
r412 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=0.56
r413 22 109 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r414 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r415 19 108 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r416 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r417 16 107 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r418 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r419 13 106 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.202
r420 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=0.56
r421 10 105 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r422 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r423 7 104 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r424 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r425 4 100 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r426 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r427 1 99 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.202
r428 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_16%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 51 52 54 55 57 58 60 61
+ 63 64 66 67 69 70 72 73 75 76 78 79 81 82 84 85 87 88 90 91 93 94 96 97 130
+ 135
r255 135 136 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=15.065 $Y=1.202
+ $X2=15.09 $Y2=1.202
r256 134 135 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=14.595 $Y=1.202
+ $X2=15.065 $Y2=1.202
r257 133 134 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=14.57 $Y=1.202
+ $X2=14.595 $Y2=1.202
r258 132 133 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=14.15 $Y=1.202
+ $X2=14.57 $Y2=1.202
r259 131 132 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=14.125 $Y=1.202
+ $X2=14.15 $Y2=1.202
r260 129 131 1.97003 $w=3.67e-07 $l=1.5e-08 $layer=POLY_cond $X=14.11 $Y=1.202
+ $X2=14.125 $Y2=1.202
r261 129 130 17.0918 $w=1.7e-07 $l=1.445e-06 $layer=licon1_POLY $count=8
+ $X=14.11 $Y=1.16 $X2=14.11 $Y2=1.16
r262 127 129 59.7575 $w=3.67e-07 $l=4.55e-07 $layer=POLY_cond $X=13.655 $Y=1.202
+ $X2=14.11 $Y2=1.202
r263 126 127 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=13.63 $Y=1.202
+ $X2=13.655 $Y2=1.202
r264 125 126 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=13.21 $Y=1.202
+ $X2=13.63 $Y2=1.202
r265 124 125 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=13.185 $Y=1.202
+ $X2=13.21 $Y2=1.202
r266 123 124 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=12.715 $Y=1.202
+ $X2=13.185 $Y2=1.202
r267 122 123 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=12.69 $Y=1.202
+ $X2=12.715 $Y2=1.202
r268 121 122 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=12.27 $Y=1.202
+ $X2=12.69 $Y2=1.202
r269 120 121 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=12.245 $Y=1.202
+ $X2=12.27 $Y2=1.202
r270 119 120 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=11.775 $Y=1.202
+ $X2=12.245 $Y2=1.202
r271 118 119 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=11.75 $Y=1.202
+ $X2=11.775 $Y2=1.202
r272 117 118 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=11.305 $Y=1.202
+ $X2=11.75 $Y2=1.202
r273 116 117 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=11.28 $Y=1.202
+ $X2=11.305 $Y2=1.202
r274 115 116 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=10.835 $Y=1.202
+ $X2=11.28 $Y2=1.202
r275 114 115 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=10.81 $Y=1.202
+ $X2=10.835 $Y2=1.202
r276 113 114 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=10.39 $Y=1.202
+ $X2=10.81 $Y2=1.202
r277 112 113 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=10.365 $Y=1.202
+ $X2=10.39 $Y2=1.202
r278 111 112 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=9.895 $Y=1.202
+ $X2=10.365 $Y2=1.202
r279 110 111 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=9.87 $Y=1.202
+ $X2=9.895 $Y2=1.202
r280 109 110 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=9.45 $Y=1.202
+ $X2=9.87 $Y2=1.202
r281 108 109 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=9.425 $Y=1.202
+ $X2=9.45 $Y2=1.202
r282 107 108 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=8.955 $Y=1.202
+ $X2=9.425 $Y2=1.202
r283 106 107 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=8.93 $Y=1.202
+ $X2=8.955 $Y2=1.202
r284 104 106 34.1471 $w=3.67e-07 $l=2.6e-07 $layer=POLY_cond $X=8.67 $Y=1.202
+ $X2=8.93 $Y2=1.202
r285 104 105 17.0918 $w=1.7e-07 $l=1.445e-06 $layer=licon1_POLY $count=8 $X=8.67
+ $Y=1.16 $X2=8.67 $Y2=1.16
r286 102 104 24.297 $w=3.67e-07 $l=1.85e-07 $layer=POLY_cond $X=8.485 $Y=1.202
+ $X2=8.67 $Y2=1.202
r287 101 102 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=8.46 $Y=1.202
+ $X2=8.485 $Y2=1.202
r288 100 101 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=8.015 $Y=1.202
+ $X2=8.46 $Y2=1.202
r289 99 100 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=7.99 $Y=1.202
+ $X2=8.015 $Y2=1.202
r290 97 130 121.22 $w=2.68e-07 $l=2.84e-06 $layer=LI1_cond $X=11.27 $Y=1.19
+ $X2=14.11 $Y2=1.19
r291 97 105 110.976 $w=2.68e-07 $l=2.6e-06 $layer=LI1_cond $X=11.27 $Y=1.19
+ $X2=8.67 $Y2=1.19
r292 94 136 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=15.09 $Y=0.995
+ $X2=15.09 $Y2=1.202
r293 94 96 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=15.09 $Y=0.995
+ $X2=15.09 $Y2=0.56
r294 91 135 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=15.065 $Y=1.41
+ $X2=15.065 $Y2=1.202
r295 91 93 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.065 $Y=1.41
+ $X2=15.065 $Y2=1.985
r296 88 134 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=14.595 $Y=1.41
+ $X2=14.595 $Y2=1.202
r297 88 90 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=14.595 $Y=1.41
+ $X2=14.595 $Y2=1.985
r298 85 133 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=14.57 $Y=0.995
+ $X2=14.57 $Y2=1.202
r299 85 87 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=14.57 $Y=0.995
+ $X2=14.57 $Y2=0.56
r300 82 132 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=14.15 $Y=0.995
+ $X2=14.15 $Y2=1.202
r301 82 84 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=14.15 $Y=0.995
+ $X2=14.15 $Y2=0.56
r302 79 131 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=14.125 $Y=1.41
+ $X2=14.125 $Y2=1.202
r303 79 81 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=14.125 $Y=1.41
+ $X2=14.125 $Y2=1.985
r304 76 127 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=13.655 $Y=1.41
+ $X2=13.655 $Y2=1.202
r305 76 78 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=13.655 $Y=1.41
+ $X2=13.655 $Y2=1.985
r306 73 126 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=13.63 $Y=0.995
+ $X2=13.63 $Y2=1.202
r307 73 75 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.63 $Y=0.995
+ $X2=13.63 $Y2=0.56
r308 70 125 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=13.21 $Y=0.995
+ $X2=13.21 $Y2=1.202
r309 70 72 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.21 $Y=0.995
+ $X2=13.21 $Y2=0.56
r310 67 124 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=13.185 $Y=1.41
+ $X2=13.185 $Y2=1.202
r311 67 69 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=13.185 $Y=1.41
+ $X2=13.185 $Y2=1.985
r312 64 123 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=12.715 $Y=1.41
+ $X2=12.715 $Y2=1.202
r313 64 66 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.715 $Y=1.41
+ $X2=12.715 $Y2=1.985
r314 61 122 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=12.69 $Y=0.995
+ $X2=12.69 $Y2=1.202
r315 61 63 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.69 $Y=0.995
+ $X2=12.69 $Y2=0.56
r316 58 121 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=12.27 $Y=0.995
+ $X2=12.27 $Y2=1.202
r317 58 60 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.27 $Y=0.995
+ $X2=12.27 $Y2=0.56
r318 55 120 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=12.245 $Y=1.41
+ $X2=12.245 $Y2=1.202
r319 55 57 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.245 $Y=1.41
+ $X2=12.245 $Y2=1.985
r320 52 119 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=11.775 $Y=1.41
+ $X2=11.775 $Y2=1.202
r321 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.775 $Y=1.41
+ $X2=11.775 $Y2=1.985
r322 49 118 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.75 $Y=0.995
+ $X2=11.75 $Y2=1.202
r323 49 51 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.75 $Y=0.995
+ $X2=11.75 $Y2=0.56
r324 46 117 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=11.305 $Y=1.41
+ $X2=11.305 $Y2=1.202
r325 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.305 $Y=1.41
+ $X2=11.305 $Y2=1.985
r326 43 116 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.28 $Y=0.995
+ $X2=11.28 $Y2=1.202
r327 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.28 $Y=0.995
+ $X2=11.28 $Y2=0.56
r328 40 115 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.835 $Y=1.41
+ $X2=10.835 $Y2=1.202
r329 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.835 $Y=1.41
+ $X2=10.835 $Y2=1.985
r330 37 114 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.81 $Y=0.995
+ $X2=10.81 $Y2=1.202
r331 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.81 $Y=0.995
+ $X2=10.81 $Y2=0.56
r332 34 113 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.39 $Y=0.995
+ $X2=10.39 $Y2=1.202
r333 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.39 $Y=0.995
+ $X2=10.39 $Y2=0.56
r334 31 112 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.365 $Y=1.41
+ $X2=10.365 $Y2=1.202
r335 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.365 $Y=1.41
+ $X2=10.365 $Y2=1.985
r336 28 111 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.895 $Y=1.41
+ $X2=9.895 $Y2=1.202
r337 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.895 $Y=1.41
+ $X2=9.895 $Y2=1.985
r338 25 110 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.87 $Y=0.995
+ $X2=9.87 $Y2=1.202
r339 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.87 $Y=0.995
+ $X2=9.87 $Y2=0.56
r340 22 109 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.45 $Y=0.995
+ $X2=9.45 $Y2=1.202
r341 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.45 $Y=0.995
+ $X2=9.45 $Y2=0.56
r342 19 108 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.425 $Y=1.41
+ $X2=9.425 $Y2=1.202
r343 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.425 $Y=1.41
+ $X2=9.425 $Y2=1.985
r344 16 107 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.955 $Y=1.41
+ $X2=8.955 $Y2=1.202
r345 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.955 $Y=1.41
+ $X2=8.955 $Y2=1.985
r346 13 106 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.93 $Y=0.995
+ $X2=8.93 $Y2=1.202
r347 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.93 $Y=0.995
+ $X2=8.93 $Y2=0.56
r348 10 102 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.485 $Y=1.41
+ $X2=8.485 $Y2=1.202
r349 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.485 $Y=1.41
+ $X2=8.485 $Y2=1.985
r350 7 101 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.46 $Y=0.995
+ $X2=8.46 $Y2=1.202
r351 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.46 $Y=0.995
+ $X2=8.46 $Y2=0.56
r352 4 100 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.015 $Y=1.41
+ $X2=8.015 $Y2=1.202
r353 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.015 $Y=1.41
+ $X2=8.015 $Y2=1.985
r354 1 99 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.99 $Y=0.995
+ $X2=7.99 $Y2=1.202
r355 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.99 $Y=0.995
+ $X2=7.99 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
+ 16 17 52 54 60 62 66 68 72 74 78 80 84 88 92 96 100 104 108 112 116 120 124
+ 126 128 133 134 136 137 139 140 142 143 145 146 148 149 151 152 154 155 157
+ 158 160 161 162 164 200 208 211 214 217 220 224
r228 223 224 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.41 $Y=2.72
+ $X2=15.41 $Y2=2.72
r229 220 221 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r230 218 221 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r231 217 218 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r232 215 218 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r233 214 215 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r234 212 215 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r235 211 212 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r236 209 212 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r237 208 209 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r238 203 224 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.95 $Y=2.72
+ $X2=15.41 $Y2=2.72
r239 202 203 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.95 $Y=2.72
+ $X2=14.95 $Y2=2.72
r240 200 223 4.07187 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=15.165 $Y=2.72
+ $X2=15.402 $Y2=2.72
r241 200 202 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=15.165 $Y=2.72
+ $X2=14.95 $Y2=2.72
r242 199 203 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=14.03 $Y=2.72
+ $X2=14.95 $Y2=2.72
r243 198 199 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.03 $Y=2.72
+ $X2=14.03 $Y2=2.72
r244 196 199 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.11 $Y=2.72
+ $X2=14.03 $Y2=2.72
r245 195 196 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r246 193 196 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.19 $Y=2.72
+ $X2=13.11 $Y2=2.72
r247 192 193 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r248 190 193 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=12.19 $Y2=2.72
r249 189 190 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r250 187 190 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=11.27 $Y2=2.72
r251 186 187 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r252 184 187 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=10.35 $Y2=2.72
r253 183 184 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r254 181 184 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r255 180 181 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r256 178 181 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r257 177 178 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r258 175 178 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r259 174 175 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r260 172 175 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r261 172 221 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=4.83 $Y2=2.72
r262 171 172 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r263 169 220 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.095 $Y=2.72
+ $X2=4.96 $Y2=2.72
r264 169 171 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.095 $Y=2.72
+ $X2=5.75 $Y2=2.72
r265 168 209 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r266 167 168 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r267 165 205 4.1687 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r268 165 167 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.69 $Y2=2.72
r269 164 208 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=1.2 $Y2=2.72
r270 164 167 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=0.69 $Y2=2.72
r271 162 168 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r272 162 205 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r273 160 198 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=14.225 $Y=2.72
+ $X2=14.03 $Y2=2.72
r274 160 161 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.225 $Y=2.72
+ $X2=14.36 $Y2=2.72
r275 159 202 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=14.495 $Y=2.72
+ $X2=14.95 $Y2=2.72
r276 159 161 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.495 $Y=2.72
+ $X2=14.36 $Y2=2.72
r277 157 195 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=13.285 $Y=2.72
+ $X2=13.11 $Y2=2.72
r278 157 158 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.285 $Y=2.72
+ $X2=13.42 $Y2=2.72
r279 156 198 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=13.555 $Y=2.72
+ $X2=14.03 $Y2=2.72
r280 156 158 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.555 $Y=2.72
+ $X2=13.42 $Y2=2.72
r281 154 192 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=12.345 $Y=2.72
+ $X2=12.19 $Y2=2.72
r282 154 155 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.345 $Y=2.72
+ $X2=12.48 $Y2=2.72
r283 153 195 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=12.615 $Y=2.72
+ $X2=13.11 $Y2=2.72
r284 153 155 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.615 $Y=2.72
+ $X2=12.48 $Y2=2.72
r285 151 189 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=11.405 $Y=2.72
+ $X2=11.27 $Y2=2.72
r286 151 152 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.405 $Y=2.72
+ $X2=11.54 $Y2=2.72
r287 150 192 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=11.675 $Y=2.72
+ $X2=12.19 $Y2=2.72
r288 150 152 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.675 $Y=2.72
+ $X2=11.54 $Y2=2.72
r289 148 186 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=10.465 $Y=2.72
+ $X2=10.35 $Y2=2.72
r290 148 149 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.465 $Y=2.72
+ $X2=10.6 $Y2=2.72
r291 147 189 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=10.735 $Y=2.72
+ $X2=11.27 $Y2=2.72
r292 147 149 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.735 $Y=2.72
+ $X2=10.6 $Y2=2.72
r293 145 183 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=9.525 $Y=2.72
+ $X2=9.43 $Y2=2.72
r294 145 146 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=9.525 $Y=2.72
+ $X2=9.66 $Y2=2.72
r295 144 186 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=9.795 $Y=2.72
+ $X2=10.35 $Y2=2.72
r296 144 146 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=9.795 $Y=2.72
+ $X2=9.66 $Y2=2.72
r297 142 180 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=8.585 $Y=2.72
+ $X2=8.51 $Y2=2.72
r298 142 143 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.585 $Y=2.72
+ $X2=8.72 $Y2=2.72
r299 141 183 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=8.855 $Y=2.72
+ $X2=9.43 $Y2=2.72
r300 141 143 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.855 $Y=2.72
+ $X2=8.72 $Y2=2.72
r301 139 177 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=7.645 $Y=2.72
+ $X2=7.59 $Y2=2.72
r302 139 140 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.645 $Y=2.72
+ $X2=7.78 $Y2=2.72
r303 138 180 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=7.915 $Y=2.72
+ $X2=8.51 $Y2=2.72
r304 138 140 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.915 $Y=2.72
+ $X2=7.78 $Y2=2.72
r305 136 174 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.705 $Y=2.72
+ $X2=6.67 $Y2=2.72
r306 136 137 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.705 $Y=2.72
+ $X2=6.84 $Y2=2.72
r307 135 177 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=6.975 $Y=2.72
+ $X2=7.59 $Y2=2.72
r308 135 137 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.975 $Y=2.72
+ $X2=6.84 $Y2=2.72
r309 133 171 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=5.765 $Y=2.72
+ $X2=5.75 $Y2=2.72
r310 133 134 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.765 $Y=2.72
+ $X2=5.9 $Y2=2.72
r311 132 174 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.035 $Y=2.72
+ $X2=6.67 $Y2=2.72
r312 132 134 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.035 $Y=2.72
+ $X2=5.9 $Y2=2.72
r313 128 131 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=15.3 $Y=1.66
+ $X2=15.3 $Y2=2.34
r314 126 223 3.21282 $w=2.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=15.3 $Y=2.635
+ $X2=15.402 $Y2=2.72
r315 126 131 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=15.3 $Y=2.635
+ $X2=15.3 $Y2=2.34
r316 122 161 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.36 $Y=2.635
+ $X2=14.36 $Y2=2.72
r317 122 124 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=14.36 $Y=2.635
+ $X2=14.36 $Y2=2
r318 118 158 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.42 $Y=2.635
+ $X2=13.42 $Y2=2.72
r319 118 120 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=13.42 $Y=2.635
+ $X2=13.42 $Y2=2
r320 114 155 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.48 $Y=2.635
+ $X2=12.48 $Y2=2.72
r321 114 116 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=12.48 $Y=2.635
+ $X2=12.48 $Y2=2
r322 110 152 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.54 $Y=2.635
+ $X2=11.54 $Y2=2.72
r323 110 112 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=11.54 $Y=2.635
+ $X2=11.54 $Y2=2
r324 106 149 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.6 $Y=2.635
+ $X2=10.6 $Y2=2.72
r325 106 108 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=10.6 $Y=2.635
+ $X2=10.6 $Y2=2
r326 102 146 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.66 $Y=2.635
+ $X2=9.66 $Y2=2.72
r327 102 104 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=9.66 $Y=2.635
+ $X2=9.66 $Y2=2
r328 98 143 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.72 $Y=2.635
+ $X2=8.72 $Y2=2.72
r329 98 100 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.72 $Y=2.635
+ $X2=8.72 $Y2=2
r330 94 140 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.78 $Y=2.635
+ $X2=7.78 $Y2=2.72
r331 94 96 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.78 $Y=2.635
+ $X2=7.78 $Y2=2
r332 90 137 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=2.635
+ $X2=6.84 $Y2=2.72
r333 90 92 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.84 $Y=2.635
+ $X2=6.84 $Y2=2
r334 86 134 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=2.635
+ $X2=5.9 $Y2=2.72
r335 86 88 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.9 $Y=2.635
+ $X2=5.9 $Y2=2
r336 82 220 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=2.72
r337 82 84 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=2
r338 81 217 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.155 $Y=2.72
+ $X2=4.02 $Y2=2.72
r339 80 220 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.825 $Y=2.72
+ $X2=4.96 $Y2=2.72
r340 80 81 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.825 $Y=2.72
+ $X2=4.155 $Y2=2.72
r341 76 217 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=2.72
r342 76 78 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=2
r343 75 214 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=3.08 $Y2=2.72
r344 74 217 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=4.02 $Y2=2.72
r345 74 75 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=3.215 $Y2=2.72
r346 70 214 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2.72
r347 70 72 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2
r348 69 211 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.14 $Y2=2.72
r349 68 214 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=3.08 $Y2=2.72
r350 68 69 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=2.275 $Y2=2.72
r351 64 211 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.72
r352 64 66 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2
r353 63 208 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.2 $Y2=2.72
r354 62 211 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=2.14 $Y2=2.72
r355 62 63 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=1.335 $Y2=2.72
r356 58 208 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.72
r357 58 60 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r358 54 57 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r359 52 205 3.116 $w=2.7e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.197 $Y2=2.72
r360 52 57 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r361 17 131 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=15.155
+ $Y=1.485 $X2=15.3 $Y2=2.34
r362 17 128 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=15.155
+ $Y=1.485 $X2=15.3 $Y2=1.66
r363 16 124 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=14.215
+ $Y=1.485 $X2=14.36 $Y2=2
r364 15 120 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=13.275
+ $Y=1.485 $X2=13.42 $Y2=2
r365 14 116 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=12.335
+ $Y=1.485 $X2=12.48 $Y2=2
r366 13 112 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=11.395
+ $Y=1.485 $X2=11.54 $Y2=2
r367 12 108 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=10.455
+ $Y=1.485 $X2=10.6 $Y2=2
r368 11 104 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=9.515
+ $Y=1.485 $X2=9.66 $Y2=2
r369 10 100 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=8.575
+ $Y=1.485 $X2=8.72 $Y2=2
r370 9 96 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=7.635
+ $Y=1.485 $X2=7.78 $Y2=2
r371 8 92 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.695
+ $Y=1.485 $X2=6.84 $Y2=2
r372 7 88 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.755
+ $Y=1.485 $X2=5.9 $Y2=2
r373 6 84 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=2
r374 5 78 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=2
r375 4 72 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2
r376 3 66 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r377 2 60 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r378 1 57 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r379 1 54 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 17 18 19 20 21 22 23 24 73 75 77 81 83 87 89 93 95 99 101 105 107 111 113 117
+ 119 121 125 127 141 145 147 151 153 157 159 163 165 169 171 175 177 181 183
+ 186 190 192 194 196 198 200 202 205 209 211 213 215 217 219 221 224 225 226
+ 232 234
r329 229 234 1.96759 $w=4.08e-07 $l=7e-08 $layer=LI1_cond $X=8.13 $Y=1.26
+ $X2=8.13 $Y2=1.19
r330 226 234 0.224867 $w=4.08e-07 $l=8e-09 $layer=LI1_cond $X=8.13 $Y=1.182
+ $X2=8.13 $Y2=1.19
r331 226 232 4.42096 $w=4.08e-07 $l=1.27e-07 $layer=LI1_cond $X=8.13 $Y=1.182
+ $X2=8.13 $Y2=1.055
r332 226 229 0.196759 $w=4.08e-07 $l=7e-09 $layer=LI1_cond $X=8.13 $Y=1.267
+ $X2=8.13 $Y2=1.26
r333 224 225 7.97845 $w=3.88e-07 $l=2.7e-07 $layer=LI1_cond $X=14.92 $Y=1.055
+ $X2=14.92 $Y2=1.325
r334 203 226 6.40871 $w=4.08e-07 $l=2.28e-07 $layer=LI1_cond $X=8.13 $Y=1.495
+ $X2=8.13 $Y2=1.267
r335 203 205 1.06026 $w=4.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=8.13 $Y=1.495
+ $X2=8.17 $Y2=1.58
r336 186 221 3.14896 $w=3e-07 $l=9.88686e-08 $layer=LI1_cond $X=14.86 $Y=1.495
+ $X2=14.83 $Y2=1.58
r337 186 225 7.25612 $w=2.68e-07 $l=1.7e-07 $layer=LI1_cond $X=14.86 $Y=1.495
+ $X2=14.86 $Y2=1.325
r338 183 223 3.28347 $w=2.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.86 $Y=0.885
+ $X2=14.86 $Y2=0.76
r339 183 224 7.25612 $w=2.68e-07 $l=1.7e-07 $layer=LI1_cond $X=14.86 $Y=0.885
+ $X2=14.86 $Y2=1.055
r340 179 221 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.83 $Y=1.665
+ $X2=14.83 $Y2=1.58
r341 179 181 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=14.83 $Y=1.665
+ $X2=14.83 $Y2=2.34
r342 178 219 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.055 $Y=1.58
+ $X2=13.89 $Y2=1.58
r343 177 221 3.44808 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.665 $Y=1.58
+ $X2=14.83 $Y2=1.58
r344 177 178 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=14.665 $Y=1.58
+ $X2=14.055 $Y2=1.58
r345 173 219 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.89 $Y=1.665
+ $X2=13.89 $Y2=1.58
r346 173 175 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=13.89 $Y=1.665
+ $X2=13.89 $Y2=2.34
r347 172 217 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.115 $Y=1.58
+ $X2=12.95 $Y2=1.58
r348 171 219 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.725 $Y=1.58
+ $X2=13.89 $Y2=1.58
r349 171 172 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=13.725 $Y=1.58
+ $X2=13.115 $Y2=1.58
r350 167 217 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.95 $Y=1.665
+ $X2=12.95 $Y2=1.58
r351 167 169 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=12.95 $Y=1.665
+ $X2=12.95 $Y2=2.34
r352 166 215 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.175 $Y=1.58
+ $X2=12.01 $Y2=1.58
r353 165 217 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.785 $Y=1.58
+ $X2=12.95 $Y2=1.58
r354 165 166 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=12.785 $Y=1.58
+ $X2=12.175 $Y2=1.58
r355 161 215 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.01 $Y=1.665
+ $X2=12.01 $Y2=1.58
r356 161 163 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=12.01 $Y=1.665
+ $X2=12.01 $Y2=2.34
r357 160 213 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.235 $Y=1.58
+ $X2=11.07 $Y2=1.58
r358 159 215 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.845 $Y=1.58
+ $X2=12.01 $Y2=1.58
r359 159 160 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=11.845 $Y=1.58
+ $X2=11.235 $Y2=1.58
r360 155 213 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.07 $Y=1.665
+ $X2=11.07 $Y2=1.58
r361 155 157 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=11.07 $Y=1.665
+ $X2=11.07 $Y2=2.34
r362 154 211 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.295 $Y=1.58
+ $X2=10.13 $Y2=1.58
r363 153 213 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.905 $Y=1.58
+ $X2=11.07 $Y2=1.58
r364 153 154 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=10.905 $Y=1.58
+ $X2=10.295 $Y2=1.58
r365 149 211 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.13 $Y=1.665
+ $X2=10.13 $Y2=1.58
r366 149 151 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=10.13 $Y=1.665
+ $X2=10.13 $Y2=2.34
r367 148 209 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.355 $Y=1.58
+ $X2=9.19 $Y2=1.58
r368 147 211 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.965 $Y=1.58
+ $X2=10.13 $Y2=1.58
r369 147 148 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=9.965 $Y=1.58
+ $X2=9.355 $Y2=1.58
r370 143 209 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.19 $Y=1.665
+ $X2=9.19 $Y2=1.58
r371 143 145 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=9.19 $Y=1.665
+ $X2=9.19 $Y2=2.34
r372 142 205 5.68638 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=8.415 $Y=1.58
+ $X2=8.17 $Y2=1.58
r373 141 209 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.025 $Y=1.58
+ $X2=9.19 $Y2=1.58
r374 141 142 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=9.025 $Y=1.58
+ $X2=8.415 $Y2=1.58
r375 138 140 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=12.95 $Y=0.76
+ $X2=13.89 $Y2=0.76
r376 136 138 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=12.01 $Y=0.76
+ $X2=12.95 $Y2=0.76
r377 134 136 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=11.07 $Y=0.76
+ $X2=12.01 $Y2=0.76
r378 132 134 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=10.13 $Y=0.76
+ $X2=11.07 $Y2=0.76
r379 130 132 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=9.19 $Y=0.76
+ $X2=10.13 $Y2=0.76
r380 128 207 3.75819 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=8.335 $Y=0.76
+ $X2=8.185 $Y2=0.76
r381 128 130 39.4136 $w=2.48e-07 $l=8.55e-07 $layer=LI1_cond $X=8.335 $Y=0.76
+ $X2=9.19 $Y2=0.76
r382 127 223 3.54615 $w=2.5e-07 $l=1.35e-07 $layer=LI1_cond $X=14.725 $Y=0.76
+ $X2=14.86 $Y2=0.76
r383 127 140 38.4916 $w=2.48e-07 $l=8.35e-07 $layer=LI1_cond $X=14.725 $Y=0.76
+ $X2=13.89 $Y2=0.76
r384 123 205 1.06026 $w=3.3e-07 $l=1.18427e-07 $layer=LI1_cond $X=8.25 $Y=1.665
+ $X2=8.17 $Y2=1.58
r385 123 125 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=8.25 $Y=1.665
+ $X2=8.25 $Y2=2.34
r386 121 207 3.13183 $w=3e-07 $l=1.25e-07 $layer=LI1_cond $X=8.185 $Y=0.885
+ $X2=8.185 $Y2=0.76
r387 121 232 6.53051 $w=2.98e-07 $l=1.7e-07 $layer=LI1_cond $X=8.185 $Y=0.885
+ $X2=8.185 $Y2=1.055
r388 120 202 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.475 $Y=1.58
+ $X2=7.31 $Y2=1.58
r389 119 205 5.68638 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=7.925 $Y=1.58
+ $X2=8.17 $Y2=1.58
r390 119 120 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=7.925 $Y=1.58
+ $X2=7.475 $Y2=1.58
r391 115 202 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.31 $Y=1.665
+ $X2=7.31 $Y2=1.58
r392 115 117 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=7.31 $Y=1.665
+ $X2=7.31 $Y2=2.34
r393 114 200 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.535 $Y=1.58
+ $X2=6.37 $Y2=1.58
r394 113 202 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.145 $Y=1.58
+ $X2=7.31 $Y2=1.58
r395 113 114 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.145 $Y=1.58
+ $X2=6.535 $Y2=1.58
r396 109 200 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.37 $Y=1.665
+ $X2=6.37 $Y2=1.58
r397 109 111 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.37 $Y=1.665
+ $X2=6.37 $Y2=2.34
r398 108 198 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.595 $Y=1.58
+ $X2=5.43 $Y2=1.58
r399 107 200 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.205 $Y=1.58
+ $X2=6.37 $Y2=1.58
r400 107 108 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.205 $Y=1.58
+ $X2=5.595 $Y2=1.58
r401 103 198 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.43 $Y=1.665
+ $X2=5.43 $Y2=1.58
r402 103 105 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.43 $Y=1.665
+ $X2=5.43 $Y2=2.34
r403 102 196 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.655 $Y=1.58
+ $X2=4.49 $Y2=1.58
r404 101 198 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.265 $Y=1.58
+ $X2=5.43 $Y2=1.58
r405 101 102 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.265 $Y=1.58
+ $X2=4.655 $Y2=1.58
r406 97 196 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=1.665
+ $X2=4.49 $Y2=1.58
r407 97 99 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.49 $Y=1.665
+ $X2=4.49 $Y2=2.34
r408 96 194 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.715 $Y=1.58
+ $X2=3.55 $Y2=1.58
r409 95 196 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.325 $Y=1.58
+ $X2=4.49 $Y2=1.58
r410 95 96 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.325 $Y=1.58
+ $X2=3.715 $Y2=1.58
r411 91 194 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=1.665
+ $X2=3.55 $Y2=1.58
r412 91 93 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.55 $Y=1.665
+ $X2=3.55 $Y2=2.34
r413 90 192 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=1.58
+ $X2=2.61 $Y2=1.58
r414 89 194 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=1.58
+ $X2=3.55 $Y2=1.58
r415 89 90 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.385 $Y=1.58
+ $X2=2.775 $Y2=1.58
r416 85 192 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=1.58
r417 85 87 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=2.34
r418 84 190 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=1.58
+ $X2=1.67 $Y2=1.58
r419 83 192 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=1.58
+ $X2=2.61 $Y2=1.58
r420 83 84 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.445 $Y=1.58
+ $X2=1.835 $Y2=1.58
r421 79 190 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=1.58
r422 79 81 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=2.34
r423 78 188 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.73 $Y2=1.58
r424 77 190 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=1.67 $Y2=1.58
r425 77 78 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=0.895 $Y2=1.58
r426 73 188 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=1.58
r427 73 75 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=2.34
r428 24 221 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=14.685
+ $Y=1.485 $X2=14.83 $Y2=1.66
r429 24 181 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=14.685
+ $Y=1.485 $X2=14.83 $Y2=2.34
r430 23 219 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=13.745
+ $Y=1.485 $X2=13.89 $Y2=1.66
r431 23 175 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=13.745
+ $Y=1.485 $X2=13.89 $Y2=2.34
r432 22 217 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=12.805
+ $Y=1.485 $X2=12.95 $Y2=1.66
r433 22 169 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=12.805
+ $Y=1.485 $X2=12.95 $Y2=2.34
r434 21 215 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=11.865
+ $Y=1.485 $X2=12.01 $Y2=1.66
r435 21 163 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=11.865
+ $Y=1.485 $X2=12.01 $Y2=2.34
r436 20 213 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=10.925
+ $Y=1.485 $X2=11.07 $Y2=1.66
r437 20 157 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.925
+ $Y=1.485 $X2=11.07 $Y2=2.34
r438 19 211 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=9.985
+ $Y=1.485 $X2=10.13 $Y2=1.66
r439 19 151 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=9.985
+ $Y=1.485 $X2=10.13 $Y2=2.34
r440 18 209 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=9.045
+ $Y=1.485 $X2=9.19 $Y2=1.66
r441 18 145 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=9.045
+ $Y=1.485 $X2=9.19 $Y2=2.34
r442 17 205 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=8.105
+ $Y=1.485 $X2=8.25 $Y2=1.66
r443 17 125 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=8.105
+ $Y=1.485 $X2=8.25 $Y2=2.34
r444 16 202 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=7.165
+ $Y=1.485 $X2=7.31 $Y2=1.66
r445 16 117 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.165
+ $Y=1.485 $X2=7.31 $Y2=2.34
r446 15 200 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=6.225
+ $Y=1.485 $X2=6.37 $Y2=1.66
r447 15 111 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.225
+ $Y=1.485 $X2=6.37 $Y2=2.34
r448 14 198 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=1.66
r449 14 105 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=2.34
r450 13 196 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=1.66
r451 13 99 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=2.34
r452 12 194 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.66
r453 12 93 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2.34
r454 11 192 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.66
r455 11 87 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.34
r456 10 190 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r457 10 81 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
r458 9 188 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r459 9 75 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r460 8 223 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=14.645
+ $Y=0.235 $X2=14.83 $Y2=0.72
r461 7 140 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=13.705
+ $Y=0.235 $X2=13.89 $Y2=0.72
r462 6 138 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=12.765
+ $Y=0.235 $X2=12.95 $Y2=0.72
r463 5 136 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=11.825
+ $Y=0.235 $X2=12.01 $Y2=0.72
r464 4 134 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=10.885
+ $Y=0.235 $X2=11.07 $Y2=0.72
r465 3 132 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=9.945
+ $Y=0.235 $X2=10.13 $Y2=0.72
r466 2 130 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=9.005
+ $Y=0.235 $X2=9.19 $Y2=0.72
r467 1 207 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=8.065
+ $Y=0.235 $X2=8.25 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_16%A_27_47# 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 54 56 57 60 62 66 68 72 74 78 80 84 86 90 92 96 98 100 101 102 118
+ 120 122 123 124 125 126 127 128
r227 118 134 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=15.34 $Y=0.465
+ $X2=15.34 $Y2=0.36
r228 118 120 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=15.34 $Y=0.465
+ $X2=15.34 $Y2=0.72
r229 115 117 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=13.42 $Y=0.36
+ $X2=14.36 $Y2=0.36
r230 113 115 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=12.48 $Y=0.36
+ $X2=13.42 $Y2=0.36
r231 111 113 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=11.54 $Y=0.36
+ $X2=12.48 $Y2=0.36
r232 109 111 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=10.6 $Y=0.36
+ $X2=11.54 $Y2=0.36
r233 107 109 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=9.66 $Y=0.36
+ $X2=10.6 $Y2=0.36
r234 105 107 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=8.72 $Y=0.36
+ $X2=9.66 $Y2=0.36
r235 103 130 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=7.865 $Y=0.36
+ $X2=7.74 $Y2=0.36
r236 103 105 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=7.865 $Y=0.36
+ $X2=8.72 $Y2=0.36
r237 102 134 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=15.215 $Y=0.36
+ $X2=15.34 $Y2=0.36
r238 102 117 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=15.215 $Y=0.36
+ $X2=14.36 $Y2=0.36
r239 101 132 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.74 $Y=0.715
+ $X2=7.74 $Y2=0.8
r240 100 130 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=7.74 $Y=0.465
+ $X2=7.74 $Y2=0.36
r241 100 101 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=7.74 $Y=0.465
+ $X2=7.74 $Y2=0.715
r242 99 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.005 $Y=0.8
+ $X2=6.84 $Y2=0.8
r243 98 132 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.615 $Y=0.8
+ $X2=7.74 $Y2=0.8
r244 98 99 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.615 $Y=0.8
+ $X2=7.005 $Y2=0.8
r245 94 128 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=0.715
+ $X2=6.84 $Y2=0.8
r246 94 96 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.84 $Y=0.715
+ $X2=6.84 $Y2=0.38
r247 93 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.065 $Y=0.8
+ $X2=5.9 $Y2=0.8
r248 92 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=0.8
+ $X2=6.84 $Y2=0.8
r249 92 93 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.675 $Y=0.8
+ $X2=6.065 $Y2=0.8
r250 88 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=0.715
+ $X2=5.9 $Y2=0.8
r251 88 90 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.9 $Y=0.715
+ $X2=5.9 $Y2=0.38
r252 87 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=0.8
+ $X2=4.96 $Y2=0.8
r253 86 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.735 $Y=0.8
+ $X2=5.9 $Y2=0.8
r254 86 87 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.735 $Y=0.8
+ $X2=5.125 $Y2=0.8
r255 82 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=0.715
+ $X2=4.96 $Y2=0.8
r256 82 84 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.96 $Y=0.715
+ $X2=4.96 $Y2=0.38
r257 81 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=0.8
+ $X2=4.02 $Y2=0.8
r258 80 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=0.8
+ $X2=4.96 $Y2=0.8
r259 80 81 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.795 $Y=0.8
+ $X2=4.185 $Y2=0.8
r260 76 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.715
+ $X2=4.02 $Y2=0.8
r261 76 78 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.02 $Y=0.715
+ $X2=4.02 $Y2=0.38
r262 75 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=0.8
+ $X2=3.08 $Y2=0.8
r263 74 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=0.8
+ $X2=4.02 $Y2=0.8
r264 74 75 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.855 $Y=0.8
+ $X2=3.245 $Y2=0.8
r265 70 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.715
+ $X2=3.08 $Y2=0.8
r266 70 72 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.08 $Y=0.715
+ $X2=3.08 $Y2=0.38
r267 69 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=0.8
+ $X2=2.14 $Y2=0.8
r268 68 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=0.8
+ $X2=3.08 $Y2=0.8
r269 68 69 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.915 $Y=0.8
+ $X2=2.305 $Y2=0.8
r270 64 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.715
+ $X2=2.14 $Y2=0.8
r271 64 66 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.14 $Y=0.715
+ $X2=2.14 $Y2=0.38
r272 63 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=0.8
+ $X2=1.2 $Y2=0.8
r273 62 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0.8
+ $X2=2.14 $Y2=0.8
r274 62 63 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.975 $Y=0.8
+ $X2=1.365 $Y2=0.8
r275 58 122 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.715
+ $X2=1.2 $Y2=0.8
r276 58 60 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.2 $Y=0.715
+ $X2=1.2 $Y2=0.38
r277 56 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0.8
+ $X2=1.2 $Y2=0.8
r278 56 57 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.035 $Y=0.8
+ $X2=0.425 $Y2=0.8
r279 52 57 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=0.715
+ $X2=0.425 $Y2=0.8
r280 52 54 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.26 $Y=0.715
+ $X2=0.26 $Y2=0.38
r281 17 134 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=15.165
+ $Y=0.235 $X2=15.3 $Y2=0.38
r282 17 120 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=15.165
+ $Y=0.235 $X2=15.3 $Y2=0.72
r283 16 117 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=14.225
+ $Y=0.235 $X2=14.36 $Y2=0.38
r284 15 115 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=13.285
+ $Y=0.235 $X2=13.42 $Y2=0.38
r285 14 113 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=12.345
+ $Y=0.235 $X2=12.48 $Y2=0.38
r286 13 111 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=11.355
+ $Y=0.235 $X2=11.54 $Y2=0.38
r287 12 109 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=10.465
+ $Y=0.235 $X2=10.6 $Y2=0.38
r288 11 107 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=9.525
+ $Y=0.235 $X2=9.66 $Y2=0.38
r289 10 105 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=8.535
+ $Y=0.235 $X2=8.72 $Y2=0.38
r290 9 132 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=7.645
+ $Y=0.235 $X2=7.78 $Y2=0.72
r291 9 130 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.645
+ $Y=0.235 $X2=7.78 $Y2=0.38
r292 8 96 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=6.705
+ $Y=0.235 $X2=6.84 $Y2=0.38
r293 7 90 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.765
+ $Y=0.235 $X2=5.9 $Y2=0.38
r294 6 84 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=4.825
+ $Y=0.235 $X2=4.96 $Y2=0.38
r295 5 78 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.885
+ $Y=0.235 $X2=4.02 $Y2=0.38
r296 4 72 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.945
+ $Y=0.235 $X2=3.08 $Y2=0.38
r297 3 66 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.38
r298 2 60 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.38
r299 1 54 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_16%VGND 1 2 3 4 5 6 7 8 27 29 33 35 39 41 45
+ 47 51 55 59 63 66 67 69 70 72 73 74 76 95 96 99 102 105 108 111
r193 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r194 109 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.37 $Y2=0
r195 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r196 106 109 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.45 $Y2=0
r197 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r198 103 106 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.53 $Y2=0
r199 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r200 100 103 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.61 $Y2=0
r201 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r202 95 96 1.03333 $w=1.7e-07 $l=1.53e-06 $layer=mcon $count=9 $X=15.41 $Y=0
+ $X2=15.41 $Y2=0
r203 93 96 2.22512 $w=4.8e-07 $l=7.82e-06 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=15.41 $Y2=0
r204 92 95 510.182 $w=1.68e-07 $l=7.82e-06 $layer=LI1_cond $X=7.59 $Y=0
+ $X2=15.41 $Y2=0
r205 92 93 1.03333 $w=1.7e-07 $l=1.53e-06 $layer=mcon $count=9 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r206 90 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=7.59
+ $Y2=0
r207 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r208 87 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r209 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r210 84 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r211 84 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=4.37 $Y2=0
r212 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r213 81 111 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.625 $Y=0
+ $X2=4.49 $Y2=0
r214 81 83 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.625 $Y=0 $X2=5.29
+ $Y2=0
r215 76 99 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.73
+ $Y2=0
r216 76 78 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0
+ $X2=0.23 $Y2=0
r217 74 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r218 74 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r219 72 89 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=7.175 $Y=0 $X2=7.13
+ $Y2=0
r220 72 73 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.175 $Y=0 $X2=7.31
+ $Y2=0
r221 71 92 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.445 $Y=0
+ $X2=7.59 $Y2=0
r222 71 73 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.445 $Y=0 $X2=7.31
+ $Y2=0
r223 69 86 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=6.235 $Y=0 $X2=6.21
+ $Y2=0
r224 69 70 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.235 $Y=0 $X2=6.37
+ $Y2=0
r225 68 89 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=6.505 $Y=0
+ $X2=7.13 $Y2=0
r226 68 70 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.505 $Y=0 $X2=6.37
+ $Y2=0
r227 66 83 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.295 $Y=0 $X2=5.29
+ $Y2=0
r228 66 67 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.295 $Y=0 $X2=5.43
+ $Y2=0
r229 65 86 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=5.565 $Y=0
+ $X2=6.21 $Y2=0
r230 65 67 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.565 $Y=0 $X2=5.43
+ $Y2=0
r231 61 73 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.31 $Y=0.085
+ $X2=7.31 $Y2=0
r232 61 63 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.31 $Y=0.085
+ $X2=7.31 $Y2=0.38
r233 57 70 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.37 $Y=0.085
+ $X2=6.37 $Y2=0
r234 57 59 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.37 $Y=0.085
+ $X2=6.37 $Y2=0.38
r235 53 67 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.43 $Y=0.085
+ $X2=5.43 $Y2=0
r236 53 55 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.43 $Y=0.085
+ $X2=5.43 $Y2=0.38
r237 49 111 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=0.085
+ $X2=4.49 $Y2=0
r238 49 51 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.49 $Y=0.085
+ $X2=4.49 $Y2=0.38
r239 48 108 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.685 $Y=0
+ $X2=3.55 $Y2=0
r240 47 111 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.355 $Y=0
+ $X2=4.49 $Y2=0
r241 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.355 $Y=0
+ $X2=3.685 $Y2=0
r242 43 108 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0
r243 43 45 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0.38
r244 42 105 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.745 $Y=0
+ $X2=2.61 $Y2=0
r245 41 108 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.415 $Y=0
+ $X2=3.55 $Y2=0
r246 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.415 $Y=0
+ $X2=2.745 $Y2=0
r247 37 105 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0
r248 37 39 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0.38
r249 36 102 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.805 $Y=0
+ $X2=1.67 $Y2=0
r250 35 105 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.475 $Y=0
+ $X2=2.61 $Y2=0
r251 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.475 $Y=0
+ $X2=1.805 $Y2=0
r252 31 102 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0
r253 31 33 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0.38
r254 30 99 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=0.73
+ $Y2=0
r255 29 102 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.535 $Y=0
+ $X2=1.67 $Y2=0
r256 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.535 $Y=0
+ $X2=0.865 $Y2=0
r257 25 99 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r258 25 27 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.38
r259 8 63 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=7.125
+ $Y=0.235 $X2=7.31 $Y2=0.38
r260 7 59 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=6.185
+ $Y=0.235 $X2=6.37 $Y2=0.38
r261 6 55 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=5.245
+ $Y=0.235 $X2=5.43 $Y2=0.38
r262 5 51 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.235 $X2=4.49 $Y2=0.38
r263 4 45 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.38
r264 3 39 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.38
r265 2 33 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.38
r266 1 27 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

