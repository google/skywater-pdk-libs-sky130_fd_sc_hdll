* NGSPICE file created from sky130_fd_sc_hdll__nor3b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__nor3b_1 A B C_N VGND VNB VPB VPWR Y
M1000 a_91_199# C_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=4.62e+11p ps=4.11e+06u
M1001 a_263_297# B a_169_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u
M1002 a_169_297# a_91_199# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.3e+11p ps=2.66e+06u
M1003 a_91_199# C_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=3.057e+11p ps=2.71e+06u
M1004 Y B VGND VNB nshort w=650000u l=150000u
+  ad=4.29e+11p pd=3.92e+06u as=0p ps=0u
M1005 VGND a_91_199# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_263_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

