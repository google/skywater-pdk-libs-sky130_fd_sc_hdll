* File: sky130_fd_sc_hdll__o21ba_2.spice
* Created: Wed Sep  2 08:43:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o21ba_2.pex.spice"
.subckt sky130_fd_sc_hdll__o21ba_2  VNB VPB B1_N A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_B1_N_M1011_g N_A_27_93#_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0869439 AS=0.1092 PD=0.812523 PS=1.36 NRD=12.852 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1011_d N_A_186_21#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.134556 AS=0.128375 PD=1.25748 PS=1.045 NRD=11.076 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_A_186_21#_M1003_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.128375 PD=1.82 PS=1.045 NRD=0 NRS=22.152 M=1 R=4.33333
+ SA=75001.1 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_518_47#_M1004_d N_A_27_93#_M1004_g N_A_186_21#_M1004_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.121875 AS=0.169 PD=1.025 PS=1.82 NRD=9.228 NRS=0 M=1
+ R=4.33333 SA=75000.2 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g N_A_518_47#_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.121875 PD=0.92 PS=1.025 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1007 N_A_518_47#_M1007_d N_A1_M1007_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_B1_N_M1005_g N_A_27_93#_M1005_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0904183 AS=0.1134 PD=0.801549 PS=1.38 NRD=75.1752 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90003.1 A=0.0756 P=1.2 MULT=1
MM1000 N_VPWR_M1005_d N_A_186_21#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.215282 AS=0.1575 PD=1.90845 PS=1.315 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.4 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A_186_21#_M1008_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.3925 AS=0.1575 PD=1.785 PS=1.315 NRD=0.9653 NRS=5.8903 M=1 R=5.55556
+ SA=90000.9 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1001 N_A_186_21#_M1001_d N_A_27_93#_M1001_g N_VPWR_M1008_d VPB PHIGHVT L=0.18
+ W=1 AD=0.1725 AS=0.3925 PD=1.345 PS=1.785 NRD=11.8003 NRS=8.8453 M=1 R=5.55556
+ SA=90001.9 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1010 A_621_297# N_A2_M1010_g N_A_186_21#_M1001_d VPB PHIGHVT L=0.18 W=1
+ AD=0.1175 AS=0.1725 PD=1.235 PS=1.345 NRD=12.2928 NRS=0.9653 M=1 R=5.55556
+ SA=90002.4 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g A_621_297# VPB PHIGHVT L=0.18 W=1 AD=0.29
+ AS=0.1175 PD=2.58 PS=1.235 NRD=0.9653 NRS=12.2928 M=1 R=5.55556 SA=90002.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
pX13_noxref noxref_13 A2 A2 PROBETYPE=1
c_69 VPB 0 1.78374e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__o21ba_2.pxi.spice"
*
.ends
*
*
