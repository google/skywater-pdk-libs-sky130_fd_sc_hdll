* File: sky130_fd_sc_hdll__dlxtn_2.spice
* Created: Wed Sep  2 08:30:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__dlxtn_2.pex.spice"
.subckt sky130_fd_sc_hdll__dlxtn_2  VNB VPB GATE_N D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* GATE_N	GATE_N
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_GATE_N_M1015_g N_A_27_47#_M1015_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1000 N_A_211_363#_M1000_d N_A_27_47#_M1000_g N_VGND_M1015_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0672 PD=1.36 PS=0.74 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_D_M1009_g N_A_319_47#_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1006 A_505_47# N_A_319_47#_M1006_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0836769 AS=0.0672 PD=0.872308 PS=0.74 NRD=41.208 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1013 N_A_608_413#_M1013_d N_A_27_47#_M1013_g A_505_47# VNB NSHORT L=0.15
+ W=0.36 AD=0.0675 AS=0.0717231 PD=0.735 PS=0.747692 NRD=14.988 NRS=48.072 M=1
+ R=2.4 SA=75001.2 SB=75001.2 A=0.054 P=1.02 MULT=1
MM1001 A_718_47# N_A_211_363#_M1001_g N_A_608_413#_M1013_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0609231 AS=0.0675 PD=0.687692 PS=0.735 NRD=38.076 NRS=16.656 M=1
+ R=2.4 SA=75001.8 SB=75000.7 A=0.054 P=1.02 MULT=1
MM1011 N_VGND_M1011_d N_A_783_21#_M1011_g A_718_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0710769 PD=1.46 PS=0.802308 NRD=12.852 NRS=32.628 M=1 R=2.8
+ SA=75001.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_608_413#_M1014_g N_A_783_21#_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.2015 PD=0.97 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1014_d N_A_783_21#_M1007_g N_Q_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A_783_21#_M1008_g N_Q_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.104 PD=1.82 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_GATE_N_M1002_g N_A_27_47#_M1002_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1016 N_A_211_363#_M1016_d N_A_27_47#_M1016_g N_VPWR_M1002_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1010 N_VPWR_M1010_d N_D_M1010_g N_A_319_47#_M1010_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90001.7 A=0.1152 P=1.64 MULT=1
MM1003 A_503_369# N_A_319_47#_M1003_g N_VPWR_M1010_d VPB PHIGHVT L=0.18 W=0.64
+ AD=0.122023 AS=0.0928 PD=1.18943 PS=0.93 NRD=41.7443 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90001.2 A=0.1152 P=1.64 MULT=1
MM1018 N_A_608_413#_M1018_d N_A_211_363#_M1018_g A_503_369# VPB PHIGHVT L=0.18
+ W=0.42 AD=0.09975 AS=0.0800774 PD=0.895 PS=0.780566 NRD=60.9715 NRS=63.631 M=1
+ R=2.33333 SA=90001.2 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1005 A_739_413# N_A_27_47#_M1005_g N_A_608_413#_M1018_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0483 AS=0.09975 PD=0.65 PS=0.895 NRD=28.1316 NRS=30.4759 M=1
+ R=2.33333 SA=90001.8 SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1019 N_VPWR_M1019_d N_A_783_21#_M1019_g A_739_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.1134 AS=0.0483 PD=1.38 PS=0.65 NRD=2.3443 NRS=28.1316 M=1 R=2.33333
+ SA=90002.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1017 N_VPWR_M1017_d N_A_608_413#_M1017_g N_A_783_21#_M1017_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.2 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1017_d N_A_783_21#_M1004_g N_Q_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_A_783_21#_M1012_g N_Q_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.9461 P=16.85
c_130 VPB 0 1.7336e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__dlxtn_2.pxi.spice"
*
.ends
*
*
