* File: sky130_fd_sc_hdll__sdfxtp_2.spice
* Created: Wed Sep  2 08:52:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__sdfxtp_2.pex.spice"
.subckt sky130_fd_sc_hdll__sdfxtp_2  VNB VPB CLK SCE D SCD VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SCD	SCD
* D	D
* SCE	SCE
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1031 N_VGND_M1031_d N_CLK_M1031_g N_A_27_47#_M1031_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1092 PD=0.74 PS=1.36 NRD=12.852 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_A_203_47#_M1009_d N_A_27_47#_M1009_g N_VGND_M1031_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1302 AS=0.0672 PD=1.46 PS=0.74 NRD=12.852 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_SCE_M1014_g N_A_319_47#_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0861 AS=0.1176 PD=0.83 PS=1.4 NRD=35.712 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1017 A_517_47# N_A_319_47#_M1017_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0714 AS=0.0861 PD=0.76 PS=0.83 NRD=32.856 NRS=1.428 M=1 R=2.8 SA=75000.8
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_608_369#_M1002_d N_D_M1002_g A_517_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.0714 PD=0.8 PS=0.76 NRD=14.28 NRS=32.856 M=1 R=2.8 SA=75001.3
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1032 A_721_47# N_SCE_M1032_g N_A_608_369#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0483 AS=0.0798 PD=0.65 PS=0.8 NRD=17.136 NRS=14.28 M=1 R=2.8 SA=75001.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_SCD_M1025_g A_721_47# VNB NSHORT L=0.15 W=0.42 AD=0.1512
+ AS=0.0483 PD=1.56 PS=0.65 NRD=21.42 NRS=17.136 M=1 R=2.8 SA=75002.2 SB=75000.3
+ A=0.063 P=1.14 MULT=1
MM1030 N_A_1011_47#_M1030_d N_A_27_47#_M1030_g N_A_608_369#_M1030_s VNB NSHORT
+ L=0.15 W=0.36 AD=0.0774 AS=0.1008 PD=0.79 PS=1.28 NRD=34.992 NRS=4.992 M=1
+ R=2.4 SA=75000.2 SB=75003.8 A=0.054 P=1.02 MULT=1
MM1018 A_1127_47# N_A_203_47#_M1018_g N_A_1011_47#_M1030_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0731077 AS=0.0774 PD=0.747692 PS=0.79 NRD=49.356 NRS=14.988 M=1
+ R=2.4 SA=75000.8 SB=75003.2 A=0.054 P=1.02 MULT=1
MM1007 N_VGND_M1007_d N_A_1189_183#_M1007_g A_1127_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.130992 AS=0.0852923 PD=1.00642 PS=0.872308 NRD=47.136 NRS=42.3 M=1 R=2.8
+ SA=75001.2 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1028 N_A_1189_183#_M1028_d N_A_1011_47#_M1028_g N_VGND_M1007_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.126592 AS=0.199608 PD=1.2736 PS=1.53358 NRD=4.68 NRS=34.68
+ M=1 R=4.26667 SA=75001.4 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1013 N_A_1474_413#_M1013_d N_A_203_47#_M1013_g N_A_1189_183#_M1028_d VNB
+ NSHORT L=0.15 W=0.36 AD=0.0927 AS=0.071208 PD=0.875 PS=0.7164 NRD=43.332
+ NRS=16.656 M=1 R=2.4 SA=75002.6 SB=75001.4 A=0.054 P=1.02 MULT=1
MM1023 A_1625_47# N_A_27_47#_M1023_g N_A_1474_413#_M1013_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0609231 AS=0.0927 PD=0.687692 PS=0.875 NRD=38.076 NRS=34.992 M=1
+ R=2.4 SA=75003.3 SB=75000.7 A=0.054 P=1.02 MULT=1
MM1006 N_VGND_M1006_d N_A_1667_315#_M1006_g A_1625_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0710769 PD=1.46 PS=0.802308 NRD=12.852 NRS=32.628 M=1 R=2.8
+ SA=75003.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_1474_413#_M1016_g N_A_1667_315#_M1016_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=8.304 M=1
+ R=4.33333 SA=75000.2 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1016_d N_A_1667_315#_M1005_g N_Q_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1015_d N_A_1667_315#_M1015_g N_Q_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.21125 AS=0.12025 PD=1.95 PS=1.02 NRD=6.456 NRS=8.304 M=1 R=4.33333
+ SA=75001.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_CLK_M1001_g N_A_27_47#_M1001_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1022 N_A_203_47#_M1022_d N_A_27_47#_M1022_g N_VPWR_M1001_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1011 N_VPWR_M1011_d N_SCE_M1011_g N_A_319_47#_M1011_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90002.2 A=0.1152 P=1.64 MULT=1
MM1008 A_504_369# N_SCE_M1008_g N_VPWR_M1011_d VPB PHIGHVT L=0.18 W=0.64
+ AD=0.1088 AS=0.0928 PD=0.98 PS=0.93 NRD=35.3812 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90001.7 A=0.1152 P=1.64 MULT=1
MM1033 N_A_608_369#_M1033_d N_D_M1033_g A_504_369# VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.1088 PD=0.93 PS=0.98 NRD=1.5366 NRS=35.3812 M=1 R=3.55556
+ SA=90001.2 SB=90001.2 A=0.1152 P=1.64 MULT=1
MM1027 A_702_369# N_A_319_47#_M1027_g N_A_608_369#_M1033_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1072 AS=0.0928 PD=0.975 PS=0.93 NRD=34.6129 NRS=1.5366 M=1
+ R=3.55556 SA=90001.6 SB=90000.7 A=0.1152 P=1.64 MULT=1
MM1024 N_VPWR_M1024_d N_SCD_M1024_g A_702_369# VPB PHIGHVT L=0.18 W=0.64
+ AD=0.1888 AS=0.1072 PD=1.87 PS=0.975 NRD=9.2196 NRS=34.6129 M=1 R=3.55556
+ SA=90002.2 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1021 N_A_1011_47#_M1021_d N_A_203_47#_M1021_g N_A_608_369#_M1021_s VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.07035 AS=0.1344 PD=0.755 PS=1.48 NRD=14.0658 NRS=25.7873
+ M=1 R=2.33333 SA=90000.2 SB=90003.7 A=0.0756 P=1.2 MULT=1
MM1012 A_1121_413# N_A_27_47#_M1012_g N_A_1011_47#_M1021_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0735 AS=0.07035 PD=0.77 PS=0.755 NRD=56.2829 NRS=11.7215 M=1
+ R=2.33333 SA=90000.7 SB=90003.2 A=0.0756 P=1.2 MULT=1
MM1000 N_VPWR_M1000_d N_A_1189_183#_M1000_g A_1121_413# VPB PHIGHVT L=0.18
+ W=0.42 AD=0.132623 AS=0.0735 PD=0.918974 PS=0.77 NRD=116.072 NRS=56.2829 M=1
+ R=2.33333 SA=90001.3 SB=90002.7 A=0.0756 P=1.2 MULT=1
MM1019 N_A_1189_183#_M1019_d N_A_1011_47#_M1019_g N_VPWR_M1000_d VPB PHIGHVT
+ L=0.18 W=0.75 AD=0.147885 AS=0.236827 PD=1.40385 PS=1.64103 NRD=1.3002
+ NRS=1.3002 M=1 R=4.16667 SA=90001.3 SB=90001.2 A=0.135 P=1.86 MULT=1
MM1003 N_A_1474_413#_M1003_d N_A_27_47#_M1003_g N_A_1189_183#_M1019_d VPB
+ PHIGHVT L=0.18 W=0.42 AD=0.0609 AS=0.0828154 PD=0.71 PS=0.786154 NRD=2.3443
+ NRS=28.1316 M=1 R=2.33333 SA=90002.5 SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1029 A_1568_413# N_A_203_47#_M1029_g N_A_1474_413#_M1003_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.10605 AS=0.0609 PD=0.925 PS=0.71 NRD=92.6294 NRS=2.3443 M=1
+ R=2.33333 SA=90003 SB=90001 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_A_1667_315#_M1010_g A_1568_413# VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1617 AS=0.10605 PD=1.61 PS=0.925 NRD=53.9386 NRS=92.6294 M=1
+ R=2.33333 SA=90003.7 SB=90000.3 A=0.0756 P=1.2 MULT=1
MM1026 N_VPWR_M1026_d N_A_1474_413#_M1026_g N_A_1667_315#_M1026_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1026_d N_A_1667_315#_M1004_g N_Q_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1020 N_VPWR_M1020_d N_A_1667_315#_M1020_g N_Q_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.33 AS=0.145 PD=2.66 PS=1.29 NRD=8.8453 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.2 A=0.18 P=2.36 MULT=1
DX34_noxref VNB VPB NWDIODE A=18.3291 P=26.05
c_103 VNB 0 4.47538e-20 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hdll__sdfxtp_2.pxi.spice"
*
.ends
*
*
