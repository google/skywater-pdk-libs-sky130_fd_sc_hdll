# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__ebufn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__ebufn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.355000 1.615000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.358200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.960000 1.075000 1.290000 1.630000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.700500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.125000 1.495000 3.585000 2.465000 ;
        RECT 3.255000 0.255000 3.585000 0.825000 ;
        RECT 3.315000 0.825000 3.585000 1.495000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT -0.005000  2.635000 3.680000 2.805000 ;
      RECT  0.000000 -0.085000 3.680000 0.085000 ;
      RECT  0.085000  0.280000 0.345000 0.615000 ;
      RECT  0.085000  0.615000 1.235000 0.825000 ;
      RECT  0.085000  1.785000 0.790000 2.005000 ;
      RECT  0.085000  2.005000 0.345000 2.465000 ;
      RECT  0.515000  0.085000 0.895000 0.445000 ;
      RECT  0.515000  2.175000 0.890000 2.635000 ;
      RECT  0.525000  0.825000 0.790000 1.785000 ;
      RECT  1.065000  0.255000 2.175000 0.465000 ;
      RECT  1.065000  0.465000 1.235000 0.615000 ;
      RECT  1.115000  1.800000 1.905000 2.005000 ;
      RECT  1.115000  2.005000 1.370000 2.460000 ;
      RECT  1.460000  0.635000 1.790000 1.075000 ;
      RECT  1.460000  1.075000 2.745000 1.325000 ;
      RECT  1.460000  1.325000 1.905000 1.800000 ;
      RECT  1.540000  2.175000 1.900000 2.635000 ;
      RECT  1.960000  0.465000 2.175000 0.735000 ;
      RECT  1.960000  0.735000 3.085000 0.905000 ;
      RECT  2.345000  0.085000 3.085000 0.565000 ;
      RECT  2.915000  0.905000 3.085000 0.995000 ;
      RECT  2.915000  0.995000 3.145000 1.325000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__ebufn_1
END LIBRARY
