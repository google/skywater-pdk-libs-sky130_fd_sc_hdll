* File: sky130_fd_sc_hdll__sdfxtp_1.pxi.spice
* Created: Wed Sep  2 08:52:21 2020
* 
x_PM_SKY130_FD_SC_HDLL__SDFXTP_1%CLK N_CLK_c_194_n N_CLK_c_198_n N_CLK_c_195_n
+ N_CLK_M1028_g N_CLK_c_199_n N_CLK_M1002_g CLK
+ PM_SKY130_FD_SC_HDLL__SDFXTP_1%CLK
x_PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_27_47# N_A_27_47#_M1028_s N_A_27_47#_M1002_s
+ N_A_27_47#_M1007_g N_A_27_47#_c_244_n N_A_27_47#_c_245_n N_A_27_47#_M1017_g
+ N_A_27_47#_M1026_g N_A_27_47#_c_234_n N_A_27_47#_c_235_n N_A_27_47#_c_248_n
+ N_A_27_47#_c_249_n N_A_27_47#_M1011_g N_A_27_47#_c_250_n N_A_27_47#_c_251_n
+ N_A_27_47#_M1004_g N_A_27_47#_c_236_n N_A_27_47#_M1027_g N_A_27_47#_c_451_p
+ N_A_27_47#_c_238_n N_A_27_47#_c_239_n N_A_27_47#_c_253_n N_A_27_47#_c_359_p
+ N_A_27_47#_c_240_n N_A_27_47#_c_255_n N_A_27_47#_c_256_n N_A_27_47#_c_257_n
+ N_A_27_47#_c_258_n N_A_27_47#_c_259_n N_A_27_47#_c_260_n N_A_27_47#_c_261_n
+ N_A_27_47#_c_241_n N_A_27_47#_c_242_n N_A_27_47#_c_243_n
+ PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__SDFXTP_1%SCE N_SCE_c_470_n N_SCE_M1009_g N_SCE_M1013_g
+ N_SCE_c_472_n N_SCE_M1006_g N_SCE_M1029_g N_SCE_c_465_n N_SCE_c_466_n SCE
+ N_SCE_c_473_n N_SCE_c_467_n N_SCE_c_468_n SCE
+ PM_SKY130_FD_SC_HDLL__SDFXTP_1%SCE
x_PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_319_47# N_A_319_47#_M1013_s
+ N_A_319_47#_M1009_s N_A_319_47#_M1021_g N_A_319_47#_c_565_n
+ N_A_319_47#_M1022_g N_A_319_47#_c_560_n N_A_319_47#_c_567_n
+ N_A_319_47#_c_573_n N_A_319_47#_c_561_n N_A_319_47#_c_575_n
+ N_A_319_47#_c_569_n N_A_319_47#_c_562_n N_A_319_47#_c_570_n
+ N_A_319_47#_c_563_n N_A_319_47#_c_564_n N_A_319_47#_c_580_n
+ PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_319_47#
x_PM_SKY130_FD_SC_HDLL__SDFXTP_1%D N_D_c_675_n N_D_M1030_g N_D_M1003_g D D
+ PM_SKY130_FD_SC_HDLL__SDFXTP_1%D
x_PM_SKY130_FD_SC_HDLL__SDFXTP_1%SCD N_SCD_M1020_g N_SCD_c_717_n N_SCD_c_718_n
+ N_SCD_M1019_g SCD N_SCD_c_716_n PM_SKY130_FD_SC_HDLL__SDFXTP_1%SCD
x_PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_203_47# N_A_203_47#_M1007_d
+ N_A_203_47#_M1017_d N_A_203_47#_c_781_n N_A_203_47#_M1014_g
+ N_A_203_47#_M1023_g N_A_203_47#_M1018_g N_A_203_47#_c_782_n
+ N_A_203_47#_M1015_g N_A_203_47#_c_767_n N_A_203_47#_c_768_n
+ N_A_203_47#_c_769_n N_A_203_47#_c_770_n N_A_203_47#_c_771_n
+ N_A_203_47#_c_772_n N_A_203_47#_c_773_n N_A_203_47#_c_774_n
+ N_A_203_47#_c_775_n N_A_203_47#_c_776_n N_A_203_47#_c_777_n
+ N_A_203_47#_c_778_n N_A_203_47#_c_779_n N_A_203_47#_c_780_n
+ PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_203_47#
x_PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_1189_21# N_A_1189_21#_M1012_d
+ N_A_1189_21#_M1025_d N_A_1189_21#_M1005_g N_A_1189_21#_c_969_n
+ N_A_1189_21#_c_975_n N_A_1189_21#_M1000_g N_A_1189_21#_c_970_n
+ N_A_1189_21#_c_971_n N_A_1189_21#_c_998_n N_A_1189_21#_c_972_n
+ N_A_1189_21#_c_1002_n N_A_1189_21#_c_973_n
+ PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_1189_21#
x_PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_1011_47# N_A_1011_47#_M1026_d
+ N_A_1011_47#_M1014_d N_A_1011_47#_c_1064_n N_A_1011_47#_M1025_g
+ N_A_1011_47#_M1012_g N_A_1011_47#_c_1061_n N_A_1011_47#_c_1062_n
+ N_A_1011_47#_c_1076_n N_A_1011_47#_c_1080_n N_A_1011_47#_c_1063_n
+ N_A_1011_47#_c_1067_n N_A_1011_47#_c_1068_n N_A_1011_47#_c_1069_n
+ PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_1011_47#
x_PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_1647_21# N_A_1647_21#_M1001_s
+ N_A_1647_21#_M1024_s N_A_1647_21#_M1008_g N_A_1647_21#_c_1170_n
+ N_A_1647_21#_M1010_g N_A_1647_21#_c_1164_n N_A_1647_21#_M1031_g
+ N_A_1647_21#_c_1165_n N_A_1647_21#_M1016_g N_A_1647_21#_c_1172_n
+ N_A_1647_21#_c_1182_p N_A_1647_21#_c_1166_n N_A_1647_21#_c_1173_n
+ N_A_1647_21#_c_1167_n N_A_1647_21#_c_1168_n N_A_1647_21#_c_1184_p
+ N_A_1647_21#_c_1192_p PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_1647_21#
x_PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_1474_413# N_A_1474_413#_M1018_d
+ N_A_1474_413#_M1004_d N_A_1474_413#_c_1253_n N_A_1474_413#_M1024_g
+ N_A_1474_413#_c_1247_n N_A_1474_413#_M1001_g N_A_1474_413#_c_1248_n
+ N_A_1474_413#_c_1249_n N_A_1474_413#_c_1258_n N_A_1474_413#_c_1261_n
+ N_A_1474_413#_c_1250_n N_A_1474_413#_c_1256_n N_A_1474_413#_c_1251_n
+ N_A_1474_413#_c_1252_n PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_1474_413#
x_PM_SKY130_FD_SC_HDLL__SDFXTP_1%VPWR N_VPWR_M1002_d N_VPWR_M1009_d
+ N_VPWR_M1019_d N_VPWR_M1000_d N_VPWR_M1010_d N_VPWR_M1024_d N_VPWR_c_1333_n
+ N_VPWR_c_1334_n N_VPWR_c_1335_n N_VPWR_c_1336_n N_VPWR_c_1337_n
+ N_VPWR_c_1338_n N_VPWR_c_1339_n N_VPWR_c_1340_n N_VPWR_c_1341_n
+ N_VPWR_c_1342_n N_VPWR_c_1343_n N_VPWR_c_1344_n VPWR N_VPWR_c_1345_n
+ N_VPWR_c_1346_n N_VPWR_c_1347_n N_VPWR_c_1348_n N_VPWR_c_1332_n
+ N_VPWR_c_1350_n N_VPWR_c_1351_n N_VPWR_c_1352_n
+ PM_SKY130_FD_SC_HDLL__SDFXTP_1%VPWR
x_PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_608_369# N_A_608_369#_M1003_d
+ N_A_608_369#_M1026_s N_A_608_369#_M1030_d N_A_608_369#_M1014_s
+ N_A_608_369#_c_1495_n N_A_608_369#_c_1507_n N_A_608_369#_c_1519_n
+ N_A_608_369#_c_1484_n N_A_608_369#_c_1491_n N_A_608_369#_c_1492_n
+ N_A_608_369#_c_1485_n N_A_608_369#_c_1486_n N_A_608_369#_c_1487_n
+ N_A_608_369#_c_1488_n N_A_608_369#_c_1489_n N_A_608_369#_c_1490_n
+ N_A_608_369#_c_1494_n PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_608_369#
x_PM_SKY130_FD_SC_HDLL__SDFXTP_1%Q N_Q_M1031_d N_Q_M1016_d N_Q_c_1607_n Q Q
+ N_Q_c_1610_n N_Q_c_1608_n PM_SKY130_FD_SC_HDLL__SDFXTP_1%Q
x_PM_SKY130_FD_SC_HDLL__SDFXTP_1%VGND N_VGND_M1028_d N_VGND_M1013_d
+ N_VGND_M1020_d N_VGND_M1005_d N_VGND_M1008_d N_VGND_M1001_d N_VGND_c_1633_n
+ N_VGND_c_1634_n N_VGND_c_1635_n N_VGND_c_1636_n N_VGND_c_1637_n
+ N_VGND_c_1638_n N_VGND_c_1639_n N_VGND_c_1640_n N_VGND_c_1641_n
+ N_VGND_c_1642_n N_VGND_c_1643_n N_VGND_c_1644_n N_VGND_c_1645_n VGND
+ N_VGND_c_1646_n N_VGND_c_1647_n N_VGND_c_1648_n N_VGND_c_1649_n
+ N_VGND_c_1650_n N_VGND_c_1651_n PM_SKY130_FD_SC_HDLL__SDFXTP_1%VGND
cc_1 VNB N_CLK_c_194_n 0.0583772f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.325
cc_2 VNB N_CLK_c_195_n 0.0176355f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_3 VNB CLK 0.0188196f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_27_47#_M1007_g 0.0375848f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_5 VNB N_A_27_47#_M1026_g 0.0532273f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_c_234_n 0.0172606f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_235_n 0.00252324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_236_n 0.0103696f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1027_g 0.0447949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_238_n 0.00363705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_239_n 0.00651432f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_240_n 0.0026153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_241_n 0.0271693f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_242_n 0.0072594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_243_n 0.00135089f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_SCE_M1013_g 0.0532415f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.74
cc_17 VNB N_SCE_M1029_g 0.0173106f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_18 VNB N_SCE_c_465_n 0.00779079f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_19 VNB N_SCE_c_466_n 0.00118673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_SCE_c_467_n 0.0324407f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_SCE_c_468_n 0.0011318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB SCE 0.00871703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_319_47#_M1021_g 0.021567f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_24 VNB N_A_319_47#_c_560_n 0.0140321f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_25 VNB N_A_319_47#_c_561_n 0.00231465f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_319_47#_c_562_n 0.0025595f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_319_47#_c_563_n 0.00277032f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_319_47#_c_564_n 0.0333689f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_D_M1003_g 0.0465924f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.74
cc_30 VNB N_SCD_M1020_g 0.0452314f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_31 VNB SCD 0.0074008f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_SCD_c_716_n 0.0152332f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_33 VNB N_A_203_47#_c_767_n 0.00343716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_203_47#_c_768_n 0.00526411f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_203_47#_c_769_n 0.00696616f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_203_47#_c_770_n 0.00523362f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_203_47#_c_771_n 0.0540748f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_203_47#_c_772_n 0.00194843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_203_47#_c_773_n 0.00182186f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_203_47#_c_774_n 0.0116233f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_203_47#_c_775_n 0.0282254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_203_47#_c_776_n 0.00514406f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_203_47#_c_777_n 0.0181899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_203_47#_c_778_n 0.0285365f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_203_47#_c_779_n 0.0182472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_203_47#_c_780_n 0.0160413f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_1189_21#_M1005_g 0.0212905f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_48 VNB N_A_1189_21#_c_969_n 0.0164066f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_1189_21#_c_970_n 0.00853932f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_50 VNB N_A_1189_21#_c_971_n 0.030045f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_1189_21#_c_972_n 0.00469491f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_1189_21#_c_973_n 0.00263218f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_1011_47#_M1012_g 0.03597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1011_47#_c_1061_n 0.00817418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_1011_47#_c_1062_n 0.00258415f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_56 VNB N_A_1011_47#_c_1063_n 0.0122681f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1647_21#_M1008_g 0.0529975f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_58 VNB N_A_1647_21#_c_1164_n 0.0196808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_1647_21#_c_1165_n 0.0231286f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_60 VNB N_A_1647_21#_c_1166_n 0.00377099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_1647_21#_c_1167_n 0.00574146f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_1647_21#_c_1168_n 0.00767738f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1474_413#_c_1247_n 0.0201839f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_1474_413#_c_1248_n 0.0410187f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.105
cc_65 VNB N_A_1474_413#_c_1249_n 0.0119893f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1474_413#_c_1250_n 0.00211001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1474_413#_c_1251_n 0.0099142f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1474_413#_c_1252_n 0.00193332f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VPWR_c_1332_n 0.440529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_608_369#_c_1484_n 2.48589e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_608_369#_c_1485_n 0.0157766f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_608_369#_c_1486_n 0.00126846f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_608_369#_c_1487_n 0.00359021f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_608_369#_c_1488_n 0.0101757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_608_369#_c_1489_n 0.00249978f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_608_369#_c_1490_n 0.0017307f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_Q_c_1607_n 0.0257579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_Q_c_1608_n 0.0248899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1633_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1634_n 0.00491179f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1635_n 0.00586751f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1636_n 0.00554283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1637_n 0.0046831f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1638_n 0.0294925f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1639_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1640_n 0.0419197f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1641_n 0.00381885f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1642_n 0.0506248f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1643_n 0.00709041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1644_n 0.0229461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1645_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1646_n 0.0154125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1647_n 0.0484085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1648_n 0.0236473f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1649_n 0.505072f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1650_n 0.0055668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1651_n 0.00603399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VPB N_CLK_c_194_n 0.00482568f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_99 VPB N_CLK_c_198_n 0.0166215f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.59
cc_100 VPB N_CLK_c_199_n 0.0478608f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.74
cc_101 VPB CLK 0.018034f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_102 VPB N_A_27_47#_c_244_n 0.0165313f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_27_47#_c_245_n 0.0251878f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_104 VPB N_A_27_47#_c_234_n 0.0157747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_27_47#_c_235_n 0.0052974f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_27_47#_c_248_n 0.011717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_27_47#_c_249_n 0.050198f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_27_47#_c_250_n 0.0170508f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_27_47#_c_251_n 0.0233159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_27_47#_c_236_n 0.0181089f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_27_47#_c_253_n 0.00135894f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_27_47#_c_240_n 0.00368748f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_27_47#_c_255_n 0.00358354f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_27_47#_c_256_n 0.00307948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_27_47#_c_257_n 0.00818052f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_27_47#_c_258_n 0.0620921f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_27_47#_c_259_n 9.26987e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_27_47#_c_260_n 0.00534134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_27_47#_c_261_n 0.00183196f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_27_47#_c_241_n 0.0120872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_27_47#_c_242_n 0.020668f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_27_47#_c_243_n 0.00540204f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_SCE_c_470_n 0.0190803f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_124 VPB N_SCE_M1013_g 0.00578264f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.74
cc_125 VPB N_SCE_c_472_n 0.0160063f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=2.135
cc_126 VPB N_SCE_c_473_n 0.0613549f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB SCE 0.00370634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_319_47#_c_565_n 0.0483351f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.665
cc_129 VPB N_A_319_47#_c_560_n 0.0110715f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.16
cc_130 VPB N_A_319_47#_c_567_n 0.00408285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_319_47#_c_561_n 0.00568384f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_319_47#_c_569_n 0.00293027f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_319_47#_c_570_n 0.00183048f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_D_c_675_n 0.0489403f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_135 VPB N_D_M1003_g 0.0052563f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.74
cc_136 VPB D 0.00834963f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=2.135
cc_137 VPB N_SCD_c_717_n 0.00922874f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.74
cc_138 VPB N_SCD_c_718_n 0.0275598f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=2.135
cc_139 VPB SCD 0.0058351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_SCD_c_716_n 0.0201164f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_141 VPB N_A_203_47#_c_781_n 0.0628983f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=2.135
cc_142 VPB N_A_203_47#_c_782_n 0.0544866f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_143 VPB N_A_203_47#_c_767_n 0.00466902f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_203_47#_c_768_n 0.00454474f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_203_47#_c_780_n 0.0177947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_1189_21#_c_969_n 0.0312088f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_1189_21#_c_975_n 0.0244868f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_148 VPB N_A_1189_21#_c_972_n 0.0085277f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_1011_47#_c_1064_n 0.01851f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=2.135
cc_150 VPB N_A_1011_47#_c_1061_n 0.0178529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_1011_47#_c_1062_n 0.018702f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.16
cc_152 VPB N_A_1011_47#_c_1067_n 0.00177935f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_1011_47#_c_1068_n 0.00549416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_1011_47#_c_1069_n 0.00538019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_1647_21#_M1008_g 0.0228521f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_156 VPB N_A_1647_21#_c_1170_n 0.0686242f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.665
cc_157 VPB N_A_1647_21#_c_1165_n 0.028706f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_158 VPB N_A_1647_21#_c_1172_n 0.0129293f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_1647_21#_c_1173_n 0.00551938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_1647_21#_c_1167_n 0.00574146f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_1474_413#_c_1253_n 0.0198033f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=2.135
cc_162 VPB N_A_1474_413#_c_1248_n 0.0147613f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_163 VPB N_A_1474_413#_c_1249_n 0.00732521f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_1474_413#_c_1256_n 0.0055098f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_1474_413#_c_1251_n 0.00407395f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_1333_n 0.00126291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_1334_n 4.89699e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_1335_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_1336_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_1337_n 0.00548992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_1338_n 0.00471485f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_1339_n 0.0429455f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1340_n 0.00324297f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1341_n 0.0551677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1342_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1343_n 0.0234195f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1344_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1345_n 0.0156572f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1346_n 0.0270443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1347_n 0.0507262f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1348_n 0.0238235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1332_n 0.0637614f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1350_n 0.0054556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1351_n 0.00502699f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1352_n 0.00584025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_608_369#_c_1491_n 0.0113352f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_608_369#_c_1492_n 5.53729e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_608_369#_c_1488_n 0.0122437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_608_369#_c_1494_n 0.00885905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB Q 0.0288181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_Q_c_1610_n 0.0126746f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_Q_c_1608_n 0.0126124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 N_CLK_c_194_n N_A_27_47#_M1007_g 0.00437311f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_194 N_CLK_c_195_n N_A_27_47#_M1007_g 0.0161772f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_195 CLK N_A_27_47#_M1007_g 3.44553e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_196 N_CLK_c_198_n N_A_27_47#_c_244_n 0.004446f $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_197 N_CLK_c_199_n N_A_27_47#_c_244_n 0.00668506f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_198 CLK N_A_27_47#_c_244_n 6.27642e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_199 N_CLK_c_199_n N_A_27_47#_c_245_n 0.0192752f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_200 N_CLK_c_194_n N_A_27_47#_c_238_n 0.00788454f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_201 N_CLK_c_195_n N_A_27_47#_c_238_n 0.00700547f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_202 CLK N_A_27_47#_c_238_n 0.00774265f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_203 N_CLK_c_194_n N_A_27_47#_c_239_n 0.00622672f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_204 CLK N_A_27_47#_c_239_n 0.0144574f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_205 N_CLK_c_199_n N_A_27_47#_c_253_n 0.0171149f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_206 CLK N_A_27_47#_c_253_n 0.00731943f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_207 N_CLK_c_194_n N_A_27_47#_c_240_n 0.0045363f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_208 N_CLK_c_198_n N_A_27_47#_c_240_n 7.61846e-19 $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_209 N_CLK_c_199_n N_A_27_47#_c_240_n 0.0042845f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_210 CLK N_A_27_47#_c_240_n 0.0429434f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_211 N_CLK_c_194_n N_A_27_47#_c_255_n 2.26313e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_212 N_CLK_c_199_n N_A_27_47#_c_255_n 0.007998f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_213 CLK N_A_27_47#_c_255_n 0.0153364f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_214 N_CLK_c_199_n N_A_27_47#_c_256_n 0.00150514f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_215 N_CLK_c_194_n N_A_27_47#_c_241_n 0.0130887f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_216 CLK N_A_27_47#_c_241_n 0.00184424f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_217 N_CLK_c_199_n N_VPWR_c_1333_n 0.0125197f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_218 N_CLK_c_199_n N_VPWR_c_1345_n 0.00304525f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_219 N_CLK_c_199_n N_VPWR_c_1332_n 0.00455272f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_220 N_CLK_c_194_n N_VGND_c_1646_n 4.61451e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_221 N_CLK_c_195_n N_VGND_c_1646_n 0.00340075f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_222 N_CLK_c_195_n N_VGND_c_1649_n 0.00497799f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_223 N_CLK_c_195_n N_VGND_c_1650_n 0.0115525f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_224 N_A_27_47#_c_258_n N_SCE_c_470_n 0.00312335f $X=5.555 $Y=1.825 $X2=-0.19
+ $Y2=-0.24
cc_225 N_A_27_47#_c_258_n N_SCE_c_472_n 0.00201569f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_258_n N_SCE_c_473_n 0.00331869f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_258_n SCE 0.00858979f $X=5.555 $Y=1.825 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_258_n N_A_319_47#_c_565_n 0.00193553f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_229 N_A_27_47#_c_258_n N_A_319_47#_c_560_n 0.012706f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_258_n N_A_319_47#_c_573_n 0.0211859f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_258_n N_A_319_47#_c_561_n 0.00964382f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_232 N_A_27_47#_c_258_n N_A_319_47#_c_575_n 0.0361285f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_258_n N_A_319_47#_c_569_n 0.0135446f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_M1007_g N_A_319_47#_c_562_n 9.20042e-19 $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_258_n N_A_319_47#_c_570_n 0.0130533f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_258_n N_A_319_47#_c_564_n 0.00293413f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_237 N_A_27_47#_c_258_n N_A_319_47#_c_580_n 0.00491135f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_238 N_A_27_47#_c_258_n N_D_c_675_n 0.00616123f $X=5.555 $Y=1.825 $X2=-0.19
+ $Y2=-0.24
cc_239 N_A_27_47#_c_258_n D 0.0102464f $X=5.555 $Y=1.825 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_258_n N_SCD_c_718_n 0.00274884f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_258_n SCD 0.00910253f $X=5.555 $Y=1.825 $X2=0 $Y2=0
cc_242 N_A_27_47#_c_258_n N_SCD_c_716_n 0.0013799f $X=5.555 $Y=1.825 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_258_n N_A_203_47#_M1017_d 7.52281e-19 $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_244 N_A_27_47#_c_235_n N_A_203_47#_c_781_n 0.0194945f $X=5.055 $Y=1.32 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_249_n N_A_203_47#_c_781_n 0.0316637f $X=5.515 $Y=1.99 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_257_n N_A_203_47#_c_781_n 0.00224123f $X=5.75 $Y=1.825 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_258_n N_A_203_47#_c_781_n 0.0095879f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_250_n N_A_203_47#_c_782_n 0.0165967f $X=7.28 $Y=1.89 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_251_n N_A_203_47#_c_782_n 0.0113242f $X=7.28 $Y=1.99 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_236_n N_A_203_47#_c_782_n 0.0164015f $X=7.755 $Y=1.32 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_260_n N_A_203_47#_c_782_n 0.00420927f $X=7.325 $Y=1.825
+ $X2=0 $Y2=0
cc_252 N_A_27_47#_c_243_n N_A_203_47#_c_782_n 0.00257462f $X=7.315 $Y=1.41 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_M1026_g N_A_203_47#_c_767_n 0.00796706f $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_234_n N_A_203_47#_c_767_n 0.00904756f $X=5.415 $Y=1.32 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_235_n N_A_203_47#_c_767_n 0.00418731f $X=5.055 $Y=1.32 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_c_248_n N_A_203_47#_c_767_n 0.00637651f $X=5.515 $Y=1.575
+ $X2=0 $Y2=0
cc_257 N_A_27_47#_c_249_n N_A_203_47#_c_767_n 7.35344e-19 $X=5.515 $Y=1.99 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_c_257_n N_A_203_47#_c_767_n 0.0169317f $X=5.75 $Y=1.825 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_258_n N_A_203_47#_c_767_n 0.0161657f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_259_n N_A_203_47#_c_767_n 4.35179e-19 $X=5.895 $Y=1.825
+ $X2=0 $Y2=0
cc_261 N_A_27_47#_c_250_n N_A_203_47#_c_768_n 4.64672e-19 $X=7.28 $Y=1.89 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_236_n N_A_203_47#_c_768_n 0.00774933f $X=7.755 $Y=1.32 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_M1027_g N_A_203_47#_c_768_n 0.00700265f $X=7.83 $Y=0.415 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_260_n N_A_203_47#_c_768_n 0.00568845f $X=7.325 $Y=1.825
+ $X2=0 $Y2=0
cc_265 N_A_27_47#_c_242_n N_A_203_47#_c_768_n 0.00113444f $X=7.315 $Y=1.32 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_c_243_n N_A_203_47#_c_768_n 0.0330587f $X=7.315 $Y=1.41 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_236_n N_A_203_47#_c_769_n 0.00853729f $X=7.755 $Y=1.32 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_M1027_g N_A_203_47#_c_769_n 0.0121341f $X=7.83 $Y=0.415 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_242_n N_A_203_47#_c_769_n 2.74628e-19 $X=7.315 $Y=1.32 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_243_n N_A_203_47#_c_769_n 0.0133202f $X=7.315 $Y=1.41 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_M1007_g N_A_203_47#_c_770_n 0.00640849f $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_238_n N_A_203_47#_c_770_n 0.00344258f $X=0.665 $Y=0.72 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_240_n N_A_203_47#_c_770_n 0.00374014f $X=0.81 $Y=1.235 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_M1026_g N_A_203_47#_c_771_n 0.00225641f $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_M1026_g N_A_203_47#_c_772_n 3.50278e-19 $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_M1027_g N_A_203_47#_c_773_n 2.47228e-19 $X=7.83 $Y=0.415 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_243_n N_A_203_47#_c_773_n 0.00207442f $X=7.315 $Y=1.41 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_234_n N_A_203_47#_c_774_n 0.00102588f $X=5.415 $Y=1.32 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_242_n N_A_203_47#_c_774_n 0.0012618f $X=7.315 $Y=1.32 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_M1026_g N_A_203_47#_c_775_n 0.016368f $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_234_n N_A_203_47#_c_775_n 0.0189929f $X=5.415 $Y=1.32 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_257_n N_A_203_47#_c_775_n 4.31662e-19 $X=5.75 $Y=1.825 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_M1026_g N_A_203_47#_c_776_n 0.0122484f $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_234_n N_A_203_47#_c_776_n 0.00609027f $X=5.415 $Y=1.32 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_257_n N_A_203_47#_c_776_n 0.00398178f $X=5.75 $Y=1.825 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_M1026_g N_A_203_47#_c_777_n 0.0140838f $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_M1027_g N_A_203_47#_c_778_n 0.0167626f $X=7.83 $Y=0.415 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_242_n N_A_203_47#_c_778_n 0.0176132f $X=7.315 $Y=1.32 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_243_n N_A_203_47#_c_778_n 9.7768e-19 $X=7.315 $Y=1.41 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_M1027_g N_A_203_47#_c_779_n 0.0145692f $X=7.83 $Y=0.415 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_M1007_g N_A_203_47#_c_780_n 0.0133504f $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_245_n N_A_203_47#_c_780_n 0.00212706f $X=0.97 $Y=1.74 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_238_n N_A_203_47#_c_780_n 0.00981189f $X=0.665 $Y=0.72 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_359_p N_A_203_47#_c_780_n 0.006717f $X=0.78 $Y=1.795 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_240_n N_A_203_47#_c_780_n 0.0584555f $X=0.81 $Y=1.235 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_256_n N_A_203_47#_c_780_n 0.00207039f $X=0.895 $Y=1.825
+ $X2=0 $Y2=0
cc_297 N_A_27_47#_c_258_n N_A_203_47#_c_780_n 0.0255099f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_241_n N_A_203_47#_c_780_n 0.0167016f $X=0.97 $Y=1.235 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_261_n N_A_1189_21#_M1025_d 0.00343409f $X=7.13 $Y=1.825
+ $X2=0 $Y2=0
cc_300 N_A_27_47#_c_234_n N_A_1189_21#_c_969_n 0.0116076f $X=5.415 $Y=1.32 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_249_n N_A_1189_21#_c_969_n 0.0209627f $X=5.515 $Y=1.99 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_257_n N_A_1189_21#_c_969_n 0.00212256f $X=5.75 $Y=1.825
+ $X2=0 $Y2=0
cc_303 N_A_27_47#_c_259_n N_A_1189_21#_c_969_n 0.00152496f $X=5.895 $Y=1.825
+ $X2=0 $Y2=0
cc_304 N_A_27_47#_c_261_n N_A_1189_21#_c_969_n 0.00150072f $X=7.13 $Y=1.825
+ $X2=0 $Y2=0
cc_305 N_A_27_47#_c_249_n N_A_1189_21#_c_975_n 0.0264165f $X=5.515 $Y=1.99 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_261_n N_A_1189_21#_c_975_n 0.00126931f $X=7.13 $Y=1.825
+ $X2=0 $Y2=0
cc_307 N_A_27_47#_c_251_n N_A_1189_21#_c_972_n 0.00848935f $X=7.28 $Y=1.99 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_M1027_g N_A_1189_21#_c_972_n 7.19355e-19 $X=7.83 $Y=0.415
+ $X2=0 $Y2=0
cc_309 N_A_27_47#_c_260_n N_A_1189_21#_c_972_n 0.00297493f $X=7.325 $Y=1.825
+ $X2=0 $Y2=0
cc_310 N_A_27_47#_c_261_n N_A_1189_21#_c_972_n 0.0235945f $X=7.13 $Y=1.825 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_242_n N_A_1189_21#_c_972_n 0.00581535f $X=7.315 $Y=1.32
+ $X2=0 $Y2=0
cc_312 N_A_27_47#_c_243_n N_A_1189_21#_c_972_n 0.0513894f $X=7.315 $Y=1.41 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_M1027_g N_A_1189_21#_c_973_n 4.17953e-19 $X=7.83 $Y=0.415
+ $X2=0 $Y2=0
cc_314 N_A_27_47#_c_250_n N_A_1011_47#_c_1064_n 0.01106f $X=7.28 $Y=1.89 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_251_n N_A_1011_47#_c_1064_n 0.0127283f $X=7.28 $Y=1.99 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_261_n N_A_1011_47#_c_1064_n 0.0108509f $X=7.13 $Y=1.825
+ $X2=0 $Y2=0
cc_317 N_A_27_47#_c_242_n N_A_1011_47#_M1012_g 0.00626018f $X=7.315 $Y=1.32
+ $X2=0 $Y2=0
cc_318 N_A_27_47#_c_250_n N_A_1011_47#_c_1062_n 0.00626018f $X=7.28 $Y=1.89
+ $X2=0 $Y2=0
cc_319 N_A_27_47#_c_261_n N_A_1011_47#_c_1062_n 5.36013e-19 $X=7.13 $Y=1.825
+ $X2=0 $Y2=0
cc_320 N_A_27_47#_c_249_n N_A_1011_47#_c_1076_n 0.0105456f $X=5.515 $Y=1.99
+ $X2=0 $Y2=0
cc_321 N_A_27_47#_c_257_n N_A_1011_47#_c_1076_n 0.0282006f $X=5.75 $Y=1.825
+ $X2=0 $Y2=0
cc_322 N_A_27_47#_c_258_n N_A_1011_47#_c_1076_n 0.00865498f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_323 N_A_27_47#_c_259_n N_A_1011_47#_c_1076_n 0.00430757f $X=5.895 $Y=1.825
+ $X2=0 $Y2=0
cc_324 N_A_27_47#_M1026_g N_A_1011_47#_c_1080_n 0.00165193f $X=4.98 $Y=0.415
+ $X2=0 $Y2=0
cc_325 N_A_27_47#_M1026_g N_A_1011_47#_c_1063_n 9.11618e-19 $X=4.98 $Y=0.415
+ $X2=0 $Y2=0
cc_326 N_A_27_47#_c_234_n N_A_1011_47#_c_1063_n 9.13335e-19 $X=5.415 $Y=1.32
+ $X2=0 $Y2=0
cc_327 N_A_27_47#_c_249_n N_A_1011_47#_c_1067_n 0.00172994f $X=5.515 $Y=1.99
+ $X2=0 $Y2=0
cc_328 N_A_27_47#_c_257_n N_A_1011_47#_c_1067_n 0.0251845f $X=5.75 $Y=1.825
+ $X2=0 $Y2=0
cc_329 N_A_27_47#_c_259_n N_A_1011_47#_c_1067_n 0.0026672f $X=5.895 $Y=1.825
+ $X2=0 $Y2=0
cc_330 N_A_27_47#_c_261_n N_A_1011_47#_c_1067_n 0.0197646f $X=7.13 $Y=1.825
+ $X2=0 $Y2=0
cc_331 N_A_27_47#_c_234_n N_A_1011_47#_c_1068_n 0.00253446f $X=5.415 $Y=1.32
+ $X2=0 $Y2=0
cc_332 N_A_27_47#_c_248_n N_A_1011_47#_c_1068_n 4.58049e-19 $X=5.515 $Y=1.575
+ $X2=0 $Y2=0
cc_333 N_A_27_47#_c_249_n N_A_1011_47#_c_1068_n 7.66691e-19 $X=5.515 $Y=1.99
+ $X2=0 $Y2=0
cc_334 N_A_27_47#_c_257_n N_A_1011_47#_c_1068_n 0.0135917f $X=5.75 $Y=1.825
+ $X2=0 $Y2=0
cc_335 N_A_27_47#_c_259_n N_A_1011_47#_c_1068_n 0.00215887f $X=5.895 $Y=1.825
+ $X2=0 $Y2=0
cc_336 N_A_27_47#_c_261_n N_A_1011_47#_c_1068_n 0.00517722f $X=7.13 $Y=1.825
+ $X2=0 $Y2=0
cc_337 N_A_27_47#_c_261_n N_A_1011_47#_c_1069_n 0.0168129f $X=7.13 $Y=1.825
+ $X2=0 $Y2=0
cc_338 N_A_27_47#_M1027_g N_A_1647_21#_M1008_g 0.0474153f $X=7.83 $Y=0.415 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_251_n N_A_1474_413#_c_1258_n 0.00640375f $X=7.28 $Y=1.99
+ $X2=0 $Y2=0
cc_340 N_A_27_47#_c_260_n N_A_1474_413#_c_1258_n 8.86193e-19 $X=7.325 $Y=1.825
+ $X2=0 $Y2=0
cc_341 N_A_27_47#_c_243_n N_A_1474_413#_c_1258_n 0.0115751f $X=7.315 $Y=1.41
+ $X2=0 $Y2=0
cc_342 N_A_27_47#_M1027_g N_A_1474_413#_c_1261_n 0.00862171f $X=7.83 $Y=0.415
+ $X2=0 $Y2=0
cc_343 N_A_27_47#_M1027_g N_A_1474_413#_c_1250_n 0.00427799f $X=7.83 $Y=0.415
+ $X2=0 $Y2=0
cc_344 N_A_27_47#_c_236_n N_A_1474_413#_c_1256_n 2.04942e-19 $X=7.755 $Y=1.32
+ $X2=0 $Y2=0
cc_345 N_A_27_47#_c_243_n N_A_1474_413#_c_1256_n 0.00153882f $X=7.315 $Y=1.41
+ $X2=0 $Y2=0
cc_346 N_A_27_47#_M1027_g N_A_1474_413#_c_1252_n 0.00124739f $X=7.83 $Y=0.415
+ $X2=0 $Y2=0
cc_347 N_A_27_47#_c_359_p N_VPWR_M1002_d 0.00171205f $X=0.78 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_348 N_A_27_47#_c_261_n N_VPWR_M1000_d 0.00710555f $X=7.13 $Y=1.825 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_245_n N_VPWR_c_1333_n 0.00955536f $X=0.97 $Y=1.74 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_253_n N_VPWR_c_1333_n 0.00629408f $X=0.665 $Y=1.88 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_359_p N_VPWR_c_1333_n 0.0135522f $X=0.78 $Y=1.795 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_255_n N_VPWR_c_1333_n 0.0246493f $X=0.265 $Y=1.96 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_256_n N_VPWR_c_1333_n 0.00146287f $X=0.895 $Y=1.825 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_c_258_n N_VPWR_c_1334_n 0.00142595f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_258_n N_VPWR_c_1335_n 8.00522e-19 $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_261_n N_VPWR_c_1336_n 0.00999501f $X=7.13 $Y=1.825 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_249_n N_VPWR_c_1341_n 0.00454633f $X=5.515 $Y=1.99 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_c_253_n N_VPWR_c_1345_n 0.00180073f $X=0.665 $Y=1.88 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_c_255_n N_VPWR_c_1345_n 0.0120313f $X=0.265 $Y=1.96 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_245_n N_VPWR_c_1346_n 0.00590576f $X=0.97 $Y=1.74 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_251_n N_VPWR_c_1347_n 0.00543513f $X=7.28 $Y=1.99 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_c_243_n N_VPWR_c_1347_n 2.64586e-19 $X=7.315 $Y=1.41 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_245_n N_VPWR_c_1332_n 0.00667006f $X=0.97 $Y=1.74 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_249_n N_VPWR_c_1332_n 0.00640619f $X=5.515 $Y=1.99 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_251_n N_VPWR_c_1332_n 0.00692642f $X=7.28 $Y=1.99 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_253_n N_VPWR_c_1332_n 0.00425497f $X=0.665 $Y=1.88 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_359_p N_VPWR_c_1332_n 5.98513e-19 $X=0.78 $Y=1.795 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_255_n N_VPWR_c_1332_n 0.00646745f $X=0.265 $Y=1.96 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_256_n N_VPWR_c_1332_n 0.32046f $X=0.895 $Y=1.825 $X2=0 $Y2=0
cc_370 N_A_27_47#_c_243_n N_VPWR_c_1332_n 6.79633e-19 $X=7.315 $Y=1.41 $X2=0
+ $Y2=0
cc_371 N_A_27_47#_c_258_n N_A_608_369#_c_1495_n 0.00670474f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_c_258_n N_A_608_369#_c_1491_n 0.0293627f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_258_n N_A_608_369#_c_1492_n 0.008435f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_374 N_A_27_47#_M1026_g N_A_608_369#_c_1487_n 0.0044467f $X=4.98 $Y=0.415
+ $X2=0 $Y2=0
cc_375 N_A_27_47#_M1026_g N_A_608_369#_c_1488_n 0.00914943f $X=4.98 $Y=0.415
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_c_258_n N_A_608_369#_c_1488_n 0.0104876f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_377 N_A_27_47#_M1026_g N_A_608_369#_c_1489_n 0.00199422f $X=4.98 $Y=0.415
+ $X2=0 $Y2=0
cc_378 N_A_27_47#_M1026_g N_A_608_369#_c_1490_n 0.00164257f $X=4.98 $Y=0.415
+ $X2=0 $Y2=0
cc_379 N_A_27_47#_c_257_n N_A_608_369#_c_1494_n 0.00293569f $X=5.75 $Y=1.825
+ $X2=0 $Y2=0
cc_380 N_A_27_47#_c_258_n N_A_608_369#_c_1494_n 0.011045f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_381 N_A_27_47#_c_258_n A_702_369# 0.00142862f $X=5.555 $Y=1.825 $X2=-0.19
+ $Y2=-0.24
cc_382 N_A_27_47#_c_238_n N_VGND_M1028_d 0.00215637f $X=0.665 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_383 N_A_27_47#_M1026_g N_VGND_c_1634_n 0.00339332f $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_M1007_g N_VGND_c_1638_n 0.00468308f $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_M1026_g N_VGND_c_1642_n 0.00431421f $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_c_451_p N_VGND_c_1646_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_c_238_n N_VGND_c_1646_n 0.00244629f $X=0.665 $Y=0.72 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_M1027_g N_VGND_c_1647_n 0.0037981f $X=7.83 $Y=0.415 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_M1028_s N_VGND_c_1649_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_M1007_g N_VGND_c_1649_n 0.00934478f $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_M1026_g N_VGND_c_1649_n 0.00732012f $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_M1027_g N_VGND_c_1649_n 0.005791f $X=7.83 $Y=0.415 $X2=0 $Y2=0
cc_393 N_A_27_47#_c_451_p N_VGND_c_1649_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_c_238_n N_VGND_c_1649_n 0.00602661f $X=0.665 $Y=0.72 $X2=0
+ $Y2=0
cc_395 N_A_27_47#_M1007_g N_VGND_c_1650_n 0.0101565f $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_c_238_n N_VGND_c_1650_n 0.0211078f $X=0.665 $Y=0.72 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_c_241_n N_VGND_c_1650_n 5.78916e-19 $X=0.97 $Y=1.235 $X2=0
+ $Y2=0
cc_398 N_SCE_M1013_g N_A_319_47#_M1021_g 0.0313276f $X=2.01 $Y=0.445 $X2=0 $Y2=0
cc_399 N_SCE_c_465_n N_A_319_47#_M1021_g 0.0112544f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_400 SCE N_A_319_47#_M1021_g 0.00326341f $X=2.07 $Y=0.84 $X2=0 $Y2=0
cc_401 N_SCE_c_466_n N_A_319_47#_c_565_n 2.11997e-19 $X=3.42 $Y=0.95 $X2=0 $Y2=0
cc_402 N_SCE_c_467_n N_A_319_47#_c_565_n 0.0157262f $X=3.53 $Y=0.95 $X2=0 $Y2=0
cc_403 N_SCE_c_470_n N_A_319_47#_c_560_n 0.00268171f $X=1.96 $Y=1.77 $X2=0 $Y2=0
cc_404 N_SCE_M1013_g N_A_319_47#_c_560_n 0.00837412f $X=2.01 $Y=0.445 $X2=0
+ $Y2=0
cc_405 N_SCE_c_473_n N_A_319_47#_c_560_n 0.0103947f $X=2.025 $Y=1.52 $X2=0 $Y2=0
cc_406 N_SCE_c_468_n N_A_319_47#_c_560_n 0.0117596f $X=2.047 $Y=0.785 $X2=0
+ $Y2=0
cc_407 SCE N_A_319_47#_c_560_n 0.0675595f $X=2.07 $Y=0.84 $X2=0 $Y2=0
cc_408 N_SCE_c_470_n N_A_319_47#_c_567_n 0.00579439f $X=1.96 $Y=1.77 $X2=0 $Y2=0
cc_409 N_SCE_c_470_n N_A_319_47#_c_573_n 0.0137048f $X=1.96 $Y=1.77 $X2=0 $Y2=0
cc_410 N_SCE_c_472_n N_A_319_47#_c_573_n 0.00528858f $X=2.43 $Y=1.77 $X2=0 $Y2=0
cc_411 N_SCE_c_473_n N_A_319_47#_c_573_n 0.0048728f $X=2.025 $Y=1.52 $X2=0 $Y2=0
cc_412 SCE N_A_319_47#_c_573_n 0.0212535f $X=2.07 $Y=0.84 $X2=0 $Y2=0
cc_413 N_SCE_c_470_n N_A_319_47#_c_561_n 6.74057e-19 $X=1.96 $Y=1.77 $X2=0 $Y2=0
cc_414 N_SCE_M1013_g N_A_319_47#_c_561_n 0.00113389f $X=2.01 $Y=0.445 $X2=0
+ $Y2=0
cc_415 N_SCE_c_472_n N_A_319_47#_c_561_n 0.00301815f $X=2.43 $Y=1.77 $X2=0 $Y2=0
cc_416 N_SCE_c_473_n N_A_319_47#_c_561_n 0.0108646f $X=2.025 $Y=1.52 $X2=0 $Y2=0
cc_417 SCE N_A_319_47#_c_561_n 0.0429654f $X=2.07 $Y=0.84 $X2=0 $Y2=0
cc_418 N_SCE_c_466_n N_A_319_47#_c_569_n 0.00960462f $X=3.42 $Y=0.95 $X2=0 $Y2=0
cc_419 N_SCE_c_467_n N_A_319_47#_c_569_n 5.10023e-19 $X=3.53 $Y=0.95 $X2=0 $Y2=0
cc_420 N_SCE_c_465_n N_A_319_47#_c_563_n 0.0198926f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_421 N_SCE_c_466_n N_A_319_47#_c_563_n 0.00387695f $X=3.42 $Y=0.95 $X2=0 $Y2=0
cc_422 SCE N_A_319_47#_c_563_n 0.0133765f $X=2.07 $Y=0.84 $X2=0 $Y2=0
cc_423 N_SCE_c_465_n N_A_319_47#_c_564_n 0.00342266f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_424 N_SCE_c_473_n N_A_319_47#_c_564_n 0.0053677f $X=2.025 $Y=1.52 $X2=0 $Y2=0
cc_425 SCE N_A_319_47#_c_564_n 9.65653e-19 $X=2.07 $Y=0.84 $X2=0 $Y2=0
cc_426 N_SCE_c_472_n N_A_319_47#_c_580_n 0.0087726f $X=2.43 $Y=1.77 $X2=0 $Y2=0
cc_427 N_SCE_c_472_n N_D_c_675_n 0.0317564f $X=2.43 $Y=1.77 $X2=-0.19 $Y2=-0.24
cc_428 N_SCE_c_465_n N_D_c_675_n 6.57582e-19 $X=3.335 $Y=0.7 $X2=-0.19 $Y2=-0.24
cc_429 N_SCE_c_473_n N_D_c_675_n 0.0163209f $X=2.025 $Y=1.52 $X2=-0.19 $Y2=-0.24
cc_430 N_SCE_M1029_g N_D_M1003_g 0.0117556f $X=3.53 $Y=0.445 $X2=0 $Y2=0
cc_431 N_SCE_c_465_n N_D_M1003_g 0.0135073f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_432 N_SCE_c_466_n N_D_M1003_g 0.00203037f $X=3.42 $Y=0.95 $X2=0 $Y2=0
cc_433 N_SCE_c_467_n N_D_M1003_g 0.0215793f $X=3.53 $Y=0.95 $X2=0 $Y2=0
cc_434 N_SCE_c_465_n D 0.00670682f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_435 N_SCE_c_473_n D 2.13317e-19 $X=2.025 $Y=1.52 $X2=0 $Y2=0
cc_436 N_SCE_M1029_g N_SCD_M1020_g 0.0574661f $X=3.53 $Y=0.445 $X2=0 $Y2=0
cc_437 N_SCE_c_466_n N_SCD_M1020_g 0.00124626f $X=3.42 $Y=0.95 $X2=0 $Y2=0
cc_438 N_SCE_c_466_n SCD 0.00503288f $X=3.42 $Y=0.95 $X2=0 $Y2=0
cc_439 N_SCE_c_467_n SCD 5.8751e-19 $X=3.53 $Y=0.95 $X2=0 $Y2=0
cc_440 N_SCE_M1029_g N_A_203_47#_c_771_n 0.00105565f $X=3.53 $Y=0.445 $X2=0
+ $Y2=0
cc_441 N_SCE_c_465_n N_A_203_47#_c_771_n 0.0429067f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_442 N_SCE_c_466_n N_A_203_47#_c_771_n 0.0110804f $X=3.42 $Y=0.95 $X2=0 $Y2=0
cc_443 N_SCE_c_473_n N_A_203_47#_c_771_n 0.0035596f $X=2.025 $Y=1.52 $X2=0 $Y2=0
cc_444 N_SCE_c_467_n N_A_203_47#_c_771_n 0.00506552f $X=3.53 $Y=0.95 $X2=0 $Y2=0
cc_445 N_SCE_c_468_n N_A_203_47#_c_771_n 0.00666037f $X=2.047 $Y=0.785 $X2=0
+ $Y2=0
cc_446 SCE N_A_203_47#_c_771_n 0.0242551f $X=2.07 $Y=0.84 $X2=0 $Y2=0
cc_447 N_SCE_c_470_n N_A_203_47#_c_780_n 0.00143269f $X=1.96 $Y=1.77 $X2=0 $Y2=0
cc_448 N_SCE_c_470_n N_VPWR_c_1334_n 0.0113766f $X=1.96 $Y=1.77 $X2=0 $Y2=0
cc_449 N_SCE_c_472_n N_VPWR_c_1334_n 0.00947361f $X=2.43 $Y=1.77 $X2=0 $Y2=0
cc_450 N_SCE_c_472_n N_VPWR_c_1339_n 0.00454152f $X=2.43 $Y=1.77 $X2=0 $Y2=0
cc_451 N_SCE_c_470_n N_VPWR_c_1346_n 0.00312096f $X=1.96 $Y=1.77 $X2=0 $Y2=0
cc_452 N_SCE_c_470_n N_VPWR_c_1332_n 0.00489637f $X=1.96 $Y=1.77 $X2=0 $Y2=0
cc_453 N_SCE_c_472_n N_VPWR_c_1332_n 0.00504866f $X=2.43 $Y=1.77 $X2=0 $Y2=0
cc_454 N_SCE_c_465_n N_A_608_369#_M1003_d 0.00271541f $X=3.335 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_455 N_SCE_c_472_n N_A_608_369#_c_1495_n 6.17318e-19 $X=2.43 $Y=1.77 $X2=0
+ $Y2=0
cc_456 N_SCE_M1029_g N_A_608_369#_c_1507_n 0.00787009f $X=3.53 $Y=0.445 $X2=0
+ $Y2=0
cc_457 N_SCE_c_465_n N_A_608_369#_c_1507_n 0.0209567f $X=3.335 $Y=0.7 $X2=0
+ $Y2=0
cc_458 N_SCE_c_467_n N_A_608_369#_c_1507_n 4.66881e-19 $X=3.53 $Y=0.95 $X2=0
+ $Y2=0
cc_459 N_SCE_M1029_g N_A_608_369#_c_1484_n 0.00410769f $X=3.53 $Y=0.445 $X2=0
+ $Y2=0
cc_460 N_SCE_c_465_n N_A_608_369#_c_1484_n 0.00517226f $X=3.335 $Y=0.7 $X2=0
+ $Y2=0
cc_461 N_SCE_M1029_g N_A_608_369#_c_1486_n 0.00111248f $X=3.53 $Y=0.445 $X2=0
+ $Y2=0
cc_462 N_SCE_c_465_n N_A_608_369#_c_1486_n 0.00650856f $X=3.335 $Y=0.7 $X2=0
+ $Y2=0
cc_463 N_SCE_c_466_n N_A_608_369#_c_1486_n 0.00423271f $X=3.42 $Y=0.95 $X2=0
+ $Y2=0
cc_464 N_SCE_c_465_n N_VGND_M1013_d 0.00114095f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_465 N_SCE_c_468_n N_VGND_M1013_d 7.7409e-19 $X=2.047 $Y=0.785 $X2=0 $Y2=0
cc_466 N_SCE_M1013_g N_VGND_c_1633_n 0.00775013f $X=2.01 $Y=0.445 $X2=0 $Y2=0
cc_467 N_SCE_c_465_n N_VGND_c_1633_n 0.00915315f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_468 N_SCE_c_468_n N_VGND_c_1633_n 0.0063553f $X=2.047 $Y=0.785 $X2=0 $Y2=0
cc_469 N_SCE_M1013_g N_VGND_c_1638_n 0.00393143f $X=2.01 $Y=0.445 $X2=0 $Y2=0
cc_470 N_SCE_c_468_n N_VGND_c_1638_n 0.00293412f $X=2.047 $Y=0.785 $X2=0 $Y2=0
cc_471 N_SCE_M1029_g N_VGND_c_1640_n 0.00362032f $X=3.53 $Y=0.445 $X2=0 $Y2=0
cc_472 N_SCE_c_465_n N_VGND_c_1640_n 0.0109339f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_473 N_SCE_M1013_g N_VGND_c_1649_n 0.00556035f $X=2.01 $Y=0.445 $X2=0 $Y2=0
cc_474 N_SCE_M1029_g N_VGND_c_1649_n 0.00537207f $X=3.53 $Y=0.445 $X2=0 $Y2=0
cc_475 N_SCE_c_465_n N_VGND_c_1649_n 0.00875593f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_476 N_SCE_c_468_n N_VGND_c_1649_n 0.00263734f $X=2.047 $Y=0.785 $X2=0 $Y2=0
cc_477 N_SCE_c_465_n A_507_47# 0.00476634f $X=3.335 $Y=0.7 $X2=-0.19 $Y2=-0.24
cc_478 N_A_319_47#_c_565_n N_D_c_675_n 0.0267545f $X=3.42 $Y=1.77 $X2=-0.19
+ $Y2=-0.24
cc_479 N_A_319_47#_c_561_n N_D_c_675_n 0.00380365f $X=2.47 $Y=1.86 $X2=-0.19
+ $Y2=-0.24
cc_480 N_A_319_47#_c_575_n N_D_c_675_n 0.0166353f $X=3.33 $Y=1.967 $X2=-0.19
+ $Y2=-0.24
cc_481 N_A_319_47#_c_569_n N_D_c_675_n 0.00129025f $X=3.455 $Y=1.52 $X2=-0.19
+ $Y2=-0.24
cc_482 N_A_319_47#_M1021_g N_D_M1003_g 0.0248729f $X=2.46 $Y=0.445 $X2=0 $Y2=0
cc_483 N_A_319_47#_c_565_n N_D_M1003_g 0.0166724f $X=3.42 $Y=1.77 $X2=0 $Y2=0
cc_484 N_A_319_47#_c_561_n N_D_M1003_g 0.00537883f $X=2.47 $Y=1.86 $X2=0 $Y2=0
cc_485 N_A_319_47#_c_569_n N_D_M1003_g 3.57045e-19 $X=3.455 $Y=1.52 $X2=0 $Y2=0
cc_486 N_A_319_47#_c_563_n N_D_M1003_g 6.95674e-19 $X=2.55 $Y=1.04 $X2=0 $Y2=0
cc_487 N_A_319_47#_c_564_n N_D_M1003_g 0.0189419f $X=2.55 $Y=1.04 $X2=0 $Y2=0
cc_488 N_A_319_47#_c_565_n D 0.00203711f $X=3.42 $Y=1.77 $X2=0 $Y2=0
cc_489 N_A_319_47#_c_561_n D 0.0232562f $X=2.47 $Y=1.86 $X2=0 $Y2=0
cc_490 N_A_319_47#_c_575_n D 0.0232233f $X=3.33 $Y=1.967 $X2=0 $Y2=0
cc_491 N_A_319_47#_c_569_n D 0.0246039f $X=3.455 $Y=1.52 $X2=0 $Y2=0
cc_492 N_A_319_47#_c_565_n N_SCD_c_718_n 0.0337327f $X=3.42 $Y=1.77 $X2=0 $Y2=0
cc_493 N_A_319_47#_c_575_n N_SCD_c_718_n 2.15603e-19 $X=3.33 $Y=1.967 $X2=0
+ $Y2=0
cc_494 N_A_319_47#_c_569_n N_SCD_c_718_n 0.0025761f $X=3.455 $Y=1.52 $X2=0 $Y2=0
cc_495 N_A_319_47#_c_565_n SCD 0.00200159f $X=3.42 $Y=1.77 $X2=0 $Y2=0
cc_496 N_A_319_47#_c_569_n SCD 0.021781f $X=3.455 $Y=1.52 $X2=0 $Y2=0
cc_497 N_A_319_47#_c_565_n N_SCD_c_716_n 0.0166742f $X=3.42 $Y=1.77 $X2=0 $Y2=0
cc_498 N_A_319_47#_c_569_n N_SCD_c_716_n 2.90907e-19 $X=3.455 $Y=1.52 $X2=0
+ $Y2=0
cc_499 N_A_319_47#_c_560_n N_A_203_47#_c_770_n 0.00266292f $X=1.62 $Y=1.86 $X2=0
+ $Y2=0
cc_500 N_A_319_47#_M1021_g N_A_203_47#_c_771_n 0.0013306f $X=2.46 $Y=0.445 $X2=0
+ $Y2=0
cc_501 N_A_319_47#_c_565_n N_A_203_47#_c_771_n 2.76438e-19 $X=3.42 $Y=1.77 $X2=0
+ $Y2=0
cc_502 N_A_319_47#_c_560_n N_A_203_47#_c_771_n 0.0181188f $X=1.62 $Y=1.86 $X2=0
+ $Y2=0
cc_503 N_A_319_47#_c_569_n N_A_203_47#_c_771_n 0.00222993f $X=3.455 $Y=1.52
+ $X2=0 $Y2=0
cc_504 N_A_319_47#_c_562_n N_A_203_47#_c_771_n 0.0047194f $X=1.74 $Y=0.36 $X2=0
+ $Y2=0
cc_505 N_A_319_47#_c_563_n N_A_203_47#_c_771_n 0.00829416f $X=2.55 $Y=1.04 $X2=0
+ $Y2=0
cc_506 N_A_319_47#_c_564_n N_A_203_47#_c_771_n 0.00516347f $X=2.55 $Y=1.04 $X2=0
+ $Y2=0
cc_507 N_A_319_47#_c_560_n N_A_203_47#_c_780_n 0.0981158f $X=1.62 $Y=1.86 $X2=0
+ $Y2=0
cc_508 N_A_319_47#_c_567_n N_A_203_47#_c_780_n 0.0273077f $X=1.725 $Y=2.175
+ $X2=0 $Y2=0
cc_509 N_A_319_47#_c_562_n N_A_203_47#_c_780_n 0.00751792f $X=1.74 $Y=0.36 $X2=0
+ $Y2=0
cc_510 N_A_319_47#_c_570_n N_A_203_47#_c_780_n 0.0159784f $X=1.672 $Y=1.967
+ $X2=0 $Y2=0
cc_511 N_A_319_47#_c_573_n N_VPWR_M1009_d 0.00351251f $X=2.385 $Y=1.967 $X2=0
+ $Y2=0
cc_512 N_A_319_47#_c_567_n N_VPWR_c_1334_n 0.0154733f $X=1.725 $Y=2.175 $X2=0
+ $Y2=0
cc_513 N_A_319_47#_c_573_n N_VPWR_c_1334_n 0.0184987f $X=2.385 $Y=1.967 $X2=0
+ $Y2=0
cc_514 N_A_319_47#_c_565_n N_VPWR_c_1339_n 0.00441747f $X=3.42 $Y=1.77 $X2=0
+ $Y2=0
cc_515 N_A_319_47#_c_573_n N_VPWR_c_1339_n 3.89445e-19 $X=2.385 $Y=1.967 $X2=0
+ $Y2=0
cc_516 N_A_319_47#_c_575_n N_VPWR_c_1339_n 0.00525224f $X=3.33 $Y=1.967 $X2=0
+ $Y2=0
cc_517 N_A_319_47#_c_580_n N_VPWR_c_1339_n 0.00269709f $X=2.47 $Y=1.967 $X2=0
+ $Y2=0
cc_518 N_A_319_47#_c_567_n N_VPWR_c_1346_n 0.0170259f $X=1.725 $Y=2.175 $X2=0
+ $Y2=0
cc_519 N_A_319_47#_c_573_n N_VPWR_c_1346_n 0.00234063f $X=2.385 $Y=1.967 $X2=0
+ $Y2=0
cc_520 N_A_319_47#_M1009_s N_VPWR_c_1332_n 0.0019314f $X=1.6 $Y=1.845 $X2=0
+ $Y2=0
cc_521 N_A_319_47#_c_565_n N_VPWR_c_1332_n 0.00617905f $X=3.42 $Y=1.77 $X2=0
+ $Y2=0
cc_522 N_A_319_47#_c_567_n N_VPWR_c_1332_n 0.00494372f $X=1.725 $Y=2.175 $X2=0
+ $Y2=0
cc_523 N_A_319_47#_c_573_n N_VPWR_c_1332_n 0.00311756f $X=2.385 $Y=1.967 $X2=0
+ $Y2=0
cc_524 N_A_319_47#_c_575_n N_VPWR_c_1332_n 0.00494869f $X=3.33 $Y=1.967 $X2=0
+ $Y2=0
cc_525 N_A_319_47#_c_580_n N_VPWR_c_1332_n 0.0020288f $X=2.47 $Y=1.967 $X2=0
+ $Y2=0
cc_526 N_A_319_47#_c_575_n A_504_369# 0.00716796f $X=3.33 $Y=1.967 $X2=-0.19
+ $Y2=-0.24
cc_527 N_A_319_47#_c_575_n N_A_608_369#_M1030_d 0.00417681f $X=3.33 $Y=1.967
+ $X2=0 $Y2=0
cc_528 N_A_319_47#_c_565_n N_A_608_369#_c_1495_n 0.0103902f $X=3.42 $Y=1.77
+ $X2=0 $Y2=0
cc_529 N_A_319_47#_c_575_n N_A_608_369#_c_1495_n 0.0324509f $X=3.33 $Y=1.967
+ $X2=0 $Y2=0
cc_530 N_A_319_47#_M1021_g N_A_608_369#_c_1507_n 5.06401e-19 $X=2.46 $Y=0.445
+ $X2=0 $Y2=0
cc_531 N_A_319_47#_c_565_n N_A_608_369#_c_1519_n 0.00369522f $X=3.42 $Y=1.77
+ $X2=0 $Y2=0
cc_532 N_A_319_47#_c_565_n N_A_608_369#_c_1492_n 5.55331e-19 $X=3.42 $Y=1.77
+ $X2=0 $Y2=0
cc_533 N_A_319_47#_c_575_n N_A_608_369#_c_1492_n 0.00647567f $X=3.33 $Y=1.967
+ $X2=0 $Y2=0
cc_534 N_A_319_47#_c_569_n N_A_608_369#_c_1492_n 0.00209567f $X=3.455 $Y=1.52
+ $X2=0 $Y2=0
cc_535 N_A_319_47#_M1021_g N_VGND_c_1633_n 0.00907666f $X=2.46 $Y=0.445 $X2=0
+ $Y2=0
cc_536 N_A_319_47#_c_562_n N_VGND_c_1638_n 0.0202133f $X=1.74 $Y=0.36 $X2=0
+ $Y2=0
cc_537 N_A_319_47#_M1021_g N_VGND_c_1640_n 0.00365142f $X=2.46 $Y=0.445 $X2=0
+ $Y2=0
cc_538 N_A_319_47#_M1013_s N_VGND_c_1649_n 0.00233134f $X=1.595 $Y=0.235 $X2=0
+ $Y2=0
cc_539 N_A_319_47#_M1021_g N_VGND_c_1649_n 0.00431635f $X=2.46 $Y=0.445 $X2=0
+ $Y2=0
cc_540 N_A_319_47#_c_562_n N_VGND_c_1649_n 0.00622938f $X=1.74 $Y=0.36 $X2=0
+ $Y2=0
cc_541 N_A_319_47#_c_562_n N_VGND_c_1650_n 0.00203921f $X=1.74 $Y=0.36 $X2=0
+ $Y2=0
cc_542 N_D_M1003_g SCD 0.00550319f $X=3 $Y=0.445 $X2=0 $Y2=0
cc_543 N_D_M1003_g N_A_203_47#_c_771_n 0.00372001f $X=3 $Y=0.445 $X2=0 $Y2=0
cc_544 D N_A_203_47#_c_771_n 0.00878071f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_545 N_D_c_675_n N_VPWR_c_1334_n 0.00170479f $X=2.95 $Y=1.77 $X2=0 $Y2=0
cc_546 N_D_c_675_n N_VPWR_c_1339_n 0.00455384f $X=2.95 $Y=1.77 $X2=0 $Y2=0
cc_547 N_D_c_675_n N_VPWR_c_1332_n 0.00628186f $X=2.95 $Y=1.77 $X2=0 $Y2=0
cc_548 N_D_c_675_n N_A_608_369#_c_1495_n 0.00796293f $X=2.95 $Y=1.77 $X2=0 $Y2=0
cc_549 N_D_M1003_g N_A_608_369#_c_1507_n 0.0031616f $X=3 $Y=0.445 $X2=0 $Y2=0
cc_550 N_D_M1003_g N_VGND_c_1633_n 0.0015803f $X=3 $Y=0.445 $X2=0 $Y2=0
cc_551 N_D_M1003_g N_VGND_c_1640_n 0.0042011f $X=3 $Y=0.445 $X2=0 $Y2=0
cc_552 N_D_M1003_g N_VGND_c_1649_n 0.00607125f $X=3 $Y=0.445 $X2=0 $Y2=0
cc_553 N_SCD_M1020_g N_A_203_47#_c_771_n 0.00245337f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_554 SCD N_A_203_47#_c_771_n 0.00958434f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_555 N_SCD_c_716_n N_A_203_47#_c_771_n 0.00138804f $X=3.97 $Y=1.355 $X2=0
+ $Y2=0
cc_556 N_SCD_c_718_n N_VPWR_c_1335_n 0.00627598f $X=3.935 $Y=1.77 $X2=0 $Y2=0
cc_557 N_SCD_c_718_n N_VPWR_c_1339_n 0.00504444f $X=3.935 $Y=1.77 $X2=0 $Y2=0
cc_558 N_SCD_c_718_n N_VPWR_c_1332_n 0.00784388f $X=3.935 $Y=1.77 $X2=0 $Y2=0
cc_559 N_SCD_c_718_n N_A_608_369#_c_1495_n 0.00520197f $X=3.935 $Y=1.77 $X2=0
+ $Y2=0
cc_560 N_SCD_M1020_g N_A_608_369#_c_1507_n 0.00468836f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_561 N_SCD_c_718_n N_A_608_369#_c_1519_n 0.0072605f $X=3.935 $Y=1.77 $X2=0
+ $Y2=0
cc_562 N_SCD_M1020_g N_A_608_369#_c_1484_n 0.00659485f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_563 N_SCD_c_718_n N_A_608_369#_c_1491_n 0.0108115f $X=3.935 $Y=1.77 $X2=0
+ $Y2=0
cc_564 SCD N_A_608_369#_c_1491_n 0.0138435f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_565 N_SCD_c_716_n N_A_608_369#_c_1491_n 0.00199327f $X=3.97 $Y=1.355 $X2=0
+ $Y2=0
cc_566 N_SCD_c_718_n N_A_608_369#_c_1492_n 0.00271587f $X=3.935 $Y=1.77 $X2=0
+ $Y2=0
cc_567 SCD N_A_608_369#_c_1492_n 0.0118154f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_568 N_SCD_M1020_g N_A_608_369#_c_1485_n 0.00830957f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_569 SCD N_A_608_369#_c_1485_n 0.0137228f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_570 N_SCD_c_716_n N_A_608_369#_c_1485_n 0.00215057f $X=3.97 $Y=1.355 $X2=0
+ $Y2=0
cc_571 N_SCD_M1020_g N_A_608_369#_c_1486_n 0.00228168f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_572 SCD N_A_608_369#_c_1486_n 0.0120393f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_573 N_SCD_M1020_g N_A_608_369#_c_1487_n 0.00233059f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_574 N_SCD_M1020_g N_A_608_369#_c_1488_n 0.00400866f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_575 N_SCD_c_717_n N_A_608_369#_c_1488_n 0.00345986f $X=3.935 $Y=1.67 $X2=0
+ $Y2=0
cc_576 N_SCD_c_718_n N_A_608_369#_c_1488_n 0.00105043f $X=3.935 $Y=1.77 $X2=0
+ $Y2=0
cc_577 SCD N_A_608_369#_c_1488_n 0.0231455f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_578 N_SCD_c_716_n N_A_608_369#_c_1488_n 0.00629503f $X=3.97 $Y=1.355 $X2=0
+ $Y2=0
cc_579 N_SCD_M1020_g N_A_608_369#_c_1489_n 4.17422e-19 $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_580 N_SCD_c_718_n N_A_608_369#_c_1494_n 0.00289044f $X=3.935 $Y=1.77 $X2=0
+ $Y2=0
cc_581 N_SCD_M1020_g N_VGND_c_1634_n 0.0104318f $X=3.91 $Y=0.445 $X2=0 $Y2=0
cc_582 N_SCD_M1020_g N_VGND_c_1640_n 0.00404961f $X=3.91 $Y=0.445 $X2=0 $Y2=0
cc_583 N_SCD_M1020_g N_VGND_c_1649_n 0.00679524f $X=3.91 $Y=0.445 $X2=0 $Y2=0
cc_584 N_A_203_47#_c_774_n N_A_1189_21#_M1012_d 2.26277e-19 $X=7.23 $Y=0.805
+ $X2=-0.19 $Y2=-0.24
cc_585 N_A_203_47#_c_774_n N_A_1189_21#_M1005_g 0.00175918f $X=7.23 $Y=0.805
+ $X2=0 $Y2=0
cc_586 N_A_203_47#_c_777_n N_A_1189_21#_M1005_g 0.0145234f $X=5.45 $Y=0.705
+ $X2=0 $Y2=0
cc_587 N_A_203_47#_c_774_n N_A_1189_21#_c_970_n 0.0370465f $X=7.23 $Y=0.805
+ $X2=0 $Y2=0
cc_588 N_A_203_47#_c_774_n N_A_1189_21#_c_971_n 0.00214522f $X=7.23 $Y=0.805
+ $X2=0 $Y2=0
cc_589 N_A_203_47#_c_775_n N_A_1189_21#_c_971_n 0.0145234f $X=5.45 $Y=0.87 $X2=0
+ $Y2=0
cc_590 N_A_203_47#_c_769_n N_A_1189_21#_c_998_n 0.00335557f $X=7.735 $Y=0.87
+ $X2=0 $Y2=0
cc_591 N_A_203_47#_c_773_n N_A_1189_21#_c_998_n 0.00225381f $X=7.395 $Y=0.805
+ $X2=0 $Y2=0
cc_592 N_A_203_47#_c_779_n N_A_1189_21#_c_998_n 0.00420064f $X=7.365 $Y=0.705
+ $X2=0 $Y2=0
cc_593 N_A_203_47#_c_768_n N_A_1189_21#_c_972_n 0.00442548f $X=7.825 $Y=1.74
+ $X2=0 $Y2=0
cc_594 N_A_203_47#_c_769_n N_A_1189_21#_c_1002_n 5.99165e-19 $X=7.735 $Y=0.87
+ $X2=0 $Y2=0
cc_595 N_A_203_47#_c_773_n N_A_1189_21#_c_1002_n 5.90931e-19 $X=7.395 $Y=0.805
+ $X2=0 $Y2=0
cc_596 N_A_203_47#_c_774_n N_A_1189_21#_c_1002_n 0.00516952f $X=7.23 $Y=0.805
+ $X2=0 $Y2=0
cc_597 N_A_203_47#_c_779_n N_A_1189_21#_c_1002_n 0.00267868f $X=7.365 $Y=0.705
+ $X2=0 $Y2=0
cc_598 N_A_203_47#_c_768_n N_A_1189_21#_c_973_n 0.00194004f $X=7.825 $Y=1.74
+ $X2=0 $Y2=0
cc_599 N_A_203_47#_c_769_n N_A_1189_21#_c_973_n 0.0189118f $X=7.735 $Y=0.87
+ $X2=0 $Y2=0
cc_600 N_A_203_47#_c_773_n N_A_1189_21#_c_973_n 3.95623e-19 $X=7.395 $Y=0.805
+ $X2=0 $Y2=0
cc_601 N_A_203_47#_c_774_n N_A_1189_21#_c_973_n 0.0258444f $X=7.23 $Y=0.805
+ $X2=0 $Y2=0
cc_602 N_A_203_47#_c_778_n N_A_1189_21#_c_973_n 0.00195749f $X=7.365 $Y=0.87
+ $X2=0 $Y2=0
cc_603 N_A_203_47#_c_769_n N_A_1011_47#_M1012_g 3.9777e-19 $X=7.735 $Y=0.87
+ $X2=0 $Y2=0
cc_604 N_A_203_47#_c_779_n N_A_1011_47#_M1012_g 0.0233325f $X=7.365 $Y=0.705
+ $X2=0 $Y2=0
cc_605 N_A_203_47#_c_781_n N_A_1011_47#_c_1076_n 0.00454283f $X=5 $Y=1.99 $X2=0
+ $Y2=0
cc_606 N_A_203_47#_c_767_n N_A_1011_47#_c_1076_n 0.00454699f $X=4.99 $Y=1.74
+ $X2=0 $Y2=0
cc_607 N_A_203_47#_c_772_n N_A_1011_47#_c_1080_n 0.0026338f $X=5.385 $Y=0.805
+ $X2=0 $Y2=0
cc_608 N_A_203_47#_c_774_n N_A_1011_47#_c_1080_n 0.00505066f $X=7.23 $Y=0.805
+ $X2=0 $Y2=0
cc_609 N_A_203_47#_c_775_n N_A_1011_47#_c_1080_n 0.00218731f $X=5.45 $Y=0.87
+ $X2=0 $Y2=0
cc_610 N_A_203_47#_c_776_n N_A_1011_47#_c_1080_n 0.0238697f $X=5.45 $Y=0.87
+ $X2=0 $Y2=0
cc_611 N_A_203_47#_c_777_n N_A_1011_47#_c_1080_n 0.00847732f $X=5.45 $Y=0.705
+ $X2=0 $Y2=0
cc_612 N_A_203_47#_c_767_n N_A_1011_47#_c_1063_n 0.00995592f $X=4.99 $Y=1.74
+ $X2=0 $Y2=0
cc_613 N_A_203_47#_c_772_n N_A_1011_47#_c_1063_n 0.00104696f $X=5.385 $Y=0.805
+ $X2=0 $Y2=0
cc_614 N_A_203_47#_c_774_n N_A_1011_47#_c_1063_n 0.0188221f $X=7.23 $Y=0.805
+ $X2=0 $Y2=0
cc_615 N_A_203_47#_c_776_n N_A_1011_47#_c_1063_n 0.0241643f $X=5.45 $Y=0.87
+ $X2=0 $Y2=0
cc_616 N_A_203_47#_c_777_n N_A_1011_47#_c_1063_n 0.00620262f $X=5.45 $Y=0.705
+ $X2=0 $Y2=0
cc_617 N_A_203_47#_c_767_n N_A_1011_47#_c_1068_n 0.00657117f $X=4.99 $Y=1.74
+ $X2=0 $Y2=0
cc_618 N_A_203_47#_c_774_n N_A_1011_47#_c_1068_n 0.0065601f $X=7.23 $Y=0.805
+ $X2=0 $Y2=0
cc_619 N_A_203_47#_c_774_n N_A_1011_47#_c_1069_n 0.00229853f $X=7.23 $Y=0.805
+ $X2=0 $Y2=0
cc_620 N_A_203_47#_c_768_n N_A_1647_21#_M1008_g 0.00204049f $X=7.825 $Y=1.74
+ $X2=0 $Y2=0
cc_621 N_A_203_47#_c_769_n N_A_1647_21#_M1008_g 0.0010356f $X=7.735 $Y=0.87
+ $X2=0 $Y2=0
cc_622 N_A_203_47#_c_782_n N_A_1647_21#_c_1170_n 0.0359061f $X=7.76 $Y=1.99
+ $X2=0 $Y2=0
cc_623 N_A_203_47#_c_768_n N_A_1647_21#_c_1170_n 3.34486e-19 $X=7.825 $Y=1.74
+ $X2=0 $Y2=0
cc_624 N_A_203_47#_c_782_n N_A_1474_413#_c_1258_n 0.014497f $X=7.76 $Y=1.99
+ $X2=0 $Y2=0
cc_625 N_A_203_47#_c_768_n N_A_1474_413#_c_1258_n 0.00940433f $X=7.825 $Y=1.74
+ $X2=0 $Y2=0
cc_626 N_A_203_47#_c_769_n N_A_1474_413#_c_1261_n 0.0320299f $X=7.735 $Y=0.87
+ $X2=0 $Y2=0
cc_627 N_A_203_47#_c_773_n N_A_1474_413#_c_1261_n 8.95493e-19 $X=7.395 $Y=0.805
+ $X2=0 $Y2=0
cc_628 N_A_203_47#_c_778_n N_A_1474_413#_c_1261_n 7.65858e-19 $X=7.365 $Y=0.87
+ $X2=0 $Y2=0
cc_629 N_A_203_47#_c_779_n N_A_1474_413#_c_1261_n 0.0015773f $X=7.365 $Y=0.705
+ $X2=0 $Y2=0
cc_630 N_A_203_47#_c_769_n N_A_1474_413#_c_1250_n 0.0240657f $X=7.735 $Y=0.87
+ $X2=0 $Y2=0
cc_631 N_A_203_47#_c_773_n N_A_1474_413#_c_1250_n 0.00122719f $X=7.395 $Y=0.805
+ $X2=0 $Y2=0
cc_632 N_A_203_47#_c_782_n N_A_1474_413#_c_1256_n 0.006274f $X=7.76 $Y=1.99
+ $X2=0 $Y2=0
cc_633 N_A_203_47#_c_768_n N_A_1474_413#_c_1256_n 0.043296f $X=7.825 $Y=1.74
+ $X2=0 $Y2=0
cc_634 N_A_203_47#_c_768_n N_A_1474_413#_c_1252_n 0.024806f $X=7.825 $Y=1.74
+ $X2=0 $Y2=0
cc_635 N_A_203_47#_c_769_n N_A_1474_413#_c_1252_n 0.003753f $X=7.735 $Y=0.87
+ $X2=0 $Y2=0
cc_636 N_A_203_47#_c_780_n N_VPWR_c_1333_n 0.0107869f $X=1.2 $Y=0.51 $X2=0 $Y2=0
cc_637 N_A_203_47#_c_780_n N_VPWR_c_1334_n 5.70469e-19 $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_638 N_A_203_47#_c_781_n N_VPWR_c_1335_n 0.00261116f $X=5 $Y=1.99 $X2=0 $Y2=0
cc_639 N_A_203_47#_c_781_n N_VPWR_c_1341_n 0.00659238f $X=5 $Y=1.99 $X2=0 $Y2=0
cc_640 N_A_203_47#_c_780_n N_VPWR_c_1346_n 0.0163465f $X=1.2 $Y=0.51 $X2=0 $Y2=0
cc_641 N_A_203_47#_c_782_n N_VPWR_c_1347_n 0.00460277f $X=7.76 $Y=1.99 $X2=0
+ $Y2=0
cc_642 N_A_203_47#_c_781_n N_VPWR_c_1332_n 0.00864761f $X=5 $Y=1.99 $X2=0 $Y2=0
cc_643 N_A_203_47#_c_782_n N_VPWR_c_1332_n 0.00654625f $X=7.76 $Y=1.99 $X2=0
+ $Y2=0
cc_644 N_A_203_47#_c_767_n N_VPWR_c_1332_n 0.00196481f $X=4.99 $Y=1.74 $X2=0
+ $Y2=0
cc_645 N_A_203_47#_c_780_n N_VPWR_c_1332_n 0.00418267f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_646 N_A_203_47#_c_771_n N_A_608_369#_c_1507_n 0.00642978f $X=5.045 $Y=0.805
+ $X2=0 $Y2=0
cc_647 N_A_203_47#_c_771_n N_A_608_369#_c_1485_n 0.0286775f $X=5.045 $Y=0.805
+ $X2=0 $Y2=0
cc_648 N_A_203_47#_c_771_n N_A_608_369#_c_1486_n 0.00791492f $X=5.045 $Y=0.805
+ $X2=0 $Y2=0
cc_649 N_A_203_47#_c_781_n N_A_608_369#_c_1488_n 0.00543259f $X=5 $Y=1.99 $X2=0
+ $Y2=0
cc_650 N_A_203_47#_c_767_n N_A_608_369#_c_1488_n 0.0594075f $X=4.99 $Y=1.74
+ $X2=0 $Y2=0
cc_651 N_A_203_47#_c_771_n N_A_608_369#_c_1488_n 0.0123751f $X=5.045 $Y=0.805
+ $X2=0 $Y2=0
cc_652 N_A_203_47#_c_776_n N_A_608_369#_c_1488_n 0.0127869f $X=5.45 $Y=0.87
+ $X2=0 $Y2=0
cc_653 N_A_203_47#_c_771_n N_A_608_369#_c_1489_n 0.00506513f $X=5.045 $Y=0.805
+ $X2=0 $Y2=0
cc_654 N_A_203_47#_c_776_n N_A_608_369#_c_1489_n 6.01474e-19 $X=5.45 $Y=0.87
+ $X2=0 $Y2=0
cc_655 N_A_203_47#_c_771_n N_A_608_369#_c_1490_n 0.00562077f $X=5.045 $Y=0.805
+ $X2=0 $Y2=0
cc_656 N_A_203_47#_c_772_n N_A_608_369#_c_1490_n 9.47294e-19 $X=5.385 $Y=0.805
+ $X2=0 $Y2=0
cc_657 N_A_203_47#_c_776_n N_A_608_369#_c_1490_n 0.0121034f $X=5.45 $Y=0.87
+ $X2=0 $Y2=0
cc_658 N_A_203_47#_c_781_n N_A_608_369#_c_1494_n 0.0110623f $X=5 $Y=1.99 $X2=0
+ $Y2=0
cc_659 N_A_203_47#_c_767_n N_A_608_369#_c_1494_n 0.00558961f $X=4.99 $Y=1.74
+ $X2=0 $Y2=0
cc_660 N_A_203_47#_c_771_n N_VGND_c_1633_n 0.00116876f $X=5.045 $Y=0.805 $X2=0
+ $Y2=0
cc_661 N_A_203_47#_c_771_n N_VGND_c_1634_n 8.73533e-19 $X=5.045 $Y=0.805 $X2=0
+ $Y2=0
cc_662 N_A_203_47#_c_774_n N_VGND_c_1635_n 0.00197442f $X=7.23 $Y=0.805 $X2=0
+ $Y2=0
cc_663 N_A_203_47#_c_770_n N_VGND_c_1638_n 4.93882e-19 $X=1.385 $Y=0.805 $X2=0
+ $Y2=0
cc_664 N_A_203_47#_c_780_n N_VGND_c_1638_n 0.0101403f $X=1.2 $Y=0.51 $X2=0 $Y2=0
cc_665 N_A_203_47#_c_772_n N_VGND_c_1642_n 4.34458e-19 $X=5.385 $Y=0.805 $X2=0
+ $Y2=0
cc_666 N_A_203_47#_c_776_n N_VGND_c_1642_n 0.00334975f $X=5.45 $Y=0.87 $X2=0
+ $Y2=0
cc_667 N_A_203_47#_c_777_n N_VGND_c_1642_n 0.0037981f $X=5.45 $Y=0.705 $X2=0
+ $Y2=0
cc_668 N_A_203_47#_c_769_n N_VGND_c_1647_n 0.00256736f $X=7.735 $Y=0.87 $X2=0
+ $Y2=0
cc_669 N_A_203_47#_c_773_n N_VGND_c_1647_n 7.48069e-19 $X=7.395 $Y=0.805 $X2=0
+ $Y2=0
cc_670 N_A_203_47#_c_778_n N_VGND_c_1647_n 6.76248e-19 $X=7.365 $Y=0.87 $X2=0
+ $Y2=0
cc_671 N_A_203_47#_c_779_n N_VGND_c_1647_n 0.00424048f $X=7.365 $Y=0.705 $X2=0
+ $Y2=0
cc_672 N_A_203_47#_M1007_d N_VGND_c_1649_n 0.00503858f $X=1.015 $Y=0.235 $X2=0
+ $Y2=0
cc_673 N_A_203_47#_c_769_n N_VGND_c_1649_n 0.00151201f $X=7.735 $Y=0.87 $X2=0
+ $Y2=0
cc_674 N_A_203_47#_c_770_n N_VGND_c_1649_n 0.0161544f $X=1.385 $Y=0.805 $X2=0
+ $Y2=0
cc_675 N_A_203_47#_c_771_n N_VGND_c_1649_n 0.169182f $X=5.045 $Y=0.805 $X2=0
+ $Y2=0
cc_676 N_A_203_47#_c_772_n N_VGND_c_1649_n 0.0202259f $X=5.385 $Y=0.805 $X2=0
+ $Y2=0
cc_677 N_A_203_47#_c_773_n N_VGND_c_1649_n 0.0182227f $X=7.395 $Y=0.805 $X2=0
+ $Y2=0
cc_678 N_A_203_47#_c_774_n N_VGND_c_1649_n 0.0851539f $X=7.23 $Y=0.805 $X2=0
+ $Y2=0
cc_679 N_A_203_47#_c_776_n N_VGND_c_1649_n 0.00195657f $X=5.45 $Y=0.87 $X2=0
+ $Y2=0
cc_680 N_A_203_47#_c_777_n N_VGND_c_1649_n 0.00579376f $X=5.45 $Y=0.705 $X2=0
+ $Y2=0
cc_681 N_A_203_47#_c_778_n N_VGND_c_1649_n 4.46961e-19 $X=7.365 $Y=0.87 $X2=0
+ $Y2=0
cc_682 N_A_203_47#_c_779_n N_VGND_c_1649_n 0.00605236f $X=7.365 $Y=0.705 $X2=0
+ $Y2=0
cc_683 N_A_203_47#_c_780_n N_VGND_c_1649_n 0.00363393f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_684 N_A_203_47#_c_780_n N_VGND_c_1650_n 0.00751197f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_685 N_A_1189_21#_c_969_n N_A_1011_47#_c_1064_n 0.00443215f $X=6.045 $Y=1.89
+ $X2=0 $Y2=0
cc_686 N_A_1189_21#_c_975_n N_A_1011_47#_c_1064_n 0.00751995f $X=6.045 $Y=1.99
+ $X2=0 $Y2=0
cc_687 N_A_1189_21#_c_972_n N_A_1011_47#_c_1064_n 0.0034626f $X=6.975 $Y=2.3
+ $X2=0 $Y2=0
cc_688 N_A_1189_21#_M1005_g N_A_1011_47#_M1012_g 0.0105723f $X=6.02 $Y=0.445
+ $X2=0 $Y2=0
cc_689 N_A_1189_21#_c_969_n N_A_1011_47#_M1012_g 0.00556587f $X=6.045 $Y=1.89
+ $X2=0 $Y2=0
cc_690 N_A_1189_21#_c_970_n N_A_1011_47#_M1012_g 0.0137737f $X=6.775 $Y=0.93
+ $X2=0 $Y2=0
cc_691 N_A_1189_21#_c_971_n N_A_1011_47#_M1012_g 0.00764307f $X=6.13 $Y=0.93
+ $X2=0 $Y2=0
cc_692 N_A_1189_21#_c_998_n N_A_1011_47#_M1012_g 0.00823318f $X=6.917 $Y=0.765
+ $X2=0 $Y2=0
cc_693 N_A_1189_21#_c_972_n N_A_1011_47#_M1012_g 0.0120894f $X=6.975 $Y=2.3
+ $X2=0 $Y2=0
cc_694 N_A_1189_21#_c_1002_n N_A_1011_47#_M1012_g 0.00587221f $X=7.095 $Y=0.45
+ $X2=0 $Y2=0
cc_695 N_A_1189_21#_c_973_n N_A_1011_47#_M1012_g 0.0094035f $X=6.917 $Y=0.93
+ $X2=0 $Y2=0
cc_696 N_A_1189_21#_c_969_n N_A_1011_47#_c_1061_n 0.0177187f $X=6.045 $Y=1.89
+ $X2=0 $Y2=0
cc_697 N_A_1189_21#_c_970_n N_A_1011_47#_c_1061_n 0.0077389f $X=6.775 $Y=0.93
+ $X2=0 $Y2=0
cc_698 N_A_1189_21#_c_969_n N_A_1011_47#_c_1062_n 0.00223289f $X=6.045 $Y=1.89
+ $X2=0 $Y2=0
cc_699 N_A_1189_21#_c_975_n N_A_1011_47#_c_1076_n 0.0108018f $X=6.045 $Y=1.99
+ $X2=0 $Y2=0
cc_700 N_A_1189_21#_M1005_g N_A_1011_47#_c_1080_n 0.00207438f $X=6.02 $Y=0.445
+ $X2=0 $Y2=0
cc_701 N_A_1189_21#_M1005_g N_A_1011_47#_c_1063_n 0.0160733f $X=6.02 $Y=0.445
+ $X2=0 $Y2=0
cc_702 N_A_1189_21#_c_970_n N_A_1011_47#_c_1063_n 0.0245772f $X=6.775 $Y=0.93
+ $X2=0 $Y2=0
cc_703 N_A_1189_21#_c_969_n N_A_1011_47#_c_1067_n 0.00843684f $X=6.045 $Y=1.89
+ $X2=0 $Y2=0
cc_704 N_A_1189_21#_c_975_n N_A_1011_47#_c_1067_n 0.00928103f $X=6.045 $Y=1.99
+ $X2=0 $Y2=0
cc_705 N_A_1189_21#_c_972_n N_A_1011_47#_c_1067_n 0.00615785f $X=6.975 $Y=2.3
+ $X2=0 $Y2=0
cc_706 N_A_1189_21#_c_969_n N_A_1011_47#_c_1068_n 0.0154376f $X=6.045 $Y=1.89
+ $X2=0 $Y2=0
cc_707 N_A_1189_21#_c_970_n N_A_1011_47#_c_1068_n 0.0116171f $X=6.775 $Y=0.93
+ $X2=0 $Y2=0
cc_708 N_A_1189_21#_c_971_n N_A_1011_47#_c_1068_n 6.09916e-19 $X=6.13 $Y=0.93
+ $X2=0 $Y2=0
cc_709 N_A_1189_21#_c_970_n N_A_1011_47#_c_1069_n 0.0272897f $X=6.775 $Y=0.93
+ $X2=0 $Y2=0
cc_710 N_A_1189_21#_c_971_n N_A_1011_47#_c_1069_n 4.18624e-19 $X=6.13 $Y=0.93
+ $X2=0 $Y2=0
cc_711 N_A_1189_21#_c_972_n N_A_1011_47#_c_1069_n 0.0208622f $X=6.975 $Y=2.3
+ $X2=0 $Y2=0
cc_712 N_A_1189_21#_c_972_n N_A_1474_413#_c_1258_n 0.01227f $X=6.975 $Y=2.3
+ $X2=0 $Y2=0
cc_713 N_A_1189_21#_c_1002_n N_A_1474_413#_c_1261_n 0.0128757f $X=7.095 $Y=0.45
+ $X2=0 $Y2=0
cc_714 N_A_1189_21#_c_969_n N_VPWR_c_1336_n 4.19095e-19 $X=6.045 $Y=1.89 $X2=0
+ $Y2=0
cc_715 N_A_1189_21#_c_975_n N_VPWR_c_1336_n 0.00562055f $X=6.045 $Y=1.99 $X2=0
+ $Y2=0
cc_716 N_A_1189_21#_c_972_n N_VPWR_c_1336_n 0.0162643f $X=6.975 $Y=2.3 $X2=0
+ $Y2=0
cc_717 N_A_1189_21#_c_975_n N_VPWR_c_1341_n 0.00457093f $X=6.045 $Y=1.99 $X2=0
+ $Y2=0
cc_718 N_A_1189_21#_c_972_n N_VPWR_c_1347_n 0.0131951f $X=6.975 $Y=2.3 $X2=0
+ $Y2=0
cc_719 N_A_1189_21#_M1025_d N_VPWR_c_1332_n 0.00356119f $X=6.83 $Y=1.735 $X2=0
+ $Y2=0
cc_720 N_A_1189_21#_c_975_n N_VPWR_c_1332_n 0.00675697f $X=6.045 $Y=1.99 $X2=0
+ $Y2=0
cc_721 N_A_1189_21#_c_972_n N_VPWR_c_1332_n 0.00372404f $X=6.975 $Y=2.3 $X2=0
+ $Y2=0
cc_722 N_A_1189_21#_c_970_n N_VGND_M1005_d 0.00306693f $X=6.775 $Y=0.93 $X2=0
+ $Y2=0
cc_723 N_A_1189_21#_M1005_g N_VGND_c_1635_n 0.00917212f $X=6.02 $Y=0.445 $X2=0
+ $Y2=0
cc_724 N_A_1189_21#_c_970_n N_VGND_c_1635_n 0.0261026f $X=6.775 $Y=0.93 $X2=0
+ $Y2=0
cc_725 N_A_1189_21#_c_971_n N_VGND_c_1635_n 4.99767e-19 $X=6.13 $Y=0.93 $X2=0
+ $Y2=0
cc_726 N_A_1189_21#_c_998_n N_VGND_c_1635_n 0.00370702f $X=6.917 $Y=0.765 $X2=0
+ $Y2=0
cc_727 N_A_1189_21#_c_1002_n N_VGND_c_1635_n 0.0130144f $X=7.095 $Y=0.45 $X2=0
+ $Y2=0
cc_728 N_A_1189_21#_M1005_g N_VGND_c_1642_n 0.00585385f $X=6.02 $Y=0.445 $X2=0
+ $Y2=0
cc_729 N_A_1189_21#_c_1002_n N_VGND_c_1647_n 0.0161142f $X=7.095 $Y=0.45 $X2=0
+ $Y2=0
cc_730 N_A_1189_21#_M1012_d N_VGND_c_1649_n 0.00269568f $X=6.84 $Y=0.235 $X2=0
+ $Y2=0
cc_731 N_A_1189_21#_M1005_g N_VGND_c_1649_n 0.00711557f $X=6.02 $Y=0.445 $X2=0
+ $Y2=0
cc_732 N_A_1189_21#_c_970_n N_VGND_c_1649_n 0.00901003f $X=6.775 $Y=0.93 $X2=0
+ $Y2=0
cc_733 N_A_1189_21#_c_1002_n N_VGND_c_1649_n 0.00733201f $X=7.095 $Y=0.45 $X2=0
+ $Y2=0
cc_734 N_A_1011_47#_c_1076_n N_VPWR_M1000_d 0.00207853f $X=6.045 $Y=2.275 $X2=0
+ $Y2=0
cc_735 N_A_1011_47#_c_1067_n N_VPWR_M1000_d 0.00430275f $X=6.137 $Y=2.19 $X2=0
+ $Y2=0
cc_736 N_A_1011_47#_c_1064_n N_VPWR_c_1336_n 0.00576644f $X=6.74 $Y=1.66 $X2=0
+ $Y2=0
cc_737 N_A_1011_47#_c_1061_n N_VPWR_c_1336_n 9.61279e-19 $X=6.64 $Y=1.41 $X2=0
+ $Y2=0
cc_738 N_A_1011_47#_c_1076_n N_VPWR_c_1336_n 0.0138308f $X=6.045 $Y=2.275 $X2=0
+ $Y2=0
cc_739 N_A_1011_47#_c_1067_n N_VPWR_c_1336_n 0.025477f $X=6.137 $Y=2.19 $X2=0
+ $Y2=0
cc_740 N_A_1011_47#_c_1069_n N_VPWR_c_1336_n 0.0073199f $X=6.52 $Y=1.41 $X2=0
+ $Y2=0
cc_741 N_A_1011_47#_c_1076_n N_VPWR_c_1341_n 0.0401946f $X=6.045 $Y=2.275 $X2=0
+ $Y2=0
cc_742 N_A_1011_47#_c_1064_n N_VPWR_c_1347_n 0.00702461f $X=6.74 $Y=1.66 $X2=0
+ $Y2=0
cc_743 N_A_1011_47#_M1014_d N_VPWR_c_1332_n 0.00230779f $X=5.09 $Y=2.065 $X2=0
+ $Y2=0
cc_744 N_A_1011_47#_c_1064_n N_VPWR_c_1332_n 0.00801852f $X=6.74 $Y=1.66 $X2=0
+ $Y2=0
cc_745 N_A_1011_47#_c_1076_n N_VPWR_c_1332_n 0.0179762f $X=6.045 $Y=2.275 $X2=0
+ $Y2=0
cc_746 N_A_1011_47#_c_1080_n N_A_608_369#_c_1489_n 0.0114634f $X=5.705 $Y=0.45
+ $X2=0 $Y2=0
cc_747 N_A_1011_47#_c_1076_n N_A_608_369#_c_1494_n 0.0102205f $X=6.045 $Y=2.275
+ $X2=0 $Y2=0
cc_748 N_A_1011_47#_c_1076_n A_1121_413# 0.00508444f $X=6.045 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_749 N_A_1011_47#_M1012_g N_VGND_c_1635_n 0.00920087f $X=6.765 $Y=0.555 $X2=0
+ $Y2=0
cc_750 N_A_1011_47#_c_1080_n N_VGND_c_1635_n 0.00855527f $X=5.705 $Y=0.45 $X2=0
+ $Y2=0
cc_751 N_A_1011_47#_c_1063_n N_VGND_c_1635_n 0.0022438f $X=5.79 $Y=1.315 $X2=0
+ $Y2=0
cc_752 N_A_1011_47#_c_1080_n N_VGND_c_1642_n 0.0261432f $X=5.705 $Y=0.45 $X2=0
+ $Y2=0
cc_753 N_A_1011_47#_M1012_g N_VGND_c_1647_n 0.00496302f $X=6.765 $Y=0.555 $X2=0
+ $Y2=0
cc_754 N_A_1011_47#_M1026_d N_VGND_c_1649_n 0.00263646f $X=5.055 $Y=0.235 $X2=0
+ $Y2=0
cc_755 N_A_1011_47#_M1012_g N_VGND_c_1649_n 0.00649763f $X=6.765 $Y=0.555 $X2=0
+ $Y2=0
cc_756 N_A_1011_47#_c_1080_n N_VGND_c_1649_n 0.011136f $X=5.705 $Y=0.45 $X2=0
+ $Y2=0
cc_757 N_A_1011_47#_c_1080_n A_1117_47# 0.00665246f $X=5.705 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_758 N_A_1011_47#_c_1063_n A_1117_47# 0.00333286f $X=5.79 $Y=1.315 $X2=-0.19
+ $Y2=-0.24
cc_759 N_A_1647_21#_c_1170_n N_A_1474_413#_c_1253_n 0.00271108f $X=8.335 $Y=1.99
+ $X2=0 $Y2=0
cc_760 N_A_1647_21#_c_1165_n N_A_1474_413#_c_1253_n 0.0182096f $X=9.91 $Y=1.41
+ $X2=0 $Y2=0
cc_761 N_A_1647_21#_c_1182_p N_A_1474_413#_c_1253_n 0.00777604f $X=9.205 $Y=1.95
+ $X2=0 $Y2=0
cc_762 N_A_1647_21#_c_1173_n N_A_1474_413#_c_1253_n 0.00606137f $X=9.312
+ $Y=1.575 $X2=0 $Y2=0
cc_763 N_A_1647_21#_c_1184_p N_A_1474_413#_c_1253_n 0.00844135f $X=9.262 $Y=1.74
+ $X2=0 $Y2=0
cc_764 N_A_1647_21#_c_1164_n N_A_1474_413#_c_1247_n 0.0211139f $X=9.885 $Y=0.995
+ $X2=0 $Y2=0
cc_765 N_A_1647_21#_c_1166_n N_A_1474_413#_c_1247_n 0.00459902f $X=9.31 $Y=0.995
+ $X2=0 $Y2=0
cc_766 N_A_1647_21#_c_1168_n N_A_1474_413#_c_1247_n 0.00597533f $X=9.205
+ $Y=0.385 $X2=0 $Y2=0
cc_767 N_A_1647_21#_M1008_g N_A_1474_413#_c_1248_n 0.00781812f $X=8.31 $Y=0.445
+ $X2=0 $Y2=0
cc_768 N_A_1647_21#_c_1172_n N_A_1474_413#_c_1248_n 0.00734699f $X=9.12 $Y=1.74
+ $X2=0 $Y2=0
cc_769 N_A_1647_21#_c_1168_n N_A_1474_413#_c_1248_n 0.00747686f $X=9.205
+ $Y=0.385 $X2=0 $Y2=0
cc_770 N_A_1647_21#_c_1184_p N_A_1474_413#_c_1248_n 0.00407845f $X=9.262 $Y=1.74
+ $X2=0 $Y2=0
cc_771 N_A_1647_21#_c_1192_p N_A_1474_413#_c_1248_n 0.0141721f $X=9.312 $Y=1.16
+ $X2=0 $Y2=0
cc_772 N_A_1647_21#_c_1165_n N_A_1474_413#_c_1249_n 0.0211139f $X=9.91 $Y=1.41
+ $X2=0 $Y2=0
cc_773 N_A_1647_21#_c_1173_n N_A_1474_413#_c_1249_n 0.00342329f $X=9.312
+ $Y=1.575 $X2=0 $Y2=0
cc_774 N_A_1647_21#_c_1167_n N_A_1474_413#_c_1249_n 0.0206668f $X=9.945 $Y=1.16
+ $X2=0 $Y2=0
cc_775 N_A_1647_21#_c_1192_p N_A_1474_413#_c_1249_n 0.00346806f $X=9.312 $Y=1.16
+ $X2=0 $Y2=0
cc_776 N_A_1647_21#_c_1170_n N_A_1474_413#_c_1258_n 0.00532082f $X=8.335 $Y=1.99
+ $X2=0 $Y2=0
cc_777 N_A_1647_21#_M1008_g N_A_1474_413#_c_1261_n 0.0050536f $X=8.31 $Y=0.445
+ $X2=0 $Y2=0
cc_778 N_A_1647_21#_M1008_g N_A_1474_413#_c_1250_n 0.020596f $X=8.31 $Y=0.445
+ $X2=0 $Y2=0
cc_779 N_A_1647_21#_M1008_g N_A_1474_413#_c_1256_n 0.0140353f $X=8.31 $Y=0.445
+ $X2=0 $Y2=0
cc_780 N_A_1647_21#_c_1170_n N_A_1474_413#_c_1256_n 0.0209368f $X=8.335 $Y=1.99
+ $X2=0 $Y2=0
cc_781 N_A_1647_21#_c_1172_n N_A_1474_413#_c_1256_n 0.0249855f $X=9.12 $Y=1.74
+ $X2=0 $Y2=0
cc_782 N_A_1647_21#_M1008_g N_A_1474_413#_c_1251_n 0.0178907f $X=8.31 $Y=0.445
+ $X2=0 $Y2=0
cc_783 N_A_1647_21#_c_1170_n N_A_1474_413#_c_1251_n 0.00752012f $X=8.335 $Y=1.99
+ $X2=0 $Y2=0
cc_784 N_A_1647_21#_c_1172_n N_A_1474_413#_c_1251_n 0.0359918f $X=9.12 $Y=1.74
+ $X2=0 $Y2=0
cc_785 N_A_1647_21#_c_1168_n N_A_1474_413#_c_1251_n 7.42989e-19 $X=9.205
+ $Y=0.385 $X2=0 $Y2=0
cc_786 N_A_1647_21#_c_1192_p N_A_1474_413#_c_1251_n 0.0277655f $X=9.312 $Y=1.16
+ $X2=0 $Y2=0
cc_787 N_A_1647_21#_M1008_g N_A_1474_413#_c_1252_n 0.004115f $X=8.31 $Y=0.445
+ $X2=0 $Y2=0
cc_788 N_A_1647_21#_c_1170_n N_VPWR_c_1337_n 0.016422f $X=8.335 $Y=1.99 $X2=0
+ $Y2=0
cc_789 N_A_1647_21#_c_1172_n N_VPWR_c_1337_n 0.018568f $X=9.12 $Y=1.74 $X2=0
+ $Y2=0
cc_790 N_A_1647_21#_c_1182_p N_VPWR_c_1337_n 0.0148444f $X=9.205 $Y=1.95 $X2=0
+ $Y2=0
cc_791 N_A_1647_21#_c_1165_n N_VPWR_c_1338_n 0.00699339f $X=9.91 $Y=1.41 $X2=0
+ $Y2=0
cc_792 N_A_1647_21#_c_1182_p N_VPWR_c_1338_n 0.0375787f $X=9.205 $Y=1.95 $X2=0
+ $Y2=0
cc_793 N_A_1647_21#_c_1167_n N_VPWR_c_1338_n 0.00968518f $X=9.945 $Y=1.16 $X2=0
+ $Y2=0
cc_794 N_A_1647_21#_c_1184_p N_VPWR_c_1338_n 0.0206045f $X=9.262 $Y=1.74 $X2=0
+ $Y2=0
cc_795 N_A_1647_21#_c_1182_p N_VPWR_c_1343_n 0.0166993f $X=9.205 $Y=1.95 $X2=0
+ $Y2=0
cc_796 N_A_1647_21#_c_1170_n N_VPWR_c_1347_n 0.00670191f $X=8.335 $Y=1.99 $X2=0
+ $Y2=0
cc_797 N_A_1647_21#_c_1165_n N_VPWR_c_1348_n 0.00604256f $X=9.91 $Y=1.41 $X2=0
+ $Y2=0
cc_798 N_A_1647_21#_M1024_s N_VPWR_c_1332_n 0.00242267f $X=9.08 $Y=1.485 $X2=0
+ $Y2=0
cc_799 N_A_1647_21#_c_1170_n N_VPWR_c_1332_n 0.0136918f $X=8.335 $Y=1.99 $X2=0
+ $Y2=0
cc_800 N_A_1647_21#_c_1165_n N_VPWR_c_1332_n 0.011153f $X=9.91 $Y=1.41 $X2=0
+ $Y2=0
cc_801 N_A_1647_21#_c_1172_n N_VPWR_c_1332_n 0.0145324f $X=9.12 $Y=1.74 $X2=0
+ $Y2=0
cc_802 N_A_1647_21#_c_1182_p N_VPWR_c_1332_n 0.0105267f $X=9.205 $Y=1.95 $X2=0
+ $Y2=0
cc_803 N_A_1647_21#_c_1164_n N_Q_c_1607_n 0.00699388f $X=9.885 $Y=0.995 $X2=0
+ $Y2=0
cc_804 N_A_1647_21#_c_1165_n N_Q_c_1607_n 0.00373637f $X=9.91 $Y=1.41 $X2=0
+ $Y2=0
cc_805 N_A_1647_21#_c_1167_n N_Q_c_1607_n 0.00529837f $X=9.945 $Y=1.16 $X2=0
+ $Y2=0
cc_806 N_A_1647_21#_c_1168_n N_Q_c_1607_n 0.00386543f $X=9.205 $Y=0.385 $X2=0
+ $Y2=0
cc_807 N_A_1647_21#_c_1165_n Q 0.00888111f $X=9.91 $Y=1.41 $X2=0 $Y2=0
cc_808 N_A_1647_21#_c_1165_n N_Q_c_1610_n 0.00735415f $X=9.91 $Y=1.41 $X2=0
+ $Y2=0
cc_809 N_A_1647_21#_c_1173_n N_Q_c_1610_n 8.77928e-19 $X=9.312 $Y=1.575 $X2=0
+ $Y2=0
cc_810 N_A_1647_21#_c_1167_n N_Q_c_1610_n 0.00536204f $X=9.945 $Y=1.16 $X2=0
+ $Y2=0
cc_811 N_A_1647_21#_c_1184_p N_Q_c_1610_n 0.00163954f $X=9.262 $Y=1.74 $X2=0
+ $Y2=0
cc_812 N_A_1647_21#_c_1164_n N_Q_c_1608_n 0.00376297f $X=9.885 $Y=0.995 $X2=0
+ $Y2=0
cc_813 N_A_1647_21#_c_1165_n N_Q_c_1608_n 0.0131747f $X=9.91 $Y=1.41 $X2=0 $Y2=0
cc_814 N_A_1647_21#_c_1167_n N_Q_c_1608_n 0.0237652f $X=9.945 $Y=1.16 $X2=0
+ $Y2=0
cc_815 N_A_1647_21#_M1008_g N_VGND_c_1636_n 0.0151621f $X=8.31 $Y=0.445 $X2=0
+ $Y2=0
cc_816 N_A_1647_21#_c_1168_n N_VGND_c_1636_n 0.0185593f $X=9.205 $Y=0.385 $X2=0
+ $Y2=0
cc_817 N_A_1647_21#_c_1164_n N_VGND_c_1637_n 0.00309623f $X=9.885 $Y=0.995 $X2=0
+ $Y2=0
cc_818 N_A_1647_21#_c_1167_n N_VGND_c_1637_n 0.00933114f $X=9.945 $Y=1.16 $X2=0
+ $Y2=0
cc_819 N_A_1647_21#_c_1168_n N_VGND_c_1644_n 0.0178335f $X=9.205 $Y=0.385 $X2=0
+ $Y2=0
cc_820 N_A_1647_21#_M1008_g N_VGND_c_1647_n 0.00516796f $X=8.31 $Y=0.445 $X2=0
+ $Y2=0
cc_821 N_A_1647_21#_c_1164_n N_VGND_c_1648_n 0.00543342f $X=9.885 $Y=0.995 $X2=0
+ $Y2=0
cc_822 N_A_1647_21#_M1001_s N_VGND_c_1649_n 0.00253533f $X=9.08 $Y=0.235 $X2=0
+ $Y2=0
cc_823 N_A_1647_21#_M1008_g N_VGND_c_1649_n 0.0104668f $X=8.31 $Y=0.445 $X2=0
+ $Y2=0
cc_824 N_A_1647_21#_c_1164_n N_VGND_c_1649_n 0.0107205f $X=9.885 $Y=0.995 $X2=0
+ $Y2=0
cc_825 N_A_1647_21#_c_1168_n N_VGND_c_1649_n 0.013314f $X=9.205 $Y=0.385 $X2=0
+ $Y2=0
cc_826 N_A_1474_413#_c_1253_n N_VPWR_c_1337_n 0.00215411f $X=9.44 $Y=1.41 $X2=0
+ $Y2=0
cc_827 N_A_1474_413#_c_1253_n N_VPWR_c_1338_n 0.00616442f $X=9.44 $Y=1.41 $X2=0
+ $Y2=0
cc_828 N_A_1474_413#_c_1253_n N_VPWR_c_1343_n 0.00621235f $X=9.44 $Y=1.41 $X2=0
+ $Y2=0
cc_829 N_A_1474_413#_c_1258_n N_VPWR_c_1347_n 0.0323122f $X=8.115 $Y=2.25 $X2=0
+ $Y2=0
cc_830 N_A_1474_413#_M1004_d N_VPWR_c_1332_n 0.00242502f $X=7.37 $Y=2.065 $X2=0
+ $Y2=0
cc_831 N_A_1474_413#_c_1253_n N_VPWR_c_1332_n 0.0119363f $X=9.44 $Y=1.41 $X2=0
+ $Y2=0
cc_832 N_A_1474_413#_c_1258_n N_VPWR_c_1332_n 0.030159f $X=8.115 $Y=2.25 $X2=0
+ $Y2=0
cc_833 N_A_1474_413#_c_1258_n A_1570_413# 0.00944908f $X=8.115 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_834 N_A_1474_413#_c_1256_n A_1570_413# 0.00123507f $X=8.2 $Y=2.165 $X2=-0.19
+ $Y2=-0.24
cc_835 N_A_1474_413#_c_1247_n N_Q_c_1607_n 4.1802e-19 $X=9.465 $Y=0.995 $X2=0
+ $Y2=0
cc_836 N_A_1474_413#_c_1253_n N_Q_c_1610_n 3.97267e-19 $X=9.44 $Y=1.41 $X2=0
+ $Y2=0
cc_837 N_A_1474_413#_c_1247_n N_VGND_c_1636_n 0.00244375f $X=9.465 $Y=0.995
+ $X2=0 $Y2=0
cc_838 N_A_1474_413#_c_1261_n N_VGND_c_1636_n 0.0139611f $X=8.115 $Y=0.45 $X2=0
+ $Y2=0
cc_839 N_A_1474_413#_c_1250_n N_VGND_c_1636_n 0.0058633f $X=8.2 $Y=0.995 $X2=0
+ $Y2=0
cc_840 N_A_1474_413#_c_1251_n N_VGND_c_1636_n 0.0152781f $X=8.965 $Y=1.16 $X2=0
+ $Y2=0
cc_841 N_A_1474_413#_c_1247_n N_VGND_c_1637_n 0.00309623f $X=9.465 $Y=0.995
+ $X2=0 $Y2=0
cc_842 N_A_1474_413#_c_1247_n N_VGND_c_1644_n 0.00572277f $X=9.465 $Y=0.995
+ $X2=0 $Y2=0
cc_843 N_A_1474_413#_c_1261_n N_VGND_c_1647_n 0.0283066f $X=8.115 $Y=0.45 $X2=0
+ $Y2=0
cc_844 N_A_1474_413#_M1018_d N_VGND_c_1649_n 0.00301738f $X=7.38 $Y=0.235 $X2=0
+ $Y2=0
cc_845 N_A_1474_413#_c_1247_n N_VGND_c_1649_n 0.0116721f $X=9.465 $Y=0.995 $X2=0
+ $Y2=0
cc_846 N_A_1474_413#_c_1261_n N_VGND_c_1649_n 0.0263339f $X=8.115 $Y=0.45 $X2=0
+ $Y2=0
cc_847 N_A_1474_413#_c_1261_n A_1581_47# 0.00834876f $X=8.115 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_848 N_A_1474_413#_c_1250_n A_1581_47# 0.00142012f $X=8.2 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_849 N_VPWR_c_1332_n A_504_369# 0.00301127f $X=10.35 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_850 N_VPWR_c_1332_n N_A_608_369#_M1030_d 0.00192656f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_851 N_VPWR_c_1332_n N_A_608_369#_M1014_s 0.002768f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_852 N_VPWR_c_1334_n N_A_608_369#_c_1495_n 0.00527813f $X=2.195 $Y=2.33 $X2=0
+ $Y2=0
cc_853 N_VPWR_c_1335_n N_A_608_369#_c_1495_n 0.0109395f $X=4.195 $Y=2.33 $X2=0
+ $Y2=0
cc_854 N_VPWR_c_1339_n N_A_608_369#_c_1495_n 0.0429697f $X=4.11 $Y=2.72 $X2=0
+ $Y2=0
cc_855 N_VPWR_c_1332_n N_A_608_369#_c_1495_n 0.0157065f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_856 N_VPWR_c_1335_n N_A_608_369#_c_1519_n 0.00457937f $X=4.195 $Y=2.33 $X2=0
+ $Y2=0
cc_857 N_VPWR_M1019_d N_A_608_369#_c_1491_n 0.00399644f $X=4.025 $Y=1.845 $X2=0
+ $Y2=0
cc_858 N_VPWR_c_1335_n N_A_608_369#_c_1491_n 0.0119067f $X=4.195 $Y=2.33 $X2=0
+ $Y2=0
cc_859 N_VPWR_c_1339_n N_A_608_369#_c_1491_n 0.00264158f $X=4.11 $Y=2.72 $X2=0
+ $Y2=0
cc_860 N_VPWR_c_1341_n N_A_608_369#_c_1491_n 0.00429797f $X=6.4 $Y=2.72 $X2=0
+ $Y2=0
cc_861 N_VPWR_c_1332_n N_A_608_369#_c_1491_n 0.00580702f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_862 N_VPWR_c_1335_n N_A_608_369#_c_1494_n 0.0144725f $X=4.195 $Y=2.33 $X2=0
+ $Y2=0
cc_863 N_VPWR_c_1341_n N_A_608_369#_c_1494_n 0.0140749f $X=6.4 $Y=2.72 $X2=0
+ $Y2=0
cc_864 N_VPWR_c_1332_n N_A_608_369#_c_1494_n 0.00421345f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_865 N_VPWR_c_1332_n A_702_369# 0.00224063f $X=10.35 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_866 N_VPWR_c_1332_n A_1121_413# 0.00241113f $X=10.35 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_867 N_VPWR_c_1332_n A_1570_413# 0.00341742f $X=10.35 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_868 N_VPWR_c_1332_n N_Q_M1016_d 0.00223285f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_869 N_VPWR_c_1348_n Q 0.0248083f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_870 N_VPWR_c_1332_n Q 0.0195789f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_871 N_VPWR_c_1338_n N_Q_c_1610_n 0.0590731f $X=9.675 $Y=1.79 $X2=0 $Y2=0
cc_872 N_A_608_369#_c_1495_n A_702_369# 0.00440371f $X=3.72 $Y=2.33 $X2=-0.19
+ $Y2=-0.24
cc_873 N_A_608_369#_c_1519_n A_702_369# 0.00269202f $X=3.805 $Y=2.245 $X2=-0.19
+ $Y2=-0.24
cc_874 N_A_608_369#_c_1492_n A_702_369# 9.64403e-19 $X=3.89 $Y=1.91 $X2=-0.19
+ $Y2=-0.24
cc_875 N_A_608_369#_c_1507_n N_VGND_c_1633_n 0.00427557f $X=3.725 $Y=0.36 $X2=0
+ $Y2=0
cc_876 N_A_608_369#_c_1507_n N_VGND_c_1634_n 0.0110659f $X=3.725 $Y=0.36 $X2=0
+ $Y2=0
cc_877 N_A_608_369#_c_1484_n N_VGND_c_1634_n 0.00463869f $X=3.81 $Y=0.695 $X2=0
+ $Y2=0
cc_878 N_A_608_369#_c_1485_n N_VGND_c_1634_n 0.0142693f $X=4.565 $Y=0.78 $X2=0
+ $Y2=0
cc_879 N_A_608_369#_c_1489_n N_VGND_c_1634_n 0.00958988f $X=4.75 $Y=0.45 $X2=0
+ $Y2=0
cc_880 N_A_608_369#_c_1507_n N_VGND_c_1640_n 0.0409414f $X=3.725 $Y=0.36 $X2=0
+ $Y2=0
cc_881 N_A_608_369#_c_1485_n N_VGND_c_1640_n 0.00337254f $X=4.565 $Y=0.78 $X2=0
+ $Y2=0
cc_882 N_A_608_369#_c_1485_n N_VGND_c_1642_n 0.00402378f $X=4.565 $Y=0.78 $X2=0
+ $Y2=0
cc_883 N_A_608_369#_c_1489_n N_VGND_c_1642_n 0.012161f $X=4.75 $Y=0.45 $X2=0
+ $Y2=0
cc_884 N_A_608_369#_M1003_d N_VGND_c_1649_n 0.00250516f $X=3.075 $Y=0.235 $X2=0
+ $Y2=0
cc_885 N_A_608_369#_M1026_s N_VGND_c_1649_n 0.00195217f $X=4.625 $Y=0.235 $X2=0
+ $Y2=0
cc_886 N_A_608_369#_c_1507_n N_VGND_c_1649_n 0.0135588f $X=3.725 $Y=0.36 $X2=0
+ $Y2=0
cc_887 N_A_608_369#_c_1485_n N_VGND_c_1649_n 0.00576196f $X=4.565 $Y=0.78 $X2=0
+ $Y2=0
cc_888 N_A_608_369#_c_1489_n N_VGND_c_1649_n 0.00544577f $X=4.75 $Y=0.45 $X2=0
+ $Y2=0
cc_889 N_A_608_369#_c_1507_n A_721_47# 0.00210886f $X=3.725 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_890 N_A_608_369#_c_1484_n A_721_47# 0.00225806f $X=3.81 $Y=0.695 $X2=-0.19
+ $Y2=-0.24
cc_891 N_Q_c_1607_n N_VGND_c_1648_n 0.0270615f $X=10.145 $Y=0.395 $X2=0 $Y2=0
cc_892 N_Q_M1031_d N_VGND_c_1649_n 0.00254123f $X=9.96 $Y=0.235 $X2=0 $Y2=0
cc_893 N_Q_c_1607_n N_VGND_c_1649_n 0.019901f $X=10.145 $Y=0.395 $X2=0 $Y2=0
cc_894 N_VGND_c_1649_n A_507_47# 0.00336446f $X=10.35 $Y=0 $X2=-0.19 $Y2=-0.24
cc_895 N_VGND_c_1649_n A_721_47# 0.00152414f $X=10.35 $Y=0 $X2=-0.19 $Y2=-0.24
cc_896 N_VGND_c_1649_n A_1117_47# 0.00301061f $X=10.35 $Y=0 $X2=-0.19 $Y2=-0.24
cc_897 N_VGND_c_1649_n A_1581_47# 0.00280389f $X=10.35 $Y=0 $X2=-0.19 $Y2=-0.24
