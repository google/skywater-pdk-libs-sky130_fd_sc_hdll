* File: sky130_fd_sc_hdll__nor2_4.pxi.spice
* Created: Thu Aug 27 19:15:36 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR2_4%A N_A_c_68_n N_A_M1002_g N_A_c_74_n N_A_M1001_g
+ N_A_c_69_n N_A_M1007_g N_A_c_75_n N_A_M1003_g N_A_c_70_n N_A_M1008_g
+ N_A_c_76_n N_A_M1006_g N_A_c_77_n N_A_M1010_g N_A_c_71_n N_A_M1013_g A A
+ N_A_c_72_n N_A_c_73_n A PM_SKY130_FD_SC_HDLL__NOR2_4%A
x_PM_SKY130_FD_SC_HDLL__NOR2_4%B N_B_c_147_n N_B_M1004_g N_B_c_152_n N_B_M1000_g
+ N_B_c_148_n N_B_M1005_g N_B_c_153_n N_B_M1009_g N_B_c_149_n N_B_M1011_g
+ N_B_c_154_n N_B_M1012_g N_B_c_155_n N_B_M1015_g N_B_c_150_n N_B_M1014_g B
+ N_B_c_159_n N_B_c_151_n B PM_SKY130_FD_SC_HDLL__NOR2_4%B
x_PM_SKY130_FD_SC_HDLL__NOR2_4%A_27_297# N_A_27_297#_M1001_s N_A_27_297#_M1003_s
+ N_A_27_297#_M1010_s N_A_27_297#_M1009_s N_A_27_297#_M1015_s
+ N_A_27_297#_c_233_n N_A_27_297#_c_234_n N_A_27_297#_c_235_n
+ N_A_27_297#_c_275_p N_A_27_297#_c_236_n N_A_27_297#_c_237_n
+ N_A_27_297#_c_252_n N_A_27_297#_c_261_n N_A_27_297#_c_263_n
+ N_A_27_297#_c_238_n N_A_27_297#_c_265_n N_A_27_297#_c_239_n
+ PM_SKY130_FD_SC_HDLL__NOR2_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__NOR2_4%VPWR N_VPWR_M1001_d N_VPWR_M1006_d N_VPWR_c_320_n
+ N_VPWR_c_321_n VPWR N_VPWR_c_322_n N_VPWR_c_323_n N_VPWR_c_324_n
+ N_VPWR_c_319_n N_VPWR_c_326_n N_VPWR_c_327_n PM_SKY130_FD_SC_HDLL__NOR2_4%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR2_4%Y N_Y_M1002_s N_Y_M1008_s N_Y_M1004_d N_Y_M1011_d
+ N_Y_M1000_d N_Y_M1012_d N_Y_c_393_n N_Y_c_379_n N_Y_c_380_n N_Y_c_404_n
+ N_Y_c_381_n N_Y_c_408_n N_Y_c_388_n N_Y_c_452_n N_Y_c_389_n N_Y_c_382_n
+ N_Y_c_428_n N_Y_c_459_n N_Y_c_390_n N_Y_c_383_n N_Y_c_384_n N_Y_c_385_n
+ N_Y_c_386_n N_Y_c_391_n Y PM_SKY130_FD_SC_HDLL__NOR2_4%Y
x_PM_SKY130_FD_SC_HDLL__NOR2_4%VGND N_VGND_M1002_d N_VGND_M1007_d N_VGND_M1013_d
+ N_VGND_M1005_s N_VGND_M1014_s N_VGND_c_504_n N_VGND_c_505_n N_VGND_c_506_n
+ N_VGND_c_507_n N_VGND_c_508_n N_VGND_c_509_n N_VGND_c_510_n N_VGND_c_511_n
+ N_VGND_c_512_n N_VGND_c_513_n N_VGND_c_514_n N_VGND_c_515_n N_VGND_c_516_n
+ VGND N_VGND_c_517_n N_VGND_c_518_n N_VGND_c_519_n
+ PM_SKY130_FD_SC_HDLL__NOR2_4%VGND
cc_1 VNB N_A_c_68_n 0.0218461f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_69_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_3 VNB N_A_c_70_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_4 VNB N_A_c_71_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_5 VNB N_A_c_72_n 0.0151855f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_6 VNB N_A_c_73_n 0.0818134f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_7 VNB N_B_c_147_n 0.0164943f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_8 VNB N_B_c_148_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_9 VNB N_B_c_149_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_10 VNB N_B_c_150_n 0.0201851f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_11 VNB N_B_c_151_n 0.0781893f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_12 VNB N_VPWR_c_319_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_13 VNB N_Y_c_379_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_14 VNB N_Y_c_380_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_15 VNB N_Y_c_381_n 0.0042799f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.202
cc_16 VNB N_Y_c_382_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_17 VNB N_Y_c_383_n 0.0165551f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Y_c_384_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_Y_c_385_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_386_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB Y 0.0245691f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_504_n 0.0103581f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.41
cc_23 VNB N_VGND_c_505_n 0.0337721f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.985
cc_24 VNB N_VGND_c_506_n 0.0198149f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.985
cc_25 VNB N_VGND_c_507_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_26 VNB N_VGND_c_508_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_509_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_28 VNB N_VGND_c_510_n 0.0185415f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=1.202
cc_29 VNB N_VGND_c_511_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_30 VNB N_VGND_c_512_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_31 VNB N_VGND_c_513_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=1.202
cc_32 VNB N_VGND_c_514_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.175
cc_33 VNB N_VGND_c_515_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.175
cc_34 VNB N_VGND_c_516_n 0.00545425f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.175
cc_35 VNB N_VGND_c_517_n 0.0126728f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_518_n 0.240661f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_519_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VPB N_A_c_74_n 0.0198936f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_39 VPB N_A_c_75_n 0.0158033f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_40 VPB N_A_c_76_n 0.015524f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_41 VPB N_A_c_77_n 0.0161001f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_42 VPB N_A_c_73_n 0.0483919f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.202
cc_43 VPB N_B_c_152_n 0.0162388f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_44 VPB N_B_c_153_n 0.0158911f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_45 VPB N_B_c_154_n 0.0158728f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_46 VPB N_B_c_155_n 0.0192164f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_47 VPB N_B_c_151_n 0.0473433f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.16
cc_48 VPB N_A_27_297#_c_233_n 0.011936f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_49 VPB N_A_27_297#_c_234_n 0.0307403f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.985
cc_50 VPB N_A_27_297#_c_235_n 0.00262139f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.985
cc_51 VPB N_A_27_297#_c_236_n 0.00210179f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_52 VPB N_A_27_297#_c_237_n 0.00441003f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_297#_c_238_n 0.00104475f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.202
cc_54 VPB N_A_27_297#_c_239_n 0.0255868f $X=-0.19 $Y=1.305 $X2=0.745 $Y2=1.175
cc_55 VPB N_VPWR_c_320_n 4.04661e-19 $X=-0.19 $Y=1.305 $X2=0.96 $Y2=0.56
cc_56 VPB N_VPWR_c_321_n 0.00229677f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=0.995
cc_57 VPB N_VPWR_c_322_n 0.015553f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.985
cc_58 VPB N_VPWR_c_323_n 0.0140826f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.995
cc_59 VPB N_VPWR_c_324_n 0.0692492f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_60 VPB N_VPWR_c_319_n 0.0538259f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_61 VPB N_VPWR_c_326_n 0.00503453f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=1.202
cc_62 VPB N_VPWR_c_327_n 0.00426137f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.16
cc_63 VPB N_Y_c_388_n 0.00136873f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_64 VPB N_Y_c_389_n 0.0024215f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.16
cc_65 VPB N_Y_c_390_n 0.00295624f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_Y_c_391_n 0.00101112f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB Y 0.0338649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 N_A_c_71_n N_B_c_147_n 0.0248003f $X=1.95 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_69 N_A_c_77_n N_B_c_152_n 0.00980578f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_70 N_A_c_72_n N_B_c_159_n 0.00892702f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_c_73_n N_B_c_159_n 8.75854e-19 $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_72 N_A_c_72_n N_B_c_151_n 7.91431e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_c_73_n N_B_c_151_n 0.0248003f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_74 N_A_c_72_n N_A_27_297#_c_233_n 0.018453f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_c_74_n N_A_27_297#_c_235_n 0.0151435f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_76 N_A_c_75_n N_A_27_297#_c_235_n 0.0164876f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A_c_72_n N_A_27_297#_c_235_n 0.0530179f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_c_73_n N_A_27_297#_c_235_n 0.00953178f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_79 N_A_c_76_n N_A_27_297#_c_236_n 0.01491f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A_c_77_n N_A_27_297#_c_236_n 0.0111858f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_c_72_n N_A_27_297#_c_236_n 0.0439319f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A_c_73_n N_A_27_297#_c_236_n 0.00905881f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_83 N_A_c_77_n N_A_27_297#_c_237_n 0.00359583f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_c_72_n N_A_27_297#_c_237_n 3.67829e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_c_73_n N_A_27_297#_c_237_n 3.8543e-19 $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_86 N_A_c_76_n N_A_27_297#_c_252_n 4.84481e-19 $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_c_77_n N_A_27_297#_c_252_n 0.0132763f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A_c_72_n N_A_27_297#_c_238_n 0.0132791f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A_c_73_n N_A_27_297#_c_238_n 0.00435155f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_90 N_A_c_74_n N_VPWR_c_320_n 0.0171285f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_91 N_A_c_75_n N_VPWR_c_320_n 0.0117009f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A_c_76_n N_VPWR_c_320_n 6.2189e-19 $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_93 N_A_c_75_n N_VPWR_c_321_n 6.52114e-19 $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_c_76_n N_VPWR_c_321_n 0.014932f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A_c_77_n N_VPWR_c_321_n 0.00519421f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A_c_74_n N_VPWR_c_322_n 0.00427505f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A_c_75_n N_VPWR_c_323_n 0.00622633f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A_c_76_n N_VPWR_c_323_n 0.00427505f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A_c_77_n N_VPWR_c_324_n 0.00596194f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A_c_74_n N_VPWR_c_319_n 0.00825932f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_c_75_n N_VPWR_c_319_n 0.0104011f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_c_76_n N_VPWR_c_319_n 0.00732977f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_c_77_n N_VPWR_c_319_n 0.0099828f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_c_68_n N_Y_c_393_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A_c_69_n N_Y_c_393_n 0.00686626f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A_c_70_n N_Y_c_393_n 5.45498e-19 $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_107 N_A_c_69_n N_Y_c_379_n 0.00901745f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A_c_70_n N_Y_c_379_n 0.00901745f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_c_72_n N_Y_c_379_n 0.0397461f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_c_73_n N_Y_c_379_n 0.00345541f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_111 N_A_c_68_n N_Y_c_380_n 0.00266157f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A_c_69_n N_Y_c_380_n 0.00116636f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A_c_72_n N_Y_c_380_n 0.0306016f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_c_73_n N_Y_c_380_n 0.00358305f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_115 N_A_c_69_n N_Y_c_404_n 5.24597e-19 $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A_c_70_n N_Y_c_404_n 0.00651696f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_117 N_A_c_71_n N_Y_c_381_n 0.01152f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A_c_72_n N_Y_c_381_n 0.00658691f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_c_71_n N_Y_c_408_n 5.32212e-19 $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A_c_70_n N_Y_c_384_n 0.00119564f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A_c_72_n N_Y_c_384_n 0.0307352f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_c_73_n N_Y_c_384_n 0.00486271f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_123 N_A_c_68_n N_VGND_c_505_n 0.00496762f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A_c_72_n N_VGND_c_505_n 0.019131f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_c_68_n N_VGND_c_506_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_c_69_n N_VGND_c_506_n 0.00423334f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_c_69_n N_VGND_c_507_n 0.00379224f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A_c_70_n N_VGND_c_507_n 0.00276126f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_c_71_n N_VGND_c_508_n 0.00268723f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_c_70_n N_VGND_c_511_n 0.00423334f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_c_71_n N_VGND_c_511_n 0.00437852f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_c_68_n N_VGND_c_518_n 0.0106014f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_c_69_n N_VGND_c_518_n 0.006093f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_c_70_n N_VGND_c_518_n 0.00608558f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_c_71_n N_VGND_c_518_n 0.00615622f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_136 N_B_c_152_n N_A_27_297#_c_237_n 0.00330119f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_137 N_B_c_159_n N_A_27_297#_c_237_n 3.67829e-19 $X=3.665 $Y=1.16 $X2=0 $Y2=0
cc_138 N_B_c_151_n N_A_27_297#_c_237_n 3.8543e-19 $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_139 N_B_c_152_n N_A_27_297#_c_252_n 0.00892871f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_140 N_B_c_153_n N_A_27_297#_c_252_n 5.45419e-19 $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_141 N_B_c_152_n N_A_27_297#_c_261_n 0.0129846f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_142 N_B_c_153_n N_A_27_297#_c_261_n 0.00812567f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_143 N_B_c_154_n N_A_27_297#_c_263_n 0.010646f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_144 N_B_c_155_n N_A_27_297#_c_263_n 0.00815214f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_145 N_B_c_152_n N_A_27_297#_c_265_n 6.08324e-19 $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_146 N_B_c_153_n N_A_27_297#_c_265_n 0.00957505f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_147 N_B_c_154_n N_A_27_297#_c_265_n 0.00659328f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_148 N_B_c_155_n N_A_27_297#_c_265_n 5.58213e-19 $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_149 N_B_c_154_n N_A_27_297#_c_239_n 6.11111e-19 $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_150 N_B_c_155_n N_A_27_297#_c_239_n 0.0098131f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_151 N_B_c_152_n N_VPWR_c_324_n 0.00429425f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_152 N_B_c_153_n N_VPWR_c_324_n 0.00430873f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_153 N_B_c_154_n N_VPWR_c_324_n 0.00430943f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_154 N_B_c_155_n N_VPWR_c_324_n 0.00430873f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_155 N_B_c_152_n N_VPWR_c_319_n 0.00609019f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_156 N_B_c_153_n N_VPWR_c_319_n 0.00605584f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_157 N_B_c_154_n N_VPWR_c_319_n 0.0060559f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_158 N_B_c_155_n N_VPWR_c_319_n 0.00715103f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_159 N_B_c_147_n N_Y_c_381_n 0.00894227f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_160 N_B_c_159_n N_Y_c_381_n 0.00651491f $X=3.665 $Y=1.16 $X2=0 $Y2=0
cc_161 N_B_c_147_n N_Y_c_408_n 0.00644736f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_162 N_B_c_148_n N_Y_c_408_n 0.00686626f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_163 N_B_c_149_n N_Y_c_408_n 5.45498e-19 $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_164 N_B_c_152_n N_Y_c_388_n 0.00184921f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_165 N_B_c_159_n N_Y_c_388_n 0.0138618f $X=3.665 $Y=1.16 $X2=0 $Y2=0
cc_166 N_B_c_151_n N_Y_c_388_n 0.00436648f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_167 N_B_c_153_n N_Y_c_389_n 0.0155165f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_168 N_B_c_154_n N_Y_c_389_n 0.0161472f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_169 N_B_c_159_n N_Y_c_389_n 0.0568026f $X=3.665 $Y=1.16 $X2=0 $Y2=0
cc_170 N_B_c_151_n N_Y_c_389_n 0.0110865f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_171 N_B_c_148_n N_Y_c_382_n 0.00901745f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B_c_149_n N_Y_c_382_n 0.00901745f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_173 N_B_c_159_n N_Y_c_382_n 0.0397461f $X=3.665 $Y=1.16 $X2=0 $Y2=0
cc_174 N_B_c_151_n N_Y_c_382_n 0.00345541f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_175 N_B_c_148_n N_Y_c_428_n 5.24597e-19 $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_176 N_B_c_149_n N_Y_c_428_n 0.00651696f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_177 N_B_c_155_n N_Y_c_390_n 0.0194908f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_178 N_B_c_159_n N_Y_c_390_n 0.013112f $X=3.665 $Y=1.16 $X2=0 $Y2=0
cc_179 N_B_c_151_n N_Y_c_390_n 0.00205167f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_180 N_B_c_150_n N_Y_c_383_n 0.013507f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_181 N_B_c_159_n N_Y_c_383_n 0.0069316f $X=3.665 $Y=1.16 $X2=0 $Y2=0
cc_182 N_B_c_147_n N_Y_c_385_n 0.00116636f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_183 N_B_c_148_n N_Y_c_385_n 0.00116636f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_184 N_B_c_159_n N_Y_c_385_n 0.0306016f $X=3.665 $Y=1.16 $X2=0 $Y2=0
cc_185 N_B_c_151_n N_Y_c_385_n 0.00358305f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_186 N_B_c_149_n N_Y_c_386_n 0.00119564f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_187 N_B_c_159_n N_Y_c_386_n 0.0307352f $X=3.665 $Y=1.16 $X2=0 $Y2=0
cc_188 N_B_c_151_n N_Y_c_386_n 0.00486271f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_189 N_B_c_159_n N_Y_c_391_n 0.0138618f $X=3.665 $Y=1.16 $X2=0 $Y2=0
cc_190 N_B_c_151_n N_Y_c_391_n 0.00419992f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_191 N_B_c_155_n Y 0.00127274f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_192 N_B_c_150_n Y 0.0178248f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_193 N_B_c_159_n Y 0.0122425f $X=3.665 $Y=1.16 $X2=0 $Y2=0
cc_194 N_B_c_147_n N_VGND_c_508_n 0.00268723f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_195 N_B_c_148_n N_VGND_c_509_n 0.00379224f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_196 N_B_c_149_n N_VGND_c_509_n 0.00276126f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_197 N_B_c_150_n N_VGND_c_510_n 0.00453359f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_198 N_B_c_147_n N_VGND_c_513_n 0.00423334f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_199 N_B_c_148_n N_VGND_c_513_n 0.00423334f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_200 N_B_c_149_n N_VGND_c_515_n 0.00423334f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_201 N_B_c_150_n N_VGND_c_515_n 0.00437852f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_202 N_B_c_147_n N_VGND_c_518_n 0.00587047f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_203 N_B_c_148_n N_VGND_c_518_n 0.006093f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_204 N_B_c_149_n N_VGND_c_518_n 0.00608558f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_205 N_B_c_150_n N_VGND_c_518_n 0.00727267f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A_27_297#_c_235_n N_VPWR_M1001_d 0.00188315f $X=1.135 $Y=1.56 $X2=-0.19
+ $Y2=1.305
cc_207 N_A_27_297#_c_236_n N_VPWR_M1006_d 0.00184035f $X=1.945 $Y=1.56 $X2=0
+ $Y2=0
cc_208 N_A_27_297#_c_234_n N_VPWR_c_320_n 0.0487409f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_209 N_A_27_297#_c_235_n N_VPWR_c_320_n 0.0212439f $X=1.135 $Y=1.56 $X2=0
+ $Y2=0
cc_210 N_A_27_297#_c_275_p N_VPWR_c_320_n 0.0385613f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_211 N_A_27_297#_c_275_p N_VPWR_c_321_n 0.0461742f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_212 N_A_27_297#_c_236_n N_VPWR_c_321_n 0.0194872f $X=1.945 $Y=1.56 $X2=0
+ $Y2=0
cc_213 N_A_27_297#_c_252_n N_VPWR_c_321_n 0.0496968f $X=2.135 $Y=2.295 $X2=0
+ $Y2=0
cc_214 N_A_27_297#_c_234_n N_VPWR_c_322_n 0.019258f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_215 N_A_27_297#_c_275_p N_VPWR_c_323_n 0.0118139f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_216 N_A_27_297#_c_252_n N_VPWR_c_324_n 0.0224921f $X=2.135 $Y=2.295 $X2=0
+ $Y2=0
cc_217 N_A_27_297#_c_261_n N_VPWR_c_324_n 0.0317606f $X=2.885 $Y=2.38 $X2=0
+ $Y2=0
cc_218 N_A_27_297#_c_263_n N_VPWR_c_324_n 0.0317869f $X=3.825 $Y=2.38 $X2=0
+ $Y2=0
cc_219 N_A_27_297#_c_265_n N_VPWR_c_324_n 0.0220286f $X=3.1 $Y=2.02 $X2=0 $Y2=0
cc_220 N_A_27_297#_c_239_n N_VPWR_c_324_n 0.030108f $X=4.04 $Y=2 $X2=0 $Y2=0
cc_221 N_A_27_297#_M1001_s N_VPWR_c_319_n 0.00442207f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_222 N_A_27_297#_M1003_s N_VPWR_c_319_n 0.00647849f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_223 N_A_27_297#_M1010_s N_VPWR_c_319_n 0.00231261f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_224 N_A_27_297#_M1009_s N_VPWR_c_319_n 0.00231261f $X=2.955 $Y=1.485 $X2=0
+ $Y2=0
cc_225 N_A_27_297#_M1015_s N_VPWR_c_319_n 0.00225715f $X=3.895 $Y=1.485 $X2=0
+ $Y2=0
cc_226 N_A_27_297#_c_234_n N_VPWR_c_319_n 0.0105137f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_227 N_A_27_297#_c_275_p N_VPWR_c_319_n 0.00646998f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_228 N_A_27_297#_c_252_n N_VPWR_c_319_n 0.014078f $X=2.135 $Y=2.295 $X2=0
+ $Y2=0
cc_229 N_A_27_297#_c_261_n N_VPWR_c_319_n 0.0196262f $X=2.885 $Y=2.38 $X2=0
+ $Y2=0
cc_230 N_A_27_297#_c_263_n N_VPWR_c_319_n 0.0196297f $X=3.825 $Y=2.38 $X2=0
+ $Y2=0
cc_231 N_A_27_297#_c_265_n N_VPWR_c_319_n 0.0139179f $X=3.1 $Y=2.02 $X2=0 $Y2=0
cc_232 N_A_27_297#_c_239_n N_VPWR_c_319_n 0.0173457f $X=4.04 $Y=2 $X2=0 $Y2=0
cc_233 N_A_27_297#_c_261_n N_Y_M1000_d 0.0034107f $X=2.885 $Y=2.38 $X2=0 $Y2=0
cc_234 N_A_27_297#_c_263_n N_Y_M1012_d 0.00343888f $X=3.825 $Y=2.38 $X2=0 $Y2=0
cc_235 N_A_27_297#_c_237_n N_Y_c_381_n 0.0131084f $X=2.135 $Y=1.665 $X2=0 $Y2=0
cc_236 N_A_27_297#_c_237_n N_Y_c_388_n 0.0150774f $X=2.135 $Y=1.665 $X2=0 $Y2=0
cc_237 N_A_27_297#_c_252_n N_Y_c_388_n 0.00543755f $X=2.135 $Y=2.295 $X2=0 $Y2=0
cc_238 N_A_27_297#_c_252_n N_Y_c_452_n 0.0232292f $X=2.135 $Y=2.295 $X2=0 $Y2=0
cc_239 N_A_27_297#_c_261_n N_Y_c_452_n 0.0128008f $X=2.885 $Y=2.38 $X2=0 $Y2=0
cc_240 N_A_27_297#_c_265_n N_Y_c_452_n 0.0141845f $X=3.1 $Y=2.02 $X2=0 $Y2=0
cc_241 N_A_27_297#_M1009_s N_Y_c_389_n 0.00199621f $X=2.955 $Y=1.485 $X2=0 $Y2=0
cc_242 N_A_27_297#_c_261_n N_Y_c_389_n 0.0030044f $X=2.885 $Y=2.38 $X2=0 $Y2=0
cc_243 N_A_27_297#_c_263_n N_Y_c_389_n 0.00435577f $X=3.825 $Y=2.38 $X2=0 $Y2=0
cc_244 N_A_27_297#_c_265_n N_Y_c_389_n 0.0196167f $X=3.1 $Y=2.02 $X2=0 $Y2=0
cc_245 N_A_27_297#_c_263_n N_Y_c_459_n 0.0128008f $X=3.825 $Y=2.38 $X2=0 $Y2=0
cc_246 N_A_27_297#_c_265_n N_Y_c_459_n 0.0116296f $X=3.1 $Y=2.02 $X2=0 $Y2=0
cc_247 N_A_27_297#_c_239_n N_Y_c_459_n 0.01593f $X=4.04 $Y=2 $X2=0 $Y2=0
cc_248 N_A_27_297#_M1015_s N_Y_c_390_n 0.00180849f $X=3.895 $Y=1.485 $X2=0 $Y2=0
cc_249 N_A_27_297#_c_263_n N_Y_c_390_n 0.0030044f $X=3.825 $Y=2.38 $X2=0 $Y2=0
cc_250 N_A_27_297#_c_239_n N_Y_c_390_n 0.0171956f $X=4.04 $Y=2 $X2=0 $Y2=0
cc_251 N_A_27_297#_M1015_s Y 0.00203659f $X=3.895 $Y=1.485 $X2=0 $Y2=0
cc_252 N_A_27_297#_c_239_n Y 0.0176151f $X=4.04 $Y=2 $X2=0 $Y2=0
cc_253 N_A_27_297#_c_233_n N_VGND_c_505_n 0.00202255f $X=0.227 $Y=1.665 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_319_n N_Y_M1000_d 0.00232895f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_255 N_VPWR_c_319_n N_Y_M1012_d 0.00232895f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_256 N_Y_c_379_n N_VGND_M1007_d 0.00251047f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_257 N_Y_c_381_n N_VGND_M1013_d 0.00162089f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_258 N_Y_c_382_n N_VGND_M1005_s 0.00251047f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_259 N_Y_c_383_n N_VGND_M1014_s 0.00282644f $X=4.095 $Y=0.815 $X2=0 $Y2=0
cc_260 N_Y_c_380_n N_VGND_c_505_n 0.00835456f $X=0.915 $Y=0.815 $X2=0 $Y2=0
cc_261 N_Y_c_393_n N_VGND_c_506_n 0.0223596f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_262 N_Y_c_379_n N_VGND_c_506_n 0.00266636f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_263 N_Y_c_393_n N_VGND_c_507_n 0.0183628f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_264 N_Y_c_379_n N_VGND_c_507_n 0.0127273f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_265 N_Y_c_381_n N_VGND_c_508_n 0.0122559f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_266 N_Y_c_408_n N_VGND_c_509_n 0.0183628f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_267 N_Y_c_382_n N_VGND_c_509_n 0.0127273f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_268 N_Y_c_383_n N_VGND_c_510_n 0.0231185f $X=4.095 $Y=0.815 $X2=0 $Y2=0
cc_269 N_Y_c_379_n N_VGND_c_511_n 0.00198695f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_270 N_Y_c_404_n N_VGND_c_511_n 0.0231806f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_271 N_Y_c_381_n N_VGND_c_511_n 0.00254521f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_272 N_Y_c_381_n N_VGND_c_513_n 0.00198695f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_273 N_Y_c_408_n N_VGND_c_513_n 0.0223596f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_274 N_Y_c_382_n N_VGND_c_513_n 0.00266636f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_275 N_Y_c_382_n N_VGND_c_515_n 0.00198695f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_276 N_Y_c_428_n N_VGND_c_515_n 0.0231806f $X=3.57 $Y=0.39 $X2=0 $Y2=0
cc_277 N_Y_c_383_n N_VGND_c_515_n 0.00254521f $X=4.095 $Y=0.815 $X2=0 $Y2=0
cc_278 N_Y_c_383_n N_VGND_c_517_n 0.00424816f $X=4.095 $Y=0.815 $X2=0 $Y2=0
cc_279 N_Y_M1002_s N_VGND_c_518_n 0.0025535f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_280 N_Y_M1008_s N_VGND_c_518_n 0.00304143f $X=1.505 $Y=0.235 $X2=0 $Y2=0
cc_281 N_Y_M1004_d N_VGND_c_518_n 0.0025535f $X=2.445 $Y=0.235 $X2=0 $Y2=0
cc_282 N_Y_M1011_d N_VGND_c_518_n 0.00304143f $X=3.385 $Y=0.235 $X2=0 $Y2=0
cc_283 N_Y_c_393_n N_VGND_c_518_n 0.0141302f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_284 N_Y_c_379_n N_VGND_c_518_n 0.00972452f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_285 N_Y_c_404_n N_VGND_c_518_n 0.0143352f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_286 N_Y_c_381_n N_VGND_c_518_n 0.0094839f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_287 N_Y_c_408_n N_VGND_c_518_n 0.0141302f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_288 N_Y_c_382_n N_VGND_c_518_n 0.00972452f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_289 N_Y_c_428_n N_VGND_c_518_n 0.0143352f $X=3.57 $Y=0.39 $X2=0 $Y2=0
cc_290 N_Y_c_383_n N_VGND_c_518_n 0.0132175f $X=4.095 $Y=0.815 $X2=0 $Y2=0
