* NGSPICE file created from sky130_fd_sc_hdll__mux2_12.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__mux2_12 A0 A1 S VGND VNB VPB VPWR X
M1000 a_119_47# S VGND VNB nshort w=650000u l=150000u
+  ad=7.02e+11p pd=7.36e+06u as=2.9705e+12p ps=2.604e+07u
M1001 VGND a_973_297# a_1163_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.02e+11p ps=7.36e+06u
M1002 a_27_47# A1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.66e+12p pd=1.532e+07u as=1.16e+12p ps=1.032e+07u
M1003 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=3.69e+12p pd=3.338e+07u as=1.74e+12p ps=1.548e+07u
M1004 a_27_47# A0 a_1163_47# VNB nshort w=650000u l=150000u
+  ad=1.287e+12p pd=1.176e+07u as=0p ps=0u
M1005 a_117_297# a_973_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR S a_597_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.16e+12p ps=1.032e+07u
M1007 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_597_297# A0 a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1163_47# a_973_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_47# A0 a_597_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1163_47# A0 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR S a_973_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1013 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.053e+12p pd=1.104e+07u as=0p ps=0u
M1015 a_597_297# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_47# A1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_597_297# A0 a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND S a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_119_47# S VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_973_297# a_1163_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_117_297# A1 a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_973_297# a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_27_47# A0 a_597_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_973_297# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_27_47# A1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_117_297# a_973_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_973_297# S VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1039 VGND S a_973_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_119_47# A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_27_47# A0 a_1163_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPWR S a_597_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_1163_47# a_973_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_1163_47# A0 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_117_297# A1 a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1049 VPWR a_973_297# a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1050 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1051 a_27_47# A1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1052 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1053 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1054 VGND S a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1055 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1056 a_597_297# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1057 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1058 a_119_47# A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1059 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

