* File: sky130_fd_sc_hdll__a32o_4.pxi.spice
* Created: Thu Aug 27 18:56:17 2020
* 
x_PM_SKY130_FD_SC_HDLL__A32O_4%A_79_21# N_A_79_21#_M1016_s N_A_79_21#_M1007_s
+ N_A_79_21#_M1000_d N_A_79_21#_M1009_s N_A_79_21#_c_99_n N_A_79_21#_M1004_g
+ N_A_79_21#_c_108_n N_A_79_21#_M1002_g N_A_79_21#_c_100_n N_A_79_21#_M1006_g
+ N_A_79_21#_c_109_n N_A_79_21#_M1008_g N_A_79_21#_c_101_n N_A_79_21#_M1018_g
+ N_A_79_21#_c_110_n N_A_79_21#_M1015_g N_A_79_21#_c_111_n N_A_79_21#_M1024_g
+ N_A_79_21#_c_102_n N_A_79_21#_M1025_g N_A_79_21#_c_103_n N_A_79_21#_c_113_n
+ N_A_79_21#_c_114_n N_A_79_21#_c_172_p N_A_79_21#_c_104_n N_A_79_21#_c_105_n
+ N_A_79_21#_c_139_p N_A_79_21#_c_140_p N_A_79_21#_c_154_p N_A_79_21#_c_106_n
+ N_A_79_21#_c_151_p N_A_79_21#_c_152_p N_A_79_21#_c_153_p N_A_79_21#_c_107_n
+ PM_SKY130_FD_SC_HDLL__A32O_4%A_79_21#
x_PM_SKY130_FD_SC_HDLL__A32O_4%A3 N_A3_c_278_n N_A3_M1022_g N_A3_c_282_n
+ N_A3_M1005_g N_A3_c_279_n N_A3_M1023_g N_A3_c_283_n N_A3_M1010_g A3 A3
+ N_A3_c_281_n A3 A3 PM_SKY130_FD_SC_HDLL__A32O_4%A3
x_PM_SKY130_FD_SC_HDLL__A32O_4%A2 N_A2_c_332_n N_A2_M1019_g N_A2_c_328_n
+ N_A2_M1001_g N_A2_c_333_n N_A2_M1027_g N_A2_c_329_n N_A2_M1020_g A2
+ N_A2_c_331_n A2 PM_SKY130_FD_SC_HDLL__A32O_4%A2
x_PM_SKY130_FD_SC_HDLL__A32O_4%A1 N_A1_M1016_g N_A1_c_378_n N_A1_M1003_g
+ N_A1_M1026_g N_A1_c_379_n N_A1_M1012_g A1 A1 N_A1_c_376_n A1 A1
+ PM_SKY130_FD_SC_HDLL__A32O_4%A1
x_PM_SKY130_FD_SC_HDLL__A32O_4%B1 N_B1_M1007_g N_B1_c_426_n N_B1_M1000_g
+ N_B1_M1017_g N_B1_c_427_n N_B1_M1021_g B1 B1 N_B1_c_425_n
+ N_B1_X29_noxref_CONDUCTOR B1 B1 PM_SKY130_FD_SC_HDLL__A32O_4%B1
x_PM_SKY130_FD_SC_HDLL__A32O_4%B2 N_B2_M1011_g N_B2_c_480_n N_B2_M1009_g
+ N_B2_M1014_g N_B2_c_481_n N_B2_M1013_g N_B2_c_477_n B2 B2 B2 N_B2_c_479_n
+ N_B2_c_497_n B2 PM_SKY130_FD_SC_HDLL__A32O_4%B2
x_PM_SKY130_FD_SC_HDLL__A32O_4%VPWR N_VPWR_M1002_d N_VPWR_M1008_d N_VPWR_M1024_d
+ N_VPWR_M1010_d N_VPWR_M1019_s N_VPWR_M1003_s N_VPWR_c_521_n N_VPWR_c_522_n
+ N_VPWR_c_523_n N_VPWR_c_524_n N_VPWR_c_525_n N_VPWR_c_526_n VPWR
+ N_VPWR_c_527_n N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_520_n
+ N_VPWR_c_532_n N_VPWR_c_533_n N_VPWR_c_534_n N_VPWR_c_535_n N_VPWR_c_536_n
+ PM_SKY130_FD_SC_HDLL__A32O_4%VPWR
x_PM_SKY130_FD_SC_HDLL__A32O_4%X N_X_M1004_d N_X_M1018_d N_X_M1002_s N_X_M1015_s
+ N_X_c_655_n N_X_c_658_n N_X_c_659_n N_X_c_660_n N_X_c_662_n N_X_c_667_n
+ N_X_c_673_n N_X_c_675_n N_X_c_677_n N_X_c_679_n X X X N_X_c_651_n N_X_c_653_n
+ X PM_SKY130_FD_SC_HDLL__A32O_4%X
x_PM_SKY130_FD_SC_HDLL__A32O_4%A_493_297# N_A_493_297#_M1005_s
+ N_A_493_297#_M1019_d N_A_493_297#_M1027_d N_A_493_297#_M1012_d
+ N_A_493_297#_M1021_s N_A_493_297#_M1013_d N_A_493_297#_c_748_n
+ N_A_493_297#_c_721_n N_A_493_297#_c_735_n N_A_493_297#_c_752_n
+ N_A_493_297#_c_736_n N_A_493_297#_c_756_n N_A_493_297#_c_737_n
+ N_A_493_297#_c_760_n N_A_493_297#_c_739_n N_A_493_297#_c_761_n
+ N_A_493_297#_c_722_n N_A_493_297#_c_723_n N_A_493_297#_c_746_n
+ N_A_493_297#_c_747_n PM_SKY130_FD_SC_HDLL__A32O_4%A_493_297#
x_PM_SKY130_FD_SC_HDLL__A32O_4%VGND N_VGND_M1004_s N_VGND_M1006_s N_VGND_M1025_s
+ N_VGND_M1023_d N_VGND_M1011_s N_VGND_c_812_n N_VGND_c_813_n VGND
+ N_VGND_c_814_n N_VGND_c_815_n N_VGND_c_816_n N_VGND_c_817_n N_VGND_c_818_n
+ N_VGND_c_819_n N_VGND_c_820_n N_VGND_c_821_n N_VGND_c_822_n N_VGND_c_823_n
+ PM_SKY130_FD_SC_HDLL__A32O_4%VGND
x_PM_SKY130_FD_SC_HDLL__A32O_4%A_485_47# N_A_485_47#_M1022_s N_A_485_47#_M1001_d
+ N_A_485_47#_c_927_n N_A_485_47#_c_928_n N_A_485_47#_c_925_n
+ PM_SKY130_FD_SC_HDLL__A32O_4%A_485_47#
x_PM_SKY130_FD_SC_HDLL__A32O_4%A_695_47# N_A_695_47#_M1001_s N_A_695_47#_M1020_s
+ N_A_695_47#_M1026_d N_A_695_47#_c_950_n PM_SKY130_FD_SC_HDLL__A32O_4%A_695_47#
x_PM_SKY130_FD_SC_HDLL__A32O_4%A_1194_47# N_A_1194_47#_M1007_d
+ N_A_1194_47#_M1017_d N_A_1194_47#_M1014_d N_A_1194_47#_c_970_n
+ N_A_1194_47#_c_992_n N_A_1194_47#_c_977_n N_A_1194_47#_c_980_n
+ N_A_1194_47#_c_978_n N_A_1194_47#_c_986_n
+ PM_SKY130_FD_SC_HDLL__A32O_4%A_1194_47#
cc_1 VNB N_A_79_21#_c_99_n 0.0187572f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_100_n 0.0167376f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_3 VNB N_A_79_21#_c_101_n 0.0171868f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_4 VNB N_A_79_21#_c_102_n 0.0166258f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_5 VNB N_A_79_21#_c_103_n 0.00499804f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=1.16
cc_6 VNB N_A_79_21#_c_104_n 0.00911532f $X=-0.19 $Y=-0.24 $X2=5.78 $Y2=0.72
cc_7 VNB N_A_79_21#_c_105_n 0.0126406f $X=-0.19 $Y=-0.24 $X2=5.865 $Y2=1.495
cc_8 VNB N_A_79_21#_c_106_n 0.00464445f $X=-0.19 $Y=-0.24 $X2=6.565 $Y2=0.72
cc_9 VNB N_A_79_21#_c_107_n 0.0764601f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_10 VNB N_A3_c_278_n 0.016461f $X=-0.19 $Y=-0.24 $X2=4.825 $Y2=0.235
cc_11 VNB N_A3_c_279_n 0.0215708f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB A3 0.00646996f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_13 VNB N_A3_c_281_n 0.0533282f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_14 VNB N_A2_c_328_n 0.022465f $X=-0.19 $Y=-0.24 $X2=7.405 $Y2=1.485
cc_15 VNB N_A2_c_329_n 0.0167331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB A2 0.00392606f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_17 VNB N_A2_c_331_n 0.0463869f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_18 VNB N_A1_M1016_g 0.0183466f $X=-0.19 $Y=-0.24 $X2=6.465 $Y2=1.485
cc_19 VNB N_A1_M1026_g 0.0216365f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A1_c_376_n 0.0501765f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_21 VNB A1 0.00186887f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_22 VNB N_B1_M1007_g 0.0218936f $X=-0.19 $Y=-0.24 $X2=6.465 $Y2=1.485
cc_23 VNB N_B1_M1017_g 0.0188099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB B1 0.00651373f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_25 VNB N_B1_c_425_n 0.043742f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_26 VNB N_B2_M1011_g 0.01858f $X=-0.19 $Y=-0.24 $X2=6.465 $Y2=1.485
cc_27 VNB N_B2_M1014_g 0.0246977f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_B2_c_477_n 0.0300932f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_29 VNB B2 0.00887859f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_30 VNB N_B2_c_479_n 0.0266804f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.56
cc_31 VNB N_VPWR_c_520_n 0.345644f $X=-0.19 $Y=-0.24 $X2=5.95 $Y2=1.99
cc_32 VNB N_X_c_651_n 0.0071443f $X=-0.19 $Y=-0.24 $X2=5.78 $Y2=1.58
cc_33 VNB X 0.0238043f $X=-0.19 $Y=-0.24 $X2=5.01 $Y2=0.72
cc_34 VNB N_VGND_c_812_n 0.010303f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_35 VNB N_VGND_c_813_n 0.0126078f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_36 VNB N_VGND_c_814_n 0.0123546f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_37 VNB N_VGND_c_815_n 0.0131442f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.56
cc_38 VNB N_VGND_c_816_n 0.0133958f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_39 VNB N_VGND_c_817_n 0.0962447f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=1.16
cc_40 VNB N_VGND_c_818_n 0.0165472f $X=-0.19 $Y=-0.24 $X2=5.78 $Y2=1.58
cc_41 VNB N_VGND_c_819_n 0.39853f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=1.58
cc_42 VNB N_VGND_c_820_n 0.00537041f $X=-0.19 $Y=-0.24 $X2=5.865 $Y2=1.665
cc_43 VNB N_VGND_c_821_n 0.00537882f $X=-0.19 $Y=-0.24 $X2=7.55 $Y2=2
cc_44 VNB N_VGND_c_822_n 0.0119695f $X=-0.19 $Y=-0.24 $X2=5.865 $Y2=1.58
cc_45 VNB N_VGND_c_823_n 0.0055668f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_46 VNB N_A_485_47#_c_925_n 0.00815884f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_47 VNB N_A_695_47#_c_950_n 0.0047211f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_48 VNB N_A_1194_47#_c_970_n 0.00248626f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VPB N_A_79_21#_c_108_n 0.0183023f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_50 VPB N_A_79_21#_c_109_n 0.0158104f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_51 VPB N_A_79_21#_c_110_n 0.0160869f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_52 VPB N_A_79_21#_c_111_n 0.0154967f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_53 VPB N_A_79_21#_c_103_n 2.19146e-19 $X=-0.19 $Y=1.305 $X2=1.95 $Y2=1.16
cc_54 VPB N_A_79_21#_c_113_n 0.00152104f $X=-0.19 $Y=1.305 $X2=2.06 $Y2=1.495
cc_55 VPB N_A_79_21#_c_114_n 0.00765505f $X=-0.19 $Y=1.305 $X2=5.78 $Y2=1.58
cc_56 VPB N_A_79_21#_c_105_n 0.00438704f $X=-0.19 $Y=1.305 $X2=5.865 $Y2=1.495
cc_57 VPB N_A_79_21#_c_107_n 0.0470623f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_58 VPB N_A3_c_282_n 0.016206f $X=-0.19 $Y=1.305 $X2=7.405 $Y2=1.485
cc_59 VPB N_A3_c_283_n 0.0199635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A3_c_281_n 0.0283026f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_61 VPB N_A2_c_332_n 0.0206372f $X=-0.19 $Y=1.305 $X2=4.825 $Y2=0.235
cc_62 VPB N_A2_c_333_n 0.0162737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB A2 0.00161492f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_64 VPB N_A2_c_331_n 0.0222782f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_65 VPB N_A1_c_378_n 0.0159944f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A1_c_379_n 0.0194127f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A1_c_376_n 0.027108f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=0.995
cc_68 VPB A1 0.00228799f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.56
cc_69 VPB N_B1_c_426_n 0.0192858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_B1_c_427_n 0.0156532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB B1 0.0030869f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_72 VPB N_B1_c_425_n 0.0204048f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_73 VPB N_B2_c_480_n 0.016393f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_B2_c_481_n 0.0210629f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_B2_c_477_n 0.0248092f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_76 VPB B2 0.002587f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_77 VPB N_B2_c_479_n 0.0092983f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=0.56
cc_78 VPB N_VPWR_c_521_n 0.0103693f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.995
cc_79 VPB N_VPWR_c_522_n 0.025861f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_80 VPB N_VPWR_c_523_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=1.41 $Y2=0.995
cc_81 VPB N_VPWR_c_524_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_82 VPB N_VPWR_c_525_n 0.0147977f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_83 VPB N_VPWR_c_526_n 0.0123761f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_84 VPB N_VPWR_c_527_n 0.0140826f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=1.16
cc_85 VPB N_VPWR_c_528_n 0.0140826f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=1.16
cc_86 VPB N_VPWR_c_529_n 0.0133404f $X=-0.19 $Y=1.305 $X2=5.78 $Y2=1.58
cc_87 VPB N_VPWR_c_530_n 0.0747109f $X=-0.19 $Y=1.305 $X2=6.445 $Y2=1.99
cc_88 VPB N_VPWR_c_520_n 0.047749f $X=-0.19 $Y=1.305 $X2=5.95 $Y2=1.99
cc_89 VPB N_VPWR_c_532_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_533_n 0.00503453f $X=-0.19 $Y=1.305 $X2=6.565 $Y2=0.72
cc_91 VPB N_VPWR_c_534_n 0.0106906f $X=-0.19 $Y=1.305 $X2=6.445 $Y2=1.995
cc_92 VPB N_VPWR_c_535_n 0.00538776f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=1.202
cc_93 VPB N_VPWR_c_536_n 0.00547281f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_X_c_653_n 0.00716948f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=1.58
cc_95 VPB X 0.00907734f $X=-0.19 $Y=1.305 $X2=5.01 $Y2=0.72
cc_96 VPB N_A_493_297#_c_721_n 0.00782002f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_97 VPB N_A_493_297#_c_722_n 0.00747984f $X=-0.19 $Y=1.305 $X2=2.06 $Y2=1.325
cc_98 VPB N_A_493_297#_c_723_n 0.0195224f $X=-0.19 $Y=1.305 $X2=5.78 $Y2=1.58
cc_99 N_A_79_21#_c_102_n N_A3_c_278_n 0.0227756f $X=1.93 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_100 N_A_79_21#_c_111_n N_A3_c_282_n 0.0226992f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_79_21#_c_113_n N_A3_c_282_n 0.00197721f $X=2.06 $Y=1.495 $X2=0 $Y2=0
cc_102 N_A_79_21#_c_114_n N_A3_c_282_n 0.0207272f $X=5.78 $Y=1.58 $X2=0 $Y2=0
cc_103 N_A_79_21#_c_114_n N_A3_c_283_n 0.0146912f $X=5.78 $Y=1.58 $X2=0 $Y2=0
cc_104 N_A_79_21#_c_103_n A3 0.0149831f $X=1.95 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_79_21#_c_114_n A3 0.0579332f $X=5.78 $Y=1.58 $X2=0 $Y2=0
cc_106 N_A_79_21#_c_103_n N_A3_c_281_n 0.00568189f $X=1.95 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_79_21#_c_113_n N_A3_c_281_n 0.00199272f $X=2.06 $Y=1.495 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_114_n N_A3_c_281_n 0.0114806f $X=5.78 $Y=1.58 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_107_n N_A3_c_281_n 0.0227756f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_114_n N_A2_c_332_n 0.0144732f $X=5.78 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_111 N_A_79_21#_c_114_n N_A2_c_333_n 0.0124303f $X=5.78 $Y=1.58 $X2=0 $Y2=0
cc_112 N_A_79_21#_c_104_n N_A2_c_329_n 5.39901e-19 $X=5.78 $Y=0.72 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_114_n A2 0.0495996f $X=5.78 $Y=1.58 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_114_n N_A2_c_331_n 0.00709873f $X=5.78 $Y=1.58 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_104_n N_A1_M1016_g 0.00400249f $X=5.78 $Y=0.72 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_114_n N_A1_c_378_n 0.0124303f $X=5.78 $Y=1.58 $X2=0 $Y2=0
cc_117 N_A_79_21#_c_104_n N_A1_M1026_g 0.0110355f $X=5.78 $Y=0.72 $X2=0 $Y2=0
cc_118 N_A_79_21#_c_105_n N_A1_M1026_g 0.00515269f $X=5.865 $Y=1.495 $X2=0 $Y2=0
cc_119 N_A_79_21#_c_114_n N_A1_c_379_n 0.0143307f $X=5.78 $Y=1.58 $X2=0 $Y2=0
cc_120 N_A_79_21#_c_105_n N_A1_c_379_n 0.00219725f $X=5.865 $Y=1.495 $X2=0 $Y2=0
cc_121 N_A_79_21#_c_139_p N_A1_c_379_n 0.0062519f $X=5.865 $Y=1.905 $X2=0 $Y2=0
cc_122 N_A_79_21#_c_140_p N_A1_c_379_n 0.00109482f $X=5.95 $Y=1.99 $X2=0 $Y2=0
cc_123 N_A_79_21#_c_114_n N_A1_c_376_n 0.00792324f $X=5.78 $Y=1.58 $X2=0 $Y2=0
cc_124 N_A_79_21#_c_104_n N_A1_c_376_n 0.00923254f $X=5.78 $Y=0.72 $X2=0 $Y2=0
cc_125 N_A_79_21#_c_105_n N_A1_c_376_n 0.00492333f $X=5.865 $Y=1.495 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_114_n A1 0.0583325f $X=5.78 $Y=1.58 $X2=0 $Y2=0
cc_127 N_A_79_21#_c_104_n A1 0.034631f $X=5.78 $Y=0.72 $X2=0 $Y2=0
cc_128 N_A_79_21#_c_105_n A1 0.0172865f $X=5.865 $Y=1.495 $X2=0 $Y2=0
cc_129 N_A_79_21#_c_105_n N_B1_M1007_g 0.00625781f $X=5.865 $Y=1.495 $X2=0 $Y2=0
cc_130 N_A_79_21#_c_106_n N_B1_M1007_g 0.0110355f $X=6.565 $Y=0.72 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_105_n N_B1_c_426_n 4.01068e-19 $X=5.865 $Y=1.495 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_139_p N_B1_c_426_n 0.00700796f $X=5.865 $Y=1.905 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_151_p N_B1_c_426_n 0.00213503f $X=5.865 $Y=1.58 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_152_p N_B1_c_426_n 0.0113702f $X=6.445 $Y=1.995 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_153_p N_B1_c_426_n 0.00132495f $X=6.51 $Y=1.995 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_154_p N_B1_c_427_n 0.0105478f $X=7.55 $Y=2 $X2=0 $Y2=0
cc_137 N_A_79_21#_M1000_d B1 0.00248603f $X=6.465 $Y=1.485 $X2=0 $Y2=0
cc_138 N_A_79_21#_c_105_n B1 0.0353181f $X=5.865 $Y=1.495 $X2=0 $Y2=0
cc_139 N_A_79_21#_c_154_p B1 0.0261351f $X=7.55 $Y=2 $X2=0 $Y2=0
cc_140 N_A_79_21#_c_106_n B1 0.0289638f $X=6.565 $Y=0.72 $X2=0 $Y2=0
cc_141 N_A_79_21#_c_151_p B1 0.0116308f $X=5.865 $Y=1.58 $X2=0 $Y2=0
cc_142 N_A_79_21#_c_152_p B1 0.0149085f $X=6.445 $Y=1.995 $X2=0 $Y2=0
cc_143 N_A_79_21#_c_105_n N_B1_c_425_n 0.00253732f $X=5.865 $Y=1.495 $X2=0 $Y2=0
cc_144 N_A_79_21#_c_154_p N_B1_c_425_n 7.53851e-19 $X=7.55 $Y=2 $X2=0 $Y2=0
cc_145 N_A_79_21#_c_106_n N_B1_c_425_n 0.00512589f $X=6.565 $Y=0.72 $X2=0 $Y2=0
cc_146 N_A_79_21#_c_152_p N_B1_c_425_n 2.74349e-19 $X=6.445 $Y=1.995 $X2=0 $Y2=0
cc_147 N_A_79_21#_c_154_p N_B2_c_480_n 0.0151952f $X=7.55 $Y=2 $X2=0 $Y2=0
cc_148 N_A_79_21#_c_154_p N_B2_c_481_n 0.00286533f $X=7.55 $Y=2 $X2=0 $Y2=0
cc_149 N_A_79_21#_c_154_p N_B2_c_477_n 0.00147402f $X=7.55 $Y=2 $X2=0 $Y2=0
cc_150 N_A_79_21#_M1009_s B2 0.00530013f $X=7.405 $Y=1.485 $X2=0 $Y2=0
cc_151 N_A_79_21#_c_154_p B2 0.00952506f $X=7.55 $Y=2 $X2=0 $Y2=0
cc_152 N_A_79_21#_c_154_p B2 0.00121372f $X=7.55 $Y=2 $X2=0 $Y2=0
cc_153 N_A_79_21#_c_114_n N_VPWR_M1024_d 0.00289491f $X=5.78 $Y=1.58 $X2=0 $Y2=0
cc_154 N_A_79_21#_c_172_p N_VPWR_M1024_d 0.0015405f $X=2.17 $Y=1.58 $X2=0 $Y2=0
cc_155 N_A_79_21#_c_114_n N_VPWR_M1010_d 0.00550381f $X=5.78 $Y=1.58 $X2=0 $Y2=0
cc_156 N_A_79_21#_c_114_n N_VPWR_M1019_s 0.00369099f $X=5.78 $Y=1.58 $X2=0 $Y2=0
cc_157 N_A_79_21#_c_114_n N_VPWR_M1003_s 0.00369099f $X=5.78 $Y=1.58 $X2=0 $Y2=0
cc_158 N_A_79_21#_c_108_n N_VPWR_c_522_n 0.0118533f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_79_21#_c_109_n N_VPWR_c_522_n 5.94114e-19 $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_160 N_A_79_21#_c_108_n N_VPWR_c_523_n 6.33692e-19 $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_161 N_A_79_21#_c_109_n N_VPWR_c_523_n 0.0144185f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_79_21#_c_110_n N_VPWR_c_523_n 0.0108266f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A_79_21#_c_111_n N_VPWR_c_523_n 5.96427e-19 $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_164 N_A_79_21#_c_110_n N_VPWR_c_524_n 6.33692e-19 $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_165 N_A_79_21#_c_111_n N_VPWR_c_524_n 0.0146295f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_79_21#_c_103_n N_VPWR_c_524_n 6.69973e-19 $X=1.95 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_79_21#_c_114_n N_VPWR_c_524_n 0.0045497f $X=5.78 $Y=1.58 $X2=0 $Y2=0
cc_168 N_A_79_21#_c_172_p N_VPWR_c_524_n 0.0106663f $X=2.17 $Y=1.58 $X2=0 $Y2=0
cc_169 N_A_79_21#_c_108_n N_VPWR_c_527_n 0.00622633f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_170 N_A_79_21#_c_109_n N_VPWR_c_527_n 0.00427505f $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_171 N_A_79_21#_c_110_n N_VPWR_c_528_n 0.00622633f $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_172 N_A_79_21#_c_111_n N_VPWR_c_528_n 0.00427505f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_173 N_A_79_21#_M1000_d N_VPWR_c_520_n 0.00235479f $X=6.465 $Y=1.485 $X2=0
+ $Y2=0
cc_174 N_A_79_21#_M1009_s N_VPWR_c_520_n 0.00235479f $X=7.405 $Y=1.485 $X2=0
+ $Y2=0
cc_175 N_A_79_21#_c_108_n N_VPWR_c_520_n 0.0104011f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A_79_21#_c_109_n N_VPWR_c_520_n 0.00732977f $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_177 N_A_79_21#_c_110_n N_VPWR_c_520_n 0.0104011f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A_79_21#_c_111_n N_VPWR_c_520_n 0.00732977f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_179 N_A_79_21#_c_99_n N_X_c_655_n 0.0176817f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_79_21#_c_103_n N_X_c_655_n 0.00166061f $X=1.95 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A_79_21#_c_107_n N_X_c_655_n 2.18975e-19 $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_182 N_A_79_21#_c_108_n N_X_c_658_n 0.0236575f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A_79_21#_c_99_n N_X_c_659_n 0.00391984f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_79_21#_c_108_n N_X_c_660_n 0.00722591f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A_79_21#_c_109_n N_X_c_660_n 0.00682765f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_186 N_A_79_21#_c_100_n N_X_c_662_n 0.0121659f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_79_21#_c_101_n N_X_c_662_n 0.011914f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_79_21#_c_102_n N_X_c_662_n 0.00527111f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_79_21#_c_103_n N_X_c_662_n 0.0566884f $X=1.95 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_79_21#_c_107_n N_X_c_662_n 0.0072055f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_191 N_A_79_21#_c_109_n N_X_c_667_n 0.0154704f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_192 N_A_79_21#_c_110_n N_X_c_667_n 0.0163986f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A_79_21#_c_111_n N_X_c_667_n 0.00149571f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A_79_21#_c_103_n N_X_c_667_n 0.0615229f $X=1.95 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A_79_21#_c_172_p N_X_c_667_n 0.0133517f $X=2.17 $Y=1.58 $X2=0 $Y2=0
cc_196 N_A_79_21#_c_107_n N_X_c_667_n 0.0103198f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_197 N_A_79_21#_c_101_n N_X_c_673_n 0.00393134f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A_79_21#_c_102_n N_X_c_673_n 0.00379089f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_79_21#_c_110_n N_X_c_675_n 0.00722591f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_200 N_A_79_21#_c_111_n N_X_c_675_n 0.00682765f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A_79_21#_c_103_n N_X_c_677_n 0.0123849f $X=1.95 $Y=1.16 $X2=0 $Y2=0
cc_202 N_A_79_21#_c_107_n N_X_c_677_n 0.00297321f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_203 N_A_79_21#_c_103_n N_X_c_679_n 0.0140387f $X=1.95 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A_79_21#_c_107_n N_X_c_679_n 0.00411803f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_205 N_A_79_21#_c_99_n X 0.0199963f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A_79_21#_c_108_n X 0.00339212f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A_79_21#_c_103_n X 0.0183389f $X=1.95 $Y=1.16 $X2=0 $Y2=0
cc_208 N_A_79_21#_c_114_n N_A_493_297#_M1005_s 0.00366194f $X=5.78 $Y=1.58
+ $X2=-0.19 $Y2=-0.24
cc_209 N_A_79_21#_c_114_n N_A_493_297#_M1019_d 0.0073112f $X=5.78 $Y=1.58 $X2=0
+ $Y2=0
cc_210 N_A_79_21#_c_114_n N_A_493_297#_M1027_d 0.00886286f $X=5.78 $Y=1.58 $X2=0
+ $Y2=0
cc_211 N_A_79_21#_c_114_n N_A_493_297#_M1012_d 0.0181463f $X=5.78 $Y=1.58 $X2=0
+ $Y2=0
cc_212 N_A_79_21#_c_105_n N_A_493_297#_M1012_d 2.95804e-19 $X=5.865 $Y=1.495
+ $X2=0 $Y2=0
cc_213 N_A_79_21#_c_139_p N_A_493_297#_M1012_d 0.00886206f $X=5.865 $Y=1.905
+ $X2=0 $Y2=0
cc_214 N_A_79_21#_c_140_p N_A_493_297#_M1012_d 0.00530018f $X=5.95 $Y=1.99 $X2=0
+ $Y2=0
cc_215 N_A_79_21#_c_151_p N_A_493_297#_M1012_d 0.0034373f $X=5.865 $Y=1.58 $X2=0
+ $Y2=0
cc_216 N_A_79_21#_c_152_p N_A_493_297#_M1012_d 0.0121667f $X=6.445 $Y=1.995
+ $X2=0 $Y2=0
cc_217 N_A_79_21#_c_154_p N_A_493_297#_M1021_s 0.00488593f $X=7.55 $Y=2 $X2=0
+ $Y2=0
cc_218 N_A_79_21#_c_114_n N_A_493_297#_c_721_n 0.0383908f $X=5.78 $Y=1.58 $X2=0
+ $Y2=0
cc_219 N_A_79_21#_c_114_n N_A_493_297#_c_735_n 0.0102182f $X=5.78 $Y=1.58 $X2=0
+ $Y2=0
cc_220 N_A_79_21#_c_114_n N_A_493_297#_c_736_n 0.0277152f $X=5.78 $Y=1.58 $X2=0
+ $Y2=0
cc_221 N_A_79_21#_c_114_n N_A_493_297#_c_737_n 0.0378695f $X=5.78 $Y=1.58 $X2=0
+ $Y2=0
cc_222 N_A_79_21#_c_140_p N_A_493_297#_c_737_n 0.0121023f $X=5.95 $Y=1.99 $X2=0
+ $Y2=0
cc_223 N_A_79_21#_M1000_d N_A_493_297#_c_739_n 0.00367601f $X=6.465 $Y=1.485
+ $X2=0 $Y2=0
cc_224 N_A_79_21#_M1009_s N_A_493_297#_c_739_n 0.00359247f $X=7.405 $Y=1.485
+ $X2=0 $Y2=0
cc_225 N_A_79_21#_c_114_n N_A_493_297#_c_739_n 0.00613779f $X=5.78 $Y=1.58 $X2=0
+ $Y2=0
cc_226 N_A_79_21#_c_140_p N_A_493_297#_c_739_n 0.0123638f $X=5.95 $Y=1.99 $X2=0
+ $Y2=0
cc_227 N_A_79_21#_c_152_p N_A_493_297#_c_739_n 0.0279546f $X=6.445 $Y=1.995
+ $X2=0 $Y2=0
cc_228 N_A_79_21#_c_153_p N_A_493_297#_c_739_n 0.0619396f $X=6.51 $Y=1.995 $X2=0
+ $Y2=0
cc_229 N_A_79_21#_c_154_p N_A_493_297#_c_723_n 0.0111115f $X=7.55 $Y=2 $X2=0
+ $Y2=0
cc_230 N_A_79_21#_c_114_n N_A_493_297#_c_746_n 0.0102182f $X=5.78 $Y=1.58 $X2=0
+ $Y2=0
cc_231 N_A_79_21#_c_114_n N_A_493_297#_c_747_n 0.0102182f $X=5.78 $Y=1.58 $X2=0
+ $Y2=0
cc_232 N_A_79_21#_c_99_n N_VGND_c_813_n 0.00812954f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_79_21#_c_100_n N_VGND_c_813_n 5.10336e-19 $X=0.94 $Y=0.995 $X2=0
+ $Y2=0
cc_234 N_A_79_21#_c_99_n N_VGND_c_814_n 0.00339367f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A_79_21#_c_100_n N_VGND_c_814_n 0.00340075f $X=0.94 $Y=0.995 $X2=0
+ $Y2=0
cc_236 N_A_79_21#_c_101_n N_VGND_c_815_n 0.00340075f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_237 N_A_79_21#_c_102_n N_VGND_c_815_n 0.00273179f $X=1.93 $Y=0.995 $X2=0
+ $Y2=0
cc_238 N_A_79_21#_c_104_n N_VGND_c_817_n 0.00520015f $X=5.78 $Y=0.72 $X2=0 $Y2=0
cc_239 N_A_79_21#_M1016_s N_VGND_c_819_n 0.00259839f $X=4.825 $Y=0.235 $X2=0
+ $Y2=0
cc_240 N_A_79_21#_M1007_s N_VGND_c_819_n 0.00259839f $X=6.43 $Y=0.235 $X2=0
+ $Y2=0
cc_241 N_A_79_21#_c_99_n N_VGND_c_819_n 0.00407103f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_79_21#_c_100_n N_VGND_c_819_n 0.00407108f $X=0.94 $Y=0.995 $X2=0
+ $Y2=0
cc_243 N_A_79_21#_c_101_n N_VGND_c_819_n 0.00418642f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_244 N_A_79_21#_c_102_n N_VGND_c_819_n 0.00513576f $X=1.93 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_A_79_21#_c_104_n N_VGND_c_819_n 0.0111591f $X=5.78 $Y=0.72 $X2=0 $Y2=0
cc_246 N_A_79_21#_c_99_n N_VGND_c_820_n 4.98468e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A_79_21#_c_100_n N_VGND_c_820_n 0.00701096f $X=0.94 $Y=0.995 $X2=0
+ $Y2=0
cc_248 N_A_79_21#_c_101_n N_VGND_c_820_n 0.00727879f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_249 N_A_79_21#_c_102_n N_VGND_c_820_n 4.78403e-19 $X=1.93 $Y=0.995 $X2=0
+ $Y2=0
cc_250 N_A_79_21#_c_101_n N_VGND_c_821_n 5.25757e-19 $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_251 N_A_79_21#_c_102_n N_VGND_c_821_n 0.010602f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A_79_21#_c_103_n N_VGND_c_821_n 0.00800756f $X=1.95 $Y=1.16 $X2=0 $Y2=0
cc_253 N_A_79_21#_c_114_n N_A_485_47#_c_925_n 0.00615854f $X=5.78 $Y=1.58 $X2=0
+ $Y2=0
cc_254 N_A_79_21#_c_104_n N_A_695_47#_M1026_d 0.00722815f $X=5.78 $Y=0.72 $X2=0
+ $Y2=0
cc_255 N_A_79_21#_M1016_s N_A_695_47#_c_950_n 0.00416045f $X=4.825 $Y=0.235
+ $X2=0 $Y2=0
cc_256 N_A_79_21#_c_104_n N_A_695_47#_c_950_n 0.0459803f $X=5.78 $Y=0.72 $X2=0
+ $Y2=0
cc_257 N_A_79_21#_c_106_n N_A_1194_47#_M1007_d 0.010741f $X=6.565 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_258 N_A_79_21#_M1007_s N_A_1194_47#_c_970_n 0.00416045f $X=6.43 $Y=0.235
+ $X2=0 $Y2=0
cc_259 N_A_79_21#_c_106_n N_A_1194_47#_c_970_n 0.0440811f $X=6.565 $Y=0.72 $X2=0
+ $Y2=0
cc_260 A3 A2 0.0154732f $X=2.915 $Y=1.105 $X2=0 $Y2=0
cc_261 N_A3_c_281_n A2 0.00100405f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_262 A3 N_A2_c_331_n 0.0010265f $X=2.915 $Y=1.105 $X2=0 $Y2=0
cc_263 N_A3_c_281_n N_A2_c_331_n 0.00764048f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_264 N_A3_c_282_n N_VPWR_c_524_n 0.0107697f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A3_c_283_n N_VPWR_c_524_n 6.67754e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A3_c_282_n N_VPWR_c_529_n 0.00622633f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_267 N_A3_c_283_n N_VPWR_c_529_n 0.00311736f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A3_c_282_n N_VPWR_c_520_n 0.0104011f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A3_c_283_n N_VPWR_c_520_n 0.00371107f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_270 N_A3_c_282_n N_VPWR_c_534_n 5.36535e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_271 N_A3_c_283_n N_VPWR_c_534_n 0.0104595f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_272 N_A3_c_282_n N_A_493_297#_c_748_n 0.00140601f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_273 N_A3_c_283_n N_A_493_297#_c_748_n 0.00397069f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_274 N_A3_c_283_n N_A_493_297#_c_721_n 0.0149699f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_275 N_A3_c_282_n N_A_493_297#_c_735_n 0.00158423f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_276 N_A3_c_283_n N_A_493_297#_c_752_n 0.00260293f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_277 N_A3_c_278_n N_VGND_c_816_n 0.00468308f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A3_c_279_n N_VGND_c_816_n 0.00342417f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A3_c_278_n N_VGND_c_819_n 0.00801881f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_280 N_A3_c_279_n N_VGND_c_819_n 0.00410992f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_281 N_A3_c_278_n N_VGND_c_821_n 0.00801067f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_282 N_A3_c_279_n N_VGND_c_821_n 5.13099e-19 $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_283 N_A3_c_278_n N_VGND_c_822_n 4.98468e-19 $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_284 N_A3_c_279_n N_VGND_c_822_n 0.00800318f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_285 N_A3_c_278_n N_A_485_47#_c_927_n 0.00438037f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_286 N_A3_c_278_n N_A_485_47#_c_928_n 0.00517315f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_287 A3 N_A_485_47#_c_928_n 0.00977463f $X=2.915 $Y=1.105 $X2=0 $Y2=0
cc_288 N_A3_c_281_n N_A_485_47#_c_928_n 0.00316718f $X=2.845 $Y=1.202 $X2=0
+ $Y2=0
cc_289 N_A3_c_279_n N_A_485_47#_c_925_n 0.0138319f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_290 A3 N_A_485_47#_c_925_n 0.0357061f $X=2.915 $Y=1.105 $X2=0 $Y2=0
cc_291 N_A3_c_281_n N_A_485_47#_c_925_n 0.00649437f $X=2.845 $Y=1.202 $X2=0
+ $Y2=0
cc_292 N_A2_c_329_n N_A1_M1016_g 0.0246742f $X=4.33 $Y=0.995 $X2=0 $Y2=0
cc_293 N_A2_c_333_n N_A1_c_378_n 0.0386055f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_294 A2 N_A1_c_376_n 0.00192062f $X=4.035 $Y=1.105 $X2=0 $Y2=0
cc_295 N_A2_c_331_n N_A1_c_376_n 0.0246742f $X=4.305 $Y=1.202 $X2=0 $Y2=0
cc_296 A2 A1 0.0165393f $X=4.035 $Y=1.105 $X2=0 $Y2=0
cc_297 N_A2_c_331_n A1 2.9754e-19 $X=4.305 $Y=1.202 $X2=0 $Y2=0
cc_298 N_A2_c_332_n N_VPWR_c_525_n 0.00311736f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_299 N_A2_c_333_n N_VPWR_c_526_n 0.00453434f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_300 N_A2_c_332_n N_VPWR_c_520_n 0.00499342f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_301 N_A2_c_333_n N_VPWR_c_520_n 0.00516277f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_302 N_A2_c_332_n N_VPWR_c_534_n 0.00187777f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_303 N_A2_c_332_n N_VPWR_c_535_n 0.00969468f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_304 N_A2_c_333_n N_VPWR_c_535_n 0.0067928f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_305 N_A2_c_333_n N_VPWR_c_536_n 5.36535e-19 $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_306 N_A2_c_332_n N_A_493_297#_c_752_n 0.0042783f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_307 N_A2_c_332_n N_A_493_297#_c_736_n 0.0154573f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_308 N_A2_c_333_n N_A_493_297#_c_736_n 0.013884f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_309 N_A2_c_333_n N_A_493_297#_c_756_n 0.00412276f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_310 N_A2_c_328_n N_VGND_c_817_n 0.00366111f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_311 N_A2_c_329_n N_VGND_c_817_n 0.00366111f $X=4.33 $Y=0.995 $X2=0 $Y2=0
cc_312 N_A2_c_328_n N_VGND_c_819_n 0.00669801f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_313 N_A2_c_329_n N_VGND_c_819_n 0.00539914f $X=4.33 $Y=0.995 $X2=0 $Y2=0
cc_314 N_A2_c_328_n N_VGND_c_822_n 0.00276567f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_315 N_A2_c_328_n N_A_485_47#_c_925_n 0.0110467f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_316 A2 N_A_485_47#_c_925_n 0.027736f $X=4.035 $Y=1.105 $X2=0 $Y2=0
cc_317 N_A2_c_331_n N_A_485_47#_c_925_n 0.00658933f $X=4.305 $Y=1.202 $X2=0
+ $Y2=0
cc_318 N_A2_c_328_n N_A_695_47#_c_950_n 0.00830874f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_319 N_A2_c_329_n N_A_695_47#_c_950_n 0.0102498f $X=4.33 $Y=0.995 $X2=0 $Y2=0
cc_320 A2 N_A_695_47#_c_950_n 0.00428441f $X=4.035 $Y=1.105 $X2=0 $Y2=0
cc_321 N_A1_c_376_n N_B1_c_425_n 0.0038527f $X=5.245 $Y=1.212 $X2=0 $Y2=0
cc_322 N_A1_c_378_n N_VPWR_c_526_n 0.00311736f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_323 N_A1_c_379_n N_VPWR_c_530_n 0.00453434f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_324 N_A1_c_378_n N_VPWR_c_520_n 0.00373628f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_325 N_A1_c_379_n N_VPWR_c_520_n 0.0065142f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_326 N_A1_c_378_n N_VPWR_c_535_n 4.88209e-19 $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_327 N_A1_c_378_n N_VPWR_c_536_n 0.00943288f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_328 N_A1_c_379_n N_VPWR_c_536_n 0.00962799f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_329 N_A1_c_378_n N_A_493_297#_c_756_n 0.00397069f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_330 N_A1_c_378_n N_A_493_297#_c_737_n 0.0133714f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_331 N_A1_c_379_n N_A_493_297#_c_737_n 0.0150429f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_332 N_A1_c_379_n N_A_493_297#_c_760_n 0.00666024f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_333 N_A1_c_379_n N_A_493_297#_c_761_n 0.00420108f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_334 N_A1_M1016_g N_VGND_c_817_n 0.00366111f $X=4.75 $Y=0.56 $X2=0 $Y2=0
cc_335 N_A1_M1026_g N_VGND_c_817_n 0.00366111f $X=5.22 $Y=0.56 $X2=0 $Y2=0
cc_336 N_A1_M1016_g N_VGND_c_819_n 0.00539914f $X=4.75 $Y=0.56 $X2=0 $Y2=0
cc_337 N_A1_M1026_g N_VGND_c_819_n 0.00669801f $X=5.22 $Y=0.56 $X2=0 $Y2=0
cc_338 N_A1_M1016_g N_A_695_47#_c_950_n 0.00972451f $X=4.75 $Y=0.56 $X2=0 $Y2=0
cc_339 N_A1_M1026_g N_A_695_47#_c_950_n 0.00818766f $X=5.22 $Y=0.56 $X2=0 $Y2=0
cc_340 A1 N_A_695_47#_c_950_n 0.00278778f $X=5.345 $Y=1.19 $X2=0 $Y2=0
cc_341 N_B1_M1017_g N_B2_M1011_g 0.0219891f $X=6.825 $Y=0.56 $X2=0 $Y2=0
cc_342 N_B1_c_427_n N_B2_c_480_n 0.0396375f $X=6.845 $Y=1.41 $X2=0 $Y2=0
cc_343 B1 N_B2_c_480_n 0.00220155f $X=6.965 $Y=1.105 $X2=0 $Y2=0
cc_344 B1 N_B2_c_477_n 0.00380573f $X=6.965 $Y=1.105 $X2=0 $Y2=0
cc_345 N_B1_c_425_n N_B2_c_477_n 0.0188298f $X=6.825 $Y=1.217 $X2=0 $Y2=0
cc_346 B1 B2 0.01481f $X=6.965 $Y=1.105 $X2=0 $Y2=0
cc_347 B1 N_B2_c_497_n 0.0127375f $X=6.965 $Y=1.105 $X2=0 $Y2=0
cc_348 N_B1_c_426_n N_VPWR_c_530_n 0.00439333f $X=6.375 $Y=1.41 $X2=0 $Y2=0
cc_349 N_B1_c_427_n N_VPWR_c_530_n 0.00439333f $X=6.845 $Y=1.41 $X2=0 $Y2=0
cc_350 N_B1_c_426_n N_VPWR_c_520_n 0.00736527f $X=6.375 $Y=1.41 $X2=0 $Y2=0
cc_351 N_B1_c_427_n N_VPWR_c_520_n 0.00610813f $X=6.845 $Y=1.41 $X2=0 $Y2=0
cc_352 B1 N_A_493_297#_M1012_d 0.00303759f $X=6.965 $Y=1.105 $X2=0 $Y2=0
cc_353 B1 N_A_493_297#_M1021_s 0.00371694f $X=6.965 $Y=1.105 $X2=0 $Y2=0
cc_354 N_B1_c_426_n N_A_493_297#_c_739_n 0.00927722f $X=6.375 $Y=1.41 $X2=0
+ $Y2=0
cc_355 N_B1_c_427_n N_A_493_297#_c_739_n 0.0092122f $X=6.845 $Y=1.41 $X2=0 $Y2=0
cc_356 N_B1_M1007_g N_VGND_c_817_n 0.00366111f $X=6.355 $Y=0.56 $X2=0 $Y2=0
cc_357 N_B1_M1017_g N_VGND_c_817_n 0.00366111f $X=6.825 $Y=0.56 $X2=0 $Y2=0
cc_358 N_B1_M1007_g N_VGND_c_819_n 0.00669801f $X=6.355 $Y=0.56 $X2=0 $Y2=0
cc_359 N_B1_M1017_g N_VGND_c_819_n 0.00550601f $X=6.825 $Y=0.56 $X2=0 $Y2=0
cc_360 N_B1_M1017_g N_VGND_c_823_n 0.00105522f $X=6.825 $Y=0.56 $X2=0 $Y2=0
cc_361 N_B1_M1007_g N_A_1194_47#_c_970_n 0.00818766f $X=6.355 $Y=0.56 $X2=0
+ $Y2=0
cc_362 N_B1_M1017_g N_A_1194_47#_c_970_n 0.0102498f $X=6.825 $Y=0.56 $X2=0 $Y2=0
cc_363 B1 N_A_1194_47#_c_970_n 0.00615043f $X=6.965 $Y=1.105 $X2=0 $Y2=0
cc_364 N_B1_M1017_g N_A_1194_47#_c_977_n 0.00335708f $X=6.825 $Y=0.56 $X2=0
+ $Y2=0
cc_365 N_B1_M1017_g N_A_1194_47#_c_978_n 0.00184846f $X=6.825 $Y=0.56 $X2=0
+ $Y2=0
cc_366 B1 N_A_1194_47#_c_978_n 0.00948197f $X=6.965 $Y=1.105 $X2=0 $Y2=0
cc_367 N_B2_c_480_n N_VPWR_c_530_n 0.00439333f $X=7.315 $Y=1.41 $X2=0 $Y2=0
cc_368 N_B2_c_481_n N_VPWR_c_530_n 0.00439333f $X=7.785 $Y=1.41 $X2=0 $Y2=0
cc_369 N_B2_c_480_n N_VPWR_c_520_n 0.00610813f $X=7.315 $Y=1.41 $X2=0 $Y2=0
cc_370 N_B2_c_481_n N_VPWR_c_520_n 0.00699435f $X=7.785 $Y=1.41 $X2=0 $Y2=0
cc_371 N_B2_c_480_n N_A_493_297#_c_739_n 0.0092122f $X=7.315 $Y=1.41 $X2=0 $Y2=0
cc_372 N_B2_c_481_n N_A_493_297#_c_739_n 0.0140683f $X=7.785 $Y=1.41 $X2=0 $Y2=0
cc_373 N_B2_c_481_n N_A_493_297#_c_723_n 0.0083028f $X=7.785 $Y=1.41 $X2=0 $Y2=0
cc_374 B2 N_A_493_297#_c_723_n 0.00874362f $X=7.96 $Y=1.105 $X2=0 $Y2=0
cc_375 N_B2_c_479_n N_A_493_297#_c_723_n 0.00442545f $X=8.005 $Y=1.16 $X2=0
+ $Y2=0
cc_376 N_B2_M1011_g N_VGND_c_817_n 0.00341252f $X=7.29 $Y=0.56 $X2=0 $Y2=0
cc_377 N_B2_M1014_g N_VGND_c_818_n 0.00341252f $X=7.76 $Y=0.56 $X2=0 $Y2=0
cc_378 N_B2_M1011_g N_VGND_c_819_n 0.00409755f $X=7.29 $Y=0.56 $X2=0 $Y2=0
cc_379 N_B2_M1014_g N_VGND_c_819_n 0.00496234f $X=7.76 $Y=0.56 $X2=0 $Y2=0
cc_380 N_B2_M1011_g N_VGND_c_823_n 0.00810717f $X=7.29 $Y=0.56 $X2=0 $Y2=0
cc_381 N_B2_M1014_g N_VGND_c_823_n 0.00887115f $X=7.76 $Y=0.56 $X2=0 $Y2=0
cc_382 N_B2_M1011_g N_A_1194_47#_c_980_n 0.0160546f $X=7.29 $Y=0.56 $X2=0 $Y2=0
cc_383 N_B2_M1014_g N_A_1194_47#_c_980_n 0.0136203f $X=7.76 $Y=0.56 $X2=0 $Y2=0
cc_384 N_B2_c_477_n N_A_1194_47#_c_980_n 0.00523729f $X=7.885 $Y=1.165 $X2=0
+ $Y2=0
cc_385 B2 N_A_1194_47#_c_980_n 0.0219147f $X=7.96 $Y=1.105 $X2=0 $Y2=0
cc_386 N_B2_c_479_n N_A_1194_47#_c_980_n 0.00384366f $X=8.005 $Y=1.16 $X2=0
+ $Y2=0
cc_387 N_B2_c_497_n N_A_1194_47#_c_980_n 0.0106783f $X=7.537 $Y=1.295 $X2=0
+ $Y2=0
cc_388 N_B2_M1014_g N_A_1194_47#_c_986_n 0.00456759f $X=7.76 $Y=0.56 $X2=0 $Y2=0
cc_389 N_VPWR_c_520_n N_X_M1002_s 0.00647849f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_390 N_VPWR_c_520_n N_X_M1015_s 0.00647849f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_391 N_VPWR_M1002_d N_X_c_658_n 3.55515e-19 $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_392 N_VPWR_c_522_n N_X_c_658_n 0.00149271f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_393 N_VPWR_c_522_n N_X_c_660_n 0.0332981f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_394 N_VPWR_c_523_n N_X_c_660_n 0.0410603f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_395 N_VPWR_c_527_n N_X_c_660_n 0.0118139f $X=0.985 $Y=2.72 $X2=0 $Y2=0
cc_396 N_VPWR_c_520_n N_X_c_660_n 0.00646998f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_397 N_VPWR_M1008_d N_X_c_667_n 0.00369624f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_398 N_VPWR_c_523_n N_X_c_667_n 0.0156171f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_399 N_VPWR_c_523_n N_X_c_675_n 0.0336646f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_400 N_VPWR_c_524_n N_X_c_675_n 0.0410603f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_401 N_VPWR_c_528_n N_X_c_675_n 0.0118139f $X=1.925 $Y=2.72 $X2=0 $Y2=0
cc_402 N_VPWR_c_520_n N_X_c_675_n 0.00646998f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_403 N_VPWR_M1002_d N_X_c_653_n 0.0035341f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_404 N_VPWR_c_522_n N_X_c_653_n 0.0148711f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_405 N_VPWR_c_520_n N_A_493_297#_M1005_s 0.00460277f $X=8.05 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_406 N_VPWR_c_520_n N_A_493_297#_M1019_d 0.00252028f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_520_n N_A_493_297#_M1027_d 0.00272704f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_520_n N_A_493_297#_M1012_d 0.00801795f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_520_n N_A_493_297#_M1021_s 0.00233855f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_520_n N_A_493_297#_M1013_d 0.00219869f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_524_n N_A_493_297#_c_748_n 0.0232292f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_412 N_VPWR_c_529_n N_A_493_297#_c_748_n 0.0116326f $X=2.865 $Y=2.72 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_520_n N_A_493_297#_c_748_n 0.00643448f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_534_n N_A_493_297#_c_748_n 0.0156776f $X=3.08 $Y=2.34 $X2=0
+ $Y2=0
cc_415 N_VPWR_M1010_d N_A_493_297#_c_721_n 0.00548945f $X=2.935 $Y=1.485 $X2=0
+ $Y2=0
cc_416 N_VPWR_c_525_n N_A_493_297#_c_721_n 0.00489589f $X=3.855 $Y=2.72 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_529_n N_A_493_297#_c_721_n 0.00238709f $X=2.865 $Y=2.72 $X2=0
+ $Y2=0
cc_418 N_VPWR_c_520_n N_A_493_297#_c_721_n 0.0135801f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_419 N_VPWR_c_534_n N_A_493_297#_c_721_n 0.0242262f $X=3.08 $Y=2.34 $X2=0
+ $Y2=0
cc_420 N_VPWR_c_524_n N_A_493_297#_c_735_n 0.0116213f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_421 N_VPWR_c_525_n N_A_493_297#_c_752_n 0.0116326f $X=3.855 $Y=2.72 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_520_n N_A_493_297#_c_752_n 0.00643448f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_423 N_VPWR_c_534_n N_A_493_297#_c_752_n 0.0119006f $X=3.08 $Y=2.34 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_535_n N_A_493_297#_c_752_n 0.0156776f $X=4.07 $Y=2.34 $X2=0
+ $Y2=0
cc_425 N_VPWR_M1019_s N_A_493_297#_c_736_n 0.00379868f $X=3.925 $Y=1.485 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_525_n N_A_493_297#_c_736_n 0.00238709f $X=3.855 $Y=2.72 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_526_n N_A_493_297#_c_736_n 0.00320526f $X=4.795 $Y=2.72 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_520_n N_A_493_297#_c_736_n 0.0112979f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_535_n N_A_493_297#_c_736_n 0.0196308f $X=4.07 $Y=2.34 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_526_n N_A_493_297#_c_756_n 0.0116326f $X=4.795 $Y=2.72 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_520_n N_A_493_297#_c_756_n 0.00643448f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_432 N_VPWR_c_535_n N_A_493_297#_c_756_n 0.0128538f $X=4.07 $Y=2.34 $X2=0
+ $Y2=0
cc_433 N_VPWR_c_536_n N_A_493_297#_c_756_n 0.0156776f $X=5.01 $Y=2.34 $X2=0
+ $Y2=0
cc_434 N_VPWR_M1003_s N_A_493_297#_c_737_n 0.00379868f $X=4.865 $Y=1.485 $X2=0
+ $Y2=0
cc_435 N_VPWR_c_526_n N_A_493_297#_c_737_n 0.00238709f $X=4.795 $Y=2.72 $X2=0
+ $Y2=0
cc_436 N_VPWR_c_530_n N_A_493_297#_c_737_n 0.00320526f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_437 N_VPWR_c_520_n N_A_493_297#_c_737_n 0.0113396f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_438 N_VPWR_c_536_n N_A_493_297#_c_737_n 0.0196308f $X=5.01 $Y=2.34 $X2=0
+ $Y2=0
cc_439 N_VPWR_c_530_n N_A_493_297#_c_739_n 0.108429f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_440 N_VPWR_c_520_n N_A_493_297#_c_739_n 0.0824872f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_441 N_VPWR_c_530_n N_A_493_297#_c_761_n 0.00931009f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_520_n N_A_493_297#_c_761_n 0.00636368f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_443 N_VPWR_c_536_n N_A_493_297#_c_761_n 0.0116213f $X=5.01 $Y=2.34 $X2=0
+ $Y2=0
cc_444 N_VPWR_c_530_n N_A_493_297#_c_722_n 0.0140118f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_445 N_VPWR_c_520_n N_A_493_297#_c_722_n 0.00943351f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_446 N_X_c_651_n N_VGND_M1004_s 0.00291379f $X=0.23 $Y=0.805 $X2=-0.19
+ $Y2=-0.24
cc_447 X N_VGND_M1004_s 3.49814e-19 $X=0.235 $Y=0.85 $X2=-0.19 $Y2=-0.24
cc_448 N_X_c_662_n N_VGND_M1006_s 0.00407492f $X=1.585 $Y=0.72 $X2=0 $Y2=0
cc_449 N_X_c_655_n N_VGND_c_813_n 0.0020301f $X=0.645 $Y=0.72 $X2=0 $Y2=0
cc_450 N_X_c_659_n N_VGND_c_813_n 0.012714f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_451 N_X_c_651_n N_VGND_c_813_n 0.018421f $X=0.23 $Y=0.805 $X2=0 $Y2=0
cc_452 N_X_c_655_n N_VGND_c_814_n 0.00325651f $X=0.645 $Y=0.72 $X2=0 $Y2=0
cc_453 N_X_c_659_n N_VGND_c_814_n 0.01143f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_454 N_X_c_662_n N_VGND_c_814_n 0.00245287f $X=1.585 $Y=0.72 $X2=0 $Y2=0
cc_455 N_X_c_662_n N_VGND_c_815_n 0.0032663f $X=1.585 $Y=0.72 $X2=0 $Y2=0
cc_456 N_X_c_673_n N_VGND_c_815_n 0.0116326f $X=1.67 $Y=0.42 $X2=0 $Y2=0
cc_457 N_X_M1004_d N_VGND_c_819_n 0.00307738f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_458 N_X_M1018_d N_VGND_c_819_n 0.00680678f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_459 N_X_c_655_n N_VGND_c_819_n 0.00598053f $X=0.645 $Y=0.72 $X2=0 $Y2=0
cc_460 N_X_c_659_n N_VGND_c_819_n 0.00643448f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_461 N_X_c_662_n N_VGND_c_819_n 0.011481f $X=1.585 $Y=0.72 $X2=0 $Y2=0
cc_462 N_X_c_673_n N_VGND_c_819_n 0.00643448f $X=1.67 $Y=0.42 $X2=0 $Y2=0
cc_463 N_X_c_651_n N_VGND_c_819_n 0.00110403f $X=0.23 $Y=0.805 $X2=0 $Y2=0
cc_464 N_X_c_662_n N_VGND_c_820_n 0.0197774f $X=1.585 $Y=0.72 $X2=0 $Y2=0
cc_465 N_X_c_673_n N_VGND_c_820_n 0.0128539f $X=1.67 $Y=0.42 $X2=0 $Y2=0
cc_466 N_X_c_673_n N_VGND_c_821_n 0.0156777f $X=1.67 $Y=0.42 $X2=0 $Y2=0
cc_467 N_VGND_c_819_n N_A_485_47#_M1022_s 0.00621001f $X=8.05 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_468 N_VGND_c_819_n N_A_485_47#_M1001_d 0.00259839f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_469 N_VGND_c_816_n N_A_485_47#_c_927_n 0.011459f $X=2.865 $Y=0 $X2=0 $Y2=0
cc_470 N_VGND_c_819_n N_A_485_47#_c_927_n 0.00644035f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_471 N_VGND_c_821_n N_A_485_47#_c_927_n 0.0128539f $X=2.07 $Y=0 $X2=0 $Y2=0
cc_472 N_VGND_M1023_d N_A_485_47#_c_925_n 0.00647497f $X=2.895 $Y=0.235 $X2=0
+ $Y2=0
cc_473 N_VGND_c_816_n N_A_485_47#_c_925_n 0.00233958f $X=2.865 $Y=0 $X2=0 $Y2=0
cc_474 N_VGND_c_817_n N_A_485_47#_c_925_n 0.00332968f $X=7.335 $Y=0 $X2=0 $Y2=0
cc_475 N_VGND_c_819_n N_A_485_47#_c_925_n 0.0127632f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_476 N_VGND_c_822_n N_A_485_47#_c_925_n 0.0222621f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_477 N_VGND_c_819_n N_A_695_47#_M1001_s 0.00253093f $X=8.05 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_478 N_VGND_c_819_n N_A_695_47#_M1020_s 0.00217615f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_479 N_VGND_c_819_n N_A_695_47#_M1026_d 0.00253093f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_480 N_VGND_c_817_n N_A_695_47#_c_950_n 0.100713f $X=7.335 $Y=0 $X2=0 $Y2=0
cc_481 N_VGND_c_819_n N_A_695_47#_c_950_n 0.0772485f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_482 N_VGND_c_822_n N_A_695_47#_c_950_n 0.0138766f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_483 N_VGND_c_819_n N_A_1194_47#_M1007_d 0.00253093f $X=8.05 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_484 N_VGND_c_819_n N_A_1194_47#_M1017_d 0.00270767f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_485 N_VGND_c_819_n N_A_1194_47#_M1014_d 0.00429389f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_486 N_VGND_c_817_n N_A_1194_47#_c_970_n 0.0483121f $X=7.335 $Y=0 $X2=0 $Y2=0
cc_487 N_VGND_c_819_n N_A_1194_47#_c_970_n 0.0371662f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_488 N_VGND_c_817_n N_A_1194_47#_c_992_n 0.0115494f $X=7.335 $Y=0 $X2=0 $Y2=0
cc_489 N_VGND_c_819_n N_A_1194_47#_c_992_n 0.00651407f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_490 N_VGND_M1011_s N_A_1194_47#_c_980_n 0.00487142f $X=7.365 $Y=0.235 $X2=0
+ $Y2=0
cc_491 N_VGND_c_817_n N_A_1194_47#_c_980_n 0.00239531f $X=7.335 $Y=0 $X2=0 $Y2=0
cc_492 N_VGND_c_818_n N_A_1194_47#_c_980_n 0.00319074f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_493 N_VGND_c_819_n N_A_1194_47#_c_980_n 0.0114047f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_494 N_VGND_c_823_n N_A_1194_47#_c_980_n 0.0188453f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_495 N_VGND_c_818_n N_A_1194_47#_c_986_n 0.0116477f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_496 N_VGND_c_819_n N_A_1194_47#_c_986_n 0.00643744f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_497 N_VGND_c_823_n N_A_1194_47#_c_986_n 0.0128539f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_498 N_A_485_47#_c_925_n N_A_695_47#_M1001_s 0.00822572f $X=4.07 $Y=0.74
+ $X2=-0.19 $Y2=-0.24
cc_499 N_A_485_47#_M1001_d N_A_695_47#_c_950_n 0.00424315f $X=3.935 $Y=0.235
+ $X2=0 $Y2=0
cc_500 N_A_485_47#_c_925_n N_A_695_47#_c_950_n 0.0401184f $X=4.07 $Y=0.74 $X2=0
+ $Y2=0
cc_501 N_A_695_47#_c_950_n N_A_1194_47#_c_970_n 0.010958f $X=5.48 $Y=0.38 $X2=0
+ $Y2=0
