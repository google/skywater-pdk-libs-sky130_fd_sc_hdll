* File: sky130_fd_sc_hdll__o211ai_2.spice
* Created: Wed Sep  2 08:42:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o211ai_2.pex.spice"
.subckt sky130_fd_sc_hdll__o211ai_2  VNB VPB C1 B1 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1007 N_A_27_47#_M1007_d N_C1_M1007_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.21775 AS=0.10725 PD=1.97 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.3
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1013 N_A_27_47#_M1013_d N_C1_M1013_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75000.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1000 N_A_316_47#_M1000_d N_B1_M1000_g N_A_27_47#_M1013_d VNB NSHORT L=0.15
+ W=0.65 AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=0 NRS=9.228 M=1 R=4.33333
+ SA=75001.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1002 N_A_316_47#_M1000_d N_B1_M1002_g N_A_27_47#_M1002_s VNB NSHORT L=0.15
+ W=0.65 AD=0.10725 AS=0.18525 PD=0.98 PS=1.87 NRD=9.228 NRS=0 M=1 R=4.33333
+ SA=75001.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_316_47#_M1004_d N_A2_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.115375 AS=0.21775 PD=1.005 PS=1.97 NRD=0 NRS=9.228 M=1 R=4.33333
+ SA=75000.3 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1011 N_A_316_47#_M1004_d N_A2_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.115375 AS=0.099125 PD=1.005 PS=0.955 NRD=13.836 NRS=0 M=1 R=4.33333
+ SA=75000.8 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1009 N_A_316_47#_M1009_d N_A1_M1009_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.108875 AS=0.099125 PD=0.985 PS=0.955 NRD=0 NRS=5.532 M=1 R=4.33333
+ SA=75001.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1010 N_A_316_47#_M1009_d N_A1_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.108875 AS=0.19825 PD=0.985 PS=1.91 NRD=10.152 NRS=3.684 M=1 R=4.33333
+ SA=75001.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_C1_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.275
+ AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1014 N_VPWR_M1014_d N_C1_M1014_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1014_d N_B1_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.1
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1015 N_VPWR_M1015_d N_B1_M1015_g N_Y_M1006_s VPB PHIGHVT L=0.18 W=1 AD=0.275
+ AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1001 N_Y_M1001_d N_A2_M1001_g N_A_527_297#_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1008 N_Y_M1001_d N_A2_M1008_g N_A_527_297#_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g N_A_527_297#_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.1
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1005_d N_A1_M1012_g N_A_527_297#_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.7312 P=14.09
*
.include "sky130_fd_sc_hdll__o211ai_2.pxi.spice"
*
.ends
*
*
