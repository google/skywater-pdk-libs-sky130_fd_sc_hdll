* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__dlxtn_4 D GATE_N VGND VNB VPB VPWR Q
X0 a_609_413# a_27_47# a_703_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X1 a_774_21# a_609_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_609_413# a_211_363# a_709_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X3 a_27_47# GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X4 a_709_47# a_774_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_319_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR a_774_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 a_503_369# a_211_363# a_609_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X8 VGND a_27_47# a_211_363# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND a_774_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND a_774_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_774_21# a_609_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 Q a_774_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 VPWR a_319_47# a_503_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X14 a_27_47# GATE_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VPWR a_774_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 VPWR a_27_47# a_211_363# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X17 Q a_774_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_505_47# a_27_47# a_609_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X19 a_319_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X20 a_703_413# a_774_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X21 VGND a_319_47# a_505_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 Q a_774_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 Q a_774_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
