* File: sky130_fd_sc_hdll__dlxtn_4.pxi.spice
* Created: Wed Sep  2 08:30:08 2020
* 
x_PM_SKY130_FD_SC_HDLL__DLXTN_4%GATE_N N_GATE_N_c_142_n N_GATE_N_c_143_n
+ N_GATE_N_M1004_g N_GATE_N_c_137_n N_GATE_N_M1016_g N_GATE_N_c_138_n GATE_N
+ GATE_N N_GATE_N_c_140_n N_GATE_N_c_141_n PM_SKY130_FD_SC_HDLL__DLXTN_4%GATE_N
x_PM_SKY130_FD_SC_HDLL__DLXTN_4%A_27_47# N_A_27_47#_M1016_s N_A_27_47#_M1004_s
+ N_A_27_47#_c_187_n N_A_27_47#_c_188_n N_A_27_47#_M1019_g N_A_27_47#_M1001_g
+ N_A_27_47#_M1008_g N_A_27_47#_c_189_n N_A_27_47#_M1015_g N_A_27_47#_c_316_p
+ N_A_27_47#_c_179_n N_A_27_47#_c_180_n N_A_27_47#_c_190_n N_A_27_47#_c_191_n
+ N_A_27_47#_c_181_n N_A_27_47#_c_182_n N_A_27_47#_c_192_n N_A_27_47#_c_193_n
+ N_A_27_47#_c_194_n N_A_27_47#_c_195_n N_A_27_47#_c_183_n N_A_27_47#_c_184_n
+ N_A_27_47#_c_185_n N_A_27_47#_c_186_n PM_SKY130_FD_SC_HDLL__DLXTN_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__DLXTN_4%D N_D_c_330_n N_D_c_335_n N_D_M1011_g
+ N_D_M1010_g D N_D_c_332_n N_D_c_333_n PM_SKY130_FD_SC_HDLL__DLXTN_4%D
x_PM_SKY130_FD_SC_HDLL__DLXTN_4%A_319_47# N_A_319_47#_M1010_s
+ N_A_319_47#_M1011_s N_A_319_47#_c_373_n N_A_319_47#_c_381_n
+ N_A_319_47#_M1006_g N_A_319_47#_M1007_g N_A_319_47#_c_382_n
+ N_A_319_47#_c_374_n N_A_319_47#_c_383_n N_A_319_47#_c_384_n
+ N_A_319_47#_c_375_n N_A_319_47#_c_376_n N_A_319_47#_c_377_n
+ N_A_319_47#_c_378_n N_A_319_47#_c_379_n
+ PM_SKY130_FD_SC_HDLL__DLXTN_4%A_319_47#
x_PM_SKY130_FD_SC_HDLL__DLXTN_4%A_211_363# N_A_211_363#_M1001_d
+ N_A_211_363#_M1019_d N_A_211_363#_c_463_n N_A_211_363#_c_468_n
+ N_A_211_363#_c_469_n N_A_211_363#_M1018_g N_A_211_363#_c_464_n
+ N_A_211_363#_M1000_g N_A_211_363#_c_471_n N_A_211_363#_c_472_n
+ N_A_211_363#_c_473_n N_A_211_363#_c_474_n N_A_211_363#_c_466_n
+ PM_SKY130_FD_SC_HDLL__DLXTN_4%A_211_363#
x_PM_SKY130_FD_SC_HDLL__DLXTN_4%A_774_21# N_A_774_21#_M1014_s
+ N_A_774_21#_M1017_s N_A_774_21#_M1009_g N_A_774_21#_c_574_n
+ N_A_774_21#_M1022_g N_A_774_21#_c_575_n N_A_774_21#_M1002_g
+ N_A_774_21#_c_566_n N_A_774_21#_M1003_g N_A_774_21#_c_576_n
+ N_A_774_21#_M1013_g N_A_774_21#_c_567_n N_A_774_21#_M1005_g
+ N_A_774_21#_c_577_n N_A_774_21#_M1020_g N_A_774_21#_c_568_n
+ N_A_774_21#_M1012_g N_A_774_21#_c_578_n N_A_774_21#_M1023_g
+ N_A_774_21#_c_569_n N_A_774_21#_M1021_g N_A_774_21#_c_579_n
+ N_A_774_21#_c_614_p N_A_774_21#_c_570_n N_A_774_21#_c_580_n
+ N_A_774_21#_c_571_n N_A_774_21#_c_596_p N_A_774_21#_c_597_p
+ N_A_774_21#_c_572_n PM_SKY130_FD_SC_HDLL__DLXTN_4%A_774_21#
x_PM_SKY130_FD_SC_HDLL__DLXTN_4%A_609_413# N_A_609_413#_M1008_d
+ N_A_609_413#_M1018_d N_A_609_413#_c_690_n N_A_609_413#_M1017_g
+ N_A_609_413#_c_684_n N_A_609_413#_M1014_g N_A_609_413#_c_685_n
+ N_A_609_413#_c_686_n N_A_609_413#_c_695_n N_A_609_413#_c_697_n
+ N_A_609_413#_c_687_n N_A_609_413#_c_693_n N_A_609_413#_c_688_n
+ N_A_609_413#_c_689_n PM_SKY130_FD_SC_HDLL__DLXTN_4%A_609_413#
x_PM_SKY130_FD_SC_HDLL__DLXTN_4%VPWR N_VPWR_M1004_d N_VPWR_M1011_d
+ N_VPWR_M1022_d N_VPWR_M1017_d N_VPWR_M1013_s N_VPWR_M1023_s N_VPWR_c_763_n
+ N_VPWR_c_764_n N_VPWR_c_765_n N_VPWR_c_766_n N_VPWR_c_767_n N_VPWR_c_768_n
+ N_VPWR_c_769_n N_VPWR_c_770_n N_VPWR_c_771_n N_VPWR_c_772_n N_VPWR_c_773_n
+ VPWR N_VPWR_c_774_n N_VPWR_c_775_n N_VPWR_c_776_n N_VPWR_c_777_n
+ N_VPWR_c_778_n N_VPWR_c_779_n N_VPWR_c_780_n N_VPWR_c_762_n
+ PM_SKY130_FD_SC_HDLL__DLXTN_4%VPWR
x_PM_SKY130_FD_SC_HDLL__DLXTN_4%Q N_Q_M1003_d N_Q_M1012_d N_Q_M1002_d
+ N_Q_M1020_d N_Q_c_882_n N_Q_c_890_n N_Q_c_885_n N_Q_c_898_n Q Q Q Q Q Q Q Q Q
+ Q N_Q_c_910_n Q Q PM_SKY130_FD_SC_HDLL__DLXTN_4%Q
x_PM_SKY130_FD_SC_HDLL__DLXTN_4%VGND N_VGND_M1016_d N_VGND_M1010_d
+ N_VGND_M1009_d N_VGND_M1014_d N_VGND_M1005_s N_VGND_M1021_s N_VGND_c_932_n
+ N_VGND_c_933_n N_VGND_c_934_n N_VGND_c_935_n N_VGND_c_936_n N_VGND_c_937_n
+ N_VGND_c_938_n VGND N_VGND_c_939_n N_VGND_c_940_n N_VGND_c_941_n
+ N_VGND_c_942_n N_VGND_c_943_n N_VGND_c_944_n N_VGND_c_945_n N_VGND_c_946_n
+ N_VGND_c_947_n N_VGND_c_948_n PM_SKY130_FD_SC_HDLL__DLXTN_4%VGND
cc_1 VNB N_GATE_N_c_137_n 0.0173562f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_2 VNB N_GATE_N_c_138_n 0.0272334f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_3 VNB GATE_N 0.0156215f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_GATE_N_c_140_n 0.0217779f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_GATE_N_c_141_n 0.0136718f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_6 VNB N_A_27_47#_M1001_g 0.0409473f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_179_n 0.00253943f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.19
cc_8 VNB N_A_27_47#_c_180_n 0.00649765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_181_n 0.0314041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_182_n 0.00433768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_183_n 0.00733671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_184_n 0.0266603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_185_n 0.0179916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_186_n 0.00507045f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_D_c_330_n 0.00677792f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.07
cc_16 VNB N_D_M1010_g 0.0261824f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_17 VNB N_D_c_332_n 0.00682796f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_D_c_333_n 0.0452157f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.665
cc_19 VNB N_A_319_47#_c_373_n 0.0143712f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_20 VNB N_A_319_47#_c_374_n 0.00320313f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_21 VNB N_A_319_47#_c_375_n 0.00579201f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_22 VNB N_A_319_47#_c_376_n 0.00340984f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_23 VNB N_A_319_47#_c_377_n 0.00287801f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_24 VNB N_A_319_47#_c_378_n 0.0307071f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_319_47#_c_379_n 0.0180872f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_211_363#_c_463_n 0.00637303f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_27 VNB N_A_211_363#_c_464_n 0.013345f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_211_363#_M1000_g 0.0465169f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_211_363#_c_466_n 0.0139676f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_774_21#_M1009_g 0.0481327f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_31 VNB N_A_774_21#_c_566_n 0.0172779f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.665
cc_32 VNB N_A_774_21#_c_567_n 0.016491f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_33 VNB N_A_774_21#_c_568_n 0.0169182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_774_21#_c_569_n 0.0223996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_774_21#_c_570_n 0.00260453f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_774_21#_c_571_n 0.00316203f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_774_21#_c_572_n 0.0824221f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_609_413#_c_684_n 0.0199931f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_39 VNB N_A_609_413#_c_685_n 0.0479719f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_40 VNB N_A_609_413#_c_686_n 0.0124501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_609_413#_c_687_n 0.00299652f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_42 VNB N_A_609_413#_c_688_n 0.00582053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_609_413#_c_689_n 0.00274485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VPWR_c_762_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_Q_c_882_n 0.00105358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB Q 0.00193786f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_47 VNB Q 0.0197851f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_932_n 0.00472484f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_933_n 0.00536307f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_50 VNB N_VGND_c_934_n 0.00516693f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_935_n 0.0113721f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_52 VNB N_VGND_c_936_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_937_n 0.0489444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_938_n 0.00324439f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_939_n 0.0154125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_940_n 0.0298657f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_941_n 0.0241012f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_942_n 0.0198444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_943_n 0.0199261f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_944_n 0.0085923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_945_n 0.00859087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_946_n 0.00548191f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_947_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_948_n 0.378435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VPB N_GATE_N_c_142_n 0.0108902f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_66 VPB N_GATE_N_c_143_n 0.0470277f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.74
cc_67 VPB GATE_N 0.0156114f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_68 VPB N_GATE_N_c_140_n 0.0110489f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_69 VPB N_A_27_47#_c_187_n 0.0189977f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_70 VPB N_A_27_47#_c_188_n 0.0258635f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_71 VPB N_A_27_47#_c_189_n 0.0513172f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_72 VPB N_A_27_47#_c_190_n 0.00132472f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_47#_c_191_n 0.00364092f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_47#_c_192_n 0.00288926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_47#_c_193_n 0.00293305f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_47#_c_194_n 0.0104382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_47#_c_195_n 0.0243318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_47#_c_183_n 0.00320855f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_27_47#_c_184_n 0.0122042f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_27_47#_c_186_n 2.1875e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_D_c_330_n 0.0240874f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.07
cc_82 VPB N_D_c_335_n 0.0271119f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.4
cc_83 VPB N_D_c_332_n 0.00328738f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_319_47#_c_373_n 0.0191153f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_85 VPB N_A_319_47#_c_381_n 0.0226052f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_86 VPB N_A_319_47#_c_382_n 0.00765308f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.665
cc_87 VPB N_A_319_47#_c_383_n 0.00424606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_319_47#_c_384_n 0.00286464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_319_47#_c_376_n 0.00369206f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_90 VPB N_A_211_363#_c_463_n 0.0314554f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_91 VPB N_A_211_363#_c_468_n 0.0111674f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_92 VPB N_A_211_363#_c_469_n 0.0230242f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_93 VPB N_A_211_363#_c_464_n 0.017856f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_211_363#_c_471_n 0.00178424f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_95 VPB N_A_211_363#_c_472_n 0.00135179f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_96 VPB N_A_211_363#_c_473_n 0.00645783f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.19
cc_97 VPB N_A_211_363#_c_474_n 0.0130463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_211_363#_c_466_n 0.011923f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_774_21#_M1009_g 0.0157135f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_100 VPB N_A_774_21#_c_574_n 0.074699f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_101 VPB N_A_774_21#_c_575_n 0.0163255f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_774_21#_c_576_n 0.0159305f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_103 VPB N_A_774_21#_c_577_n 0.0160611f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_104 VPB N_A_774_21#_c_578_n 0.0207606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_774_21#_c_579_n 0.00729205f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_774_21#_c_580_n 0.00379503f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_774_21#_c_571_n 0.00281539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_774_21#_c_572_n 0.0562593f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_609_413#_c_690_n 0.0194297f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_110 VPB N_A_609_413#_c_685_n 0.0158736f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.805
cc_111 VPB N_A_609_413#_c_686_n 0.00700558f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_609_413#_c_693_n 0.0057329f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_113 VPB N_A_609_413#_c_688_n 0.00221288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_763_n 0.00126291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_764_n 0.00367613f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_116 VPB N_VPWR_c_765_n 0.00470153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_766_n 0.00260949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_767_n 0.00238371f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_768_n 0.0113462f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_769_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_770_n 0.0332128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_771_n 0.00446482f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_772_n 0.043878f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_773_n 0.00324376f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_774_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_775_n 0.0234599f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_776_n 0.0180975f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_777_n 0.0183743f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_778_n 0.0054556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_779_n 0.00427244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_780_n 0.00359922f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_762_n 0.061069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_Q_c_885_n 0.00154178f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB Q 0.00133662f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_135 VPB Q 0.00657623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 N_GATE_N_c_143_n N_A_27_47#_c_187_n 0.00668506f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_137 GATE_N N_A_27_47#_c_187_n 3.7104e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_138 N_GATE_N_c_140_n N_A_27_47#_c_187_n 0.00242709f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_139 N_GATE_N_c_143_n N_A_27_47#_c_188_n 0.0192779f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_140 N_GATE_N_c_137_n N_A_27_47#_M1001_g 0.0154184f $X=0.52 $Y=0.73 $X2=0
+ $Y2=0
cc_141 N_GATE_N_c_141_n N_A_27_47#_M1001_g 0.00177708f $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_142 N_GATE_N_c_137_n N_A_27_47#_c_179_n 0.00643492f $X=0.52 $Y=0.73 $X2=0
+ $Y2=0
cc_143 N_GATE_N_c_138_n N_A_27_47#_c_179_n 0.0137188f $X=0.52 $Y=0.805 $X2=0
+ $Y2=0
cc_144 N_GATE_N_c_138_n N_A_27_47#_c_180_n 0.00657185f $X=0.52 $Y=0.805 $X2=0
+ $Y2=0
cc_145 GATE_N N_A_27_47#_c_180_n 0.0125186f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_146 N_GATE_N_c_140_n N_A_27_47#_c_180_n 3.35813e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_147 N_GATE_N_c_143_n N_A_27_47#_c_190_n 0.0189751f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_148 N_GATE_N_c_143_n N_A_27_47#_c_191_n 0.00836964f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_149 GATE_N N_A_27_47#_c_191_n 0.0139005f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_150 N_GATE_N_c_140_n N_A_27_47#_c_191_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_151 N_GATE_N_c_143_n N_A_27_47#_c_192_n 2.26411e-19 $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_152 GATE_N N_A_27_47#_c_192_n 0.00684198f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_153 N_GATE_N_c_140_n N_A_27_47#_c_192_n 0.00225027f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_154 N_GATE_N_c_143_n N_A_27_47#_c_183_n 0.00465299f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_155 N_GATE_N_c_138_n N_A_27_47#_c_183_n 0.00196813f $X=0.52 $Y=0.805 $X2=0
+ $Y2=0
cc_156 GATE_N N_A_27_47#_c_183_n 0.0249872f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_157 N_GATE_N_c_140_n N_A_27_47#_c_183_n 0.00189147f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_158 N_GATE_N_c_141_n N_A_27_47#_c_183_n 0.00128063f $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_159 GATE_N N_A_27_47#_c_184_n 0.00100538f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_160 N_GATE_N_c_140_n N_A_27_47#_c_184_n 0.0129544f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_161 N_GATE_N_c_143_n N_VPWR_c_763_n 0.0125197f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_162 N_GATE_N_c_143_n N_VPWR_c_774_n 0.00304525f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_163 N_GATE_N_c_143_n N_VPWR_c_762_n 0.00454898f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_164 N_GATE_N_c_137_n N_VGND_c_939_n 0.00198377f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_165 N_GATE_N_c_138_n N_VGND_c_939_n 6.41851e-19 $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_166 N_GATE_N_c_137_n N_VGND_c_944_n 0.0142867f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_167 N_GATE_N_c_137_n N_VGND_c_948_n 0.00367064f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_195_n N_D_c_330_n 0.00789696f $X=3.115 $Y=1.485 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_195_n N_D_c_332_n 0.012909f $X=3.115 $Y=1.485 $X2=0 $Y2=0
cc_170 N_A_27_47#_M1001_g N_D_c_333_n 0.00523969f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_195_n N_A_319_47#_c_373_n 0.00625272f $X=3.115 $Y=1.485
+ $X2=0 $Y2=0
cc_172 N_A_27_47#_c_186_n N_A_319_47#_c_373_n 0.00363102f $X=3.37 $Y=1.415 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_c_195_n N_A_319_47#_c_383_n 0.0135374f $X=3.115 $Y=1.485 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_c_195_n N_A_319_47#_c_384_n 0.0114021f $X=3.115 $Y=1.485 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_c_181_n N_A_319_47#_c_375_n 9.85912e-19 $X=3 $Y=0.87 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_c_182_n N_A_319_47#_c_375_n 0.0130183f $X=3.26 $Y=0.87 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_195_n N_A_319_47#_c_375_n 0.00840141f $X=3.115 $Y=1.485
+ $X2=0 $Y2=0
cc_178 N_A_27_47#_c_186_n N_A_319_47#_c_375_n 0.00168439f $X=3.37 $Y=1.415 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_195_n N_A_319_47#_c_376_n 0.0109087f $X=3.115 $Y=1.485 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_181_n N_A_319_47#_c_378_n 0.0120615f $X=3 $Y=0.87 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_182_n N_A_319_47#_c_378_n 9.79877e-19 $X=3.26 $Y=0.87 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_195_n N_A_319_47#_c_378_n 0.00107604f $X=3.115 $Y=1.485
+ $X2=0 $Y2=0
cc_183 N_A_27_47#_c_186_n N_A_319_47#_c_378_n 9.85161e-19 $X=3.37 $Y=1.415 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_181_n N_A_319_47#_c_379_n 0.0020564f $X=3 $Y=0.87 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_182_n N_A_319_47#_c_379_n 2.08303e-19 $X=3.26 $Y=0.87 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_185_n N_A_319_47#_c_379_n 0.0174883f $X=3.025 $Y=0.705 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_189_n N_A_211_363#_c_463_n 0.0123807f $X=3.425 $Y=1.99 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_181_n N_A_211_363#_c_463_n 0.0221963f $X=3 $Y=0.87 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_182_n N_A_211_363#_c_463_n 0.00174975f $X=3.26 $Y=0.87 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_193_n N_A_211_363#_c_463_n 0.00185365f $X=3.26 $Y=1.485
+ $X2=0 $Y2=0
cc_191 N_A_27_47#_c_195_n N_A_211_363#_c_463_n 0.00700268f $X=3.115 $Y=1.485
+ $X2=0 $Y2=0
cc_192 N_A_27_47#_c_186_n N_A_211_363#_c_463_n 0.00360536f $X=3.37 $Y=1.415
+ $X2=0 $Y2=0
cc_193 N_A_27_47#_c_189_n N_A_211_363#_c_468_n 0.00494294f $X=3.425 $Y=1.99
+ $X2=0 $Y2=0
cc_194 N_A_27_47#_c_194_n N_A_211_363#_c_468_n 0.00360536f $X=3.26 $Y=1.485
+ $X2=0 $Y2=0
cc_195 N_A_27_47#_c_189_n N_A_211_363#_c_469_n 0.0140166f $X=3.425 $Y=1.99 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_189_n N_A_211_363#_c_464_n 0.0151523f $X=3.425 $Y=1.99 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_182_n N_A_211_363#_c_464_n 7.03475e-19 $X=3.26 $Y=0.87 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_193_n N_A_211_363#_c_464_n 0.00437354f $X=3.26 $Y=1.485
+ $X2=0 $Y2=0
cc_199 N_A_27_47#_c_194_n N_A_211_363#_c_464_n 0.00589636f $X=3.26 $Y=1.485
+ $X2=0 $Y2=0
cc_200 N_A_27_47#_c_195_n N_A_211_363#_c_464_n 0.00133008f $X=3.115 $Y=1.485
+ $X2=0 $Y2=0
cc_201 N_A_27_47#_c_186_n N_A_211_363#_c_464_n 0.0137322f $X=3.37 $Y=1.415 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_181_n N_A_211_363#_M1000_g 0.0192996f $X=3 $Y=0.87 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_182_n N_A_211_363#_M1000_g 0.00367077f $X=3.26 $Y=0.87 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_185_n N_A_211_363#_M1000_g 0.0127891f $X=3.025 $Y=0.705
+ $X2=0 $Y2=0
cc_205 N_A_27_47#_c_186_n N_A_211_363#_M1000_g 0.0053616f $X=3.37 $Y=1.415 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_188_n N_A_211_363#_c_471_n 0.00228048f $X=0.965 $Y=1.74
+ $X2=0 $Y2=0
cc_207 N_A_27_47#_c_190_n N_A_211_363#_c_471_n 0.00571095f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_c_195_n N_A_211_363#_c_471_n 0.0274397f $X=3.115 $Y=1.485
+ $X2=0 $Y2=0
cc_209 N_A_27_47#_c_183_n N_A_211_363#_c_471_n 0.00136602f $X=0.805 $Y=1.235
+ $X2=0 $Y2=0
cc_210 N_A_27_47#_c_194_n N_A_211_363#_c_472_n 0.00157421f $X=3.26 $Y=1.485
+ $X2=0 $Y2=0
cc_211 N_A_27_47#_c_195_n N_A_211_363#_c_472_n 0.0267994f $X=3.115 $Y=1.485
+ $X2=0 $Y2=0
cc_212 N_A_27_47#_c_195_n N_A_211_363#_c_473_n 0.0996761f $X=3.115 $Y=1.485
+ $X2=0 $Y2=0
cc_213 N_A_27_47#_c_189_n N_A_211_363#_c_474_n 3.94094e-19 $X=3.425 $Y=1.99
+ $X2=0 $Y2=0
cc_214 N_A_27_47#_c_181_n N_A_211_363#_c_474_n 3.90521e-19 $X=3 $Y=0.87 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_182_n N_A_211_363#_c_474_n 0.00161882f $X=3.26 $Y=0.87 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_193_n N_A_211_363#_c_474_n 0.00256606f $X=3.26 $Y=1.485
+ $X2=0 $Y2=0
cc_217 N_A_27_47#_c_195_n N_A_211_363#_c_474_n 0.0244544f $X=3.115 $Y=1.485
+ $X2=0 $Y2=0
cc_218 N_A_27_47#_c_186_n N_A_211_363#_c_474_n 0.0364655f $X=3.37 $Y=1.415 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_c_188_n N_A_211_363#_c_466_n 0.0065629f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_M1001_g N_A_211_363#_c_466_n 0.0217846f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_c_179_n N_A_211_363#_c_466_n 0.0103633f $X=0.66 $Y=0.72 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_c_190_n N_A_211_363#_c_466_n 0.0085487f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_192_n N_A_211_363#_c_466_n 0.00212801f $X=0.89 $Y=1.485
+ $X2=0 $Y2=0
cc_224 N_A_27_47#_c_195_n N_A_211_363#_c_466_n 0.0182722f $X=3.115 $Y=1.485
+ $X2=0 $Y2=0
cc_225 N_A_27_47#_c_183_n N_A_211_363#_c_466_n 0.0567523f $X=0.805 $Y=1.235
+ $X2=0 $Y2=0
cc_226 N_A_27_47#_c_194_n N_A_774_21#_M1009_g 0.0011227f $X=3.26 $Y=1.485 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_186_n N_A_774_21#_M1009_g 2.24311e-19 $X=3.37 $Y=1.415 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_c_189_n N_A_774_21#_c_574_n 0.0395287f $X=3.425 $Y=1.99 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_c_194_n N_A_774_21#_c_574_n 6.47236e-19 $X=3.26 $Y=1.485 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_189_n N_A_609_413#_c_695_n 0.0124489f $X=3.425 $Y=1.99 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_194_n N_A_609_413#_c_695_n 0.0172324f $X=3.26 $Y=1.485 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_181_n N_A_609_413#_c_697_n 0.00144439f $X=3 $Y=0.87 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_182_n N_A_609_413#_c_697_n 0.0162478f $X=3.26 $Y=0.87 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_185_n N_A_609_413#_c_697_n 0.00440823f $X=3.025 $Y=0.705
+ $X2=0 $Y2=0
cc_235 N_A_27_47#_c_182_n N_A_609_413#_c_687_n 0.0121655f $X=3.26 $Y=0.87 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_189_n N_A_609_413#_c_693_n 0.00712699f $X=3.425 $Y=1.99
+ $X2=0 $Y2=0
cc_237 N_A_27_47#_c_193_n N_A_609_413#_c_693_n 0.00202292f $X=3.26 $Y=1.485
+ $X2=0 $Y2=0
cc_238 N_A_27_47#_c_194_n N_A_609_413#_c_693_n 0.0373254f $X=3.26 $Y=1.485 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_186_n N_A_609_413#_c_693_n 0.00258815f $X=3.37 $Y=1.415
+ $X2=0 $Y2=0
cc_240 N_A_27_47#_c_182_n N_A_609_413#_c_689_n 0.00183439f $X=3.26 $Y=0.87 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_186_n N_A_609_413#_c_689_n 0.0124639f $X=3.37 $Y=1.415 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_190_n N_VPWR_M1004_d 0.001889f $X=0.66 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_243 N_A_27_47#_c_188_n N_VPWR_c_763_n 0.00960416f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_c_190_n N_VPWR_c_763_n 0.0208334f $X=0.66 $Y=1.88 $X2=0 $Y2=0
cc_245 N_A_27_47#_c_191_n N_VPWR_c_763_n 0.0246493f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_246 N_A_27_47#_c_192_n N_VPWR_c_763_n 0.00106399f $X=0.89 $Y=1.485 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_195_n N_VPWR_c_764_n 0.0018348f $X=3.115 $Y=1.485 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_188_n N_VPWR_c_770_n 0.00590576f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_189_n N_VPWR_c_772_n 0.00439333f $X=3.425 $Y=1.99 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_190_n N_VPWR_c_774_n 0.00180073f $X=0.66 $Y=1.88 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_191_n N_VPWR_c_774_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_188_n N_VPWR_c_762_n 0.0113647f $X=0.965 $Y=1.74 $X2=0 $Y2=0
cc_253 N_A_27_47#_c_189_n N_VPWR_c_762_n 0.0063084f $X=3.425 $Y=1.99 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_190_n N_VPWR_c_762_n 0.00528325f $X=0.66 $Y=1.88 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_191_n N_VPWR_c_762_n 0.00646745f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_256 N_A_27_47#_c_179_n N_VGND_M1016_d 0.00227127f $X=0.66 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_257 N_A_27_47#_c_181_n N_VGND_c_937_n 0.00166672f $X=3 $Y=0.87 $X2=0 $Y2=0
cc_258 N_A_27_47#_c_182_n N_VGND_c_937_n 0.00255568f $X=3.26 $Y=0.87 $X2=0 $Y2=0
cc_259 N_A_27_47#_c_185_n N_VGND_c_937_n 0.00425892f $X=3.025 $Y=0.705 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_316_p N_VGND_c_939_n 0.00725596f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_261 N_A_27_47#_c_179_n N_VGND_c_939_n 0.00244154f $X=0.66 $Y=0.72 $X2=0 $Y2=0
cc_262 N_A_27_47#_M1001_g N_VGND_c_940_n 0.00585385f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_M1001_g N_VGND_c_944_n 0.00317372f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_316_p N_VGND_c_944_n 0.00895866f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_179_n N_VGND_c_944_n 0.0228644f $X=0.66 $Y=0.72 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_184_n N_VGND_c_944_n 6.84207e-19 $X=0.99 $Y=1.235 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_M1016_s N_VGND_c_948_n 0.00437169f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_M1001_g N_VGND_c_948_n 0.0120602f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_269 N_A_27_47#_c_316_p N_VGND_c_948_n 0.00608739f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_270 N_A_27_47#_c_179_n N_VGND_c_948_n 0.00625251f $X=0.66 $Y=0.72 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_181_n N_VGND_c_948_n 0.00243808f $X=3 $Y=0.87 $X2=0 $Y2=0
cc_272 N_A_27_47#_c_182_n N_VGND_c_948_n 0.0046064f $X=3.26 $Y=0.87 $X2=0 $Y2=0
cc_273 N_A_27_47#_c_185_n N_VGND_c_948_n 0.00638862f $X=3.025 $Y=0.705 $X2=0
+ $Y2=0
cc_274 N_D_c_333_n N_A_319_47#_c_373_n 0.0145035f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_275 N_D_c_330_n N_A_319_47#_c_381_n 0.0145035f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_276 N_D_c_335_n N_A_319_47#_c_381_n 0.00935018f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_277 N_D_c_335_n N_A_319_47#_c_382_n 0.0136011f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_278 N_D_M1010_g N_A_319_47#_c_374_n 0.0153745f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_279 N_D_c_332_n N_A_319_47#_c_374_n 0.00639931f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_280 N_D_c_333_n N_A_319_47#_c_374_n 0.0029398f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_281 N_D_c_330_n N_A_319_47#_c_383_n 0.0106635f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_282 N_D_c_330_n N_A_319_47#_c_384_n 0.00412429f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_283 N_D_c_332_n N_A_319_47#_c_384_n 0.0233961f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_284 N_D_c_333_n N_A_319_47#_c_384_n 0.00131849f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_285 N_D_M1010_g N_A_319_47#_c_375_n 0.00591272f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_286 N_D_c_332_n N_A_319_47#_c_375_n 0.00919404f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_287 N_D_c_332_n N_A_319_47#_c_376_n 0.0139605f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_288 N_D_c_333_n N_A_319_47#_c_376_n 0.0057769f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_289 N_D_M1010_g N_A_319_47#_c_377_n 8.59557e-19 $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_290 N_D_c_332_n N_A_319_47#_c_377_n 0.0138491f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_291 N_D_c_333_n N_A_319_47#_c_377_n 0.0042466f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_292 N_D_M1010_g N_A_319_47#_c_378_n 0.0198512f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_293 N_D_M1010_g N_A_319_47#_c_379_n 0.0127335f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_294 N_D_c_335_n N_A_211_363#_c_473_n 0.00420236f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_295 N_D_c_330_n N_A_211_363#_c_466_n 0.00494044f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_296 N_D_c_335_n N_A_211_363#_c_466_n 0.00105075f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_297 N_D_M1010_g N_A_211_363#_c_466_n 0.00193515f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_298 N_D_c_332_n N_A_211_363#_c_466_n 0.0276277f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_299 N_D_c_333_n N_A_211_363#_c_466_n 0.00238672f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_300 N_D_c_335_n N_VPWR_c_764_n 0.00664063f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_301 N_D_c_335_n N_VPWR_c_770_n 0.00674916f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_302 N_D_c_335_n N_VPWR_c_762_n 0.00848136f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_303 N_D_M1010_g N_VGND_c_940_n 0.00196986f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_304 N_D_M1010_g N_VGND_c_945_n 0.0139983f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_305 N_D_M1010_g N_VGND_c_948_n 0.00398772f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_306 N_D_c_333_n N_VGND_c_948_n 0.00103829f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_307 N_A_319_47#_c_373_n N_A_211_363#_c_463_n 0.0253561f $X=2.425 $Y=1.67
+ $X2=0 $Y2=0
cc_308 N_A_319_47#_c_381_n N_A_211_363#_c_468_n 0.0105715f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_309 N_A_319_47#_c_381_n N_A_211_363#_c_469_n 0.022499f $X=2.425 $Y=1.77 $X2=0
+ $Y2=0
cc_310 N_A_319_47#_c_382_n N_A_211_363#_c_471_n 0.00264542f $X=1.72 $Y=1.99
+ $X2=0 $Y2=0
cc_311 N_A_319_47#_c_381_n N_A_211_363#_c_472_n 0.00150338f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_312 N_A_319_47#_c_381_n N_A_211_363#_c_473_n 0.00506867f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_313 N_A_319_47#_c_382_n N_A_211_363#_c_473_n 0.0233342f $X=1.72 $Y=1.99 $X2=0
+ $Y2=0
cc_314 N_A_319_47#_c_383_n N_A_211_363#_c_473_n 0.00667484f $X=2.12 $Y=1.58
+ $X2=0 $Y2=0
cc_315 N_A_319_47#_c_373_n N_A_211_363#_c_474_n 0.004659f $X=2.425 $Y=1.67 $X2=0
+ $Y2=0
cc_316 N_A_319_47#_c_381_n N_A_211_363#_c_474_n 0.00233669f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_317 N_A_319_47#_c_383_n N_A_211_363#_c_474_n 0.00664087f $X=2.12 $Y=1.58
+ $X2=0 $Y2=0
cc_318 N_A_319_47#_c_376_n N_A_211_363#_c_474_n 0.00578855f $X=2.205 $Y=1.495
+ $X2=0 $Y2=0
cc_319 N_A_319_47#_c_382_n N_A_211_363#_c_466_n 0.0392174f $X=1.72 $Y=1.99 $X2=0
+ $Y2=0
cc_320 N_A_319_47#_c_384_n N_A_211_363#_c_466_n 0.00880329f $X=1.885 $Y=1.58
+ $X2=0 $Y2=0
cc_321 N_A_319_47#_c_377_n N_A_211_363#_c_466_n 0.0191835f $X=1.72 $Y=0.51 $X2=0
+ $Y2=0
cc_322 N_A_319_47#_c_381_n N_A_609_413#_c_695_n 4.98758e-19 $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_323 N_A_319_47#_c_379_n N_A_609_413#_c_697_n 7.53078e-19 $X=2.43 $Y=0.765
+ $X2=0 $Y2=0
cc_324 N_A_319_47#_c_381_n N_VPWR_c_764_n 0.0227809f $X=2.425 $Y=1.77 $X2=0
+ $Y2=0
cc_325 N_A_319_47#_c_382_n N_VPWR_c_764_n 0.0355228f $X=1.72 $Y=1.99 $X2=0 $Y2=0
cc_326 N_A_319_47#_c_383_n N_VPWR_c_764_n 0.013562f $X=2.12 $Y=1.58 $X2=0 $Y2=0
cc_327 N_A_319_47#_c_382_n N_VPWR_c_770_n 0.0159613f $X=1.72 $Y=1.99 $X2=0 $Y2=0
cc_328 N_A_319_47#_c_381_n N_VPWR_c_772_n 0.00368966f $X=2.425 $Y=1.77 $X2=0
+ $Y2=0
cc_329 N_A_319_47#_M1011_s N_VPWR_c_762_n 0.00181388f $X=1.595 $Y=1.845 $X2=0
+ $Y2=0
cc_330 N_A_319_47#_c_381_n N_VPWR_c_762_n 0.00386434f $X=2.425 $Y=1.77 $X2=0
+ $Y2=0
cc_331 N_A_319_47#_c_382_n N_VPWR_c_762_n 0.0057885f $X=1.72 $Y=1.99 $X2=0 $Y2=0
cc_332 N_A_319_47#_c_375_n N_VGND_M1010_d 0.00229352f $X=2.205 $Y=1.095 $X2=0
+ $Y2=0
cc_333 N_A_319_47#_c_378_n N_VGND_c_937_n 0.00112938f $X=2.405 $Y=0.93 $X2=0
+ $Y2=0
cc_334 N_A_319_47#_c_379_n N_VGND_c_937_n 0.00585385f $X=2.43 $Y=0.765 $X2=0
+ $Y2=0
cc_335 N_A_319_47#_c_374_n N_VGND_c_940_n 0.00256875f $X=2.12 $Y=0.7 $X2=0 $Y2=0
cc_336 N_A_319_47#_c_377_n N_VGND_c_940_n 0.00723406f $X=1.72 $Y=0.51 $X2=0
+ $Y2=0
cc_337 N_A_319_47#_c_374_n N_VGND_c_945_n 0.00613814f $X=2.12 $Y=0.7 $X2=0 $Y2=0
cc_338 N_A_319_47#_c_375_n N_VGND_c_945_n 0.0161158f $X=2.205 $Y=1.095 $X2=0
+ $Y2=0
cc_339 N_A_319_47#_c_377_n N_VGND_c_945_n 0.00746555f $X=1.72 $Y=0.51 $X2=0
+ $Y2=0
cc_340 N_A_319_47#_c_378_n N_VGND_c_945_n 4.19595e-19 $X=2.405 $Y=0.93 $X2=0
+ $Y2=0
cc_341 N_A_319_47#_c_379_n N_VGND_c_945_n 0.00317372f $X=2.43 $Y=0.765 $X2=0
+ $Y2=0
cc_342 N_A_319_47#_M1010_s N_VGND_c_948_n 0.00343585f $X=1.595 $Y=0.235 $X2=0
+ $Y2=0
cc_343 N_A_319_47#_c_374_n N_VGND_c_948_n 0.0051978f $X=2.12 $Y=0.7 $X2=0 $Y2=0
cc_344 N_A_319_47#_c_375_n N_VGND_c_948_n 0.00710218f $X=2.205 $Y=1.095 $X2=0
+ $Y2=0
cc_345 N_A_319_47#_c_377_n N_VGND_c_948_n 0.00607883f $X=1.72 $Y=0.51 $X2=0
+ $Y2=0
cc_346 N_A_319_47#_c_378_n N_VGND_c_948_n 0.00117722f $X=2.405 $Y=0.93 $X2=0
+ $Y2=0
cc_347 N_A_319_47#_c_379_n N_VGND_c_948_n 0.0065019f $X=2.43 $Y=0.765 $X2=0
+ $Y2=0
cc_348 N_A_211_363#_M1000_g N_A_774_21#_M1009_g 0.0465716f $X=3.47 $Y=0.415
+ $X2=0 $Y2=0
cc_349 N_A_211_363#_c_469_n N_A_609_413#_c_695_n 0.00431285f $X=2.955 $Y=1.99
+ $X2=0 $Y2=0
cc_350 N_A_211_363#_M1000_g N_A_609_413#_c_697_n 0.0131523f $X=3.47 $Y=0.415
+ $X2=0 $Y2=0
cc_351 N_A_211_363#_M1000_g N_A_609_413#_c_687_n 0.00558087f $X=3.47 $Y=0.415
+ $X2=0 $Y2=0
cc_352 N_A_211_363#_c_464_n N_A_609_413#_c_693_n 6.43727e-19 $X=3.395 $Y=1.32
+ $X2=0 $Y2=0
cc_353 N_A_211_363#_M1000_g N_A_609_413#_c_689_n 0.00329131f $X=3.47 $Y=0.415
+ $X2=0 $Y2=0
cc_354 N_A_211_363#_c_473_n N_VPWR_M1011_d 8.51638e-19 $X=2.61 $Y=1.855 $X2=0
+ $Y2=0
cc_355 N_A_211_363#_c_466_n N_VPWR_c_763_n 0.0202126f $X=1.2 $Y=0.51 $X2=0 $Y2=0
cc_356 N_A_211_363#_c_469_n N_VPWR_c_764_n 0.00314538f $X=2.955 $Y=1.99 $X2=0
+ $Y2=0
cc_357 N_A_211_363#_c_472_n N_VPWR_c_764_n 8.70426e-19 $X=2.755 $Y=1.855 $X2=0
+ $Y2=0
cc_358 N_A_211_363#_c_473_n N_VPWR_c_764_n 0.017675f $X=2.61 $Y=1.855 $X2=0
+ $Y2=0
cc_359 N_A_211_363#_c_474_n N_VPWR_c_764_n 0.00794167f $X=2.87 $Y=1.52 $X2=0
+ $Y2=0
cc_360 N_A_211_363#_c_466_n N_VPWR_c_770_n 0.0120448f $X=1.2 $Y=0.51 $X2=0 $Y2=0
cc_361 N_A_211_363#_c_469_n N_VPWR_c_772_n 0.00588257f $X=2.955 $Y=1.99 $X2=0
+ $Y2=0
cc_362 N_A_211_363#_c_474_n N_VPWR_c_772_n 0.00458985f $X=2.87 $Y=1.52 $X2=0
+ $Y2=0
cc_363 N_A_211_363#_c_469_n N_VPWR_c_762_n 0.00926841f $X=2.955 $Y=1.99 $X2=0
+ $Y2=0
cc_364 N_A_211_363#_c_471_n N_VPWR_c_762_n 0.0151917f $X=1.345 $Y=1.855 $X2=0
+ $Y2=0
cc_365 N_A_211_363#_c_472_n N_VPWR_c_762_n 0.0147851f $X=2.755 $Y=1.855 $X2=0
+ $Y2=0
cc_366 N_A_211_363#_c_473_n N_VPWR_c_762_n 0.0597289f $X=2.61 $Y=1.855 $X2=0
+ $Y2=0
cc_367 N_A_211_363#_c_474_n N_VPWR_c_762_n 0.00409402f $X=2.87 $Y=1.52 $X2=0
+ $Y2=0
cc_368 N_A_211_363#_c_466_n N_VPWR_c_762_n 0.00298632f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_369 N_A_211_363#_c_472_n A_503_369# 0.00110422f $X=2.755 $Y=1.855 $X2=-0.19
+ $Y2=-0.24
cc_370 N_A_211_363#_c_473_n A_503_369# 0.00150032f $X=2.61 $Y=1.855 $X2=-0.19
+ $Y2=-0.24
cc_371 N_A_211_363#_c_474_n A_503_369# 0.00329968f $X=2.87 $Y=1.52 $X2=-0.19
+ $Y2=-0.24
cc_372 N_A_211_363#_M1000_g N_VGND_c_937_n 0.0037981f $X=3.47 $Y=0.415 $X2=0
+ $Y2=0
cc_373 N_A_211_363#_c_466_n N_VGND_c_940_n 0.00732874f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_374 N_A_211_363#_M1001_d N_VGND_c_948_n 0.00535012f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_375 N_A_211_363#_M1000_g N_VGND_c_948_n 0.00555936f $X=3.47 $Y=0.415 $X2=0
+ $Y2=0
cc_376 N_A_211_363#_c_466_n N_VGND_c_948_n 0.00616598f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_377 N_A_774_21#_c_574_n N_A_609_413#_c_690_n 0.00329184f $X=3.97 $Y=1.99
+ $X2=0 $Y2=0
cc_378 N_A_774_21#_c_575_n N_A_609_413#_c_690_n 0.0181794f $X=5.445 $Y=1.41
+ $X2=0 $Y2=0
cc_379 N_A_774_21#_c_580_n N_A_609_413#_c_690_n 0.00417068f $X=4.765 $Y=1.535
+ $X2=0 $Y2=0
cc_380 N_A_774_21#_c_566_n N_A_609_413#_c_684_n 0.0173169f $X=5.47 $Y=0.995
+ $X2=0 $Y2=0
cc_381 N_A_774_21#_c_570_n N_A_609_413#_c_684_n 0.00640823f $X=4.755 $Y=0.58
+ $X2=0 $Y2=0
cc_382 N_A_774_21#_M1009_g N_A_609_413#_c_685_n 0.01646f $X=3.945 $Y=0.445 $X2=0
+ $Y2=0
cc_383 N_A_774_21#_c_574_n N_A_609_413#_c_685_n 0.00487525f $X=3.97 $Y=1.99
+ $X2=0 $Y2=0
cc_384 N_A_774_21#_c_579_n N_A_609_413#_c_685_n 0.00879412f $X=4.64 $Y=1.7 $X2=0
+ $Y2=0
cc_385 N_A_774_21#_c_596_p N_A_609_413#_c_685_n 0.00127702f $X=4.725 $Y=1.755
+ $X2=0 $Y2=0
cc_386 N_A_774_21#_c_597_p N_A_609_413#_c_685_n 0.0194877f $X=4.765 $Y=1.16
+ $X2=0 $Y2=0
cc_387 N_A_774_21#_c_580_n N_A_609_413#_c_686_n 0.0036478f $X=4.765 $Y=1.535
+ $X2=0 $Y2=0
cc_388 N_A_774_21#_c_571_n N_A_609_413#_c_686_n 0.0276191f $X=5.405 $Y=1.16
+ $X2=0 $Y2=0
cc_389 N_A_774_21#_c_572_n N_A_609_413#_c_686_n 0.0253766f $X=6.855 $Y=1.202
+ $X2=0 $Y2=0
cc_390 N_A_774_21#_c_574_n N_A_609_413#_c_695_n 0.00565077f $X=3.97 $Y=1.99
+ $X2=0 $Y2=0
cc_391 N_A_774_21#_M1009_g N_A_609_413#_c_697_n 0.00576368f $X=3.945 $Y=0.445
+ $X2=0 $Y2=0
cc_392 N_A_774_21#_M1009_g N_A_609_413#_c_687_n 0.0213862f $X=3.945 $Y=0.445
+ $X2=0 $Y2=0
cc_393 N_A_774_21#_M1009_g N_A_609_413#_c_693_n 0.0120161f $X=3.945 $Y=0.445
+ $X2=0 $Y2=0
cc_394 N_A_774_21#_c_574_n N_A_609_413#_c_693_n 0.0264208f $X=3.97 $Y=1.99 $X2=0
+ $Y2=0
cc_395 N_A_774_21#_c_579_n N_A_609_413#_c_693_n 0.022954f $X=4.64 $Y=1.7 $X2=0
+ $Y2=0
cc_396 N_A_774_21#_M1009_g N_A_609_413#_c_688_n 0.0123103f $X=3.945 $Y=0.445
+ $X2=0 $Y2=0
cc_397 N_A_774_21#_c_574_n N_A_609_413#_c_688_n 0.00820473f $X=3.97 $Y=1.99
+ $X2=0 $Y2=0
cc_398 N_A_774_21#_c_579_n N_A_609_413#_c_688_n 0.02399f $X=4.64 $Y=1.7 $X2=0
+ $Y2=0
cc_399 N_A_774_21#_c_597_p N_A_609_413#_c_688_n 0.0278868f $X=4.765 $Y=1.16
+ $X2=0 $Y2=0
cc_400 N_A_774_21#_M1009_g N_A_609_413#_c_689_n 0.00472825f $X=3.945 $Y=0.445
+ $X2=0 $Y2=0
cc_401 N_A_774_21#_c_574_n N_VPWR_c_765_n 0.0103025f $X=3.97 $Y=1.99 $X2=0 $Y2=0
cc_402 N_A_774_21#_c_579_n N_VPWR_c_765_n 0.00806355f $X=4.64 $Y=1.7 $X2=0 $Y2=0
cc_403 N_A_774_21#_c_614_p N_VPWR_c_765_n 0.013068f $X=4.725 $Y=2.27 $X2=0 $Y2=0
cc_404 N_A_774_21#_c_575_n N_VPWR_c_766_n 0.0192228f $X=5.445 $Y=1.41 $X2=0
+ $Y2=0
cc_405 N_A_774_21#_c_576_n N_VPWR_c_766_n 0.00140509f $X=5.915 $Y=1.41 $X2=0
+ $Y2=0
cc_406 N_A_774_21#_c_571_n N_VPWR_c_766_n 0.0207774f $X=5.405 $Y=1.16 $X2=0
+ $Y2=0
cc_407 N_A_774_21#_c_572_n N_VPWR_c_766_n 0.00160396f $X=6.855 $Y=1.202 $X2=0
+ $Y2=0
cc_408 N_A_774_21#_c_576_n N_VPWR_c_767_n 0.0071945f $X=5.915 $Y=1.41 $X2=0
+ $Y2=0
cc_409 N_A_774_21#_c_577_n N_VPWR_c_767_n 0.0184093f $X=6.385 $Y=1.41 $X2=0
+ $Y2=0
cc_410 N_A_774_21#_c_578_n N_VPWR_c_767_n 0.00139722f $X=6.855 $Y=1.41 $X2=0
+ $Y2=0
cc_411 N_A_774_21#_c_572_n N_VPWR_c_767_n 0.00527012f $X=6.855 $Y=1.202 $X2=0
+ $Y2=0
cc_412 N_A_774_21#_c_578_n N_VPWR_c_769_n 0.0121267f $X=6.855 $Y=1.41 $X2=0
+ $Y2=0
cc_413 N_A_774_21#_c_574_n N_VPWR_c_772_n 0.00621666f $X=3.97 $Y=1.99 $X2=0
+ $Y2=0
cc_414 N_A_774_21#_c_614_p N_VPWR_c_775_n 0.0115253f $X=4.725 $Y=2.27 $X2=0
+ $Y2=0
cc_415 N_A_774_21#_c_575_n N_VPWR_c_776_n 0.00622633f $X=5.445 $Y=1.41 $X2=0
+ $Y2=0
cc_416 N_A_774_21#_c_576_n N_VPWR_c_776_n 0.00598673f $X=5.915 $Y=1.41 $X2=0
+ $Y2=0
cc_417 N_A_774_21#_c_577_n N_VPWR_c_777_n 0.00622633f $X=6.385 $Y=1.41 $X2=0
+ $Y2=0
cc_418 N_A_774_21#_c_578_n N_VPWR_c_777_n 0.00643798f $X=6.855 $Y=1.41 $X2=0
+ $Y2=0
cc_419 N_A_774_21#_M1017_s N_VPWR_c_762_n 0.00284579f $X=4.6 $Y=1.485 $X2=0
+ $Y2=0
cc_420 N_A_774_21#_c_574_n N_VPWR_c_762_n 0.0144537f $X=3.97 $Y=1.99 $X2=0 $Y2=0
cc_421 N_A_774_21#_c_575_n N_VPWR_c_762_n 0.0104011f $X=5.445 $Y=1.41 $X2=0
+ $Y2=0
cc_422 N_A_774_21#_c_576_n N_VPWR_c_762_n 0.00999552f $X=5.915 $Y=1.41 $X2=0
+ $Y2=0
cc_423 N_A_774_21#_c_577_n N_VPWR_c_762_n 0.0104011f $X=6.385 $Y=1.41 $X2=0
+ $Y2=0
cc_424 N_A_774_21#_c_578_n N_VPWR_c_762_n 0.0120253f $X=6.855 $Y=1.41 $X2=0
+ $Y2=0
cc_425 N_A_774_21#_c_579_n N_VPWR_c_762_n 0.0129053f $X=4.64 $Y=1.7 $X2=0 $Y2=0
cc_426 N_A_774_21#_c_614_p N_VPWR_c_762_n 0.00827281f $X=4.725 $Y=2.27 $X2=0
+ $Y2=0
cc_427 N_A_774_21#_c_566_n N_Q_c_882_n 0.00524009f $X=5.47 $Y=0.995 $X2=0 $Y2=0
cc_428 N_A_774_21#_c_567_n N_Q_c_882_n 0.00602488f $X=5.94 $Y=0.995 $X2=0 $Y2=0
cc_429 N_A_774_21#_c_575_n N_Q_c_890_n 0.00473677f $X=5.445 $Y=1.41 $X2=0 $Y2=0
cc_430 N_A_774_21#_c_576_n N_Q_c_890_n 0.00346986f $X=5.915 $Y=1.41 $X2=0 $Y2=0
cc_431 N_A_774_21#_c_577_n N_Q_c_890_n 3.75009e-19 $X=6.385 $Y=1.41 $X2=0 $Y2=0
cc_432 N_A_774_21#_c_572_n N_Q_c_890_n 0.00522013f $X=6.855 $Y=1.202 $X2=0 $Y2=0
cc_433 N_A_774_21#_c_575_n N_Q_c_885_n 0.00177605f $X=5.445 $Y=1.41 $X2=0 $Y2=0
cc_434 N_A_774_21#_c_576_n N_Q_c_885_n 0.00247675f $X=5.915 $Y=1.41 $X2=0 $Y2=0
cc_435 N_A_774_21#_c_577_n N_Q_c_885_n 2.75106e-19 $X=6.385 $Y=1.41 $X2=0 $Y2=0
cc_436 N_A_774_21#_c_572_n N_Q_c_885_n 0.00485245f $X=6.855 $Y=1.202 $X2=0 $Y2=0
cc_437 N_A_774_21#_c_571_n N_Q_c_898_n 0.0225433f $X=5.405 $Y=1.16 $X2=0 $Y2=0
cc_438 N_A_774_21#_c_572_n N_Q_c_898_n 0.0151066f $X=6.855 $Y=1.202 $X2=0 $Y2=0
cc_439 N_A_774_21#_c_567_n Q 0.00389878f $X=5.94 $Y=0.995 $X2=0 $Y2=0
cc_440 N_A_774_21#_c_568_n Q 6.37256e-19 $X=6.41 $Y=0.995 $X2=0 $Y2=0
cc_441 N_A_774_21#_c_572_n Q 0.00278736f $X=6.855 $Y=1.202 $X2=0 $Y2=0
cc_442 N_A_774_21#_c_576_n Q 0.0125305f $X=5.915 $Y=1.41 $X2=0 $Y2=0
cc_443 N_A_774_21#_c_568_n Q 0.0022241f $X=6.41 $Y=0.995 $X2=0 $Y2=0
cc_444 N_A_774_21#_c_569_n Q 0.00383003f $X=6.88 $Y=0.995 $X2=0 $Y2=0
cc_445 N_A_774_21#_c_577_n Q 0.00582467f $X=6.385 $Y=1.41 $X2=0 $Y2=0
cc_446 N_A_774_21#_c_578_n Q 0.0195168f $X=6.855 $Y=1.41 $X2=0 $Y2=0
cc_447 N_A_774_21#_c_572_n Q 0.00595439f $X=6.855 $Y=1.202 $X2=0 $Y2=0
cc_448 N_A_774_21#_c_572_n Q 0.017113f $X=6.855 $Y=1.202 $X2=0 $Y2=0
cc_449 N_A_774_21#_c_572_n N_Q_c_910_n 0.059537f $X=6.855 $Y=1.202 $X2=0 $Y2=0
cc_450 N_A_774_21#_c_572_n Q 0.025259f $X=6.855 $Y=1.202 $X2=0 $Y2=0
cc_451 N_A_774_21#_M1009_g N_VGND_c_932_n 0.00727714f $X=3.945 $Y=0.445 $X2=0
+ $Y2=0
cc_452 N_A_774_21#_c_570_n N_VGND_c_932_n 0.00790442f $X=4.755 $Y=0.58 $X2=0
+ $Y2=0
cc_453 N_A_774_21#_c_566_n N_VGND_c_933_n 0.00373785f $X=5.47 $Y=0.995 $X2=0
+ $Y2=0
cc_454 N_A_774_21#_c_571_n N_VGND_c_933_n 0.0147682f $X=5.405 $Y=1.16 $X2=0
+ $Y2=0
cc_455 N_A_774_21#_c_572_n N_VGND_c_933_n 0.00221294f $X=6.855 $Y=1.202 $X2=0
+ $Y2=0
cc_456 N_A_774_21#_c_567_n N_VGND_c_934_n 0.00382269f $X=5.94 $Y=0.995 $X2=0
+ $Y2=0
cc_457 N_A_774_21#_c_568_n N_VGND_c_934_n 0.00405678f $X=6.41 $Y=0.995 $X2=0
+ $Y2=0
cc_458 N_A_774_21#_c_572_n N_VGND_c_934_n 0.00326139f $X=6.855 $Y=1.202 $X2=0
+ $Y2=0
cc_459 N_A_774_21#_c_569_n N_VGND_c_936_n 0.0066844f $X=6.88 $Y=0.995 $X2=0
+ $Y2=0
cc_460 N_A_774_21#_M1009_g N_VGND_c_937_n 0.00475644f $X=3.945 $Y=0.445 $X2=0
+ $Y2=0
cc_461 N_A_774_21#_c_570_n N_VGND_c_941_n 0.00635207f $X=4.755 $Y=0.58 $X2=0
+ $Y2=0
cc_462 N_A_774_21#_c_566_n N_VGND_c_942_n 0.00585385f $X=5.47 $Y=0.995 $X2=0
+ $Y2=0
cc_463 N_A_774_21#_c_567_n N_VGND_c_942_n 0.00547395f $X=5.94 $Y=0.995 $X2=0
+ $Y2=0
cc_464 N_A_774_21#_c_568_n N_VGND_c_943_n 0.00585385f $X=6.41 $Y=0.995 $X2=0
+ $Y2=0
cc_465 N_A_774_21#_c_569_n N_VGND_c_943_n 0.00585385f $X=6.88 $Y=0.995 $X2=0
+ $Y2=0
cc_466 N_A_774_21#_M1014_s N_VGND_c_948_n 0.00691214f $X=4.6 $Y=0.235 $X2=0
+ $Y2=0
cc_467 N_A_774_21#_M1009_g N_VGND_c_948_n 0.00943411f $X=3.945 $Y=0.445 $X2=0
+ $Y2=0
cc_468 N_A_774_21#_c_566_n N_VGND_c_948_n 0.0109309f $X=5.47 $Y=0.995 $X2=0
+ $Y2=0
cc_469 N_A_774_21#_c_567_n N_VGND_c_948_n 0.00990847f $X=5.94 $Y=0.995 $X2=0
+ $Y2=0
cc_470 N_A_774_21#_c_568_n N_VGND_c_948_n 0.0108771f $X=6.41 $Y=0.995 $X2=0
+ $Y2=0
cc_471 N_A_774_21#_c_569_n N_VGND_c_948_n 0.0118212f $X=6.88 $Y=0.995 $X2=0
+ $Y2=0
cc_472 N_A_774_21#_c_570_n N_VGND_c_948_n 0.0066044f $X=4.755 $Y=0.58 $X2=0
+ $Y2=0
cc_473 N_A_609_413#_c_695_n N_VPWR_c_764_n 0.00465685f $X=3.78 $Y=2.34 $X2=0
+ $Y2=0
cc_474 N_A_609_413#_c_690_n N_VPWR_c_765_n 0.00308741f $X=4.96 $Y=1.41 $X2=0
+ $Y2=0
cc_475 N_A_609_413#_c_695_n N_VPWR_c_765_n 0.0133617f $X=3.78 $Y=2.34 $X2=0
+ $Y2=0
cc_476 N_A_609_413#_c_693_n N_VPWR_c_765_n 0.00839059f $X=3.865 $Y=2.255 $X2=0
+ $Y2=0
cc_477 N_A_609_413#_c_690_n N_VPWR_c_766_n 0.00419888f $X=4.96 $Y=1.41 $X2=0
+ $Y2=0
cc_478 N_A_609_413#_c_695_n N_VPWR_c_772_n 0.0417852f $X=3.78 $Y=2.34 $X2=0
+ $Y2=0
cc_479 N_A_609_413#_c_690_n N_VPWR_c_775_n 0.00702461f $X=4.96 $Y=1.41 $X2=0
+ $Y2=0
cc_480 N_A_609_413#_M1018_d N_VPWR_c_762_n 0.00233855f $X=3.045 $Y=2.065 $X2=0
+ $Y2=0
cc_481 N_A_609_413#_c_690_n N_VPWR_c_762_n 0.0139295f $X=4.96 $Y=1.41 $X2=0
+ $Y2=0
cc_482 N_A_609_413#_c_695_n N_VPWR_c_762_n 0.0324445f $X=3.78 $Y=2.34 $X2=0
+ $Y2=0
cc_483 N_A_609_413#_c_695_n A_703_413# 0.00873394f $X=3.78 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_484 N_A_609_413#_c_693_n A_703_413# 0.00235785f $X=3.865 $Y=2.255 $X2=-0.19
+ $Y2=-0.24
cc_485 N_A_609_413#_c_684_n N_VGND_c_932_n 0.00549625f $X=4.985 $Y=0.995 $X2=0
+ $Y2=0
cc_486 N_A_609_413#_c_697_n N_VGND_c_932_n 0.0133617f $X=3.78 $Y=0.45 $X2=0
+ $Y2=0
cc_487 N_A_609_413#_c_687_n N_VGND_c_932_n 0.00523144f $X=3.865 $Y=0.995 $X2=0
+ $Y2=0
cc_488 N_A_609_413#_c_688_n N_VGND_c_932_n 0.00808131f $X=4.415 $Y=1.16 $X2=0
+ $Y2=0
cc_489 N_A_609_413#_c_684_n N_VGND_c_933_n 0.0036647f $X=4.985 $Y=0.995 $X2=0
+ $Y2=0
cc_490 N_A_609_413#_c_697_n N_VGND_c_937_n 0.0284302f $X=3.78 $Y=0.45 $X2=0
+ $Y2=0
cc_491 N_A_609_413#_c_684_n N_VGND_c_941_n 0.00585385f $X=4.985 $Y=0.995 $X2=0
+ $Y2=0
cc_492 N_A_609_413#_M1008_d N_VGND_c_948_n 0.00237979f $X=3.115 $Y=0.235 $X2=0
+ $Y2=0
cc_493 N_A_609_413#_c_684_n N_VGND_c_948_n 0.0122012f $X=4.985 $Y=0.995 $X2=0
+ $Y2=0
cc_494 N_A_609_413#_c_697_n N_VGND_c_948_n 0.0288414f $X=3.78 $Y=0.45 $X2=0
+ $Y2=0
cc_495 N_A_609_413#_c_697_n A_709_47# 0.00922888f $X=3.78 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_496 N_A_609_413#_c_687_n A_709_47# 0.00144817f $X=3.865 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_497 N_VPWR_c_762_n A_503_369# 0.00402004f $X=7.13 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_498 N_VPWR_c_762_n A_703_413# 0.00296345f $X=7.13 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_499 N_VPWR_c_762_n N_Q_M1002_d 0.00439839f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_500 N_VPWR_c_762_n N_Q_M1020_d 0.00439839f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_501 N_VPWR_c_766_n N_Q_c_890_n 0.0599927f $X=5.21 $Y=1.735 $X2=0 $Y2=0
cc_502 N_VPWR_c_767_n N_Q_c_890_n 0.0723968f $X=6.15 $Y=1.835 $X2=0 $Y2=0
cc_503 N_VPWR_c_776_n Q 0.017659f $X=6.065 $Y=2.72 $X2=0 $Y2=0
cc_504 N_VPWR_c_762_n Q 0.0110326f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_505 N_VPWR_c_767_n Q 0.0589656f $X=6.15 $Y=1.835 $X2=0 $Y2=0
cc_506 N_VPWR_c_769_n Q 0.0615738f $X=7.09 $Y=1.835 $X2=0 $Y2=0
cc_507 N_VPWR_c_777_n Q 0.0157397f $X=7.005 $Y=2.72 $X2=0 $Y2=0
cc_508 N_VPWR_c_762_n Q 0.0100208f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_509 N_VPWR_c_767_n N_Q_c_910_n 0.0178695f $X=6.15 $Y=1.835 $X2=0 $Y2=0
cc_510 N_VPWR_c_769_n Q 0.0145641f $X=7.09 $Y=1.835 $X2=0 $Y2=0
cc_511 N_Q_c_910_n N_VGND_c_934_n 0.0185952f $X=6.535 $Y=1.16 $X2=0 $Y2=0
cc_512 Q N_VGND_c_936_n 0.00998619f $X=7.125 $Y=1.19 $X2=0 $Y2=0
cc_513 Q N_VGND_c_942_n 0.00897751f $X=5.645 $Y=0.425 $X2=0 $Y2=0
cc_514 Q N_VGND_c_943_n 0.0090872f $X=6.595 $Y=0.425 $X2=0 $Y2=0
cc_515 N_Q_M1003_d N_VGND_c_948_n 0.00457716f $X=5.545 $Y=0.235 $X2=0 $Y2=0
cc_516 N_Q_M1012_d N_VGND_c_948_n 0.0044972f $X=6.485 $Y=0.235 $X2=0 $Y2=0
cc_517 Q N_VGND_c_948_n 0.0102095f $X=5.645 $Y=0.425 $X2=0 $Y2=0
cc_518 Q N_VGND_c_948_n 0.00959809f $X=6.595 $Y=0.425 $X2=0 $Y2=0
cc_519 N_VGND_c_948_n A_505_47# 0.0145643f $X=7.13 $Y=0 $X2=-0.19 $Y2=-0.24
cc_520 N_VGND_c_948_n A_709_47# 0.00276161f $X=7.13 $Y=0 $X2=-0.19 $Y2=-0.24
