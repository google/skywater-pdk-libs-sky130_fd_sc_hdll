* File: sky130_fd_sc_hdll__mux2i_4.pxi.spice
* Created: Thu Aug 27 19:11:15 2020
* 
x_PM_SKY130_FD_SC_HDLL__MUX2I_4%A0 N_A0_c_106_n N_A0_M1010_g N_A0_c_111_n
+ N_A0_M1002_g N_A0_c_107_n N_A0_M1012_g N_A0_c_112_n N_A0_M1015_g N_A0_c_108_n
+ N_A0_M1025_g N_A0_c_113_n N_A0_M1022_g N_A0_c_114_n N_A0_M1030_g N_A0_c_109_n
+ N_A0_M1032_g A0 A0 N_A0_c_110_n A0 A0 PM_SKY130_FD_SC_HDLL__MUX2I_4%A0
x_PM_SKY130_FD_SC_HDLL__MUX2I_4%A1 N_A1_c_168_n N_A1_M1013_g N_A1_c_174_n
+ N_A1_M1000_g N_A1_c_169_n N_A1_M1019_g N_A1_c_175_n N_A1_M1007_g N_A1_c_170_n
+ N_A1_M1026_g N_A1_c_176_n N_A1_M1011_g N_A1_c_177_n N_A1_M1017_g N_A1_c_171_n
+ N_A1_M1027_g A1 A1 A1 A1 N_A1_c_172_n A1 A1 A1 A1
+ PM_SKY130_FD_SC_HDLL__MUX2I_4%A1
x_PM_SKY130_FD_SC_HDLL__MUX2I_4%S N_S_c_247_n N_S_M1005_g N_S_c_238_n
+ N_S_M1006_g N_S_c_248_n N_S_M1009_g N_S_c_239_n N_S_M1008_g N_S_c_249_n
+ N_S_M1020_g N_S_c_240_n N_S_M1016_g N_S_c_250_n N_S_M1031_g N_S_c_241_n
+ N_S_M1024_g N_S_c_242_n N_S_M1033_g N_S_c_243_n N_S_M1029_g N_S_c_252_n
+ N_S_c_244_n N_S_c_245_n S S S S S N_S_c_246_n S S S S S
+ PM_SKY130_FD_SC_HDLL__MUX2I_4%S
x_PM_SKY130_FD_SC_HDLL__MUX2I_4%A_1311_21# N_A_1311_21#_M1029_d
+ N_A_1311_21#_M1033_d N_A_1311_21#_c_370_n N_A_1311_21#_M1001_g
+ N_A_1311_21#_c_380_n N_A_1311_21#_M1003_g N_A_1311_21#_c_371_n
+ N_A_1311_21#_M1004_g N_A_1311_21#_c_381_n N_A_1311_21#_M1014_g
+ N_A_1311_21#_c_372_n N_A_1311_21#_M1021_g N_A_1311_21#_c_382_n
+ N_A_1311_21#_M1018_g N_A_1311_21#_c_383_n N_A_1311_21#_M1023_g
+ N_A_1311_21#_c_373_n N_A_1311_21#_M1028_g N_A_1311_21#_c_374_n
+ N_A_1311_21#_c_375_n N_A_1311_21#_c_404_n N_A_1311_21#_c_450_p
+ N_A_1311_21#_c_376_n N_A_1311_21#_c_384_n N_A_1311_21#_c_385_n
+ N_A_1311_21#_c_377_n N_A_1311_21#_c_378_n N_A_1311_21#_c_379_n
+ PM_SKY130_FD_SC_HDLL__MUX2I_4%A_1311_21#
x_PM_SKY130_FD_SC_HDLL__MUX2I_4%Y N_Y_M1010_s N_Y_M1012_s N_Y_M1032_s
+ N_Y_M1019_d N_Y_M1027_d N_Y_M1002_d N_Y_M1015_d N_Y_M1030_d N_Y_M1007_d
+ N_Y_M1017_d N_Y_c_484_n N_Y_c_487_n N_Y_c_485_n Y Y Y Y Y N_Y_c_489_n Y
+ PM_SKY130_FD_SC_HDLL__MUX2I_4%Y
x_PM_SKY130_FD_SC_HDLL__MUX2I_4%A_117_297# N_A_117_297#_M1002_s
+ N_A_117_297#_M1022_s N_A_117_297#_M1005_d N_A_117_297#_M1020_d
+ N_A_117_297#_c_556_n PM_SKY130_FD_SC_HDLL__MUX2I_4%A_117_297#
x_PM_SKY130_FD_SC_HDLL__MUX2I_4%A_493_297# N_A_493_297#_M1000_s
+ N_A_493_297#_M1011_s N_A_493_297#_M1003_s N_A_493_297#_M1018_s
+ N_A_493_297#_c_597_n N_A_493_297#_c_637_p N_A_493_297#_c_611_n
+ N_A_493_297#_c_612_n N_A_493_297#_c_618_n N_A_493_297#_c_613_n
+ PM_SKY130_FD_SC_HDLL__MUX2I_4%A_493_297#
x_PM_SKY130_FD_SC_HDLL__MUX2I_4%VPWR N_VPWR_M1005_s N_VPWR_M1009_s
+ N_VPWR_M1031_s N_VPWR_M1014_d N_VPWR_M1023_d N_VPWR_c_657_n N_VPWR_c_658_n
+ N_VPWR_c_659_n N_VPWR_c_660_n N_VPWR_c_661_n N_VPWR_c_662_n N_VPWR_c_663_n
+ N_VPWR_c_664_n N_VPWR_c_665_n N_VPWR_c_666_n VPWR N_VPWR_c_667_n
+ N_VPWR_c_656_n N_VPWR_c_669_n N_VPWR_c_670_n
+ PM_SKY130_FD_SC_HDLL__MUX2I_4%VPWR
x_PM_SKY130_FD_SC_HDLL__MUX2I_4%A_109_47# N_A_109_47#_M1010_d
+ N_A_109_47#_M1025_d N_A_109_47#_M1001_s N_A_109_47#_M1021_s
+ N_A_109_47#_c_811_n N_A_109_47#_c_773_n N_A_109_47#_c_774_n
+ N_A_109_47#_c_775_n N_A_109_47#_c_776_n N_A_109_47#_c_777_n
+ N_A_109_47#_c_778_n N_A_109_47#_c_788_n N_A_109_47#_c_779_n
+ PM_SKY130_FD_SC_HDLL__MUX2I_4%A_109_47#
x_PM_SKY130_FD_SC_HDLL__MUX2I_4%A_485_47# N_A_485_47#_M1013_s
+ N_A_485_47#_M1026_s N_A_485_47#_M1006_s N_A_485_47#_M1016_s
+ N_A_485_47#_c_867_n N_A_485_47#_c_878_n N_A_485_47#_c_879_n
+ N_A_485_47#_c_884_n N_A_485_47#_c_885_n
+ PM_SKY130_FD_SC_HDLL__MUX2I_4%A_485_47#
x_PM_SKY130_FD_SC_HDLL__MUX2I_4%VGND N_VGND_M1006_d N_VGND_M1008_d
+ N_VGND_M1024_d N_VGND_M1004_d N_VGND_M1028_d N_VGND_c_918_n N_VGND_c_919_n
+ N_VGND_c_920_n N_VGND_c_921_n N_VGND_c_922_n N_VGND_c_923_n N_VGND_c_924_n
+ N_VGND_c_925_n N_VGND_c_926_n N_VGND_c_927_n N_VGND_c_928_n N_VGND_c_929_n
+ VGND N_VGND_c_930_n N_VGND_c_931_n N_VGND_c_932_n N_VGND_c_933_n
+ PM_SKY130_FD_SC_HDLL__MUX2I_4%VGND
cc_1 VNB N_A0_c_106_n 0.0196633f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A0_c_107_n 0.016964f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_3 VNB N_A0_c_108_n 0.0171836f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_4 VNB N_A0_c_109_n 0.0166592f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_5 VNB N_A0_c_110_n 0.07794f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_6 VNB N_A1_c_168_n 0.0164026f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_7 VNB N_A1_c_169_n 0.0166886f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_8 VNB N_A1_c_170_n 0.0171301f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_9 VNB N_A1_c_171_n 0.0222991f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_10 VNB N_A1_c_172_n 0.0766807f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.16
cc_11 VNB A1 0.00395037f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_S_c_238_n 0.0218576f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_13 VNB N_S_c_239_n 0.0161794f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_14 VNB N_S_c_240_n 0.0166886f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_15 VNB N_S_c_241_n 0.0158516f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_16 VNB N_S_c_242_n 0.0275122f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_17 VNB N_S_c_243_n 0.0202819f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_S_c_244_n 9.74523e-19 $X=-0.19 $Y=-0.24 $X2=1.035 $Y2=1.16
cc_19 VNB N_S_c_245_n 0.0116739f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.202
cc_20 VNB N_S_c_246_n 0.092385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_1311_21#_c_370_n 0.0159768f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_22 VNB N_A_1311_21#_c_371_n 0.0165154f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_23 VNB N_A_1311_21#_c_372_n 0.0175938f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_24 VNB N_A_1311_21#_c_373_n 0.0177677f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_1311_21#_c_374_n 0.00188285f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.202
cc_26 VNB N_A_1311_21#_c_375_n 0.00142015f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.202
cc_27 VNB N_A_1311_21#_c_376_n 0.0155218f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.16
cc_28 VNB N_A_1311_21#_c_377_n 0.00723806f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_1311_21#_c_378_n 0.0219794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_1311_21#_c_379_n 0.0783619f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_Y_c_484_n 0.00233266f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.202
cc_32 VNB N_Y_c_485_n 0.00749881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB Y 0.0362988f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_656_n 0.383598f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_109_47#_c_773_n 0.00444967f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_36 VNB N_A_109_47#_c_774_n 0.00118342f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_37 VNB N_A_109_47#_c_775_n 0.0355593f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_109_47#_c_776_n 0.00331514f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.202
cc_39 VNB N_A_109_47#_c_777_n 0.00329117f $X=-0.19 $Y=-0.24 $X2=1.035 $Y2=1.16
cc_40 VNB N_A_109_47#_c_778_n 0.00496916f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.202
cc_41 VNB N_A_109_47#_c_779_n 0.00247078f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.16
cc_42 VNB N_A_485_47#_c_867_n 0.0069465f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_43 VNB N_VGND_c_918_n 0.0078084f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_44 VNB N_VGND_c_919_n 0.0134688f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_45 VNB N_VGND_c_920_n 0.0142091f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_46 VNB N_VGND_c_921_n 3.35731e-19 $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.105
cc_47 VNB N_VGND_c_922_n 0.00464512f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_48 VNB N_VGND_c_923_n 0.00561497f $X=-0.19 $Y=-0.24 $X2=1.035 $Y2=1.16
cc_49 VNB N_VGND_c_924_n 0.106403f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=1.202
cc_50 VNB N_VGND_c_925_n 0.00631443f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.202
cc_51 VNB N_VGND_c_926_n 0.0173881f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.202
cc_52 VNB N_VGND_c_927_n 0.00478085f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.16
cc_53 VNB N_VGND_c_928_n 0.0209545f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.16
cc_54 VNB N_VGND_c_929_n 0.00631443f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_55 VNB N_VGND_c_930_n 0.0189752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_931_n 0.433396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_932_n 0.00781014f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_933_n 0.00496766f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VPB N_A0_c_111_n 0.019155f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_60 VPB N_A0_c_112_n 0.0162614f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_61 VPB N_A0_c_113_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_62 VPB N_A0_c_114_n 0.016445f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_63 VPB N_A0_c_110_n 0.0473912f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_64 VPB N_A1_c_174_n 0.016445f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_65 VPB N_A1_c_175_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_66 VPB N_A1_c_176_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_67 VPB N_A1_c_177_n 0.0210879f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_68 VPB N_A1_c_172_n 0.0492565f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.16
cc_69 VPB A1 0.00201667f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_S_c_247_n 0.0202445f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_71 VPB N_S_c_248_n 0.0158129f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.995
cc_72 VPB N_S_c_249_n 0.01609f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=0.995
cc_73 VPB N_S_c_250_n 0.0159251f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_74 VPB N_S_c_242_n 0.0298017f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_75 VPB N_S_c_252_n 0.0101694f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.202
cc_76 VPB N_S_c_244_n 0.00102033f $X=-0.19 $Y=1.305 $X2=1.035 $Y2=1.16
cc_77 VPB N_S_c_245_n 0.00286228f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=1.202
cc_78 VPB N_S_c_246_n 0.0573763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_1311_21#_c_380_n 0.0155843f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_80 VPB N_A_1311_21#_c_381_n 0.0152727f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_81 VPB N_A_1311_21#_c_382_n 0.015982f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.995
cc_82 VPB N_A_1311_21#_c_383_n 0.0165514f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_83 VPB N_A_1311_21#_c_384_n 0.00494099f $X=-0.19 $Y=1.305 $X2=1.035 $Y2=1.16
cc_84 VPB N_A_1311_21#_c_385_n 0.0208429f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.16
cc_85 VPB N_A_1311_21#_c_378_n 0.019721f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_1311_21#_c_379_n 0.0467262f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_Y_c_487_n 0.00219582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB Y 0.0379835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_Y_c_489_n 0.00747992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_117_297#_c_556_n 0.00939914f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_91 VPB N_A_493_297#_c_597_n 0.00721458f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=0.995
cc_92 VPB N_VPWR_c_657_n 0.00558805f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_93 VPB N_VPWR_c_658_n 0.0132054f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_94 VPB N_VPWR_c_659_n 0.0132269f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.995
cc_95 VPB N_VPWR_c_660_n 0.00285945f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.105
cc_96 VPB N_VPWR_c_661_n 0.104999f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_662_n 0.00513086f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.202
cc_98 VPB N_VPWR_c_663_n 0.00547281f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.202
cc_99 VPB N_VPWR_c_664_n 0.0123761f $X=-0.19 $Y=1.305 $X2=1.035 $Y2=1.16
cc_100 VPB N_VPWR_c_665_n 0.0189384f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_101 VPB N_VPWR_c_666_n 0.00513086f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=1.202
cc_102 VPB N_VPWR_c_667_n 0.0188763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_656_n 0.0501609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_669_n 0.00537041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_670_n 0.00537882f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 N_A0_c_109_n N_A1_c_168_n 0.0253282f $X=1.93 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_107 N_A0_c_114_n N_A1_c_174_n 0.041284f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A0_c_110_n N_A1_c_172_n 0.0253282f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_109 N_A0_c_110_n A1 0.00206219f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_110 N_A0_c_106_n N_Y_c_484_n 0.0119518f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A0_c_107_n N_Y_c_484_n 0.00831741f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A0_c_108_n N_Y_c_484_n 0.00857637f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A0_c_109_n N_Y_c_484_n 0.0091452f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A0_c_111_n N_Y_c_487_n 0.0133352f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A0_c_112_n N_Y_c_487_n 0.0112427f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A0_c_113_n N_Y_c_487_n 0.0112427f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A0_c_114_n N_Y_c_487_n 0.0112427f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A0_c_106_n Y 0.0287485f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A0_c_111_n Y 0.0284248f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_120 A0 Y 0.018802f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_121 N_A0_c_111_n N_A_117_297#_c_556_n 0.0073309f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A0_c_112_n N_A_117_297#_c_556_n 0.0123901f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A0_c_113_n N_A_117_297#_c_556_n 0.0161919f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A0_c_114_n N_A_117_297#_c_556_n 0.0154983f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A0_c_110_n N_A_117_297#_c_556_n 0.0189547f $X=1.905 $Y=1.202 $X2=0
+ $Y2=0
cc_126 A0 N_A_117_297#_c_556_n 0.0304133f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_127 N_A0_c_114_n N_A_493_297#_c_597_n 8.47478e-19 $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_128 N_A0_c_111_n N_VPWR_c_661_n 0.00439333f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A0_c_112_n N_VPWR_c_661_n 0.00439333f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A0_c_113_n N_VPWR_c_661_n 0.00439333f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A0_c_114_n N_VPWR_c_661_n 0.00439333f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A0_c_111_n N_VPWR_c_656_n 0.00699435f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A0_c_112_n N_VPWR_c_656_n 0.00608292f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A0_c_113_n N_VPWR_c_656_n 0.00608292f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A0_c_114_n N_VPWR_c_656_n 0.00610813f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A0_c_109_n N_A_109_47#_c_775_n 0.00598557f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A0_c_108_n N_A_109_47#_c_776_n 5.03517e-19 $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A0_c_109_n N_A_109_47#_c_776_n 0.00299356f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A0_c_110_n N_A_109_47#_c_776_n 0.00407598f $X=1.905 $Y=1.202 $X2=0
+ $Y2=0
cc_140 N_A0_c_107_n N_A_109_47#_c_778_n 5.26678e-19 $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A0_c_108_n N_A_109_47#_c_778_n 0.00451504f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A0_c_109_n N_A_109_47#_c_778_n 0.00225375f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A0_c_110_n N_A_109_47#_c_778_n 0.00586298f $X=1.905 $Y=1.202 $X2=0
+ $Y2=0
cc_144 N_A0_c_106_n N_A_109_47#_c_788_n 0.00363882f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A0_c_107_n N_A_109_47#_c_788_n 0.00865599f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A0_c_108_n N_A_109_47#_c_788_n 0.01098f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A0_c_110_n N_A_109_47#_c_788_n 0.00642921f $X=1.905 $Y=1.202 $X2=0
+ $Y2=0
cc_148 A0 N_A_109_47#_c_788_n 0.042652f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_149 N_A0_c_109_n N_A_485_47#_c_867_n 5.23135e-19 $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A0_c_106_n N_VGND_c_924_n 0.00370116f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A0_c_107_n N_VGND_c_924_n 0.00370116f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A0_c_108_n N_VGND_c_924_n 0.00370116f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A0_c_109_n N_VGND_c_924_n 0.00370116f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A0_c_106_n N_VGND_c_931_n 0.00633963f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A0_c_107_n N_VGND_c_931_n 0.00551239f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A0_c_108_n N_VGND_c_931_n 0.00563217f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A0_c_109_n N_VGND_c_931_n 0.00545403f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A1_c_172_n N_S_c_245_n 6.88572e-19 $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_159 A1 N_S_c_245_n 0.0181001f $X=3.925 $Y=1.19 $X2=0 $Y2=0
cc_160 N_A1_c_172_n N_S_c_246_n 0.00647224f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_161 A1 N_S_c_246_n 0.00370997f $X=3.925 $Y=1.19 $X2=0 $Y2=0
cc_162 N_A1_c_168_n N_Y_c_484_n 0.00902847f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A1_c_169_n N_Y_c_484_n 0.00827443f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A1_c_170_n N_Y_c_484_n 0.00853339f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A1_c_171_n N_Y_c_484_n 0.00853339f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_166 A1 N_Y_c_484_n 5.12982e-19 $X=3.925 $Y=1.19 $X2=0 $Y2=0
cc_167 N_A1_c_174_n N_Y_c_487_n 0.0104486f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A1_c_175_n N_Y_c_487_n 0.0092122f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A1_c_176_n N_Y_c_487_n 0.0092122f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A1_c_177_n N_Y_c_487_n 0.0092122f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A1_c_174_n N_A_117_297#_c_556_n 0.0155969f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A1_c_175_n N_A_117_297#_c_556_n 0.0124734f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A1_c_176_n N_A_117_297#_c_556_n 0.0124734f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A1_c_177_n N_A_117_297#_c_556_n 0.0144732f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A1_c_172_n N_A_117_297#_c_556_n 0.0176759f $X=3.785 $Y=1.202 $X2=0
+ $Y2=0
cc_176 A1 N_A_117_297#_c_556_n 0.0812793f $X=3.925 $Y=1.19 $X2=0 $Y2=0
cc_177 N_A1_c_174_n N_A_493_297#_c_597_n 0.00588483f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_178 N_A1_c_175_n N_A_493_297#_c_597_n 0.00977137f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_179 N_A1_c_176_n N_A_493_297#_c_597_n 0.00977137f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_180 N_A1_c_177_n N_A_493_297#_c_597_n 0.0117712f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A1_c_177_n N_VPWR_c_657_n 0.00291855f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A1_c_174_n N_VPWR_c_661_n 0.00439333f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A1_c_175_n N_VPWR_c_661_n 0.00439333f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A1_c_176_n N_VPWR_c_661_n 0.00439333f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A1_c_177_n N_VPWR_c_661_n 0.00439333f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_186 N_A1_c_174_n N_VPWR_c_656_n 0.00610813f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_187 N_A1_c_175_n N_VPWR_c_656_n 0.00608292f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A1_c_176_n N_VPWR_c_656_n 0.00608292f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A1_c_177_n N_VPWR_c_656_n 0.00736527f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_190 N_A1_c_168_n N_A_109_47#_c_775_n 0.00627598f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A1_c_169_n N_A_109_47#_c_775_n 0.00212165f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A1_c_170_n N_A_109_47#_c_775_n 0.00215271f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A1_c_171_n N_A_109_47#_c_775_n 0.00301975f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A1_c_172_n N_A_109_47#_c_775_n 0.0120003f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_195 A1 N_A_109_47#_c_775_n 0.045905f $X=3.925 $Y=1.19 $X2=0 $Y2=0
cc_196 N_A1_c_168_n N_A_109_47#_c_776_n 4.23023e-19 $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A1_c_168_n N_A_485_47#_c_867_n 0.00342584f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A1_c_169_n N_A_485_47#_c_867_n 0.0077424f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A1_c_170_n N_A_485_47#_c_867_n 0.0077424f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A1_c_171_n N_A_485_47#_c_867_n 0.00954923f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A1_c_172_n N_A_485_47#_c_867_n 0.0103179f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_202 A1 N_A_485_47#_c_867_n 0.0985243f $X=3.925 $Y=1.19 $X2=0 $Y2=0
cc_203 N_A1_c_171_n N_VGND_c_918_n 0.00323055f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A1_c_168_n N_VGND_c_924_n 0.00370116f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A1_c_169_n N_VGND_c_924_n 0.00370116f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A1_c_170_n N_VGND_c_924_n 0.00370116f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A1_c_171_n N_VGND_c_924_n 0.00370116f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A1_c_168_n N_VGND_c_931_n 0.00535232f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A1_c_169_n N_VGND_c_931_n 0.00545208f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A1_c_170_n N_VGND_c_931_n 0.00557186f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A1_c_171_n N_VGND_c_931_n 0.00677096f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_212 N_S_c_241_n N_A_1311_21#_c_370_n 0.0223656f $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_213 N_S_c_250_n N_A_1311_21#_c_380_n 0.0376944f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_214 N_S_c_252_n N_A_1311_21#_c_380_n 0.0130584f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_215 N_S_c_245_n N_A_1311_21#_c_380_n 8.1953e-19 $X=6.36 $Y=1.182 $X2=0 $Y2=0
cc_216 N_S_c_252_n N_A_1311_21#_c_381_n 0.0149152f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_217 N_S_c_252_n N_A_1311_21#_c_382_n 0.0133014f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_218 N_S_c_242_n N_A_1311_21#_c_383_n 0.0322661f $X=8.635 $Y=1.41 $X2=0 $Y2=0
cc_219 N_S_c_252_n N_A_1311_21#_c_383_n 0.0179858f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_220 N_S_c_244_n N_A_1311_21#_c_383_n 2.65369e-19 $X=8.565 $Y=1.16 $X2=0 $Y2=0
cc_221 N_S_c_243_n N_A_1311_21#_c_373_n 0.0176195f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_222 N_S_c_242_n N_A_1311_21#_c_374_n 0.00114887f $X=8.635 $Y=1.41 $X2=0 $Y2=0
cc_223 N_S_c_252_n N_A_1311_21#_c_374_n 0.0608377f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_224 N_S_c_244_n N_A_1311_21#_c_374_n 0.0137152f $X=8.565 $Y=1.16 $X2=0 $Y2=0
cc_225 N_S_c_242_n N_A_1311_21#_c_375_n 4.73878e-19 $X=8.635 $Y=1.41 $X2=0 $Y2=0
cc_226 N_S_c_243_n N_A_1311_21#_c_375_n 0.00150278f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_227 N_S_c_244_n N_A_1311_21#_c_375_n 0.00580268f $X=8.565 $Y=1.16 $X2=0 $Y2=0
cc_228 N_S_c_242_n N_A_1311_21#_c_404_n 0.00198062f $X=8.635 $Y=1.41 $X2=0 $Y2=0
cc_229 N_S_c_243_n N_A_1311_21#_c_404_n 0.0163692f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_230 N_S_c_252_n N_A_1311_21#_c_404_n 0.00502258f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_231 N_S_c_244_n N_A_1311_21#_c_404_n 0.0108369f $X=8.565 $Y=1.16 $X2=0 $Y2=0
cc_232 N_S_c_242_n N_A_1311_21#_c_378_n 0.0203828f $X=8.635 $Y=1.41 $X2=0 $Y2=0
cc_233 N_S_c_243_n N_A_1311_21#_c_378_n 0.00409123f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_234 N_S_c_252_n N_A_1311_21#_c_378_n 0.0110463f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_235 N_S_c_244_n N_A_1311_21#_c_378_n 0.0253668f $X=8.565 $Y=1.16 $X2=0 $Y2=0
cc_236 N_S_c_242_n N_A_1311_21#_c_379_n 0.0243722f $X=8.635 $Y=1.41 $X2=0 $Y2=0
cc_237 N_S_c_252_n N_A_1311_21#_c_379_n 0.0279865f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_238 N_S_c_244_n N_A_1311_21#_c_379_n 0.00241591f $X=8.565 $Y=1.16 $X2=0 $Y2=0
cc_239 N_S_c_245_n N_A_1311_21#_c_379_n 0.00875208f $X=6.36 $Y=1.182 $X2=0 $Y2=0
cc_240 N_S_c_246_n N_A_1311_21#_c_379_n 0.0223656f $X=6.185 $Y=1.202 $X2=0 $Y2=0
cc_241 N_S_c_247_n N_A_117_297#_c_556_n 0.012587f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_242 N_S_c_248_n N_A_117_297#_c_556_n 0.0105872f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_243 N_S_c_249_n N_A_117_297#_c_556_n 0.0105872f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_244 N_S_c_250_n N_A_117_297#_c_556_n 0.00449112f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_245 N_S_c_245_n N_A_117_297#_c_556_n 0.0812614f $X=6.36 $Y=1.182 $X2=0 $Y2=0
cc_246 N_S_c_246_n N_A_117_297#_c_556_n 0.0240387f $X=6.185 $Y=1.202 $X2=0 $Y2=0
cc_247 N_S_c_252_n N_A_493_297#_M1003_s 0.00193761f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_248 N_S_c_252_n N_A_493_297#_M1018_s 0.00415063f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_249 N_S_c_247_n N_A_493_297#_c_597_n 0.0153636f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_250 N_S_c_248_n N_A_493_297#_c_597_n 0.0128942f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_251 N_S_c_249_n N_A_493_297#_c_597_n 0.0133638f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_252 N_S_c_250_n N_A_493_297#_c_597_n 0.0149083f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_253 N_S_c_252_n N_A_493_297#_c_597_n 0.00740135f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_254 N_S_c_245_n N_A_493_297#_c_597_n 0.0124166f $X=6.36 $Y=1.182 $X2=0 $Y2=0
cc_255 N_S_c_252_n N_A_493_297#_c_611_n 0.0226965f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_256 N_S_c_252_n N_A_493_297#_c_612_n 0.0122384f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_257 N_S_c_252_n N_A_493_297#_c_613_n 0.0122384f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_258 N_S_c_245_n N_VPWR_M1031_s 0.00350501f $X=6.36 $Y=1.182 $X2=0 $Y2=0
cc_259 N_S_c_252_n N_VPWR_M1014_d 0.00251566f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_260 N_S_c_252_n N_VPWR_M1023_d 0.00458846f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_261 N_S_c_247_n N_VPWR_c_657_n 0.00923392f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_262 N_S_c_248_n N_VPWR_c_657_n 0.00106266f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_263 N_S_c_247_n N_VPWR_c_658_n 0.00452725f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_264 N_S_c_248_n N_VPWR_c_658_n 0.00311736f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_265 N_S_c_249_n N_VPWR_c_659_n 0.00453434f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_266 N_S_c_250_n N_VPWR_c_659_n 0.00311736f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_267 N_S_c_242_n N_VPWR_c_660_n 0.00857191f $X=8.635 $Y=1.41 $X2=0 $Y2=0
cc_268 N_S_c_252_n N_VPWR_c_660_n 0.00684744f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_269 N_S_c_242_n N_VPWR_c_667_n 0.00622633f $X=8.635 $Y=1.41 $X2=0 $Y2=0
cc_270 N_S_c_247_n N_VPWR_c_656_n 0.00518249f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_271 N_S_c_248_n N_VPWR_c_656_n 0.00375605f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_272 N_S_c_249_n N_VPWR_c_656_n 0.00518254f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_273 N_S_c_250_n N_VPWR_c_656_n 0.00375605f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_274 N_S_c_242_n N_VPWR_c_656_n 0.0113715f $X=8.635 $Y=1.41 $X2=0 $Y2=0
cc_275 N_S_c_247_n N_VPWR_c_669_n 0.00118604f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_276 N_S_c_248_n N_VPWR_c_669_n 0.011082f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_277 N_S_c_249_n N_VPWR_c_669_n 0.00820729f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_278 N_S_c_250_n N_VPWR_c_669_n 0.00106505f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_279 N_S_c_249_n N_VPWR_c_670_n 0.00118604f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_280 N_S_c_250_n N_VPWR_c_670_n 0.0110489f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_281 N_S_c_252_n N_A_109_47#_c_773_n 0.0107545f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_282 N_S_c_238_n N_A_109_47#_c_775_n 0.00347579f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_283 N_S_c_239_n N_A_109_47#_c_775_n 0.00260874f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_284 N_S_c_240_n N_A_109_47#_c_775_n 0.00260874f $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_285 N_S_c_241_n N_A_109_47#_c_775_n 0.00598499f $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_286 N_S_c_252_n N_A_109_47#_c_775_n 0.00437043f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_287 N_S_c_245_n N_A_109_47#_c_775_n 0.0625972f $X=6.36 $Y=1.182 $X2=0 $Y2=0
cc_288 N_S_c_246_n N_A_109_47#_c_775_n 0.019445f $X=6.185 $Y=1.202 $X2=0 $Y2=0
cc_289 N_S_c_241_n N_A_109_47#_c_777_n 4.06927e-19 $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_290 N_S_c_252_n N_A_109_47#_c_777_n 0.00902051f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_291 N_S_c_252_n N_A_109_47#_c_779_n 0.0071147f $X=8.48 $Y=1.51 $X2=0 $Y2=0
cc_292 N_S_c_238_n N_A_485_47#_c_867_n 0.0138196f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_293 N_S_c_245_n N_A_485_47#_c_867_n 0.0266009f $X=6.36 $Y=1.182 $X2=0 $Y2=0
cc_294 N_S_c_246_n N_A_485_47#_c_867_n 0.00769628f $X=6.185 $Y=1.202 $X2=0 $Y2=0
cc_295 N_S_c_239_n N_A_485_47#_c_878_n 0.00423992f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_296 N_S_c_239_n N_A_485_47#_c_879_n 0.0112105f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_297 N_S_c_240_n N_A_485_47#_c_879_n 0.0114317f $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_298 N_S_c_241_n N_A_485_47#_c_879_n 0.00479851f $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_299 N_S_c_245_n N_A_485_47#_c_879_n 0.0350088f $X=6.36 $Y=1.182 $X2=0 $Y2=0
cc_300 N_S_c_246_n N_A_485_47#_c_879_n 0.00640214f $X=6.185 $Y=1.202 $X2=0 $Y2=0
cc_301 N_S_c_241_n N_A_485_47#_c_884_n 0.00221725f $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_302 N_S_c_245_n N_A_485_47#_c_885_n 0.00692589f $X=6.36 $Y=1.182 $X2=0 $Y2=0
cc_303 N_S_c_246_n N_A_485_47#_c_885_n 0.00300262f $X=6.185 $Y=1.202 $X2=0 $Y2=0
cc_304 N_S_c_238_n N_VGND_c_918_n 0.00330805f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_305 N_S_c_238_n N_VGND_c_919_n 0.00428022f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_306 N_S_c_239_n N_VGND_c_919_n 0.00199743f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_307 N_S_c_240_n N_VGND_c_920_n 0.00428022f $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_308 N_S_c_241_n N_VGND_c_920_n 0.00271402f $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_309 N_S_c_240_n N_VGND_c_921_n 6.00933e-19 $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_310 N_S_c_241_n N_VGND_c_921_n 0.0120654f $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_311 N_S_c_245_n N_VGND_c_921_n 0.0048265f $X=6.36 $Y=1.182 $X2=0 $Y2=0
cc_312 N_S_c_243_n N_VGND_c_923_n 0.00319783f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_313 N_S_c_243_n N_VGND_c_930_n 0.00428022f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_314 N_S_c_238_n N_VGND_c_931_n 0.00680412f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_315 N_S_c_239_n N_VGND_c_931_n 0.00260317f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_316 N_S_c_240_n N_VGND_c_931_n 0.00560507f $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_317 N_S_c_241_n N_VGND_c_931_n 0.00297927f $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_318 N_S_c_243_n N_VGND_c_931_n 0.00689881f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_319 N_S_c_238_n N_VGND_c_932_n 5.64511e-19 $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_320 N_S_c_239_n N_VGND_c_932_n 0.00964409f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_321 N_S_c_240_n N_VGND_c_932_n 0.00162962f $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_322 N_A_1311_21#_c_380_n N_A_117_297#_c_556_n 7.07233e-19 $X=6.655 $Y=1.41
+ $X2=0 $Y2=0
cc_323 N_A_1311_21#_c_380_n N_A_493_297#_c_597_n 0.0122063f $X=6.655 $Y=1.41
+ $X2=0 $Y2=0
cc_324 N_A_1311_21#_c_381_n N_A_493_297#_c_611_n 0.0117368f $X=7.125 $Y=1.41
+ $X2=0 $Y2=0
cc_325 N_A_1311_21#_c_382_n N_A_493_297#_c_611_n 0.0122494f $X=7.595 $Y=1.41
+ $X2=0 $Y2=0
cc_326 N_A_1311_21#_c_383_n N_A_493_297#_c_612_n 0.00793745f $X=8.12 $Y=1.41
+ $X2=0 $Y2=0
cc_327 N_A_1311_21#_c_383_n N_A_493_297#_c_618_n 0.00578962f $X=8.12 $Y=1.41
+ $X2=0 $Y2=0
cc_328 N_A_1311_21#_c_383_n N_VPWR_c_660_n 0.00313517f $X=8.12 $Y=1.41 $X2=0
+ $Y2=0
cc_329 N_A_1311_21#_c_385_n N_VPWR_c_660_n 0.0131278f $X=8.87 $Y=1.96 $X2=0
+ $Y2=0
cc_330 N_A_1311_21#_c_380_n N_VPWR_c_663_n 5.36535e-19 $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_331 N_A_1311_21#_c_381_n N_VPWR_c_663_n 0.00943288f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_332 N_A_1311_21#_c_382_n N_VPWR_c_663_n 0.00788671f $X=7.595 $Y=1.41 $X2=0
+ $Y2=0
cc_333 N_A_1311_21#_c_383_n N_VPWR_c_663_n 0.00103264f $X=8.12 $Y=1.41 $X2=0
+ $Y2=0
cc_334 N_A_1311_21#_c_380_n N_VPWR_c_664_n 0.00453434f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_335 N_A_1311_21#_c_381_n N_VPWR_c_664_n 0.00311736f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_336 N_A_1311_21#_c_382_n N_VPWR_c_665_n 0.00453434f $X=7.595 $Y=1.41 $X2=0
+ $Y2=0
cc_337 N_A_1311_21#_c_383_n N_VPWR_c_665_n 0.00702461f $X=8.12 $Y=1.41 $X2=0
+ $Y2=0
cc_338 N_A_1311_21#_c_385_n N_VPWR_c_667_n 0.0182037f $X=8.87 $Y=1.96 $X2=0
+ $Y2=0
cc_339 N_A_1311_21#_M1033_d N_VPWR_c_656_n 0.00425811f $X=8.725 $Y=1.485 $X2=0
+ $Y2=0
cc_340 N_A_1311_21#_c_380_n N_VPWR_c_656_n 0.00513756f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_341 N_A_1311_21#_c_381_n N_VPWR_c_656_n 0.00371107f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_342 N_A_1311_21#_c_382_n N_VPWR_c_656_n 0.00527133f $X=7.595 $Y=1.41 $X2=0
+ $Y2=0
cc_343 N_A_1311_21#_c_383_n N_VPWR_c_656_n 0.012767f $X=8.12 $Y=1.41 $X2=0 $Y2=0
cc_344 N_A_1311_21#_c_385_n N_VPWR_c_656_n 0.00993477f $X=8.87 $Y=1.96 $X2=0
+ $Y2=0
cc_345 N_A_1311_21#_c_380_n N_VPWR_c_670_n 0.00675973f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_346 N_A_1311_21#_c_381_n N_VPWR_c_670_n 4.88209e-19 $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_347 N_A_1311_21#_c_370_n N_A_109_47#_c_811_n 0.00389287f $X=6.63 $Y=0.995
+ $X2=0 $Y2=0
cc_348 N_A_1311_21#_c_371_n N_A_109_47#_c_773_n 0.00749341f $X=7.1 $Y=0.995
+ $X2=0 $Y2=0
cc_349 N_A_1311_21#_c_372_n N_A_109_47#_c_773_n 0.0111949f $X=7.57 $Y=0.995
+ $X2=0 $Y2=0
cc_350 N_A_1311_21#_c_374_n N_A_109_47#_c_773_n 0.0221647f $X=8.09 $Y=1.16 $X2=0
+ $Y2=0
cc_351 N_A_1311_21#_c_379_n N_A_109_47#_c_773_n 0.00431283f $X=8.12 $Y=1.202
+ $X2=0 $Y2=0
cc_352 N_A_1311_21#_c_373_n N_A_109_47#_c_774_n 0.00508525f $X=8.145 $Y=0.995
+ $X2=0 $Y2=0
cc_353 N_A_1311_21#_c_374_n N_A_109_47#_c_774_n 0.012939f $X=8.09 $Y=1.16 $X2=0
+ $Y2=0
cc_354 N_A_1311_21#_c_375_n N_A_109_47#_c_774_n 0.00559134f $X=8.2 $Y=1.075
+ $X2=0 $Y2=0
cc_355 N_A_1311_21#_c_450_p N_A_109_47#_c_774_n 0.0130631f $X=8.31 $Y=0.74 $X2=0
+ $Y2=0
cc_356 N_A_1311_21#_c_379_n N_A_109_47#_c_774_n 0.00423644f $X=8.12 $Y=1.202
+ $X2=0 $Y2=0
cc_357 N_A_1311_21#_c_370_n N_A_109_47#_c_775_n 0.00551547f $X=6.63 $Y=0.995
+ $X2=0 $Y2=0
cc_358 N_A_1311_21#_c_370_n N_A_109_47#_c_777_n 0.00372235f $X=6.63 $Y=0.995
+ $X2=0 $Y2=0
cc_359 N_A_1311_21#_c_371_n N_A_109_47#_c_777_n 8.34829e-19 $X=7.1 $Y=0.995
+ $X2=0 $Y2=0
cc_360 N_A_1311_21#_c_379_n N_A_109_47#_c_777_n 0.00393542f $X=8.12 $Y=1.202
+ $X2=0 $Y2=0
cc_361 N_A_1311_21#_c_370_n N_A_109_47#_c_779_n 0.00496768f $X=6.63 $Y=0.995
+ $X2=0 $Y2=0
cc_362 N_A_1311_21#_c_371_n N_A_109_47#_c_779_n 0.00785442f $X=7.1 $Y=0.995
+ $X2=0 $Y2=0
cc_363 N_A_1311_21#_c_379_n N_A_109_47#_c_779_n 0.00389072f $X=8.12 $Y=1.202
+ $X2=0 $Y2=0
cc_364 N_A_1311_21#_c_375_n N_VGND_M1028_d 7.9502e-19 $X=8.2 $Y=1.075 $X2=0
+ $Y2=0
cc_365 N_A_1311_21#_c_404_n N_VGND_M1028_d 0.0058436f $X=8.785 $Y=0.74 $X2=0
+ $Y2=0
cc_366 N_A_1311_21#_c_450_p N_VGND_M1028_d 3.67444e-19 $X=8.31 $Y=0.74 $X2=0
+ $Y2=0
cc_367 N_A_1311_21#_c_370_n N_VGND_c_921_n 0.00844855f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_368 N_A_1311_21#_c_371_n N_VGND_c_921_n 5.83912e-19 $X=7.1 $Y=0.995 $X2=0
+ $Y2=0
cc_369 N_A_1311_21#_c_371_n N_VGND_c_922_n 0.0029572f $X=7.1 $Y=0.995 $X2=0
+ $Y2=0
cc_370 N_A_1311_21#_c_372_n N_VGND_c_922_n 0.0031255f $X=7.57 $Y=0.995 $X2=0
+ $Y2=0
cc_371 N_A_1311_21#_c_373_n N_VGND_c_923_n 0.00322931f $X=8.145 $Y=0.995 $X2=0
+ $Y2=0
cc_372 N_A_1311_21#_c_404_n N_VGND_c_923_n 0.0151325f $X=8.785 $Y=0.74 $X2=0
+ $Y2=0
cc_373 N_A_1311_21#_c_450_p N_VGND_c_923_n 0.00250582f $X=8.31 $Y=0.74 $X2=0
+ $Y2=0
cc_374 N_A_1311_21#_c_370_n N_VGND_c_926_n 0.00486043f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_375 N_A_1311_21#_c_371_n N_VGND_c_926_n 0.00436487f $X=7.1 $Y=0.995 $X2=0
+ $Y2=0
cc_376 N_A_1311_21#_c_372_n N_VGND_c_928_n 0.00435702f $X=7.57 $Y=0.995 $X2=0
+ $Y2=0
cc_377 N_A_1311_21#_c_373_n N_VGND_c_928_n 0.00448878f $X=8.145 $Y=0.995 $X2=0
+ $Y2=0
cc_378 N_A_1311_21#_c_450_p N_VGND_c_928_n 0.0023405f $X=8.31 $Y=0.74 $X2=0
+ $Y2=0
cc_379 N_A_1311_21#_c_404_n N_VGND_c_930_n 0.00298484f $X=8.785 $Y=0.74 $X2=0
+ $Y2=0
cc_380 N_A_1311_21#_c_376_n N_VGND_c_930_n 0.0179308f $X=8.87 $Y=0.42 $X2=0
+ $Y2=0
cc_381 N_A_1311_21#_M1029_d N_VGND_c_931_n 0.00227813f $X=8.735 $Y=0.235 $X2=0
+ $Y2=0
cc_382 N_A_1311_21#_c_370_n N_VGND_c_931_n 0.00466975f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_383 N_A_1311_21#_c_371_n N_VGND_c_931_n 0.00610838f $X=7.1 $Y=0.995 $X2=0
+ $Y2=0
cc_384 N_A_1311_21#_c_372_n N_VGND_c_931_n 0.00627182f $X=7.57 $Y=0.995 $X2=0
+ $Y2=0
cc_385 N_A_1311_21#_c_373_n N_VGND_c_931_n 0.00693478f $X=8.145 $Y=0.995 $X2=0
+ $Y2=0
cc_386 N_A_1311_21#_c_404_n N_VGND_c_931_n 0.00643535f $X=8.785 $Y=0.74 $X2=0
+ $Y2=0
cc_387 N_A_1311_21#_c_450_p N_VGND_c_931_n 0.00393914f $X=8.31 $Y=0.74 $X2=0
+ $Y2=0
cc_388 N_A_1311_21#_c_376_n N_VGND_c_931_n 0.00992122f $X=8.87 $Y=0.42 $X2=0
+ $Y2=0
cc_389 N_Y_c_487_n N_A_117_297#_M1002_s 0.00501331f $X=4.02 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_390 N_Y_c_487_n N_A_117_297#_M1022_s 0.00501331f $X=4.02 $Y=2.34 $X2=0 $Y2=0
cc_391 N_Y_M1015_d N_A_117_297#_c_556_n 0.00510345f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_392 N_Y_M1030_d N_A_117_297#_c_556_n 0.00992815f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_393 N_Y_M1007_d N_A_117_297#_c_556_n 0.00364655f $X=2.935 $Y=1.485 $X2=0
+ $Y2=0
cc_394 N_Y_M1017_d N_A_117_297#_c_556_n 0.00822488f $X=3.875 $Y=1.485 $X2=0
+ $Y2=0
cc_395 N_Y_c_487_n N_A_117_297#_c_556_n 0.0424407f $X=4.02 $Y=2.34 $X2=0 $Y2=0
cc_396 Y N_A_117_297#_c_556_n 0.0121051f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_397 N_Y_c_487_n N_A_493_297#_M1000_s 0.00367601f $X=4.02 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_398 N_Y_c_487_n N_A_493_297#_M1011_s 0.00367601f $X=4.02 $Y=2.34 $X2=0 $Y2=0
cc_399 N_Y_M1007_d N_A_493_297#_c_597_n 0.00351463f $X=2.935 $Y=1.485 $X2=0
+ $Y2=0
cc_400 N_Y_M1017_d N_A_493_297#_c_597_n 0.00529004f $X=3.875 $Y=1.485 $X2=0
+ $Y2=0
cc_401 N_Y_c_487_n N_A_493_297#_c_597_n 0.0929488f $X=4.02 $Y=2.34 $X2=0 $Y2=0
cc_402 N_Y_c_487_n N_VPWR_c_657_n 0.0137365f $X=4.02 $Y=2.34 $X2=0 $Y2=0
cc_403 N_Y_c_487_n N_VPWR_c_661_n 0.17281f $X=4.02 $Y=2.34 $X2=0 $Y2=0
cc_404 N_Y_c_489_n N_VPWR_c_661_n 0.0125737f $X=0.207 $Y=2.255 $X2=0 $Y2=0
cc_405 N_Y_M1002_d N_VPWR_c_656_n 0.00219877f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_406 N_Y_M1015_d N_VPWR_c_656_n 0.00233855f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_407 N_Y_M1030_d N_VPWR_c_656_n 0.00233855f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_408 N_Y_M1007_d N_VPWR_c_656_n 0.00233855f $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_409 N_Y_M1017_d N_VPWR_c_656_n 0.0021994f $X=3.875 $Y=1.485 $X2=0 $Y2=0
cc_410 N_Y_c_487_n N_VPWR_c_656_n 0.133209f $X=4.02 $Y=2.34 $X2=0 $Y2=0
cc_411 N_Y_c_489_n N_VPWR_c_656_n 0.00848224f $X=0.207 $Y=2.255 $X2=0 $Y2=0
cc_412 N_Y_c_484_n N_A_109_47#_M1010_d 0.00422721f $X=4.02 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_413 N_Y_c_484_n N_A_109_47#_M1025_d 0.00520516f $X=4.02 $Y=0.4 $X2=0 $Y2=0
cc_414 N_Y_M1032_s N_A_109_47#_c_775_n 0.00213469f $X=2.005 $Y=0.235 $X2=0 $Y2=0
cc_415 N_Y_c_484_n N_A_109_47#_c_775_n 0.0171891f $X=4.02 $Y=0.4 $X2=0 $Y2=0
cc_416 N_Y_c_484_n N_A_109_47#_c_776_n 0.00224225f $X=4.02 $Y=0.4 $X2=0 $Y2=0
cc_417 N_Y_M1012_s N_A_109_47#_c_788_n 0.00493404f $X=1.015 $Y=0.235 $X2=0 $Y2=0
cc_418 N_Y_c_484_n N_A_109_47#_c_788_n 0.0670205f $X=4.02 $Y=0.4 $X2=0 $Y2=0
cc_419 Y N_A_109_47#_c_788_n 0.0121051f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_420 N_Y_c_484_n N_A_485_47#_M1013_s 0.00410643f $X=4.02 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_421 N_Y_c_484_n N_A_485_47#_M1026_s 0.0051787f $X=4.02 $Y=0.4 $X2=0 $Y2=0
cc_422 N_Y_M1019_d N_A_485_47#_c_867_n 0.00309592f $X=2.895 $Y=0.235 $X2=0 $Y2=0
cc_423 N_Y_M1027_d N_A_485_47#_c_867_n 0.00496297f $X=3.885 $Y=0.235 $X2=0 $Y2=0
cc_424 N_Y_c_484_n N_A_485_47#_c_867_n 0.0870091f $X=4.02 $Y=0.4 $X2=0 $Y2=0
cc_425 N_Y_c_484_n N_VGND_c_918_n 0.012183f $X=4.02 $Y=0.4 $X2=0 $Y2=0
cc_426 N_Y_c_484_n N_VGND_c_924_n 0.157323f $X=4.02 $Y=0.4 $X2=0 $Y2=0
cc_427 N_Y_c_485_n N_VGND_c_924_n 0.0114485f $X=0.207 $Y=0.485 $X2=0 $Y2=0
cc_428 N_Y_M1010_s N_VGND_c_931_n 0.00213654f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_429 N_Y_M1012_s N_VGND_c_931_n 0.00260777f $X=1.015 $Y=0.235 $X2=0 $Y2=0
cc_430 N_Y_M1032_s N_VGND_c_931_n 0.00180037f $X=2.005 $Y=0.235 $X2=0 $Y2=0
cc_431 N_Y_M1019_d N_VGND_c_931_n 0.00213626f $X=2.895 $Y=0.235 $X2=0 $Y2=0
cc_432 N_Y_M1027_d N_VGND_c_931_n 0.00175336f $X=3.885 $Y=0.235 $X2=0 $Y2=0
cc_433 N_Y_c_484_n N_VGND_c_931_n 0.0841512f $X=4.02 $Y=0.4 $X2=0 $Y2=0
cc_434 N_Y_c_485_n N_VGND_c_931_n 0.00840192f $X=0.207 $Y=0.485 $X2=0 $Y2=0
cc_435 N_A_117_297#_c_556_n N_A_493_297#_M1000_s 0.00364655f $X=5.95 $Y=1.66
+ $X2=-0.19 $Y2=1.305
cc_436 N_A_117_297#_c_556_n N_A_493_297#_M1011_s 0.00364655f $X=5.95 $Y=1.66
+ $X2=0 $Y2=0
cc_437 N_A_117_297#_M1005_d N_A_493_297#_c_597_n 0.00478012f $X=4.865 $Y=1.485
+ $X2=0 $Y2=0
cc_438 N_A_117_297#_M1020_d N_A_493_297#_c_597_n 0.00478012f $X=5.805 $Y=1.485
+ $X2=0 $Y2=0
cc_439 N_A_117_297#_c_556_n N_A_493_297#_c_597_n 0.208022f $X=5.95 $Y=1.66 $X2=0
+ $Y2=0
cc_440 N_A_117_297#_c_556_n N_VPWR_M1005_s 0.00537349f $X=5.95 $Y=1.66 $X2=-0.19
+ $Y2=1.305
cc_441 N_A_117_297#_c_556_n N_VPWR_M1009_s 0.00374855f $X=5.95 $Y=1.66 $X2=0
+ $Y2=0
cc_442 N_A_117_297#_M1002_s N_VPWR_c_656_n 0.00235479f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_443 N_A_117_297#_M1022_s N_VPWR_c_656_n 0.00235479f $X=1.525 $Y=1.485 $X2=0
+ $Y2=0
cc_444 N_A_117_297#_M1005_d N_VPWR_c_656_n 0.00338665f $X=4.865 $Y=1.485 $X2=0
+ $Y2=0
cc_445 N_A_117_297#_M1020_d N_VPWR_c_656_n 0.00338665f $X=5.805 $Y=1.485 $X2=0
+ $Y2=0
cc_446 N_A_117_297#_c_556_n N_A_109_47#_c_776_n 0.00623829f $X=5.95 $Y=1.66
+ $X2=0 $Y2=0
cc_447 N_A_117_297#_c_556_n N_A_109_47#_c_778_n 0.00686595f $X=5.95 $Y=1.66
+ $X2=0 $Y2=0
cc_448 N_A_493_297#_c_597_n N_VPWR_M1005_s 0.00508531f $X=6.805 $Y=2 $X2=-0.19
+ $Y2=1.305
cc_449 N_A_493_297#_c_597_n N_VPWR_M1009_s 0.00351043f $X=6.805 $Y=2 $X2=0 $Y2=0
cc_450 N_A_493_297#_c_597_n N_VPWR_M1031_s 0.00446737f $X=6.805 $Y=2 $X2=0 $Y2=0
cc_451 N_A_493_297#_c_611_n N_VPWR_M1014_d 0.00404868f $X=7.745 $Y=2 $X2=0 $Y2=0
cc_452 N_A_493_297#_c_597_n N_VPWR_c_657_n 0.0206557f $X=6.805 $Y=2 $X2=0 $Y2=0
cc_453 N_A_493_297#_c_597_n N_VPWR_c_658_n 0.00860446f $X=6.805 $Y=2 $X2=0 $Y2=0
cc_454 N_A_493_297#_c_597_n N_VPWR_c_659_n 0.00861424f $X=6.805 $Y=2 $X2=0 $Y2=0
cc_455 N_A_493_297#_c_597_n N_VPWR_c_661_n 0.00346265f $X=6.805 $Y=2 $X2=0 $Y2=0
cc_456 N_A_493_297#_c_637_p N_VPWR_c_663_n 0.0156776f $X=6.89 $Y=2.3 $X2=0 $Y2=0
cc_457 N_A_493_297#_c_611_n N_VPWR_c_663_n 0.0196308f $X=7.745 $Y=2 $X2=0 $Y2=0
cc_458 N_A_493_297#_c_618_n N_VPWR_c_663_n 0.0128538f $X=7.83 $Y=2.3 $X2=0 $Y2=0
cc_459 N_A_493_297#_c_597_n N_VPWR_c_664_n 0.00319869f $X=6.805 $Y=2 $X2=0 $Y2=0
cc_460 N_A_493_297#_c_637_p N_VPWR_c_664_n 0.011801f $X=6.89 $Y=2.3 $X2=0 $Y2=0
cc_461 N_A_493_297#_c_611_n N_VPWR_c_664_n 0.00238051f $X=7.745 $Y=2 $X2=0 $Y2=0
cc_462 N_A_493_297#_c_611_n N_VPWR_c_665_n 0.00319869f $X=7.745 $Y=2 $X2=0 $Y2=0
cc_463 N_A_493_297#_c_618_n N_VPWR_c_665_n 0.011801f $X=7.83 $Y=2.3 $X2=0 $Y2=0
cc_464 N_A_493_297#_M1000_s N_VPWR_c_656_n 0.00235479f $X=2.465 $Y=1.485 $X2=0
+ $Y2=0
cc_465 N_A_493_297#_M1011_s N_VPWR_c_656_n 0.00235479f $X=3.405 $Y=1.485 $X2=0
+ $Y2=0
cc_466 N_A_493_297#_M1003_s N_VPWR_c_656_n 0.00272704f $X=6.745 $Y=1.485 $X2=0
+ $Y2=0
cc_467 N_A_493_297#_M1018_s N_VPWR_c_656_n 0.00699652f $X=7.685 $Y=1.485 $X2=0
+ $Y2=0
cc_468 N_A_493_297#_c_597_n N_VPWR_c_656_n 0.0479794f $X=6.805 $Y=2 $X2=0 $Y2=0
cc_469 N_A_493_297#_c_637_p N_VPWR_c_656_n 0.00646745f $X=6.89 $Y=2.3 $X2=0
+ $Y2=0
cc_470 N_A_493_297#_c_611_n N_VPWR_c_656_n 0.0114411f $X=7.745 $Y=2 $X2=0 $Y2=0
cc_471 N_A_493_297#_c_618_n N_VPWR_c_656_n 0.00646745f $X=7.83 $Y=2.3 $X2=0
+ $Y2=0
cc_472 N_A_493_297#_c_597_n N_VPWR_c_669_n 0.0196308f $X=6.805 $Y=2 $X2=0 $Y2=0
cc_473 N_A_493_297#_c_597_n N_VPWR_c_670_n 0.0196307f $X=6.805 $Y=2 $X2=0 $Y2=0
cc_474 N_A_493_297#_c_637_p N_VPWR_c_670_n 0.0128538f $X=6.89 $Y=2.3 $X2=0 $Y2=0
cc_475 N_A_109_47#_c_775_n N_A_485_47#_M1016_s 0.0014194f $X=6.69 $Y=0.85 $X2=0
+ $Y2=0
cc_476 N_A_109_47#_c_775_n N_A_485_47#_c_867_n 0.0739797f $X=6.69 $Y=0.85 $X2=0
+ $Y2=0
cc_477 N_A_109_47#_c_776_n N_A_485_47#_c_867_n 9.22088e-19 $X=1.91 $Y=0.85 $X2=0
+ $Y2=0
cc_478 N_A_109_47#_c_778_n N_A_485_47#_c_867_n 0.00244004f $X=1.67 $Y=0.74 $X2=0
+ $Y2=0
cc_479 N_A_109_47#_c_775_n N_A_485_47#_c_879_n 0.031146f $X=6.69 $Y=0.85 $X2=0
+ $Y2=0
cc_480 N_A_109_47#_c_775_n N_A_485_47#_c_885_n 0.00672766f $X=6.69 $Y=0.85 $X2=0
+ $Y2=0
cc_481 N_A_109_47#_c_775_n N_VGND_M1024_d 0.0019359f $X=6.69 $Y=0.85 $X2=0 $Y2=0
cc_482 N_A_109_47#_c_773_n N_VGND_M1004_d 0.00224377f $X=7.745 $Y=0.81 $X2=0
+ $Y2=0
cc_483 N_A_109_47#_c_775_n N_VGND_c_918_n 0.00135173f $X=6.69 $Y=0.85 $X2=0
+ $Y2=0
cc_484 N_A_109_47#_c_811_n N_VGND_c_921_n 0.0205277f $X=6.89 $Y=0.42 $X2=0 $Y2=0
cc_485 N_A_109_47#_c_775_n N_VGND_c_921_n 0.00688907f $X=6.69 $Y=0.85 $X2=0
+ $Y2=0
cc_486 N_A_109_47#_c_773_n N_VGND_c_922_n 0.0150984f $X=7.745 $Y=0.81 $X2=0
+ $Y2=0
cc_487 N_A_109_47#_c_774_n N_VGND_c_922_n 0.0020224f $X=7.83 $Y=0.675 $X2=0
+ $Y2=0
cc_488 N_A_109_47#_c_811_n N_VGND_c_926_n 0.0116287f $X=6.89 $Y=0.42 $X2=0 $Y2=0
cc_489 N_A_109_47#_c_779_n N_VGND_c_926_n 0.00313081f $X=7.1 $Y=0.825 $X2=0
+ $Y2=0
cc_490 N_A_109_47#_c_773_n N_VGND_c_928_n 0.00314682f $X=7.745 $Y=0.81 $X2=0
+ $Y2=0
cc_491 N_A_109_47#_c_774_n N_VGND_c_928_n 0.00420686f $X=7.83 $Y=0.675 $X2=0
+ $Y2=0
cc_492 N_A_109_47#_M1010_d N_VGND_c_931_n 0.00262417f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_493 N_A_109_47#_M1025_d N_VGND_c_931_n 0.00263016f $X=1.485 $Y=0.235 $X2=0
+ $Y2=0
cc_494 N_A_109_47#_M1001_s N_VGND_c_931_n 0.00284605f $X=6.705 $Y=0.235 $X2=0
+ $Y2=0
cc_495 N_A_109_47#_M1021_s N_VGND_c_931_n 0.00963868f $X=7.645 $Y=0.235 $X2=0
+ $Y2=0
cc_496 N_A_109_47#_c_811_n N_VGND_c_931_n 0.00295874f $X=6.89 $Y=0.42 $X2=0
+ $Y2=0
cc_497 N_A_109_47#_c_773_n N_VGND_c_931_n 0.00689674f $X=7.745 $Y=0.81 $X2=0
+ $Y2=0
cc_498 N_A_109_47#_c_774_n N_VGND_c_931_n 0.00540999f $X=7.83 $Y=0.675 $X2=0
+ $Y2=0
cc_499 N_A_109_47#_c_775_n N_VGND_c_931_n 0.217422f $X=6.69 $Y=0.85 $X2=0 $Y2=0
cc_500 N_A_109_47#_c_776_n N_VGND_c_931_n 0.0146935f $X=1.91 $Y=0.85 $X2=0 $Y2=0
cc_501 N_A_109_47#_c_777_n N_VGND_c_931_n 0.0176392f $X=6.885 $Y=0.85 $X2=0
+ $Y2=0
cc_502 N_A_109_47#_c_779_n N_VGND_c_931_n 0.00565548f $X=7.1 $Y=0.825 $X2=0
+ $Y2=0
cc_503 N_A_109_47#_c_775_n N_VGND_c_932_n 0.00151302f $X=6.69 $Y=0.85 $X2=0
+ $Y2=0
cc_504 N_A_485_47#_c_867_n N_VGND_M1006_d 0.00564723f $X=4.925 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_505 N_A_485_47#_c_879_n N_VGND_M1008_d 0.00361385f $X=5.865 $Y=0.74 $X2=0
+ $Y2=0
cc_506 N_A_485_47#_c_867_n N_VGND_c_918_n 0.0185297f $X=4.925 $Y=0.74 $X2=0
+ $Y2=0
cc_507 N_A_485_47#_c_867_n N_VGND_c_919_n 0.00298484f $X=4.925 $Y=0.74 $X2=0
+ $Y2=0
cc_508 N_A_485_47#_c_878_n N_VGND_c_919_n 0.011459f $X=5.01 $Y=0.42 $X2=0 $Y2=0
cc_509 N_A_485_47#_c_879_n N_VGND_c_919_n 0.00233622f $X=5.865 $Y=0.74 $X2=0
+ $Y2=0
cc_510 N_A_485_47#_c_879_n N_VGND_c_920_n 0.00299413f $X=5.865 $Y=0.74 $X2=0
+ $Y2=0
cc_511 N_A_485_47#_c_884_n N_VGND_c_920_n 0.011459f $X=5.95 $Y=0.42 $X2=0 $Y2=0
cc_512 N_A_485_47#_c_884_n N_VGND_c_921_n 0.0249836f $X=5.95 $Y=0.42 $X2=0 $Y2=0
cc_513 N_A_485_47#_c_867_n N_VGND_c_924_n 0.00332039f $X=4.925 $Y=0.74 $X2=0
+ $Y2=0
cc_514 N_A_485_47#_M1013_s N_VGND_c_931_n 0.0021497f $X=2.425 $Y=0.235 $X2=0
+ $Y2=0
cc_515 N_A_485_47#_M1026_s N_VGND_c_931_n 0.00248559f $X=3.365 $Y=0.235 $X2=0
+ $Y2=0
cc_516 N_A_485_47#_M1006_s N_VGND_c_931_n 0.00245057f $X=4.875 $Y=0.235 $X2=0
+ $Y2=0
cc_517 N_A_485_47#_M1016_s N_VGND_c_931_n 0.00300458f $X=5.815 $Y=0.235 $X2=0
+ $Y2=0
cc_518 N_A_485_47#_c_867_n N_VGND_c_931_n 0.0087015f $X=4.925 $Y=0.74 $X2=0
+ $Y2=0
cc_519 N_A_485_47#_c_878_n N_VGND_c_931_n 0.00305234f $X=5.01 $Y=0.42 $X2=0
+ $Y2=0
cc_520 N_A_485_47#_c_879_n N_VGND_c_931_n 0.00520815f $X=5.865 $Y=0.74 $X2=0
+ $Y2=0
cc_521 N_A_485_47#_c_884_n N_VGND_c_931_n 0.00305234f $X=5.95 $Y=0.42 $X2=0
+ $Y2=0
cc_522 N_A_485_47#_c_878_n N_VGND_c_932_n 0.0156777f $X=5.01 $Y=0.42 $X2=0 $Y2=0
cc_523 N_A_485_47#_c_879_n N_VGND_c_932_n 0.0176018f $X=5.865 $Y=0.74 $X2=0
+ $Y2=0
