* File: sky130_fd_sc_hdll__nor4bb_2.pex.spice
* Created: Thu Aug 27 19:17:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_2%D_N 3 5 6 8 9 10 14 15 16
c33 15 0 3.26347e-20 $X=0.53 $Y=1.16
c34 14 0 7.12326e-20 $X=0.53 $Y=1.16
r35 14 17 39.6736 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.16
+ $X2=0.545 $Y2=1.325
r36 14 16 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.16
+ $X2=0.545 $Y2=0.995
r37 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.16 $X2=0.53 $Y2=1.16
r38 9 10 9.67483 $w=4.03e-07 $l=3.4e-07 $layer=LI1_cond $X=0.627 $Y=1.19
+ $X2=0.627 $Y2=1.53
r39 9 15 0.853661 $w=4.03e-07 $l=3e-08 $layer=LI1_cond $X=0.627 $Y=1.19
+ $X2=0.627 $Y2=1.16
r40 6 8 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.975
+ $X2=0.495 $Y2=2.26
r41 5 6 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.875 $X2=0.495
+ $Y2=1.975
r42 5 17 182.367 $w=2e-07 $l=5.5e-07 $layer=POLY_cond $X=0.495 $Y=1.875
+ $X2=0.495 $Y2=1.325
r43 3 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.47 $Y=0.675
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_2%C_N 1 3 4 6 7 15
c31 15 0 1.69374e-19 $X=1.155 $Y=1.19
r32 7 15 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=1.085 $Y=1.16 $X2=1.155
+ $Y2=1.16
r33 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.085
+ $Y=1.16 $X2=1.085 $Y2=1.16
r34 4 10 46.2237 $w=3.35e-07 $l=2.89396e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.115 $Y2=1.16
r35 4 6 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.03 $Y=1.41 $X2=1.03
+ $Y2=1.695
r36 1 10 38.6365 $w=3.35e-07 $l=2.13014e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.115 $Y2=1.16
r37 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_2%A_216_93# 1 2 7 9 10 12 13 15 16 18 19 24
+ 26 29 33 35 39
c77 39 0 1.69374e-19 $X=2.545 $Y=1.202
c78 29 0 1.18672e-19 $X=2.31 $Y=1.16
c79 24 0 3.26347e-20 $X=1.525 $Y=1.075
c80 13 0 9.6109e-20 $X=2.545 $Y=1.41
r81 39 40 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=2.545 $Y=1.202
+ $X2=2.57 $Y2=1.202
r82 36 37 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=2.075 $Y=1.202
+ $X2=2.1 $Y2=1.202
r83 33 34 13.5292 $w=2.57e-07 $l=2.85e-07 $layer=LI1_cond $X=1.24 $Y=0.655
+ $X2=1.525 $Y2=0.655
r84 30 39 30.6965 $w=3.69e-07 $l=2.35e-07 $layer=POLY_cond $X=2.31 $Y=1.202
+ $X2=2.545 $Y2=1.202
r85 30 37 27.4309 $w=3.69e-07 $l=2.1e-07 $layer=POLY_cond $X=2.31 $Y=1.202
+ $X2=2.1 $Y2=1.202
r86 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.31
+ $Y=1.16 $X2=2.31 $Y2=1.16
r87 27 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=1.16
+ $X2=1.525 $Y2=1.16
r88 27 29 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.61 $Y=1.16 $X2=2.31
+ $Y2=1.16
r89 25 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=1.245
+ $X2=1.525 $Y2=1.16
r90 25 26 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.525 $Y=1.245
+ $X2=1.525 $Y2=1.525
r91 24 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=1.075
+ $X2=1.525 $Y2=1.16
r92 23 34 3.1561 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.525 $Y=0.825
+ $X2=1.525 $Y2=0.655
r93 23 24 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.525 $Y=0.825
+ $X2=1.525 $Y2=1.075
r94 19 26 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.44 $Y=1.62
+ $X2=1.525 $Y2=1.525
r95 19 21 10.2153 $w=1.88e-07 $l=1.75e-07 $layer=LI1_cond $X=1.44 $Y=1.62
+ $X2=1.265 $Y2=1.62
r96 16 40 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=1.202
r97 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=0.56
r98 13 39 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.545 $Y=1.41
+ $X2=2.545 $Y2=1.202
r99 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.545 $Y=1.41
+ $X2=2.545 $Y2=1.985
r100 10 37 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.1 $Y=0.995
+ $X2=2.1 $Y2=1.202
r101 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.1 $Y=0.995
+ $X2=2.1 $Y2=0.56
r102 7 36 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.075 $Y=1.41
+ $X2=2.075 $Y2=1.202
r103 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.075 $Y=1.41
+ $X2=2.075 $Y2=1.985
r104 2 21 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.485 $X2=1.265 $Y2=1.63
r105 1 33 182 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.465 $X2=1.24 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_2%A_27_93# 1 2 7 9 10 12 13 15 16 18 20 23
+ 25 28 29 30 32 33 35 41 43 47
c100 47 0 1.18672e-19 $X=3.485 $Y=1.202
c101 32 0 9.6109e-20 $X=2.78 $Y=1.415
r102 47 48 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.485 $Y=1.202
+ $X2=3.51 $Y2=1.202
r103 44 45 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=2.99 $Y=1.202
+ $X2=3.015 $Y2=1.202
r104 38 41 2.76586 $w=3.73e-07 $l=9e-08 $layer=LI1_cond $X=0.17 $Y=0.637
+ $X2=0.26 $Y2=0.637
r105 36 47 5.70789 $w=3.8e-07 $l=4.5e-08 $layer=POLY_cond $X=3.44 $Y=1.202
+ $X2=3.485 $Y2=1.202
r106 36 45 53.9079 $w=3.8e-07 $l=4.25e-07 $layer=POLY_cond $X=3.44 $Y=1.202
+ $X2=3.015 $Y2=1.202
r107 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.44
+ $Y=1.16 $X2=3.44 $Y2=1.16
r108 33 35 31.8864 $w=1.98e-07 $l=5.75e-07 $layer=LI1_cond $X=2.865 $Y=1.175
+ $X2=3.44 $Y2=1.175
r109 31 33 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.78 $Y=1.275
+ $X2=2.865 $Y2=1.175
r110 31 32 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.78 $Y=1.275
+ $X2=2.78 $Y2=1.415
r111 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.695 $Y=1.5
+ $X2=2.78 $Y2=1.415
r112 29 30 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.695 $Y=1.5
+ $X2=1.95 $Y2=1.5
r113 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.865 $Y=1.585
+ $X2=1.95 $Y2=1.5
r114 27 28 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.865 $Y=1.585
+ $X2=1.865 $Y2=1.885
r115 26 43 2.20034 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.97
+ $X2=0.215 $Y2=1.97
r116 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.78 $Y=1.97
+ $X2=1.865 $Y2=1.885
r117 25 26 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=1.78 $Y=1.97
+ $X2=0.345 $Y2=1.97
r118 21 43 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.215 $Y=2.055
+ $X2=0.215 $Y2=1.97
r119 21 23 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=0.215 $Y=2.055
+ $X2=0.215 $Y2=2.29
r120 20 43 4.23118 $w=2.15e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.17 $Y=1.885
+ $X2=0.215 $Y2=1.97
r121 19 38 5.38787 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=0.637
r122 19 20 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=1.885
r123 16 48 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=1.202
r124 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=0.56
r125 13 47 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.485 $Y=1.41
+ $X2=3.485 $Y2=1.202
r126 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.485 $Y=1.41
+ $X2=3.485 $Y2=1.985
r127 10 45 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.015 $Y=1.41
+ $X2=3.015 $Y2=1.202
r128 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.015 $Y=1.41
+ $X2=3.015 $Y2=1.985
r129 7 44 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=1.202
r130 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=0.56
r131 2 23 600 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.05 $X2=0.26 $Y2=2.29
r132 1 41 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_2%B 1 3 4 6 7 9 10 12 13 19 20 23
c45 20 0 1.40272e-19 $X=4.965 $Y=1.202
r46 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.965 $Y=1.202
+ $X2=4.99 $Y2=1.202
r47 18 20 27.9053 $w=3.8e-07 $l=2.2e-07 $layer=POLY_cond $X=4.745 $Y=1.202
+ $X2=4.965 $Y2=1.202
r48 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.745
+ $Y=1.16 $X2=4.745 $Y2=1.16
r49 16 18 31.7105 $w=3.8e-07 $l=2.5e-07 $layer=POLY_cond $X=4.495 $Y=1.202
+ $X2=4.745 $Y2=1.202
r50 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.47 $Y=1.202
+ $X2=4.495 $Y2=1.202
r51 13 19 4.99091 $w=1.98e-07 $l=9e-08 $layer=LI1_cond $X=4.655 $Y=1.175
+ $X2=4.745 $Y2=1.175
r52 13 23 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=4.655 $Y=1.175
+ $X2=4.645 $Y2=1.175
r53 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.99 $Y=0.995
+ $X2=4.99 $Y2=1.202
r54 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.99 $Y=0.995
+ $X2=4.99 $Y2=0.56
r55 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.965 $Y=1.41
+ $X2=4.965 $Y2=1.202
r56 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.965 $Y=1.41
+ $X2=4.965 $Y2=1.985
r57 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.495 $Y=1.41
+ $X2=4.495 $Y2=1.202
r58 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.495 $Y=1.41
+ $X2=4.495 $Y2=1.985
r59 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.47 $Y=0.995
+ $X2=4.47 $Y2=1.202
r60 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.47 $Y=0.995 $X2=4.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_2%A 1 3 4 6 7 9 10 12 13 20
c36 13 0 1.40272e-19 $X=5.67 $Y=1.19
c37 4 0 6.56464e-20 $X=5.435 $Y=1.41
r38 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=5.905 $Y=1.202
+ $X2=5.93 $Y2=1.202
r39 18 20 28.5395 $w=3.8e-07 $l=2.25e-07 $layer=POLY_cond $X=5.68 $Y=1.202
+ $X2=5.905 $Y2=1.202
r40 16 18 31.0763 $w=3.8e-07 $l=2.45e-07 $layer=POLY_cond $X=5.435 $Y=1.202
+ $X2=5.68 $Y2=1.202
r41 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=5.41 $Y=1.202
+ $X2=5.435 $Y2=1.202
r42 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.68
+ $Y=1.16 $X2=5.68 $Y2=1.16
r43 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.93 $Y=0.995
+ $X2=5.93 $Y2=1.202
r44 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.93 $Y=0.995
+ $X2=5.93 $Y2=0.56
r45 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.905 $Y=1.41
+ $X2=5.905 $Y2=1.202
r46 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.905 $Y=1.41
+ $X2=5.905 $Y2=1.985
r47 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.435 $Y=1.41
+ $X2=5.435 $Y2=1.202
r48 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.435 $Y=1.41
+ $X2=5.435 $Y2=1.985
r49 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.41 $Y=0.995
+ $X2=5.41 $Y2=1.202
r50 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.41 $Y=0.995 $X2=5.41
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_2%VPWR 1 2 9 13 16 17 18 20 33 34 37
r62 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r63 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r64 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r65 30 31 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r66 28 31 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=1.15 $Y=2.72 $X2=5.29
+ $Y2=2.72
r67 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r68 27 30 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=5.29 $Y2=2.72
r69 27 28 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r70 25 37 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r71 25 27 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r72 20 37 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r73 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r74 18 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r75 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r76 16 30 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.545 $Y=2.72
+ $X2=5.29 $Y2=2.72
r77 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.545 $Y=2.72
+ $X2=5.65 $Y2=2.72
r78 15 33 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=5.755 $Y=2.72
+ $X2=6.21 $Y2=2.72
r79 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.755 $Y=2.72
+ $X2=5.65 $Y2=2.72
r80 11 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.65 $Y=2.635
+ $X2=5.65 $Y2=2.72
r81 11 13 35.6493 $w=2.08e-07 $l=6.75e-07 $layer=LI1_cond $X=5.65 $Y=2.635
+ $X2=5.65 $Y2=1.96
r82 7 37 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r83 7 9 9.40151 $w=3.78e-07 $l=3.1e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.325
r84 2 13 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.525
+ $Y=1.485 $X2=5.67 $Y2=1.96
r85 1 9 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.05 $X2=0.73 $Y2=2.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_2%A_343_297# 1 2 3 16
r24 14 16 45.1374 $w=2.38e-07 $l=9.4e-07 $layer=LI1_cond $X=2.78 $Y=2.345
+ $X2=3.72 $Y2=2.345
r25 11 14 45.1374 $w=2.38e-07 $l=9.4e-07 $layer=LI1_cond $X=1.84 $Y=2.345
+ $X2=2.78 $Y2=2.345
r26 3 16 600 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=3.575
+ $Y=1.485 $X2=3.72 $Y2=2.31
r27 2 14 600 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=1.485 $X2=2.78 $Y2=2.31
r28 1 11 600 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=1.715
+ $Y=1.485 $X2=1.84 $Y2=2.31
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_2%A_433_297# 1 2 7 11 13
c35 13 0 6.56464e-20 $X=4.73 $Y=1.62
r36 11 16 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=1.875
+ $X2=4.75 $Y2=1.96
r37 11 13 10.1336 $w=2.88e-07 $l=2.55e-07 $layer=LI1_cond $X=4.75 $Y=1.875
+ $X2=4.75 $Y2=1.62
r38 7 16 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.605 $Y=1.96
+ $X2=4.75 $Y2=1.96
r39 7 9 149.727 $w=1.68e-07 $l=2.295e-06 $layer=LI1_cond $X=4.605 $Y=1.96
+ $X2=2.31 $Y2=1.96
r40 2 16 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=4.585
+ $Y=1.485 $X2=4.73 $Y2=1.96
r41 2 13 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.585
+ $Y=1.485 $X2=4.73 $Y2=1.62
r42 1 9 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=2.165
+ $Y=1.485 $X2=2.31 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_2%Y 1 2 3 4 5 18 20 21 24 26 28 32 34 38 40
+ 42 43 44 45 49 55
r104 49 55 4.87572 $w=2.58e-07 $l=1.1e-07 $layer=LI1_cond $X=3.81 $Y=1.575
+ $X2=3.7 $Y2=1.575
r105 45 49 4.52065 $w=2.6e-07 $l=2.1e-07 $layer=LI1_cond $X=4.02 $Y=1.575
+ $X2=3.81 $Y2=1.575
r106 44 55 0.664871 $w=2.58e-07 $l=1.5e-08 $layer=LI1_cond $X=3.685 $Y=1.575
+ $X2=3.7 $Y2=1.575
r107 44 51 19.2813 $w=2.58e-07 $l=4.35e-07 $layer=LI1_cond $X=3.685 $Y=1.575
+ $X2=3.25 $Y2=1.575
r108 41 45 11.9572 $w=5.88e-07 $l=5.4e-07 $layer=LI1_cond $X=4.02 $Y=0.905
+ $X2=4.02 $Y2=1.445
r109 41 42 1.44414 $w=4.2e-07 $l=9e-08 $layer=LI1_cond $X=4.02 $Y=0.905 $X2=4.02
+ $Y2=0.815
r110 36 38 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.645 $Y=0.725
+ $X2=5.645 $Y2=0.39
r111 35 43 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.895 $Y=0.815
+ $X2=4.705 $Y2=0.815
r112 34 36 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=5.455 $Y=0.815
+ $X2=5.645 $Y2=0.725
r113 34 35 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=5.455 $Y=0.815
+ $X2=4.895 $Y2=0.815
r114 30 43 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=4.705 $Y=0.725
+ $X2=4.705 $Y2=0.815
r115 30 32 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.705 $Y=0.725
+ $X2=4.705 $Y2=0.39
r116 29 42 9.75736 $w=1.8e-07 $l=2.1e-07 $layer=LI1_cond $X=4.23 $Y=0.815
+ $X2=4.02 $Y2=0.815
r117 28 43 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.515 $Y=0.815
+ $X2=4.705 $Y2=0.815
r118 28 29 17.5606 $w=1.78e-07 $l=2.85e-07 $layer=LI1_cond $X=4.515 $Y=0.815
+ $X2=4.23 $Y2=0.815
r119 27 40 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.415 $Y=0.815
+ $X2=3.225 $Y2=0.815
r120 26 42 9.75736 $w=1.8e-07 $l=2.1e-07 $layer=LI1_cond $X=3.81 $Y=0.815
+ $X2=4.02 $Y2=0.815
r121 26 27 24.3384 $w=1.78e-07 $l=3.95e-07 $layer=LI1_cond $X=3.81 $Y=0.815
+ $X2=3.415 $Y2=0.815
r122 22 40 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=3.225 $Y=0.725
+ $X2=3.225 $Y2=0.815
r123 22 24 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.225 $Y=0.725
+ $X2=3.225 $Y2=0.39
r124 20 40 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.035 $Y=0.815
+ $X2=3.225 $Y2=0.815
r125 20 21 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.035 $Y=0.815
+ $X2=2.475 $Y2=0.815
r126 16 21 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=2.285 $Y=0.725
+ $X2=2.475 $Y2=0.815
r127 16 18 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.285 $Y=0.725
+ $X2=2.285 $Y2=0.39
r128 5 51 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.105
+ $Y=1.485 $X2=3.25 $Y2=1.62
r129 4 38 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=5.485
+ $Y=0.235 $X2=5.67 $Y2=0.39
r130 3 32 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.545
+ $Y=0.235 $X2=4.73 $Y2=0.39
r131 2 24 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.065
+ $Y=0.235 $X2=3.25 $Y2=0.39
r132 1 18 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.175
+ $Y=0.235 $X2=2.31 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_2%A_823_297# 1 2 3 10 14 15 16 20
r37 20 22 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=6.115 $Y=1.63
+ $X2=6.115 $Y2=2.31
r38 18 20 0.151637 $w=3.78e-07 $l=5e-09 $layer=LI1_cond $X=6.115 $Y=1.625
+ $X2=6.115 $Y2=1.63
r39 17 25 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.325 $Y=1.54
+ $X2=5.22 $Y2=1.54
r40 16 18 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=5.925 $Y=1.54
+ $X2=6.115 $Y2=1.625
r41 16 17 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.925 $Y=1.54
+ $X2=5.325 $Y2=1.54
r42 15 27 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=5.22 $Y=2.215
+ $X2=5.22 $Y2=2.34
r43 14 25 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.22 $Y=1.625
+ $X2=5.22 $Y2=1.54
r44 14 15 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=5.22 $Y=1.625
+ $X2=5.22 $Y2=2.215
r45 10 27 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=5.115 $Y=2.34
+ $X2=5.22 $Y2=2.34
r46 10 12 39.4136 $w=2.48e-07 $l=8.55e-07 $layer=LI1_cond $X=5.115 $Y=2.34
+ $X2=4.26 $Y2=2.34
r47 3 22 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=5.995
+ $Y=1.485 $X2=6.14 $Y2=2.31
r48 3 20 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.995
+ $Y=1.485 $X2=6.14 $Y2=1.63
r49 2 27 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.055
+ $Y=1.485 $X2=5.2 $Y2=2.3
r50 2 25 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=5.055
+ $Y=1.485 $X2=5.2 $Y2=1.62
r51 1 12 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.115
+ $Y=1.485 $X2=4.26 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4BB_2%VGND 1 2 3 4 5 6 7 26 28 32 36 40 42 44
+ 47 48 50 51 52 66 71 74 78 84 87
c95 26 0 7.12326e-20 $X=0.77 $Y=0.66
r96 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r97 83 84 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=4.26 $Y=0.235
+ $X2=4.345 $Y2=0.235
r98 80 83 6.54105 $w=6.38e-07 $l=3.5e-07 $layer=LI1_cond $X=3.91 $Y=0.235
+ $X2=4.26 $Y2=0.235
r99 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r100 77 80 3.55086 $w=6.38e-07 $l=1.9e-07 $layer=LI1_cond $X=3.72 $Y=0.235
+ $X2=3.91 $Y2=0.235
r101 77 78 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=0.235
+ $X2=3.635 $Y2=0.235
r102 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r103 72 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r104 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r105 69 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r106 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r107 66 86 4.23443 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=6.055 $Y=0
+ $X2=6.247 $Y2=0
r108 66 68 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.055 $Y=0
+ $X2=5.75 $Y2=0
r109 65 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r110 65 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=3.91
+ $Y2=0
r111 64 84 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.83 $Y=0
+ $X2=4.345 $Y2=0
r112 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r113 61 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r114 60 78 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.45 $Y=0
+ $X2=3.635 $Y2=0
r115 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r116 57 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r117 57 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r118 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r119 54 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.925 $Y=0 $X2=1.76
+ $Y2=0
r120 54 56 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.925 $Y=0
+ $X2=2.53 $Y2=0
r121 52 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r122 50 64 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.115 $Y=0
+ $X2=4.83 $Y2=0
r123 50 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.115 $Y=0 $X2=5.2
+ $Y2=0
r124 49 68 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=5.285 $Y=0
+ $X2=5.75 $Y2=0
r125 49 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.285 $Y=0 $X2=5.2
+ $Y2=0
r126 47 56 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=0
+ $X2=2.53 $Y2=0
r127 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.78
+ $Y2=0
r128 46 60 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.865 $Y=0
+ $X2=3.45 $Y2=0
r129 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.78
+ $Y2=0
r130 42 86 3.08761 $w=2.75e-07 $l=1.09087e-07 $layer=LI1_cond $X=6.192 $Y=0.085
+ $X2=6.247 $Y2=0
r131 42 44 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=6.192 $Y=0.085
+ $X2=6.192 $Y2=0.39
r132 38 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.2 $Y=0.085 $X2=5.2
+ $Y2=0
r133 38 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.2 $Y=0.085
+ $X2=5.2 $Y2=0.39
r134 34 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0
r135 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0.39
r136 30 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.76 $Y=0.085
+ $X2=1.76 $Y2=0
r137 30 32 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.76 $Y=0.085
+ $X2=1.76 $Y2=0.39
r138 29 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.77
+ $Y2=0
r139 28 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.595 $Y=0 $X2=1.76
+ $Y2=0
r140 28 29 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.595 $Y=0
+ $X2=0.855 $Y2=0
r141 24 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=0.085
+ $X2=0.77 $Y2=0
r142 24 26 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.77 $Y=0.085
+ $X2=0.77 $Y2=0.66
r143 7 44 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.005
+ $Y=0.235 $X2=6.14 $Y2=0.39
r144 6 40 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.065
+ $Y=0.235 $X2=5.2 $Y2=0.39
r145 5 83 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=4.115
+ $Y=0.235 $X2=4.26 $Y2=0.39
r146 4 77 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.39
r147 3 36 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.39
r148 2 32 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.635
+ $Y=0.235 $X2=1.76 $Y2=0.39
r149 1 26 182 $w=1.7e-07 $l=3.07409e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.465 $X2=0.77 $Y2=0.66
.ends

