* File: sky130_fd_sc_hdll__a2bb2o_2.pex.spice
* Created: Thu Aug 27 18:54:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_2%A_82_21# 1 2 7 9 10 12 13 15 16 18 20 21
+ 22 24 25 26 28 31 34 39 43 48
c115 39 0 1.72109e-19 $X=2.785 $Y=2.275
c116 34 0 1.32963e-19 $X=1 $Y=1.16
r117 47 48 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=0.955 $Y=1.202
+ $X2=0.98 $Y2=1.202
r118 46 47 57.504 $w=3.73e-07 $l=4.45e-07 $layer=POLY_cond $X=0.51 $Y=1.202
+ $X2=0.955 $Y2=1.202
r119 45 46 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=0.485 $Y=1.202
+ $X2=0.51 $Y2=1.202
r120 39 40 0.423611 $w=2.88e-07 $l=1e-08 $layer=LI1_cond $X=2.87 $Y=2.275
+ $X2=2.87 $Y2=2.285
r121 35 48 2.58445 $w=3.73e-07 $l=2e-08 $layer=POLY_cond $X=1 $Y=1.202 $X2=0.98
+ $Y2=1.202
r122 34 37 7.14859 $w=3.03e-07 $l=1.65e-07 $layer=LI1_cond $X=1.067 $Y=1.16
+ $X2=1.067 $Y2=1.325
r123 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.16
+ $X2=1 $Y2=1.16
r124 29 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.195 $Y=0.7
+ $X2=3.195 $Y2=0.785
r125 29 31 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.195 $Y=0.7
+ $X2=3.195 $Y2=0.445
r126 28 39 16.8076 $w=2.88e-07 $l=4.3589e-07 $layer=LI1_cond $X=2.99 $Y=1.895
+ $X2=2.87 $Y2=2.275
r127 27 43 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.99 $Y=0.785
+ $X2=3.195 $Y2=0.785
r128 27 28 53.6934 $w=2.18e-07 $l=1.025e-06 $layer=LI1_cond $X=2.99 $Y=0.87
+ $X2=2.99 $Y2=1.895
r129 25 40 3.82142 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.64 $Y=2.285
+ $X2=2.87 $Y2=2.285
r130 25 26 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=2.64 $Y=2.285
+ $X2=1.86 $Y2=2.285
r131 24 26 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.75 $Y=2.2
+ $X2=1.86 $Y2=2.285
r132 23 24 11.7863 $w=2.18e-07 $l=2.25e-07 $layer=LI1_cond $X=1.75 $Y=1.975
+ $X2=1.75 $Y2=2.2
r133 21 23 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.64 $Y=1.89
+ $X2=1.75 $Y2=1.975
r134 21 22 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.64 $Y=1.89
+ $X2=1.22 $Y2=1.89
r135 20 22 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.11 $Y=1.805
+ $X2=1.22 $Y2=1.89
r136 20 37 25.1442 $w=2.18e-07 $l=4.8e-07 $layer=LI1_cond $X=1.11 $Y=1.805
+ $X2=1.11 $Y2=1.325
r137 16 48 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.98 $Y2=1.202
r138 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.98 $Y2=1.985
r139 13 47 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=1.202
r140 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=0.56
r141 10 46 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.41
+ $X2=0.51 $Y2=1.202
r142 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.51 $Y=1.41
+ $X2=0.51 $Y2=1.985
r143 7 45 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=1.202
r144 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=0.56
r145 2 39 600 $w=1.7e-07 $l=4.88518e-07 $layer=licon1_PDIFF $count=1 $X=2.66
+ $Y=1.845 $X2=2.785 $Y2=2.275
r146 1 31 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.06
+ $Y=0.235 $X2=3.195 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_2%A1_N 1 3 6 8 9
c35 1 0 1.9249e-19 $X=1.615 $Y=1.41
r36 8 9 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.63 $Y=1.16 $X2=1.63
+ $Y2=1.53
r37 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.53
+ $Y=1.16 $X2=1.53 $Y2=1.16
r38 4 13 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.64 $Y=0.995
+ $X2=1.555 $Y2=1.16
r39 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.64 $Y=0.995 $X2=1.64
+ $Y2=0.445
r40 1 13 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=1.615 $Y=1.41
+ $X2=1.555 $Y2=1.16
r41 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.615 $Y=1.41
+ $X2=1.615 $Y2=1.805
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_2%A2_N 1 3 6 8
r32 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.08
+ $Y=1.16 $X2=2.08 $Y2=1.16
r33 4 11 38.532 $w=3.11e-07 $l=1.72337e-07 $layer=POLY_cond $X=2.11 $Y=0.995
+ $X2=2.095 $Y2=1.16
r34 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.11 $Y=0.995 $X2=2.11
+ $Y2=0.445
r35 1 11 47.2262 $w=3.11e-07 $l=2.82843e-07 $layer=POLY_cond $X=2.025 $Y=1.41
+ $X2=2.095 $Y2=1.16
r36 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.025 $Y=1.41
+ $X2=2.025 $Y2=1.805
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_2%A_343_47# 1 2 7 9 10 11 12 14 17 19 20 21
+ 26 30
c65 26 0 4.12944e-20 $X=2.625 $Y=1.155
c66 10 0 6.26351e-20 $X=3.02 $Y=1.435
r67 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.625
+ $Y=1.155 $X2=2.625 $Y2=1.155
r68 24 26 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.625 $Y=1.545
+ $X2=2.625 $Y2=1.155
r69 23 26 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.625 $Y=0.825
+ $X2=2.625 $Y2=1.155
r70 22 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.345 $Y=1.63
+ $X2=2.26 $Y2=1.63
r71 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.54 $Y=1.63
+ $X2=2.625 $Y2=1.545
r72 21 22 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.54 $Y=1.63
+ $X2=2.345 $Y2=1.63
r73 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.54 $Y=0.74
+ $X2=2.625 $Y2=0.825
r74 19 20 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.54 $Y=0.74
+ $X2=1.935 $Y2=0.74
r75 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.85 $Y=0.655
+ $X2=1.935 $Y2=0.74
r76 15 17 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.85 $Y=0.655
+ $X2=1.85 $Y2=0.445
r77 12 14 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.02 $Y=1.77
+ $X2=3.02 $Y2=2.165
r78 11 12 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.02 $Y=1.67 $X2=3.02
+ $Y2=1.77
r79 10 27 45.54 $w=6.04e-07 $l=3.7229e-07 $layer=POLY_cond $X=3.02 $Y=1.435
+ $X2=2.805 $Y2=1.155
r80 10 11 77.9206 $w=2e-07 $l=2.35e-07 $layer=POLY_cond $X=3.02 $Y=1.435
+ $X2=3.02 $Y2=1.67
r81 7 27 62.6463 $w=6.04e-07 $l=4.71487e-07 $layer=POLY_cond $X=2.985 $Y=0.765
+ $X2=2.805 $Y2=1.155
r82 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.985 $Y=0.765
+ $X2=2.985 $Y2=0.445
r83 2 30 600 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=1.485 $X2=2.26 $Y2=1.71
r84 1 17 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.715
+ $Y=0.235 $X2=1.85 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_2%B2 3 5 7 8
c36 5 0 1.72109e-19 $X=3.525 $Y=1.77
c37 3 0 4.12944e-20 $X=3.405 $Y=0.445
r38 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.465
+ $Y=1.47 $X2=3.465 $Y2=1.47
r39 5 11 57.2494 $w=2.85e-07 $l=3.17017e-07 $layer=POLY_cond $X=3.525 $Y=1.77
+ $X2=3.49 $Y2=1.47
r40 5 7 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.525 $Y=1.77
+ $X2=3.525 $Y2=2.165
r41 1 11 38.666 $w=2.85e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.405 $Y=1.305
+ $X2=3.49 $Y2=1.47
r42 1 3 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.405 $Y=1.305
+ $X2=3.405 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_2%B1 3 6 7 9 10 11 12 17
r31 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.165
+ $Y=1.16 $X2=4.165 $Y2=1.16
r32 17 19 27.7763 $w=2.95e-07 $l=1.7e-07 $layer=POLY_cond $X=3.995 $Y=1.16
+ $X2=4.165 $Y2=1.16
r33 11 12 10.4488 $w=3.73e-07 $l=3.4e-07 $layer=LI1_cond $X=4.267 $Y=1.19
+ $X2=4.267 $Y2=1.53
r34 11 20 0.921954 $w=3.73e-07 $l=3e-08 $layer=LI1_cond $X=4.267 $Y=1.19
+ $X2=4.267 $Y2=1.16
r35 10 20 9.52686 $w=3.73e-07 $l=3.1e-07 $layer=LI1_cond $X=4.267 $Y=0.85
+ $X2=4.267 $Y2=1.16
r36 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.995 $Y=1.77
+ $X2=3.995 $Y2=2.165
r37 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.995 $Y=1.67 $X2=3.995
+ $Y2=1.77
r38 5 17 11.9023 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.325
+ $X2=3.995 $Y2=1.16
r39 5 6 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=3.995 $Y=1.325
+ $X2=3.995 $Y2=1.67
r40 1 17 19.6068 $w=2.95e-07 $l=2.16852e-07 $layer=POLY_cond $X=3.875 $Y=0.995
+ $X2=3.995 $Y2=1.16
r41 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.875 $Y=0.995
+ $X2=3.875 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_2%VPWR 1 2 3 12 16 19 20 21 24 26 39 40 48
+ 51 59
c66 12 0 1.9249e-19 $X=1.215 $Y=2.32
r67 51 54 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.27 $Y=1.64
+ $X2=0.27 $Y2=2.32
r68 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r69 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r70 37 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r71 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r72 34 37 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r73 34 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r74 33 36 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r75 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r76 31 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.38 $Y=2.72 $X2=1.19
+ $Y2=2.72
r77 31 33 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.38 $Y=2.72
+ $X2=1.61 $Y2=2.72
r78 30 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r79 30 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r80 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r81 27 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.355 $Y=2.72
+ $X2=0.69 $Y2=2.72
r82 26 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1 $Y=2.72 $X2=1.19
+ $Y2=2.72
r83 26 29 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1 $Y=2.72 $X2=0.69
+ $Y2=2.72
r84 24 59 0.00569083 $w=4.8e-07 $l=2e-08 $layer=MET1_cond $X=0.21 $Y=2.72
+ $X2=0.23 $Y2=2.72
r85 21 54 14.7307 $w=2.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.27 $Y=2.635
+ $X2=0.27 $Y2=2.32
r86 21 27 3.40825 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.177 $Y=2.72
+ $X2=0.355 $Y2=2.72
r87 21 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r88 19 36 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.675 $Y=2.72
+ $X2=3.45 $Y2=2.72
r89 19 20 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.675 $Y=2.72
+ $X2=3.8 $Y2=2.72
r90 18 39 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.925 $Y=2.72
+ $X2=4.37 $Y2=2.72
r91 18 20 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.925 $Y=2.72
+ $X2=3.8 $Y2=2.72
r92 14 20 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.8 $Y=2.635
+ $X2=3.8 $Y2=2.72
r93 14 16 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.8 $Y=2.635
+ $X2=3.8 $Y2=2.34
r94 10 48 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=2.635
+ $X2=1.19 $Y2=2.72
r95 10 12 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=1.19 $Y=2.635
+ $X2=1.19 $Y2=2.32
r96 3 16 600 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=1 $X=3.615
+ $Y=1.845 $X2=3.76 $Y2=2.34
r97 2 12 600 $w=1.7e-07 $l=9.04599e-07 $layer=licon1_PDIFF $count=1 $X=1.07
+ $Y=1.485 $X2=1.215 $Y2=2.32
r98 1 54 400 $w=1.7e-07 $l=8.95321e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=2.32
r99 1 51 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=1.64
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_2%X 1 2 10 11 12 13 14 15 24
r27 14 15 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=0.677 $Y=1.87
+ $X2=0.677 $Y2=2.21
r28 14 24 4.15635 $w=3.03e-07 $l=1.1e-07 $layer=LI1_cond $X=0.677 $Y=1.87
+ $X2=0.677 $Y2=1.76
r29 11 24 3.13616 $w=3.03e-07 $l=8.3e-08 $layer=LI1_cond $X=0.677 $Y=1.677
+ $X2=0.677 $Y2=1.76
r30 11 12 6.65738 $w=3.03e-07 $l=1.52e-07 $layer=LI1_cond $X=0.677 $Y=1.677
+ $X2=0.677 $Y2=1.525
r31 10 12 37.4544 $w=2.18e-07 $l=7.15e-07 $layer=LI1_cond $X=0.635 $Y=0.81
+ $X2=0.635 $Y2=1.525
r32 9 13 5.59218 $w=3.03e-07 $l=1.48e-07 $layer=LI1_cond $X=0.677 $Y=0.658
+ $X2=0.677 $Y2=0.51
r33 9 10 6.65738 $w=3.03e-07 $l=1.52e-07 $layer=LI1_cond $X=0.677 $Y=0.658
+ $X2=0.677 $Y2=0.81
r34 2 24 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.6
+ $Y=1.485 $X2=0.745 $Y2=1.76
r35 1 13 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.235 $X2=0.745 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_2%A_622_369# 1 2 8 9 10 13 16
r32 11 13 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.23 $Y=2.005
+ $X2=4.23 $Y2=2.275
r33 9 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.145 $Y=1.92
+ $X2=4.23 $Y2=2.005
r34 9 10 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.145 $Y=1.92
+ $X2=3.455 $Y2=1.92
r35 8 16 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.37 $Y=2.255
+ $X2=3.29 $Y2=2.34
r36 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.37 $Y=2.005
+ $X2=3.455 $Y2=1.92
r37 7 8 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.37 $Y=2.005 $X2=3.37
+ $Y2=2.255
r38 2 13 600 $w=1.7e-07 $l=4.97242e-07 $layer=licon1_PDIFF $count=1 $X=4.085
+ $Y=1.845 $X2=4.23 $Y2=2.275
r39 1 16 600 $w=1.7e-07 $l=5.78035e-07 $layer=licon1_PDIFF $count=1 $X=3.11
+ $Y=1.845 $X2=3.29 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2O_2%VGND 1 2 3 4 13 15 17 20 22 32 44 52 55
+ 58 62 68
c61 32 0 6.26351e-20 $X=3.905 $Y=0
r62 58 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r63 57 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r64 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r65 54 55 9.96101 $w=5.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=0.2
+ $X2=2.89 $Y2=0.2
r66 50 54 4.09185 $w=5.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.53 $Y=0.2
+ $X2=2.725 $Y2=0.2
r67 50 52 14.3676 $w=5.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.53 $Y=0.2
+ $X2=2.155 $Y2=0.2
r68 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r69 44 47 11.0886 $w=4.78e-07 $l=4.45e-07 $layer=LI1_cond $X=1.24 $Y=0 $X2=1.24
+ $Y2=0.445
r70 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r71 36 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r72 36 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r73 35 55 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=2.89
+ $Y2=0
r74 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r75 32 57 5.5149 $w=1.7e-07 $l=3.47e-07 $layer=LI1_cond $X=3.905 $Y=0 $X2=4.252
+ $Y2=0
r76 32 35 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=3.905 $Y=0 $X2=2.99
+ $Y2=0
r77 31 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r78 31 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r79 30 52 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.155
+ $Y2=0
r80 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r81 28 44 6.90116 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=1.48 $Y=0 $X2=1.24
+ $Y2=0
r82 28 30 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.48 $Y=0 $X2=2.07
+ $Y2=0
r83 26 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r84 26 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r85 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r86 23 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.69
+ $Y2=0
r87 22 44 6.90116 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=1 $Y=0 $X2=1.24 $Y2=0
r88 22 25 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1 $Y=0 $X2=0.69
+ $Y2=0
r89 20 68 0.00569083 $w=4.8e-07 $l=2e-08 $layer=MET1_cond $X=0.21 $Y=0 $X2=0.23
+ $Y2=0
r90 17 62 13.9075 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.38
r91 17 23 3.40825 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.177 $Y=0 $X2=0.355
+ $Y2=0
r92 17 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r93 13 57 3.28987 $w=4.5e-07 $l=1.58915e-07 $layer=LI1_cond $X=4.13 $Y=0.085
+ $X2=4.252 $Y2=0
r94 13 15 9.16993 $w=4.48e-07 $l=3.45e-07 $layer=LI1_cond $X=4.13 $Y=0.085
+ $X2=4.13 $Y2=0.43
r95 4 15 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=3.95
+ $Y=0.235 $X2=4.135 $Y2=0.43
r96 3 54 91 $w=1.7e-07 $l=6.17009e-07 $layer=licon1_NDIFF $count=2 $X=2.185
+ $Y=0.235 $X2=2.725 $Y2=0.4
r97 2 47 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.235 $X2=1.215 $Y2=0.445
r98 1 62 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.235 $X2=0.27 $Y2=0.38
.ends

