* File: sky130_fd_sc_hdll__muxb8to1_2.spice
* Created: Thu Aug 27 19:12:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__muxb8to1_2.pex.spice"
.subckt sky130_fd_sc_hdll__muxb8to1_2  VNB VPB D[0] S[0] S[1] D[1] D[2] S[2]
+ S[3] D[3] D[4] S[4] S[5] D[5] D[6] S[6] S[7] D[7] VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* D[7]	D[7]
* S[7]	S[7]
* S[6]	S[6]
* D[6]	D[6]
* D[5]	D[5]
* S[5]	S[5]
* S[4]	S[4]
* D[4]	D[4]
* D[3]	D[3]
* S[3]	S[3]
* S[2]	S[2]
* D[2]	D[2]
* D[1]	D[1]
* S[1]	S[1]
* S[0]	S[0]
* D[0]	D[0]
* VPB	VPB
* VNB	VNB
MM1019 N_A_27_47#_M1019_d N_D[0]_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1053 N_A_27_47#_M1053_d N_D[0]_M1053_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.128194 AS=0.08775 PD=1.13333 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1017 N_A_27_47#_M1053_d N_S[0]_M1017_g N_Z_M1017_s VNB NSHORT L=0.15 W=0.52
+ AD=0.102556 AS=0.0702 PD=0.906667 PS=0.79 NRD=16.728 NRS=0 M=1 R=3.46667
+ SA=75001.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1020 N_A_27_47#_M1020_d N_S[0]_M1020_g N_Z_M1017_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1043 N_VGND_M1043_d N_S[0]_M1043_g N_A_278_265#_M1043_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1035 N_A_701_47#_M1035_d N_S[1]_M1035_g N_VGND_M1043_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1015 N_A_845_69#_M1015_d N_S[1]_M1015_g N_Z_M1015_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.6 A=0.078 P=1.34 MULT=1
MM1018 N_A_845_69#_M1018_d N_S[1]_M1018_g N_Z_M1015_s VNB NSHORT L=0.15 W=0.52
+ AD=0.102556 AS=0.0702 PD=0.906667 PS=0.79 NRD=16.728 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75001.2 A=0.078 P=1.34 MULT=1
MM1036 N_VGND_M1036_d N_D[1]_M1036_g N_A_845_69#_M1018_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.128194 PD=0.92 PS=1.13333 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75000.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1051 N_VGND_M1036_d N_D[1]_M1051_g N_A_845_69#_M1051_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1057 N_A_1315_47#_M1057_d N_D[2]_M1057_g N_VGND_M1057_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1063 N_A_1315_47#_M1063_d N_D[2]_M1063_g N_VGND_M1057_s VNB NSHORT L=0.15
+ W=0.65 AD=0.128194 AS=0.08775 PD=1.13333 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1058 N_Z_M1058_d N_S[2]_M1058_g N_A_1315_47#_M1063_d VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1 R=3.46667
+ SA=75001.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1076 N_Z_M1058_d N_S[2]_M1076_g N_A_1315_47#_M1076_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1077 N_VGND_M1077_d N_S[2]_M1077_g N_A_1566_265#_M1077_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1009 N_A_1989_47#_M1009_d N_S[3]_M1009_g N_VGND_M1077_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1052 N_Z_M1052_d N_S[3]_M1052_g N_A_2133_69#_M1052_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.6 A=0.078 P=1.34 MULT=1
MM1065 N_Z_M1052_d N_S[3]_M1065_g N_A_2133_69#_M1065_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1 R=3.46667
+ SA=75000.6 SB=75001.2 A=0.078 P=1.34 MULT=1
MM1012 N_A_2133_69#_M1065_s N_D[3]_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15
+ W=0.65 AD=0.128194 AS=0.08775 PD=1.13333 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1078 N_A_2133_69#_M1078_d N_D[3]_M1078_g N_VGND_M1012_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1031 N_VGND_M1031_d N_D[4]_M1031_g N_A_2603_47#_M1031_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1048 N_VGND_M1031_d N_D[4]_M1048_g N_A_2603_47#_M1048_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.128194 PD=0.92 PS=1.13333 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75000.7 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1021 N_Z_M1021_d N_S[4]_M1021_g N_A_2603_47#_M1048_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1 R=3.46667
+ SA=75001.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1044 N_Z_M1021_d N_S[4]_M1044_g N_A_2603_47#_M1044_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1032 N_VGND_M1032_d N_S[4]_M1032_g N_A_2854_265#_M1032_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1050 N_A_3277_47#_M1050_d N_S[5]_M1050_g N_VGND_M1032_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1010 N_Z_M1010_d N_S[5]_M1010_g N_A_3421_69#_M1010_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.6 A=0.078 P=1.34 MULT=1
MM1026 N_Z_M1010_d N_S[5]_M1026_g N_A_3421_69#_M1026_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1 R=3.46667
+ SA=75000.6 SB=75001.2 A=0.078 P=1.34 MULT=1
MM1047 N_VGND_M1047_d N_D[5]_M1047_g N_A_3421_69#_M1026_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.128194 PD=0.92 PS=1.13333 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75000.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1054 N_VGND_M1047_d N_D[5]_M1054_g N_A_3421_69#_M1054_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1070 N_VGND_M1070_d N_D[6]_M1070_g N_A_3891_47#_M1070_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1079 N_VGND_M1070_d N_D[6]_M1079_g N_A_3891_47#_M1079_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.128194 PD=0.92 PS=1.13333 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75000.7 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1059 N_Z_M1059_d N_S[6]_M1059_g N_A_3891_47#_M1079_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1 R=3.46667
+ SA=75001.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1074 N_Z_M1059_d N_S[6]_M1074_g N_A_3891_47#_M1074_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1075 N_VGND_M1075_d N_S[6]_M1075_g N_A_4142_265#_M1075_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1007 N_A_4565_47#_M1007_d N_S[7]_M1007_g N_VGND_M1075_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1055 N_Z_M1055_d N_S[7]_M1055_g N_A_4709_69#_M1055_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.6 A=0.078 P=1.34 MULT=1
MM1071 N_Z_M1055_d N_S[7]_M1071_g N_A_4709_69#_M1071_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1 R=3.46667
+ SA=75000.6 SB=75001.2 A=0.078 P=1.34 MULT=1
MM1011 N_A_4709_69#_M1071_s N_D[7]_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.128194 AS=0.08775 PD=1.13333 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1027 N_A_4709_69#_M1027_d N_D[7]_M1027_g N_VGND_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_A_27_297#_M1003_d N_D[0]_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1034 N_A_27_297#_M1034_d N_D[0]_M1034_g N_VPWR_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001 A=0.18 P=2.36 MULT=1
MM1006 N_A_27_297#_M1034_d N_A_278_265#_M1006_g N_Z_M1006_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182 M=1
+ R=4.55556 SA=90001.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1013 N_A_27_297#_M1013_d N_A_278_265#_M1013_g N_Z_M1006_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1008 N_VPWR_M1008_d N_S[0]_M1008_g N_A_278_265#_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.18 AS=0.27 PD=1.36 PS=2.54 NRD=7.8603 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1045 N_A_701_47#_M1045_d N_S[1]_M1045_g N_VPWR_M1008_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.18 PD=2.54 PS=1.36 NRD=0.9653 NRS=7.8603 M=1 R=5.55556 SA=90000.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1040 N_A_824_333#_M1040_d N_A_701_47#_M1040_g N_Z_M1040_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1056 N_A_824_333#_M1056_d N_A_701_47#_M1056_g N_Z_M1040_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.2 A=0.1476 P=2 MULT=1
MM1022 N_A_824_333#_M1056_d N_D[1]_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1049 N_A_824_333#_M1049_d N_D[1]_M1049_g N_VPWR_M1022_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_D[2]_M1000_g N_A_1315_297#_M1000_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1060 N_VPWR_M1000_d N_D[2]_M1060_g N_A_1315_297#_M1060_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.181154 PD=1.29 PS=1.47802 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.6 SB=90001 A=0.18 P=2.36 MULT=1
MM1004 N_Z_M1004_d N_A_1566_265#_M1004_g N_A_1315_297#_M1060_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.148546 PD=1.11 PS=1.21198 NRD=1.182 NRS=14.4007
+ M=1 R=4.55556 SA=90001.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1061 N_Z_M1004_d N_A_1566_265#_M1061_g N_A_1315_297#_M1061_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1067 N_VPWR_M1067_d N_S[2]_M1067_g N_A_1566_265#_M1067_s VPB PHIGHVT L=0.18
+ W=1 AD=0.18 AS=0.27 PD=1.36 PS=2.54 NRD=7.8603 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1023 N_A_1989_47#_M1023_d N_S[3]_M1023_g N_VPWR_M1067_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.18 PD=2.54 PS=1.36 NRD=0.9653 NRS=7.8603 M=1 R=5.55556 SA=90000.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1005 N_Z_M1005_d N_A_1989_47#_M1005_g N_A_2112_333#_M1005_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1062 N_Z_M1005_d N_A_1989_47#_M1062_g N_A_2112_333#_M1062_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.148546 PD=1.11 PS=1.21198 NRD=1.182 NRS=14.4007 M=1
+ R=4.55556 SA=90000.6 SB=90001.2 A=0.1476 P=2 MULT=1
MM1001 N_VPWR_M1001_d N_D[3]_M1001_g N_A_2112_333#_M1062_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.181154 PD=1.29 PS=1.47802 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1068 N_VPWR_M1001_d N_D[3]_M1068_g N_A_2112_333#_M1068_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1014 N_A_2603_297#_M1014_d N_D[4]_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1037 N_A_2603_297#_M1037_d N_D[4]_M1037_g N_VPWR_M1014_s VPB PHIGHVT L=0.18
+ W=1 AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.6 SB=90001 A=0.18 P=2.36 MULT=1
MM1016 N_A_2603_297#_M1037_d N_A_2854_265#_M1016_g N_Z_M1016_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182
+ M=1 R=4.55556 SA=90001.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1041 N_A_2603_297#_M1041_d N_A_2854_265#_M1041_g N_Z_M1016_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1002 N_VPWR_M1002_d N_S[4]_M1002_g N_A_2854_265#_M1002_s VPB PHIGHVT L=0.18
+ W=1 AD=0.18 AS=0.27 PD=1.36 PS=2.54 NRD=7.8603 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1028 N_A_3277_47#_M1028_d N_S[5]_M1028_g N_VPWR_M1002_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.18 PD=2.54 PS=1.36 NRD=0.9653 NRS=7.8603 M=1 R=5.55556 SA=90000.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1024 N_A_3400_333#_M1024_d N_A_3277_47#_M1024_g N_Z_M1024_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1042 N_A_3400_333#_M1042_d N_A_3277_47#_M1042_g N_Z_M1024_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.2 A=0.1476 P=2 MULT=1
MM1025 N_A_3400_333#_M1042_d N_D[5]_M1025_g N_VPWR_M1025_s VPB PHIGHVT L=0.18
+ W=1 AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1038 N_A_3400_333#_M1038_d N_D[5]_M1038_g N_VPWR_M1025_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1029 N_A_3891_297#_M1029_d N_D[6]_M1029_g N_VPWR_M1029_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1072 N_A_3891_297#_M1072_d N_D[6]_M1072_g N_VPWR_M1029_s VPB PHIGHVT L=0.18
+ W=1 AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.6 SB=90001 A=0.18 P=2.36 MULT=1
MM1033 N_A_3891_297#_M1072_d N_A_4142_265#_M1033_g N_Z_M1033_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182
+ M=1 R=4.55556 SA=90001.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1046 N_A_3891_297#_M1046_d N_A_4142_265#_M1046_g N_Z_M1033_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1039 N_VPWR_M1039_d N_S[6]_M1039_g N_A_4142_265#_M1039_s VPB PHIGHVT L=0.18
+ W=1 AD=0.18 AS=0.27 PD=1.36 PS=2.54 NRD=7.8603 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1066 N_A_4565_47#_M1066_d N_S[7]_M1066_g N_VPWR_M1039_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.18 PD=2.54 PS=1.36 NRD=0.9653 NRS=7.8603 M=1 R=5.55556 SA=90000.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1064 N_A_4688_333#_M1064_d N_A_4565_47#_M1064_g N_Z_M1064_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1073 N_A_4688_333#_M1073_d N_A_4565_47#_M1073_g N_Z_M1064_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.2 A=0.1476 P=2 MULT=1
MM1030 N_A_4688_333#_M1073_d N_D[7]_M1030_g N_VPWR_M1030_s VPB PHIGHVT L=0.18
+ W=1 AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1069 N_A_4688_333#_M1069_d N_D[7]_M1069_g N_VPWR_M1030_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.5 SB=90000.2 A=0.18 P=2.36 MULT=1
DX80_noxref VNB VPB NWDIODE A=41.9547 P=55.49
c_255 VNB 0 0.00145591f $X=25.445 $Y=-0.085
*
.include "sky130_fd_sc_hdll__muxb8to1_2.pxi.spice"
*
.ends
*
*
