* File: sky130_fd_sc_hdll__xnor3_4.pxi.spice
* Created: Thu Aug 27 19:29:37 2020
* 
x_PM_SKY130_FD_SC_HDLL__XNOR3_4%A_101_21# N_A_101_21#_M1023_d
+ N_A_101_21#_M1019_d N_A_101_21#_c_168_n N_A_101_21#_M1005_g
+ N_A_101_21#_c_177_n N_A_101_21#_M1000_g N_A_101_21#_c_169_n
+ N_A_101_21#_M1007_g N_A_101_21#_c_178_n N_A_101_21#_M1012_g
+ N_A_101_21#_c_170_n N_A_101_21#_M1009_g N_A_101_21#_c_179_n
+ N_A_101_21#_M1022_g N_A_101_21#_c_171_n N_A_101_21#_M1017_g
+ N_A_101_21#_c_180_n N_A_101_21#_M1024_g N_A_101_21#_c_172_n
+ N_A_101_21#_c_181_n N_A_101_21#_c_188_p N_A_101_21#_c_193_p
+ N_A_101_21#_c_224_p N_A_101_21#_c_173_n N_A_101_21#_c_182_n
+ N_A_101_21#_c_174_n N_A_101_21#_c_183_n N_A_101_21#_c_184_n
+ N_A_101_21#_c_197_p N_A_101_21#_c_208_p N_A_101_21#_c_175_n
+ N_A_101_21#_c_176_n PM_SKY130_FD_SC_HDLL__XNOR3_4%A_101_21#
x_PM_SKY130_FD_SC_HDLL__XNOR3_4%C N_C_c_310_n N_C_M1026_g N_C_M1002_g
+ N_C_c_311_n N_C_M1019_g N_C_c_312_n N_C_M1023_g N_C_c_313_n N_C_c_314_n C
+ N_C_c_335_n C PM_SKY130_FD_SC_HDLL__XNOR3_4%C
x_PM_SKY130_FD_SC_HDLL__XNOR3_4%A_532_93# N_A_532_93#_M1026_d
+ N_A_532_93#_M1002_d N_A_532_93#_c_370_n N_A_532_93#_M1025_g
+ N_A_532_93#_c_371_n N_A_532_93#_M1020_g N_A_532_93#_c_386_n
+ N_A_532_93#_c_372_n N_A_532_93#_c_376_n N_A_532_93#_c_377_n
+ N_A_532_93#_c_378_n N_A_532_93#_c_373_n
+ PM_SKY130_FD_SC_HDLL__XNOR3_4%A_532_93#
x_PM_SKY130_FD_SC_HDLL__XNOR3_4%A_1089_297# N_A_1089_297#_M1004_d
+ N_A_1089_297#_M1027_d N_A_1089_297#_c_456_n N_A_1089_297#_M1021_g
+ N_A_1089_297#_M1011_g N_A_1089_297#_c_443_n N_A_1089_297#_c_444_n
+ N_A_1089_297#_c_458_n N_A_1089_297#_M1010_g N_A_1089_297#_c_445_n
+ N_A_1089_297#_M1015_g N_A_1089_297#_c_446_n N_A_1089_297#_c_447_n
+ N_A_1089_297#_c_461_n N_A_1089_297#_c_448_n N_A_1089_297#_c_449_n
+ N_A_1089_297#_c_465_p N_A_1089_297#_c_450_n N_A_1089_297#_c_451_n
+ N_A_1089_297#_c_452_n N_A_1089_297#_c_453_n N_A_1089_297#_c_454_n
+ N_A_1089_297#_c_455_n PM_SKY130_FD_SC_HDLL__XNOR3_4%A_1089_297#
x_PM_SKY130_FD_SC_HDLL__XNOR3_4%B N_B_c_630_n N_B_M1027_g N_B_M1004_g
+ N_B_c_623_n N_B_c_624_n N_B_M1008_g N_B_M1006_g N_B_c_633_n N_B_c_634_n
+ N_B_M1014_g N_B_c_635_n N_B_c_636_n N_B_M1016_g N_B_c_626_n N_B_c_627_n
+ N_B_c_628_n N_B_c_641_n B N_B_c_629_n B PM_SKY130_FD_SC_HDLL__XNOR3_4%B
x_PM_SKY130_FD_SC_HDLL__XNOR3_4%A N_A_c_756_n N_A_M1018_g N_A_c_757_n
+ N_A_M1003_g A PM_SKY130_FD_SC_HDLL__XNOR3_4%A
x_PM_SKY130_FD_SC_HDLL__XNOR3_4%A_1207_297# N_A_1207_297#_M1006_s
+ N_A_1207_297#_M1015_d N_A_1207_297#_M1008_s N_A_1207_297#_M1010_d
+ N_A_1207_297#_c_794_n N_A_1207_297#_M1013_g N_A_1207_297#_c_795_n
+ N_A_1207_297#_M1001_g N_A_1207_297#_c_796_n N_A_1207_297#_c_809_n
+ N_A_1207_297#_c_803_n N_A_1207_297#_c_797_n N_A_1207_297#_c_798_n
+ N_A_1207_297#_c_799_n N_A_1207_297#_c_805_n N_A_1207_297#_c_814_n
+ N_A_1207_297#_c_800_n N_A_1207_297#_c_801_n N_A_1207_297#_c_829_n
+ N_A_1207_297#_c_830_n PM_SKY130_FD_SC_HDLL__XNOR3_4%A_1207_297#
x_PM_SKY130_FD_SC_HDLL__XNOR3_4%VPWR N_VPWR_M1000_s N_VPWR_M1012_s
+ N_VPWR_M1024_s N_VPWR_M1027_s N_VPWR_M1018_d N_VPWR_c_930_n N_VPWR_c_931_n
+ N_VPWR_c_932_n N_VPWR_c_933_n N_VPWR_c_934_n N_VPWR_c_935_n N_VPWR_c_936_n
+ N_VPWR_c_937_n N_VPWR_c_938_n N_VPWR_c_939_n N_VPWR_c_940_n VPWR
+ N_VPWR_c_941_n N_VPWR_c_942_n N_VPWR_c_929_n N_VPWR_c_944_n N_VPWR_c_945_n
+ PM_SKY130_FD_SC_HDLL__XNOR3_4%VPWR
x_PM_SKY130_FD_SC_HDLL__XNOR3_4%X N_X_M1005_s N_X_M1009_s N_X_M1000_d
+ N_X_M1022_d N_X_c_1046_n N_X_c_1051_n N_X_c_1055_n N_X_c_1056_n N_X_c_1057_n
+ N_X_c_1047_n X N_X_c_1067_n PM_SKY130_FD_SC_HDLL__XNOR3_4%X
x_PM_SKY130_FD_SC_HDLL__XNOR3_4%A_657_325# N_A_657_325#_M1020_d
+ N_A_657_325#_M1006_d N_A_657_325#_M1019_s N_A_657_325#_M1016_d
+ N_A_657_325#_c_1095_n N_A_657_325#_c_1090_n N_A_657_325#_c_1091_n
+ N_A_657_325#_c_1092_n N_A_657_325#_c_1097_n N_A_657_325#_c_1098_n
+ N_A_657_325#_c_1099_n N_A_657_325#_c_1100_n N_A_657_325#_c_1093_n
+ N_A_657_325#_c_1102_n N_A_657_325#_c_1139_n N_A_657_325#_c_1094_n
+ N_A_657_325#_c_1103_n N_A_657_325#_c_1142_n N_A_657_325#_c_1104_n
+ PM_SKY130_FD_SC_HDLL__XNOR3_4%A_657_325#
x_PM_SKY130_FD_SC_HDLL__XNOR3_4%A_681_49# N_A_681_49#_M1023_s
+ N_A_681_49#_M1014_d N_A_681_49#_M1025_d N_A_681_49#_M1008_d
+ N_A_681_49#_c_1257_n N_A_681_49#_c_1245_n N_A_681_49#_c_1249_n
+ N_A_681_49#_c_1286_n N_A_681_49#_c_1250_n N_A_681_49#_c_1246_n
+ N_A_681_49#_c_1364_p N_A_681_49#_c_1299_n N_A_681_49#_c_1300_n
+ N_A_681_49#_c_1247_n N_A_681_49#_c_1321_n N_A_681_49#_c_1252_n
+ N_A_681_49#_c_1253_n N_A_681_49#_c_1254_n N_A_681_49#_c_1255_n
+ PM_SKY130_FD_SC_HDLL__XNOR3_4%A_681_49#
x_PM_SKY130_FD_SC_HDLL__XNOR3_4%A_1490_297# N_A_1490_297#_M1011_d
+ N_A_1490_297#_M1001_d N_A_1490_297#_M1021_d N_A_1490_297#_M1013_d
+ N_A_1490_297#_c_1380_n N_A_1490_297#_c_1392_n N_A_1490_297#_c_1384_n
+ N_A_1490_297#_c_1381_n N_A_1490_297#_c_1393_n N_A_1490_297#_c_1386_n
+ N_A_1490_297#_c_1382_n PM_SKY130_FD_SC_HDLL__XNOR3_4%A_1490_297#
x_PM_SKY130_FD_SC_HDLL__XNOR3_4%VGND N_VGND_M1005_d N_VGND_M1007_d
+ N_VGND_M1017_d N_VGND_M1004_s N_VGND_M1003_d N_VGND_c_1446_n N_VGND_c_1447_n
+ N_VGND_c_1448_n N_VGND_c_1449_n N_VGND_c_1450_n N_VGND_c_1451_n
+ N_VGND_c_1452_n N_VGND_c_1453_n N_VGND_c_1454_n N_VGND_c_1455_n
+ N_VGND_c_1456_n N_VGND_c_1457_n VGND N_VGND_c_1458_n N_VGND_c_1459_n
+ N_VGND_c_1460_n N_VGND_c_1461_n N_VGND_c_1462_n
+ PM_SKY130_FD_SC_HDLL__XNOR3_4%VGND
cc_1 VNB N_A_101_21#_c_168_n 0.0219887f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.995
cc_2 VNB N_A_101_21#_c_169_n 0.0170092f $X=-0.19 $Y=-0.24 $X2=1.05 $Y2=0.995
cc_3 VNB N_A_101_21#_c_170_n 0.0165817f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=0.995
cc_4 VNB N_A_101_21#_c_171_n 0.0183996f $X=-0.19 $Y=-0.24 $X2=2 $Y2=0.995
cc_5 VNB N_A_101_21#_c_172_n 0.00109516f $X=-0.19 $Y=-0.24 $X2=2.175 $Y2=1.325
cc_6 VNB N_A_101_21#_c_173_n 0.00138296f $X=-0.19 $Y=-0.24 $X2=2.625 $Y2=0.695
cc_7 VNB N_A_101_21#_c_174_n 0.00216705f $X=-0.19 $Y=-0.24 $X2=2.735 $Y2=0.34
cc_8 VNB N_A_101_21#_c_175_n 0.0163051f $X=-0.19 $Y=-0.24 $X2=3.7 $Y2=0.355
cc_9 VNB N_A_101_21#_c_176_n 0.0999705f $X=-0.19 $Y=-0.24 $X2=2.045 $Y2=1.202
cc_10 VNB N_C_c_310_n 0.0199971f $X=-0.19 $Y=-0.24 $X2=3.875 $Y2=0.245
cc_11 VNB N_C_c_311_n 0.0145755f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.56
cc_12 VNB N_C_c_312_n 0.0221238f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.985
cc_13 VNB N_C_c_313_n 0.011843f $X=-0.19 $Y=-0.24 $X2=1.05 $Y2=0.56
cc_14 VNB N_C_c_314_n 0.0544628f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=1.985
cc_15 VNB N_A_532_93#_c_370_n 0.0252997f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.995
cc_16 VNB N_A_532_93#_c_371_n 0.0211819f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.41
cc_17 VNB N_A_532_93#_c_372_n 0.00260551f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=1.985
cc_18 VNB N_A_532_93#_c_373_n 0.00274123f $X=-0.19 $Y=-0.24 $X2=2.045 $Y2=1.41
cc_19 VNB N_A_1089_297#_M1011_g 0.0360077f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.985
cc_20 VNB N_A_1089_297#_c_443_n 0.029369f $X=-0.19 $Y=-0.24 $X2=1.05 $Y2=0.56
cc_21 VNB N_A_1089_297#_c_444_n 0.001407f $X=-0.19 $Y=-0.24 $X2=1.05 $Y2=0.56
cc_22 VNB N_A_1089_297#_c_445_n 0.0195477f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=0.995
cc_23 VNB N_A_1089_297#_c_446_n 0.0288128f $X=-0.19 $Y=-0.24 $X2=1.575 $Y2=1.41
cc_24 VNB N_A_1089_297#_c_447_n 0.0176837f $X=-0.19 $Y=-0.24 $X2=1.575 $Y2=1.985
cc_25 VNB N_A_1089_297#_c_448_n 0.00239787f $X=-0.19 $Y=-0.24 $X2=2.63 $Y2=1.96
cc_26 VNB N_A_1089_297#_c_449_n 0.00773632f $X=-0.19 $Y=-0.24 $X2=2.625
+ $Y2=0.425
cc_27 VNB N_A_1089_297#_c_450_n 0.0128101f $X=-0.19 $Y=-0.24 $X2=2.74 $Y2=2.045
cc_28 VNB N_A_1089_297#_c_451_n 0.00136794f $X=-0.19 $Y=-0.24 $X2=2.74 $Y2=2.235
cc_29 VNB N_A_1089_297#_c_452_n 0.00305675f $X=-0.19 $Y=-0.24 $X2=3.9 $Y2=0.355
cc_30 VNB N_A_1089_297#_c_453_n 0.00216739f $X=-0.19 $Y=-0.24 $X2=4.02 $Y2=0.37
cc_31 VNB N_A_1089_297#_c_454_n 0.00620483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_1089_297#_c_455_n 0.00259923f $X=-0.19 $Y=-0.24 $X2=1.05 $Y2=1.202
cc_33 VNB N_B_M1004_g 0.0300439f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_B_c_623_n 0.0595974f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.56
cc_35 VNB N_B_c_624_n 0.0273885f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.56
cc_36 VNB N_B_M1006_g 0.0290181f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=1.41
cc_37 VNB N_B_c_626_n 0.010365f $X=-0.19 $Y=-0.24 $X2=2.175 $Y2=1.325
cc_38 VNB N_B_c_627_n 0.00131136f $X=-0.19 $Y=-0.24 $X2=2.63 $Y2=1.96
cc_39 VNB N_B_c_628_n 0.0298429f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=1.96
cc_40 VNB N_B_c_629_n 0.021241f $X=-0.19 $Y=-0.24 $X2=2.735 $Y2=0.34
cc_41 VNB N_A_c_756_n 0.0230531f $X=-0.19 $Y=-0.24 $X2=3.875 $Y2=0.245
cc_42 VNB N_A_c_757_n 0.0182223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB A 0.00406657f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.995
cc_44 VNB N_A_1207_297#_c_794_n 0.0267203f $X=-0.19 $Y=-0.24 $X2=1.05 $Y2=0.995
cc_45 VNB N_A_1207_297#_c_795_n 0.0198808f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=1.41
cc_46 VNB N_A_1207_297#_c_796_n 0.00430585f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=0.995
cc_47 VNB N_A_1207_297#_c_797_n 0.00275527f $X=-0.19 $Y=-0.24 $X2=2 $Y2=0.56
cc_48 VNB N_A_1207_297#_c_798_n 0.0020163f $X=-0.19 $Y=-0.24 $X2=2.045 $Y2=1.41
cc_49 VNB N_A_1207_297#_c_799_n 0.00350271f $X=-0.19 $Y=-0.24 $X2=2.045
+ $Y2=1.985
cc_50 VNB N_A_1207_297#_c_800_n 0.00247723f $X=-0.19 $Y=-0.24 $X2=2.625
+ $Y2=0.695
cc_51 VNB N_A_1207_297#_c_801_n 0.00732735f $X=-0.19 $Y=-0.24 $X2=3.7 $Y2=0.34
cc_52 VNB N_VPWR_c_929_n 0.440529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_X_c_1046_n 9.06365e-19 $X=-0.19 $Y=-0.24 $X2=1.05 $Y2=0.56
cc_54 VNB N_X_c_1047_n 8.41723e-19 $X=-0.19 $Y=-0.24 $X2=2.045 $Y2=1.985
cc_55 VNB N_A_657_325#_c_1090_n 0.0107286f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=1.985
cc_56 VNB N_A_657_325#_c_1091_n 0.0135137f $X=-0.19 $Y=-0.24 $X2=1.575 $Y2=1.41
cc_57 VNB N_A_657_325#_c_1092_n 0.00281469f $X=-0.19 $Y=-0.24 $X2=1.575
+ $Y2=1.985
cc_58 VNB N_A_657_325#_c_1093_n 0.00225677f $X=-0.19 $Y=-0.24 $X2=2.175
+ $Y2=1.875
cc_59 VNB N_A_657_325#_c_1094_n 0.0104433f $X=-0.19 $Y=-0.24 $X2=2.85 $Y2=2.32
cc_60 VNB N_A_681_49#_c_1245_n 0.00873334f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=1.41
cc_61 VNB N_A_681_49#_c_1246_n 0.0097913f $X=-0.19 $Y=-0.24 $X2=1.575 $Y2=1.985
cc_62 VNB N_A_681_49#_c_1247_n 0.00622338f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.78
cc_63 VNB N_A_1490_297#_c_1380_n 0.00788636f $X=-0.19 $Y=-0.24 $X2=1.05 $Y2=0.56
cc_64 VNB N_A_1490_297#_c_1381_n 0.0307904f $X=-0.19 $Y=-0.24 $X2=2 $Y2=0.56
cc_65 VNB N_A_1490_297#_c_1382_n 0.0135316f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=1.96
cc_66 VNB N_VGND_c_1446_n 0.00471684f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=1.985
cc_67 VNB N_VGND_c_1447_n 0.00417754f $X=-0.19 $Y=-0.24 $X2=1.575 $Y2=1.41
cc_68 VNB N_VGND_c_1448_n 0.0171678f $X=-0.19 $Y=-0.24 $X2=1.575 $Y2=1.985
cc_69 VNB N_VGND_c_1449_n 0.00255418f $X=-0.19 $Y=-0.24 $X2=2.045 $Y2=1.41
cc_70 VNB N_VGND_c_1450_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=2.175 $Y2=1.875
cc_71 VNB N_VGND_c_1451_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=1.96
cc_72 VNB N_VGND_c_1452_n 0.0112126f $X=-0.19 $Y=-0.24 $X2=2.74 $Y2=2.045
cc_73 VNB N_VGND_c_1453_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=2.74 $Y2=2.235
cc_74 VNB N_VGND_c_1454_n 0.0222227f $X=-0.19 $Y=-0.24 $X2=3.7 $Y2=0.34
cc_75 VNB N_VGND_c_1455_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=2.735 $Y2=0.34
cc_76 VNB N_VGND_c_1456_n 0.108747f $X=-0.19 $Y=-0.24 $X2=3.945 $Y2=2.32
cc_77 VNB N_VGND_c_1457_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=3.945 $Y2=2.32
cc_78 VNB N_VGND_c_1458_n 0.0678678f $X=-0.19 $Y=-0.24 $X2=2.115 $Y2=1.16
cc_79 VNB N_VGND_c_1459_n 0.0259875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1460_n 0.532607f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1461_n 0.00449846f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1462_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VPB N_A_101_21#_c_177_n 0.0207574f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.41
cc_84 VPB N_A_101_21#_c_178_n 0.0161737f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=1.41
cc_85 VPB N_A_101_21#_c_179_n 0.0161684f $X=-0.19 $Y=1.305 $X2=1.575 $Y2=1.41
cc_86 VPB N_A_101_21#_c_180_n 0.0176334f $X=-0.19 $Y=1.305 $X2=2.045 $Y2=1.41
cc_87 VPB N_A_101_21#_c_181_n 0.00158809f $X=-0.19 $Y=1.305 $X2=2.175 $Y2=1.875
cc_88 VPB N_A_101_21#_c_182_n 0.0038652f $X=-0.19 $Y=1.305 $X2=2.74 $Y2=2.235
cc_89 VPB N_A_101_21#_c_183_n 0.00112766f $X=-0.19 $Y=1.305 $X2=2.85 $Y2=2.32
cc_90 VPB N_A_101_21#_c_184_n 0.0124849f $X=-0.19 $Y=1.305 $X2=3.945 $Y2=2.32
cc_91 VPB N_A_101_21#_c_176_n 0.0615756f $X=-0.19 $Y=1.305 $X2=2.045 $Y2=1.202
cc_92 VPB N_C_M1002_g 0.0314008f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=0.995
cc_93 VPB N_C_c_311_n 0.0408591f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=0.56
cc_94 VPB N_C_c_313_n 0.00696928f $X=-0.19 $Y=1.305 $X2=1.05 $Y2=0.56
cc_95 VPB N_C_c_314_n 0.0248178f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=1.985
cc_96 VPB N_A_532_93#_c_370_n 0.0345528f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=0.995
cc_97 VPB N_A_532_93#_c_372_n 0.00441836f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=1.985
cc_98 VPB N_A_532_93#_c_376_n 0.00959494f $X=-0.19 $Y=1.305 $X2=1.53 $Y2=0.56
cc_99 VPB N_A_532_93#_c_377_n 0.00173389f $X=-0.19 $Y=1.305 $X2=1.575 $Y2=1.985
cc_100 VPB N_A_532_93#_c_378_n 0.00184072f $X=-0.19 $Y=1.305 $X2=1.575 $Y2=1.985
cc_101 VPB N_A_532_93#_c_373_n 2.68423e-19 $X=-0.19 $Y=1.305 $X2=2.045 $Y2=1.41
cc_102 VPB N_A_1089_297#_c_456_n 0.0204513f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=0.995
cc_103 VPB N_A_1089_297#_c_444_n 0.0104627f $X=-0.19 $Y=1.305 $X2=1.05 $Y2=0.56
cc_104 VPB N_A_1089_297#_c_458_n 0.0241571f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=1.41
cc_105 VPB N_A_1089_297#_c_446_n 0.0104543f $X=-0.19 $Y=1.305 $X2=1.575 $Y2=1.41
cc_106 VPB N_A_1089_297#_c_447_n 0.00765838f $X=-0.19 $Y=1.305 $X2=1.575
+ $Y2=1.985
cc_107 VPB N_A_1089_297#_c_461_n 0.00601461f $X=-0.19 $Y=1.305 $X2=2 $Y2=0.56
cc_108 VPB N_A_1089_297#_c_455_n 0.00321756f $X=-0.19 $Y=1.305 $X2=1.05
+ $Y2=1.202
cc_109 VPB N_B_c_630_n 0.0216593f $X=-0.19 $Y=1.305 $X2=3.875 $Y2=0.245
cc_110 VPB N_B_c_624_n 0.00748587f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=0.56
cc_111 VPB N_B_M1008_g 0.0155244f $X=-0.19 $Y=1.305 $X2=1.05 $Y2=0.995
cc_112 VPB N_B_c_633_n 0.124505f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=1.985
cc_113 VPB N_B_c_634_n 0.0170126f $X=-0.19 $Y=1.305 $X2=1.53 $Y2=0.995
cc_114 VPB N_B_c_635_n 0.0101708f $X=-0.19 $Y=1.305 $X2=1.575 $Y2=1.985
cc_115 VPB N_B_c_636_n 0.00717497f $X=-0.19 $Y=1.305 $X2=2 $Y2=0.995
cc_116 VPB N_B_M1016_g 0.0130994f $X=-0.19 $Y=1.305 $X2=2.045 $Y2=1.41
cc_117 VPB N_B_c_626_n 0.00875008f $X=-0.19 $Y=1.305 $X2=2.175 $Y2=1.325
cc_118 VPB N_B_c_627_n 9.77983e-19 $X=-0.19 $Y=1.305 $X2=2.63 $Y2=1.96
cc_119 VPB N_B_c_628_n 0.0052573f $X=-0.19 $Y=1.305 $X2=2.285 $Y2=1.96
cc_120 VPB N_B_c_641_n 0.00204456f $X=-0.19 $Y=1.305 $X2=2.625 $Y2=0.695
cc_121 VPB B 0.00802749f $X=-0.19 $Y=1.305 $X2=2.74 $Y2=2.045
cc_122 VPB N_A_c_756_n 0.02697f $X=-0.19 $Y=1.305 $X2=3.875 $Y2=0.245
cc_123 VPB A 0.00142645f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=0.995
cc_124 VPB N_A_1207_297#_c_794_n 0.0291085f $X=-0.19 $Y=1.305 $X2=1.05 $Y2=0.995
cc_125 VPB N_A_1207_297#_c_803_n 0.00189028f $X=-0.19 $Y=1.305 $X2=1.575
+ $Y2=1.985
cc_126 VPB N_A_1207_297#_c_799_n 2.7046e-19 $X=-0.19 $Y=1.305 $X2=2.045
+ $Y2=1.985
cc_127 VPB N_A_1207_297#_c_805_n 0.00156472f $X=-0.19 $Y=1.305 $X2=2.045
+ $Y2=1.985
cc_128 VPB N_A_1207_297#_c_801_n 0.00274744f $X=-0.19 $Y=1.305 $X2=3.7 $Y2=0.34
cc_129 VPB N_VPWR_c_930_n 0.00470597f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=1.985
cc_130 VPB N_VPWR_c_931_n 0.00417454f $X=-0.19 $Y=1.305 $X2=1.575 $Y2=1.985
cc_131 VPB N_VPWR_c_932_n 0.0169755f $X=-0.19 $Y=1.305 $X2=2.045 $Y2=1.41
cc_132 VPB N_VPWR_c_933_n 0.00686977f $X=-0.19 $Y=1.305 $X2=2.175 $Y2=1.875
cc_133 VPB N_VPWR_c_934_n 0.00743637f $X=-0.19 $Y=1.305 $X2=2.285 $Y2=1.96
cc_134 VPB N_VPWR_c_935_n 0.0112126f $X=-0.19 $Y=1.305 $X2=2.74 $Y2=2.045
cc_135 VPB N_VPWR_c_936_n 0.00324402f $X=-0.19 $Y=1.305 $X2=2.74 $Y2=2.235
cc_136 VPB N_VPWR_c_937_n 0.0211506f $X=-0.19 $Y=1.305 $X2=3.7 $Y2=0.34
cc_137 VPB N_VPWR_c_938_n 0.00324069f $X=-0.19 $Y=1.305 $X2=2.735 $Y2=0.34
cc_138 VPB N_VPWR_c_939_n 0.0625838f $X=-0.19 $Y=1.305 $X2=3.945 $Y2=2.32
cc_139 VPB N_VPWR_c_940_n 0.00513206f $X=-0.19 $Y=1.305 $X2=3.945 $Y2=2.32
cc_140 VPB N_VPWR_c_941_n 0.0960788f $X=-0.19 $Y=1.305 $X2=1.575 $Y2=1.202
cc_141 VPB N_VPWR_c_942_n 0.0218344f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_929_n 0.0839116f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_944_n 0.00589444f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_945_n 0.00563188f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_X_c_1047_n 0.00131358f $X=-0.19 $Y=1.305 $X2=2.045 $Y2=1.985
cc_146 VPB N_A_657_325#_c_1095_n 0.0110171f $X=-0.19 $Y=1.305 $X2=1.05 $Y2=0.995
cc_147 VPB N_A_657_325#_c_1092_n 0.00805098f $X=-0.19 $Y=1.305 $X2=1.575
+ $Y2=1.985
cc_148 VPB N_A_657_325#_c_1097_n 0.00296592f $X=-0.19 $Y=1.305 $X2=2 $Y2=0.995
cc_149 VPB N_A_657_325#_c_1098_n 0.00293344f $X=-0.19 $Y=1.305 $X2=2.045
+ $Y2=1.41
cc_150 VPB N_A_657_325#_c_1099_n 0.0106403f $X=-0.19 $Y=1.305 $X2=2.045
+ $Y2=1.985
cc_151 VPB N_A_657_325#_c_1100_n 0.00172555f $X=-0.19 $Y=1.305 $X2=2.045
+ $Y2=1.985
cc_152 VPB N_A_657_325#_c_1093_n 0.00149669f $X=-0.19 $Y=1.305 $X2=2.175
+ $Y2=1.875
cc_153 VPB N_A_657_325#_c_1102_n 0.024643f $X=-0.19 $Y=1.305 $X2=2.63 $Y2=1.96
cc_154 VPB N_A_657_325#_c_1103_n 3.60787e-19 $X=-0.19 $Y=1.305 $X2=3.945
+ $Y2=2.32
cc_155 VPB N_A_657_325#_c_1104_n 3.41339e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_681_49#_c_1245_n 0.00148953f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=1.41
cc_157 VPB N_A_681_49#_c_1249_n 0.00271739f $X=-0.19 $Y=1.305 $X2=1.075
+ $Y2=1.985
cc_158 VPB N_A_681_49#_c_1250_n 8.62277e-19 $X=-0.19 $Y=1.305 $X2=1.53 $Y2=0.56
cc_159 VPB N_A_681_49#_c_1246_n 0.0021572f $X=-0.19 $Y=1.305 $X2=1.575 $Y2=1.985
cc_160 VPB N_A_681_49#_c_1252_n 0.0148602f $X=-0.19 $Y=1.305 $X2=2.285 $Y2=1.96
cc_161 VPB N_A_681_49#_c_1253_n 0.00333347f $X=-0.19 $Y=1.305 $X2=2.625
+ $Y2=0.425
cc_162 VPB N_A_681_49#_c_1254_n 0.008761f $X=-0.19 $Y=1.305 $X2=2.74 $Y2=2.235
cc_163 VPB N_A_681_49#_c_1255_n 0.00154407f $X=-0.19 $Y=1.305 $X2=2.85 $Y2=2.32
cc_164 VPB N_A_1490_297#_c_1380_n 0.00468751f $X=-0.19 $Y=1.305 $X2=1.05
+ $Y2=0.56
cc_165 VPB N_A_1490_297#_c_1384_n 0.0147295f $X=-0.19 $Y=1.305 $X2=1.575
+ $Y2=1.985
cc_166 VPB N_A_1490_297#_c_1381_n 0.0229927f $X=-0.19 $Y=1.305 $X2=2 $Y2=0.56
cc_167 VPB N_A_1490_297#_c_1386_n 0.0101148f $X=-0.19 $Y=1.305 $X2=2.175
+ $Y2=1.325
cc_168 N_A_101_21#_c_171_n N_C_c_310_n 0.0124123f $X=2 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_169 N_A_101_21#_c_172_n N_C_c_310_n 0.00141454f $X=2.175 $Y=1.325 $X2=-0.19
+ $Y2=-0.24
cc_170 N_A_101_21#_c_188_p N_C_c_310_n 0.0121806f $X=2.515 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_171 N_A_101_21#_c_173_n N_C_c_310_n 0.0106989f $X=2.625 $Y=0.695 $X2=-0.19
+ $Y2=-0.24
cc_172 N_A_101_21#_c_174_n N_C_c_310_n 0.00609706f $X=2.735 $Y=0.34 $X2=-0.19
+ $Y2=-0.24
cc_173 N_A_101_21#_c_180_n N_C_M1002_g 0.0216907f $X=2.045 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_101_21#_c_181_n N_C_M1002_g 0.00555142f $X=2.175 $Y=1.875 $X2=0 $Y2=0
cc_175 N_A_101_21#_c_193_p N_C_M1002_g 0.0132115f $X=2.63 $Y=1.96 $X2=0 $Y2=0
cc_176 N_A_101_21#_c_182_n N_C_M1002_g 0.00742917f $X=2.74 $Y=2.235 $X2=0 $Y2=0
cc_177 N_A_101_21#_c_183_n N_C_M1002_g 0.00743853f $X=2.85 $Y=2.32 $X2=0 $Y2=0
cc_178 N_A_101_21#_c_184_n N_C_c_311_n 0.0112964f $X=3.945 $Y=2.32 $X2=0 $Y2=0
cc_179 N_A_101_21#_c_197_p N_C_c_312_n 0.0106037f $X=3.9 $Y=0.355 $X2=0 $Y2=0
cc_180 N_A_101_21#_c_172_n N_C_c_313_n 0.0016003f $X=2.175 $Y=1.325 $X2=0 $Y2=0
cc_181 N_A_101_21#_c_181_n N_C_c_313_n 8.85809e-19 $X=2.175 $Y=1.875 $X2=0 $Y2=0
cc_182 N_A_101_21#_c_176_n N_C_c_313_n 0.0266772f $X=2.045 $Y=1.202 $X2=0 $Y2=0
cc_183 N_A_101_21#_c_175_n N_C_c_314_n 0.0111296f $X=3.7 $Y=0.355 $X2=0 $Y2=0
cc_184 N_A_101_21#_c_175_n N_C_c_335_n 0.00344638f $X=3.7 $Y=0.355 $X2=0 $Y2=0
cc_185 N_A_101_21#_c_188_p N_A_532_93#_M1026_d 0.00226086f $X=2.515 $Y=0.78
+ $X2=-0.19 $Y2=-0.24
cc_186 N_A_101_21#_c_173_n N_A_532_93#_M1026_d 0.00618081f $X=2.625 $Y=0.695
+ $X2=-0.19 $Y2=-0.24
cc_187 N_A_101_21#_c_193_p N_A_532_93#_M1002_d 0.00416203f $X=2.63 $Y=1.96 $X2=0
+ $Y2=0
cc_188 N_A_101_21#_c_182_n N_A_532_93#_M1002_d 0.00266846f $X=2.74 $Y=2.235
+ $X2=0 $Y2=0
cc_189 N_A_101_21#_c_184_n N_A_532_93#_c_370_n 0.0116412f $X=3.945 $Y=2.32 $X2=0
+ $Y2=0
cc_190 N_A_101_21#_c_208_p N_A_532_93#_c_371_n 0.00264322f $X=4.02 $Y=0.37 $X2=0
+ $Y2=0
cc_191 N_A_101_21#_c_188_p N_A_532_93#_c_386_n 0.00409956f $X=2.515 $Y=0.78
+ $X2=0 $Y2=0
cc_192 N_A_101_21#_c_193_p N_A_532_93#_c_386_n 0.0200253f $X=2.63 $Y=1.96 $X2=0
+ $Y2=0
cc_193 N_A_101_21#_c_184_n N_A_532_93#_c_386_n 0.00176797f $X=3.945 $Y=2.32
+ $X2=0 $Y2=0
cc_194 N_A_101_21#_c_172_n N_A_532_93#_c_372_n 0.0118646f $X=2.175 $Y=1.325
+ $X2=0 $Y2=0
cc_195 N_A_101_21#_c_181_n N_A_532_93#_c_372_n 0.00630296f $X=2.175 $Y=1.875
+ $X2=0 $Y2=0
cc_196 N_A_101_21#_c_188_p N_A_532_93#_c_372_n 0.0138225f $X=2.515 $Y=0.78 $X2=0
+ $Y2=0
cc_197 N_A_101_21#_c_173_n N_A_532_93#_c_372_n 0.00736858f $X=2.625 $Y=0.695
+ $X2=0 $Y2=0
cc_198 N_A_101_21#_c_175_n N_A_532_93#_c_372_n 0.0130244f $X=3.7 $Y=0.355 $X2=0
+ $Y2=0
cc_199 N_A_101_21#_c_176_n N_A_532_93#_c_372_n 7.41983e-19 $X=2.045 $Y=1.202
+ $X2=0 $Y2=0
cc_200 N_A_101_21#_M1019_d N_A_532_93#_c_376_n 0.00779963f $X=3.8 $Y=1.625 $X2=0
+ $Y2=0
cc_201 N_A_101_21#_c_184_n N_A_532_93#_c_376_n 0.0039224f $X=3.945 $Y=2.32 $X2=0
+ $Y2=0
cc_202 N_A_101_21#_M1019_d N_A_532_93#_c_377_n 5.89264e-19 $X=3.8 $Y=1.625 $X2=0
+ $Y2=0
cc_203 N_A_101_21#_c_184_n N_A_532_93#_c_378_n 0.00633062f $X=3.945 $Y=2.32
+ $X2=0 $Y2=0
cc_204 N_A_101_21#_c_181_n N_VPWR_M1024_s 0.00451219f $X=2.175 $Y=1.875 $X2=0
+ $Y2=0
cc_205 N_A_101_21#_c_193_p N_VPWR_M1024_s 0.00859265f $X=2.63 $Y=1.96 $X2=0
+ $Y2=0
cc_206 N_A_101_21#_c_224_p N_VPWR_M1024_s 9.86211e-19 $X=2.285 $Y=1.96 $X2=0
+ $Y2=0
cc_207 N_A_101_21#_c_177_n N_VPWR_c_930_n 0.00805332f $X=0.605 $Y=1.41 $X2=0
+ $Y2=0
cc_208 N_A_101_21#_c_178_n N_VPWR_c_931_n 0.00707507f $X=1.075 $Y=1.41 $X2=0
+ $Y2=0
cc_209 N_A_101_21#_c_179_n N_VPWR_c_931_n 0.00404416f $X=1.575 $Y=1.41 $X2=0
+ $Y2=0
cc_210 N_A_101_21#_c_176_n N_VPWR_c_931_n 0.00402805f $X=2.045 $Y=1.202 $X2=0
+ $Y2=0
cc_211 N_A_101_21#_c_179_n N_VPWR_c_932_n 0.00552168f $X=1.575 $Y=1.41 $X2=0
+ $Y2=0
cc_212 N_A_101_21#_c_180_n N_VPWR_c_932_n 0.00427505f $X=2.045 $Y=1.41 $X2=0
+ $Y2=0
cc_213 N_A_101_21#_c_179_n N_VPWR_c_933_n 5.19858e-19 $X=1.575 $Y=1.41 $X2=0
+ $Y2=0
cc_214 N_A_101_21#_c_180_n N_VPWR_c_933_n 0.0112695f $X=2.045 $Y=1.41 $X2=0
+ $Y2=0
cc_215 N_A_101_21#_c_193_p N_VPWR_c_933_n 0.0126548f $X=2.63 $Y=1.96 $X2=0 $Y2=0
cc_216 N_A_101_21#_c_224_p N_VPWR_c_933_n 0.0133756f $X=2.285 $Y=1.96 $X2=0
+ $Y2=0
cc_217 N_A_101_21#_c_182_n N_VPWR_c_933_n 0.00145799f $X=2.74 $Y=2.235 $X2=0
+ $Y2=0
cc_218 N_A_101_21#_c_183_n N_VPWR_c_933_n 0.0137789f $X=2.85 $Y=2.32 $X2=0 $Y2=0
cc_219 N_A_101_21#_c_177_n N_VPWR_c_937_n 0.00601503f $X=0.605 $Y=1.41 $X2=0
+ $Y2=0
cc_220 N_A_101_21#_c_178_n N_VPWR_c_937_n 0.00674661f $X=1.075 $Y=1.41 $X2=0
+ $Y2=0
cc_221 N_A_101_21#_c_193_p N_VPWR_c_939_n 0.00233941f $X=2.63 $Y=1.96 $X2=0
+ $Y2=0
cc_222 N_A_101_21#_c_183_n N_VPWR_c_939_n 0.0109705f $X=2.85 $Y=2.32 $X2=0 $Y2=0
cc_223 N_A_101_21#_c_184_n N_VPWR_c_939_n 0.0597844f $X=3.945 $Y=2.32 $X2=0
+ $Y2=0
cc_224 N_A_101_21#_c_177_n N_VPWR_c_929_n 0.011f $X=0.605 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A_101_21#_c_178_n N_VPWR_c_929_n 0.0119203f $X=1.075 $Y=1.41 $X2=0
+ $Y2=0
cc_226 N_A_101_21#_c_179_n N_VPWR_c_929_n 0.00903501f $X=1.575 $Y=1.41 $X2=0
+ $Y2=0
cc_227 N_A_101_21#_c_180_n N_VPWR_c_929_n 0.00732977f $X=2.045 $Y=1.41 $X2=0
+ $Y2=0
cc_228 N_A_101_21#_c_193_p N_VPWR_c_929_n 0.00553584f $X=2.63 $Y=1.96 $X2=0
+ $Y2=0
cc_229 N_A_101_21#_c_224_p N_VPWR_c_929_n 9.98534e-19 $X=2.285 $Y=1.96 $X2=0
+ $Y2=0
cc_230 N_A_101_21#_c_183_n N_VPWR_c_929_n 0.00809357f $X=2.85 $Y=2.32 $X2=0
+ $Y2=0
cc_231 N_A_101_21#_c_184_n N_VPWR_c_929_n 0.0473531f $X=3.945 $Y=2.32 $X2=0
+ $Y2=0
cc_232 N_A_101_21#_c_168_n N_X_c_1046_n 0.0181573f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_101_21#_c_169_n N_X_c_1046_n 0.00220043f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A_101_21#_c_177_n N_X_c_1051_n 0.0189644f $X=0.605 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A_101_21#_c_178_n N_X_c_1051_n 0.0135707f $X=1.075 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A_101_21#_c_179_n N_X_c_1051_n 4.9651e-19 $X=1.575 $Y=1.41 $X2=0 $Y2=0
cc_237 N_A_101_21#_c_176_n N_X_c_1051_n 0.00848497f $X=2.045 $Y=1.202 $X2=0
+ $Y2=0
cc_238 N_A_101_21#_c_176_n N_X_c_1055_n 0.0554438f $X=2.045 $Y=1.202 $X2=0 $Y2=0
cc_239 N_A_101_21#_c_170_n N_X_c_1056_n 0.00582185f $X=1.53 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A_101_21#_c_176_n N_X_c_1057_n 0.0407158f $X=2.045 $Y=1.202 $X2=0 $Y2=0
cc_241 N_A_101_21#_c_169_n N_X_c_1047_n 7.174e-19 $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_101_21#_c_178_n N_X_c_1047_n 2.91505e-19 $X=1.075 $Y=1.41 $X2=0 $Y2=0
cc_243 N_A_101_21#_c_170_n N_X_c_1047_n 0.00701394f $X=1.53 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_101_21#_c_179_n N_X_c_1047_n 0.00445754f $X=1.575 $Y=1.41 $X2=0 $Y2=0
cc_245 N_A_101_21#_c_171_n N_X_c_1047_n 0.00144676f $X=2 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_101_21#_c_180_n N_X_c_1047_n 9.53684e-19 $X=2.045 $Y=1.41 $X2=0 $Y2=0
cc_247 N_A_101_21#_c_172_n N_X_c_1047_n 0.0380181f $X=2.175 $Y=1.325 $X2=0 $Y2=0
cc_248 N_A_101_21#_c_181_n N_X_c_1047_n 0.0201514f $X=2.175 $Y=1.875 $X2=0 $Y2=0
cc_249 N_A_101_21#_c_176_n N_X_c_1047_n 0.0272364f $X=2.045 $Y=1.202 $X2=0 $Y2=0
cc_250 N_A_101_21#_c_179_n N_X_c_1067_n 0.014604f $X=1.575 $Y=1.41 $X2=0 $Y2=0
cc_251 N_A_101_21#_c_181_n N_X_c_1067_n 0.0202726f $X=2.175 $Y=1.875 $X2=0 $Y2=0
cc_252 N_A_101_21#_c_224_p N_X_c_1067_n 0.0140085f $X=2.285 $Y=1.96 $X2=0 $Y2=0
cc_253 N_A_101_21#_c_184_n N_A_657_325#_M1019_s 0.00736441f $X=3.945 $Y=2.32
+ $X2=0 $Y2=0
cc_254 N_A_101_21#_M1019_d N_A_657_325#_c_1095_n 0.00509381f $X=3.8 $Y=1.625
+ $X2=0 $Y2=0
cc_255 N_A_101_21#_c_193_p N_A_657_325#_c_1095_n 0.00831987f $X=2.63 $Y=1.96
+ $X2=0 $Y2=0
cc_256 N_A_101_21#_c_182_n N_A_657_325#_c_1095_n 9.56599e-19 $X=2.74 $Y=2.235
+ $X2=0 $Y2=0
cc_257 N_A_101_21#_c_184_n N_A_657_325#_c_1095_n 0.0571361f $X=3.945 $Y=2.32
+ $X2=0 $Y2=0
cc_258 N_A_101_21#_c_208_p N_A_657_325#_c_1090_n 0.0126757f $X=4.02 $Y=0.37
+ $X2=0 $Y2=0
cc_259 N_A_101_21#_c_175_n N_A_681_49#_M1023_s 0.00652268f $X=3.7 $Y=0.355
+ $X2=-0.19 $Y2=-0.24
cc_260 N_A_101_21#_M1023_d N_A_681_49#_c_1257_n 0.00837215f $X=3.875 $Y=0.245
+ $X2=0 $Y2=0
cc_261 N_A_101_21#_c_208_p N_A_681_49#_c_1257_n 0.0136844f $X=4.02 $Y=0.37 $X2=0
+ $Y2=0
cc_262 N_A_101_21#_c_197_p N_A_681_49#_c_1247_n 0.0136844f $X=3.9 $Y=0.355 $X2=0
+ $Y2=0
cc_263 N_A_101_21#_c_175_n N_A_681_49#_c_1247_n 0.0181831f $X=3.7 $Y=0.355 $X2=0
+ $Y2=0
cc_264 N_A_101_21#_c_172_n N_VGND_M1017_d 0.00214092f $X=2.175 $Y=1.325 $X2=0
+ $Y2=0
cc_265 N_A_101_21#_c_188_p N_VGND_M1017_d 0.00889686f $X=2.515 $Y=0.78 $X2=0
+ $Y2=0
cc_266 N_A_101_21#_c_168_n N_VGND_c_1446_n 0.00687701f $X=0.58 $Y=0.995 $X2=0
+ $Y2=0
cc_267 N_A_101_21#_c_169_n N_VGND_c_1447_n 0.00717939f $X=1.05 $Y=0.995 $X2=0
+ $Y2=0
cc_268 N_A_101_21#_c_170_n N_VGND_c_1447_n 0.00413278f $X=1.53 $Y=0.995 $X2=0
+ $Y2=0
cc_269 N_A_101_21#_c_176_n N_VGND_c_1447_n 0.00308104f $X=2.045 $Y=1.202 $X2=0
+ $Y2=0
cc_270 N_A_101_21#_c_170_n N_VGND_c_1448_n 0.00531141f $X=1.53 $Y=0.995 $X2=0
+ $Y2=0
cc_271 N_A_101_21#_c_171_n N_VGND_c_1448_n 0.0046653f $X=2 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A_101_21#_c_170_n N_VGND_c_1449_n 8.64053e-19 $X=1.53 $Y=0.995 $X2=0
+ $Y2=0
cc_273 N_A_101_21#_c_171_n N_VGND_c_1449_n 0.00969109f $X=2 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A_101_21#_c_172_n N_VGND_c_1449_n 0.0147747f $X=2.175 $Y=1.325 $X2=0
+ $Y2=0
cc_275 N_A_101_21#_c_188_p N_VGND_c_1449_n 0.0045481f $X=2.515 $Y=0.78 $X2=0
+ $Y2=0
cc_276 N_A_101_21#_c_173_n N_VGND_c_1449_n 0.00744451f $X=2.625 $Y=0.695 $X2=0
+ $Y2=0
cc_277 N_A_101_21#_c_174_n N_VGND_c_1449_n 0.0142743f $X=2.735 $Y=0.34 $X2=0
+ $Y2=0
cc_278 N_A_101_21#_c_176_n N_VGND_c_1449_n 7.5828e-19 $X=2.045 $Y=1.202 $X2=0
+ $Y2=0
cc_279 N_A_101_21#_c_168_n N_VGND_c_1454_n 0.00545968f $X=0.58 $Y=0.995 $X2=0
+ $Y2=0
cc_280 N_A_101_21#_c_169_n N_VGND_c_1454_n 0.00585385f $X=1.05 $Y=0.995 $X2=0
+ $Y2=0
cc_281 N_A_101_21#_c_188_p N_VGND_c_1458_n 0.00219715f $X=2.515 $Y=0.78 $X2=0
+ $Y2=0
cc_282 N_A_101_21#_c_174_n N_VGND_c_1458_n 0.0156439f $X=2.735 $Y=0.34 $X2=0
+ $Y2=0
cc_283 N_A_101_21#_c_175_n N_VGND_c_1458_n 0.0893431f $X=3.7 $Y=0.355 $X2=0
+ $Y2=0
cc_284 N_A_101_21#_c_168_n N_VGND_c_1460_n 0.0108498f $X=0.58 $Y=0.995 $X2=0
+ $Y2=0
cc_285 N_A_101_21#_c_169_n N_VGND_c_1460_n 0.0111002f $X=1.05 $Y=0.995 $X2=0
+ $Y2=0
cc_286 N_A_101_21#_c_170_n N_VGND_c_1460_n 0.00957564f $X=1.53 $Y=0.995 $X2=0
+ $Y2=0
cc_287 N_A_101_21#_c_171_n N_VGND_c_1460_n 0.00809951f $X=2 $Y=0.995 $X2=0 $Y2=0
cc_288 N_A_101_21#_c_172_n N_VGND_c_1460_n 0.00101551f $X=2.175 $Y=1.325 $X2=0
+ $Y2=0
cc_289 N_A_101_21#_c_188_p N_VGND_c_1460_n 0.00486078f $X=2.515 $Y=0.78 $X2=0
+ $Y2=0
cc_290 N_A_101_21#_c_174_n N_VGND_c_1460_n 0.00844855f $X=2.735 $Y=0.34 $X2=0
+ $Y2=0
cc_291 N_A_101_21#_c_175_n N_VGND_c_1460_n 0.0533662f $X=3.7 $Y=0.355 $X2=0
+ $Y2=0
cc_292 N_C_c_311_n N_A_532_93#_c_370_n 0.0592216f $X=3.71 $Y=1.55 $X2=0 $Y2=0
cc_293 N_C_c_335_n N_A_532_93#_c_370_n 2.68329e-19 $X=3.545 $Y=1.16 $X2=0 $Y2=0
cc_294 N_C_c_312_n N_A_532_93#_c_371_n 0.0232388f $X=3.8 $Y=0.995 $X2=0 $Y2=0
cc_295 N_C_M1002_g N_A_532_93#_c_386_n 0.011319f $X=2.61 $Y=1.805 $X2=0 $Y2=0
cc_296 N_C_c_314_n N_A_532_93#_c_386_n 0.00634718f $X=3.61 $Y=1.16 $X2=0 $Y2=0
cc_297 N_C_c_310_n N_A_532_93#_c_372_n 0.00436363f $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_298 N_C_M1002_g N_A_532_93#_c_372_n 0.00203559f $X=2.61 $Y=1.805 $X2=0 $Y2=0
cc_299 N_C_c_311_n N_A_532_93#_c_372_n 0.00508695f $X=3.71 $Y=1.55 $X2=0 $Y2=0
cc_300 N_C_c_312_n N_A_532_93#_c_372_n 0.00235914f $X=3.8 $Y=0.995 $X2=0 $Y2=0
cc_301 N_C_c_313_n N_A_532_93#_c_372_n 0.0020376f $X=2.61 $Y=1.202 $X2=0 $Y2=0
cc_302 N_C_c_314_n N_A_532_93#_c_372_n 0.0266322f $X=3.61 $Y=1.16 $X2=0 $Y2=0
cc_303 N_C_c_335_n N_A_532_93#_c_372_n 0.018733f $X=3.545 $Y=1.16 $X2=0 $Y2=0
cc_304 N_C_c_311_n N_A_532_93#_c_376_n 0.017213f $X=3.71 $Y=1.55 $X2=0 $Y2=0
cc_305 N_C_c_314_n N_A_532_93#_c_376_n 0.0140512f $X=3.61 $Y=1.16 $X2=0 $Y2=0
cc_306 N_C_c_335_n N_A_532_93#_c_376_n 0.0378363f $X=3.545 $Y=1.16 $X2=0 $Y2=0
cc_307 N_C_c_311_n N_A_532_93#_c_377_n 0.00427971f $X=3.71 $Y=1.55 $X2=0 $Y2=0
cc_308 N_C_c_311_n N_A_532_93#_c_373_n 0.00353238f $X=3.71 $Y=1.55 $X2=0 $Y2=0
cc_309 N_C_c_335_n N_A_532_93#_c_373_n 0.0207305f $X=3.545 $Y=1.16 $X2=0 $Y2=0
cc_310 N_C_M1002_g N_VPWR_c_933_n 0.00202848f $X=2.61 $Y=1.805 $X2=0 $Y2=0
cc_311 N_C_M1002_g N_VPWR_c_939_n 0.00514356f $X=2.61 $Y=1.805 $X2=0 $Y2=0
cc_312 N_C_c_311_n N_VPWR_c_939_n 0.00427564f $X=3.71 $Y=1.55 $X2=0 $Y2=0
cc_313 N_C_M1002_g N_VPWR_c_929_n 0.00682402f $X=2.61 $Y=1.805 $X2=0 $Y2=0
cc_314 N_C_c_311_n N_VPWR_c_929_n 0.00784458f $X=3.71 $Y=1.55 $X2=0 $Y2=0
cc_315 N_C_M1002_g N_A_657_325#_c_1095_n 9.4239e-19 $X=2.61 $Y=1.805 $X2=0 $Y2=0
cc_316 N_C_c_311_n N_A_657_325#_c_1095_n 0.0102234f $X=3.71 $Y=1.55 $X2=0 $Y2=0
cc_317 N_C_c_312_n N_A_681_49#_c_1257_n 0.00846885f $X=3.8 $Y=0.995 $X2=0 $Y2=0
cc_318 N_C_c_335_n N_A_681_49#_c_1257_n 0.00489958f $X=3.545 $Y=1.16 $X2=0 $Y2=0
cc_319 N_C_c_312_n N_A_681_49#_c_1247_n 0.00389299f $X=3.8 $Y=0.995 $X2=0 $Y2=0
cc_320 N_C_c_314_n N_A_681_49#_c_1247_n 0.00656019f $X=3.61 $Y=1.16 $X2=0 $Y2=0
cc_321 N_C_c_335_n N_A_681_49#_c_1247_n 0.028934f $X=3.545 $Y=1.16 $X2=0 $Y2=0
cc_322 N_C_c_310_n N_VGND_c_1449_n 0.00141765f $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_323 N_C_c_310_n N_VGND_c_1458_n 8.79444e-19 $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_324 N_C_c_312_n N_VGND_c_1458_n 0.00357877f $X=3.8 $Y=0.995 $X2=0 $Y2=0
cc_325 N_C_c_312_n N_VGND_c_1460_n 0.00692546f $X=3.8 $Y=0.995 $X2=0 $Y2=0
cc_326 N_A_532_93#_c_370_n N_VPWR_c_934_n 0.00632978f $X=4.245 $Y=1.41 $X2=0
+ $Y2=0
cc_327 N_A_532_93#_c_370_n N_VPWR_c_939_n 0.00412251f $X=4.245 $Y=1.41 $X2=0
+ $Y2=0
cc_328 N_A_532_93#_c_370_n N_VPWR_c_929_n 0.00595559f $X=4.245 $Y=1.41 $X2=0
+ $Y2=0
cc_329 N_A_532_93#_c_376_n N_A_657_325#_M1019_s 0.00373918f $X=4.03 $Y=1.62
+ $X2=0 $Y2=0
cc_330 N_A_532_93#_c_370_n N_A_657_325#_c_1095_n 0.0184006f $X=4.245 $Y=1.41
+ $X2=0 $Y2=0
cc_331 N_A_532_93#_c_376_n N_A_657_325#_c_1095_n 0.0556467f $X=4.03 $Y=1.62
+ $X2=0 $Y2=0
cc_332 N_A_532_93#_c_373_n N_A_657_325#_c_1095_n 0.00386917f $X=4.22 $Y=1.16
+ $X2=0 $Y2=0
cc_333 N_A_532_93#_c_371_n N_A_657_325#_c_1091_n 0.00387381f $X=4.33 $Y=0.995
+ $X2=0 $Y2=0
cc_334 N_A_532_93#_c_370_n N_A_657_325#_c_1092_n 0.00449957f $X=4.245 $Y=1.41
+ $X2=0 $Y2=0
cc_335 N_A_532_93#_c_370_n N_A_681_49#_c_1257_n 0.00399242f $X=4.245 $Y=1.41
+ $X2=0 $Y2=0
cc_336 N_A_532_93#_c_371_n N_A_681_49#_c_1257_n 0.0151871f $X=4.33 $Y=0.995
+ $X2=0 $Y2=0
cc_337 N_A_532_93#_c_373_n N_A_681_49#_c_1257_n 0.0193226f $X=4.22 $Y=1.16 $X2=0
+ $Y2=0
cc_338 N_A_532_93#_c_370_n N_A_681_49#_c_1245_n 0.00108145f $X=4.245 $Y=1.41
+ $X2=0 $Y2=0
cc_339 N_A_532_93#_c_371_n N_A_681_49#_c_1245_n 0.0150189f $X=4.33 $Y=0.995
+ $X2=0 $Y2=0
cc_340 N_A_532_93#_c_377_n N_A_681_49#_c_1245_n 0.00218396f $X=4.115 $Y=1.535
+ $X2=0 $Y2=0
cc_341 N_A_532_93#_c_373_n N_A_681_49#_c_1245_n 0.0247426f $X=4.22 $Y=1.16 $X2=0
+ $Y2=0
cc_342 N_A_532_93#_c_371_n N_A_681_49#_c_1247_n 5.11968e-19 $X=4.33 $Y=0.995
+ $X2=0 $Y2=0
cc_343 N_A_532_93#_c_372_n N_A_681_49#_c_1247_n 0.0151384f $X=2.99 $Y=0.76 $X2=0
+ $Y2=0
cc_344 N_A_532_93#_c_376_n N_A_681_49#_c_1253_n 5.94479e-19 $X=4.03 $Y=1.62
+ $X2=0 $Y2=0
cc_345 N_A_532_93#_c_377_n N_A_681_49#_c_1253_n 6.54862e-19 $X=4.115 $Y=1.535
+ $X2=0 $Y2=0
cc_346 N_A_532_93#_c_370_n N_A_681_49#_c_1254_n 0.00719438f $X=4.245 $Y=1.41
+ $X2=0 $Y2=0
cc_347 N_A_532_93#_c_376_n N_A_681_49#_c_1254_n 0.0102953f $X=4.03 $Y=1.62 $X2=0
+ $Y2=0
cc_348 N_A_532_93#_c_377_n N_A_681_49#_c_1254_n 0.00669828f $X=4.115 $Y=1.535
+ $X2=0 $Y2=0
cc_349 N_A_532_93#_c_371_n N_VGND_c_1458_n 0.0042361f $X=4.33 $Y=0.995 $X2=0
+ $Y2=0
cc_350 N_A_532_93#_c_371_n N_VGND_c_1460_n 0.0075143f $X=4.33 $Y=0.995 $X2=0
+ $Y2=0
cc_351 N_A_1089_297#_c_461_n N_B_c_630_n 0.00852064f $X=5.75 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_352 N_A_1089_297#_c_455_n N_B_c_630_n 8.18494e-19 $X=5.81 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_353 N_A_1089_297#_c_465_p N_B_M1004_g 0.00383107f $X=5.835 $Y=0.85 $X2=0
+ $Y2=0
cc_354 N_A_1089_297#_c_455_n N_B_M1004_g 0.0151084f $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_355 N_A_1089_297#_c_449_n N_B_c_623_n 0.0050801f $X=7.025 $Y=0.85 $X2=0 $Y2=0
cc_356 N_A_1089_297#_c_455_n N_B_c_623_n 0.0150884f $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_357 N_A_1089_297#_c_461_n N_B_c_624_n 0.00784394f $X=5.75 $Y=1.58 $X2=0 $Y2=0
cc_358 N_A_1089_297#_c_455_n N_B_c_624_n 0.00791542f $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_359 N_A_1089_297#_c_456_n N_B_M1008_g 0.0119272f $X=7.36 $Y=1.41 $X2=0 $Y2=0
cc_360 N_A_1089_297#_M1011_g N_B_M1006_g 0.0104686f $X=7.385 $Y=0.455 $X2=0
+ $Y2=0
cc_361 N_A_1089_297#_c_446_n N_B_M1006_g 0.021209f $X=7.26 $Y=1.16 $X2=0 $Y2=0
cc_362 N_A_1089_297#_c_448_n N_B_M1006_g 0.00188578f $X=7.15 $Y=0.995 $X2=0
+ $Y2=0
cc_363 N_A_1089_297#_c_449_n N_B_M1006_g 0.00221468f $X=7.025 $Y=0.85 $X2=0
+ $Y2=0
cc_364 N_A_1089_297#_c_451_n N_B_M1006_g 6.75018e-19 $X=7.315 $Y=0.85 $X2=0
+ $Y2=0
cc_365 N_A_1089_297#_c_452_n N_B_M1006_g 0.00140598f $X=7.17 $Y=0.85 $X2=0 $Y2=0
cc_366 N_A_1089_297#_c_456_n N_B_c_633_n 0.0105804f $X=7.36 $Y=1.41 $X2=0 $Y2=0
cc_367 N_A_1089_297#_c_458_n N_B_c_633_n 0.00616735f $X=8.85 $Y=1.57 $X2=0 $Y2=0
cc_368 N_A_1089_297#_c_444_n N_B_c_635_n 0.00407979f $X=8.85 $Y=1.47 $X2=0 $Y2=0
cc_369 N_A_1089_297#_c_458_n N_B_c_636_n 0.00407979f $X=8.85 $Y=1.57 $X2=0 $Y2=0
cc_370 N_A_1089_297#_c_458_n N_B_M1016_g 0.0249809f $X=8.85 $Y=1.57 $X2=0 $Y2=0
cc_371 N_A_1089_297#_c_447_n N_B_c_626_n 0.00181049f $X=7.36 $Y=1.202 $X2=0
+ $Y2=0
cc_372 N_A_1089_297#_c_443_n N_B_c_627_n 0.001267f $X=8.85 $Y=1.28 $X2=0 $Y2=0
cc_373 N_A_1089_297#_c_450_n N_B_c_627_n 0.00731236f $X=8.505 $Y=0.85 $X2=0
+ $Y2=0
cc_374 N_A_1089_297#_c_454_n N_B_c_627_n 0.021521f $X=8.65 $Y=0.85 $X2=0 $Y2=0
cc_375 N_A_1089_297#_c_443_n N_B_c_628_n 0.0192205f $X=8.85 $Y=1.28 $X2=0 $Y2=0
cc_376 N_A_1089_297#_c_447_n N_B_c_628_n 0.00774709f $X=7.36 $Y=1.202 $X2=0
+ $Y2=0
cc_377 N_A_1089_297#_c_450_n N_B_c_628_n 0.00133312f $X=8.505 $Y=0.85 $X2=0
+ $Y2=0
cc_378 N_A_1089_297#_c_454_n N_B_c_628_n 0.00172718f $X=8.65 $Y=0.85 $X2=0 $Y2=0
cc_379 N_A_1089_297#_c_443_n B 8.1069e-19 $X=8.85 $Y=1.28 $X2=0 $Y2=0
cc_380 N_A_1089_297#_c_444_n B 0.00133275f $X=8.85 $Y=1.47 $X2=0 $Y2=0
cc_381 N_A_1089_297#_c_458_n B 0.00483815f $X=8.85 $Y=1.57 $X2=0 $Y2=0
cc_382 N_A_1089_297#_c_450_n B 0.00414594f $X=8.505 $Y=0.85 $X2=0 $Y2=0
cc_383 N_A_1089_297#_c_453_n B 0.00235209f $X=8.65 $Y=0.85 $X2=0 $Y2=0
cc_384 N_A_1089_297#_c_454_n B 0.0183366f $X=8.65 $Y=0.85 $X2=0 $Y2=0
cc_385 N_A_1089_297#_M1011_g N_B_c_629_n 0.00774709f $X=7.385 $Y=0.455 $X2=0
+ $Y2=0
cc_386 N_A_1089_297#_c_443_n N_B_c_629_n 0.00135777f $X=8.85 $Y=1.28 $X2=0 $Y2=0
cc_387 N_A_1089_297#_c_445_n N_B_c_629_n 0.0134808f $X=8.88 $Y=0.945 $X2=0 $Y2=0
cc_388 N_A_1089_297#_c_450_n N_B_c_629_n 0.00740121f $X=8.505 $Y=0.85 $X2=0
+ $Y2=0
cc_389 N_A_1089_297#_c_453_n N_B_c_629_n 0.0014125f $X=8.65 $Y=0.85 $X2=0 $Y2=0
cc_390 N_A_1089_297#_c_454_n N_B_c_629_n 0.00207369f $X=8.65 $Y=0.85 $X2=0 $Y2=0
cc_391 N_A_1089_297#_c_443_n N_A_c_756_n 0.0181958f $X=8.85 $Y=1.28 $X2=-0.19
+ $Y2=-0.24
cc_392 N_A_1089_297#_c_444_n N_A_c_756_n 0.0102542f $X=8.85 $Y=1.47 $X2=-0.19
+ $Y2=-0.24
cc_393 N_A_1089_297#_c_458_n N_A_c_756_n 0.0315533f $X=8.85 $Y=1.57 $X2=-0.19
+ $Y2=-0.24
cc_394 N_A_1089_297#_c_454_n N_A_c_756_n 6.45074e-19 $X=8.65 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_395 N_A_1089_297#_c_445_n N_A_c_757_n 0.0188577f $X=8.88 $Y=0.945 $X2=0 $Y2=0
cc_396 N_A_1089_297#_c_454_n N_A_c_757_n 2.38541e-19 $X=8.65 $Y=0.85 $X2=0 $Y2=0
cc_397 N_A_1089_297#_c_443_n A 0.0015686f $X=8.85 $Y=1.28 $X2=0 $Y2=0
cc_398 N_A_1089_297#_c_444_n A 0.00114147f $X=8.85 $Y=1.47 $X2=0 $Y2=0
cc_399 N_A_1089_297#_c_454_n A 0.0133858f $X=8.65 $Y=0.85 $X2=0 $Y2=0
cc_400 N_A_1089_297#_c_449_n N_A_1207_297#_M1006_s 8.89732e-19 $X=7.025 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_401 N_A_1089_297#_c_455_n N_A_1207_297#_c_796_n 0.00447674f $X=5.81 $Y=0.74
+ $X2=0 $Y2=0
cc_402 N_A_1089_297#_c_449_n N_A_1207_297#_c_809_n 0.001069f $X=7.025 $Y=0.85
+ $X2=0 $Y2=0
cc_403 N_A_1089_297#_c_458_n N_A_1207_297#_c_803_n 0.00416703f $X=8.85 $Y=1.57
+ $X2=0 $Y2=0
cc_404 N_A_1089_297#_c_445_n N_A_1207_297#_c_798_n 0.00187335f $X=8.88 $Y=0.945
+ $X2=0 $Y2=0
cc_405 N_A_1089_297#_c_453_n N_A_1207_297#_c_798_n 0.00537182f $X=8.65 $Y=0.85
+ $X2=0 $Y2=0
cc_406 N_A_1089_297#_c_454_n N_A_1207_297#_c_798_n 0.00520032f $X=8.65 $Y=0.85
+ $X2=0 $Y2=0
cc_407 N_A_1089_297#_M1011_g N_A_1207_297#_c_814_n 0.00613906f $X=7.385 $Y=0.455
+ $X2=0 $Y2=0
cc_408 N_A_1089_297#_c_445_n N_A_1207_297#_c_814_n 0.0087978f $X=8.88 $Y=0.945
+ $X2=0 $Y2=0
cc_409 N_A_1089_297#_c_448_n N_A_1207_297#_c_814_n 3.69046e-19 $X=7.15 $Y=0.995
+ $X2=0 $Y2=0
cc_410 N_A_1089_297#_c_449_n N_A_1207_297#_c_814_n 0.0554529f $X=7.025 $Y=0.85
+ $X2=0 $Y2=0
cc_411 N_A_1089_297#_c_450_n N_A_1207_297#_c_814_n 0.0955498f $X=8.505 $Y=0.85
+ $X2=0 $Y2=0
cc_412 N_A_1089_297#_c_451_n N_A_1207_297#_c_814_n 0.026662f $X=7.315 $Y=0.85
+ $X2=0 $Y2=0
cc_413 N_A_1089_297#_c_452_n N_A_1207_297#_c_814_n 0.00310602f $X=7.17 $Y=0.85
+ $X2=0 $Y2=0
cc_414 N_A_1089_297#_c_453_n N_A_1207_297#_c_814_n 0.0266136f $X=8.65 $Y=0.85
+ $X2=0 $Y2=0
cc_415 N_A_1089_297#_c_454_n N_A_1207_297#_c_814_n 0.00475288f $X=8.65 $Y=0.85
+ $X2=0 $Y2=0
cc_416 N_A_1089_297#_c_449_n N_A_1207_297#_c_800_n 0.0271297f $X=7.025 $Y=0.85
+ $X2=0 $Y2=0
cc_417 N_A_1089_297#_c_455_n N_A_1207_297#_c_800_n 0.00716303f $X=5.81 $Y=0.74
+ $X2=0 $Y2=0
cc_418 N_A_1089_297#_c_461_n N_A_1207_297#_c_801_n 0.0194501f $X=5.75 $Y=1.58
+ $X2=0 $Y2=0
cc_419 N_A_1089_297#_c_449_n N_A_1207_297#_c_801_n 0.0123942f $X=7.025 $Y=0.85
+ $X2=0 $Y2=0
cc_420 N_A_1089_297#_c_465_p N_A_1207_297#_c_801_n 5.77119e-19 $X=5.835 $Y=0.85
+ $X2=0 $Y2=0
cc_421 N_A_1089_297#_c_455_n N_A_1207_297#_c_801_n 0.0672745f $X=5.81 $Y=0.74
+ $X2=0 $Y2=0
cc_422 N_A_1089_297#_c_445_n N_A_1207_297#_c_829_n 0.00156626f $X=8.88 $Y=0.945
+ $X2=0 $Y2=0
cc_423 N_A_1089_297#_c_445_n N_A_1207_297#_c_830_n 0.00809859f $X=8.88 $Y=0.945
+ $X2=0 $Y2=0
cc_424 N_A_1089_297#_c_458_n N_VPWR_c_941_n 0.00434439f $X=8.85 $Y=1.57 $X2=0
+ $Y2=0
cc_425 N_A_1089_297#_M1027_d N_VPWR_c_929_n 0.00367747f $X=5.445 $Y=1.485 $X2=0
+ $Y2=0
cc_426 N_A_1089_297#_c_458_n N_VPWR_c_929_n 0.00650675f $X=8.85 $Y=1.57 $X2=0
+ $Y2=0
cc_427 N_A_1089_297#_c_458_n N_VPWR_c_945_n 0.00129998f $X=8.85 $Y=1.57 $X2=0
+ $Y2=0
cc_428 N_A_1089_297#_c_449_n N_A_657_325#_M1006_d 0.00134889f $X=7.025 $Y=0.85
+ $X2=0 $Y2=0
cc_429 N_A_1089_297#_c_451_n N_A_657_325#_M1006_d 5.4759e-19 $X=7.315 $Y=0.85
+ $X2=0 $Y2=0
cc_430 N_A_1089_297#_c_452_n N_A_657_325#_M1006_d 0.00657455f $X=7.17 $Y=0.85
+ $X2=0 $Y2=0
cc_431 N_A_1089_297#_c_465_p N_A_657_325#_c_1091_n 0.0023462f $X=5.835 $Y=0.85
+ $X2=0 $Y2=0
cc_432 N_A_1089_297#_c_455_n N_A_657_325#_c_1091_n 0.00358462f $X=5.81 $Y=0.74
+ $X2=0 $Y2=0
cc_433 N_A_1089_297#_c_461_n N_A_657_325#_c_1092_n 0.0144171f $X=5.75 $Y=1.58
+ $X2=0 $Y2=0
cc_434 N_A_1089_297#_c_455_n N_A_657_325#_c_1092_n 0.00928178f $X=5.81 $Y=0.74
+ $X2=0 $Y2=0
cc_435 N_A_1089_297#_M1027_d N_A_657_325#_c_1097_n 0.00767171f $X=5.445 $Y=1.485
+ $X2=0 $Y2=0
cc_436 N_A_1089_297#_c_461_n N_A_657_325#_c_1097_n 0.0315546f $X=5.75 $Y=1.58
+ $X2=0 $Y2=0
cc_437 N_A_1089_297#_M1027_d N_A_657_325#_c_1098_n 0.00313827f $X=5.445 $Y=1.485
+ $X2=0 $Y2=0
cc_438 N_A_1089_297#_M1027_d N_A_657_325#_c_1100_n 0.00318432f $X=5.445 $Y=1.485
+ $X2=0 $Y2=0
cc_439 N_A_1089_297#_c_456_n N_A_657_325#_c_1093_n 0.00131578f $X=7.36 $Y=1.41
+ $X2=0 $Y2=0
cc_440 N_A_1089_297#_c_446_n N_A_657_325#_c_1093_n 6.52616e-19 $X=7.26 $Y=1.16
+ $X2=0 $Y2=0
cc_441 N_A_1089_297#_c_447_n N_A_657_325#_c_1093_n 3.9697e-19 $X=7.36 $Y=1.202
+ $X2=0 $Y2=0
cc_442 N_A_1089_297#_c_448_n N_A_657_325#_c_1093_n 0.0160828f $X=7.15 $Y=0.995
+ $X2=0 $Y2=0
cc_443 N_A_1089_297#_c_449_n N_A_657_325#_c_1093_n 0.0093317f $X=7.025 $Y=0.85
+ $X2=0 $Y2=0
cc_444 N_A_1089_297#_c_451_n N_A_657_325#_c_1093_n 0.00105141f $X=7.315 $Y=0.85
+ $X2=0 $Y2=0
cc_445 N_A_1089_297#_c_452_n N_A_657_325#_c_1093_n 0.0039699f $X=7.17 $Y=0.85
+ $X2=0 $Y2=0
cc_446 N_A_1089_297#_c_456_n N_A_657_325#_c_1102_n 0.00258134f $X=7.36 $Y=1.41
+ $X2=0 $Y2=0
cc_447 N_A_1089_297#_c_458_n N_A_657_325#_c_1102_n 0.00822576f $X=8.85 $Y=1.57
+ $X2=0 $Y2=0
cc_448 N_A_1089_297#_M1011_g N_A_657_325#_c_1139_n 0.00223265f $X=7.385 $Y=0.455
+ $X2=0 $Y2=0
cc_449 N_A_1089_297#_c_452_n N_A_657_325#_c_1139_n 0.00184505f $X=7.17 $Y=0.85
+ $X2=0 $Y2=0
cc_450 N_A_1089_297#_c_455_n N_A_657_325#_c_1094_n 0.00616264f $X=5.81 $Y=0.74
+ $X2=0 $Y2=0
cc_451 N_A_1089_297#_c_446_n N_A_657_325#_c_1142_n 2.19531e-19 $X=7.26 $Y=1.16
+ $X2=0 $Y2=0
cc_452 N_A_1089_297#_c_448_n N_A_657_325#_c_1142_n 0.00294425f $X=7.15 $Y=0.995
+ $X2=0 $Y2=0
cc_453 N_A_1089_297#_c_449_n N_A_657_325#_c_1142_n 0.0126621f $X=7.025 $Y=0.85
+ $X2=0 $Y2=0
cc_454 N_A_1089_297#_c_451_n N_A_657_325#_c_1142_n 0.00134696f $X=7.315 $Y=0.85
+ $X2=0 $Y2=0
cc_455 N_A_1089_297#_c_452_n N_A_657_325#_c_1142_n 0.0125043f $X=7.17 $Y=0.85
+ $X2=0 $Y2=0
cc_456 N_A_1089_297#_c_450_n N_A_681_49#_M1014_d 0.00140408f $X=8.505 $Y=0.85
+ $X2=0 $Y2=0
cc_457 N_A_1089_297#_c_453_n N_A_681_49#_M1014_d 0.00214439f $X=8.65 $Y=0.85
+ $X2=0 $Y2=0
cc_458 N_A_1089_297#_c_454_n N_A_681_49#_M1014_d 0.00513165f $X=8.65 $Y=0.85
+ $X2=0 $Y2=0
cc_459 N_A_1089_297#_c_446_n N_A_681_49#_c_1249_n 0.00881942f $X=7.26 $Y=1.16
+ $X2=0 $Y2=0
cc_460 N_A_1089_297#_c_448_n N_A_681_49#_c_1249_n 0.0271004f $X=7.15 $Y=0.995
+ $X2=0 $Y2=0
cc_461 N_A_1089_297#_c_449_n N_A_681_49#_c_1249_n 5.63776e-19 $X=7.025 $Y=0.85
+ $X2=0 $Y2=0
cc_462 N_A_1089_297#_c_456_n N_A_681_49#_c_1286_n 0.00383389f $X=7.36 $Y=1.41
+ $X2=0 $Y2=0
cc_463 N_A_1089_297#_c_456_n N_A_681_49#_c_1250_n 0.0175777f $X=7.36 $Y=1.41
+ $X2=0 $Y2=0
cc_464 N_A_1089_297#_c_446_n N_A_681_49#_c_1250_n 7.42472e-19 $X=7.26 $Y=1.16
+ $X2=0 $Y2=0
cc_465 N_A_1089_297#_c_447_n N_A_681_49#_c_1250_n 9.0109e-19 $X=7.36 $Y=1.202
+ $X2=0 $Y2=0
cc_466 N_A_1089_297#_c_448_n N_A_681_49#_c_1250_n 0.00152864f $X=7.15 $Y=0.995
+ $X2=0 $Y2=0
cc_467 N_A_1089_297#_c_450_n N_A_681_49#_c_1250_n 0.00419686f $X=8.505 $Y=0.85
+ $X2=0 $Y2=0
cc_468 N_A_1089_297#_c_451_n N_A_681_49#_c_1250_n 6.55203e-19 $X=7.315 $Y=0.85
+ $X2=0 $Y2=0
cc_469 N_A_1089_297#_c_456_n N_A_681_49#_c_1246_n 0.00139259f $X=7.36 $Y=1.41
+ $X2=0 $Y2=0
cc_470 N_A_1089_297#_M1011_g N_A_681_49#_c_1246_n 0.0164012f $X=7.385 $Y=0.455
+ $X2=0 $Y2=0
cc_471 N_A_1089_297#_c_448_n N_A_681_49#_c_1246_n 0.0173003f $X=7.15 $Y=0.995
+ $X2=0 $Y2=0
cc_472 N_A_1089_297#_c_450_n N_A_681_49#_c_1246_n 0.0173494f $X=8.505 $Y=0.85
+ $X2=0 $Y2=0
cc_473 N_A_1089_297#_c_451_n N_A_681_49#_c_1246_n 0.00232583f $X=7.315 $Y=0.85
+ $X2=0 $Y2=0
cc_474 N_A_1089_297#_c_452_n N_A_681_49#_c_1246_n 0.0185267f $X=7.17 $Y=0.85
+ $X2=0 $Y2=0
cc_475 N_A_1089_297#_c_450_n N_A_681_49#_c_1299_n 0.00166303f $X=8.505 $Y=0.85
+ $X2=0 $Y2=0
cc_476 N_A_1089_297#_c_445_n N_A_681_49#_c_1300_n 0.00333256f $X=8.88 $Y=0.945
+ $X2=0 $Y2=0
cc_477 N_A_1089_297#_c_453_n N_A_681_49#_c_1300_n 3.55136e-19 $X=8.65 $Y=0.85
+ $X2=0 $Y2=0
cc_478 N_A_1089_297#_c_454_n N_A_681_49#_c_1300_n 0.00528249f $X=8.65 $Y=0.85
+ $X2=0 $Y2=0
cc_479 N_A_1089_297#_c_461_n N_A_681_49#_c_1252_n 0.0275977f $X=5.75 $Y=1.58
+ $X2=0 $Y2=0
cc_480 N_A_1089_297#_c_448_n N_A_681_49#_c_1252_n 8.40027e-19 $X=7.15 $Y=0.995
+ $X2=0 $Y2=0
cc_481 N_A_1089_297#_c_449_n N_A_681_49#_c_1252_n 0.0525142f $X=7.025 $Y=0.85
+ $X2=0 $Y2=0
cc_482 N_A_1089_297#_c_465_p N_A_681_49#_c_1252_n 0.0124731f $X=5.835 $Y=0.85
+ $X2=0 $Y2=0
cc_483 N_A_1089_297#_c_455_n N_A_681_49#_c_1252_n 0.00234688f $X=5.81 $Y=0.74
+ $X2=0 $Y2=0
cc_484 N_A_1089_297#_c_456_n N_A_681_49#_c_1255_n 0.00348376f $X=7.36 $Y=1.41
+ $X2=0 $Y2=0
cc_485 N_A_1089_297#_c_446_n N_A_681_49#_c_1255_n 0.00431105f $X=7.26 $Y=1.16
+ $X2=0 $Y2=0
cc_486 N_A_1089_297#_c_447_n N_A_681_49#_c_1255_n 2.0806e-19 $X=7.36 $Y=1.202
+ $X2=0 $Y2=0
cc_487 N_A_1089_297#_c_448_n N_A_681_49#_c_1255_n 0.00243787f $X=7.15 $Y=0.995
+ $X2=0 $Y2=0
cc_488 N_A_1089_297#_c_451_n N_A_681_49#_c_1255_n 0.015476f $X=7.315 $Y=0.85
+ $X2=0 $Y2=0
cc_489 N_A_1089_297#_c_450_n N_A_1490_297#_M1011_d 0.00166227f $X=8.505 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_490 N_A_1089_297#_c_456_n N_A_1490_297#_c_1380_n 0.00686704f $X=7.36 $Y=1.41
+ $X2=0 $Y2=0
cc_491 N_A_1089_297#_c_450_n N_A_1490_297#_c_1380_n 0.0181022f $X=8.505 $Y=0.85
+ $X2=0 $Y2=0
cc_492 N_A_1089_297#_c_453_n N_A_1490_297#_c_1380_n 0.0020738f $X=8.65 $Y=0.85
+ $X2=0 $Y2=0
cc_493 N_A_1089_297#_c_454_n N_A_1490_297#_c_1380_n 0.00517339f $X=8.65 $Y=0.85
+ $X2=0 $Y2=0
cc_494 N_A_1089_297#_c_456_n N_A_1490_297#_c_1392_n 0.00431165f $X=7.36 $Y=1.41
+ $X2=0 $Y2=0
cc_495 N_A_1089_297#_c_458_n N_A_1490_297#_c_1393_n 0.0165035f $X=8.85 $Y=1.57
+ $X2=0 $Y2=0
cc_496 N_A_1089_297#_c_454_n N_A_1490_297#_c_1393_n 0.00161448f $X=8.65 $Y=0.85
+ $X2=0 $Y2=0
cc_497 N_A_1089_297#_c_465_p N_VGND_c_1450_n 0.00371415f $X=5.835 $Y=0.85 $X2=0
+ $Y2=0
cc_498 N_A_1089_297#_c_455_n N_VGND_c_1450_n 0.0242422f $X=5.81 $Y=0.74 $X2=0
+ $Y2=0
cc_499 N_A_1089_297#_M1011_g N_VGND_c_1456_n 0.00575161f $X=7.385 $Y=0.455 $X2=0
+ $Y2=0
cc_500 N_A_1089_297#_c_445_n N_VGND_c_1456_n 0.00585385f $X=8.88 $Y=0.945 $X2=0
+ $Y2=0
cc_501 N_A_1089_297#_c_452_n N_VGND_c_1456_n 0.00340751f $X=7.17 $Y=0.85 $X2=0
+ $Y2=0
cc_502 N_A_1089_297#_c_454_n N_VGND_c_1456_n 0.00104987f $X=8.65 $Y=0.85 $X2=0
+ $Y2=0
cc_503 N_A_1089_297#_c_455_n N_VGND_c_1456_n 0.00893636f $X=5.81 $Y=0.74 $X2=0
+ $Y2=0
cc_504 N_A_1089_297#_M1004_d N_VGND_c_1460_n 0.00248802f $X=5.625 $Y=0.235 $X2=0
+ $Y2=0
cc_505 N_A_1089_297#_M1011_g N_VGND_c_1460_n 0.00668858f $X=7.385 $Y=0.455 $X2=0
+ $Y2=0
cc_506 N_A_1089_297#_c_445_n N_VGND_c_1460_n 0.00635456f $X=8.88 $Y=0.945 $X2=0
+ $Y2=0
cc_507 N_A_1089_297#_c_449_n N_VGND_c_1460_n 0.00910735f $X=7.025 $Y=0.85 $X2=0
+ $Y2=0
cc_508 N_A_1089_297#_c_465_p N_VGND_c_1460_n 0.0148686f $X=5.835 $Y=0.85 $X2=0
+ $Y2=0
cc_509 N_A_1089_297#_c_455_n N_VGND_c_1460_n 0.00459762f $X=5.81 $Y=0.74 $X2=0
+ $Y2=0
cc_510 N_B_M1004_g N_A_1207_297#_c_796_n 0.00442504f $X=5.55 $Y=0.56 $X2=0 $Y2=0
cc_511 N_B_c_623_n N_A_1207_297#_c_809_n 0.00295958f $X=6.455 $Y=1.16 $X2=0
+ $Y2=0
cc_512 N_B_M1006_g N_A_1207_297#_c_809_n 0.00414932f $X=6.58 $Y=0.565 $X2=0
+ $Y2=0
cc_513 B N_A_1207_297#_c_803_n 0.008575f $X=8.445 $Y=1.445 $X2=0 $Y2=0
cc_514 N_B_M1006_g N_A_1207_297#_c_814_n 0.00178436f $X=6.58 $Y=0.565 $X2=0
+ $Y2=0
cc_515 N_B_c_629_n N_A_1207_297#_c_814_n 0.00325658f $X=8.265 $Y=0.995 $X2=0
+ $Y2=0
cc_516 N_B_M1004_g N_A_1207_297#_c_800_n 4.2117e-19 $X=5.55 $Y=0.56 $X2=0 $Y2=0
cc_517 N_B_M1006_g N_A_1207_297#_c_800_n 9.07111e-19 $X=6.58 $Y=0.565 $X2=0
+ $Y2=0
cc_518 N_B_c_630_n N_A_1207_297#_c_801_n 0.003607f $X=5.355 $Y=1.41 $X2=0 $Y2=0
cc_519 N_B_M1004_g N_A_1207_297#_c_801_n 0.00134479f $X=5.55 $Y=0.56 $X2=0 $Y2=0
cc_520 N_B_c_623_n N_A_1207_297#_c_801_n 0.014573f $X=6.455 $Y=1.16 $X2=0 $Y2=0
cc_521 N_B_M1008_g N_A_1207_297#_c_801_n 0.00424996f $X=6.555 $Y=1.905 $X2=0
+ $Y2=0
cc_522 N_B_M1006_g N_A_1207_297#_c_801_n 0.00389371f $X=6.58 $Y=0.565 $X2=0
+ $Y2=0
cc_523 N_B_c_626_n N_A_1207_297#_c_801_n 0.0011146f $X=6.555 $Y=1.16 $X2=0 $Y2=0
cc_524 N_B_c_630_n N_VPWR_c_934_n 0.0113699f $X=5.355 $Y=1.41 $X2=0 $Y2=0
cc_525 N_B_c_630_n N_VPWR_c_941_n 0.00455828f $X=5.355 $Y=1.41 $X2=0 $Y2=0
cc_526 N_B_c_634_n N_VPWR_c_941_n 0.0407088f $X=6.655 $Y=2.54 $X2=0 $Y2=0
cc_527 N_B_c_630_n N_VPWR_c_929_n 0.00656627f $X=5.355 $Y=1.41 $X2=0 $Y2=0
cc_528 N_B_c_633_n N_VPWR_c_929_n 0.0412005f $X=8.185 $Y=2.54 $X2=0 $Y2=0
cc_529 N_B_c_634_n N_VPWR_c_929_n 0.0071208f $X=6.655 $Y=2.54 $X2=0 $Y2=0
cc_530 N_B_M1004_g N_A_657_325#_c_1091_n 0.003112f $X=5.55 $Y=0.56 $X2=0 $Y2=0
cc_531 N_B_c_630_n N_A_657_325#_c_1092_n 0.0127882f $X=5.355 $Y=1.41 $X2=0 $Y2=0
cc_532 N_B_c_624_n N_A_657_325#_c_1092_n 0.00535881f $X=5.625 $Y=1.16 $X2=0
+ $Y2=0
cc_533 N_B_c_630_n N_A_657_325#_c_1097_n 0.0175458f $X=5.355 $Y=1.41 $X2=0 $Y2=0
cc_534 N_B_c_630_n N_A_657_325#_c_1098_n 0.00608631f $X=5.355 $Y=1.41 $X2=0
+ $Y2=0
cc_535 N_B_M1008_g N_A_657_325#_c_1098_n 8.94333e-19 $X=6.555 $Y=1.905 $X2=0
+ $Y2=0
cc_536 N_B_c_630_n N_A_657_325#_c_1100_n 0.00366198f $X=5.355 $Y=1.41 $X2=0
+ $Y2=0
cc_537 N_B_c_623_n N_A_657_325#_c_1093_n 0.00354518f $X=6.455 $Y=1.16 $X2=0
+ $Y2=0
cc_538 N_B_M1008_g N_A_657_325#_c_1093_n 0.0315935f $X=6.555 $Y=1.905 $X2=0
+ $Y2=0
cc_539 N_B_M1006_g N_A_657_325#_c_1093_n 0.0086054f $X=6.58 $Y=0.565 $X2=0 $Y2=0
cc_540 N_B_c_626_n N_A_657_325#_c_1093_n 0.0105369f $X=6.555 $Y=1.16 $X2=0 $Y2=0
cc_541 N_B_M1008_g N_A_657_325#_c_1102_n 0.00817171f $X=6.555 $Y=1.905 $X2=0
+ $Y2=0
cc_542 N_B_c_633_n N_A_657_325#_c_1102_n 0.0364604f $X=8.185 $Y=2.54 $X2=0 $Y2=0
cc_543 N_B_c_634_n N_A_657_325#_c_1102_n 2.38151e-19 $X=6.655 $Y=2.54 $X2=0
+ $Y2=0
cc_544 N_B_M1016_g N_A_657_325#_c_1102_n 0.0102069f $X=8.285 $Y=1.965 $X2=0
+ $Y2=0
cc_545 N_B_M1006_g N_A_657_325#_c_1139_n 5.90705e-19 $X=6.58 $Y=0.565 $X2=0
+ $Y2=0
cc_546 N_B_M1004_g N_A_657_325#_c_1094_n 9.01698e-19 $X=5.55 $Y=0.56 $X2=0 $Y2=0
cc_547 N_B_c_624_n N_A_657_325#_c_1094_n 0.0038653f $X=5.625 $Y=1.16 $X2=0 $Y2=0
cc_548 N_B_M1006_g N_A_657_325#_c_1142_n 0.0110774f $X=6.58 $Y=0.565 $X2=0 $Y2=0
cc_549 N_B_M1008_g N_A_657_325#_c_1104_n 0.00716396f $X=6.555 $Y=1.905 $X2=0
+ $Y2=0
cc_550 N_B_c_634_n N_A_657_325#_c_1104_n 2.51585e-19 $X=6.655 $Y=2.54 $X2=0
+ $Y2=0
cc_551 N_B_c_624_n N_A_681_49#_c_1245_n 4.44674e-19 $X=5.625 $Y=1.16 $X2=0 $Y2=0
cc_552 N_B_M1008_g N_A_681_49#_c_1249_n 0.00145677f $X=6.555 $Y=1.905 $X2=0
+ $Y2=0
cc_553 N_B_M1008_g N_A_681_49#_c_1286_n 0.00446449f $X=6.555 $Y=1.905 $X2=0
+ $Y2=0
cc_554 N_B_c_629_n N_A_681_49#_c_1246_n 0.0026019f $X=8.265 $Y=0.995 $X2=0 $Y2=0
cc_555 N_B_c_627_n N_A_681_49#_c_1299_n 0.0029291f $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_556 N_B_c_628_n N_A_681_49#_c_1299_n 4.30216e-19 $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_557 N_B_c_629_n N_A_681_49#_c_1299_n 0.00498906f $X=8.265 $Y=0.995 $X2=0
+ $Y2=0
cc_558 N_B_c_628_n N_A_681_49#_c_1300_n 0.00110831f $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_559 N_B_c_629_n N_A_681_49#_c_1321_n 0.00521263f $X=8.265 $Y=0.995 $X2=0
+ $Y2=0
cc_560 N_B_c_630_n N_A_681_49#_c_1252_n 0.00469456f $X=5.355 $Y=1.41 $X2=0 $Y2=0
cc_561 N_B_c_623_n N_A_681_49#_c_1252_n 0.00486395f $X=6.455 $Y=1.16 $X2=0 $Y2=0
cc_562 N_B_c_624_n N_A_681_49#_c_1252_n 2.58451e-19 $X=5.625 $Y=1.16 $X2=0 $Y2=0
cc_563 N_B_M1008_g N_A_681_49#_c_1252_n 0.00507147f $X=6.555 $Y=1.905 $X2=0
+ $Y2=0
cc_564 N_B_c_626_n N_A_681_49#_c_1252_n 2.29578e-19 $X=6.555 $Y=1.16 $X2=0 $Y2=0
cc_565 N_B_M1008_g N_A_681_49#_c_1255_n 4.48588e-19 $X=6.555 $Y=1.905 $X2=0
+ $Y2=0
cc_566 N_B_c_635_n N_A_1490_297#_c_1380_n 0.00160527f $X=8.285 $Y=1.47 $X2=0
+ $Y2=0
cc_567 N_B_M1016_g N_A_1490_297#_c_1380_n 0.00912353f $X=8.285 $Y=1.965 $X2=0
+ $Y2=0
cc_568 N_B_c_627_n N_A_1490_297#_c_1380_n 0.0332296f $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_569 N_B_c_641_n N_A_1490_297#_c_1380_n 0.0142666f $X=8.375 $Y=1.53 $X2=0
+ $Y2=0
cc_570 N_B_c_629_n N_A_1490_297#_c_1380_n 0.0105486f $X=8.265 $Y=0.995 $X2=0
+ $Y2=0
cc_571 N_B_M1016_g N_A_1490_297#_c_1393_n 0.011211f $X=8.285 $Y=1.965 $X2=0
+ $Y2=0
cc_572 N_B_c_628_n N_A_1490_297#_c_1393_n 0.00114355f $X=8.24 $Y=1.16 $X2=0
+ $Y2=0
cc_573 N_B_c_641_n N_A_1490_297#_c_1393_n 0.00934779f $X=8.375 $Y=1.53 $X2=0
+ $Y2=0
cc_574 B N_A_1490_297#_c_1393_n 0.0165342f $X=8.445 $Y=1.445 $X2=0 $Y2=0
cc_575 N_B_M1004_g N_VGND_c_1450_n 0.00883459f $X=5.55 $Y=0.56 $X2=0 $Y2=0
cc_576 N_B_c_624_n N_VGND_c_1450_n 0.00541821f $X=5.625 $Y=1.16 $X2=0 $Y2=0
cc_577 N_B_M1004_g N_VGND_c_1456_n 0.00560495f $X=5.55 $Y=0.56 $X2=0 $Y2=0
cc_578 N_B_M1006_g N_VGND_c_1456_n 0.00421216f $X=6.58 $Y=0.565 $X2=0 $Y2=0
cc_579 N_B_c_629_n N_VGND_c_1456_n 0.00357877f $X=8.265 $Y=0.995 $X2=0 $Y2=0
cc_580 N_B_M1004_g N_VGND_c_1460_n 0.0109084f $X=5.55 $Y=0.56 $X2=0 $Y2=0
cc_581 N_B_M1006_g N_VGND_c_1460_n 0.0071589f $X=6.58 $Y=0.565 $X2=0 $Y2=0
cc_582 N_B_c_629_n N_VGND_c_1460_n 0.00613199f $X=8.265 $Y=0.995 $X2=0 $Y2=0
cc_583 N_A_c_756_n N_A_1207_297#_c_794_n 0.0637929f $X=9.405 $Y=1.41 $X2=0 $Y2=0
cc_584 A N_A_1207_297#_c_794_n 8.4217e-19 $X=9.295 $Y=1.105 $X2=0 $Y2=0
cc_585 N_A_c_757_n N_A_1207_297#_c_795_n 0.0202318f $X=9.43 $Y=0.995 $X2=0 $Y2=0
cc_586 N_A_c_756_n N_A_1207_297#_c_803_n 0.0144336f $X=9.405 $Y=1.41 $X2=0 $Y2=0
cc_587 A N_A_1207_297#_c_803_n 0.0301432f $X=9.295 $Y=1.105 $X2=0 $Y2=0
cc_588 N_A_c_756_n N_A_1207_297#_c_797_n 5.76324e-19 $X=9.405 $Y=1.41 $X2=0
+ $Y2=0
cc_589 N_A_c_757_n N_A_1207_297#_c_797_n 0.0114592f $X=9.43 $Y=0.995 $X2=0 $Y2=0
cc_590 A N_A_1207_297#_c_797_n 0.0142387f $X=9.295 $Y=1.105 $X2=0 $Y2=0
cc_591 N_A_c_756_n N_A_1207_297#_c_798_n 0.00444032f $X=9.405 $Y=1.41 $X2=0
+ $Y2=0
cc_592 A N_A_1207_297#_c_798_n 0.0205785f $X=9.295 $Y=1.105 $X2=0 $Y2=0
cc_593 N_A_c_756_n N_A_1207_297#_c_799_n 7.33895e-19 $X=9.405 $Y=1.41 $X2=0
+ $Y2=0
cc_594 N_A_c_757_n N_A_1207_297#_c_799_n 0.00359979f $X=9.43 $Y=0.995 $X2=0
+ $Y2=0
cc_595 A N_A_1207_297#_c_799_n 0.021115f $X=9.295 $Y=1.105 $X2=0 $Y2=0
cc_596 N_A_c_756_n N_A_1207_297#_c_805_n 0.00336141f $X=9.405 $Y=1.41 $X2=0
+ $Y2=0
cc_597 A N_A_1207_297#_c_829_n 9.51454e-19 $X=9.295 $Y=1.105 $X2=0 $Y2=0
cc_598 N_A_c_756_n N_VPWR_c_941_n 0.00309549f $X=9.405 $Y=1.41 $X2=0 $Y2=0
cc_599 N_A_c_756_n N_VPWR_c_929_n 0.00394227f $X=9.405 $Y=1.41 $X2=0 $Y2=0
cc_600 N_A_c_756_n N_VPWR_c_945_n 0.0113659f $X=9.405 $Y=1.41 $X2=0 $Y2=0
cc_601 N_A_c_756_n N_A_657_325#_c_1102_n 0.00147672f $X=9.405 $Y=1.41 $X2=0
+ $Y2=0
cc_602 N_A_c_756_n N_A_1490_297#_c_1393_n 0.0136104f $X=9.405 $Y=1.41 $X2=0
+ $Y2=0
cc_603 N_A_c_756_n N_A_1490_297#_c_1386_n 3.68126e-19 $X=9.405 $Y=1.41 $X2=0
+ $Y2=0
cc_604 N_A_c_757_n N_VGND_c_1451_n 0.00276126f $X=9.43 $Y=0.995 $X2=0 $Y2=0
cc_605 N_A_c_757_n N_VGND_c_1456_n 0.00439206f $X=9.43 $Y=0.995 $X2=0 $Y2=0
cc_606 N_A_c_757_n N_VGND_c_1460_n 0.00642697f $X=9.43 $Y=0.995 $X2=0 $Y2=0
cc_607 N_A_1207_297#_c_803_n N_VPWR_M1018_d 0.00495492f $X=9.705 $Y=1.6 $X2=0
+ $Y2=0
cc_608 N_A_1207_297#_c_794_n N_VPWR_c_942_n 0.00436183f $X=9.875 $Y=1.41 $X2=0
+ $Y2=0
cc_609 N_A_1207_297#_M1010_d N_VPWR_c_929_n 0.00402227f $X=8.94 $Y=1.645 $X2=0
+ $Y2=0
cc_610 N_A_1207_297#_c_794_n N_VPWR_c_929_n 0.00600176f $X=9.875 $Y=1.41 $X2=0
+ $Y2=0
cc_611 N_A_1207_297#_c_794_n N_VPWR_c_945_n 0.00837545f $X=9.875 $Y=1.41 $X2=0
+ $Y2=0
cc_612 N_A_1207_297#_c_814_n N_A_657_325#_M1006_d 0.00599208f $X=9.015 $Y=0.51
+ $X2=0 $Y2=0
cc_613 N_A_1207_297#_c_801_n N_A_657_325#_c_1097_n 0.0132911f $X=6.16 $Y=0.51
+ $X2=0 $Y2=0
cc_614 N_A_1207_297#_c_801_n N_A_657_325#_c_1098_n 0.00274773f $X=6.16 $Y=0.51
+ $X2=0 $Y2=0
cc_615 N_A_1207_297#_M1008_s N_A_657_325#_c_1099_n 0.0102858f $X=6.035 $Y=1.485
+ $X2=0 $Y2=0
cc_616 N_A_1207_297#_c_801_n N_A_657_325#_c_1099_n 0.0128549f $X=6.16 $Y=0.51
+ $X2=0 $Y2=0
cc_617 N_A_1207_297#_M1006_s N_A_657_325#_c_1093_n 2.84455e-19 $X=6.205 $Y=0.245
+ $X2=0 $Y2=0
cc_618 N_A_1207_297#_c_801_n N_A_657_325#_c_1093_n 0.072119f $X=6.16 $Y=0.51
+ $X2=0 $Y2=0
cc_619 N_A_1207_297#_M1010_d N_A_657_325#_c_1102_n 0.00261136f $X=8.94 $Y=1.645
+ $X2=0 $Y2=0
cc_620 N_A_1207_297#_c_809_n N_A_657_325#_c_1139_n 0.00646194f $X=6.355 $Y=0.4
+ $X2=0 $Y2=0
cc_621 N_A_1207_297#_c_814_n N_A_657_325#_c_1139_n 0.0112439f $X=9.015 $Y=0.51
+ $X2=0 $Y2=0
cc_622 N_A_1207_297#_c_800_n N_A_657_325#_c_1139_n 0.00136926f $X=6.315 $Y=0.51
+ $X2=0 $Y2=0
cc_623 N_A_1207_297#_c_801_n N_A_657_325#_c_1139_n 0.00265819f $X=6.16 $Y=0.51
+ $X2=0 $Y2=0
cc_624 N_A_1207_297#_M1006_s N_A_657_325#_c_1142_n 0.00187185f $X=6.205 $Y=0.245
+ $X2=0 $Y2=0
cc_625 N_A_1207_297#_c_809_n N_A_657_325#_c_1142_n 0.00399903f $X=6.355 $Y=0.4
+ $X2=0 $Y2=0
cc_626 N_A_1207_297#_c_814_n N_A_657_325#_c_1142_n 0.0032462f $X=9.015 $Y=0.51
+ $X2=0 $Y2=0
cc_627 N_A_1207_297#_c_801_n N_A_657_325#_c_1142_n 0.012754f $X=6.16 $Y=0.51
+ $X2=0 $Y2=0
cc_628 N_A_1207_297#_c_814_n N_A_681_49#_M1014_d 0.00427772f $X=9.015 $Y=0.51
+ $X2=0 $Y2=0
cc_629 N_A_1207_297#_c_814_n N_A_681_49#_c_1246_n 0.0147234f $X=9.015 $Y=0.51
+ $X2=0 $Y2=0
cc_630 N_A_1207_297#_c_814_n N_A_681_49#_c_1299_n 0.00610486f $X=9.015 $Y=0.51
+ $X2=0 $Y2=0
cc_631 N_A_1207_297#_c_814_n N_A_681_49#_c_1300_n 0.00980954f $X=9.015 $Y=0.51
+ $X2=0 $Y2=0
cc_632 N_A_1207_297#_c_829_n N_A_681_49#_c_1300_n 0.0012274f $X=9.16 $Y=0.51
+ $X2=0 $Y2=0
cc_633 N_A_1207_297#_c_830_n N_A_681_49#_c_1300_n 0.00676874f $X=9.16 $Y=0.51
+ $X2=0 $Y2=0
cc_634 N_A_1207_297#_c_814_n N_A_681_49#_c_1321_n 0.0119237f $X=9.015 $Y=0.51
+ $X2=0 $Y2=0
cc_635 N_A_1207_297#_M1008_s N_A_681_49#_c_1252_n 0.00802537f $X=6.035 $Y=1.485
+ $X2=0 $Y2=0
cc_636 N_A_1207_297#_c_801_n N_A_681_49#_c_1252_n 0.0183124f $X=6.16 $Y=0.51
+ $X2=0 $Y2=0
cc_637 N_A_1207_297#_c_814_n N_A_1490_297#_M1011_d 0.00653094f $X=9.015 $Y=0.51
+ $X2=-0.19 $Y2=-0.24
cc_638 N_A_1207_297#_c_814_n N_A_1490_297#_c_1380_n 0.00162336f $X=9.015 $Y=0.51
+ $X2=0 $Y2=0
cc_639 N_A_1207_297#_c_794_n N_A_1490_297#_c_1381_n 0.0195627f $X=9.875 $Y=1.41
+ $X2=0 $Y2=0
cc_640 N_A_1207_297#_c_795_n N_A_1490_297#_c_1381_n 0.0097849f $X=9.9 $Y=0.995
+ $X2=0 $Y2=0
cc_641 N_A_1207_297#_c_803_n N_A_1490_297#_c_1381_n 0.0112214f $X=9.705 $Y=1.6
+ $X2=0 $Y2=0
cc_642 N_A_1207_297#_c_799_n N_A_1490_297#_c_1381_n 0.0381742f $X=9.79 $Y=1.325
+ $X2=0 $Y2=0
cc_643 N_A_1207_297#_c_805_n N_A_1490_297#_c_1381_n 0.00830381f $X=9.79 $Y=1.495
+ $X2=0 $Y2=0
cc_644 N_A_1207_297#_M1010_d N_A_1490_297#_c_1393_n 0.00774465f $X=8.94 $Y=1.645
+ $X2=0 $Y2=0
cc_645 N_A_1207_297#_c_794_n N_A_1490_297#_c_1393_n 0.00221849f $X=9.875 $Y=1.41
+ $X2=0 $Y2=0
cc_646 N_A_1207_297#_c_803_n N_A_1490_297#_c_1393_n 0.0353842f $X=9.705 $Y=1.6
+ $X2=0 $Y2=0
cc_647 N_A_1207_297#_c_794_n N_A_1490_297#_c_1386_n 0.0126341f $X=9.875 $Y=1.41
+ $X2=0 $Y2=0
cc_648 N_A_1207_297#_c_803_n N_A_1490_297#_c_1386_n 0.00653478f $X=9.705 $Y=1.6
+ $X2=0 $Y2=0
cc_649 N_A_1207_297#_c_799_n N_A_1490_297#_c_1386_n 0.00278512f $X=9.79 $Y=1.325
+ $X2=0 $Y2=0
cc_650 N_A_1207_297#_c_794_n N_A_1490_297#_c_1382_n 2.03932e-19 $X=9.875 $Y=1.41
+ $X2=0 $Y2=0
cc_651 N_A_1207_297#_c_797_n N_VGND_M1003_d 0.00147467f $X=9.705 $Y=0.82 $X2=0
+ $Y2=0
cc_652 N_A_1207_297#_c_799_n N_VGND_M1003_d 0.00108061f $X=9.79 $Y=1.325 $X2=0
+ $Y2=0
cc_653 N_A_1207_297#_c_795_n N_VGND_c_1451_n 0.00414899f $X=9.9 $Y=0.995 $X2=0
+ $Y2=0
cc_654 N_A_1207_297#_c_797_n N_VGND_c_1451_n 0.0111874f $X=9.705 $Y=0.82 $X2=0
+ $Y2=0
cc_655 N_A_1207_297#_c_799_n N_VGND_c_1451_n 0.00164729f $X=9.79 $Y=1.325 $X2=0
+ $Y2=0
cc_656 N_A_1207_297#_c_829_n N_VGND_c_1451_n 0.00112928f $X=9.16 $Y=0.51 $X2=0
+ $Y2=0
cc_657 N_A_1207_297#_c_796_n N_VGND_c_1456_n 0.0114103f $X=6.245 $Y=0.375 $X2=0
+ $Y2=0
cc_658 N_A_1207_297#_c_809_n N_VGND_c_1456_n 0.0150413f $X=6.355 $Y=0.4 $X2=0
+ $Y2=0
cc_659 N_A_1207_297#_c_797_n N_VGND_c_1456_n 0.00248202f $X=9.705 $Y=0.82 $X2=0
+ $Y2=0
cc_660 N_A_1207_297#_c_814_n N_VGND_c_1456_n 0.00568764f $X=9.015 $Y=0.51 $X2=0
+ $Y2=0
cc_661 N_A_1207_297#_c_800_n N_VGND_c_1456_n 4.91623e-19 $X=6.315 $Y=0.51 $X2=0
+ $Y2=0
cc_662 N_A_1207_297#_c_829_n N_VGND_c_1456_n 3.63685e-19 $X=9.16 $Y=0.51 $X2=0
+ $Y2=0
cc_663 N_A_1207_297#_c_830_n N_VGND_c_1456_n 0.0149689f $X=9.16 $Y=0.51 $X2=0
+ $Y2=0
cc_664 N_A_1207_297#_c_795_n N_VGND_c_1459_n 0.00536613f $X=9.9 $Y=0.995 $X2=0
+ $Y2=0
cc_665 N_A_1207_297#_c_799_n N_VGND_c_1459_n 0.00182428f $X=9.79 $Y=1.325 $X2=0
+ $Y2=0
cc_666 N_A_1207_297#_M1015_d N_VGND_c_1460_n 0.00240207f $X=8.955 $Y=0.235 $X2=0
+ $Y2=0
cc_667 N_A_1207_297#_c_795_n N_VGND_c_1460_n 0.0103767f $X=9.9 $Y=0.995 $X2=0
+ $Y2=0
cc_668 N_A_1207_297#_c_796_n N_VGND_c_1460_n 0.00165885f $X=6.245 $Y=0.375 $X2=0
+ $Y2=0
cc_669 N_A_1207_297#_c_809_n N_VGND_c_1460_n 0.00259517f $X=6.355 $Y=0.4 $X2=0
+ $Y2=0
cc_670 N_A_1207_297#_c_797_n N_VGND_c_1460_n 0.00552122f $X=9.705 $Y=0.82 $X2=0
+ $Y2=0
cc_671 N_A_1207_297#_c_799_n N_VGND_c_1460_n 0.00402105f $X=9.79 $Y=1.325 $X2=0
+ $Y2=0
cc_672 N_A_1207_297#_c_814_n N_VGND_c_1460_n 0.235445f $X=9.015 $Y=0.51 $X2=0
+ $Y2=0
cc_673 N_A_1207_297#_c_800_n N_VGND_c_1460_n 0.0297997f $X=6.315 $Y=0.51 $X2=0
+ $Y2=0
cc_674 N_A_1207_297#_c_829_n N_VGND_c_1460_n 0.0285254f $X=9.16 $Y=0.51 $X2=0
+ $Y2=0
cc_675 N_A_1207_297#_c_830_n N_VGND_c_1460_n 0.0036194f $X=9.16 $Y=0.51 $X2=0
+ $Y2=0
cc_676 N_VPWR_c_929_n N_X_M1000_d 0.00233757f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_677 N_VPWR_c_929_n N_X_M1022_d 0.00439555f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_678 N_VPWR_c_930_n N_X_c_1051_n 0.0698025f $X=0.37 $Y=1.66 $X2=0 $Y2=0
cc_679 N_VPWR_c_931_n N_X_c_1051_n 0.0569238f $X=1.31 $Y=1.66 $X2=0 $Y2=0
cc_680 N_VPWR_c_937_n N_X_c_1051_n 0.0178128f $X=1.225 $Y=2.72 $X2=0 $Y2=0
cc_681 N_VPWR_c_929_n N_X_c_1051_n 0.0137157f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_682 N_VPWR_c_931_n N_X_c_1055_n 0.0138735f $X=1.31 $Y=1.66 $X2=0 $Y2=0
cc_683 N_VPWR_c_931_n N_X_c_1047_n 0.00816305f $X=1.31 $Y=1.66 $X2=0 $Y2=0
cc_684 N_VPWR_c_931_n N_X_c_1067_n 0.0634618f $X=1.31 $Y=1.66 $X2=0 $Y2=0
cc_685 N_VPWR_c_932_n N_X_c_1067_n 0.0208347f $X=2.065 $Y=2.72 $X2=0 $Y2=0
cc_686 N_VPWR_c_933_n N_X_c_1067_n 0.01963f $X=2.285 $Y=2.3 $X2=0 $Y2=0
cc_687 N_VPWR_c_929_n N_X_c_1067_n 0.0121067f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_688 N_VPWR_c_929_n N_A_657_325#_M1016_d 0.00241089f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_689 N_VPWR_c_934_n N_A_657_325#_c_1095_n 0.00147971f $X=5.12 $Y=2.32 $X2=0
+ $Y2=0
cc_690 N_VPWR_c_939_n N_A_657_325#_c_1095_n 0.012236f $X=4.955 $Y=2.72 $X2=0
+ $Y2=0
cc_691 N_VPWR_c_929_n N_A_657_325#_c_1095_n 0.0223233f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_692 N_VPWR_M1027_s N_A_657_325#_c_1092_n 0.00648603f $X=4.995 $Y=2.175 $X2=0
+ $Y2=0
cc_693 N_VPWR_M1027_s N_A_657_325#_c_1097_n 0.00155527f $X=4.995 $Y=2.175 $X2=0
+ $Y2=0
cc_694 N_VPWR_c_934_n N_A_657_325#_c_1097_n 0.00612755f $X=5.12 $Y=2.32 $X2=0
+ $Y2=0
cc_695 N_VPWR_c_941_n N_A_657_325#_c_1097_n 0.00666556f $X=9.425 $Y=2.72 $X2=0
+ $Y2=0
cc_696 N_VPWR_c_929_n N_A_657_325#_c_1097_n 0.0119497f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_697 N_VPWR_c_934_n N_A_657_325#_c_1098_n 0.00140976f $X=5.12 $Y=2.32 $X2=0
+ $Y2=0
cc_698 N_VPWR_c_941_n N_A_657_325#_c_1099_n 0.0300226f $X=9.425 $Y=2.72 $X2=0
+ $Y2=0
cc_699 N_VPWR_c_929_n N_A_657_325#_c_1099_n 0.0193106f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_700 N_VPWR_c_934_n N_A_657_325#_c_1100_n 0.00679194f $X=5.12 $Y=2.32 $X2=0
+ $Y2=0
cc_701 N_VPWR_c_941_n N_A_657_325#_c_1100_n 0.0105925f $X=9.425 $Y=2.72 $X2=0
+ $Y2=0
cc_702 N_VPWR_c_929_n N_A_657_325#_c_1100_n 0.00644598f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_703 N_VPWR_c_941_n N_A_657_325#_c_1102_n 0.134682f $X=9.425 $Y=2.72 $X2=0
+ $Y2=0
cc_704 N_VPWR_c_929_n N_A_657_325#_c_1102_n 0.0811181f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_705 N_VPWR_c_945_n N_A_657_325#_c_1102_n 0.00711003f $X=9.64 $Y=2.36 $X2=0
+ $Y2=0
cc_706 N_VPWR_M1027_s N_A_657_325#_c_1103_n 0.00233831f $X=4.995 $Y=2.175 $X2=0
+ $Y2=0
cc_707 N_VPWR_c_934_n N_A_657_325#_c_1103_n 0.0144069f $X=5.12 $Y=2.32 $X2=0
+ $Y2=0
cc_708 N_VPWR_c_929_n N_A_657_325#_c_1103_n 8.22076e-19 $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_709 N_VPWR_c_941_n N_A_657_325#_c_1104_n 0.0103509f $X=9.425 $Y=2.72 $X2=0
+ $Y2=0
cc_710 N_VPWR_c_929_n N_A_657_325#_c_1104_n 0.00587789f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_711 N_VPWR_M1027_s N_A_681_49#_c_1252_n 0.00109947f $X=4.995 $Y=2.175 $X2=0
+ $Y2=0
cc_712 N_VPWR_c_929_n N_A_1490_297#_M1013_d 0.00259864f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_713 N_VPWR_c_942_n N_A_1490_297#_c_1384_n 0.0197624f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_714 N_VPWR_c_929_n N_A_1490_297#_c_1384_n 0.0111058f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_715 N_VPWR_c_945_n N_A_1490_297#_c_1384_n 0.0121318f $X=9.64 $Y=2.36 $X2=0
+ $Y2=0
cc_716 N_VPWR_M1018_d N_A_1490_297#_c_1393_n 0.00390782f $X=9.495 $Y=1.485 $X2=0
+ $Y2=0
cc_717 N_VPWR_c_941_n N_A_1490_297#_c_1393_n 0.00692236f $X=9.425 $Y=2.72 $X2=0
+ $Y2=0
cc_718 N_VPWR_c_929_n N_A_1490_297#_c_1393_n 0.0149452f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_719 N_VPWR_c_945_n N_A_1490_297#_c_1393_n 0.0198562f $X=9.64 $Y=2.36 $X2=0
+ $Y2=0
cc_720 N_VPWR_c_942_n N_A_1490_297#_c_1386_n 0.00346082f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_721 N_VPWR_c_929_n N_A_1490_297#_c_1386_n 0.00566025f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_722 N_X_c_1055_n N_VGND_c_1447_n 0.0100081f $X=1.565 $Y=1.16 $X2=0 $Y2=0
cc_723 N_X_c_1056_n N_VGND_c_1447_n 0.0282893f $X=1.79 $Y=0.56 $X2=0 $Y2=0
cc_724 N_X_c_1056_n N_VGND_c_1448_n 0.0120203f $X=1.79 $Y=0.56 $X2=0 $Y2=0
cc_725 N_X_c_1046_n N_VGND_c_1454_n 0.0105213f $X=0.84 $Y=0.56 $X2=0 $Y2=0
cc_726 N_X_M1005_s N_VGND_c_1460_n 0.00448447f $X=0.655 $Y=0.235 $X2=0 $Y2=0
cc_727 N_X_M1009_s N_VGND_c_1460_n 0.00443674f $X=1.605 $Y=0.235 $X2=0 $Y2=0
cc_728 N_X_c_1046_n N_VGND_c_1460_n 0.010586f $X=0.84 $Y=0.56 $X2=0 $Y2=0
cc_729 N_X_c_1056_n N_VGND_c_1460_n 0.0110799f $X=1.79 $Y=0.56 $X2=0 $Y2=0
cc_730 N_A_657_325#_c_1095_n N_A_681_49#_M1025_d 0.012215f $X=4.975 $Y=1.98
+ $X2=0 $Y2=0
cc_731 N_A_657_325#_c_1102_n N_A_681_49#_M1008_d 0.00924946f $X=8.605 $Y=2.36
+ $X2=0 $Y2=0
cc_732 N_A_657_325#_M1020_d N_A_681_49#_c_1257_n 0.00773142f $X=4.405 $Y=0.245
+ $X2=0 $Y2=0
cc_733 N_A_657_325#_c_1090_n N_A_681_49#_c_1257_n 0.0173367f $X=4.865 $Y=0.37
+ $X2=0 $Y2=0
cc_734 N_A_657_325#_c_1091_n N_A_681_49#_c_1257_n 0.0140571f $X=4.95 $Y=1.035
+ $X2=0 $Y2=0
cc_735 N_A_657_325#_M1020_d N_A_681_49#_c_1245_n 0.00248769f $X=4.405 $Y=0.245
+ $X2=0 $Y2=0
cc_736 N_A_657_325#_c_1091_n N_A_681_49#_c_1245_n 0.0179156f $X=4.95 $Y=1.035
+ $X2=0 $Y2=0
cc_737 N_A_657_325#_c_1092_n N_A_681_49#_c_1245_n 0.00902524f $X=5.06 $Y=1.895
+ $X2=0 $Y2=0
cc_738 N_A_657_325#_c_1094_n N_A_681_49#_c_1245_n 0.0132103f $X=5.06 $Y=1.12
+ $X2=0 $Y2=0
cc_739 N_A_657_325#_c_1093_n N_A_681_49#_c_1249_n 0.00870819f $X=6.5 $Y=2.275
+ $X2=0 $Y2=0
cc_740 N_A_657_325#_c_1142_n N_A_681_49#_c_1249_n 2.50678e-19 $X=6.79 $Y=0.74
+ $X2=0 $Y2=0
cc_741 N_A_657_325#_c_1093_n N_A_681_49#_c_1286_n 0.0255541f $X=6.5 $Y=2.275
+ $X2=0 $Y2=0
cc_742 N_A_657_325#_c_1102_n N_A_681_49#_c_1286_n 0.0238103f $X=8.605 $Y=2.36
+ $X2=0 $Y2=0
cc_743 N_A_657_325#_c_1102_n N_A_681_49#_c_1250_n 0.0100462f $X=8.605 $Y=2.36
+ $X2=0 $Y2=0
cc_744 N_A_657_325#_c_1139_n N_A_681_49#_c_1246_n 0.00253431f $X=6.79 $Y=0.545
+ $X2=0 $Y2=0
cc_745 N_A_657_325#_c_1095_n N_A_681_49#_c_1252_n 0.00437461f $X=4.975 $Y=1.98
+ $X2=0 $Y2=0
cc_746 N_A_657_325#_c_1092_n N_A_681_49#_c_1252_n 0.0161183f $X=5.06 $Y=1.895
+ $X2=0 $Y2=0
cc_747 N_A_657_325#_c_1097_n N_A_681_49#_c_1252_n 0.01149f $X=5.72 $Y=1.98 $X2=0
+ $Y2=0
cc_748 N_A_657_325#_c_1093_n N_A_681_49#_c_1252_n 0.0194408f $X=6.5 $Y=2.275
+ $X2=0 $Y2=0
cc_749 N_A_657_325#_c_1094_n N_A_681_49#_c_1252_n 0.0052436f $X=5.06 $Y=1.12
+ $X2=0 $Y2=0
cc_750 N_A_657_325#_c_1095_n N_A_681_49#_c_1253_n 0.00415423f $X=4.975 $Y=1.98
+ $X2=0 $Y2=0
cc_751 N_A_657_325#_c_1092_n N_A_681_49#_c_1253_n 0.00275249f $X=5.06 $Y=1.895
+ $X2=0 $Y2=0
cc_752 N_A_657_325#_c_1095_n N_A_681_49#_c_1254_n 0.0251846f $X=4.975 $Y=1.98
+ $X2=0 $Y2=0
cc_753 N_A_657_325#_c_1092_n N_A_681_49#_c_1254_n 0.0231767f $X=5.06 $Y=1.895
+ $X2=0 $Y2=0
cc_754 N_A_657_325#_c_1093_n N_A_681_49#_c_1255_n 0.00127808f $X=6.5 $Y=2.275
+ $X2=0 $Y2=0
cc_755 N_A_657_325#_c_1102_n N_A_1490_297#_M1021_d 0.00563686f $X=8.605 $Y=2.36
+ $X2=0 $Y2=0
cc_756 N_A_657_325#_c_1102_n N_A_1490_297#_c_1392_n 0.0129278f $X=8.605 $Y=2.36
+ $X2=0 $Y2=0
cc_757 N_A_657_325#_M1016_d N_A_1490_297#_c_1393_n 0.00678674f $X=8.375 $Y=1.645
+ $X2=0 $Y2=0
cc_758 N_A_657_325#_c_1102_n N_A_1490_297#_c_1393_n 0.0533312f $X=8.605 $Y=2.36
+ $X2=0 $Y2=0
cc_759 N_A_657_325#_c_1090_n N_VGND_c_1450_n 0.0140422f $X=4.865 $Y=0.37 $X2=0
+ $Y2=0
cc_760 N_A_657_325#_c_1091_n N_VGND_c_1450_n 0.0299543f $X=4.95 $Y=1.035 $X2=0
+ $Y2=0
cc_761 N_A_657_325#_c_1139_n N_VGND_c_1456_n 0.00778982f $X=6.79 $Y=0.545 $X2=0
+ $Y2=0
cc_762 N_A_657_325#_c_1142_n N_VGND_c_1456_n 0.00236041f $X=6.79 $Y=0.74 $X2=0
+ $Y2=0
cc_763 N_A_657_325#_c_1090_n N_VGND_c_1458_n 0.0335486f $X=4.865 $Y=0.37 $X2=0
+ $Y2=0
cc_764 N_A_657_325#_c_1090_n N_VGND_c_1460_n 0.0232648f $X=4.865 $Y=0.37 $X2=0
+ $Y2=0
cc_765 N_A_657_325#_c_1139_n N_VGND_c_1460_n 0.00172658f $X=6.79 $Y=0.545 $X2=0
+ $Y2=0
cc_766 N_A_657_325#_c_1142_n N_VGND_c_1460_n 4.40711e-19 $X=6.79 $Y=0.74 $X2=0
+ $Y2=0
cc_767 N_A_681_49#_c_1246_n N_A_1490_297#_M1011_d 0.00729398f $X=7.56 $Y=1.445
+ $X2=-0.19 $Y2=-0.24
cc_768 N_A_681_49#_c_1364_p N_A_1490_297#_M1011_d 0.0024562f $X=7.645 $Y=0.34
+ $X2=-0.19 $Y2=-0.24
cc_769 N_A_681_49#_c_1321_n N_A_1490_297#_M1011_d 0.0107136f $X=8.155 $Y=0.36
+ $X2=-0.19 $Y2=-0.24
cc_770 N_A_681_49#_c_1250_n N_A_1490_297#_M1021_d 0.00444096f $X=7.475 $Y=1.53
+ $X2=0 $Y2=0
cc_771 N_A_681_49#_c_1286_n N_A_1490_297#_c_1380_n 0.00453141f $X=6.99 $Y=1.62
+ $X2=0 $Y2=0
cc_772 N_A_681_49#_c_1250_n N_A_1490_297#_c_1380_n 0.013519f $X=7.475 $Y=1.53
+ $X2=0 $Y2=0
cc_773 N_A_681_49#_c_1246_n N_A_1490_297#_c_1380_n 0.062318f $X=7.56 $Y=1.445
+ $X2=0 $Y2=0
cc_774 N_A_681_49#_c_1321_n N_A_1490_297#_c_1380_n 0.0106102f $X=8.155 $Y=0.36
+ $X2=0 $Y2=0
cc_775 N_A_681_49#_c_1255_n N_A_1490_297#_c_1380_n 0.00130235f $X=7.17 $Y=1.53
+ $X2=0 $Y2=0
cc_776 N_A_681_49#_c_1252_n N_VGND_c_1450_n 0.00557009f $X=7.025 $Y=1.53 $X2=0
+ $Y2=0
cc_777 N_A_681_49#_c_1364_p N_VGND_c_1456_n 0.0104913f $X=7.645 $Y=0.34 $X2=0
+ $Y2=0
cc_778 N_A_681_49#_c_1321_n N_VGND_c_1456_n 0.0617902f $X=8.155 $Y=0.36 $X2=0
+ $Y2=0
cc_779 N_A_681_49#_c_1257_n N_VGND_c_1458_n 0.00331785f $X=4.525 $Y=0.71 $X2=0
+ $Y2=0
cc_780 N_A_681_49#_M1014_d N_VGND_c_1460_n 0.00231474f $X=8.255 $Y=0.245 $X2=0
+ $Y2=0
cc_781 N_A_681_49#_c_1364_p N_VGND_c_1460_n 0.00184693f $X=7.645 $Y=0.34 $X2=0
+ $Y2=0
cc_782 N_A_681_49#_c_1247_n N_VGND_c_1460_n 0.00750432f $X=3.755 $Y=0.765 $X2=0
+ $Y2=0
cc_783 N_A_681_49#_c_1321_n N_VGND_c_1460_n 0.00974346f $X=8.155 $Y=0.36 $X2=0
+ $Y2=0
cc_784 N_A_1490_297#_c_1382_n N_VGND_c_1459_n 0.0197576f $X=10.24 $Y=0.42 $X2=0
+ $Y2=0
cc_785 N_A_1490_297#_M1001_d N_VGND_c_1460_n 0.00399944f $X=9.975 $Y=0.235 $X2=0
+ $Y2=0
cc_786 N_A_1490_297#_c_1382_n N_VGND_c_1460_n 0.0113402f $X=10.24 $Y=0.42 $X2=0
+ $Y2=0
