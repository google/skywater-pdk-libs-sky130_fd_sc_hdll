* File: sky130_fd_sc_hdll__a211oi_1.pxi.spice
* Created: Wed Sep  2 08:16:02 2020
* 
x_PM_SKY130_FD_SC_HDLL__A211OI_1%A2 N_A2_c_40_n N_A2_M1000_g N_A2_c_41_n
+ N_A2_M1002_g A2 A2 PM_SKY130_FD_SC_HDLL__A211OI_1%A2
x_PM_SKY130_FD_SC_HDLL__A211OI_1%A1 N_A1_c_66_n N_A1_M1006_g N_A1_c_67_n
+ N_A1_M1003_g A1 A1 A1 A1 N_A1_c_70_n A1 PM_SKY130_FD_SC_HDLL__A211OI_1%A1
x_PM_SKY130_FD_SC_HDLL__A211OI_1%B1 N_B1_c_103_n N_B1_M1004_g N_B1_c_104_n
+ N_B1_M1005_g B1 B1 B1 B1 PM_SKY130_FD_SC_HDLL__A211OI_1%B1
x_PM_SKY130_FD_SC_HDLL__A211OI_1%C1 N_C1_c_139_n N_C1_M1007_g N_C1_c_140_n
+ N_C1_M1001_g C1 C1 PM_SKY130_FD_SC_HDLL__A211OI_1%C1
x_PM_SKY130_FD_SC_HDLL__A211OI_1%A_27_297# N_A_27_297#_M1000_s
+ N_A_27_297#_M1003_d N_A_27_297#_c_164_n N_A_27_297#_c_166_n
+ N_A_27_297#_c_165_n N_A_27_297#_c_175_n
+ PM_SKY130_FD_SC_HDLL__A211OI_1%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A211OI_1%VPWR N_VPWR_M1000_d N_VPWR_c_186_n VPWR
+ N_VPWR_c_187_n N_VPWR_c_188_n N_VPWR_c_185_n N_VPWR_c_190_n
+ PM_SKY130_FD_SC_HDLL__A211OI_1%VPWR
x_PM_SKY130_FD_SC_HDLL__A211OI_1%Y N_Y_M1006_d N_Y_M1007_d N_Y_M1001_d
+ N_Y_c_222_n N_Y_c_229_n N_Y_c_224_n N_Y_c_239_n Y Y Y Y Y N_Y_c_218_n Y Y Y
+ N_Y_c_221_n PM_SKY130_FD_SC_HDLL__A211OI_1%Y
x_PM_SKY130_FD_SC_HDLL__A211OI_1%VGND N_VGND_M1002_s N_VGND_M1004_d
+ N_VGND_c_261_n N_VGND_c_262_n VGND N_VGND_c_263_n N_VGND_c_264_n
+ N_VGND_c_265_n N_VGND_c_266_n PM_SKY130_FD_SC_HDLL__A211OI_1%VGND
cc_1 VNB N_A2_c_40_n 0.0341439f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_2 VNB N_A2_c_41_n 0.0188967f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_3 VNB A2 0.0212481f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_4 VNB N_A1_c_66_n 0.0169847f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_5 VNB N_A1_c_67_n 0.0252735f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_6 VNB A1 0.00256584f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_B1_c_103_n 0.017853f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_8 VNB N_B1_c_104_n 0.0214878f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_9 VNB B1 0.00390232f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_10 VNB N_C1_c_139_n 0.0205131f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_11 VNB N_C1_c_140_n 0.0289013f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_12 VNB C1 0.0017591f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_13 VNB N_VPWR_c_185_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_Y_c_218_n 0.0114896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB Y 0.0245525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_261_n 0.0114263f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_17 VNB N_VGND_c_262_n 0.0204545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_263_n 0.0292988f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_19 VNB N_VGND_c_264_n 0.0242776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_265_n 0.163467f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_266_n 0.00910682f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VPB N_A2_c_40_n 0.0364252f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_23 VPB A2 0.00477054f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_24 VPB N_A1_c_67_n 0.0270266f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_25 VPB N_A1_c_70_n 0.00283353f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.19
cc_26 VPB A1 6.65681e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_B1_c_104_n 0.026042f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_28 VPB B1 0.00110563f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_29 VPB N_C1_c_140_n 0.0320404f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_30 VPB C1 0.00148303f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_31 VPB N_A_27_297#_c_164_n 0.0265691f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_A_27_297#_c_165_n 0.00831871f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.16
cc_33 VPB N_VPWR_c_186_n 4.89699e-19 $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.56
cc_34 VPB N_VPWR_c_187_n 0.0161515f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_188_n 0.0487876f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_185_n 0.0469647f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_190_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB Y 0.0218549f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_Y_c_221_n 0.0331674f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 N_A2_c_41_n N_A1_c_66_n 0.0294911f $X=0.54 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_41 N_A2_c_40_n N_A1_c_67_n 0.0523054f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_42 A2 N_A1_c_67_n 2.07167e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_43 N_A2_c_41_n A1 0.0213264f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_44 A2 A1 0.0130235f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_45 N_A2_c_40_n N_A1_c_70_n 0.00908991f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_46 A2 N_A1_c_70_n 0.0263836f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_47 N_A2_c_40_n N_A_27_297#_c_166_n 0.0224457f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_48 A2 N_A_27_297#_c_166_n 0.00239276f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_49 N_A2_c_40_n N_A_27_297#_c_165_n 0.00121736f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_50 A2 N_A_27_297#_c_165_n 0.0191291f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_51 N_A2_c_40_n N_VPWR_c_186_n 0.015683f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_52 N_A2_c_40_n N_VPWR_c_187_n 0.0046653f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_53 N_A2_c_40_n N_VPWR_c_185_n 0.00898723f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_54 A2 N_VGND_M1002_s 0.00369942f $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_55 N_A2_c_40_n N_VGND_c_262_n 9.47949e-19 $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_56 N_A2_c_41_n N_VGND_c_262_n 0.0116654f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_57 A2 N_VGND_c_262_n 0.0270041f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_58 N_A2_c_41_n N_VGND_c_263_n 0.00571847f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_59 N_A2_c_41_n N_VGND_c_265_n 0.011451f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_60 A2 N_VGND_c_265_n 0.00167448f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_61 N_A1_c_66_n N_B1_c_103_n 0.0153237f $X=0.975 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_62 A1 N_B1_c_103_n 9.02406e-19 $X=0.605 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_63 N_A1_c_67_n N_B1_c_104_n 0.0489878f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_64 A1 N_B1_c_104_n 0.00229471f $X=1.15 $Y=1.19 $X2=0 $Y2=0
cc_65 N_A1_c_67_n B1 0.00155593f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_66 A1 B1 0.0226186f $X=1.15 $Y=1.19 $X2=0 $Y2=0
cc_67 N_A1_c_67_n N_A_27_297#_c_166_n 0.0194185f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_68 N_A1_c_70_n N_A_27_297#_c_166_n 0.0187334f $X=0.755 $Y=0.995 $X2=0 $Y2=0
cc_69 A1 N_A_27_297#_c_166_n 0.0233502f $X=1.15 $Y=1.19 $X2=0 $Y2=0
cc_70 N_A1_c_67_n N_VPWR_c_186_n 0.0117288f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_71 N_A1_c_67_n N_VPWR_c_188_n 0.00642146f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A1_c_67_n N_VPWR_c_185_n 0.0109646f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_73 N_A1_c_66_n N_Y_c_222_n 0.00164999f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_74 A1 N_Y_c_222_n 0.0197166f $X=0.605 $Y=0.425 $X2=0 $Y2=0
cc_75 N_A1_c_66_n N_Y_c_224_n 0.0013902f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_76 N_A1_c_67_n N_Y_c_224_n 0.00160971f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_77 A1 N_Y_c_224_n 0.0115859f $X=0.605 $Y=0.425 $X2=0 $Y2=0
cc_78 A1 N_Y_c_224_n 0.00993836f $X=1.15 $Y=1.19 $X2=0 $Y2=0
cc_79 N_A1_c_66_n N_VGND_c_263_n 0.00579368f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_80 A1 N_VGND_c_263_n 0.0159504f $X=0.605 $Y=0.425 $X2=0 $Y2=0
cc_81 N_A1_c_66_n N_VGND_c_265_n 0.0109884f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_82 A1 N_VGND_c_265_n 0.0113624f $X=0.605 $Y=0.425 $X2=0 $Y2=0
cc_83 N_A1_c_66_n N_VGND_c_266_n 0.00109909f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_84 A1 A_123_47# 0.00171f $X=0.605 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_85 N_B1_c_103_n N_C1_c_139_n 0.0212462f $X=1.51 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_86 N_B1_c_104_n N_C1_c_140_n 0.0674145f $X=1.535 $Y=1.41 $X2=0 $Y2=0
cc_87 B1 N_C1_c_140_n 0.0106193f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_88 N_B1_c_104_n C1 5.99344e-19 $X=1.535 $Y=1.41 $X2=0 $Y2=0
cc_89 B1 C1 0.0449238f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_90 N_B1_c_104_n N_A_27_297#_c_166_n 0.00163857f $X=1.535 $Y=1.41 $X2=0 $Y2=0
cc_91 B1 N_A_27_297#_c_166_n 0.0163876f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_92 N_B1_c_104_n N_A_27_297#_c_175_n 0.0053103f $X=1.535 $Y=1.41 $X2=0 $Y2=0
cc_93 B1 N_A_27_297#_c_175_n 0.0537361f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_94 N_B1_c_104_n N_VPWR_c_186_n 0.001145f $X=1.535 $Y=1.41 $X2=0 $Y2=0
cc_95 N_B1_c_104_n N_VPWR_c_188_n 0.00515942f $X=1.535 $Y=1.41 $X2=0 $Y2=0
cc_96 B1 N_VPWR_c_188_n 0.0172433f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_97 N_B1_c_104_n N_VPWR_c_185_n 0.00844384f $X=1.535 $Y=1.41 $X2=0 $Y2=0
cc_98 B1 N_VPWR_c_185_n 0.0106598f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_99 B1 A_325_297# 0.0103747f $X=1.625 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_100 N_B1_c_103_n N_Y_c_222_n 0.00419984f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_101 N_B1_c_103_n N_Y_c_229_n 0.0134907f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_102 N_B1_c_104_n N_Y_c_229_n 8.12006e-19 $X=1.535 $Y=1.41 $X2=0 $Y2=0
cc_103 B1 N_Y_c_229_n 0.0203048f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_104 B1 Y 0.0048114f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_105 N_B1_c_104_n N_Y_c_221_n 6.2616e-19 $X=1.535 $Y=1.41 $X2=0 $Y2=0
cc_106 B1 N_Y_c_221_n 0.0546307f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_107 N_B1_c_103_n N_VGND_c_263_n 0.00324768f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_108 N_B1_c_103_n N_VGND_c_265_n 0.00412062f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_109 N_B1_c_103_n N_VGND_c_266_n 0.00849822f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_110 N_C1_c_140_n N_VPWR_c_188_n 0.00469527f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_111 N_C1_c_140_n N_VPWR_c_185_n 0.00822901f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_112 C1 N_Y_M1001_d 0.00236994f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_113 N_C1_c_139_n N_Y_c_229_n 0.0166356f $X=2.005 $Y=0.995 $X2=0 $Y2=0
cc_114 N_C1_c_140_n N_Y_c_229_n 0.00115372f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_115 C1 N_Y_c_229_n 0.0189773f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_116 N_C1_c_139_n N_Y_c_239_n 0.00996699f $X=2.005 $Y=0.995 $X2=0 $Y2=0
cc_117 N_C1_c_139_n Y 0.00519106f $X=2.005 $Y=0.995 $X2=0 $Y2=0
cc_118 N_C1_c_140_n Y 0.0124586f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_119 C1 Y 0.0477265f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_120 N_C1_c_140_n N_Y_c_221_n 0.0331006f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_121 C1 N_Y_c_221_n 0.019359f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_122 N_C1_c_139_n N_VGND_c_264_n 0.0042361f $X=2.005 $Y=0.995 $X2=0 $Y2=0
cc_123 N_C1_c_139_n N_VGND_c_265_n 0.00693655f $X=2.005 $Y=0.995 $X2=0 $Y2=0
cc_124 N_C1_c_139_n N_VGND_c_266_n 0.00329965f $X=2.005 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_27_297#_c_166_n N_VPWR_M1000_d 0.00427817f $X=1.145 $Y=1.625
+ $X2=-0.19 $Y2=1.305
cc_126 N_A_27_297#_c_166_n N_VPWR_c_186_n 0.0203436f $X=1.145 $Y=1.625 $X2=0
+ $Y2=0
cc_127 N_A_27_297#_c_164_n N_VPWR_c_187_n 0.0162044f $X=0.28 $Y=1.85 $X2=0 $Y2=0
cc_128 N_A_27_297#_c_175_n N_VPWR_c_188_n 0.0120599f $X=1.24 $Y=1.85 $X2=0 $Y2=0
cc_129 N_A_27_297#_M1000_s N_VPWR_c_185_n 0.00412064f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_130 N_A_27_297#_M1003_d N_VPWR_c_185_n 0.00882399f $X=1.09 $Y=1.485 $X2=0
+ $Y2=0
cc_131 N_A_27_297#_c_164_n N_VPWR_c_185_n 0.00950576f $X=0.28 $Y=1.85 $X2=0
+ $Y2=0
cc_132 N_A_27_297#_c_175_n N_VPWR_c_185_n 0.00700894f $X=1.24 $Y=1.85 $X2=0
+ $Y2=0
cc_133 N_VPWR_c_185_n A_325_297# 0.00760001f $X=2.53 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_134 N_VPWR_c_185_n N_Y_M1001_d 0.00292607f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_135 N_VPWR_c_188_n N_Y_c_221_n 0.0429653f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_136 N_VPWR_c_185_n N_Y_c_221_n 0.025511f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_137 N_Y_c_229_n N_VGND_M1004_d 0.00689988f $X=2.255 $Y=0.72 $X2=0 $Y2=0
cc_138 N_Y_c_222_n N_VGND_c_263_n 0.0119078f $X=1.24 $Y=0.53 $X2=0 $Y2=0
cc_139 N_Y_c_229_n N_VGND_c_263_n 0.00318253f $X=2.255 $Y=0.72 $X2=0 $Y2=0
cc_140 N_Y_c_229_n N_VGND_c_264_n 0.0084571f $X=2.255 $Y=0.72 $X2=0 $Y2=0
cc_141 N_Y_c_239_n N_VGND_c_264_n 0.0140817f $X=2.355 $Y=0.53 $X2=0 $Y2=0
cc_142 N_Y_M1006_d N_VGND_c_265_n 0.00709856f $X=1.05 $Y=0.235 $X2=0 $Y2=0
cc_143 N_Y_M1007_d N_VGND_c_265_n 0.00386049f $X=2.08 $Y=0.235 $X2=0 $Y2=0
cc_144 N_Y_c_222_n N_VGND_c_265_n 0.00697444f $X=1.24 $Y=0.53 $X2=0 $Y2=0
cc_145 N_Y_c_229_n N_VGND_c_265_n 0.0206748f $X=2.255 $Y=0.72 $X2=0 $Y2=0
cc_146 N_Y_c_239_n N_VGND_c_265_n 0.00840761f $X=2.355 $Y=0.53 $X2=0 $Y2=0
cc_147 N_Y_c_222_n N_VGND_c_266_n 0.0121277f $X=1.24 $Y=0.53 $X2=0 $Y2=0
cc_148 N_Y_c_229_n N_VGND_c_266_n 0.020093f $X=2.255 $Y=0.72 $X2=0 $Y2=0
cc_149 N_Y_c_239_n N_VGND_c_266_n 0.00960872f $X=2.355 $Y=0.53 $X2=0 $Y2=0
cc_150 N_VGND_c_265_n A_123_47# 0.00229207f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24
