* File: sky130_fd_sc_hdll__a21boi_4.pex.spice
* Created: Wed Sep  2 08:16:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A21BOI_4%B1_N 1 3 4 6 7
r32 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.535
+ $Y=1.16 $X2=0.535 $Y2=1.16
r33 7 11 8.83366 $w=5.11e-07 $l=3.7e-07 $layer=LI1_cond $X=0.392 $Y=1.53
+ $X2=0.392 $Y2=1.16
r34 4 10 38.5462 $w=3.19e-07 $l=2.09105e-07 $layer=POLY_cond $X=0.675 $Y=0.995
+ $X2=0.575 $Y2=1.16
r35 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.675 $Y=0.995
+ $X2=0.675 $Y2=0.56
r36 1 10 46.8511 $w=3.19e-07 $l=2.85044e-07 $layer=POLY_cond $X=0.5 $Y=1.41
+ $X2=0.575 $Y2=1.16
r37 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_4%A_27_47# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 31 33 37 39 42 44 50 56 57 66
c118 10 0 3.22468e-20 $X=1.55 $Y=1.41
r119 66 67 45.6841 $w=3.64e-07 $l=3.45e-07 $layer=POLY_cond $X=2.645 $Y=1.202
+ $X2=2.99 $Y2=1.202
r120 65 66 17.8764 $w=3.64e-07 $l=1.35e-07 $layer=POLY_cond $X=2.51 $Y=1.202
+ $X2=2.645 $Y2=1.202
r121 62 63 17.8764 $w=3.64e-07 $l=1.35e-07 $layer=POLY_cond $X=2.03 $Y=1.202
+ $X2=2.165 $Y2=1.202
r122 61 62 45.6841 $w=3.64e-07 $l=3.45e-07 $layer=POLY_cond $X=1.685 $Y=1.202
+ $X2=2.03 $Y2=1.202
r123 60 61 17.8764 $w=3.64e-07 $l=1.35e-07 $layer=POLY_cond $X=1.55 $Y=1.202
+ $X2=1.685 $Y2=1.202
r124 51 65 24.4973 $w=3.64e-07 $l=1.85e-07 $layer=POLY_cond $X=2.325 $Y=1.202
+ $X2=2.51 $Y2=1.202
r125 51 63 21.1868 $w=3.64e-07 $l=1.6e-07 $layer=POLY_cond $X=2.325 $Y=1.202
+ $X2=2.165 $Y2=1.202
r126 50 51 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.325
+ $Y=1.16 $X2=2.325 $Y2=1.16
r127 48 60 0.662088 $w=3.64e-07 $l=5e-09 $layer=POLY_cond $X=1.545 $Y=1.202
+ $X2=1.55 $Y2=1.202
r128 48 58 45.022 $w=3.64e-07 $l=3.4e-07 $layer=POLY_cond $X=1.545 $Y=1.202
+ $X2=1.205 $Y2=1.202
r129 47 50 28.997 $w=3.08e-07 $l=7.8e-07 $layer=LI1_cond $X=1.545 $Y=1.19
+ $X2=2.325 $Y2=1.19
r130 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.545
+ $Y=1.16 $X2=1.545 $Y2=1.16
r131 45 57 0.475111 $w=3.1e-07 $l=1.58e-07 $layer=LI1_cond $X=1.155 $Y=1.19
+ $X2=0.997 $Y2=1.19
r132 45 47 14.4985 $w=3.08e-07 $l=3.9e-07 $layer=LI1_cond $X=1.155 $Y=1.19
+ $X2=1.545 $Y2=1.19
r133 43 57 6.30487 $w=2.42e-07 $l=1.87577e-07 $layer=LI1_cond $X=0.925 $Y=1.345
+ $X2=0.997 $Y2=1.19
r134 43 44 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=0.925 $Y=1.345
+ $X2=0.925 $Y2=1.785
r135 42 57 6.30487 $w=2.42e-07 $l=1.55e-07 $layer=LI1_cond $X=0.997 $Y=1.035
+ $X2=0.997 $Y2=1.19
r136 41 42 8.78052 $w=3.13e-07 $l=2.4e-07 $layer=LI1_cond $X=0.997 $Y=0.795
+ $X2=0.997 $Y2=1.035
r137 40 54 5.18785 $w=1.8e-07 $l=1.78e-07 $layer=LI1_cond $X=0.445 $Y=0.705
+ $X2=0.267 $Y2=0.705
r138 39 41 7.49754 $w=1.8e-07 $l=1.96924e-07 $layer=LI1_cond $X=0.84 $Y=0.705
+ $X2=0.997 $Y2=0.795
r139 39 40 24.3384 $w=1.78e-07 $l=3.95e-07 $layer=LI1_cond $X=0.84 $Y=0.705
+ $X2=0.445 $Y2=0.705
r140 38 56 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=1.895
+ $X2=0.26 $Y2=1.895
r141 37 44 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.84 $Y=1.895
+ $X2=0.925 $Y2=1.785
r142 37 38 21.7393 $w=2.18e-07 $l=4.15e-07 $layer=LI1_cond $X=0.84 $Y=1.895
+ $X2=0.425 $Y2=1.895
r143 31 54 2.62307 $w=3.55e-07 $l=9e-08 $layer=LI1_cond $X=0.267 $Y=0.615
+ $X2=0.267 $Y2=0.705
r144 31 33 8.27811 $w=3.53e-07 $l=2.55e-07 $layer=LI1_cond $X=0.267 $Y=0.615
+ $X2=0.267 $Y2=0.36
r145 28 67 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.99 $Y=1.41
+ $X2=2.99 $Y2=1.202
r146 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.99 $Y=1.41
+ $X2=2.99 $Y2=1.985
r147 25 66 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.645 $Y=0.995
+ $X2=2.645 $Y2=1.202
r148 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.645 $Y=0.995
+ $X2=2.645 $Y2=0.56
r149 22 65 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.51 $Y=1.41
+ $X2=2.51 $Y2=1.202
r150 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.51 $Y=1.41
+ $X2=2.51 $Y2=1.985
r151 19 63 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.165 $Y=0.995
+ $X2=2.165 $Y2=1.202
r152 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.165 $Y=0.995
+ $X2=2.165 $Y2=0.56
r153 16 62 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.03 $Y=1.41
+ $X2=2.03 $Y2=1.202
r154 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.03 $Y=1.41
+ $X2=2.03 $Y2=1.985
r155 13 61 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.685 $Y=0.995
+ $X2=1.685 $Y2=1.202
r156 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.685 $Y=0.995
+ $X2=1.685 $Y2=0.56
r157 10 60 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.55 $Y=1.41
+ $X2=1.55 $Y2=1.202
r158 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.55 $Y=1.41
+ $X2=1.55 $Y2=1.985
r159 7 58 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.205 $Y=0.995
+ $X2=1.205 $Y2=1.202
r160 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.205 $Y=0.995
+ $X2=1.205 $Y2=0.56
r161 2 56 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
r162 1 54 182 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.7
r163 1 33 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_4%A2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 27 31 32 33 34 48 51 54
c125 31 0 3.14505e-20 $X=3.695 $Y=1.592
c126 7 0 1.69574e-19 $X=5.875 $Y=0.995
r127 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.905
+ $Y=1.16 $X2=6.905 $Y2=1.16
r128 48 50 3.9187 $w=3.69e-07 $l=3e-08 $layer=POLY_cond $X=6.875 $Y=1.202
+ $X2=6.905 $Y2=1.202
r129 47 48 4.57182 $w=3.69e-07 $l=3.5e-08 $layer=POLY_cond $X=6.84 $Y=1.202
+ $X2=6.875 $Y2=1.202
r130 46 54 6.3601 $w=6.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.515 $Y=1.39
+ $X2=6.18 $Y2=1.39
r131 45 47 42.4526 $w=3.69e-07 $l=3.25e-07 $layer=POLY_cond $X=6.515 $Y=1.202
+ $X2=6.84 $Y2=1.202
r132 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.515
+ $Y=1.16 $X2=6.515 $Y2=1.16
r133 43 45 15.6748 $w=3.69e-07 $l=1.2e-07 $layer=POLY_cond $X=6.395 $Y=1.202
+ $X2=6.515 $Y2=1.202
r134 42 43 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=6.37 $Y=1.202
+ $X2=6.395 $Y2=1.202
r135 41 54 0.0949269 $w=6.28e-07 $l=5e-09 $layer=LI1_cond $X=6.175 $Y=1.39
+ $X2=6.18 $Y2=1.39
r136 40 42 25.4715 $w=3.69e-07 $l=1.95e-07 $layer=POLY_cond $X=6.175 $Y=1.202
+ $X2=6.37 $Y2=1.202
r137 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.175
+ $Y=1.16 $X2=6.175 $Y2=1.16
r138 38 40 35.9214 $w=3.69e-07 $l=2.75e-07 $layer=POLY_cond $X=5.9 $Y=1.202
+ $X2=6.175 $Y2=1.202
r139 37 38 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=5.875 $Y=1.202
+ $X2=5.9 $Y2=1.202
r140 34 51 4.84127 $w=6.28e-07 $l=2.55e-07 $layer=LI1_cond $X=6.65 $Y=1.39
+ $X2=6.905 $Y2=1.39
r141 34 46 2.56303 $w=6.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6.65 $Y=1.39
+ $X2=6.515 $Y2=1.39
r142 32 41 2.56303 $w=6.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6.04 $Y=1.39
+ $X2=6.175 $Y2=1.39
r143 32 33 11.207 $w=6.28e-07 $l=3.15e-07 $layer=LI1_cond $X=6.04 $Y=1.39
+ $X2=5.725 $Y2=1.39
r144 31 33 103.976 $w=2.23e-07 $l=2.03e-06 $layer=LI1_cond $X=3.695 $Y=1.592
+ $X2=5.725 $Y2=1.592
r145 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.465
+ $Y=1.16 $X2=3.465 $Y2=1.16
r146 25 31 7.50513 $w=2.25e-07 $l=2.4775e-07 $layer=LI1_cond $X=3.497 $Y=1.48
+ $X2=3.695 $Y2=1.592
r147 25 27 9.33625 $w=3.93e-07 $l=3.2e-07 $layer=LI1_cond $X=3.497 $Y=1.48
+ $X2=3.497 $Y2=1.16
r148 22 48 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.875 $Y=0.995
+ $X2=6.875 $Y2=1.202
r149 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.875 $Y=0.995
+ $X2=6.875 $Y2=0.56
r150 19 47 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.84 $Y=1.41
+ $X2=6.84 $Y2=1.202
r151 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.84 $Y=1.41
+ $X2=6.84 $Y2=1.985
r152 16 43 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.395 $Y=0.995
+ $X2=6.395 $Y2=1.202
r153 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.395 $Y=0.995
+ $X2=6.395 $Y2=0.56
r154 13 42 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.37 $Y=1.41
+ $X2=6.37 $Y2=1.202
r155 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.37 $Y=1.41
+ $X2=6.37 $Y2=1.985
r156 10 38 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.9 $Y=1.41 $X2=5.9
+ $Y2=1.202
r157 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.9 $Y=1.41
+ $X2=5.9 $Y2=1.985
r158 7 37 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.875 $Y=0.995
+ $X2=5.875 $Y2=1.202
r159 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.875 $Y=0.995
+ $X2=5.875 $Y2=0.56
r160 4 28 38.7084 $w=3.43e-07 $l=1.90526e-07 $layer=POLY_cond $X=3.545 $Y=0.995
+ $X2=3.49 $Y2=1.16
r161 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.545 $Y=0.995
+ $X2=3.545 $Y2=0.56
r162 1 28 45.964 $w=3.43e-07 $l=2.54951e-07 $layer=POLY_cond $X=3.5 $Y=1.41
+ $X2=3.49 $Y2=1.16
r163 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.5 $Y=1.41 $X2=3.5
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_4%A1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 44 45 52
r73 45 46 3.33795 $w=3.61e-07 $l=2.5e-08 $layer=POLY_cond $X=5.43 $Y=1.2
+ $X2=5.455 $Y2=1.2
r74 44 52 21.8729 $w=2.43e-07 $l=4.65e-07 $layer=LI1_cond $X=5.265 $Y=1.187
+ $X2=4.8 $Y2=1.187
r75 43 45 22.0305 $w=3.61e-07 $l=1.65e-07 $layer=POLY_cond $X=5.265 $Y=1.2
+ $X2=5.43 $Y2=1.2
r76 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.265
+ $Y=1.16 $X2=5.265 $Y2=1.16
r77 41 43 41.3906 $w=3.61e-07 $l=3.1e-07 $layer=POLY_cond $X=4.955 $Y=1.2
+ $X2=5.265 $Y2=1.2
r78 40 41 0.66759 $w=3.61e-07 $l=5e-09 $layer=POLY_cond $X=4.95 $Y=1.2 $X2=4.955
+ $Y2=1.2
r79 38 40 10.0139 $w=3.61e-07 $l=7.5e-08 $layer=POLY_cond $X=4.875 $Y=1.2
+ $X2=4.95 $Y2=1.2
r80 38 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.875
+ $Y=1.16 $X2=4.875 $Y2=1.16
r81 35 38 52.072 $w=3.61e-07 $l=3.9e-07 $layer=POLY_cond $X=4.485 $Y=1.2
+ $X2=4.875 $Y2=1.2
r82 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.485
+ $Y=1.16 $X2=4.485 $Y2=1.16
r83 33 35 1.33518 $w=3.61e-07 $l=1e-08 $layer=POLY_cond $X=4.475 $Y=1.2
+ $X2=4.485 $Y2=1.2
r84 32 33 0.66759 $w=3.61e-07 $l=5e-09 $layer=POLY_cond $X=4.47 $Y=1.2 $X2=4.475
+ $Y2=1.2
r85 31 36 18.345 $w=2.43e-07 $l=3.9e-07 $layer=LI1_cond $X=4.095 $Y=1.187
+ $X2=4.485 $Y2=1.187
r86 30 32 50.0693 $w=3.61e-07 $l=3.75e-07 $layer=POLY_cond $X=4.095 $Y=1.2
+ $X2=4.47 $Y2=1.2
r87 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.095
+ $Y=1.16 $X2=4.095 $Y2=1.16
r88 28 30 14.0194 $w=3.61e-07 $l=1.05e-07 $layer=POLY_cond $X=3.99 $Y=1.2
+ $X2=4.095 $Y2=1.2
r89 27 28 3.33795 $w=3.61e-07 $l=2.5e-08 $layer=POLY_cond $X=3.965 $Y=1.2
+ $X2=3.99 $Y2=1.2
r90 25 52 0.235192 $w=2.43e-07 $l=5e-09 $layer=LI1_cond $X=4.795 $Y=1.187
+ $X2=4.8 $Y2=1.187
r91 25 36 14.5819 $w=2.43e-07 $l=3.1e-07 $layer=LI1_cond $X=4.795 $Y=1.187
+ $X2=4.485 $Y2=1.187
r92 22 46 23.3725 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.455 $Y=0.99
+ $X2=5.455 $Y2=1.2
r93 22 24 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.455 $Y=0.99
+ $X2=5.455 $Y2=0.56
r94 19 45 19.0337 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=5.43 $Y=1.41
+ $X2=5.43 $Y2=1.2
r95 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.43 $Y=1.41
+ $X2=5.43 $Y2=1.985
r96 16 41 23.3725 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.955 $Y=0.99
+ $X2=4.955 $Y2=1.2
r97 16 18 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.955 $Y=0.99
+ $X2=4.955 $Y2=0.56
r98 13 40 19.0337 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=4.95 $Y=1.41
+ $X2=4.95 $Y2=1.2
r99 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.95 $Y=1.41
+ $X2=4.95 $Y2=1.985
r100 10 33 23.3725 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.475 $Y=0.99
+ $X2=4.475 $Y2=1.2
r101 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.475 $Y=0.99
+ $X2=4.475 $Y2=0.56
r102 7 32 19.0337 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=4.47 $Y=1.41
+ $X2=4.47 $Y2=1.2
r103 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.47 $Y=1.41
+ $X2=4.47 $Y2=1.985
r104 4 28 19.0337 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=3.99 $Y=1.41
+ $X2=3.99 $Y2=1.2
r105 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.99 $Y=1.41
+ $X2=3.99 $Y2=1.985
r106 1 27 23.3725 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.965 $Y=0.99
+ $X2=3.965 $Y2=1.2
r107 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.965 $Y=0.99
+ $X2=3.965 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_4%VPWR 1 2 3 4 5 20 23 26 30 33 36 48 52 59
+ 60 63 66 73
r115 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r116 73 76 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=6.605 $Y=2.36
+ $X2=6.605 $Y2=2.72
r117 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r118 66 69 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=5.645 $Y=2.36
+ $X2=5.645 $Y2=2.72
r119 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r120 60 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=6.67 $Y2=2.72
r121 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r122 57 76 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.795 $Y=2.72
+ $X2=6.605 $Y2=2.72
r123 57 59 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.795 $Y=2.72
+ $X2=7.13 $Y2=2.72
r124 56 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r125 56 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r126 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r127 53 69 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.835 $Y=2.72
+ $X2=5.645 $Y2=2.72
r128 53 55 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.835 $Y=2.72
+ $X2=6.21 $Y2=2.72
r129 52 76 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.415 $Y=2.72
+ $X2=6.605 $Y2=2.72
r130 52 55 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.415 $Y=2.72
+ $X2=6.21 $Y2=2.72
r131 51 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r132 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r133 48 69 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.455 $Y=2.72
+ $X2=5.645 $Y2=2.72
r134 48 50 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.455 $Y=2.72
+ $X2=5.29 $Y2=2.72
r135 47 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r136 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r137 44 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r138 43 44 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r139 41 44 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r140 41 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r141 40 43 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r142 40 41 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r143 38 63 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.905 $Y=2.72
+ $X2=0.775 $Y2=2.72
r144 38 40 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.905 $Y=2.72
+ $X2=1.15 $Y2=2.72
r145 36 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r146 34 50 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.875 $Y=2.72
+ $X2=5.29 $Y2=2.72
r147 33 46 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.495 $Y=2.72
+ $X2=4.37 $Y2=2.72
r148 32 34 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.685 $Y=2.72
+ $X2=4.875 $Y2=2.72
r149 32 33 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.685 $Y=2.72
+ $X2=4.495 $Y2=2.72
r150 30 32 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=4.685 $Y=2.36
+ $X2=4.685 $Y2=2.72
r151 27 46 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.915 $Y=2.72
+ $X2=4.37 $Y2=2.72
r152 26 43 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=2.72
+ $X2=3.45 $Y2=2.72
r153 25 27 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.725 $Y=2.72
+ $X2=3.915 $Y2=2.72
r154 25 26 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.725 $Y=2.72
+ $X2=3.535 $Y2=2.72
r155 23 25 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.725 $Y=2.36
+ $X2=3.725 $Y2=2.72
r156 18 63 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=2.635
+ $X2=0.775 $Y2=2.72
r157 18 20 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.775 $Y=2.635
+ $X2=0.775 $Y2=2.34
r158 5 73 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=6.46
+ $Y=1.485 $X2=6.605 $Y2=2.36
r159 4 66 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=5.52
+ $Y=1.485 $X2=5.665 $Y2=2.36
r160 3 30 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=4.56
+ $Y=1.485 $X2=4.71 $Y2=2.36
r161 2 23 600 $w=1.7e-07 $l=9.51643e-07 $layer=licon1_PDIFF $count=1 $X=3.59
+ $Y=1.485 $X2=3.75 $Y2=2.36
r162 1 20 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.485 $X2=0.74 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_4%A_227_297# 1 2 3 4 5 6 7 22 24 26 28 29
+ 34 36 40 42 44 46 55 56
c82 29 0 3.22468e-20 $X=3.365 $Y=1.99
r83 51 53 38.9613 $w=3.1e-07 $l=9.9e-07 $layer=LI1_cond $X=2.27 $Y=2.205
+ $X2=3.26 $Y2=2.205
r84 44 58 3.27362 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=7.115 $Y=2.105
+ $X2=7.115 $Y2=1.99
r85 44 46 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=7.115 $Y=2.105
+ $X2=7.115 $Y2=2.3
r86 43 56 4.29433 $w=2.3e-07 $l=9.3e-08 $layer=LI1_cond $X=6.235 $Y=1.99
+ $X2=6.142 $Y2=1.99
r87 42 58 3.55828 $w=2.3e-07 $l=1.25e-07 $layer=LI1_cond $X=6.99 $Y=1.99
+ $X2=7.115 $Y2=1.99
r88 42 43 37.8302 $w=2.28e-07 $l=7.55e-07 $layer=LI1_cond $X=6.99 $Y=1.99
+ $X2=6.235 $Y2=1.99
r89 38 56 2.13709 $w=1.85e-07 $l=1.15e-07 $layer=LI1_cond $X=6.142 $Y=2.105
+ $X2=6.142 $Y2=1.99
r90 38 40 11.6904 $w=1.83e-07 $l=1.95e-07 $layer=LI1_cond $X=6.142 $Y=2.105
+ $X2=6.142 $Y2=2.3
r91 37 55 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=5.285 $Y=1.99
+ $X2=5.19 $Y2=1.99
r92 36 56 4.29433 $w=2.3e-07 $l=9.2e-08 $layer=LI1_cond $X=6.05 $Y=1.99
+ $X2=6.142 $Y2=1.99
r93 36 37 38.3313 $w=2.28e-07 $l=7.65e-07 $layer=LI1_cond $X=6.05 $Y=1.99
+ $X2=5.285 $Y2=1.99
r94 32 55 2.03875 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=5.19 $Y=2.105
+ $X2=5.19 $Y2=1.99
r95 32 34 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=5.19 $Y=2.105
+ $X2=5.19 $Y2=2.3
r96 29 53 4.97025 $w=3.1e-07 $l=2.62298e-07 $layer=LI1_cond $X=3.365 $Y=1.99
+ $X2=3.26 $Y2=2.205
r97 29 31 43.3419 $w=2.28e-07 $l=8.65e-07 $layer=LI1_cond $X=3.365 $Y=1.99
+ $X2=4.23 $Y2=1.99
r98 28 55 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=5.095 $Y=1.99
+ $X2=5.19 $Y2=1.99
r99 28 31 43.3419 $w=2.28e-07 $l=8.65e-07 $layer=LI1_cond $X=5.095 $Y=1.99
+ $X2=4.23 $Y2=1.99
r100 27 49 3.38121 $w=2.5e-07 $l=1.23e-07 $layer=LI1_cond $X=1.425 $Y=2.34
+ $X2=1.302 $Y2=2.34
r101 26 51 8.95388 $w=3.1e-07 $l=2.74317e-07 $layer=LI1_cond $X=2.055 $Y=2.34
+ $X2=2.27 $Y2=2.205
r102 26 27 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=2.055 $Y=2.34
+ $X2=1.425 $Y2=2.34
r103 22 49 3.43619 $w=2.45e-07 $l=1.25e-07 $layer=LI1_cond $X=1.302 $Y=2.215
+ $X2=1.302 $Y2=2.34
r104 22 24 11.9948 $w=2.43e-07 $l=2.55e-07 $layer=LI1_cond $X=1.302 $Y=2.215
+ $X2=1.302 $Y2=1.96
r105 7 58 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=6.93
+ $Y=1.485 $X2=7.075 $Y2=1.96
r106 7 46 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=6.93
+ $Y=1.485 $X2=7.075 $Y2=2.3
r107 6 40 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.99
+ $Y=1.485 $X2=6.135 $Y2=2.3
r108 5 55 600 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=1 $X=5.04
+ $Y=1.485 $X2=5.19 $Y2=1.96
r109 5 34 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=5.04
+ $Y=1.485 $X2=5.19 $Y2=2.3
r110 4 31 600 $w=1.7e-07 $l=5.7513e-07 $layer=licon1_PDIFF $count=1 $X=4.08
+ $Y=1.485 $X2=4.23 $Y2=1.99
r111 3 53 600 $w=1.7e-07 $l=9.00514e-07 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=1.485 $X2=3.26 $Y2=2.3
r112 2 51 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=2.12
+ $Y=1.485 $X2=2.27 $Y2=2.36
r113 1 49 600 $w=1.7e-07 $l=8.77596e-07 $layer=licon1_PDIFF $count=1 $X=1.135
+ $Y=1.485 $X2=1.265 $Y2=2.3
r114 1 24 600 $w=1.7e-07 $l=5.36074e-07 $layer=licon1_PDIFF $count=1 $X=1.135
+ $Y=1.485 $X2=1.265 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_4%Y 1 2 3 4 5 6 19 23 25 28 31 35 38 43 44
+ 45 46 47 53
c88 44 0 1.09328e-19 $X=2.975 $Y=0.795
c89 35 0 1.69574e-19 $X=5.22 $Y=0.76
c90 31 0 1.51849e-19 $X=3.665 $Y=0.785
r91 50 53 18.8715 $w=4.48e-07 $l=7.1e-07 $layer=LI1_cond $X=1.79 $Y=1.81 $X2=2.5
+ $Y2=1.81
r92 47 56 6.51198 $w=4.48e-07 $l=2.45e-07 $layer=LI1_cond $X=2.505 $Y=1.81
+ $X2=2.75 $Y2=1.81
r93 47 53 0.132898 $w=4.48e-07 $l=5e-09 $layer=LI1_cond $X=2.505 $Y=1.81 $X2=2.5
+ $Y2=1.81
r94 45 56 1.86057 $w=4.48e-07 $l=7e-08 $layer=LI1_cond $X=2.82 $Y=1.81 $X2=2.75
+ $Y2=1.81
r95 33 35 50.2884 $w=2.18e-07 $l=9.6e-07 $layer=LI1_cond $X=4.26 $Y=0.785
+ $X2=5.22 $Y2=0.785
r96 31 46 5.8804 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=3.665 $Y=0.785
+ $X2=3.555 $Y2=0.785
r97 31 33 31.1683 $w=2.18e-07 $l=5.95e-07 $layer=LI1_cond $X=3.665 $Y=0.785
+ $X2=4.26 $Y2=0.785
r98 30 44 7.74863 $w=1.85e-07 $l=1.55e-07 $layer=LI1_cond $X=3.13 $Y=0.795
+ $X2=2.975 $Y2=0.795
r99 30 46 23.5682 $w=1.98e-07 $l=4.25e-07 $layer=LI1_cond $X=3.13 $Y=0.795
+ $X2=3.555 $Y2=0.795
r100 28 45 8.72399 $w=3.1e-07 $l=2.92404e-07 $layer=LI1_cond $X=2.975 $Y=1.585
+ $X2=2.82 $Y2=1.81
r101 27 44 0.431444 $w=3.1e-07 $l=1e-07 $layer=LI1_cond $X=2.975 $Y=0.895
+ $X2=2.975 $Y2=0.795
r102 27 28 25.6511 $w=3.08e-07 $l=6.9e-07 $layer=LI1_cond $X=2.975 $Y=0.895
+ $X2=2.975 $Y2=1.585
r103 26 43 4.74942 $w=2.1e-07 $l=1.13248e-07 $layer=LI1_cond $X=2.525 $Y=0.78
+ $X2=2.43 $Y2=0.74
r104 25 44 7.74863 $w=1.85e-07 $l=1.62327e-07 $layer=LI1_cond $X=2.82 $Y=0.78
+ $X2=2.975 $Y2=0.795
r105 25 26 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.82 $Y=0.78
+ $X2=2.525 $Y2=0.78
r106 21 43 1.70532 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=2.43 $Y=0.615
+ $X2=2.43 $Y2=0.74
r107 21 23 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=2.43 $Y=0.615
+ $X2=2.43 $Y2=0.42
r108 20 38 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=1.47 $Y=0.74
+ $X2=1.47 $Y2=0.535
r109 19 43 4.74942 $w=2.1e-07 $l=9.5e-08 $layer=LI1_cond $X=2.335 $Y=0.74
+ $X2=2.43 $Y2=0.74
r110 19 20 35.4952 $w=2.48e-07 $l=7.7e-07 $layer=LI1_cond $X=2.335 $Y=0.74
+ $X2=1.565 $Y2=0.74
r111 6 56 600 $w=1.7e-07 $l=4.74104e-07 $layer=licon1_PDIFF $count=1 $X=2.6
+ $Y=1.485 $X2=2.75 $Y2=1.89
r112 5 50 600 $w=1.7e-07 $l=4.33561e-07 $layer=licon1_PDIFF $count=1 $X=1.64
+ $Y=1.485 $X2=1.79 $Y2=1.85
r113 4 35 182 $w=1.7e-07 $l=6.12679e-07 $layer=licon1_NDIFF $count=1 $X=5.03
+ $Y=0.235 $X2=5.22 $Y2=0.76
r114 3 33 182 $w=1.7e-07 $l=6.254e-07 $layer=licon1_NDIFF $count=1 $X=4.04
+ $Y=0.235 $X2=4.26 $Y2=0.76
r115 2 43 182 $w=1.7e-07 $l=6.12679e-07 $layer=licon1_NDIFF $count=1 $X=2.24
+ $Y=0.235 $X2=2.43 $Y2=0.76
r116 2 23 182 $w=1.7e-07 $l=2.66927e-07 $layer=licon1_NDIFF $count=1 $X=2.24
+ $Y=0.235 $X2=2.43 $Y2=0.42
r117 1 38 182 $w=1.7e-07 $l=3.83406e-07 $layer=licon1_NDIFF $count=1 $X=1.28
+ $Y=0.235 $X2=1.47 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_4%VGND 1 2 3 4 5 18 20 22 25 32 33 34 40 56
+ 62 70 73 76
c103 32 0 1.51849e-19 $X=6.085 $Y=0
r104 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r105 72 73 8.65265 $w=6.08e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=0.22
+ $X2=3.385 $Y2=0.22
r106 68 72 6.07843 $w=6.08e-07 $l=3.1e-07 $layer=LI1_cond $X=2.99 $Y=0.22
+ $X2=3.3 $Y2=0.22
r107 68 70 11.7899 $w=6.08e-07 $l=2.45e-07 $layer=LI1_cond $X=2.99 $Y=0.22
+ $X2=2.745 $Y2=0.22
r108 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r109 62 65 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=1.975 $Y=0
+ $X2=1.975 $Y2=0.36
r110 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r111 59 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r112 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r113 56 75 3.9202 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=7 $Y=0 $X2=7.18 $Y2=0
r114 56 58 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7 $Y=0 $X2=6.67
+ $Y2=0
r115 55 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.67
+ $Y2=0
r116 54 55 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r117 52 55 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=3.45 $Y=0 $X2=5.75
+ $Y2=0
r118 52 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r119 51 54 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=3.45 $Y=0 $X2=5.75
+ $Y2=0
r120 51 73 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.45 $Y=0 $X2=3.385
+ $Y2=0
r121 51 52 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r122 48 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r123 48 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r124 47 70 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.53 $Y=0
+ $X2=2.745 $Y2=0
r125 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r126 45 62 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.165 $Y=0 $X2=1.975
+ $Y2=0
r127 45 47 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.165 $Y=0
+ $X2=2.53 $Y2=0
r128 43 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r129 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r130 40 62 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.975
+ $Y2=0
r131 40 42 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=1.61 $Y2=0
r132 38 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r133 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r134 34 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r135 32 54 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.085 $Y=0
+ $X2=5.75 $Y2=0
r136 32 33 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.085 $Y=0 $X2=6.18
+ $Y2=0
r137 31 58 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.275 $Y=0
+ $X2=6.67 $Y2=0
r138 31 33 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.275 $Y=0 $X2=6.18
+ $Y2=0
r139 27 42 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.155 $Y=0
+ $X2=1.61 $Y2=0
r140 25 37 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.77 $Y=0 $X2=0.69
+ $Y2=0
r141 25 29 10.7761 $w=3.83e-07 $l=3.6e-07 $layer=LI1_cond $X=0.962 $Y=0
+ $X2=0.962 $Y2=0.36
r142 25 27 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.962 $Y=0
+ $X2=1.155 $Y2=0
r143 20 75 3.15794 $w=2.4e-07 $l=1.11018e-07 $layer=LI1_cond $X=7.12 $Y=0.085
+ $X2=7.18 $Y2=0
r144 20 22 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=7.12 $Y=0.085
+ $X2=7.12 $Y2=0.38
r145 16 33 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.18 $Y=0.085
+ $X2=6.18 $Y2=0
r146 16 18 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=6.18 $Y=0.085
+ $X2=6.18 $Y2=0.4
r147 5 22 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=6.95
+ $Y=0.235 $X2=7.085 $Y2=0.38
r148 4 18 182 $w=1.7e-07 $l=3.01413e-07 $layer=licon1_NDIFF $count=1 $X=5.95
+ $Y=0.235 $X2=6.18 $Y2=0.4
r149 3 72 91 $w=1.7e-07 $l=6.39453e-07 $layer=licon1_NDIFF $count=2 $X=2.72
+ $Y=0.235 $X2=3.3 $Y2=0.36
r150 2 65 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=1.76
+ $Y=0.235 $X2=1.95 $Y2=0.36
r151 1 29 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=0.75
+ $Y=0.235 $X2=0.95 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_4%A_724_47# 1 2 3 4 13 19 20 21 22 25
r50 23 25 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=6.635 $Y=0.735
+ $X2=6.635 $Y2=0.395
r51 21 23 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=6.445 $Y=0.82
+ $X2=6.635 $Y2=0.735
r52 21 22 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=6.445 $Y=0.82
+ $X2=5.865 $Y2=0.82
r53 20 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.735 $Y=0.735
+ $X2=5.865 $Y2=0.82
r54 19 28 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=5.735 $Y=0.505
+ $X2=5.735 $Y2=0.38
r55 19 20 10.1947 $w=2.58e-07 $l=2.3e-07 $layer=LI1_cond $X=5.735 $Y=0.505
+ $X2=5.735 $Y2=0.735
r56 15 18 45.4063 $w=2.48e-07 $l=9.85e-07 $layer=LI1_cond $X=3.755 $Y=0.38
+ $X2=4.74 $Y2=0.38
r57 13 28 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=5.605 $Y=0.38
+ $X2=5.735 $Y2=0.38
r58 13 18 39.8745 $w=2.48e-07 $l=8.65e-07 $layer=LI1_cond $X=5.605 $Y=0.38
+ $X2=4.74 $Y2=0.38
r59 4 25 91 $w=1.7e-07 $l=2.57876e-07 $layer=licon1_NDIFF $count=2 $X=6.47
+ $Y=0.235 $X2=6.66 $Y2=0.395
r60 3 28 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.53
+ $Y=0.235 $X2=5.665 $Y2=0.36
r61 2 18 182 $w=1.7e-07 $l=2.66927e-07 $layer=licon1_NDIFF $count=1 $X=4.55
+ $Y=0.235 $X2=4.74 $Y2=0.42
r62 1 15 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.62
+ $Y=0.235 $X2=3.755 $Y2=0.42
.ends

