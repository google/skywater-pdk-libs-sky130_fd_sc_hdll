# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nand4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.300000 0.725000 3.710000 1.615000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 1.075000 0.825000 1.655000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495000 0.735000 1.760000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 1.075000 1.325000 1.325000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.901500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.155000 1.495000 2.680000 1.665000 ;
        RECT 1.155000 1.665000 1.485000 2.465000 ;
        RECT 2.190000 1.665000 2.680000 2.005000 ;
        RECT 2.190000 2.005000 2.580000 2.465000 ;
        RECT 2.410000 0.255000 3.000000 0.825000 ;
        RECT 2.410000 0.825000 2.680000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.485000 0.425000 0.715000 ;
      RECT 0.085000  0.715000 1.220000 0.905000 ;
      RECT 0.085000  0.905000 0.260000 2.065000 ;
      RECT 0.085000  2.065000 0.425000 2.465000 ;
      RECT 0.645000  0.085000 0.880000 0.545000 ;
      RECT 0.645000  1.835000 0.975000 2.635000 ;
      RECT 1.050000  0.365000 2.240000 0.555000 ;
      RECT 1.050000  0.555000 1.220000 0.715000 ;
      RECT 1.695000  1.835000 2.015000 2.635000 ;
      RECT 1.990000  0.555000 2.240000 1.325000 ;
      RECT 2.750000  2.175000 3.520000 2.635000 ;
      RECT 2.850000  0.995000 3.125000 1.835000 ;
      RECT 2.850000  1.835000 4.055000 2.005000 ;
      RECT 3.190000  0.085000 3.540000 0.545000 ;
      RECT 3.710000  0.255000 4.055000 0.545000 ;
      RECT 3.740000  2.005000 4.055000 2.465000 ;
      RECT 3.885000  0.545000 4.055000 1.835000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4bb_1
END LIBRARY
