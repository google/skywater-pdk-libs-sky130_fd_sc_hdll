# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__dfrtp_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  10.12000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.615000 1.905000 1.665000 ;
        RECT 1.455000 1.665000 1.770000 2.005000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.530500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.150000 0.255000  9.530000 0.735000 ;
        RECT 9.150000 0.735000 10.010000 0.905000 ;
        RECT 9.240000 1.455000 10.010000 1.625000 ;
        RECT 9.240000 1.625000  9.530000 2.465000 ;
        RECT 9.625000 0.905000 10.010000 1.455000 ;
    END
  END Q
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3.995000 0.735000 4.745000 0.780000 ;
        RECT 3.995000 0.780000 7.865000 0.920000 ;
        RECT 3.995000 0.920000 4.745000 0.965000 ;
        RECT 7.575000 0.735000 7.865000 0.780000 ;
        RECT 7.575000 0.920000 7.865000 0.965000 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.090000  0.345000  0.345000 0.635000 ;
      RECT 0.090000  0.635000  0.890000 0.805000 ;
      RECT 0.090000  1.795000  0.890000 1.965000 ;
      RECT 0.090000  1.965000  0.345000 2.465000 ;
      RECT 0.515000  0.085000  0.895000 0.465000 ;
      RECT 0.515000  2.135000  0.895000 2.635000 ;
      RECT 0.660000  0.805000  0.890000 1.795000 ;
      RECT 1.115000  0.345000  1.285000 2.465000 ;
      RECT 1.575000  0.085000  1.905000 0.445000 ;
      RECT 1.770000  2.175000  1.940000 2.635000 ;
      RECT 2.075000  0.305000  2.495000 0.475000 ;
      RECT 2.075000  0.475000  2.245000 1.835000 ;
      RECT 2.075000  1.835000  2.340000 2.005000 ;
      RECT 2.170000  2.005000  2.340000 2.135000 ;
      RECT 2.170000  2.135000  2.420000 2.465000 ;
      RECT 2.425000  0.765000  2.685000 1.385000 ;
      RECT 2.510000  1.575000  3.025000 1.965000 ;
      RECT 2.685000  2.135000  3.365000 2.465000 ;
      RECT 2.695000  0.305000  3.600000 0.475000 ;
      RECT 2.855000  0.765000  3.210000 0.985000 ;
      RECT 2.855000  0.985000  3.025000 1.575000 ;
      RECT 3.195000  1.185000  4.985000 1.355000 ;
      RECT 3.195000  1.355000  3.365000 2.135000 ;
      RECT 3.430000  0.475000  3.600000 1.185000 ;
      RECT 3.535000  1.865000  4.710000 2.035000 ;
      RECT 3.535000  2.035000  3.705000 2.375000 ;
      RECT 3.725000  1.525000  5.325000 1.695000 ;
      RECT 3.805000  0.765000  4.645000 1.015000 ;
      RECT 3.990000  2.205000  4.320000 2.635000 ;
      RECT 4.525000  0.085000  4.855000 0.545000 ;
      RECT 4.540000  2.035000  4.710000 2.375000 ;
      RECT 4.815000  1.005000  4.985000 1.185000 ;
      RECT 5.005000  2.175000  5.425000 2.635000 ;
      RECT 5.065000  0.275000  5.465000 0.445000 ;
      RECT 5.065000  0.445000  5.325000 0.835000 ;
      RECT 5.155000  0.835000  5.325000 1.525000 ;
      RECT 5.155000  1.695000  5.325000 1.835000 ;
      RECT 5.155000  1.835000  5.815000 2.005000 ;
      RECT 5.605000  0.705000  5.775000 1.495000 ;
      RECT 5.605000  1.495000  6.315000 1.655000 ;
      RECT 5.605000  1.655000  6.660000 1.665000 ;
      RECT 5.645000  2.005000  5.815000 2.465000 ;
      RECT 5.735000  0.255000  6.655000 0.535000 ;
      RECT 5.945000  0.705000  6.315000 1.325000 ;
      RECT 6.050000  2.125000  7.005000 2.465000 ;
      RECT 6.145000  1.665000  6.660000 1.955000 ;
      RECT 6.485000  0.535000  6.655000 1.315000 ;
      RECT 6.485000  1.315000  7.055000 1.485000 ;
      RECT 6.825000  0.085000  6.995000 0.525000 ;
      RECT 6.835000  1.485000  7.055000 1.575000 ;
      RECT 6.835000  1.575000  8.270000 1.745000 ;
      RECT 6.835000  1.745000  7.005000 2.125000 ;
      RECT 6.955000  0.695000  7.335000 0.865000 ;
      RECT 6.955000  0.865000  7.225000 1.145000 ;
      RECT 7.165000  0.295000  8.635000 0.465000 ;
      RECT 7.165000  0.465000  7.335000 0.695000 ;
      RECT 7.340000  2.175000  7.590000 2.635000 ;
      RECT 7.505000  0.635000  7.905000 1.405000 ;
      RECT 7.810000  1.915000  8.610000 2.085000 ;
      RECT 7.810000  2.085000  7.980000 2.375000 ;
      RECT 8.160000  2.255000  8.540000 2.635000 ;
      RECT 8.290000  0.465000  8.635000 1.075000 ;
      RECT 8.290000  1.075000  9.335000 1.285000 ;
      RECT 8.290000  1.285000  8.610000 1.295000 ;
      RECT 8.440000  1.295000  8.610000 1.915000 ;
      RECT 8.810000  0.085000  8.980000 0.895000 ;
      RECT 8.810000  1.575000  8.980000 2.635000 ;
      RECT 9.750000  0.085000  9.920000 0.555000 ;
      RECT 9.750000  1.795000  9.920000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.660000  1.105000 0.830000 1.275000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.115000  1.785000 1.285000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.480000  1.105000 2.650000 1.275000 ;
      RECT 2.725000  1.785000 2.895000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.105000  0.765000 4.275000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.465000  0.765000 4.635000 0.935000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.020000  1.105000 6.190000 1.275000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.470000  1.785000 6.640000 1.955000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.635000  0.765000 7.805000 0.935000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
    LAYER met1 ;
      RECT 0.600000 1.075000 0.890000 1.120000 ;
      RECT 0.600000 1.120000 6.250000 1.260000 ;
      RECT 0.600000 1.260000 0.890000 1.305000 ;
      RECT 1.005000 1.755000 1.345000 1.800000 ;
      RECT 1.005000 1.800000 6.700000 1.940000 ;
      RECT 1.005000 1.940000 1.345000 1.985000 ;
      RECT 2.420000 1.075000 2.710000 1.120000 ;
      RECT 2.420000 1.260000 2.710000 1.305000 ;
      RECT 2.665000 1.755000 2.955000 1.800000 ;
      RECT 2.665000 1.940000 2.955000 1.985000 ;
      RECT 5.960000 1.075000 6.250000 1.120000 ;
      RECT 5.960000 1.260000 6.250000 1.305000 ;
      RECT 6.410000 1.755000 6.700000 1.800000 ;
      RECT 6.410000 1.940000 6.700000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dfrtp_2
